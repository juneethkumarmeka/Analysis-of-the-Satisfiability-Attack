module basic_2500_25000_3000_125_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_1780,In_1366);
nor U1 (N_1,In_2476,In_2482);
nand U2 (N_2,In_1777,In_2139);
xnor U3 (N_3,In_6,In_343);
or U4 (N_4,In_1224,In_1052);
nand U5 (N_5,In_1056,In_2444);
xnor U6 (N_6,In_709,In_246);
nand U7 (N_7,In_1707,In_2023);
xor U8 (N_8,In_102,In_809);
or U9 (N_9,In_458,In_2156);
or U10 (N_10,In_2009,In_1611);
xor U11 (N_11,In_1197,In_715);
nor U12 (N_12,In_1772,In_1727);
xnor U13 (N_13,In_266,In_2248);
or U14 (N_14,In_2279,In_2170);
and U15 (N_15,In_1220,In_31);
nand U16 (N_16,In_321,In_2358);
or U17 (N_17,In_2126,In_2343);
xnor U18 (N_18,In_678,In_72);
nand U19 (N_19,In_1495,In_1553);
or U20 (N_20,In_1905,In_2127);
and U21 (N_21,In_1344,In_1942);
and U22 (N_22,In_846,In_479);
or U23 (N_23,In_1983,In_543);
nor U24 (N_24,In_535,In_508);
nor U25 (N_25,In_1512,In_29);
xnor U26 (N_26,In_931,In_837);
nand U27 (N_27,In_2218,In_1926);
xor U28 (N_28,In_2108,In_2056);
xor U29 (N_29,In_728,In_316);
nor U30 (N_30,In_2202,In_1944);
and U31 (N_31,In_1746,In_1524);
xnor U32 (N_32,In_1639,In_432);
nor U33 (N_33,In_672,In_1744);
and U34 (N_34,In_580,In_1878);
or U35 (N_35,In_869,In_779);
nand U36 (N_36,In_2407,In_326);
and U37 (N_37,In_1219,In_664);
and U38 (N_38,In_1827,In_1102);
nand U39 (N_39,In_104,In_905);
and U40 (N_40,In_2008,In_1800);
xor U41 (N_41,In_1462,In_330);
nor U42 (N_42,In_844,In_2376);
nor U43 (N_43,In_1418,In_2001);
xor U44 (N_44,In_288,In_1149);
xor U45 (N_45,In_514,In_1889);
xnor U46 (N_46,In_2445,In_465);
nand U47 (N_47,In_2200,In_530);
xor U48 (N_48,In_2016,In_47);
nand U49 (N_49,In_82,In_1069);
xor U50 (N_50,In_1797,In_2256);
nor U51 (N_51,In_2437,In_35);
and U52 (N_52,In_2125,In_973);
nor U53 (N_53,In_2349,In_793);
and U54 (N_54,In_1864,In_2154);
xnor U55 (N_55,In_413,In_1377);
or U56 (N_56,In_1533,In_1216);
and U57 (N_57,In_1323,In_2346);
nor U58 (N_58,In_1372,In_2371);
and U59 (N_59,In_303,In_1924);
nor U60 (N_60,In_34,In_441);
or U61 (N_61,In_1764,In_1218);
or U62 (N_62,In_2182,In_1615);
and U63 (N_63,In_200,In_52);
nand U64 (N_64,In_2081,In_1696);
and U65 (N_65,In_696,In_1534);
nor U66 (N_66,In_798,In_1013);
and U67 (N_67,In_981,In_740);
xnor U68 (N_68,In_1730,In_1790);
nor U69 (N_69,In_477,In_1552);
xor U70 (N_70,In_311,In_1045);
or U71 (N_71,In_1527,In_2423);
or U72 (N_72,In_355,In_1342);
xnor U73 (N_73,In_1661,In_1572);
and U74 (N_74,In_1683,In_970);
and U75 (N_75,In_399,In_1310);
nor U76 (N_76,In_1805,In_559);
xnor U77 (N_77,In_1325,In_1291);
and U78 (N_78,In_467,In_1675);
or U79 (N_79,In_1206,In_969);
or U80 (N_80,In_1318,In_2057);
and U81 (N_81,In_989,In_1311);
nor U82 (N_82,In_99,In_1813);
nor U83 (N_83,In_1733,In_1469);
nand U84 (N_84,In_2378,In_2196);
nand U85 (N_85,In_742,In_1968);
xnor U86 (N_86,In_2325,In_175);
xnor U87 (N_87,In_1974,In_1411);
nand U88 (N_88,In_211,In_2152);
nor U89 (N_89,In_1851,In_13);
and U90 (N_90,In_915,In_1460);
nor U91 (N_91,In_1369,In_1811);
and U92 (N_92,In_615,In_1448);
and U93 (N_93,In_1574,In_2354);
and U94 (N_94,In_86,In_207);
and U95 (N_95,In_77,In_1082);
xor U96 (N_96,In_462,In_611);
nor U97 (N_97,In_1681,In_1336);
or U98 (N_98,In_2067,In_1380);
xor U99 (N_99,In_2496,In_357);
nor U100 (N_100,In_692,In_2278);
or U101 (N_101,In_1894,In_1278);
and U102 (N_102,In_481,In_1163);
or U103 (N_103,In_471,In_2122);
nor U104 (N_104,In_2165,In_734);
nand U105 (N_105,In_762,In_2168);
and U106 (N_106,In_1374,In_2043);
xnor U107 (N_107,In_1061,In_2400);
xor U108 (N_108,In_1303,In_1221);
nor U109 (N_109,In_1128,In_493);
nor U110 (N_110,In_993,In_1105);
xor U111 (N_111,In_89,In_1641);
and U112 (N_112,In_939,In_1637);
and U113 (N_113,In_1605,In_95);
or U114 (N_114,In_1845,In_731);
nor U115 (N_115,In_1592,In_2348);
and U116 (N_116,In_2485,In_1545);
or U117 (N_117,In_219,In_1656);
nand U118 (N_118,In_2051,In_1701);
and U119 (N_119,In_588,In_383);
nor U120 (N_120,In_788,In_757);
and U121 (N_121,In_2250,In_1531);
nor U122 (N_122,In_1956,In_1496);
and U123 (N_123,In_901,In_1951);
or U124 (N_124,In_1319,In_187);
and U125 (N_125,In_1277,In_1329);
xnor U126 (N_126,In_547,In_1523);
nand U127 (N_127,In_126,In_2092);
or U128 (N_128,In_2387,In_2073);
nor U129 (N_129,In_784,In_431);
nand U130 (N_130,In_299,In_92);
xnor U131 (N_131,In_1914,In_725);
or U132 (N_132,In_243,In_1255);
xnor U133 (N_133,In_622,In_36);
or U134 (N_134,In_1732,In_2069);
or U135 (N_135,In_1608,In_2306);
xor U136 (N_136,In_230,In_1063);
xnor U137 (N_137,In_1423,In_1565);
nor U138 (N_138,In_1778,In_522);
xor U139 (N_139,In_1171,In_1111);
or U140 (N_140,In_2106,In_2411);
xnor U141 (N_141,In_2300,In_1185);
nand U142 (N_142,In_2041,In_1826);
or U143 (N_143,In_1153,In_277);
nor U144 (N_144,In_1401,In_1486);
or U145 (N_145,In_1022,In_1834);
xnor U146 (N_146,In_928,In_2148);
and U147 (N_147,In_1824,In_1991);
nand U148 (N_148,In_662,In_668);
and U149 (N_149,In_747,In_645);
nand U150 (N_150,In_2266,In_1581);
xor U151 (N_151,In_278,In_2052);
nor U152 (N_152,In_169,In_2227);
nand U153 (N_153,In_65,In_1700);
and U154 (N_154,In_199,In_712);
or U155 (N_155,In_286,In_1433);
or U156 (N_156,In_240,In_2247);
nand U157 (N_157,In_1023,In_867);
xnor U158 (N_158,In_2132,In_1282);
xor U159 (N_159,In_1376,In_1839);
and U160 (N_160,In_2146,In_879);
and U161 (N_161,In_576,In_205);
nand U162 (N_162,In_2426,In_595);
or U163 (N_163,In_2380,In_1576);
and U164 (N_164,In_500,In_2345);
or U165 (N_165,In_2374,In_1210);
nand U166 (N_166,In_283,In_242);
nor U167 (N_167,In_2186,In_1745);
xor U168 (N_168,In_1540,In_135);
nor U169 (N_169,In_1396,In_1502);
nand U170 (N_170,In_623,In_1000);
nor U171 (N_171,In_297,In_674);
or U172 (N_172,In_745,In_132);
and U173 (N_173,In_2025,In_1912);
xor U174 (N_174,In_1668,In_2184);
nor U175 (N_175,In_1722,In_587);
xnor U176 (N_176,In_1646,In_2177);
xor U177 (N_177,In_1341,In_930);
nand U178 (N_178,In_1961,In_875);
and U179 (N_179,In_2157,In_1492);
and U180 (N_180,In_332,In_1934);
xnor U181 (N_181,In_1254,In_967);
or U182 (N_182,In_1907,In_1823);
and U183 (N_183,In_2006,In_2195);
xor U184 (N_184,In_1434,In_494);
or U185 (N_185,In_1066,In_1020);
nor U186 (N_186,In_279,In_1194);
nand U187 (N_187,In_393,In_2397);
xnor U188 (N_188,In_2351,In_1556);
and U189 (N_189,In_1750,In_1741);
or U190 (N_190,In_693,In_564);
nor U191 (N_191,In_667,In_1665);
nand U192 (N_192,In_107,In_158);
nand U193 (N_193,In_1697,In_1994);
xnor U194 (N_194,In_2448,In_1966);
nor U195 (N_195,In_1062,In_1886);
nor U196 (N_196,In_2101,In_67);
xor U197 (N_197,In_2240,In_1724);
and U198 (N_198,In_483,In_222);
and U199 (N_199,In_1513,In_215);
nor U200 (N_200,In_600,In_868);
or U201 (N_201,In_1193,In_1978);
nor U202 (N_202,In_637,In_201);
and U203 (N_203,In_1798,In_453);
or U204 (N_204,In_478,In_1383);
nand U205 (N_205,In_765,In_1122);
or U206 (N_206,In_1161,In_2313);
and U207 (N_207,In_1753,In_774);
xnor U208 (N_208,In_314,In_683);
or U209 (N_209,In_1893,In_2347);
xnor U210 (N_210,In_2276,In_872);
and U211 (N_211,In_1833,In_2271);
nand U212 (N_212,N_19,In_743);
or U213 (N_213,In_1782,In_817);
or U214 (N_214,In_220,N_31);
xor U215 (N_215,In_1755,In_659);
nand U216 (N_216,In_835,In_1184);
nand U217 (N_217,In_1234,In_1166);
or U218 (N_218,In_961,In_444);
nor U219 (N_219,In_142,In_801);
nor U220 (N_220,In_1259,In_1387);
nor U221 (N_221,In_1737,In_2026);
or U222 (N_222,In_1347,In_1628);
or U223 (N_223,In_1067,In_2047);
xnor U224 (N_224,In_2307,In_1268);
and U225 (N_225,In_1612,In_2415);
nand U226 (N_226,In_885,In_329);
nor U227 (N_227,In_94,In_166);
xnor U228 (N_228,In_882,In_308);
xor U229 (N_229,In_1580,In_719);
nor U230 (N_230,In_454,In_598);
xor U231 (N_231,N_42,In_2334);
and U232 (N_232,In_2490,In_2438);
nor U233 (N_233,In_2457,In_2329);
or U234 (N_234,In_348,In_50);
nand U235 (N_235,In_233,In_1686);
and U236 (N_236,In_1620,In_408);
xnor U237 (N_237,In_2024,In_620);
or U238 (N_238,In_519,In_515);
or U239 (N_239,In_244,In_1494);
and U240 (N_240,In_1126,In_632);
nand U241 (N_241,In_2396,In_1666);
and U242 (N_242,In_937,In_310);
nor U243 (N_243,In_565,In_1807);
or U244 (N_244,In_379,N_47);
nand U245 (N_245,In_1487,In_60);
and U246 (N_246,In_1053,In_1522);
xnor U247 (N_247,In_1980,N_60);
nor U248 (N_248,In_2275,In_2392);
nand U249 (N_249,In_298,In_2046);
nand U250 (N_250,In_1480,In_579);
xnor U251 (N_251,In_571,In_88);
xnor U252 (N_252,In_1039,In_2213);
xor U253 (N_253,In_862,In_995);
nor U254 (N_254,In_190,In_1840);
xnor U255 (N_255,In_778,N_188);
nand U256 (N_256,In_1058,In_2239);
xor U257 (N_257,In_344,In_979);
or U258 (N_258,In_639,In_1573);
and U259 (N_259,In_628,In_475);
xnor U260 (N_260,In_1627,In_573);
nor U261 (N_261,In_80,N_58);
and U262 (N_262,In_1624,In_2040);
and U263 (N_263,In_934,In_2499);
and U264 (N_264,In_1408,In_1518);
nor U265 (N_265,In_97,In_1470);
nand U266 (N_266,In_572,In_424);
nand U267 (N_267,In_1332,In_2443);
or U268 (N_268,N_176,In_2489);
nor U269 (N_269,In_1759,In_1493);
nand U270 (N_270,N_80,In_2179);
xnor U271 (N_271,In_133,In_2431);
xor U272 (N_272,In_677,In_2124);
and U273 (N_273,In_1871,In_1997);
nor U274 (N_274,In_1678,N_126);
xor U275 (N_275,In_2174,In_1725);
and U276 (N_276,In_886,In_1571);
or U277 (N_277,In_2064,N_29);
and U278 (N_278,N_63,In_1252);
nand U279 (N_279,In_392,In_2446);
or U280 (N_280,In_1442,In_704);
or U281 (N_281,In_2068,In_1676);
nand U282 (N_282,In_1728,In_2188);
nor U283 (N_283,In_1352,In_223);
nand U284 (N_284,In_660,In_1662);
nand U285 (N_285,In_1348,In_1959);
nand U286 (N_286,In_1528,In_657);
or U287 (N_287,In_2361,In_1904);
xnor U288 (N_288,In_1284,In_239);
and U289 (N_289,In_838,In_2285);
nor U290 (N_290,In_1577,In_155);
nor U291 (N_291,In_259,In_372);
nor U292 (N_292,N_108,In_1005);
and U293 (N_293,In_2493,In_485);
and U294 (N_294,In_518,In_305);
nand U295 (N_295,In_1972,In_74);
or U296 (N_296,In_2497,In_1866);
or U297 (N_297,In_952,In_1337);
nand U298 (N_298,In_1139,N_6);
xor U299 (N_299,N_193,In_491);
or U300 (N_300,In_713,In_1240);
nand U301 (N_301,In_1954,In_1316);
and U302 (N_302,N_28,In_643);
and U303 (N_303,In_476,In_1919);
or U304 (N_304,N_167,In_1884);
xor U305 (N_305,In_425,In_1300);
nand U306 (N_306,In_262,In_2100);
xnor U307 (N_307,N_49,In_193);
nand U308 (N_308,In_68,In_143);
or U309 (N_309,In_331,In_2093);
nor U310 (N_310,In_503,In_1660);
or U311 (N_311,In_1140,In_1481);
nand U312 (N_312,In_698,In_1444);
xnor U313 (N_313,In_2416,In_840);
or U314 (N_314,In_1706,In_1621);
nand U315 (N_315,N_197,In_1963);
or U316 (N_316,In_1869,In_1890);
and U317 (N_317,In_957,N_66);
xor U318 (N_318,In_1175,In_1425);
nand U319 (N_319,In_1355,In_352);
and U320 (N_320,In_1152,In_2091);
or U321 (N_321,In_2031,In_2197);
nor U322 (N_322,In_1525,In_975);
or U323 (N_323,In_2447,In_926);
nor U324 (N_324,In_2190,In_1542);
nor U325 (N_325,In_1575,In_90);
and U326 (N_326,In_1603,In_1091);
nor U327 (N_327,In_828,In_359);
nand U328 (N_328,N_161,In_37);
nand U329 (N_329,N_0,In_2301);
and U330 (N_330,In_129,N_180);
and U331 (N_331,In_263,In_1016);
or U332 (N_332,In_1916,In_1693);
nor U333 (N_333,In_2262,In_1041);
and U334 (N_334,In_1087,In_1743);
nor U335 (N_335,In_871,In_1838);
or U336 (N_336,In_2198,In_2153);
xnor U337 (N_337,In_1454,In_1749);
xor U338 (N_338,In_406,In_2037);
and U339 (N_339,N_21,In_1485);
xnor U340 (N_340,In_404,In_1617);
nor U341 (N_341,In_971,In_922);
nor U342 (N_342,In_1735,In_960);
or U343 (N_343,In_218,In_767);
and U344 (N_344,In_2230,In_280);
and U345 (N_345,In_1776,In_629);
nor U346 (N_346,In_1570,In_1768);
and U347 (N_347,In_70,In_1048);
or U348 (N_348,In_1132,In_2012);
nand U349 (N_349,In_857,In_984);
nor U350 (N_350,In_412,In_2074);
xnor U351 (N_351,In_729,In_2035);
xnor U352 (N_352,In_691,In_2370);
xor U353 (N_353,N_104,In_1245);
nand U354 (N_354,In_2096,In_1483);
and U355 (N_355,In_1642,In_106);
nor U356 (N_356,In_1214,In_845);
nand U357 (N_357,In_1602,In_1949);
nor U358 (N_358,In_2163,In_2063);
nand U359 (N_359,In_1995,In_1189);
and U360 (N_360,In_504,In_2113);
nor U361 (N_361,In_986,In_927);
nor U362 (N_362,In_1883,In_541);
and U363 (N_363,In_428,In_217);
nor U364 (N_364,In_1888,In_20);
and U365 (N_365,In_91,In_1964);
or U366 (N_366,In_427,In_1114);
nand U367 (N_367,In_1710,In_603);
nor U368 (N_368,N_111,In_1283);
or U369 (N_369,In_669,In_499);
xnor U370 (N_370,In_407,N_194);
nand U371 (N_371,In_732,In_1816);
xnor U372 (N_372,In_386,In_338);
xnor U373 (N_373,In_1862,In_796);
and U374 (N_374,In_1162,N_128);
and U375 (N_375,In_1097,In_631);
nand U376 (N_376,In_1721,In_1507);
nand U377 (N_377,In_2357,In_1673);
and U378 (N_378,In_1740,In_908);
nor U379 (N_379,In_2280,In_2102);
nor U380 (N_380,In_722,In_2171);
xnor U381 (N_381,In_532,In_1996);
xor U382 (N_382,In_912,In_295);
or U383 (N_383,N_131,In_1929);
xor U384 (N_384,In_1705,In_955);
or U385 (N_385,In_2070,In_1124);
nor U386 (N_386,In_1739,In_1795);
nor U387 (N_387,In_387,In_2462);
or U388 (N_388,In_1850,N_98);
nor U389 (N_389,In_2269,In_1625);
nand U390 (N_390,In_54,In_2481);
xnor U391 (N_391,In_2222,N_101);
nand U392 (N_392,In_1409,In_2097);
xnor U393 (N_393,In_1451,In_2045);
nand U394 (N_394,In_2389,In_415);
nor U395 (N_395,In_1723,In_555);
and U396 (N_396,N_94,In_1208);
nor U397 (N_397,In_258,In_4);
nand U398 (N_398,In_794,In_2495);
nor U399 (N_399,In_1583,In_118);
and U400 (N_400,In_1936,In_1330);
and U401 (N_401,In_932,In_227);
or U402 (N_402,N_266,In_1748);
nor U403 (N_403,In_489,N_383);
xnor U404 (N_404,In_1447,In_735);
nand U405 (N_405,In_2390,In_168);
nand U406 (N_406,N_241,In_1367);
and U407 (N_407,N_115,In_214);
and U408 (N_408,In_897,N_76);
and U409 (N_409,N_173,In_964);
and U410 (N_410,In_791,In_914);
nand U411 (N_411,N_337,In_1110);
nand U412 (N_412,In_516,In_866);
nor U413 (N_413,N_210,In_1123);
nand U414 (N_414,N_370,In_1671);
or U415 (N_415,N_78,In_2302);
nand U416 (N_416,In_172,In_1249);
nor U417 (N_417,In_2429,In_1456);
and U418 (N_418,N_25,In_2027);
nor U419 (N_419,In_1466,In_1364);
nor U420 (N_420,In_1880,In_2032);
xnor U421 (N_421,In_2456,In_1267);
and U422 (N_422,In_1385,In_1360);
and U423 (N_423,In_1455,N_187);
nor U424 (N_424,In_1351,In_1322);
xnor U425 (N_425,In_2162,In_1923);
or U426 (N_426,In_2014,In_1510);
nor U427 (N_427,In_2083,In_2164);
or U428 (N_428,N_85,In_1276);
and U429 (N_429,In_1560,In_2055);
nor U430 (N_430,In_1940,In_1475);
xnor U431 (N_431,In_1664,In_1498);
nand U432 (N_432,In_10,In_906);
and U433 (N_433,In_397,In_627);
and U434 (N_434,In_2394,In_1808);
nor U435 (N_435,In_1416,In_2455);
nor U436 (N_436,N_335,In_839);
or U437 (N_437,In_1815,N_119);
nor U438 (N_438,In_388,In_766);
and U439 (N_439,In_847,In_2341);
and U440 (N_440,In_1847,In_71);
xor U441 (N_441,In_1855,In_2463);
nor U442 (N_442,In_650,In_703);
xor U443 (N_443,In_1298,In_354);
and U444 (N_444,In_695,N_152);
nor U445 (N_445,In_2422,In_1196);
nor U446 (N_446,In_2298,In_1155);
or U447 (N_447,In_673,In_1537);
xor U448 (N_448,N_40,N_309);
xnor U449 (N_449,N_186,In_333);
or U450 (N_450,In_755,N_62);
nor U451 (N_451,In_1312,In_16);
nor U452 (N_452,In_781,In_1130);
nor U453 (N_453,In_1821,In_2315);
nand U454 (N_454,In_1384,In_430);
nand U455 (N_455,In_2142,In_688);
or U456 (N_456,In_599,In_1195);
and U457 (N_457,In_1948,In_1716);
or U458 (N_458,In_1358,In_852);
nor U459 (N_459,N_61,In_1856);
nor U460 (N_460,In_826,In_1939);
nand U461 (N_461,In_1597,In_877);
and U462 (N_462,In_1841,N_247);
nand U463 (N_463,In_1500,In_1947);
and U464 (N_464,In_583,N_374);
or U465 (N_465,In_340,In_1731);
nor U466 (N_466,In_1065,N_292);
xnor U467 (N_467,In_62,In_1587);
xnor U468 (N_468,In_2464,In_1412);
xor U469 (N_469,In_221,In_276);
nor U470 (N_470,In_1654,In_1586);
nand U471 (N_471,In_1897,In_2194);
nand U472 (N_472,N_319,In_1457);
or U473 (N_473,In_1848,In_1173);
and U474 (N_474,In_120,In_473);
nor U475 (N_475,N_148,N_116);
xor U476 (N_476,N_226,N_325);
or U477 (N_477,In_1302,In_1179);
nand U478 (N_478,In_1227,In_2238);
and U479 (N_479,In_2060,In_1539);
and U480 (N_480,N_264,In_2473);
and U481 (N_481,In_800,In_887);
or U482 (N_482,In_684,In_435);
and U483 (N_483,In_505,In_1598);
and U484 (N_484,In_531,In_255);
xor U485 (N_485,In_1561,N_350);
and U486 (N_486,In_507,In_2461);
nor U487 (N_487,In_12,In_1692);
and U488 (N_488,In_2449,N_312);
nand U489 (N_489,In_2318,N_99);
or U490 (N_490,In_1037,In_96);
and U491 (N_491,In_117,In_968);
nor U492 (N_492,In_245,In_1085);
or U493 (N_493,In_1340,In_946);
and U494 (N_494,In_1299,In_2044);
and U495 (N_495,N_196,In_2309);
or U496 (N_496,N_300,In_2183);
or U497 (N_497,In_1882,In_289);
nor U498 (N_498,In_1075,In_1429);
nand U499 (N_499,N_284,N_362);
nor U500 (N_500,In_966,N_228);
and U501 (N_501,In_284,N_240);
nand U502 (N_502,In_2362,In_25);
or U503 (N_503,In_93,In_312);
nor U504 (N_504,In_1747,In_1096);
nor U505 (N_505,In_281,In_759);
nor U506 (N_506,In_456,N_288);
xor U507 (N_507,In_501,In_2252);
nor U508 (N_508,In_551,In_112);
and U509 (N_509,In_192,In_194);
or U510 (N_510,In_893,In_985);
and U511 (N_511,In_982,In_815);
and U512 (N_512,N_347,In_1168);
and U513 (N_513,In_271,In_250);
or U514 (N_514,In_1382,In_2166);
nor U515 (N_515,In_1021,In_438);
or U516 (N_516,In_1178,In_378);
xor U517 (N_517,In_2377,In_1078);
nand U518 (N_518,In_1094,N_324);
nor U519 (N_519,N_75,In_1160);
and U520 (N_520,In_1089,In_2468);
nor U521 (N_521,N_380,In_450);
nand U522 (N_522,In_2226,N_181);
xnor U523 (N_523,In_417,In_394);
or U524 (N_524,In_2319,In_497);
nand U525 (N_525,In_1177,N_382);
nand U526 (N_526,In_63,In_381);
or U527 (N_527,In_26,In_33);
nor U528 (N_528,In_2135,In_1958);
nor U529 (N_529,In_2365,In_337);
or U530 (N_530,N_209,N_340);
or U531 (N_531,In_2465,In_1354);
and U532 (N_532,In_2283,In_1950);
nand U533 (N_533,In_2007,In_274);
xnor U534 (N_534,In_1713,In_1986);
or U535 (N_535,In_410,In_1314);
nand U536 (N_536,In_1915,In_983);
nor U537 (N_537,N_107,In_2338);
nor U538 (N_538,In_550,In_2267);
and U539 (N_539,In_1109,In_1215);
xor U540 (N_540,N_139,In_1594);
nor U541 (N_541,In_1047,In_1018);
xor U542 (N_542,In_2058,In_2114);
xor U543 (N_543,N_330,In_40);
xnor U544 (N_544,In_53,In_938);
nor U545 (N_545,In_290,In_2062);
xor U546 (N_546,In_2369,N_136);
and U547 (N_547,In_157,In_849);
nand U548 (N_548,In_1346,In_2129);
or U549 (N_549,In_1775,N_171);
nor U550 (N_550,N_93,N_110);
or U551 (N_551,In_1092,In_761);
and U552 (N_552,In_272,In_708);
xnor U553 (N_553,In_2020,In_2199);
nand U554 (N_554,In_1898,In_2216);
or U555 (N_555,In_2088,In_1802);
nor U556 (N_556,In_249,In_2150);
or U557 (N_557,N_331,In_1911);
nand U558 (N_558,In_1590,In_1280);
and U559 (N_559,In_923,In_1402);
and U560 (N_560,In_1622,In_726);
and U561 (N_561,In_681,N_253);
xnor U562 (N_562,In_1719,In_1829);
xnor U563 (N_563,In_1010,In_1394);
nand U564 (N_564,In_1685,N_358);
xor U565 (N_565,In_2308,In_655);
nand U566 (N_566,N_367,In_1362);
xnor U567 (N_567,In_942,N_44);
xor U568 (N_568,In_889,In_2224);
and U569 (N_569,In_14,In_805);
and U570 (N_570,In_619,In_342);
nand U571 (N_571,In_851,In_334);
nand U572 (N_572,N_211,N_314);
xor U573 (N_573,N_163,N_150);
nor U574 (N_574,In_618,In_2160);
xor U575 (N_575,In_216,In_293);
xor U576 (N_576,N_304,In_2478);
nand U577 (N_577,In_2085,In_8);
nand U578 (N_578,In_1117,In_2412);
and U579 (N_579,In_1293,N_221);
or U580 (N_580,In_109,In_749);
or U581 (N_581,N_384,In_2381);
nor U582 (N_582,In_721,N_237);
nor U583 (N_583,In_209,In_495);
or U584 (N_584,In_1718,In_468);
nor U585 (N_585,In_1024,In_2207);
nand U586 (N_586,In_122,In_1115);
xor U587 (N_587,N_316,In_940);
xor U588 (N_588,N_183,In_2115);
or U589 (N_589,N_333,In_1555);
nand U590 (N_590,In_604,In_1489);
xnor U591 (N_591,In_1116,In_482);
nor U592 (N_592,In_2454,N_271);
or U593 (N_593,In_705,In_752);
and U594 (N_594,In_2355,N_151);
nor U595 (N_595,In_1640,In_1957);
xnor U596 (N_596,In_229,In_823);
xnor U597 (N_597,In_870,In_1651);
nand U598 (N_598,In_569,In_2178);
and U599 (N_599,In_1859,N_122);
nor U600 (N_600,In_635,N_160);
nor U601 (N_601,In_1960,In_2273);
xor U602 (N_602,N_385,In_1752);
nand U603 (N_603,In_2428,In_1814);
nand U604 (N_604,In_773,N_411);
nand U605 (N_605,In_1012,In_451);
or U606 (N_606,N_399,In_1273);
nor U607 (N_607,In_900,In_1499);
nand U608 (N_608,N_256,N_120);
nor U609 (N_609,In_162,In_977);
and U610 (N_610,In_1181,N_109);
or U611 (N_611,In_2292,In_2488);
nand U612 (N_612,In_361,In_224);
xnor U613 (N_613,In_402,In_540);
nand U614 (N_614,In_591,In_1538);
xor U615 (N_615,In_212,In_119);
xnor U616 (N_616,N_218,In_607);
xor U617 (N_617,In_1709,In_17);
and U618 (N_618,In_1464,N_364);
or U619 (N_619,N_418,In_506);
nand U620 (N_620,In_916,In_699);
nor U621 (N_621,In_405,N_334);
and U622 (N_622,N_82,N_43);
and U623 (N_623,In_1857,In_830);
or U624 (N_624,In_234,In_1324);
nor U625 (N_625,In_1262,In_1095);
nand U626 (N_626,In_1192,In_795);
or U627 (N_627,In_694,In_1445);
nor U628 (N_628,N_212,In_1150);
xor U629 (N_629,In_1432,In_130);
xnor U630 (N_630,N_528,In_1801);
or U631 (N_631,N_145,In_1688);
and U632 (N_632,N_165,N_287);
and U633 (N_633,In_1453,In_1903);
or U634 (N_634,In_2137,In_1854);
xor U635 (N_635,In_509,In_1271);
or U636 (N_636,In_527,In_524);
nor U637 (N_637,In_1120,In_2367);
or U638 (N_638,In_1708,In_1672);
and U639 (N_639,In_1222,N_321);
and U640 (N_640,In_275,In_461);
nor U641 (N_641,In_1137,In_2466);
or U642 (N_642,In_2452,In_1424);
xnor U643 (N_643,In_2326,In_1151);
nand U644 (N_644,N_232,In_1684);
and U645 (N_645,In_785,In_1029);
or U646 (N_646,N_515,In_1769);
nand U647 (N_647,In_2241,In_1373);
and U648 (N_648,In_2111,In_2486);
and U649 (N_649,In_1881,In_2260);
and U650 (N_650,In_1506,In_666);
xor U651 (N_651,In_2310,N_426);
and U652 (N_652,In_2352,In_1446);
nand U653 (N_653,In_636,In_1989);
xor U654 (N_654,In_153,In_1532);
nand U655 (N_655,In_842,In_1690);
and U656 (N_656,N_96,N_533);
nor U657 (N_657,N_338,In_1359);
nor U658 (N_658,N_591,In_521);
nor U659 (N_659,In_445,In_1872);
or U660 (N_660,In_1371,In_921);
nor U661 (N_661,In_2382,In_1209);
nand U662 (N_662,N_585,N_302);
or U663 (N_663,In_87,In_701);
nand U664 (N_664,In_28,In_1616);
nor U665 (N_665,In_1313,In_2080);
and U666 (N_666,In_1381,In_1543);
xnor U667 (N_667,N_305,In_315);
nor U668 (N_668,N_468,N_466);
xnor U669 (N_669,In_1632,N_421);
nand U670 (N_670,N_213,In_1763);
and U671 (N_671,In_948,N_354);
nor U672 (N_672,N_249,In_770);
or U673 (N_673,In_1633,In_1548);
nor U674 (N_674,In_2089,In_1762);
and U675 (N_675,N_484,In_1521);
or U676 (N_676,In_533,In_2420);
nor U677 (N_677,In_1970,N_134);
or U678 (N_678,N_582,N_493);
or U679 (N_679,In_429,In_123);
or U680 (N_680,In_414,In_1043);
nor U681 (N_681,In_1853,In_2155);
and U682 (N_682,N_439,In_2483);
and U683 (N_683,In_907,In_204);
nand U684 (N_684,In_2299,In_1530);
xnor U685 (N_685,In_890,In_1909);
and U686 (N_686,In_1001,N_198);
or U687 (N_687,In_1682,In_1042);
nor U688 (N_688,N_548,In_663);
nor U689 (N_689,N_71,N_496);
or U690 (N_690,N_225,N_381);
nor U691 (N_691,N_23,In_1256);
and U692 (N_692,N_149,In_2427);
or U693 (N_693,In_1858,In_1865);
xnor U694 (N_694,In_282,N_344);
and U695 (N_695,In_69,In_1551);
xor U696 (N_696,In_810,In_2128);
or U697 (N_697,In_2399,N_257);
xnor U698 (N_698,In_920,In_1027);
xor U699 (N_699,N_248,In_1172);
nand U700 (N_700,In_546,N_233);
xor U701 (N_701,In_32,In_237);
nand U702 (N_702,In_1084,In_2147);
xor U703 (N_703,In_739,In_2187);
and U704 (N_704,In_1225,In_2344);
or U705 (N_705,N_563,In_860);
nor U706 (N_706,In_1073,N_204);
nor U707 (N_707,In_2236,In_484);
nor U708 (N_708,In_2004,In_1503);
xnor U709 (N_709,In_2245,In_1771);
nand U710 (N_710,In_2140,In_2296);
and U711 (N_711,In_746,In_1406);
and U712 (N_712,In_446,In_807);
xor U713 (N_713,In_974,In_2072);
and U714 (N_714,In_792,In_738);
xor U715 (N_715,In_751,N_377);
or U716 (N_716,N_138,In_1514);
nor U717 (N_717,N_452,In_374);
and U718 (N_718,In_167,In_1080);
nand U719 (N_719,In_1953,In_2253);
nor U720 (N_720,In_1026,N_262);
xnor U721 (N_721,In_1417,N_471);
nor U722 (N_722,N_282,In_1201);
nand U723 (N_723,In_1379,In_1121);
xor U724 (N_724,In_945,In_1930);
and U725 (N_725,In_1789,N_89);
xnor U726 (N_726,In_789,In_1145);
and U727 (N_727,In_1081,In_2005);
xor U728 (N_728,N_164,N_65);
nand U729 (N_729,In_39,N_595);
nor U730 (N_730,N_135,N_14);
nor U731 (N_731,In_128,In_377);
xnor U732 (N_732,N_297,N_580);
xnor U733 (N_733,In_1345,In_1754);
xor U734 (N_734,N_589,In_2249);
or U735 (N_735,N_378,In_652);
nor U736 (N_736,N_419,In_2474);
and U737 (N_737,N_222,In_1088);
xor U738 (N_738,In_1286,In_1962);
and U739 (N_739,N_1,In_578);
or U740 (N_740,N_500,N_425);
or U741 (N_741,In_1007,In_896);
and U742 (N_742,In_3,In_228);
nor U743 (N_743,In_1035,In_137);
xor U744 (N_744,In_818,In_772);
xnor U745 (N_745,In_1712,In_633);
or U746 (N_746,In_1263,In_2270);
and U747 (N_747,In_1773,In_1275);
or U748 (N_748,In_41,In_2393);
and U749 (N_749,In_2327,In_996);
nor U750 (N_750,In_486,In_1226);
nor U751 (N_751,In_459,In_816);
xor U752 (N_752,In_1652,In_75);
or U753 (N_753,In_1562,In_2098);
xor U754 (N_754,In_287,N_558);
xnor U755 (N_755,In_2251,In_888);
and U756 (N_756,In_30,In_48);
nand U757 (N_757,In_2000,In_1334);
and U758 (N_758,N_443,In_2320);
nand U759 (N_759,In_1479,In_1188);
nand U760 (N_760,In_2087,In_1786);
or U761 (N_761,N_523,In_806);
nand U762 (N_762,In_1761,N_159);
xor U763 (N_763,In_1820,In_512);
xnor U764 (N_764,In_1207,N_162);
nand U765 (N_765,In_2366,N_192);
or U766 (N_766,In_241,In_944);
nand U767 (N_767,In_2243,N_77);
and U768 (N_768,In_1051,In_2470);
xor U769 (N_769,In_686,In_2324);
or U770 (N_770,N_285,In_2065);
nor U771 (N_771,In_449,N_268);
nor U772 (N_772,In_1104,In_422);
nor U773 (N_773,In_648,In_717);
nor U774 (N_774,In_1817,In_300);
and U775 (N_775,In_1634,In_1567);
nor U776 (N_776,In_360,In_716);
or U777 (N_777,In_1867,In_291);
or U778 (N_778,In_1248,N_303);
nor U779 (N_779,In_1619,In_1647);
nor U780 (N_780,In_997,In_786);
or U781 (N_781,In_61,In_641);
nor U782 (N_782,In_1241,In_2010);
and U783 (N_783,In_1515,In_1357);
or U784 (N_784,In_1796,In_1900);
nand U785 (N_785,In_1535,N_37);
nand U786 (N_786,In_1736,In_2282);
nor U787 (N_787,In_1331,In_1694);
or U788 (N_788,In_710,In_125);
nand U789 (N_789,In_804,In_720);
nor U790 (N_790,In_972,N_544);
and U791 (N_791,In_1459,In_656);
or U792 (N_792,In_2235,N_91);
or U793 (N_793,In_1321,In_987);
xnor U794 (N_794,In_1529,In_605);
nor U795 (N_795,In_727,In_853);
and U796 (N_796,N_432,N_356);
and U797 (N_797,N_177,In_812);
and U798 (N_798,N_422,N_84);
xor U799 (N_799,N_456,N_575);
or U800 (N_800,In_7,In_1317);
or U801 (N_801,In_273,In_1136);
and U802 (N_802,In_1431,N_600);
and U803 (N_803,In_909,N_322);
or U804 (N_804,In_1032,In_1635);
nand U805 (N_805,In_1250,In_1426);
and U806 (N_806,In_1861,In_1198);
nand U807 (N_807,In_366,In_584);
and U808 (N_808,In_115,In_1653);
xnor U809 (N_809,In_1971,N_414);
and U810 (N_810,In_1019,In_1536);
or U811 (N_811,N_236,In_1014);
xnor U812 (N_812,In_2305,N_487);
and U813 (N_813,In_1505,In_1333);
and U814 (N_814,In_1251,In_2254);
nand U815 (N_815,In_469,In_2233);
nor U816 (N_816,In_2430,In_2321);
nor U817 (N_817,N_751,In_1593);
and U818 (N_818,In_1421,N_619);
nand U819 (N_819,N_51,N_341);
or U820 (N_820,In_730,In_2498);
nand U821 (N_821,In_1465,N_766);
xor U822 (N_822,N_406,N_762);
or U823 (N_823,In_1977,In_910);
nand U824 (N_824,In_1405,In_585);
nor U825 (N_825,N_737,In_24);
nand U826 (N_826,In_373,In_2103);
xnor U827 (N_827,In_1478,In_247);
nor U828 (N_828,In_2232,In_707);
or U829 (N_829,In_294,N_450);
xnor U830 (N_830,In_1474,N_651);
and U831 (N_831,In_1589,In_1301);
nor U832 (N_832,In_1093,In_998);
or U833 (N_833,In_256,In_1610);
xnor U834 (N_834,In_1679,In_1973);
nor U835 (N_835,N_118,In_248);
or U836 (N_836,N_670,In_452);
xnor U837 (N_837,N_258,In_38);
and U838 (N_838,In_1591,N_488);
xnor U839 (N_839,In_1182,N_125);
nand U840 (N_840,In_78,In_790);
and U841 (N_841,In_1015,In_174);
xor U842 (N_842,In_2143,N_254);
nand U843 (N_843,In_1204,N_455);
xnor U844 (N_844,In_750,In_113);
and U845 (N_845,In_186,In_416);
or U846 (N_846,In_1835,In_1596);
or U847 (N_847,In_861,In_827);
or U848 (N_848,N_195,N_799);
nor U849 (N_849,In_1272,In_1397);
nand U850 (N_850,In_950,In_526);
and U851 (N_851,In_1200,In_1326);
or U852 (N_852,In_2435,N_654);
xor U853 (N_853,N_442,In_714);
or U854 (N_854,N_546,In_1667);
nand U855 (N_855,In_2002,In_23);
or U856 (N_856,In_2368,In_1338);
xnor U857 (N_857,N_69,N_332);
nor U858 (N_858,N_780,N_396);
or U859 (N_859,In_2360,In_919);
xor U860 (N_860,In_1046,N_779);
xnor U861 (N_861,N_429,In_1335);
and U862 (N_862,N_361,N_207);
nand U863 (N_863,In_2339,N_200);
xnor U864 (N_864,N_718,N_783);
nor U865 (N_865,N_458,In_197);
nor U866 (N_866,N_642,N_641);
nor U867 (N_867,N_627,N_534);
nand U868 (N_868,In_1167,N_656);
and U869 (N_869,In_2353,In_903);
or U870 (N_870,N_514,N_566);
xor U871 (N_871,In_1484,N_764);
and U872 (N_872,In_1517,In_1670);
and U873 (N_873,N_478,In_1618);
nor U874 (N_874,In_947,In_492);
xor U875 (N_875,In_2337,N_798);
xnor U876 (N_876,In_2405,N_415);
xor U877 (N_877,N_463,In_2484);
or U878 (N_878,In_617,In_1698);
nand U879 (N_879,N_86,In_1669);
xnor U880 (N_880,In_1711,In_114);
nand U881 (N_881,In_1164,In_457);
nor U882 (N_882,N_147,N_614);
nor U883 (N_883,N_721,N_208);
xnor U884 (N_884,In_2049,In_1832);
or U885 (N_885,In_841,In_2268);
nor U886 (N_886,In_2119,N_239);
or U887 (N_887,In_675,In_1558);
nand U888 (N_888,In_1147,N_613);
nand U889 (N_889,In_764,In_1793);
nor U890 (N_890,N_525,In_2215);
or U891 (N_891,In_1025,In_1738);
nand U892 (N_892,N_655,In_164);
nand U893 (N_893,N_497,In_895);
and U894 (N_894,N_26,N_782);
nand U895 (N_895,In_1264,In_2460);
or U896 (N_896,N_535,N_676);
nor U897 (N_897,N_388,N_473);
nand U898 (N_898,In_2017,In_1261);
or U899 (N_899,In_2471,N_573);
nor U900 (N_900,N_39,In_2458);
xnor U901 (N_901,N_773,In_753);
xnor U902 (N_902,N_765,In_391);
and U903 (N_903,In_630,In_2145);
nor U904 (N_904,N_663,In_647);
nor U905 (N_905,In_2109,N_677);
nor U906 (N_906,N_681,N_244);
or U907 (N_907,In_385,In_443);
nand U908 (N_908,In_1601,In_1645);
and U909 (N_909,In_2050,N_311);
nand U910 (N_910,In_554,In_1141);
nor U911 (N_911,In_1265,N_4);
or U912 (N_912,In_58,In_365);
and U913 (N_913,N_662,In_2221);
nand U914 (N_914,In_1887,In_210);
xnor U915 (N_915,In_1674,N_598);
and U916 (N_916,In_833,N_569);
or U917 (N_917,N_142,In_2013);
and U918 (N_918,In_183,In_2304);
xor U919 (N_919,In_1158,N_18);
nor U920 (N_920,N_440,N_592);
nand U921 (N_921,In_322,N_434);
or U922 (N_922,N_579,In_2117);
and U923 (N_923,N_52,N_554);
and U924 (N_924,In_1473,In_1287);
nand U925 (N_925,In_2204,In_1232);
nand U926 (N_926,In_644,In_2261);
or U927 (N_927,N_631,In_1269);
nor U928 (N_928,N_644,In_66);
or U929 (N_929,N_172,In_1050);
nor U930 (N_930,N_754,In_904);
xor U931 (N_931,In_1190,N_602);
or U932 (N_932,In_1629,N_386);
and U933 (N_933,In_336,In_1508);
xor U934 (N_934,N_769,N_658);
xor U935 (N_935,N_540,N_216);
and U936 (N_936,In_11,In_1393);
nand U937 (N_937,N_615,N_720);
xor U938 (N_938,In_2330,In_1578);
and U939 (N_939,In_1774,N_526);
nor U940 (N_940,N_270,In_594);
nand U941 (N_941,N_81,N_608);
or U942 (N_942,N_79,In_423);
and U943 (N_943,In_936,In_894);
xnor U944 (N_944,In_999,In_238);
or U945 (N_945,N_294,N_492);
nor U946 (N_946,In_589,In_1742);
xnor U947 (N_947,In_1952,In_1781);
or U948 (N_948,In_1569,In_2475);
nand U949 (N_949,In_1497,N_276);
nor U950 (N_950,In_2459,N_327);
nand U951 (N_951,In_188,In_57);
nor U952 (N_952,In_46,In_1606);
xor U953 (N_953,In_1320,In_163);
and U954 (N_954,N_121,N_791);
or U955 (N_955,In_1235,N_103);
nor U956 (N_956,N_395,In_1588);
nor U957 (N_957,In_1908,In_384);
or U958 (N_958,N_112,In_1308);
xor U959 (N_959,In_2112,In_2383);
nor U960 (N_960,N_155,N_481);
and U961 (N_961,In_1017,In_152);
xnor U962 (N_962,In_1076,N_482);
xnor U963 (N_963,In_2167,N_508);
nand U964 (N_964,N_570,N_323);
xnor U965 (N_965,In_105,N_273);
nand U966 (N_966,In_1427,In_189);
and U967 (N_967,N_743,N_612);
nand U968 (N_968,In_2419,In_2316);
nor U969 (N_969,In_606,In_1482);
nand U970 (N_970,In_642,In_1246);
and U971 (N_971,In_1984,In_1305);
nand U972 (N_972,In_1842,In_1004);
or U973 (N_973,N_74,In_1990);
or U974 (N_974,In_1242,N_223);
nor U975 (N_975,In_2094,N_472);
nand U976 (N_976,N_410,In_1009);
and U977 (N_977,In_1877,N_738);
and U978 (N_978,In_653,In_363);
nor U979 (N_979,N_467,In_2003);
nand U980 (N_980,In_191,In_2172);
nand U981 (N_981,N_190,In_2287);
nor U982 (N_982,In_1757,In_375);
and U983 (N_983,In_2201,In_2028);
nor U984 (N_984,In_320,N_260);
or U985 (N_985,In_1837,In_1392);
or U986 (N_986,In_1343,N_348);
nor U987 (N_987,N_683,In_1399);
nand U988 (N_988,In_511,N_562);
nand U989 (N_989,In_1304,N_697);
or U990 (N_990,N_506,In_2151);
and U991 (N_991,In_2294,N_565);
xnor U992 (N_992,In_685,N_313);
xor U993 (N_993,In_1306,In_2229);
nor U994 (N_994,In_455,In_2469);
or U995 (N_995,N_140,N_480);
xnor U996 (N_996,N_182,In_783);
or U997 (N_997,In_103,N_345);
nand U998 (N_998,N_694,In_2144);
or U999 (N_999,N_553,N_521);
nand U1000 (N_1000,N_923,N_457);
xnor U1001 (N_1001,N_597,In_2149);
nand U1002 (N_1002,N_951,In_318);
or U1003 (N_1003,N_840,In_121);
nor U1004 (N_1004,In_1386,N_34);
or U1005 (N_1005,N_872,In_235);
nand U1006 (N_1006,N_794,N_664);
xor U1007 (N_1007,In_1142,In_1921);
nand U1008 (N_1008,In_723,In_2274);
and U1009 (N_1009,N_555,In_776);
and U1010 (N_1010,In_880,In_1390);
and U1011 (N_1011,N_760,In_582);
nor U1012 (N_1012,N_483,N_693);
and U1013 (N_1013,In_147,In_803);
nor U1014 (N_1014,N_46,In_376);
and U1015 (N_1015,In_1295,In_949);
or U1016 (N_1016,In_2192,N_174);
xor U1017 (N_1017,In_1799,N_932);
or U1018 (N_1018,In_101,N_242);
nand U1019 (N_1019,N_214,N_464);
xor U1020 (N_1020,N_252,N_574);
nand U1021 (N_1021,In_380,In_590);
and U1022 (N_1022,In_127,In_1638);
xnor U1023 (N_1023,In_2193,N_846);
nor U1024 (N_1024,N_680,N_907);
xnor U1025 (N_1025,In_1825,In_1107);
or U1026 (N_1026,N_369,N_255);
nor U1027 (N_1027,N_301,In_586);
xor U1028 (N_1028,In_2259,In_560);
or U1029 (N_1029,N_637,In_98);
nand U1030 (N_1030,In_1770,In_1439);
xor U1031 (N_1031,In_181,In_2011);
nand U1032 (N_1032,N_184,In_1165);
xor U1033 (N_1033,N_969,In_1028);
nor U1034 (N_1034,N_827,N_417);
or U1035 (N_1035,In_1563,N_360);
nor U1036 (N_1036,In_825,In_1875);
or U1037 (N_1037,In_1410,In_1309);
and U1038 (N_1038,N_775,In_654);
nor U1039 (N_1039,In_1751,In_2131);
xor U1040 (N_1040,N_757,N_869);
and U1041 (N_1041,In_418,In_1547);
and U1042 (N_1042,In_836,In_1233);
xnor U1043 (N_1043,N_156,In_1788);
or U1044 (N_1044,In_2409,N_715);
and U1045 (N_1045,N_624,In_1803);
and U1046 (N_1046,In_858,In_182);
nor U1047 (N_1047,N_157,N_963);
nor U1048 (N_1048,In_1365,N_874);
or U1049 (N_1049,N_408,In_736);
xor U1050 (N_1050,In_859,N_516);
and U1051 (N_1051,In_593,In_542);
xnor U1052 (N_1052,N_661,In_2363);
xor U1053 (N_1053,In_165,N_857);
nor U1054 (N_1054,In_1467,N_632);
or U1055 (N_1055,In_1356,In_202);
nor U1056 (N_1056,In_898,N_960);
or U1057 (N_1057,N_365,In_883);
nand U1058 (N_1058,N_296,In_563);
and U1059 (N_1059,N_88,N_717);
nor U1060 (N_1060,N_9,N_185);
or U1061 (N_1061,In_581,N_286);
or U1062 (N_1062,In_364,In_1285);
or U1063 (N_1063,N_441,N_752);
xnor U1064 (N_1064,In_76,In_1702);
or U1065 (N_1065,N_918,In_398);
xnor U1066 (N_1066,In_116,In_265);
nand U1067 (N_1067,N_700,In_285);
xnor U1068 (N_1068,N_618,N_445);
nand U1069 (N_1069,In_918,N_416);
nor U1070 (N_1070,In_536,N_507);
or U1071 (N_1071,N_407,In_1511);
xnor U1072 (N_1072,In_876,In_976);
nand U1073 (N_1073,In_178,N_931);
xor U1074 (N_1074,In_2169,N_902);
nor U1075 (N_1075,N_56,In_680);
nor U1076 (N_1076,N_27,In_261);
and U1077 (N_1077,N_146,In_951);
or U1078 (N_1078,N_234,In_2219);
or U1079 (N_1079,N_5,In_440);
and U1080 (N_1080,In_1981,N_986);
and U1081 (N_1081,In_1938,In_2413);
or U1082 (N_1082,N_290,In_741);
nor U1083 (N_1083,In_171,N_696);
nand U1084 (N_1084,N_852,In_1658);
and U1085 (N_1085,N_501,N_475);
and U1086 (N_1086,In_502,In_81);
xnor U1087 (N_1087,In_538,N_54);
xor U1088 (N_1088,In_1471,N_2);
xnor U1089 (N_1089,N_943,In_1657);
xor U1090 (N_1090,In_843,In_2018);
nand U1091 (N_1091,N_379,In_1756);
nand U1092 (N_1092,In_902,N_454);
nand U1093 (N_1093,In_1794,In_1238);
nand U1094 (N_1094,N_485,In_208);
and U1095 (N_1095,N_48,N_403);
nand U1096 (N_1096,In_403,N_636);
nor U1097 (N_1097,N_424,N_901);
nand U1098 (N_1098,N_934,In_1034);
nor U1099 (N_1099,In_2434,In_2386);
and U1100 (N_1100,In_1229,In_1239);
nand U1101 (N_1101,In_301,In_1070);
or U1102 (N_1102,N_495,N_293);
nor U1103 (N_1103,N_771,In_646);
xor U1104 (N_1104,N_24,N_803);
and U1105 (N_1105,In_1490,In_1604);
nand U1106 (N_1106,N_908,N_144);
xor U1107 (N_1107,In_1353,In_487);
xnor U1108 (N_1108,N_729,N_527);
nand U1109 (N_1109,N_731,In_758);
or U1110 (N_1110,N_746,In_1804);
and U1111 (N_1111,In_110,N_245);
nand U1112 (N_1112,N_476,In_420);
nand U1113 (N_1113,In_2,In_2048);
and U1114 (N_1114,In_980,N_16);
nor U1115 (N_1115,In_254,N_557);
nor U1116 (N_1116,N_645,In_813);
nand U1117 (N_1117,In_2255,In_1339);
nor U1118 (N_1118,N_166,In_954);
nand U1119 (N_1119,N_275,In_1103);
and U1120 (N_1120,In_389,In_2206);
nand U1121 (N_1121,In_2205,N_948);
xnor U1122 (N_1122,N_50,In_146);
nor U1123 (N_1123,In_43,In_2281);
nor U1124 (N_1124,In_356,N_859);
nand U1125 (N_1125,In_1146,In_1368);
or U1126 (N_1126,In_309,In_748);
nor U1127 (N_1127,In_108,In_2212);
nor U1128 (N_1128,N_537,In_179);
nor U1129 (N_1129,In_2209,N_606);
or U1130 (N_1130,N_837,In_1223);
and U1131 (N_1131,In_544,In_2450);
or U1132 (N_1132,In_1979,In_2104);
nor U1133 (N_1133,In_2342,In_480);
and U1134 (N_1134,N_675,In_819);
nand U1135 (N_1135,N_987,In_433);
or U1136 (N_1136,N_884,N_994);
or U1137 (N_1137,In_676,In_27);
nand U1138 (N_1138,In_1378,In_177);
nor U1139 (N_1139,In_1289,In_1935);
nor U1140 (N_1140,N_572,In_991);
xor U1141 (N_1141,In_362,In_679);
nor U1142 (N_1142,In_382,N_469);
nor U1143 (N_1143,N_905,In_963);
and U1144 (N_1144,N_477,N_959);
and U1145 (N_1145,N_845,In_2176);
nand U1146 (N_1146,N_352,In_2033);
nor U1147 (N_1147,N_730,In_2421);
nand U1148 (N_1148,N_622,N_863);
nor U1149 (N_1149,In_268,N_447);
or U1150 (N_1150,N_938,In_2244);
nand U1151 (N_1151,N_545,N_714);
and U1152 (N_1152,In_831,In_612);
nor U1153 (N_1153,N_684,In_151);
xnor U1154 (N_1154,In_1792,N_531);
nor U1155 (N_1155,In_1557,In_1079);
nor U1156 (N_1156,In_1071,In_510);
or U1157 (N_1157,In_2331,In_953);
xor U1158 (N_1158,N_984,In_1290);
or U1159 (N_1159,In_614,N_950);
and U1160 (N_1160,In_1975,N_511);
nor U1161 (N_1161,N_616,In_1307);
nor U1162 (N_1162,In_42,N_881);
or U1163 (N_1163,In_2208,In_775);
nand U1164 (N_1164,N_502,N_889);
or U1165 (N_1165,N_688,In_1040);
nand U1166 (N_1166,N_267,N_811);
nor U1167 (N_1167,N_643,N_988);
nor U1168 (N_1168,In_1436,N_646);
or U1169 (N_1169,N_530,N_92);
xor U1170 (N_1170,In_1931,In_401);
or U1171 (N_1171,In_45,In_1134);
nand U1172 (N_1172,N_339,In_2375);
nand U1173 (N_1173,N_224,In_1413);
and U1174 (N_1174,N_784,N_583);
and U1175 (N_1175,In_1407,In_1691);
xor U1176 (N_1176,In_79,In_2472);
or U1177 (N_1177,N_13,N_123);
xor U1178 (N_1178,N_979,In_2388);
or U1179 (N_1179,In_347,In_1585);
or U1180 (N_1180,In_1112,In_2417);
and U1181 (N_1181,In_18,N_702);
nand U1182 (N_1182,In_1680,In_159);
and U1183 (N_1183,In_601,N_689);
nand U1184 (N_1184,In_1699,In_1849);
xor U1185 (N_1185,In_1895,N_836);
nand U1186 (N_1186,In_2336,In_2203);
or U1187 (N_1187,In_1943,In_671);
nor U1188 (N_1188,In_411,N_105);
or U1189 (N_1189,In_2116,In_64);
xor U1190 (N_1190,In_649,In_464);
nor U1191 (N_1191,N_617,In_1902);
or U1192 (N_1192,N_529,N_824);
xnor U1193 (N_1193,In_2408,In_956);
nor U1194 (N_1194,In_592,In_1729);
nand U1195 (N_1195,In_661,In_2487);
nand U1196 (N_1196,N_787,In_395);
nand U1197 (N_1197,In_2289,In_2082);
nand U1198 (N_1198,In_1154,N_132);
nand U1199 (N_1199,In_574,In_2123);
nor U1200 (N_1200,In_253,In_1086);
and U1201 (N_1201,In_1247,N_728);
nor U1202 (N_1202,N_590,In_1982);
xor U1203 (N_1203,N_1044,N_220);
and U1204 (N_1204,N_756,N_53);
nor U1205 (N_1205,N_848,N_801);
or U1206 (N_1206,N_1181,N_512);
xnor U1207 (N_1207,In_2418,N_459);
nand U1208 (N_1208,In_609,In_1873);
nor U1209 (N_1209,N_113,In_1274);
and U1210 (N_1210,In_1422,N_668);
or U1211 (N_1211,N_711,N_510);
nand U1212 (N_1212,In_1129,N_790);
or U1213 (N_1213,In_124,In_1819);
or U1214 (N_1214,N_1135,N_289);
nor U1215 (N_1215,In_690,In_1999);
or U1216 (N_1216,In_2015,N_898);
nor U1217 (N_1217,N_1158,In_2030);
or U1218 (N_1218,N_430,N_581);
nor U1219 (N_1219,In_140,N_357);
nor U1220 (N_1220,N_733,In_621);
and U1221 (N_1221,N_542,In_994);
nand U1222 (N_1222,N_911,In_1370);
nand U1223 (N_1223,N_117,In_1055);
and U1224 (N_1224,N_626,In_2373);
and U1225 (N_1225,In_1138,N_315);
nand U1226 (N_1226,N_277,In_2311);
or U1227 (N_1227,In_367,N_318);
nand U1228 (N_1228,In_1477,In_1281);
nand U1229 (N_1229,In_1212,In_863);
nand U1230 (N_1230,N_832,N_623);
and U1231 (N_1231,In_865,In_1437);
nand U1232 (N_1232,In_1985,In_1363);
or U1233 (N_1233,N_559,In_339);
or U1234 (N_1234,N_1192,In_2158);
nand U1235 (N_1235,N_903,N_1050);
and U1236 (N_1236,N_517,In_2272);
or U1237 (N_1237,N_363,N_509);
and U1238 (N_1238,In_1463,In_1440);
nand U1239 (N_1239,In_1113,In_2257);
or U1240 (N_1240,In_1231,In_346);
nand U1241 (N_1241,In_196,In_231);
or U1242 (N_1242,In_1648,N_1095);
or U1243 (N_1243,N_1165,N_759);
nand U1244 (N_1244,In_490,N_470);
or U1245 (N_1245,In_1550,In_924);
xnor U1246 (N_1246,In_1520,N_770);
or U1247 (N_1247,N_133,N_825);
nand U1248 (N_1248,N_561,N_67);
nand U1249 (N_1249,N_826,In_1965);
nand U1250 (N_1250,In_1119,In_2295);
nand U1251 (N_1251,In_2332,In_929);
nand U1252 (N_1252,In_1099,In_1202);
nand U1253 (N_1253,In_1659,N_73);
or U1254 (N_1254,N_230,In_2312);
and U1255 (N_1255,N_1185,N_1051);
xor U1256 (N_1256,N_956,In_1100);
or U1257 (N_1257,In_1415,N_1056);
and U1258 (N_1258,N_763,In_2076);
nand U1259 (N_1259,N_767,In_665);
or U1260 (N_1260,N_1164,N_914);
xor U1261 (N_1261,In_1831,In_306);
xnor U1262 (N_1262,N_1005,In_1791);
nand U1263 (N_1263,N_682,N_1048);
nand U1264 (N_1264,N_143,N_451);
nor U1265 (N_1265,N_701,In_2095);
nand U1266 (N_1266,In_1174,In_173);
xnor U1267 (N_1267,N_604,In_138);
xor U1268 (N_1268,N_1009,N_815);
xor U1269 (N_1269,In_2398,In_1626);
and U1270 (N_1270,N_970,N_1120);
or U1271 (N_1271,N_1163,In_1554);
xnor U1272 (N_1272,In_2340,N_596);
xor U1273 (N_1273,In_537,N_996);
nor U1274 (N_1274,N_1085,N_387);
nor U1275 (N_1275,In_777,N_1151);
nor U1276 (N_1276,N_936,N_778);
and U1277 (N_1277,N_279,In_1720);
and U1278 (N_1278,In_496,In_296);
or U1279 (N_1279,In_1403,In_85);
nor U1280 (N_1280,N_983,N_1182);
or U1281 (N_1281,In_1928,N_274);
nor U1282 (N_1282,N_412,In_2480);
nor U1283 (N_1283,In_602,In_2084);
or U1284 (N_1284,N_427,In_1564);
nand U1285 (N_1285,In_539,N_522);
xor U1286 (N_1286,In_567,N_251);
and U1287 (N_1287,In_1810,N_838);
or U1288 (N_1288,N_710,N_741);
or U1289 (N_1289,In_962,In_313);
xor U1290 (N_1290,N_1003,In_534);
nor U1291 (N_1291,N_547,In_434);
and U1292 (N_1292,In_2054,N_991);
nor U1293 (N_1293,N_892,In_1501);
and U1294 (N_1294,N_796,In_566);
and U1295 (N_1295,In_1244,N_1033);
nand U1296 (N_1296,In_824,N_1076);
or U1297 (N_1297,In_1183,In_2436);
nand U1298 (N_1298,In_1579,N_818);
nand U1299 (N_1299,In_545,In_1987);
nand U1300 (N_1300,In_1230,N_460);
xor U1301 (N_1301,N_448,In_2439);
nor U1302 (N_1302,N_691,In_1036);
or U1303 (N_1303,N_894,N_1114);
nor U1304 (N_1304,In_1398,N_328);
nor U1305 (N_1305,In_832,In_1785);
nand U1306 (N_1306,N_215,In_1933);
xnor U1307 (N_1307,N_625,In_21);
and U1308 (N_1308,N_1038,In_2433);
xnor U1309 (N_1309,In_206,In_2217);
xor U1310 (N_1310,In_2303,In_195);
or U1311 (N_1311,In_2066,N_1117);
or U1312 (N_1312,In_2118,N_1132);
or U1313 (N_1313,N_922,In_706);
nand U1314 (N_1314,In_850,N_945);
xnor U1315 (N_1315,In_570,N_882);
xor U1316 (N_1316,In_1449,In_1191);
nand U1317 (N_1317,In_2328,In_634);
nand U1318 (N_1318,N_394,In_1033);
or U1319 (N_1319,In_1812,N_1052);
nor U1320 (N_1320,N_992,N_409);
or U1321 (N_1321,In_1476,In_1187);
or U1322 (N_1322,In_5,N_611);
nor U1323 (N_1323,In_2293,In_513);
nor U1324 (N_1324,N_897,In_1443);
nor U1325 (N_1325,N_1017,N_1016);
nor U1326 (N_1326,In_2333,In_856);
nor U1327 (N_1327,N_1188,In_270);
nor U1328 (N_1328,In_2029,N_748);
and U1329 (N_1329,In_2286,In_1917);
nor U1330 (N_1330,N_744,In_520);
and U1331 (N_1331,N_833,In_2335);
nand U1332 (N_1332,N_278,In_51);
xor U1333 (N_1333,N_705,In_697);
xnor U1334 (N_1334,N_740,N_706);
xnor U1335 (N_1335,In_83,N_659);
nor U1336 (N_1336,In_978,N_587);
or U1337 (N_1337,In_640,N_667);
nor U1338 (N_1338,N_906,In_577);
xor U1339 (N_1339,N_712,N_758);
nand U1340 (N_1340,N_390,In_2425);
nor U1341 (N_1341,In_760,N_1070);
nor U1342 (N_1342,In_558,N_1079);
nand U1343 (N_1343,In_2036,In_1297);
nor U1344 (N_1344,N_692,In_232);
nor U1345 (N_1345,N_261,In_2364);
xor U1346 (N_1346,N_1014,N_609);
xnor U1347 (N_1347,N_976,N_70);
nor U1348 (N_1348,N_199,In_2277);
nand U1349 (N_1349,N_1144,N_1059);
nand U1350 (N_1350,N_83,N_1035);
and U1351 (N_1351,In_2442,In_2492);
nor U1352 (N_1352,In_1253,N_652);
nand U1353 (N_1353,In_1127,In_409);
or U1354 (N_1354,In_822,N_153);
or U1355 (N_1355,In_1148,In_658);
and U1356 (N_1356,In_1,N_941);
nor U1357 (N_1357,In_2356,N_405);
nand U1358 (N_1358,In_2022,In_2105);
xor U1359 (N_1359,N_935,In_226);
nand U1360 (N_1360,In_1910,In_1031);
nand U1361 (N_1361,N_1139,N_1175);
nor U1362 (N_1362,N_137,N_568);
xor U1363 (N_1363,N_402,In_2265);
xor U1364 (N_1364,N_1110,In_251);
nor U1365 (N_1365,N_1154,N_1145);
nor U1366 (N_1366,N_830,In_687);
xnor U1367 (N_1367,In_608,In_1419);
nor U1368 (N_1368,N_20,In_2385);
nor U1369 (N_1369,N_1065,In_1714);
xor U1370 (N_1370,In_1068,In_176);
xor U1371 (N_1371,In_787,N_834);
and U1372 (N_1372,In_1074,In_1236);
xnor U1373 (N_1373,N_431,In_737);
or U1374 (N_1374,In_1695,In_1844);
nor U1375 (N_1375,N_813,N_974);
nand U1376 (N_1376,N_453,N_939);
and U1377 (N_1377,N_666,In_1003);
or U1378 (N_1378,In_1631,N_87);
nand U1379 (N_1379,N_673,N_971);
nand U1380 (N_1380,N_873,In_769);
and U1381 (N_1381,N_1086,In_1976);
xnor U1382 (N_1382,N_713,In_2133);
or U1383 (N_1383,N_1006,In_225);
and U1384 (N_1384,In_1941,N_839);
or U1385 (N_1385,N_1129,In_1090);
nand U1386 (N_1386,In_2231,N_660);
or U1387 (N_1387,In_756,N_913);
or U1388 (N_1388,In_1064,N_841);
and U1389 (N_1389,In_1967,N_891);
and U1390 (N_1390,In_1993,N_1046);
nand U1391 (N_1391,In_328,N_353);
xor U1392 (N_1392,In_148,In_768);
and U1393 (N_1393,In_2099,In_624);
or U1394 (N_1394,In_1133,In_1260);
or U1395 (N_1395,N_735,N_489);
and U1396 (N_1396,In_319,In_2237);
xor U1397 (N_1397,N_479,In_2322);
or U1398 (N_1398,In_1870,In_2220);
or U1399 (N_1399,In_267,N_203);
nor U1400 (N_1400,N_578,N_808);
and U1401 (N_1401,N_95,N_202);
or U1402 (N_1402,N_1314,N_909);
nor U1403 (N_1403,In_782,N_648);
or U1404 (N_1404,N_867,N_1041);
nand U1405 (N_1405,In_1509,N_806);
or U1406 (N_1406,In_1186,N_449);
nor U1407 (N_1407,N_639,N_686);
or U1408 (N_1408,N_499,N_33);
nor U1409 (N_1409,In_1892,N_628);
nand U1410 (N_1410,In_323,In_2441);
xor U1411 (N_1411,In_1491,In_597);
xor U1412 (N_1412,N_1353,In_1765);
nor U1413 (N_1413,In_2395,N_1028);
or U1414 (N_1414,In_2141,N_462);
xor U1415 (N_1415,In_447,In_488);
nand U1416 (N_1416,In_1644,In_1057);
xor U1417 (N_1417,In_1504,In_2173);
and U1418 (N_1418,N_1209,N_373);
and U1419 (N_1419,N_1385,N_310);
nor U1420 (N_1420,In_1296,N_797);
and U1421 (N_1421,N_1273,N_1354);
or U1422 (N_1422,In_1217,In_1879);
and U1423 (N_1423,N_1111,In_1294);
or U1424 (N_1424,N_634,N_1072);
nor U1425 (N_1425,N_15,N_685);
or U1426 (N_1426,N_1243,N_1219);
nor U1427 (N_1427,N_17,N_870);
and U1428 (N_1428,N_1160,N_1107);
and U1429 (N_1429,In_22,In_1288);
nand U1430 (N_1430,N_102,N_630);
nor U1431 (N_1431,N_896,N_893);
xnor U1432 (N_1432,N_842,In_808);
nor U1433 (N_1433,N_653,N_1069);
nand U1434 (N_1434,N_947,N_1310);
or U1435 (N_1435,In_198,N_1172);
or U1436 (N_1436,N_972,N_154);
nand U1437 (N_1437,In_562,In_529);
nor U1438 (N_1438,N_1390,N_1123);
nand U1439 (N_1439,N_560,N_1251);
or U1440 (N_1440,N_1288,In_913);
xor U1441 (N_1441,N_1242,N_1078);
nand U1442 (N_1442,N_657,In_1054);
nor U1443 (N_1443,In_1784,In_1176);
nor U1444 (N_1444,N_817,N_1352);
or U1445 (N_1445,N_788,In_341);
or U1446 (N_1446,N_1327,In_1863);
xnor U1447 (N_1447,N_36,In_873);
nand U1448 (N_1448,In_1918,N_35);
xnor U1449 (N_1449,In_625,In_568);
and U1450 (N_1450,N_755,N_1091);
nor U1451 (N_1451,N_1349,N_1036);
nand U1452 (N_1452,N_980,In_1143);
and U1453 (N_1453,N_1268,N_205);
nor U1454 (N_1454,In_911,N_342);
nand U1455 (N_1455,N_130,N_1128);
and U1456 (N_1456,N_930,In_2359);
xnor U1457 (N_1457,N_633,In_1349);
and U1458 (N_1458,In_2019,N_1373);
or U1459 (N_1459,N_946,In_1461);
nor U1460 (N_1460,In_2180,In_959);
nor U1461 (N_1461,N_1292,In_1541);
xnor U1462 (N_1462,In_145,In_436);
xnor U1463 (N_1463,N_961,N_1034);
nand U1464 (N_1464,N_1159,N_858);
nor U1465 (N_1465,N_1203,N_789);
nand U1466 (N_1466,N_206,N_929);
nand U1467 (N_1467,N_1319,N_1066);
nor U1468 (N_1468,N_359,N_998);
nand U1469 (N_1469,N_41,In_1677);
xor U1470 (N_1470,N_1092,N_1320);
nor U1471 (N_1471,N_1204,N_1021);
xor U1472 (N_1472,N_854,N_1348);
nor U1473 (N_1473,N_1187,N_1378);
or U1474 (N_1474,N_505,In_811);
and U1475 (N_1475,In_134,N_704);
or U1476 (N_1476,N_949,In_160);
nor U1477 (N_1477,In_396,In_1077);
and U1478 (N_1478,N_1074,In_351);
and U1479 (N_1479,In_878,N_1356);
nor U1480 (N_1480,N_1105,In_1420);
and U1481 (N_1481,In_1846,N_1346);
or U1482 (N_1482,N_599,N_1269);
nand U1483 (N_1483,N_1226,In_421);
or U1484 (N_1484,In_556,N_1272);
nor U1485 (N_1485,In_1809,In_682);
and U1486 (N_1486,N_736,In_1734);
or U1487 (N_1487,In_1704,In_802);
nand U1488 (N_1488,N_1365,In_439);
xnor U1489 (N_1489,In_1549,N_1316);
nand U1490 (N_1490,N_1064,In_1059);
nor U1491 (N_1491,In_1516,In_1932);
nor U1492 (N_1492,N_549,N_1071);
xor U1493 (N_1493,N_1037,In_317);
xor U1494 (N_1494,In_1205,In_1108);
nor U1495 (N_1495,N_1098,N_687);
nor U1496 (N_1496,N_1263,In_470);
nand U1497 (N_1497,N_1282,N_498);
xor U1498 (N_1498,N_1218,In_260);
or U1499 (N_1499,N_1326,N_1257);
and U1500 (N_1500,N_1233,In_1279);
nor U1501 (N_1501,In_2406,N_1029);
and U1502 (N_1502,In_891,N_849);
nor U1503 (N_1503,In_1655,In_2317);
nor U1504 (N_1504,N_219,N_749);
nor U1505 (N_1505,N_1293,N_124);
and U1506 (N_1506,N_1377,N_1077);
and U1507 (N_1507,In_1913,In_100);
or U1508 (N_1508,N_141,N_722);
nand U1509 (N_1509,N_490,N_1255);
or U1510 (N_1510,In_1703,N_665);
and U1511 (N_1511,In_2314,N_265);
nor U1512 (N_1512,In_2191,In_2372);
xnor U1513 (N_1513,N_1113,In_1717);
xor U1514 (N_1514,N_649,In_1636);
and U1515 (N_1515,N_1088,N_1171);
and U1516 (N_1516,N_800,N_610);
xor U1517 (N_1517,N_1053,In_370);
nand U1518 (N_1518,N_1162,N_1388);
nor U1519 (N_1519,In_1375,N_1321);
and U1520 (N_1520,In_744,N_346);
nand U1521 (N_1521,N_993,In_1237);
nand U1522 (N_1522,In_1328,N_1230);
and U1523 (N_1523,N_1323,N_375);
or U1524 (N_1524,N_1104,N_1362);
nor U1525 (N_1525,In_1435,N_1081);
and U1526 (N_1526,N_1278,N_1100);
nand U1527 (N_1527,N_804,N_1109);
xnor U1528 (N_1528,N_320,In_474);
nor U1529 (N_1529,In_1544,In_2288);
nand U1530 (N_1530,N_880,N_1386);
xor U1531 (N_1531,In_2402,In_2214);
or U1532 (N_1532,N_1315,N_263);
xor U1533 (N_1533,N_1026,In_881);
nand U1534 (N_1534,In_1599,N_1130);
xor U1535 (N_1535,N_1178,N_1155);
nand U1536 (N_1536,N_1027,N_1342);
and U1537 (N_1537,N_1068,N_1367);
or U1538 (N_1538,N_64,N_678);
and U1539 (N_1539,N_1061,N_1089);
and U1540 (N_1540,In_463,N_246);
and U1541 (N_1541,N_298,In_988);
and U1542 (N_1542,N_1329,N_1015);
xnor U1543 (N_1543,In_1566,In_2079);
and U1544 (N_1544,In_150,N_1020);
xnor U1545 (N_1545,In_754,N_1283);
or U1546 (N_1546,N_904,N_1240);
nand U1547 (N_1547,N_539,In_1852);
xor U1548 (N_1548,In_2059,N_1191);
and U1549 (N_1549,N_1131,In_149);
and U1550 (N_1550,In_2225,In_1006);
xor U1551 (N_1551,In_2234,In_2189);
or U1552 (N_1552,N_603,N_1004);
xor U1553 (N_1553,N_571,N_888);
or U1554 (N_1554,N_343,N_398);
nand U1555 (N_1555,N_7,In_1101);
nand U1556 (N_1556,In_390,N_1331);
nand U1557 (N_1557,N_1290,In_899);
nand U1558 (N_1558,N_1375,In_1400);
xnor U1559 (N_1559,In_2453,N_1260);
nor U1560 (N_1560,N_486,N_605);
or U1561 (N_1561,In_2297,N_952);
nand U1562 (N_1562,In_2242,N_981);
nor U1563 (N_1563,N_1142,In_1901);
or U1564 (N_1564,N_1058,N_127);
xor U1565 (N_1565,In_1920,In_1584);
or U1566 (N_1566,In_2414,N_1183);
nor U1567 (N_1567,In_1546,In_943);
xor U1568 (N_1568,N_866,N_975);
nand U1569 (N_1569,N_1252,In_1906);
or U1570 (N_1570,N_822,N_1001);
nor U1571 (N_1571,N_1232,N_1166);
or U1572 (N_1572,N_175,N_937);
nor U1573 (N_1573,N_1380,N_169);
or U1574 (N_1574,N_1202,N_1244);
nor U1575 (N_1575,N_1099,N_1221);
and U1576 (N_1576,In_400,In_2185);
nand U1577 (N_1577,In_2086,N_885);
nand U1578 (N_1578,In_2042,N_336);
or U1579 (N_1579,N_1124,In_525);
nand U1580 (N_1580,N_1054,In_2228);
xnor U1581 (N_1581,In_1428,In_184);
or U1582 (N_1582,N_1366,N_1045);
nor U1583 (N_1583,N_404,In_2130);
nor U1584 (N_1584,In_548,N_851);
or U1585 (N_1585,N_1368,In_1072);
nor U1586 (N_1586,In_2290,N_707);
or U1587 (N_1587,N_1190,N_593);
and U1588 (N_1588,In_884,In_1559);
nand U1589 (N_1589,N_985,N_1339);
or U1590 (N_1590,N_1250,In_2021);
and U1591 (N_1591,N_1082,N_1138);
nor U1592 (N_1592,N_444,N_491);
or U1593 (N_1593,In_1472,N_201);
xor U1594 (N_1594,In_1806,N_635);
xnor U1595 (N_1595,N_823,In_610);
nor U1596 (N_1596,In_1649,N_781);
nand U1597 (N_1597,In_84,N_1126);
or U1598 (N_1598,N_543,N_1258);
nor U1599 (N_1599,In_2258,In_141);
or U1600 (N_1600,N_217,N_716);
xor U1601 (N_1601,N_10,In_2210);
xnor U1602 (N_1602,N_724,N_1463);
and U1603 (N_1603,N_179,N_1167);
xor U1604 (N_1604,In_1106,N_920);
and U1605 (N_1605,N_1567,N_921);
nor U1606 (N_1606,N_1141,N_999);
or U1607 (N_1607,N_281,N_1022);
xnor U1608 (N_1608,N_957,N_1442);
and U1609 (N_1609,N_1444,N_1376);
xor U1610 (N_1610,N_1341,In_2159);
and U1611 (N_1611,N_1528,N_1545);
nand U1612 (N_1612,In_2264,N_990);
xor U1613 (N_1613,N_1469,N_1428);
xnor U1614 (N_1614,N_57,N_1309);
or U1615 (N_1615,N_1103,N_1177);
nand U1616 (N_1616,In_368,N_446);
nand U1617 (N_1617,N_392,N_1225);
nand U1618 (N_1618,In_1600,N_954);
or U1619 (N_1619,N_594,N_1451);
nand U1620 (N_1620,N_1197,N_1411);
xor U1621 (N_1621,In_1876,N_955);
xnor U1622 (N_1622,N_1168,N_795);
nand U1623 (N_1623,N_368,N_1464);
nor U1624 (N_1624,N_1345,N_742);
or U1625 (N_1625,N_1208,In_1391);
or U1626 (N_1626,N_1277,In_552);
nor U1627 (N_1627,N_1583,N_168);
or U1628 (N_1628,N_1296,N_944);
and U1629 (N_1629,N_1468,In_711);
xnor U1630 (N_1630,N_928,N_1270);
nand U1631 (N_1631,N_829,N_1170);
nand U1632 (N_1632,In_1726,N_915);
or U1633 (N_1633,N_413,In_820);
nand U1634 (N_1634,N_1482,N_191);
and U1635 (N_1635,N_1237,N_1419);
nand U1636 (N_1636,N_1307,In_2440);
nand U1637 (N_1637,N_1011,In_2451);
nor U1638 (N_1638,In_1389,N_1593);
nand U1639 (N_1639,N_850,N_1577);
nor U1640 (N_1640,N_1460,In_1767);
or U1641 (N_1641,In_517,In_2284);
or U1642 (N_1642,In_170,N_916);
nand U1643 (N_1643,In_1135,N_1304);
xnor U1644 (N_1644,In_161,N_1063);
or U1645 (N_1645,N_1090,N_1222);
or U1646 (N_1646,N_1457,N_1355);
or U1647 (N_1647,In_1899,In_1787);
xnor U1648 (N_1648,In_1868,N_1297);
nand U1649 (N_1649,In_616,N_844);
or U1650 (N_1650,N_820,N_1223);
nand U1651 (N_1651,N_1384,N_1446);
and U1652 (N_1652,In_718,N_819);
or U1653 (N_1653,N_878,In_1203);
or U1654 (N_1654,N_1122,N_1582);
and U1655 (N_1655,In_848,In_252);
nand U1656 (N_1656,N_1420,N_725);
nor U1657 (N_1657,N_428,N_438);
xor U1658 (N_1658,In_1760,N_1289);
nor U1659 (N_1659,N_1449,In_2077);
or U1660 (N_1660,N_1456,N_1499);
xnor U1661 (N_1661,N_32,N_964);
nor U1662 (N_1662,N_1134,N_1106);
xor U1663 (N_1663,N_129,N_1332);
nor U1664 (N_1664,N_1563,N_231);
xnor U1665 (N_1665,In_2379,N_1410);
or U1666 (N_1666,N_805,N_1097);
xor U1667 (N_1667,In_1488,N_1439);
xnor U1668 (N_1668,N_372,N_538);
and U1669 (N_1669,N_1275,N_1118);
and U1670 (N_1670,In_1519,N_1389);
xnor U1671 (N_1671,N_1284,N_11);
xor U1672 (N_1672,N_843,N_861);
nor U1673 (N_1673,In_1388,N_953);
or U1674 (N_1674,N_1264,N_243);
or U1675 (N_1675,N_317,N_1570);
nor U1676 (N_1676,N_695,N_886);
and U1677 (N_1677,N_1302,N_1487);
and U1678 (N_1678,In_2138,N_1083);
nand U1679 (N_1679,In_302,N_940);
nand U1680 (N_1680,N_556,N_1437);
nand U1681 (N_1681,N_1402,In_466);
and U1682 (N_1682,N_1589,N_989);
and U1683 (N_1683,N_1369,N_1517);
nor U1684 (N_1684,N_1459,N_1504);
nor U1685 (N_1685,N_674,N_1347);
nand U1686 (N_1686,In_353,N_1150);
nor U1687 (N_1687,N_1478,In_1891);
nand U1688 (N_1688,N_672,In_180);
nand U1689 (N_1689,In_1243,N_835);
nand U1690 (N_1690,N_461,N_1328);
or U1691 (N_1691,In_2432,In_2071);
nor U1692 (N_1692,N_552,N_1303);
xor U1693 (N_1693,N_1207,N_1513);
or U1694 (N_1694,N_1325,In_2263);
or U1695 (N_1695,N_1093,N_1043);
or U1696 (N_1696,In_19,N_671);
and U1697 (N_1697,N_1581,N_1212);
nor U1698 (N_1698,N_1529,N_1337);
and U1699 (N_1699,N_1568,N_1560);
or U1700 (N_1700,In_596,N_927);
nand U1701 (N_1701,In_1758,N_1245);
nor U1702 (N_1702,N_1075,In_442);
nand U1703 (N_1703,N_1477,N_1440);
and U1704 (N_1704,N_1372,In_56);
and U1705 (N_1705,N_1573,In_1038);
nand U1706 (N_1706,N_1200,In_1144);
nand U1707 (N_1707,N_1102,N_1133);
and U1708 (N_1708,N_640,N_576);
nand U1709 (N_1709,In_702,N_59);
nor U1710 (N_1710,In_821,N_966);
nor U1711 (N_1711,N_1108,N_1569);
or U1712 (N_1712,In_958,N_588);
nand U1713 (N_1713,N_349,N_629);
and U1714 (N_1714,N_1450,In_1458);
or U1715 (N_1715,In_651,N_1174);
xor U1716 (N_1716,N_965,In_1118);
nand U1717 (N_1717,N_860,In_1969);
nor U1718 (N_1718,N_1173,N_1317);
nor U1719 (N_1719,N_1584,In_935);
nand U1720 (N_1720,N_1008,N_1579);
and U1721 (N_1721,In_2410,N_1060);
xnor U1722 (N_1722,N_1350,In_0);
nor U1723 (N_1723,N_1357,N_1519);
nand U1724 (N_1724,N_1476,N_1306);
nor U1725 (N_1725,N_1447,In_1885);
nand U1726 (N_1726,N_1301,N_1580);
xor U1727 (N_1727,N_1497,N_1261);
and U1728 (N_1728,N_810,N_1228);
nor U1729 (N_1729,N_1180,In_1783);
or U1730 (N_1730,N_1246,N_541);
or U1731 (N_1731,N_158,In_2404);
or U1732 (N_1732,In_131,In_523);
and U1733 (N_1733,N_912,In_1258);
or U1734 (N_1734,N_38,N_1518);
or U1735 (N_1735,N_1343,N_1465);
nor U1736 (N_1736,N_1024,In_292);
and U1737 (N_1737,N_1543,N_391);
and U1738 (N_1738,N_1422,In_2467);
nand U1739 (N_1739,In_1595,N_1548);
and U1740 (N_1740,N_435,In_1211);
xor U1741 (N_1741,In_1170,In_2350);
xnor U1742 (N_1742,In_1663,N_1470);
nand U1743 (N_1743,N_3,N_1433);
and U1744 (N_1744,N_1501,N_1473);
nor U1745 (N_1745,N_647,In_613);
nand U1746 (N_1746,In_2161,N_550);
or U1747 (N_1747,In_829,N_1031);
nand U1748 (N_1748,In_2107,In_144);
xor U1749 (N_1749,In_1945,In_448);
or U1750 (N_1750,N_828,N_22);
and U1751 (N_1751,N_1023,N_831);
xnor U1752 (N_1752,N_1351,N_1279);
or U1753 (N_1753,In_1614,N_1259);
xor U1754 (N_1754,N_1299,N_1551);
nand U1755 (N_1755,In_1395,N_1406);
nor U1756 (N_1756,N_389,In_307);
and U1757 (N_1757,In_2391,N_1530);
xnor U1758 (N_1758,N_1340,N_1229);
xnor U1759 (N_1759,N_1364,N_1591);
nor U1760 (N_1760,N_1318,N_917);
xor U1761 (N_1761,N_1550,In_1414);
nor U1762 (N_1762,N_1040,In_2078);
and U1763 (N_1763,In_371,N_1018);
and U1764 (N_1764,N_793,N_532);
nand U1765 (N_1765,In_335,N_366);
nand U1766 (N_1766,In_2223,N_977);
nand U1767 (N_1767,N_1472,N_1042);
or U1768 (N_1768,N_900,In_557);
xnor U1769 (N_1769,N_295,N_812);
and U1770 (N_1770,In_638,N_536);
nand U1771 (N_1771,N_1572,N_1391);
or U1772 (N_1772,In_1650,N_1578);
xor U1773 (N_1773,N_1313,In_1213);
xor U1774 (N_1774,N_8,N_1556);
nor U1775 (N_1775,N_1546,N_1213);
and U1776 (N_1776,N_997,N_1555);
nor U1777 (N_1777,N_1534,N_1596);
nor U1778 (N_1778,In_9,N_178);
xor U1779 (N_1779,N_1067,In_1131);
nand U1780 (N_1780,In_2403,N_1234);
and U1781 (N_1781,N_1336,N_503);
xor U1782 (N_1782,N_1281,In_1836);
nand U1783 (N_1783,N_1407,N_1361);
nand U1784 (N_1784,In_917,In_1468);
nor U1785 (N_1785,N_1479,N_926);
nand U1786 (N_1786,N_807,N_1415);
nand U1787 (N_1787,N_1189,N_1405);
nand U1788 (N_1788,N_1414,N_1112);
xnor U1789 (N_1789,N_1324,N_307);
or U1790 (N_1790,N_1383,N_1503);
nor U1791 (N_1791,N_1535,In_1438);
xnor U1792 (N_1792,In_575,In_561);
nand U1793 (N_1793,In_369,In_1843);
nand U1794 (N_1794,N_1585,N_1539);
nor U1795 (N_1795,N_925,N_229);
xnor U1796 (N_1796,N_1412,In_1687);
nor U1797 (N_1797,N_1480,N_1169);
nand U1798 (N_1798,N_1115,N_1184);
xnor U1799 (N_1799,N_1143,In_2039);
nand U1800 (N_1800,N_1761,N_726);
xnor U1801 (N_1801,N_1619,N_1740);
or U1802 (N_1802,N_1335,N_1678);
and U1803 (N_1803,N_862,N_420);
and U1804 (N_1804,N_1708,In_2494);
and U1805 (N_1805,N_326,In_472);
and U1806 (N_1806,N_1496,N_1489);
xnor U1807 (N_1807,N_1655,N_1484);
xnor U1808 (N_1808,N_1571,N_1540);
nand U1809 (N_1809,In_1643,N_1179);
xor U1810 (N_1810,N_1682,N_669);
xor U1811 (N_1811,N_1693,N_1485);
nand U1812 (N_1812,N_1665,In_139);
nor U1813 (N_1813,N_1757,N_1421);
xor U1814 (N_1814,N_1722,N_1712);
and U1815 (N_1815,N_1711,N_924);
nor U1816 (N_1816,N_1552,N_875);
nor U1817 (N_1817,N_1505,N_1156);
xor U1818 (N_1818,N_761,N_933);
or U1819 (N_1819,N_1656,N_1698);
nor U1820 (N_1820,In_1822,N_1671);
nor U1821 (N_1821,N_1305,N_1586);
and U1822 (N_1822,N_855,N_1597);
nor U1823 (N_1823,N_1012,In_1315);
nand U1824 (N_1824,In_1266,N_1455);
nand U1825 (N_1825,In_771,N_1153);
and U1826 (N_1826,N_1322,N_1498);
and U1827 (N_1827,In_1159,N_1737);
xor U1828 (N_1828,N_564,N_1670);
xor U1829 (N_1829,N_1736,N_1595);
nor U1830 (N_1830,N_1770,N_1434);
xor U1831 (N_1831,N_235,In_855);
xnor U1832 (N_1832,N_1648,N_114);
and U1833 (N_1833,N_1694,In_1860);
nor U1834 (N_1834,N_1285,N_1492);
and U1835 (N_1835,N_1623,N_1672);
and U1836 (N_1836,In_1257,In_498);
and U1837 (N_1837,N_1312,N_1300);
and U1838 (N_1838,In_1430,In_1830);
nor U1839 (N_1839,N_1728,N_1647);
and U1840 (N_1840,N_45,N_1239);
nand U1841 (N_1841,N_1767,N_1751);
nand U1842 (N_1842,N_393,N_1461);
nor U1843 (N_1843,N_853,N_1236);
xnor U1844 (N_1844,N_1723,N_1206);
and U1845 (N_1845,N_1749,N_1731);
nand U1846 (N_1846,N_1640,N_1755);
or U1847 (N_1847,N_753,N_1205);
nor U1848 (N_1848,N_1462,In_15);
xor U1849 (N_1849,In_549,N_90);
xor U1850 (N_1850,N_1787,In_2477);
or U1851 (N_1851,N_786,N_1137);
nor U1852 (N_1852,N_973,N_329);
nand U1853 (N_1853,N_1587,In_49);
xor U1854 (N_1854,N_1049,N_1280);
and U1855 (N_1855,N_1311,N_919);
or U1856 (N_1856,N_1686,N_1265);
xor U1857 (N_1857,N_1084,N_1762);
or U1858 (N_1858,N_1000,N_1798);
and U1859 (N_1859,N_1564,N_1227);
or U1860 (N_1860,In_1199,N_1641);
nand U1861 (N_1861,N_504,N_1739);
and U1862 (N_1862,N_1758,N_1554);
and U1863 (N_1863,N_1620,In_1818);
or U1864 (N_1864,N_1592,In_626);
or U1865 (N_1865,In_1327,N_1653);
nor U1866 (N_1866,In_2090,N_1025);
or U1867 (N_1867,N_792,In_1896);
and U1868 (N_1868,In_1270,N_1149);
or U1869 (N_1869,N_1742,N_1195);
and U1870 (N_1870,N_698,N_1625);
nand U1871 (N_1871,In_358,N_1481);
nor U1872 (N_1872,In_236,In_733);
or U1873 (N_1873,N_1466,N_856);
nand U1874 (N_1874,N_524,N_1643);
nand U1875 (N_1875,N_1661,N_465);
nor U1876 (N_1876,In_1157,In_1350);
nor U1877 (N_1877,In_700,N_1719);
xnor U1878 (N_1878,N_871,N_1679);
xor U1879 (N_1879,N_1448,N_1645);
and U1880 (N_1880,N_1231,N_1423);
and U1881 (N_1881,N_1438,N_601);
nor U1882 (N_1882,N_170,N_772);
or U1883 (N_1883,In_854,N_1703);
nand U1884 (N_1884,N_1668,In_2034);
or U1885 (N_1885,N_1248,N_1198);
nand U1886 (N_1886,N_1675,N_1710);
xnor U1887 (N_1887,N_1286,In_1452);
or U1888 (N_1888,N_1295,N_355);
and U1889 (N_1889,N_868,N_1654);
and U1890 (N_1890,In_1083,N_1705);
xnor U1891 (N_1891,N_1330,In_2134);
or U1892 (N_1892,N_519,N_1396);
nand U1893 (N_1893,N_1400,In_327);
xnor U1894 (N_1894,N_1408,In_55);
nor U1895 (N_1895,N_1333,N_1062);
nor U1896 (N_1896,N_1121,N_1766);
and U1897 (N_1897,N_1690,N_1436);
and U1898 (N_1898,N_283,N_1454);
and U1899 (N_1899,N_1520,In_1228);
or U1900 (N_1900,N_978,N_1734);
nor U1901 (N_1901,N_30,N_864);
nand U1902 (N_1902,N_1633,N_785);
xor U1903 (N_1903,N_1522,N_1680);
or U1904 (N_1904,In_154,In_1630);
and U1905 (N_1905,N_1768,In_1582);
xnor U1906 (N_1906,N_1617,N_1073);
nor U1907 (N_1907,N_238,N_1636);
xor U1908 (N_1908,N_1689,N_1512);
xor U1909 (N_1909,In_1955,N_1709);
nor U1910 (N_1910,N_1397,In_1609);
xnor U1911 (N_1911,N_1741,N_1417);
nand U1912 (N_1912,N_259,N_586);
or U1913 (N_1913,In_1011,N_1605);
or U1914 (N_1914,N_1788,N_967);
xnor U1915 (N_1915,N_877,N_1635);
nor U1916 (N_1916,N_942,N_1669);
and U1917 (N_1917,N_437,N_899);
xnor U1918 (N_1918,N_1795,In_426);
xnor U1919 (N_1919,In_304,N_567);
nor U1920 (N_1920,N_1194,N_1294);
nand U1921 (N_1921,N_250,N_1013);
nand U1922 (N_1922,N_1666,N_816);
and U1923 (N_1923,In_2291,N_1684);
or U1924 (N_1924,In_1988,N_1541);
nand U1925 (N_1925,In_460,N_1358);
xnor U1926 (N_1926,N_1657,N_1566);
and U1927 (N_1927,N_1720,N_1471);
xor U1928 (N_1928,In_1613,In_2136);
nor U1929 (N_1929,N_1786,In_1992);
nor U1930 (N_1930,N_1793,N_865);
and U1931 (N_1931,In_990,N_1510);
and U1932 (N_1932,N_1603,N_1615);
nand U1933 (N_1933,N_1796,In_2491);
xor U1934 (N_1934,N_1532,N_351);
or U1935 (N_1935,N_1558,N_1776);
and U1936 (N_1936,N_747,N_280);
and U1937 (N_1937,N_723,N_739);
and U1938 (N_1938,N_1638,N_1435);
xor U1939 (N_1939,N_750,N_518);
or U1940 (N_1940,N_1395,In_1044);
and U1941 (N_1941,N_1594,N_12);
and U1942 (N_1942,In_2401,N_1216);
or U1943 (N_1943,In_345,N_1659);
and U1944 (N_1944,N_1370,N_768);
nor U1945 (N_1945,N_1673,N_1561);
xor U1946 (N_1946,N_1360,In_892);
or U1947 (N_1947,N_1542,N_1658);
and U1948 (N_1948,N_1521,N_1214);
and U1949 (N_1949,N_1101,N_732);
nand U1950 (N_1950,In_1030,In_111);
xnor U1951 (N_1951,N_1744,N_1701);
nand U1952 (N_1952,N_189,In_992);
nand U1953 (N_1953,N_607,N_809);
nor U1954 (N_1954,N_1096,In_1526);
or U1955 (N_1955,N_1531,N_1392);
nand U1956 (N_1956,N_1609,N_1007);
and U1957 (N_1957,N_494,N_1490);
xnor U1958 (N_1958,N_1667,N_895);
or U1959 (N_1959,N_814,N_1637);
and U1960 (N_1960,N_1715,N_577);
and U1961 (N_1961,N_1217,N_1600);
and U1962 (N_1962,In_941,N_1624);
or U1963 (N_1963,In_670,N_708);
xor U1964 (N_1964,N_1201,In_799);
and U1965 (N_1965,N_1298,In_2110);
and U1966 (N_1966,N_1474,N_968);
xor U1967 (N_1967,N_1394,N_97);
xnor U1968 (N_1968,N_299,N_1611);
or U1969 (N_1969,N_1618,N_1381);
nor U1970 (N_1970,N_1760,N_1254);
and U1971 (N_1971,N_1769,N_1750);
and U1972 (N_1972,N_1702,In_1156);
nor U1973 (N_1973,N_1738,N_1544);
and U1974 (N_1974,In_1689,N_1161);
and U1975 (N_1975,N_1634,N_1745);
and U1976 (N_1976,In_864,N_1256);
or U1977 (N_1977,N_1629,In_2121);
nor U1978 (N_1978,In_1779,N_1186);
or U1979 (N_1979,N_1127,N_1502);
nand U1980 (N_1980,N_1613,N_995);
and U1981 (N_1981,In_1925,N_1427);
xnor U1982 (N_1982,N_1500,N_1726);
or U1983 (N_1983,N_621,N_1537);
nand U1984 (N_1984,In_1922,N_1536);
xor U1985 (N_1985,In_349,In_2424);
or U1986 (N_1986,N_1443,In_797);
nand U1987 (N_1987,N_1429,In_1998);
xnor U1988 (N_1988,In_2384,N_1775);
nand U1989 (N_1989,In_2181,In_780);
or U1990 (N_1990,In_1568,N_1379);
xor U1991 (N_1991,N_883,N_1147);
or U1992 (N_1992,N_1783,N_1559);
nor U1993 (N_1993,N_1700,N_1714);
xnor U1994 (N_1994,N_1308,N_1549);
or U1995 (N_1995,N_1538,In_874);
or U1996 (N_1996,N_1628,N_1262);
xor U1997 (N_1997,N_1445,N_1622);
nand U1998 (N_1998,N_1002,In_1361);
or U1999 (N_1999,N_1418,N_1425);
nor U2000 (N_2000,N_1363,N_1920);
or U2001 (N_2001,In_689,N_1486);
nand U2002 (N_2002,N_620,N_1772);
nand U2003 (N_2003,N_962,N_1748);
or U2004 (N_2004,In_1937,N_1789);
xnor U2005 (N_2005,N_1506,N_1890);
nor U2006 (N_2006,N_513,N_1627);
nand U2007 (N_2007,N_1884,N_1964);
or U2008 (N_2008,N_1458,N_1733);
and U2009 (N_2009,N_1724,N_1557);
and U2010 (N_2010,N_777,N_1146);
and U2011 (N_2011,In_213,N_1646);
xor U2012 (N_2012,N_1957,N_821);
and U2013 (N_2013,N_1598,In_2323);
or U2014 (N_2014,N_1958,In_1715);
and U2015 (N_2015,N_1784,N_1630);
nor U2016 (N_2016,N_1382,N_1432);
nand U2017 (N_2017,N_1871,N_1876);
nor U2018 (N_2018,N_1047,N_1852);
or U2019 (N_2019,N_423,N_1664);
and U2020 (N_2020,N_1057,N_1974);
nor U2021 (N_2021,N_1805,N_1993);
or U2022 (N_2022,N_1649,N_1885);
nor U2023 (N_2023,N_1763,N_1836);
nand U2024 (N_2024,N_1404,N_1870);
or U2025 (N_2025,In_1927,N_1946);
and U2026 (N_2026,N_1483,N_1371);
and U2027 (N_2027,N_1831,In_203);
xor U2028 (N_2028,In_269,N_1963);
and U2029 (N_2029,N_734,N_1819);
xnor U2030 (N_2030,N_1511,N_1969);
nor U2031 (N_2031,N_1862,N_1508);
xnor U2032 (N_2032,In_553,N_106);
nor U2033 (N_2033,In_2075,N_1916);
or U2034 (N_2034,N_1116,N_1809);
and U2035 (N_2035,N_1516,N_1951);
nor U2036 (N_2036,N_1984,N_1687);
and U2037 (N_2037,N_1971,N_1746);
xor U2038 (N_2038,N_1813,N_1817);
or U2039 (N_2039,N_1893,In_324);
xor U2040 (N_2040,N_1562,N_1721);
and U2041 (N_2041,N_690,N_1843);
xor U2042 (N_2042,N_1621,N_1923);
and U2043 (N_2043,N_1868,N_1773);
xor U2044 (N_2044,N_1495,N_1055);
xnor U2045 (N_2045,N_1393,N_1691);
nand U2046 (N_2046,N_1612,In_2120);
and U2047 (N_2047,N_72,N_1249);
xor U2048 (N_2048,N_1291,N_1965);
and U2049 (N_2049,N_1730,N_1892);
nand U2050 (N_2050,N_1759,N_1921);
nand U2051 (N_2051,In_156,N_1610);
or U2052 (N_2052,N_401,N_1475);
nand U2053 (N_2053,N_1880,In_1180);
or U2054 (N_2054,N_1922,N_1780);
nand U2055 (N_2055,N_1879,N_1955);
xnor U2056 (N_2056,N_879,In_1607);
nand U2057 (N_2057,In_1828,N_551);
and U2058 (N_2058,N_397,N_1947);
xnor U2059 (N_2059,N_1891,N_1851);
or U2060 (N_2060,N_520,N_1507);
or U2061 (N_2061,N_719,N_1696);
xnor U2062 (N_2062,N_1590,N_1977);
xor U2063 (N_2063,N_1846,N_1452);
nor U2064 (N_2064,N_1631,N_1887);
and U2065 (N_2065,N_1695,N_1801);
or U2066 (N_2066,N_1639,N_1867);
and U2067 (N_2067,N_1925,N_1954);
and U2068 (N_2068,N_1962,N_291);
nand U2069 (N_2069,N_376,N_1662);
or U2070 (N_2070,N_1525,In_933);
xor U2071 (N_2071,N_1941,N_55);
nand U2072 (N_2072,N_1895,N_1883);
nand U2073 (N_2073,N_776,N_1844);
nand U2074 (N_2074,N_1674,N_269);
nand U2075 (N_2075,N_1764,In_1404);
nand U2076 (N_2076,N_1864,N_1509);
nand U2077 (N_2077,N_1241,N_1238);
xnor U2078 (N_2078,N_1953,N_1856);
nor U2079 (N_2079,N_1944,N_1790);
nand U2080 (N_2080,N_1901,N_1825);
nand U2081 (N_2081,N_802,In_1623);
xor U2082 (N_2082,N_1820,N_1881);
nor U2083 (N_2083,N_1681,In_1098);
or U2084 (N_2084,N_1812,N_1990);
nor U2085 (N_2085,N_847,N_1910);
or U2086 (N_2086,N_1688,N_1827);
xnor U2087 (N_2087,N_1338,N_1806);
nand U2088 (N_2088,N_1685,N_1677);
nor U2089 (N_2089,N_1882,N_1913);
or U2090 (N_2090,N_1829,N_1799);
nor U2091 (N_2091,N_1911,N_1929);
nor U2092 (N_2092,N_1842,N_1995);
xnor U2093 (N_2093,N_306,N_1287);
and U2094 (N_2094,In_257,N_1431);
nand U2095 (N_2095,In_1002,N_1950);
xor U2096 (N_2096,N_1952,N_1140);
nand U2097 (N_2097,N_1792,N_1948);
or U2098 (N_2098,N_1533,N_1752);
and U2099 (N_2099,N_1735,In_264);
nand U2100 (N_2100,N_1811,N_1903);
and U2101 (N_2101,N_1575,N_1663);
nor U2102 (N_2102,N_1979,In_2246);
or U2103 (N_2103,N_1215,N_1794);
and U2104 (N_2104,N_1938,N_1945);
and U2105 (N_2105,N_1830,N_100);
or U2106 (N_2106,N_745,N_272);
nor U2107 (N_2107,N_1837,N_1608);
xnor U2108 (N_2108,N_1565,N_1514);
nor U2109 (N_2109,N_1899,N_1441);
nor U2110 (N_2110,N_1898,N_679);
and U2111 (N_2111,N_1526,N_1973);
xor U2112 (N_2112,In_59,N_1835);
nand U2113 (N_2113,N_1968,N_1524);
or U2114 (N_2114,N_1344,N_1918);
nor U2115 (N_2115,N_1599,N_699);
and U2116 (N_2116,N_1854,N_1814);
nor U2117 (N_2117,N_1271,N_584);
nand U2118 (N_2118,N_1547,N_1896);
nand U2119 (N_2119,N_1606,N_1998);
xnor U2120 (N_2120,N_1626,N_1912);
xnor U2121 (N_2121,N_1199,N_1992);
or U2122 (N_2122,N_1157,N_371);
and U2123 (N_2123,N_1861,N_1902);
nor U2124 (N_2124,N_1897,N_1939);
nand U2125 (N_2125,N_1616,N_887);
nor U2126 (N_2126,N_650,N_1845);
or U2127 (N_2127,N_1942,N_1777);
xor U2128 (N_2128,N_1915,N_1906);
xnor U2129 (N_2129,N_1676,N_1527);
nor U2130 (N_2130,N_1267,N_1833);
and U2131 (N_2131,N_1220,N_1401);
nor U2132 (N_2132,In_2479,N_1976);
nand U2133 (N_2133,N_982,N_1574);
or U2134 (N_2134,N_1997,N_1779);
nor U2135 (N_2135,N_1934,N_1888);
xor U2136 (N_2136,N_1988,N_1224);
and U2137 (N_2137,N_1889,N_1176);
or U2138 (N_2138,N_436,In_2038);
nor U2139 (N_2139,N_1771,In_724);
and U2140 (N_2140,N_1900,N_958);
nand U2141 (N_2141,N_1136,N_1860);
nand U2142 (N_2142,N_1826,N_1960);
nor U2143 (N_2143,N_1834,In_44);
xnor U2144 (N_2144,In_1450,N_1430);
nor U2145 (N_2145,N_1859,N_638);
nand U2146 (N_2146,In_437,N_1274);
and U2147 (N_2147,N_1816,N_1276);
xor U2148 (N_2148,N_1704,N_1914);
nor U2149 (N_2149,N_1754,N_1838);
nor U2150 (N_2150,N_1211,N_1716);
nand U2151 (N_2151,N_1774,In_1292);
nand U2152 (N_2152,N_1908,N_1119);
or U2153 (N_2153,N_1717,N_1602);
nor U2154 (N_2154,N_1247,In_1169);
and U2155 (N_2155,N_1909,N_890);
or U2156 (N_2156,N_1824,N_1718);
nand U2157 (N_2157,In_965,N_1810);
xnor U2158 (N_2158,N_1607,N_1874);
nor U2159 (N_2159,In_1766,N_1800);
nor U2160 (N_2160,N_1869,N_1930);
nand U2161 (N_2161,N_1576,N_1850);
nand U2162 (N_2162,N_1919,N_1943);
nor U2163 (N_2163,N_1933,N_1797);
and U2164 (N_2164,N_1994,N_1936);
nor U2165 (N_2165,In_73,N_1985);
nor U2166 (N_2166,N_1865,N_1651);
and U2167 (N_2167,N_1697,N_1927);
nor U2168 (N_2168,N_1935,In_185);
and U2169 (N_2169,N_1907,N_308);
or U2170 (N_2170,In_1441,N_1937);
nand U2171 (N_2171,N_1847,N_1713);
xnor U2172 (N_2172,N_1818,N_1359);
or U2173 (N_2173,N_1193,N_1148);
nor U2174 (N_2174,N_1875,N_1409);
nand U2175 (N_2175,N_1039,N_1857);
nor U2176 (N_2176,N_1828,N_1975);
and U2177 (N_2177,N_1152,In_2211);
and U2178 (N_2178,N_1706,N_474);
nand U2179 (N_2179,N_1785,N_1832);
xor U2180 (N_2180,N_400,N_1196);
nor U2181 (N_2181,N_1644,N_1235);
nand U2182 (N_2182,N_1822,N_1683);
xnor U2183 (N_2183,In_834,N_1949);
nand U2184 (N_2184,N_703,N_1981);
or U2185 (N_2185,N_1878,N_1804);
or U2186 (N_2186,N_1999,N_727);
xnor U2187 (N_2187,N_1987,N_1699);
nand U2188 (N_2188,N_1991,N_1523);
nor U2189 (N_2189,N_1210,N_1399);
or U2190 (N_2190,In_325,N_1904);
and U2191 (N_2191,N_1094,N_1940);
and U2192 (N_2192,N_1853,N_1926);
xnor U2193 (N_2193,N_910,N_1970);
nand U2194 (N_2194,N_1614,N_1849);
and U2195 (N_2195,N_1894,N_1966);
or U2196 (N_2196,N_1886,N_1453);
or U2197 (N_2197,N_1928,N_1747);
nor U2198 (N_2198,N_1841,N_1403);
xor U2199 (N_2199,N_1266,In_1060);
xnor U2200 (N_2200,N_2106,N_2133);
xnor U2201 (N_2201,N_1863,N_1515);
xor U2202 (N_2202,N_1996,N_2045);
or U2203 (N_2203,N_2055,N_2159);
or U2204 (N_2204,N_2130,N_2198);
and U2205 (N_2205,N_2164,N_2054);
nor U2206 (N_2206,N_2094,In_763);
and U2207 (N_2207,N_2113,N_2043);
or U2208 (N_2208,In_925,N_1808);
nand U2209 (N_2209,N_1756,N_2049);
and U2210 (N_2210,N_2158,N_2074);
and U2211 (N_2211,N_2044,N_1807);
nor U2212 (N_2212,N_2097,In_419);
or U2213 (N_2213,N_2003,N_2110);
xor U2214 (N_2214,N_2051,N_2041);
nor U2215 (N_2215,N_2131,N_2023);
nand U2216 (N_2216,In_1125,In_2053);
and U2217 (N_2217,N_1032,In_2061);
nand U2218 (N_2218,N_2128,N_2191);
and U2219 (N_2219,N_2121,N_1080);
or U2220 (N_2220,N_2180,N_1729);
or U2221 (N_2221,N_2085,N_1803);
and U2222 (N_2222,N_2013,N_2040);
and U2223 (N_2223,N_2009,N_1983);
and U2224 (N_2224,N_2114,In_2175);
nand U2225 (N_2225,N_2033,N_2143);
and U2226 (N_2226,N_1494,N_1961);
xor U2227 (N_2227,N_2064,N_2194);
nand U2228 (N_2228,N_2118,N_2095);
or U2229 (N_2229,N_2098,N_1858);
nand U2230 (N_2230,N_2101,N_1732);
xor U2231 (N_2231,N_2070,N_1743);
or U2232 (N_2232,N_2122,N_1781);
nand U2233 (N_2233,N_2160,N_2112);
xor U2234 (N_2234,N_2026,N_774);
xor U2235 (N_2235,N_2080,N_1956);
nor U2236 (N_2236,N_1931,N_2192);
xor U2237 (N_2237,N_2039,N_2020);
nor U2238 (N_2238,N_2116,N_2109);
nor U2239 (N_2239,N_1334,N_2069);
nor U2240 (N_2240,N_1692,N_2005);
or U2241 (N_2241,N_709,N_2156);
xor U2242 (N_2242,N_2058,N_2030);
nand U2243 (N_2243,N_227,N_1398);
xnor U2244 (N_2244,N_2000,N_2016);
and U2245 (N_2245,N_2084,N_2086);
nor U2246 (N_2246,N_2042,N_2048);
xor U2247 (N_2247,N_2150,N_2066);
or U2248 (N_2248,N_2171,N_2186);
xor U2249 (N_2249,N_1642,N_2136);
nor U2250 (N_2250,N_2050,N_1982);
or U2251 (N_2251,N_2135,N_2183);
or U2252 (N_2252,N_2125,N_2149);
nand U2253 (N_2253,N_2021,N_2142);
nand U2254 (N_2254,N_2046,N_2001);
nor U2255 (N_2255,N_2178,N_1839);
or U2256 (N_2256,N_2068,N_2185);
nor U2257 (N_2257,N_1978,N_1980);
nor U2258 (N_2258,In_1049,N_2134);
nor U2259 (N_2259,N_1840,N_2197);
nand U2260 (N_2260,N_1707,N_2129);
nor U2261 (N_2261,In_1946,N_1823);
xor U2262 (N_2262,N_1791,N_2189);
nand U2263 (N_2263,N_2190,N_2062);
and U2264 (N_2264,In_136,N_2088);
and U2265 (N_2265,N_1924,N_2014);
and U2266 (N_2266,N_1601,N_1778);
and U2267 (N_2267,N_2004,N_1125);
xnor U2268 (N_2268,N_1604,N_2127);
nor U2269 (N_2269,N_2019,N_1553);
and U2270 (N_2270,N_2120,N_2154);
or U2271 (N_2271,N_876,N_2092);
or U2272 (N_2272,N_2187,N_2123);
and U2273 (N_2273,N_2162,N_1253);
or U2274 (N_2274,N_2018,N_2163);
nand U2275 (N_2275,N_2061,N_2107);
and U2276 (N_2276,N_2139,N_2093);
xnor U2277 (N_2277,N_2083,N_2007);
nand U2278 (N_2278,N_2132,N_2047);
xnor U2279 (N_2279,N_2027,N_2028);
or U2280 (N_2280,N_2024,N_2029);
nor U2281 (N_2281,N_2105,N_1802);
nor U2282 (N_2282,N_1972,N_2071);
and U2283 (N_2283,N_1632,N_1855);
nor U2284 (N_2284,N_2111,In_1874);
xnor U2285 (N_2285,N_2165,N_1873);
or U2286 (N_2286,N_2034,N_2168);
or U2287 (N_2287,N_1866,N_2052);
xor U2288 (N_2288,N_1917,N_1989);
and U2289 (N_2289,N_2072,N_2090);
or U2290 (N_2290,N_2148,N_2182);
and U2291 (N_2291,N_2091,N_1491);
or U2292 (N_2292,N_2119,N_2184);
nor U2293 (N_2293,N_2059,In_350);
and U2294 (N_2294,N_2181,N_2126);
nor U2295 (N_2295,N_2144,N_1821);
xor U2296 (N_2296,N_2137,N_1725);
xnor U2297 (N_2297,N_2177,N_2169);
or U2298 (N_2298,N_2002,N_2032);
and U2299 (N_2299,N_2057,N_2108);
xor U2300 (N_2300,N_2141,N_2195);
xnor U2301 (N_2301,N_2012,N_2117);
nand U2302 (N_2302,N_1010,N_2031);
nand U2303 (N_2303,N_2008,N_2087);
and U2304 (N_2304,In_814,In_528);
xnor U2305 (N_2305,N_1905,N_1932);
or U2306 (N_2306,N_2081,N_2124);
and U2307 (N_2307,N_2060,N_2166);
nor U2308 (N_2308,N_1588,N_2151);
nand U2309 (N_2309,N_2179,N_2076);
xnor U2310 (N_2310,N_2010,N_68);
xor U2311 (N_2311,N_2073,N_1488);
xnor U2312 (N_2312,N_1019,N_1493);
xor U2313 (N_2313,N_2146,N_2065);
or U2314 (N_2314,N_2152,N_1087);
and U2315 (N_2315,N_2025,N_2056);
xor U2316 (N_2316,N_2196,N_2036);
and U2317 (N_2317,N_2038,N_1877);
and U2318 (N_2318,N_2145,N_2063);
or U2319 (N_2319,N_2103,N_2089);
or U2320 (N_2320,N_1967,N_433);
nor U2321 (N_2321,N_1387,N_2102);
and U2322 (N_2322,N_2167,N_1652);
or U2323 (N_2323,N_2078,N_2174);
nor U2324 (N_2324,N_2157,N_2006);
or U2325 (N_2325,N_1765,N_1753);
xnor U2326 (N_2326,N_2172,N_1848);
or U2327 (N_2327,N_2140,N_2115);
xnor U2328 (N_2328,N_2138,N_1467);
xor U2329 (N_2329,N_2175,N_2082);
xor U2330 (N_2330,N_2096,N_1650);
or U2331 (N_2331,N_2147,N_2075);
or U2332 (N_2332,N_2104,N_1782);
or U2333 (N_2333,N_1660,N_2176);
nor U2334 (N_2334,N_2022,N_2193);
nor U2335 (N_2335,N_1424,N_2100);
or U2336 (N_2336,N_1986,N_1416);
nand U2337 (N_2337,N_2199,N_2099);
xor U2338 (N_2338,N_1030,N_2067);
nor U2339 (N_2339,N_1374,N_2079);
nand U2340 (N_2340,N_1872,N_2037);
xor U2341 (N_2341,N_2053,N_1426);
or U2342 (N_2342,N_2153,N_2035);
xor U2343 (N_2343,N_1413,N_2017);
nand U2344 (N_2344,N_2155,In_1008);
or U2345 (N_2345,N_2170,N_2015);
and U2346 (N_2346,N_2077,N_2188);
and U2347 (N_2347,N_1959,N_2161);
nand U2348 (N_2348,N_2011,N_1727);
xor U2349 (N_2349,N_2173,N_1815);
nor U2350 (N_2350,N_2072,N_2076);
nand U2351 (N_2351,N_2083,N_2163);
nor U2352 (N_2352,N_2194,N_1125);
and U2353 (N_2353,N_1334,N_876);
nand U2354 (N_2354,N_2021,N_2061);
xor U2355 (N_2355,N_2072,N_2097);
and U2356 (N_2356,N_1632,N_2069);
nor U2357 (N_2357,N_1765,N_2085);
nor U2358 (N_2358,N_2029,N_2116);
and U2359 (N_2359,N_2080,N_1978);
nor U2360 (N_2360,N_2143,N_1642);
nor U2361 (N_2361,N_1732,N_1493);
xor U2362 (N_2362,N_2065,N_2132);
or U2363 (N_2363,N_2160,N_2053);
nor U2364 (N_2364,N_2114,In_1049);
nand U2365 (N_2365,N_2027,N_2186);
xor U2366 (N_2366,N_2173,N_2068);
nand U2367 (N_2367,N_2123,N_2177);
or U2368 (N_2368,N_2189,N_1413);
or U2369 (N_2369,N_1125,N_1387);
xnor U2370 (N_2370,N_2074,N_2129);
nand U2371 (N_2371,N_2164,N_2072);
xnor U2372 (N_2372,N_2048,N_2137);
and U2373 (N_2373,N_1978,N_2086);
or U2374 (N_2374,N_2005,N_709);
xnor U2375 (N_2375,N_2006,N_2047);
or U2376 (N_2376,N_2117,N_1652);
and U2377 (N_2377,N_2159,In_925);
nor U2378 (N_2378,N_2049,N_1398);
nand U2379 (N_2379,N_2036,N_1972);
and U2380 (N_2380,N_2193,N_2138);
nor U2381 (N_2381,N_2192,N_1917);
nand U2382 (N_2382,N_1725,N_2157);
and U2383 (N_2383,N_2154,N_1967);
and U2384 (N_2384,N_2117,N_2067);
nor U2385 (N_2385,N_1765,N_2185);
xor U2386 (N_2386,N_2117,In_2175);
nand U2387 (N_2387,N_2031,N_2009);
and U2388 (N_2388,N_1839,N_1488);
nor U2389 (N_2389,N_2086,N_1743);
xor U2390 (N_2390,N_2150,N_2008);
and U2391 (N_2391,N_2146,N_2152);
nor U2392 (N_2392,N_1823,N_1808);
nand U2393 (N_2393,N_2092,N_1601);
or U2394 (N_2394,In_1008,N_2046);
nand U2395 (N_2395,N_2008,N_1467);
and U2396 (N_2396,N_1729,N_2031);
nor U2397 (N_2397,In_763,N_227);
xor U2398 (N_2398,N_2105,N_2189);
or U2399 (N_2399,N_68,N_1426);
or U2400 (N_2400,N_2322,N_2397);
and U2401 (N_2401,N_2362,N_2393);
nor U2402 (N_2402,N_2355,N_2279);
or U2403 (N_2403,N_2334,N_2251);
nand U2404 (N_2404,N_2384,N_2388);
and U2405 (N_2405,N_2260,N_2232);
xnor U2406 (N_2406,N_2220,N_2230);
or U2407 (N_2407,N_2309,N_2285);
nand U2408 (N_2408,N_2201,N_2207);
xnor U2409 (N_2409,N_2371,N_2369);
nor U2410 (N_2410,N_2329,N_2389);
nor U2411 (N_2411,N_2200,N_2209);
nor U2412 (N_2412,N_2244,N_2270);
and U2413 (N_2413,N_2205,N_2265);
nand U2414 (N_2414,N_2304,N_2312);
xor U2415 (N_2415,N_2375,N_2242);
nand U2416 (N_2416,N_2229,N_2317);
and U2417 (N_2417,N_2239,N_2331);
nand U2418 (N_2418,N_2213,N_2296);
or U2419 (N_2419,N_2225,N_2315);
and U2420 (N_2420,N_2337,N_2376);
or U2421 (N_2421,N_2214,N_2233);
nor U2422 (N_2422,N_2372,N_2287);
nor U2423 (N_2423,N_2215,N_2257);
nand U2424 (N_2424,N_2380,N_2347);
nor U2425 (N_2425,N_2301,N_2367);
and U2426 (N_2426,N_2221,N_2396);
nor U2427 (N_2427,N_2321,N_2250);
xnor U2428 (N_2428,N_2210,N_2390);
nand U2429 (N_2429,N_2306,N_2327);
and U2430 (N_2430,N_2359,N_2264);
and U2431 (N_2431,N_2202,N_2267);
nand U2432 (N_2432,N_2252,N_2256);
and U2433 (N_2433,N_2330,N_2311);
xnor U2434 (N_2434,N_2275,N_2349);
or U2435 (N_2435,N_2262,N_2392);
nand U2436 (N_2436,N_2368,N_2382);
nand U2437 (N_2437,N_2395,N_2236);
nor U2438 (N_2438,N_2356,N_2273);
nor U2439 (N_2439,N_2297,N_2295);
nor U2440 (N_2440,N_2268,N_2383);
or U2441 (N_2441,N_2386,N_2319);
or U2442 (N_2442,N_2364,N_2303);
nor U2443 (N_2443,N_2313,N_2370);
xor U2444 (N_2444,N_2222,N_2294);
nor U2445 (N_2445,N_2269,N_2217);
nand U2446 (N_2446,N_2219,N_2240);
xnor U2447 (N_2447,N_2248,N_2344);
or U2448 (N_2448,N_2208,N_2353);
xnor U2449 (N_2449,N_2212,N_2308);
nand U2450 (N_2450,N_2282,N_2211);
nand U2451 (N_2451,N_2288,N_2358);
nor U2452 (N_2452,N_2290,N_2379);
nand U2453 (N_2453,N_2351,N_2314);
and U2454 (N_2454,N_2292,N_2340);
or U2455 (N_2455,N_2223,N_2276);
nor U2456 (N_2456,N_2326,N_2332);
nand U2457 (N_2457,N_2398,N_2298);
and U2458 (N_2458,N_2310,N_2307);
and U2459 (N_2459,N_2373,N_2305);
or U2460 (N_2460,N_2231,N_2255);
nand U2461 (N_2461,N_2366,N_2234);
xor U2462 (N_2462,N_2399,N_2226);
or U2463 (N_2463,N_2289,N_2258);
or U2464 (N_2464,N_2357,N_2235);
nor U2465 (N_2465,N_2228,N_2352);
xor U2466 (N_2466,N_2254,N_2291);
nor U2467 (N_2467,N_2339,N_2361);
nand U2468 (N_2468,N_2363,N_2272);
nor U2469 (N_2469,N_2378,N_2391);
and U2470 (N_2470,N_2284,N_2342);
xnor U2471 (N_2471,N_2227,N_2320);
and U2472 (N_2472,N_2224,N_2323);
nor U2473 (N_2473,N_2274,N_2237);
and U2474 (N_2474,N_2374,N_2336);
nand U2475 (N_2475,N_2281,N_2266);
nand U2476 (N_2476,N_2238,N_2206);
or U2477 (N_2477,N_2316,N_2385);
nor U2478 (N_2478,N_2299,N_2345);
and U2479 (N_2479,N_2247,N_2338);
nand U2480 (N_2480,N_2377,N_2325);
nor U2481 (N_2481,N_2216,N_2354);
nand U2482 (N_2482,N_2271,N_2245);
xnor U2483 (N_2483,N_2203,N_2335);
or U2484 (N_2484,N_2394,N_2300);
nand U2485 (N_2485,N_2249,N_2293);
nand U2486 (N_2486,N_2253,N_2218);
xnor U2487 (N_2487,N_2318,N_2241);
nand U2488 (N_2488,N_2278,N_2324);
and U2489 (N_2489,N_2350,N_2341);
or U2490 (N_2490,N_2387,N_2343);
nor U2491 (N_2491,N_2204,N_2328);
nor U2492 (N_2492,N_2365,N_2346);
xor U2493 (N_2493,N_2360,N_2261);
nor U2494 (N_2494,N_2246,N_2348);
nor U2495 (N_2495,N_2283,N_2259);
and U2496 (N_2496,N_2333,N_2263);
or U2497 (N_2497,N_2381,N_2286);
or U2498 (N_2498,N_2277,N_2243);
xor U2499 (N_2499,N_2280,N_2302);
and U2500 (N_2500,N_2385,N_2389);
xor U2501 (N_2501,N_2393,N_2286);
nor U2502 (N_2502,N_2275,N_2336);
nand U2503 (N_2503,N_2397,N_2363);
xnor U2504 (N_2504,N_2313,N_2321);
and U2505 (N_2505,N_2309,N_2248);
or U2506 (N_2506,N_2272,N_2332);
or U2507 (N_2507,N_2270,N_2351);
nor U2508 (N_2508,N_2212,N_2399);
nor U2509 (N_2509,N_2384,N_2350);
and U2510 (N_2510,N_2250,N_2387);
nand U2511 (N_2511,N_2236,N_2324);
nor U2512 (N_2512,N_2328,N_2311);
xnor U2513 (N_2513,N_2383,N_2261);
nor U2514 (N_2514,N_2217,N_2385);
nand U2515 (N_2515,N_2249,N_2266);
nand U2516 (N_2516,N_2384,N_2252);
xor U2517 (N_2517,N_2389,N_2276);
and U2518 (N_2518,N_2293,N_2367);
or U2519 (N_2519,N_2236,N_2282);
and U2520 (N_2520,N_2390,N_2290);
xnor U2521 (N_2521,N_2353,N_2228);
and U2522 (N_2522,N_2223,N_2337);
nand U2523 (N_2523,N_2338,N_2361);
xor U2524 (N_2524,N_2218,N_2397);
nor U2525 (N_2525,N_2244,N_2227);
xor U2526 (N_2526,N_2371,N_2256);
nand U2527 (N_2527,N_2366,N_2237);
xor U2528 (N_2528,N_2285,N_2245);
xnor U2529 (N_2529,N_2289,N_2204);
nor U2530 (N_2530,N_2280,N_2354);
xnor U2531 (N_2531,N_2384,N_2361);
or U2532 (N_2532,N_2294,N_2202);
nor U2533 (N_2533,N_2382,N_2248);
xor U2534 (N_2534,N_2279,N_2220);
nor U2535 (N_2535,N_2303,N_2291);
nor U2536 (N_2536,N_2380,N_2377);
and U2537 (N_2537,N_2241,N_2215);
nand U2538 (N_2538,N_2246,N_2329);
xor U2539 (N_2539,N_2330,N_2322);
and U2540 (N_2540,N_2274,N_2365);
nand U2541 (N_2541,N_2390,N_2332);
nand U2542 (N_2542,N_2272,N_2311);
and U2543 (N_2543,N_2369,N_2379);
nand U2544 (N_2544,N_2274,N_2297);
or U2545 (N_2545,N_2244,N_2398);
and U2546 (N_2546,N_2230,N_2228);
xor U2547 (N_2547,N_2381,N_2262);
nor U2548 (N_2548,N_2246,N_2275);
nor U2549 (N_2549,N_2283,N_2202);
xor U2550 (N_2550,N_2347,N_2217);
or U2551 (N_2551,N_2264,N_2323);
nor U2552 (N_2552,N_2372,N_2351);
nor U2553 (N_2553,N_2240,N_2367);
xor U2554 (N_2554,N_2326,N_2343);
nor U2555 (N_2555,N_2351,N_2368);
and U2556 (N_2556,N_2391,N_2305);
or U2557 (N_2557,N_2223,N_2366);
or U2558 (N_2558,N_2336,N_2265);
or U2559 (N_2559,N_2212,N_2299);
nor U2560 (N_2560,N_2368,N_2333);
nor U2561 (N_2561,N_2243,N_2225);
nand U2562 (N_2562,N_2245,N_2372);
and U2563 (N_2563,N_2334,N_2280);
xor U2564 (N_2564,N_2246,N_2303);
or U2565 (N_2565,N_2258,N_2315);
nand U2566 (N_2566,N_2226,N_2338);
or U2567 (N_2567,N_2352,N_2218);
nand U2568 (N_2568,N_2269,N_2353);
xnor U2569 (N_2569,N_2363,N_2222);
and U2570 (N_2570,N_2271,N_2264);
and U2571 (N_2571,N_2233,N_2224);
xnor U2572 (N_2572,N_2301,N_2249);
nor U2573 (N_2573,N_2328,N_2220);
or U2574 (N_2574,N_2223,N_2310);
nor U2575 (N_2575,N_2200,N_2284);
or U2576 (N_2576,N_2370,N_2291);
and U2577 (N_2577,N_2359,N_2251);
and U2578 (N_2578,N_2326,N_2206);
and U2579 (N_2579,N_2201,N_2217);
xnor U2580 (N_2580,N_2398,N_2206);
or U2581 (N_2581,N_2377,N_2399);
nand U2582 (N_2582,N_2266,N_2263);
nand U2583 (N_2583,N_2315,N_2285);
nand U2584 (N_2584,N_2219,N_2242);
nor U2585 (N_2585,N_2213,N_2255);
and U2586 (N_2586,N_2320,N_2288);
nor U2587 (N_2587,N_2316,N_2202);
xor U2588 (N_2588,N_2372,N_2318);
and U2589 (N_2589,N_2332,N_2366);
and U2590 (N_2590,N_2379,N_2323);
nand U2591 (N_2591,N_2268,N_2294);
and U2592 (N_2592,N_2244,N_2248);
nor U2593 (N_2593,N_2305,N_2287);
and U2594 (N_2594,N_2387,N_2238);
nand U2595 (N_2595,N_2235,N_2367);
or U2596 (N_2596,N_2362,N_2279);
and U2597 (N_2597,N_2267,N_2326);
nand U2598 (N_2598,N_2301,N_2354);
or U2599 (N_2599,N_2256,N_2331);
xor U2600 (N_2600,N_2400,N_2423);
nand U2601 (N_2601,N_2461,N_2505);
nor U2602 (N_2602,N_2441,N_2490);
and U2603 (N_2603,N_2426,N_2555);
or U2604 (N_2604,N_2554,N_2494);
or U2605 (N_2605,N_2513,N_2429);
or U2606 (N_2606,N_2553,N_2476);
and U2607 (N_2607,N_2497,N_2526);
nor U2608 (N_2608,N_2598,N_2542);
nor U2609 (N_2609,N_2449,N_2539);
nand U2610 (N_2610,N_2547,N_2588);
and U2611 (N_2611,N_2503,N_2491);
nor U2612 (N_2612,N_2499,N_2557);
and U2613 (N_2613,N_2474,N_2436);
xor U2614 (N_2614,N_2550,N_2482);
nand U2615 (N_2615,N_2402,N_2584);
nor U2616 (N_2616,N_2487,N_2463);
nor U2617 (N_2617,N_2439,N_2469);
and U2618 (N_2618,N_2475,N_2480);
nor U2619 (N_2619,N_2521,N_2485);
nand U2620 (N_2620,N_2498,N_2484);
xor U2621 (N_2621,N_2415,N_2442);
nand U2622 (N_2622,N_2473,N_2405);
xnor U2623 (N_2623,N_2593,N_2465);
xor U2624 (N_2624,N_2577,N_2541);
nor U2625 (N_2625,N_2417,N_2431);
and U2626 (N_2626,N_2430,N_2551);
nor U2627 (N_2627,N_2586,N_2447);
nand U2628 (N_2628,N_2422,N_2510);
or U2629 (N_2629,N_2414,N_2424);
or U2630 (N_2630,N_2599,N_2454);
nand U2631 (N_2631,N_2434,N_2570);
nor U2632 (N_2632,N_2457,N_2483);
and U2633 (N_2633,N_2408,N_2536);
xor U2634 (N_2634,N_2517,N_2410);
nand U2635 (N_2635,N_2563,N_2578);
xor U2636 (N_2636,N_2500,N_2466);
or U2637 (N_2637,N_2444,N_2501);
nor U2638 (N_2638,N_2428,N_2495);
or U2639 (N_2639,N_2573,N_2595);
and U2640 (N_2640,N_2549,N_2488);
and U2641 (N_2641,N_2458,N_2558);
or U2642 (N_2642,N_2425,N_2589);
and U2643 (N_2643,N_2443,N_2464);
or U2644 (N_2644,N_2533,N_2411);
and U2645 (N_2645,N_2560,N_2478);
nand U2646 (N_2646,N_2546,N_2416);
or U2647 (N_2647,N_2519,N_2534);
or U2648 (N_2648,N_2496,N_2508);
xnor U2649 (N_2649,N_2479,N_2568);
or U2650 (N_2650,N_2445,N_2587);
nor U2651 (N_2651,N_2407,N_2515);
xnor U2652 (N_2652,N_2453,N_2512);
nor U2653 (N_2653,N_2562,N_2531);
and U2654 (N_2654,N_2597,N_2530);
nor U2655 (N_2655,N_2520,N_2420);
and U2656 (N_2656,N_2450,N_2544);
or U2657 (N_2657,N_2507,N_2446);
nand U2658 (N_2658,N_2537,N_2418);
or U2659 (N_2659,N_2489,N_2459);
nor U2660 (N_2660,N_2566,N_2471);
and U2661 (N_2661,N_2561,N_2528);
xor U2662 (N_2662,N_2413,N_2427);
xor U2663 (N_2663,N_2467,N_2419);
xor U2664 (N_2664,N_2516,N_2506);
xnor U2665 (N_2665,N_2421,N_2511);
xor U2666 (N_2666,N_2460,N_2567);
nand U2667 (N_2667,N_2472,N_2559);
and U2668 (N_2668,N_2435,N_2532);
xnor U2669 (N_2669,N_2583,N_2452);
nor U2670 (N_2670,N_2575,N_2540);
nand U2671 (N_2671,N_2581,N_2451);
nor U2672 (N_2672,N_2590,N_2406);
nor U2673 (N_2673,N_2432,N_2509);
or U2674 (N_2674,N_2409,N_2455);
nand U2675 (N_2675,N_2569,N_2486);
or U2676 (N_2676,N_2504,N_2493);
and U2677 (N_2677,N_2574,N_2523);
xor U2678 (N_2678,N_2412,N_2535);
nor U2679 (N_2679,N_2582,N_2518);
xor U2680 (N_2680,N_2477,N_2448);
nand U2681 (N_2681,N_2545,N_2552);
or U2682 (N_2682,N_2456,N_2580);
nor U2683 (N_2683,N_2440,N_2524);
nor U2684 (N_2684,N_2522,N_2543);
nor U2685 (N_2685,N_2529,N_2538);
nor U2686 (N_2686,N_2591,N_2556);
nand U2687 (N_2687,N_2564,N_2492);
or U2688 (N_2688,N_2548,N_2579);
and U2689 (N_2689,N_2481,N_2571);
xnor U2690 (N_2690,N_2438,N_2594);
or U2691 (N_2691,N_2502,N_2404);
nand U2692 (N_2692,N_2514,N_2576);
nand U2693 (N_2693,N_2565,N_2433);
nand U2694 (N_2694,N_2527,N_2468);
nand U2695 (N_2695,N_2592,N_2437);
xnor U2696 (N_2696,N_2596,N_2403);
and U2697 (N_2697,N_2585,N_2470);
nand U2698 (N_2698,N_2525,N_2401);
and U2699 (N_2699,N_2572,N_2462);
and U2700 (N_2700,N_2565,N_2557);
or U2701 (N_2701,N_2500,N_2553);
nor U2702 (N_2702,N_2487,N_2537);
nand U2703 (N_2703,N_2465,N_2430);
xor U2704 (N_2704,N_2407,N_2439);
xor U2705 (N_2705,N_2427,N_2536);
or U2706 (N_2706,N_2561,N_2576);
nand U2707 (N_2707,N_2530,N_2589);
or U2708 (N_2708,N_2594,N_2490);
nor U2709 (N_2709,N_2431,N_2520);
nand U2710 (N_2710,N_2585,N_2514);
and U2711 (N_2711,N_2410,N_2452);
nand U2712 (N_2712,N_2433,N_2422);
and U2713 (N_2713,N_2514,N_2535);
nand U2714 (N_2714,N_2582,N_2413);
or U2715 (N_2715,N_2450,N_2429);
or U2716 (N_2716,N_2531,N_2509);
and U2717 (N_2717,N_2549,N_2538);
and U2718 (N_2718,N_2412,N_2425);
nand U2719 (N_2719,N_2414,N_2548);
nand U2720 (N_2720,N_2481,N_2585);
or U2721 (N_2721,N_2585,N_2510);
nand U2722 (N_2722,N_2582,N_2577);
nand U2723 (N_2723,N_2413,N_2491);
and U2724 (N_2724,N_2563,N_2400);
nand U2725 (N_2725,N_2570,N_2552);
xor U2726 (N_2726,N_2501,N_2550);
nor U2727 (N_2727,N_2536,N_2545);
nor U2728 (N_2728,N_2404,N_2589);
nand U2729 (N_2729,N_2400,N_2485);
nand U2730 (N_2730,N_2490,N_2476);
xnor U2731 (N_2731,N_2508,N_2469);
and U2732 (N_2732,N_2488,N_2490);
nand U2733 (N_2733,N_2518,N_2583);
and U2734 (N_2734,N_2469,N_2522);
or U2735 (N_2735,N_2451,N_2495);
and U2736 (N_2736,N_2458,N_2437);
nor U2737 (N_2737,N_2484,N_2405);
nand U2738 (N_2738,N_2536,N_2589);
nor U2739 (N_2739,N_2482,N_2513);
xnor U2740 (N_2740,N_2510,N_2579);
nand U2741 (N_2741,N_2468,N_2404);
or U2742 (N_2742,N_2445,N_2426);
or U2743 (N_2743,N_2474,N_2437);
nor U2744 (N_2744,N_2458,N_2577);
or U2745 (N_2745,N_2424,N_2437);
nand U2746 (N_2746,N_2484,N_2434);
or U2747 (N_2747,N_2408,N_2529);
xnor U2748 (N_2748,N_2500,N_2521);
xor U2749 (N_2749,N_2573,N_2552);
xor U2750 (N_2750,N_2483,N_2480);
and U2751 (N_2751,N_2505,N_2576);
xnor U2752 (N_2752,N_2496,N_2565);
or U2753 (N_2753,N_2517,N_2463);
xnor U2754 (N_2754,N_2459,N_2577);
or U2755 (N_2755,N_2495,N_2508);
or U2756 (N_2756,N_2434,N_2585);
or U2757 (N_2757,N_2429,N_2570);
or U2758 (N_2758,N_2536,N_2403);
xnor U2759 (N_2759,N_2591,N_2464);
or U2760 (N_2760,N_2571,N_2428);
or U2761 (N_2761,N_2566,N_2542);
nand U2762 (N_2762,N_2537,N_2477);
nor U2763 (N_2763,N_2471,N_2533);
xor U2764 (N_2764,N_2543,N_2479);
nand U2765 (N_2765,N_2455,N_2595);
nor U2766 (N_2766,N_2555,N_2453);
and U2767 (N_2767,N_2405,N_2465);
or U2768 (N_2768,N_2599,N_2504);
xor U2769 (N_2769,N_2448,N_2561);
nand U2770 (N_2770,N_2559,N_2597);
nand U2771 (N_2771,N_2434,N_2441);
and U2772 (N_2772,N_2428,N_2461);
or U2773 (N_2773,N_2464,N_2471);
nor U2774 (N_2774,N_2592,N_2508);
xor U2775 (N_2775,N_2473,N_2488);
xnor U2776 (N_2776,N_2593,N_2437);
nand U2777 (N_2777,N_2458,N_2568);
and U2778 (N_2778,N_2555,N_2586);
nand U2779 (N_2779,N_2506,N_2412);
xor U2780 (N_2780,N_2451,N_2458);
nor U2781 (N_2781,N_2586,N_2464);
xor U2782 (N_2782,N_2426,N_2576);
and U2783 (N_2783,N_2585,N_2519);
and U2784 (N_2784,N_2507,N_2598);
or U2785 (N_2785,N_2494,N_2599);
and U2786 (N_2786,N_2500,N_2537);
or U2787 (N_2787,N_2500,N_2410);
xnor U2788 (N_2788,N_2515,N_2477);
and U2789 (N_2789,N_2464,N_2469);
and U2790 (N_2790,N_2575,N_2439);
nand U2791 (N_2791,N_2550,N_2588);
or U2792 (N_2792,N_2494,N_2408);
or U2793 (N_2793,N_2463,N_2486);
and U2794 (N_2794,N_2534,N_2455);
nor U2795 (N_2795,N_2485,N_2445);
and U2796 (N_2796,N_2511,N_2428);
and U2797 (N_2797,N_2423,N_2586);
xor U2798 (N_2798,N_2518,N_2508);
xor U2799 (N_2799,N_2583,N_2537);
nor U2800 (N_2800,N_2640,N_2724);
nand U2801 (N_2801,N_2672,N_2702);
xor U2802 (N_2802,N_2666,N_2773);
and U2803 (N_2803,N_2678,N_2617);
xnor U2804 (N_2804,N_2782,N_2708);
nor U2805 (N_2805,N_2777,N_2710);
xnor U2806 (N_2806,N_2712,N_2696);
xor U2807 (N_2807,N_2654,N_2604);
or U2808 (N_2808,N_2607,N_2749);
and U2809 (N_2809,N_2648,N_2693);
xnor U2810 (N_2810,N_2774,N_2615);
and U2811 (N_2811,N_2659,N_2759);
xor U2812 (N_2812,N_2677,N_2722);
or U2813 (N_2813,N_2704,N_2688);
and U2814 (N_2814,N_2653,N_2691);
xnor U2815 (N_2815,N_2682,N_2755);
nand U2816 (N_2816,N_2786,N_2713);
and U2817 (N_2817,N_2625,N_2668);
and U2818 (N_2818,N_2753,N_2634);
and U2819 (N_2819,N_2725,N_2621);
xnor U2820 (N_2820,N_2630,N_2729);
and U2821 (N_2821,N_2742,N_2697);
nand U2822 (N_2822,N_2798,N_2757);
and U2823 (N_2823,N_2718,N_2747);
nand U2824 (N_2824,N_2737,N_2767);
or U2825 (N_2825,N_2680,N_2783);
nand U2826 (N_2826,N_2730,N_2790);
nor U2827 (N_2827,N_2658,N_2652);
xor U2828 (N_2828,N_2735,N_2733);
or U2829 (N_2829,N_2768,N_2601);
and U2830 (N_2830,N_2665,N_2623);
nor U2831 (N_2831,N_2611,N_2674);
nor U2832 (N_2832,N_2631,N_2639);
nand U2833 (N_2833,N_2632,N_2787);
and U2834 (N_2834,N_2602,N_2720);
nor U2835 (N_2835,N_2663,N_2613);
xor U2836 (N_2836,N_2778,N_2703);
or U2837 (N_2837,N_2751,N_2647);
nand U2838 (N_2838,N_2771,N_2721);
xnor U2839 (N_2839,N_2740,N_2731);
xor U2840 (N_2840,N_2741,N_2627);
and U2841 (N_2841,N_2746,N_2662);
or U2842 (N_2842,N_2770,N_2709);
nor U2843 (N_2843,N_2637,N_2775);
nand U2844 (N_2844,N_2606,N_2707);
xor U2845 (N_2845,N_2656,N_2734);
and U2846 (N_2846,N_2686,N_2745);
nor U2847 (N_2847,N_2685,N_2792);
xor U2848 (N_2848,N_2761,N_2608);
or U2849 (N_2849,N_2797,N_2669);
xnor U2850 (N_2850,N_2781,N_2684);
nand U2851 (N_2851,N_2629,N_2732);
or U2852 (N_2852,N_2779,N_2650);
xnor U2853 (N_2853,N_2776,N_2641);
xor U2854 (N_2854,N_2766,N_2605);
nand U2855 (N_2855,N_2673,N_2785);
nand U2856 (N_2856,N_2603,N_2716);
xor U2857 (N_2857,N_2717,N_2763);
and U2858 (N_2858,N_2694,N_2645);
xor U2859 (N_2859,N_2743,N_2676);
nand U2860 (N_2860,N_2624,N_2799);
and U2861 (N_2861,N_2714,N_2610);
xor U2862 (N_2862,N_2679,N_2612);
xnor U2863 (N_2863,N_2633,N_2784);
or U2864 (N_2864,N_2618,N_2794);
or U2865 (N_2865,N_2657,N_2600);
or U2866 (N_2866,N_2636,N_2643);
and U2867 (N_2867,N_2628,N_2642);
nor U2868 (N_2868,N_2762,N_2681);
and U2869 (N_2869,N_2793,N_2796);
nand U2870 (N_2870,N_2614,N_2700);
nor U2871 (N_2871,N_2609,N_2698);
or U2872 (N_2872,N_2644,N_2736);
xnor U2873 (N_2873,N_2715,N_2620);
nand U2874 (N_2874,N_2789,N_2651);
xnor U2875 (N_2875,N_2769,N_2758);
xnor U2876 (N_2876,N_2754,N_2764);
xnor U2877 (N_2877,N_2728,N_2752);
and U2878 (N_2878,N_2727,N_2619);
or U2879 (N_2879,N_2780,N_2705);
xnor U2880 (N_2880,N_2711,N_2687);
or U2881 (N_2881,N_2664,N_2646);
and U2882 (N_2882,N_2756,N_2626);
or U2883 (N_2883,N_2791,N_2695);
and U2884 (N_2884,N_2671,N_2661);
nor U2885 (N_2885,N_2744,N_2788);
nor U2886 (N_2886,N_2748,N_2675);
nor U2887 (N_2887,N_2772,N_2765);
nor U2888 (N_2888,N_2706,N_2638);
nor U2889 (N_2889,N_2701,N_2616);
xnor U2890 (N_2890,N_2683,N_2649);
and U2891 (N_2891,N_2795,N_2670);
nor U2892 (N_2892,N_2738,N_2622);
or U2893 (N_2893,N_2739,N_2692);
nand U2894 (N_2894,N_2667,N_2660);
nor U2895 (N_2895,N_2655,N_2699);
or U2896 (N_2896,N_2723,N_2760);
or U2897 (N_2897,N_2726,N_2689);
xnor U2898 (N_2898,N_2635,N_2719);
xnor U2899 (N_2899,N_2750,N_2690);
and U2900 (N_2900,N_2635,N_2613);
xnor U2901 (N_2901,N_2698,N_2782);
xnor U2902 (N_2902,N_2659,N_2697);
or U2903 (N_2903,N_2727,N_2729);
nor U2904 (N_2904,N_2792,N_2791);
nand U2905 (N_2905,N_2799,N_2768);
and U2906 (N_2906,N_2704,N_2792);
or U2907 (N_2907,N_2685,N_2600);
or U2908 (N_2908,N_2602,N_2726);
xnor U2909 (N_2909,N_2679,N_2660);
xor U2910 (N_2910,N_2651,N_2688);
and U2911 (N_2911,N_2624,N_2720);
xor U2912 (N_2912,N_2707,N_2704);
and U2913 (N_2913,N_2774,N_2797);
and U2914 (N_2914,N_2612,N_2656);
or U2915 (N_2915,N_2663,N_2618);
nor U2916 (N_2916,N_2780,N_2799);
or U2917 (N_2917,N_2669,N_2692);
xnor U2918 (N_2918,N_2733,N_2706);
or U2919 (N_2919,N_2679,N_2673);
nand U2920 (N_2920,N_2725,N_2747);
nand U2921 (N_2921,N_2779,N_2700);
and U2922 (N_2922,N_2615,N_2690);
nor U2923 (N_2923,N_2774,N_2766);
nor U2924 (N_2924,N_2733,N_2621);
and U2925 (N_2925,N_2605,N_2785);
or U2926 (N_2926,N_2768,N_2681);
or U2927 (N_2927,N_2738,N_2617);
and U2928 (N_2928,N_2623,N_2631);
nand U2929 (N_2929,N_2787,N_2727);
or U2930 (N_2930,N_2608,N_2703);
or U2931 (N_2931,N_2605,N_2665);
and U2932 (N_2932,N_2783,N_2692);
and U2933 (N_2933,N_2706,N_2773);
nand U2934 (N_2934,N_2690,N_2777);
nand U2935 (N_2935,N_2733,N_2711);
and U2936 (N_2936,N_2778,N_2742);
nand U2937 (N_2937,N_2746,N_2644);
or U2938 (N_2938,N_2744,N_2648);
nor U2939 (N_2939,N_2796,N_2790);
xor U2940 (N_2940,N_2725,N_2695);
and U2941 (N_2941,N_2764,N_2725);
and U2942 (N_2942,N_2734,N_2617);
and U2943 (N_2943,N_2664,N_2727);
or U2944 (N_2944,N_2632,N_2600);
nor U2945 (N_2945,N_2774,N_2656);
and U2946 (N_2946,N_2680,N_2635);
nand U2947 (N_2947,N_2724,N_2617);
nor U2948 (N_2948,N_2626,N_2786);
or U2949 (N_2949,N_2772,N_2650);
and U2950 (N_2950,N_2644,N_2741);
and U2951 (N_2951,N_2680,N_2696);
and U2952 (N_2952,N_2776,N_2699);
nor U2953 (N_2953,N_2712,N_2737);
nor U2954 (N_2954,N_2703,N_2755);
and U2955 (N_2955,N_2744,N_2619);
and U2956 (N_2956,N_2777,N_2702);
nor U2957 (N_2957,N_2600,N_2787);
and U2958 (N_2958,N_2790,N_2731);
xnor U2959 (N_2959,N_2699,N_2607);
and U2960 (N_2960,N_2691,N_2724);
nand U2961 (N_2961,N_2626,N_2679);
nor U2962 (N_2962,N_2769,N_2625);
nand U2963 (N_2963,N_2615,N_2650);
xnor U2964 (N_2964,N_2642,N_2629);
xor U2965 (N_2965,N_2771,N_2655);
xor U2966 (N_2966,N_2662,N_2675);
nand U2967 (N_2967,N_2756,N_2760);
and U2968 (N_2968,N_2656,N_2748);
xnor U2969 (N_2969,N_2677,N_2736);
xnor U2970 (N_2970,N_2799,N_2735);
nor U2971 (N_2971,N_2792,N_2739);
nand U2972 (N_2972,N_2789,N_2719);
or U2973 (N_2973,N_2617,N_2770);
or U2974 (N_2974,N_2729,N_2746);
nand U2975 (N_2975,N_2741,N_2612);
or U2976 (N_2976,N_2723,N_2797);
nor U2977 (N_2977,N_2677,N_2600);
and U2978 (N_2978,N_2745,N_2644);
and U2979 (N_2979,N_2741,N_2795);
nand U2980 (N_2980,N_2775,N_2665);
and U2981 (N_2981,N_2602,N_2717);
or U2982 (N_2982,N_2614,N_2609);
nand U2983 (N_2983,N_2619,N_2609);
nand U2984 (N_2984,N_2635,N_2790);
xnor U2985 (N_2985,N_2621,N_2671);
nand U2986 (N_2986,N_2621,N_2607);
or U2987 (N_2987,N_2703,N_2610);
nor U2988 (N_2988,N_2723,N_2719);
nor U2989 (N_2989,N_2705,N_2753);
xnor U2990 (N_2990,N_2687,N_2688);
xnor U2991 (N_2991,N_2768,N_2731);
nand U2992 (N_2992,N_2681,N_2714);
nand U2993 (N_2993,N_2644,N_2627);
xor U2994 (N_2994,N_2789,N_2778);
nor U2995 (N_2995,N_2622,N_2709);
nand U2996 (N_2996,N_2717,N_2691);
or U2997 (N_2997,N_2653,N_2697);
nand U2998 (N_2998,N_2775,N_2757);
xor U2999 (N_2999,N_2792,N_2669);
xor U3000 (N_3000,N_2909,N_2876);
and U3001 (N_3001,N_2962,N_2916);
xnor U3002 (N_3002,N_2813,N_2931);
nand U3003 (N_3003,N_2827,N_2957);
nand U3004 (N_3004,N_2851,N_2852);
or U3005 (N_3005,N_2988,N_2854);
or U3006 (N_3006,N_2881,N_2999);
and U3007 (N_3007,N_2867,N_2899);
nand U3008 (N_3008,N_2950,N_2858);
nor U3009 (N_3009,N_2823,N_2966);
or U3010 (N_3010,N_2947,N_2832);
xor U3011 (N_3011,N_2904,N_2803);
nand U3012 (N_3012,N_2976,N_2846);
and U3013 (N_3013,N_2898,N_2971);
or U3014 (N_3014,N_2840,N_2831);
nor U3015 (N_3015,N_2958,N_2952);
and U3016 (N_3016,N_2835,N_2834);
and U3017 (N_3017,N_2955,N_2839);
nand U3018 (N_3018,N_2896,N_2942);
nor U3019 (N_3019,N_2856,N_2812);
nor U3020 (N_3020,N_2990,N_2845);
nand U3021 (N_3021,N_2948,N_2900);
or U3022 (N_3022,N_2967,N_2818);
nor U3023 (N_3023,N_2871,N_2833);
nor U3024 (N_3024,N_2883,N_2953);
or U3025 (N_3025,N_2879,N_2903);
and U3026 (N_3026,N_2945,N_2930);
nor U3027 (N_3027,N_2933,N_2862);
or U3028 (N_3028,N_2907,N_2892);
xnor U3029 (N_3029,N_2857,N_2875);
xnor U3030 (N_3030,N_2848,N_2984);
nand U3031 (N_3031,N_2949,N_2960);
xnor U3032 (N_3032,N_2995,N_2913);
xnor U3033 (N_3033,N_2925,N_2901);
nor U3034 (N_3034,N_2937,N_2894);
or U3035 (N_3035,N_2959,N_2932);
and U3036 (N_3036,N_2998,N_2935);
nor U3037 (N_3037,N_2979,N_2927);
or U3038 (N_3038,N_2843,N_2910);
nor U3039 (N_3039,N_2895,N_2810);
and U3040 (N_3040,N_2954,N_2946);
nor U3041 (N_3041,N_2880,N_2873);
xnor U3042 (N_3042,N_2970,N_2822);
nand U3043 (N_3043,N_2987,N_2837);
xor U3044 (N_3044,N_2824,N_2817);
and U3045 (N_3045,N_2847,N_2978);
or U3046 (N_3046,N_2980,N_2921);
xnor U3047 (N_3047,N_2819,N_2826);
nor U3048 (N_3048,N_2997,N_2868);
nor U3049 (N_3049,N_2864,N_2891);
nor U3050 (N_3050,N_2986,N_2943);
nand U3051 (N_3051,N_2882,N_2866);
or U3052 (N_3052,N_2929,N_2956);
xor U3053 (N_3053,N_2815,N_2830);
nand U3054 (N_3054,N_2924,N_2825);
or U3055 (N_3055,N_2884,N_2805);
nor U3056 (N_3056,N_2939,N_2861);
nor U3057 (N_3057,N_2992,N_2806);
or U3058 (N_3058,N_2961,N_2915);
and U3059 (N_3059,N_2991,N_2897);
xor U3060 (N_3060,N_2841,N_2938);
or U3061 (N_3061,N_2985,N_2968);
xor U3062 (N_3062,N_2919,N_2829);
xnor U3063 (N_3063,N_2863,N_2923);
xnor U3064 (N_3064,N_2936,N_2972);
xor U3065 (N_3065,N_2885,N_2977);
or U3066 (N_3066,N_2941,N_2877);
nand U3067 (N_3067,N_2888,N_2874);
xnor U3068 (N_3068,N_2905,N_2911);
and U3069 (N_3069,N_2902,N_2940);
xor U3070 (N_3070,N_2965,N_2944);
or U3071 (N_3071,N_2994,N_2973);
nor U3072 (N_3072,N_2842,N_2807);
and U3073 (N_3073,N_2820,N_2993);
xor U3074 (N_3074,N_2872,N_2914);
nand U3075 (N_3075,N_2850,N_2975);
nor U3076 (N_3076,N_2926,N_2918);
nand U3077 (N_3077,N_2969,N_2983);
nor U3078 (N_3078,N_2838,N_2853);
nand U3079 (N_3079,N_2928,N_2982);
xor U3080 (N_3080,N_2800,N_2814);
nand U3081 (N_3081,N_2855,N_2844);
nand U3082 (N_3082,N_2934,N_2878);
nor U3083 (N_3083,N_2922,N_2836);
and U3084 (N_3084,N_2828,N_2917);
nor U3085 (N_3085,N_2865,N_2893);
nand U3086 (N_3086,N_2974,N_2912);
xor U3087 (N_3087,N_2951,N_2886);
nand U3088 (N_3088,N_2809,N_2869);
or U3089 (N_3089,N_2808,N_2908);
nor U3090 (N_3090,N_2996,N_2889);
nand U3091 (N_3091,N_2964,N_2802);
xnor U3092 (N_3092,N_2801,N_2811);
nor U3093 (N_3093,N_2816,N_2906);
or U3094 (N_3094,N_2887,N_2920);
nor U3095 (N_3095,N_2963,N_2859);
nor U3096 (N_3096,N_2821,N_2890);
and U3097 (N_3097,N_2981,N_2989);
or U3098 (N_3098,N_2804,N_2870);
nor U3099 (N_3099,N_2860,N_2849);
and U3100 (N_3100,N_2845,N_2897);
and U3101 (N_3101,N_2908,N_2911);
or U3102 (N_3102,N_2940,N_2805);
nand U3103 (N_3103,N_2978,N_2892);
nand U3104 (N_3104,N_2897,N_2912);
and U3105 (N_3105,N_2849,N_2829);
xor U3106 (N_3106,N_2958,N_2975);
or U3107 (N_3107,N_2833,N_2956);
and U3108 (N_3108,N_2850,N_2885);
or U3109 (N_3109,N_2838,N_2873);
and U3110 (N_3110,N_2942,N_2980);
nand U3111 (N_3111,N_2822,N_2881);
or U3112 (N_3112,N_2810,N_2899);
xnor U3113 (N_3113,N_2966,N_2852);
or U3114 (N_3114,N_2830,N_2978);
or U3115 (N_3115,N_2854,N_2945);
nor U3116 (N_3116,N_2900,N_2925);
or U3117 (N_3117,N_2842,N_2893);
nor U3118 (N_3118,N_2867,N_2884);
nand U3119 (N_3119,N_2958,N_2907);
xnor U3120 (N_3120,N_2982,N_2976);
or U3121 (N_3121,N_2975,N_2910);
and U3122 (N_3122,N_2961,N_2856);
xnor U3123 (N_3123,N_2908,N_2896);
nand U3124 (N_3124,N_2891,N_2955);
nand U3125 (N_3125,N_2999,N_2937);
nor U3126 (N_3126,N_2818,N_2974);
xor U3127 (N_3127,N_2946,N_2956);
nor U3128 (N_3128,N_2979,N_2896);
xor U3129 (N_3129,N_2829,N_2857);
nor U3130 (N_3130,N_2801,N_2938);
or U3131 (N_3131,N_2899,N_2932);
nor U3132 (N_3132,N_2827,N_2833);
and U3133 (N_3133,N_2863,N_2854);
nand U3134 (N_3134,N_2899,N_2826);
or U3135 (N_3135,N_2928,N_2915);
nor U3136 (N_3136,N_2910,N_2832);
nor U3137 (N_3137,N_2905,N_2938);
xnor U3138 (N_3138,N_2991,N_2988);
or U3139 (N_3139,N_2816,N_2825);
xor U3140 (N_3140,N_2843,N_2831);
nand U3141 (N_3141,N_2807,N_2981);
or U3142 (N_3142,N_2973,N_2970);
or U3143 (N_3143,N_2835,N_2965);
xnor U3144 (N_3144,N_2924,N_2916);
and U3145 (N_3145,N_2997,N_2938);
nor U3146 (N_3146,N_2909,N_2963);
nand U3147 (N_3147,N_2814,N_2867);
nor U3148 (N_3148,N_2869,N_2802);
xor U3149 (N_3149,N_2877,N_2859);
or U3150 (N_3150,N_2868,N_2825);
nand U3151 (N_3151,N_2864,N_2975);
xnor U3152 (N_3152,N_2841,N_2981);
nor U3153 (N_3153,N_2864,N_2840);
nand U3154 (N_3154,N_2911,N_2819);
xor U3155 (N_3155,N_2908,N_2974);
and U3156 (N_3156,N_2881,N_2810);
nor U3157 (N_3157,N_2823,N_2820);
xnor U3158 (N_3158,N_2978,N_2855);
nand U3159 (N_3159,N_2934,N_2827);
xor U3160 (N_3160,N_2847,N_2919);
nor U3161 (N_3161,N_2935,N_2954);
or U3162 (N_3162,N_2900,N_2919);
xor U3163 (N_3163,N_2820,N_2950);
nand U3164 (N_3164,N_2910,N_2969);
or U3165 (N_3165,N_2844,N_2908);
xor U3166 (N_3166,N_2893,N_2926);
and U3167 (N_3167,N_2964,N_2852);
nand U3168 (N_3168,N_2950,N_2915);
xnor U3169 (N_3169,N_2906,N_2827);
nand U3170 (N_3170,N_2829,N_2940);
and U3171 (N_3171,N_2836,N_2941);
nor U3172 (N_3172,N_2838,N_2875);
xor U3173 (N_3173,N_2805,N_2933);
or U3174 (N_3174,N_2948,N_2889);
xnor U3175 (N_3175,N_2963,N_2896);
and U3176 (N_3176,N_2950,N_2844);
or U3177 (N_3177,N_2859,N_2990);
or U3178 (N_3178,N_2961,N_2868);
or U3179 (N_3179,N_2935,N_2914);
nor U3180 (N_3180,N_2940,N_2815);
and U3181 (N_3181,N_2974,N_2988);
xor U3182 (N_3182,N_2853,N_2855);
xnor U3183 (N_3183,N_2850,N_2962);
xor U3184 (N_3184,N_2896,N_2922);
nand U3185 (N_3185,N_2871,N_2805);
xor U3186 (N_3186,N_2806,N_2901);
nand U3187 (N_3187,N_2839,N_2968);
xor U3188 (N_3188,N_2830,N_2967);
nand U3189 (N_3189,N_2916,N_2931);
nor U3190 (N_3190,N_2896,N_2969);
xor U3191 (N_3191,N_2920,N_2878);
nand U3192 (N_3192,N_2830,N_2820);
nor U3193 (N_3193,N_2955,N_2919);
nor U3194 (N_3194,N_2951,N_2885);
xnor U3195 (N_3195,N_2903,N_2828);
and U3196 (N_3196,N_2869,N_2828);
and U3197 (N_3197,N_2862,N_2809);
or U3198 (N_3198,N_2888,N_2895);
nand U3199 (N_3199,N_2964,N_2922);
nand U3200 (N_3200,N_3098,N_3169);
or U3201 (N_3201,N_3097,N_3008);
and U3202 (N_3202,N_3114,N_3153);
nand U3203 (N_3203,N_3035,N_3156);
and U3204 (N_3204,N_3082,N_3023);
nand U3205 (N_3205,N_3150,N_3083);
and U3206 (N_3206,N_3044,N_3089);
and U3207 (N_3207,N_3032,N_3055);
or U3208 (N_3208,N_3028,N_3104);
nor U3209 (N_3209,N_3136,N_3030);
nor U3210 (N_3210,N_3056,N_3096);
xnor U3211 (N_3211,N_3140,N_3046);
and U3212 (N_3212,N_3119,N_3170);
nand U3213 (N_3213,N_3086,N_3011);
xnor U3214 (N_3214,N_3027,N_3058);
xor U3215 (N_3215,N_3163,N_3190);
nand U3216 (N_3216,N_3176,N_3193);
nor U3217 (N_3217,N_3021,N_3135);
nand U3218 (N_3218,N_3101,N_3080);
or U3219 (N_3219,N_3192,N_3103);
nor U3220 (N_3220,N_3145,N_3014);
and U3221 (N_3221,N_3100,N_3185);
xor U3222 (N_3222,N_3149,N_3079);
nand U3223 (N_3223,N_3078,N_3129);
and U3224 (N_3224,N_3117,N_3039);
nor U3225 (N_3225,N_3189,N_3178);
nand U3226 (N_3226,N_3105,N_3041);
or U3227 (N_3227,N_3053,N_3102);
nand U3228 (N_3228,N_3075,N_3141);
xnor U3229 (N_3229,N_3123,N_3005);
nand U3230 (N_3230,N_3081,N_3099);
or U3231 (N_3231,N_3088,N_3187);
nor U3232 (N_3232,N_3057,N_3157);
or U3233 (N_3233,N_3191,N_3111);
and U3234 (N_3234,N_3143,N_3165);
nor U3235 (N_3235,N_3184,N_3073);
or U3236 (N_3236,N_3132,N_3049);
xnor U3237 (N_3237,N_3077,N_3125);
xor U3238 (N_3238,N_3188,N_3133);
or U3239 (N_3239,N_3183,N_3009);
nor U3240 (N_3240,N_3012,N_3148);
nor U3241 (N_3241,N_3107,N_3002);
and U3242 (N_3242,N_3066,N_3164);
nor U3243 (N_3243,N_3061,N_3019);
and U3244 (N_3244,N_3121,N_3158);
xnor U3245 (N_3245,N_3122,N_3162);
or U3246 (N_3246,N_3142,N_3174);
nor U3247 (N_3247,N_3040,N_3043);
nor U3248 (N_3248,N_3197,N_3171);
or U3249 (N_3249,N_3167,N_3137);
xnor U3250 (N_3250,N_3024,N_3139);
xnor U3251 (N_3251,N_3175,N_3004);
or U3252 (N_3252,N_3147,N_3177);
or U3253 (N_3253,N_3180,N_3144);
and U3254 (N_3254,N_3025,N_3070);
and U3255 (N_3255,N_3069,N_3045);
xnor U3256 (N_3256,N_3050,N_3003);
nor U3257 (N_3257,N_3036,N_3076);
or U3258 (N_3258,N_3060,N_3010);
xnor U3259 (N_3259,N_3116,N_3013);
or U3260 (N_3260,N_3064,N_3092);
nand U3261 (N_3261,N_3186,N_3034);
nor U3262 (N_3262,N_3062,N_3026);
xor U3263 (N_3263,N_3154,N_3196);
nand U3264 (N_3264,N_3068,N_3128);
nand U3265 (N_3265,N_3106,N_3160);
or U3266 (N_3266,N_3020,N_3047);
nand U3267 (N_3267,N_3130,N_3052);
xnor U3268 (N_3268,N_3090,N_3195);
nor U3269 (N_3269,N_3048,N_3168);
or U3270 (N_3270,N_3094,N_3109);
nor U3271 (N_3271,N_3059,N_3072);
nand U3272 (N_3272,N_3134,N_3006);
xor U3273 (N_3273,N_3110,N_3085);
xor U3274 (N_3274,N_3087,N_3198);
xor U3275 (N_3275,N_3112,N_3131);
and U3276 (N_3276,N_3029,N_3007);
or U3277 (N_3277,N_3001,N_3182);
xor U3278 (N_3278,N_3074,N_3152);
nand U3279 (N_3279,N_3018,N_3091);
nor U3280 (N_3280,N_3000,N_3146);
xnor U3281 (N_3281,N_3161,N_3038);
nand U3282 (N_3282,N_3016,N_3194);
xnor U3283 (N_3283,N_3063,N_3033);
and U3284 (N_3284,N_3022,N_3118);
nand U3285 (N_3285,N_3124,N_3173);
xnor U3286 (N_3286,N_3095,N_3199);
and U3287 (N_3287,N_3108,N_3054);
xnor U3288 (N_3288,N_3093,N_3127);
nand U3289 (N_3289,N_3067,N_3120);
nor U3290 (N_3290,N_3151,N_3015);
xor U3291 (N_3291,N_3179,N_3065);
nor U3292 (N_3292,N_3037,N_3071);
or U3293 (N_3293,N_3084,N_3155);
nor U3294 (N_3294,N_3172,N_3181);
and U3295 (N_3295,N_3113,N_3031);
xor U3296 (N_3296,N_3138,N_3126);
nand U3297 (N_3297,N_3051,N_3166);
nor U3298 (N_3298,N_3042,N_3017);
nor U3299 (N_3299,N_3159,N_3115);
and U3300 (N_3300,N_3054,N_3113);
or U3301 (N_3301,N_3077,N_3161);
or U3302 (N_3302,N_3125,N_3054);
or U3303 (N_3303,N_3021,N_3001);
and U3304 (N_3304,N_3072,N_3079);
and U3305 (N_3305,N_3079,N_3159);
or U3306 (N_3306,N_3007,N_3120);
xor U3307 (N_3307,N_3096,N_3128);
or U3308 (N_3308,N_3059,N_3106);
or U3309 (N_3309,N_3126,N_3010);
nand U3310 (N_3310,N_3171,N_3085);
nand U3311 (N_3311,N_3103,N_3186);
nor U3312 (N_3312,N_3054,N_3182);
xor U3313 (N_3313,N_3085,N_3176);
nor U3314 (N_3314,N_3177,N_3009);
nor U3315 (N_3315,N_3059,N_3001);
xnor U3316 (N_3316,N_3197,N_3138);
nand U3317 (N_3317,N_3192,N_3017);
and U3318 (N_3318,N_3144,N_3172);
nand U3319 (N_3319,N_3023,N_3056);
or U3320 (N_3320,N_3191,N_3104);
nand U3321 (N_3321,N_3061,N_3073);
xnor U3322 (N_3322,N_3122,N_3102);
and U3323 (N_3323,N_3036,N_3012);
nand U3324 (N_3324,N_3151,N_3145);
xnor U3325 (N_3325,N_3006,N_3103);
xor U3326 (N_3326,N_3189,N_3057);
nor U3327 (N_3327,N_3077,N_3043);
nor U3328 (N_3328,N_3179,N_3182);
nor U3329 (N_3329,N_3021,N_3038);
nand U3330 (N_3330,N_3100,N_3124);
and U3331 (N_3331,N_3169,N_3189);
nor U3332 (N_3332,N_3153,N_3090);
nand U3333 (N_3333,N_3092,N_3152);
nand U3334 (N_3334,N_3005,N_3136);
nand U3335 (N_3335,N_3015,N_3033);
nand U3336 (N_3336,N_3126,N_3090);
xor U3337 (N_3337,N_3121,N_3096);
or U3338 (N_3338,N_3032,N_3122);
nor U3339 (N_3339,N_3106,N_3007);
xnor U3340 (N_3340,N_3110,N_3045);
nand U3341 (N_3341,N_3098,N_3007);
nand U3342 (N_3342,N_3010,N_3018);
and U3343 (N_3343,N_3124,N_3014);
nor U3344 (N_3344,N_3199,N_3144);
xor U3345 (N_3345,N_3000,N_3178);
or U3346 (N_3346,N_3143,N_3167);
nor U3347 (N_3347,N_3090,N_3161);
nand U3348 (N_3348,N_3134,N_3129);
xnor U3349 (N_3349,N_3187,N_3085);
or U3350 (N_3350,N_3022,N_3062);
nand U3351 (N_3351,N_3049,N_3158);
xor U3352 (N_3352,N_3112,N_3031);
xor U3353 (N_3353,N_3148,N_3069);
nand U3354 (N_3354,N_3192,N_3037);
xnor U3355 (N_3355,N_3130,N_3008);
or U3356 (N_3356,N_3122,N_3134);
and U3357 (N_3357,N_3164,N_3050);
or U3358 (N_3358,N_3017,N_3145);
and U3359 (N_3359,N_3158,N_3169);
xnor U3360 (N_3360,N_3095,N_3001);
and U3361 (N_3361,N_3127,N_3148);
nand U3362 (N_3362,N_3028,N_3003);
and U3363 (N_3363,N_3156,N_3180);
nand U3364 (N_3364,N_3186,N_3080);
and U3365 (N_3365,N_3148,N_3160);
and U3366 (N_3366,N_3005,N_3035);
and U3367 (N_3367,N_3018,N_3118);
nand U3368 (N_3368,N_3005,N_3019);
and U3369 (N_3369,N_3164,N_3128);
xnor U3370 (N_3370,N_3122,N_3002);
nor U3371 (N_3371,N_3011,N_3052);
nor U3372 (N_3372,N_3128,N_3011);
nor U3373 (N_3373,N_3197,N_3193);
or U3374 (N_3374,N_3113,N_3175);
and U3375 (N_3375,N_3137,N_3155);
and U3376 (N_3376,N_3037,N_3119);
and U3377 (N_3377,N_3126,N_3062);
nand U3378 (N_3378,N_3108,N_3178);
nor U3379 (N_3379,N_3146,N_3150);
xnor U3380 (N_3380,N_3129,N_3018);
nor U3381 (N_3381,N_3062,N_3131);
and U3382 (N_3382,N_3015,N_3093);
xnor U3383 (N_3383,N_3186,N_3167);
and U3384 (N_3384,N_3090,N_3167);
nand U3385 (N_3385,N_3148,N_3075);
xnor U3386 (N_3386,N_3102,N_3064);
and U3387 (N_3387,N_3139,N_3175);
xnor U3388 (N_3388,N_3102,N_3116);
xor U3389 (N_3389,N_3038,N_3184);
or U3390 (N_3390,N_3031,N_3186);
or U3391 (N_3391,N_3174,N_3018);
and U3392 (N_3392,N_3025,N_3162);
or U3393 (N_3393,N_3190,N_3092);
xor U3394 (N_3394,N_3079,N_3182);
nor U3395 (N_3395,N_3136,N_3163);
or U3396 (N_3396,N_3139,N_3134);
nor U3397 (N_3397,N_3022,N_3196);
xor U3398 (N_3398,N_3146,N_3190);
or U3399 (N_3399,N_3112,N_3037);
nor U3400 (N_3400,N_3389,N_3242);
nor U3401 (N_3401,N_3273,N_3327);
nand U3402 (N_3402,N_3299,N_3343);
xor U3403 (N_3403,N_3349,N_3254);
and U3404 (N_3404,N_3325,N_3376);
nand U3405 (N_3405,N_3338,N_3229);
xor U3406 (N_3406,N_3388,N_3214);
nor U3407 (N_3407,N_3352,N_3390);
nor U3408 (N_3408,N_3257,N_3233);
or U3409 (N_3409,N_3313,N_3228);
and U3410 (N_3410,N_3385,N_3329);
or U3411 (N_3411,N_3356,N_3206);
xnor U3412 (N_3412,N_3275,N_3235);
nor U3413 (N_3413,N_3296,N_3317);
or U3414 (N_3414,N_3239,N_3305);
or U3415 (N_3415,N_3282,N_3341);
nor U3416 (N_3416,N_3201,N_3223);
xnor U3417 (N_3417,N_3397,N_3374);
or U3418 (N_3418,N_3297,N_3365);
xnor U3419 (N_3419,N_3340,N_3219);
xor U3420 (N_3420,N_3298,N_3210);
xor U3421 (N_3421,N_3240,N_3392);
or U3422 (N_3422,N_3360,N_3333);
and U3423 (N_3423,N_3256,N_3301);
nand U3424 (N_3424,N_3372,N_3344);
or U3425 (N_3425,N_3217,N_3270);
and U3426 (N_3426,N_3318,N_3363);
nor U3427 (N_3427,N_3276,N_3312);
nand U3428 (N_3428,N_3287,N_3267);
nor U3429 (N_3429,N_3322,N_3227);
and U3430 (N_3430,N_3308,N_3319);
or U3431 (N_3431,N_3260,N_3358);
nor U3432 (N_3432,N_3336,N_3247);
or U3433 (N_3433,N_3387,N_3359);
and U3434 (N_3434,N_3354,N_3241);
and U3435 (N_3435,N_3357,N_3248);
and U3436 (N_3436,N_3268,N_3218);
nor U3437 (N_3437,N_3335,N_3203);
and U3438 (N_3438,N_3394,N_3249);
nor U3439 (N_3439,N_3259,N_3367);
and U3440 (N_3440,N_3232,N_3253);
and U3441 (N_3441,N_3368,N_3314);
xor U3442 (N_3442,N_3245,N_3280);
xor U3443 (N_3443,N_3293,N_3212);
xnor U3444 (N_3444,N_3309,N_3290);
nand U3445 (N_3445,N_3291,N_3252);
nand U3446 (N_3446,N_3382,N_3320);
or U3447 (N_3447,N_3220,N_3284);
nor U3448 (N_3448,N_3215,N_3236);
and U3449 (N_3449,N_3213,N_3264);
and U3450 (N_3450,N_3364,N_3351);
and U3451 (N_3451,N_3378,N_3216);
nand U3452 (N_3452,N_3353,N_3304);
or U3453 (N_3453,N_3208,N_3251);
or U3454 (N_3454,N_3209,N_3258);
nand U3455 (N_3455,N_3226,N_3285);
and U3456 (N_3456,N_3279,N_3274);
nor U3457 (N_3457,N_3377,N_3277);
and U3458 (N_3458,N_3332,N_3316);
and U3459 (N_3459,N_3345,N_3288);
or U3460 (N_3460,N_3234,N_3255);
and U3461 (N_3461,N_3399,N_3231);
or U3462 (N_3462,N_3391,N_3261);
or U3463 (N_3463,N_3361,N_3211);
or U3464 (N_3464,N_3283,N_3339);
or U3465 (N_3465,N_3225,N_3230);
or U3466 (N_3466,N_3331,N_3295);
nand U3467 (N_3467,N_3315,N_3263);
nor U3468 (N_3468,N_3265,N_3386);
xor U3469 (N_3469,N_3222,N_3266);
or U3470 (N_3470,N_3200,N_3307);
and U3471 (N_3471,N_3396,N_3362);
nand U3472 (N_3472,N_3334,N_3292);
and U3473 (N_3473,N_3224,N_3347);
xnor U3474 (N_3474,N_3381,N_3379);
nor U3475 (N_3475,N_3237,N_3286);
or U3476 (N_3476,N_3348,N_3207);
or U3477 (N_3477,N_3269,N_3337);
and U3478 (N_3478,N_3346,N_3369);
xnor U3479 (N_3479,N_3324,N_3205);
xor U3480 (N_3480,N_3272,N_3294);
and U3481 (N_3481,N_3375,N_3321);
nor U3482 (N_3482,N_3373,N_3243);
nand U3483 (N_3483,N_3202,N_3383);
nand U3484 (N_3484,N_3278,N_3326);
nand U3485 (N_3485,N_3366,N_3330);
xor U3486 (N_3486,N_3328,N_3323);
nor U3487 (N_3487,N_3289,N_3204);
nor U3488 (N_3488,N_3302,N_3303);
or U3489 (N_3489,N_3244,N_3371);
or U3490 (N_3490,N_3395,N_3262);
nor U3491 (N_3491,N_3355,N_3380);
or U3492 (N_3492,N_3271,N_3250);
nand U3493 (N_3493,N_3384,N_3281);
nor U3494 (N_3494,N_3238,N_3393);
and U3495 (N_3495,N_3306,N_3342);
nor U3496 (N_3496,N_3300,N_3311);
nor U3497 (N_3497,N_3310,N_3350);
nand U3498 (N_3498,N_3221,N_3370);
or U3499 (N_3499,N_3246,N_3398);
nand U3500 (N_3500,N_3358,N_3246);
and U3501 (N_3501,N_3271,N_3386);
nor U3502 (N_3502,N_3270,N_3324);
and U3503 (N_3503,N_3275,N_3294);
xor U3504 (N_3504,N_3351,N_3224);
nand U3505 (N_3505,N_3247,N_3258);
nor U3506 (N_3506,N_3287,N_3248);
nand U3507 (N_3507,N_3379,N_3243);
xor U3508 (N_3508,N_3224,N_3287);
or U3509 (N_3509,N_3309,N_3251);
nand U3510 (N_3510,N_3210,N_3244);
nor U3511 (N_3511,N_3393,N_3204);
nor U3512 (N_3512,N_3311,N_3301);
nand U3513 (N_3513,N_3371,N_3364);
nand U3514 (N_3514,N_3207,N_3220);
and U3515 (N_3515,N_3233,N_3321);
and U3516 (N_3516,N_3257,N_3303);
xnor U3517 (N_3517,N_3367,N_3269);
or U3518 (N_3518,N_3306,N_3265);
nor U3519 (N_3519,N_3287,N_3368);
and U3520 (N_3520,N_3258,N_3300);
and U3521 (N_3521,N_3382,N_3343);
and U3522 (N_3522,N_3312,N_3225);
and U3523 (N_3523,N_3283,N_3243);
or U3524 (N_3524,N_3345,N_3252);
nand U3525 (N_3525,N_3265,N_3267);
and U3526 (N_3526,N_3254,N_3308);
and U3527 (N_3527,N_3292,N_3392);
or U3528 (N_3528,N_3230,N_3367);
xnor U3529 (N_3529,N_3390,N_3267);
nand U3530 (N_3530,N_3210,N_3326);
nor U3531 (N_3531,N_3210,N_3384);
xor U3532 (N_3532,N_3387,N_3208);
xor U3533 (N_3533,N_3261,N_3316);
nand U3534 (N_3534,N_3335,N_3209);
or U3535 (N_3535,N_3241,N_3337);
or U3536 (N_3536,N_3329,N_3388);
xnor U3537 (N_3537,N_3224,N_3312);
or U3538 (N_3538,N_3381,N_3254);
nor U3539 (N_3539,N_3300,N_3367);
nand U3540 (N_3540,N_3228,N_3305);
and U3541 (N_3541,N_3316,N_3287);
nand U3542 (N_3542,N_3357,N_3322);
or U3543 (N_3543,N_3359,N_3300);
nand U3544 (N_3544,N_3327,N_3346);
nand U3545 (N_3545,N_3395,N_3274);
or U3546 (N_3546,N_3231,N_3296);
and U3547 (N_3547,N_3394,N_3379);
nor U3548 (N_3548,N_3325,N_3309);
or U3549 (N_3549,N_3249,N_3259);
xnor U3550 (N_3550,N_3271,N_3354);
and U3551 (N_3551,N_3298,N_3208);
and U3552 (N_3552,N_3207,N_3294);
xor U3553 (N_3553,N_3326,N_3364);
nor U3554 (N_3554,N_3216,N_3392);
or U3555 (N_3555,N_3348,N_3250);
xor U3556 (N_3556,N_3260,N_3270);
xnor U3557 (N_3557,N_3270,N_3395);
xor U3558 (N_3558,N_3230,N_3208);
and U3559 (N_3559,N_3303,N_3310);
nand U3560 (N_3560,N_3342,N_3292);
or U3561 (N_3561,N_3228,N_3312);
nand U3562 (N_3562,N_3312,N_3202);
xor U3563 (N_3563,N_3256,N_3285);
xnor U3564 (N_3564,N_3254,N_3279);
nand U3565 (N_3565,N_3255,N_3335);
nand U3566 (N_3566,N_3266,N_3215);
nor U3567 (N_3567,N_3336,N_3318);
or U3568 (N_3568,N_3287,N_3347);
nand U3569 (N_3569,N_3327,N_3229);
xnor U3570 (N_3570,N_3238,N_3380);
nor U3571 (N_3571,N_3336,N_3397);
nand U3572 (N_3572,N_3339,N_3266);
nor U3573 (N_3573,N_3360,N_3366);
or U3574 (N_3574,N_3206,N_3284);
xor U3575 (N_3575,N_3239,N_3312);
and U3576 (N_3576,N_3251,N_3283);
xnor U3577 (N_3577,N_3344,N_3245);
nand U3578 (N_3578,N_3349,N_3226);
nand U3579 (N_3579,N_3355,N_3217);
and U3580 (N_3580,N_3307,N_3277);
or U3581 (N_3581,N_3298,N_3367);
and U3582 (N_3582,N_3249,N_3201);
xor U3583 (N_3583,N_3269,N_3333);
and U3584 (N_3584,N_3292,N_3397);
or U3585 (N_3585,N_3374,N_3394);
and U3586 (N_3586,N_3273,N_3221);
or U3587 (N_3587,N_3398,N_3365);
and U3588 (N_3588,N_3383,N_3200);
xnor U3589 (N_3589,N_3241,N_3298);
nand U3590 (N_3590,N_3347,N_3383);
and U3591 (N_3591,N_3386,N_3325);
xor U3592 (N_3592,N_3203,N_3228);
or U3593 (N_3593,N_3398,N_3298);
or U3594 (N_3594,N_3335,N_3201);
and U3595 (N_3595,N_3299,N_3230);
and U3596 (N_3596,N_3266,N_3350);
or U3597 (N_3597,N_3264,N_3311);
nor U3598 (N_3598,N_3336,N_3352);
nand U3599 (N_3599,N_3341,N_3229);
and U3600 (N_3600,N_3486,N_3493);
nor U3601 (N_3601,N_3522,N_3548);
or U3602 (N_3602,N_3440,N_3477);
xor U3603 (N_3603,N_3457,N_3588);
xnor U3604 (N_3604,N_3451,N_3545);
nor U3605 (N_3605,N_3501,N_3557);
nand U3606 (N_3606,N_3469,N_3584);
xor U3607 (N_3607,N_3455,N_3491);
nor U3608 (N_3608,N_3526,N_3555);
xor U3609 (N_3609,N_3485,N_3513);
nor U3610 (N_3610,N_3506,N_3434);
nor U3611 (N_3611,N_3516,N_3567);
xnor U3612 (N_3612,N_3468,N_3420);
or U3613 (N_3613,N_3542,N_3412);
nand U3614 (N_3614,N_3497,N_3479);
xnor U3615 (N_3615,N_3456,N_3424);
or U3616 (N_3616,N_3460,N_3443);
nand U3617 (N_3617,N_3494,N_3461);
nor U3618 (N_3618,N_3464,N_3599);
or U3619 (N_3619,N_3484,N_3425);
nand U3620 (N_3620,N_3439,N_3546);
or U3621 (N_3621,N_3541,N_3419);
nand U3622 (N_3622,N_3589,N_3467);
and U3623 (N_3623,N_3433,N_3598);
or U3624 (N_3624,N_3438,N_3561);
xor U3625 (N_3625,N_3530,N_3437);
xor U3626 (N_3626,N_3576,N_3404);
xnor U3627 (N_3627,N_3577,N_3586);
and U3628 (N_3628,N_3532,N_3511);
xnor U3629 (N_3629,N_3518,N_3524);
xnor U3630 (N_3630,N_3538,N_3582);
or U3631 (N_3631,N_3475,N_3558);
nand U3632 (N_3632,N_3591,N_3566);
and U3633 (N_3633,N_3432,N_3495);
xnor U3634 (N_3634,N_3595,N_3521);
or U3635 (N_3635,N_3590,N_3596);
nand U3636 (N_3636,N_3471,N_3431);
and U3637 (N_3637,N_3403,N_3459);
nor U3638 (N_3638,N_3565,N_3447);
and U3639 (N_3639,N_3579,N_3527);
nor U3640 (N_3640,N_3406,N_3429);
nand U3641 (N_3641,N_3413,N_3448);
or U3642 (N_3642,N_3593,N_3427);
and U3643 (N_3643,N_3507,N_3481);
nand U3644 (N_3644,N_3517,N_3415);
and U3645 (N_3645,N_3523,N_3550);
and U3646 (N_3646,N_3492,N_3552);
nand U3647 (N_3647,N_3504,N_3417);
or U3648 (N_3648,N_3587,N_3408);
xor U3649 (N_3649,N_3500,N_3400);
xnor U3650 (N_3650,N_3410,N_3533);
and U3651 (N_3651,N_3428,N_3496);
nand U3652 (N_3652,N_3580,N_3583);
nand U3653 (N_3653,N_3462,N_3449);
and U3654 (N_3654,N_3515,N_3536);
and U3655 (N_3655,N_3525,N_3594);
xor U3656 (N_3656,N_3421,N_3528);
nand U3657 (N_3657,N_3411,N_3592);
nor U3658 (N_3658,N_3529,N_3559);
and U3659 (N_3659,N_3564,N_3444);
xor U3660 (N_3660,N_3482,N_3418);
xnor U3661 (N_3661,N_3499,N_3409);
or U3662 (N_3662,N_3597,N_3514);
and U3663 (N_3663,N_3436,N_3551);
nand U3664 (N_3664,N_3537,N_3474);
or U3665 (N_3665,N_3407,N_3535);
xnor U3666 (N_3666,N_3543,N_3480);
or U3667 (N_3667,N_3571,N_3458);
and U3668 (N_3668,N_3473,N_3476);
xnor U3669 (N_3669,N_3503,N_3569);
or U3670 (N_3670,N_3470,N_3401);
nand U3671 (N_3671,N_3405,N_3423);
and U3672 (N_3672,N_3453,N_3553);
xnor U3673 (N_3673,N_3573,N_3442);
and U3674 (N_3674,N_3512,N_3572);
nand U3675 (N_3675,N_3450,N_3563);
and U3676 (N_3676,N_3489,N_3549);
or U3677 (N_3677,N_3560,N_3416);
or U3678 (N_3678,N_3472,N_3547);
xor U3679 (N_3679,N_3556,N_3466);
nand U3680 (N_3680,N_3465,N_3570);
or U3681 (N_3681,N_3446,N_3488);
or U3682 (N_3682,N_3509,N_3441);
or U3683 (N_3683,N_3510,N_3575);
and U3684 (N_3684,N_3463,N_3519);
xor U3685 (N_3685,N_3581,N_3478);
nor U3686 (N_3686,N_3531,N_3578);
and U3687 (N_3687,N_3487,N_3445);
or U3688 (N_3688,N_3435,N_3554);
and U3689 (N_3689,N_3454,N_3490);
xor U3690 (N_3690,N_3534,N_3498);
and U3691 (N_3691,N_3568,N_3502);
nor U3692 (N_3692,N_3585,N_3574);
or U3693 (N_3693,N_3414,N_3540);
xor U3694 (N_3694,N_3483,N_3505);
or U3695 (N_3695,N_3520,N_3452);
or U3696 (N_3696,N_3426,N_3508);
or U3697 (N_3697,N_3402,N_3562);
or U3698 (N_3698,N_3544,N_3539);
and U3699 (N_3699,N_3422,N_3430);
xnor U3700 (N_3700,N_3580,N_3533);
and U3701 (N_3701,N_3438,N_3529);
nand U3702 (N_3702,N_3465,N_3401);
nand U3703 (N_3703,N_3520,N_3416);
or U3704 (N_3704,N_3565,N_3594);
or U3705 (N_3705,N_3425,N_3429);
nor U3706 (N_3706,N_3495,N_3520);
nor U3707 (N_3707,N_3559,N_3487);
and U3708 (N_3708,N_3584,N_3550);
nand U3709 (N_3709,N_3420,N_3444);
and U3710 (N_3710,N_3431,N_3456);
xnor U3711 (N_3711,N_3512,N_3456);
nor U3712 (N_3712,N_3448,N_3547);
xnor U3713 (N_3713,N_3437,N_3466);
nor U3714 (N_3714,N_3459,N_3568);
nor U3715 (N_3715,N_3559,N_3566);
nor U3716 (N_3716,N_3425,N_3496);
and U3717 (N_3717,N_3452,N_3402);
or U3718 (N_3718,N_3576,N_3555);
xor U3719 (N_3719,N_3473,N_3549);
or U3720 (N_3720,N_3520,N_3516);
and U3721 (N_3721,N_3452,N_3456);
xor U3722 (N_3722,N_3545,N_3462);
xnor U3723 (N_3723,N_3451,N_3555);
xor U3724 (N_3724,N_3490,N_3561);
or U3725 (N_3725,N_3402,N_3547);
nand U3726 (N_3726,N_3497,N_3408);
and U3727 (N_3727,N_3485,N_3561);
xnor U3728 (N_3728,N_3497,N_3460);
nor U3729 (N_3729,N_3462,N_3557);
and U3730 (N_3730,N_3593,N_3466);
and U3731 (N_3731,N_3487,N_3413);
or U3732 (N_3732,N_3564,N_3452);
and U3733 (N_3733,N_3471,N_3545);
nand U3734 (N_3734,N_3531,N_3500);
and U3735 (N_3735,N_3576,N_3456);
nor U3736 (N_3736,N_3495,N_3420);
xor U3737 (N_3737,N_3422,N_3451);
nand U3738 (N_3738,N_3471,N_3597);
and U3739 (N_3739,N_3443,N_3588);
or U3740 (N_3740,N_3591,N_3557);
nand U3741 (N_3741,N_3405,N_3477);
or U3742 (N_3742,N_3491,N_3411);
or U3743 (N_3743,N_3515,N_3522);
or U3744 (N_3744,N_3533,N_3500);
nor U3745 (N_3745,N_3492,N_3554);
or U3746 (N_3746,N_3507,N_3570);
nand U3747 (N_3747,N_3503,N_3483);
xnor U3748 (N_3748,N_3463,N_3593);
and U3749 (N_3749,N_3510,N_3469);
nor U3750 (N_3750,N_3466,N_3526);
nor U3751 (N_3751,N_3423,N_3543);
and U3752 (N_3752,N_3543,N_3448);
nor U3753 (N_3753,N_3540,N_3462);
and U3754 (N_3754,N_3492,N_3413);
nor U3755 (N_3755,N_3514,N_3542);
and U3756 (N_3756,N_3401,N_3543);
nand U3757 (N_3757,N_3497,N_3489);
nand U3758 (N_3758,N_3536,N_3408);
nand U3759 (N_3759,N_3438,N_3410);
nand U3760 (N_3760,N_3476,N_3405);
and U3761 (N_3761,N_3559,N_3415);
xnor U3762 (N_3762,N_3469,N_3578);
or U3763 (N_3763,N_3478,N_3586);
or U3764 (N_3764,N_3514,N_3425);
xor U3765 (N_3765,N_3597,N_3431);
nand U3766 (N_3766,N_3492,N_3407);
and U3767 (N_3767,N_3494,N_3455);
xor U3768 (N_3768,N_3503,N_3529);
nor U3769 (N_3769,N_3553,N_3440);
nor U3770 (N_3770,N_3502,N_3527);
and U3771 (N_3771,N_3445,N_3498);
xor U3772 (N_3772,N_3423,N_3463);
nand U3773 (N_3773,N_3560,N_3516);
nand U3774 (N_3774,N_3419,N_3503);
xor U3775 (N_3775,N_3467,N_3420);
or U3776 (N_3776,N_3440,N_3512);
nand U3777 (N_3777,N_3401,N_3509);
xnor U3778 (N_3778,N_3522,N_3519);
xor U3779 (N_3779,N_3412,N_3575);
or U3780 (N_3780,N_3469,N_3490);
or U3781 (N_3781,N_3504,N_3405);
nand U3782 (N_3782,N_3453,N_3564);
nor U3783 (N_3783,N_3533,N_3532);
xnor U3784 (N_3784,N_3461,N_3437);
xor U3785 (N_3785,N_3598,N_3492);
nor U3786 (N_3786,N_3450,N_3515);
nand U3787 (N_3787,N_3461,N_3430);
and U3788 (N_3788,N_3551,N_3405);
and U3789 (N_3789,N_3483,N_3530);
and U3790 (N_3790,N_3479,N_3553);
nand U3791 (N_3791,N_3465,N_3515);
or U3792 (N_3792,N_3590,N_3568);
nor U3793 (N_3793,N_3507,N_3557);
or U3794 (N_3794,N_3436,N_3580);
and U3795 (N_3795,N_3532,N_3463);
xor U3796 (N_3796,N_3586,N_3481);
and U3797 (N_3797,N_3417,N_3479);
and U3798 (N_3798,N_3566,N_3419);
and U3799 (N_3799,N_3459,N_3542);
nand U3800 (N_3800,N_3790,N_3776);
and U3801 (N_3801,N_3781,N_3784);
xor U3802 (N_3802,N_3788,N_3693);
xor U3803 (N_3803,N_3741,N_3748);
and U3804 (N_3804,N_3626,N_3711);
or U3805 (N_3805,N_3658,N_3656);
nand U3806 (N_3806,N_3634,N_3617);
nand U3807 (N_3807,N_3663,N_3641);
and U3808 (N_3808,N_3676,N_3631);
and U3809 (N_3809,N_3616,N_3620);
xor U3810 (N_3810,N_3760,N_3678);
and U3811 (N_3811,N_3712,N_3689);
nor U3812 (N_3812,N_3691,N_3779);
nand U3813 (N_3813,N_3684,N_3766);
and U3814 (N_3814,N_3791,N_3787);
or U3815 (N_3815,N_3612,N_3661);
or U3816 (N_3816,N_3664,N_3733);
or U3817 (N_3817,N_3774,N_3671);
nand U3818 (N_3818,N_3708,N_3715);
nor U3819 (N_3819,N_3724,N_3746);
nor U3820 (N_3820,N_3710,N_3602);
and U3821 (N_3821,N_3627,N_3719);
xnor U3822 (N_3822,N_3694,N_3725);
nor U3823 (N_3823,N_3730,N_3754);
and U3824 (N_3824,N_3624,N_3759);
and U3825 (N_3825,N_3644,N_3610);
nand U3826 (N_3826,N_3669,N_3613);
nor U3827 (N_3827,N_3756,N_3652);
and U3828 (N_3828,N_3734,N_3655);
nand U3829 (N_3829,N_3793,N_3637);
and U3830 (N_3830,N_3687,N_3639);
nor U3831 (N_3831,N_3723,N_3640);
nand U3832 (N_3832,N_3778,N_3780);
and U3833 (N_3833,N_3607,N_3645);
xor U3834 (N_3834,N_3798,N_3773);
nor U3835 (N_3835,N_3785,N_3762);
and U3836 (N_3836,N_3628,N_3622);
xor U3837 (N_3837,N_3685,N_3717);
or U3838 (N_3838,N_3747,N_3750);
xnor U3839 (N_3839,N_3648,N_3647);
nor U3840 (N_3840,N_3764,N_3603);
or U3841 (N_3841,N_3621,N_3743);
or U3842 (N_3842,N_3770,N_3795);
or U3843 (N_3843,N_3775,N_3728);
or U3844 (N_3844,N_3635,N_3739);
nand U3845 (N_3845,N_3767,N_3799);
or U3846 (N_3846,N_3698,N_3681);
nor U3847 (N_3847,N_3769,N_3660);
xor U3848 (N_3848,N_3662,N_3713);
and U3849 (N_3849,N_3755,N_3782);
xnor U3850 (N_3850,N_3732,N_3757);
and U3851 (N_3851,N_3745,N_3736);
and U3852 (N_3852,N_3636,N_3704);
nand U3853 (N_3853,N_3797,N_3675);
nand U3854 (N_3854,N_3777,N_3625);
nor U3855 (N_3855,N_3646,N_3619);
or U3856 (N_3856,N_3789,N_3601);
and U3857 (N_3857,N_3649,N_3615);
xnor U3858 (N_3858,N_3659,N_3673);
nor U3859 (N_3859,N_3657,N_3792);
nor U3860 (N_3860,N_3674,N_3742);
xor U3861 (N_3861,N_3772,N_3683);
xor U3862 (N_3862,N_3630,N_3618);
nand U3863 (N_3863,N_3672,N_3716);
xor U3864 (N_3864,N_3642,N_3722);
nand U3865 (N_3865,N_3765,N_3729);
nor U3866 (N_3866,N_3706,N_3680);
nor U3867 (N_3867,N_3606,N_3703);
or U3868 (N_3868,N_3726,N_3668);
and U3869 (N_3869,N_3633,N_3771);
nand U3870 (N_3870,N_3608,N_3692);
and U3871 (N_3871,N_3702,N_3696);
and U3872 (N_3872,N_3749,N_3709);
nand U3873 (N_3873,N_3731,N_3651);
xor U3874 (N_3874,N_3718,N_3720);
and U3875 (N_3875,N_3679,N_3707);
nor U3876 (N_3876,N_3786,N_3697);
nor U3877 (N_3877,N_3721,N_3753);
nor U3878 (N_3878,N_3751,N_3768);
or U3879 (N_3879,N_3714,N_3600);
xnor U3880 (N_3880,N_3758,N_3737);
and U3881 (N_3881,N_3761,N_3700);
and U3882 (N_3882,N_3763,N_3643);
nor U3883 (N_3883,N_3604,N_3738);
and U3884 (N_3884,N_3611,N_3688);
nand U3885 (N_3885,N_3752,N_3653);
and U3886 (N_3886,N_3654,N_3632);
nand U3887 (N_3887,N_3796,N_3650);
and U3888 (N_3888,N_3727,N_3744);
xor U3889 (N_3889,N_3699,N_3665);
nor U3890 (N_3890,N_3690,N_3638);
xor U3891 (N_3891,N_3677,N_3686);
and U3892 (N_3892,N_3682,N_3614);
nand U3893 (N_3893,N_3695,N_3667);
or U3894 (N_3894,N_3701,N_3609);
nor U3895 (N_3895,N_3740,N_3629);
nor U3896 (N_3896,N_3705,N_3623);
xnor U3897 (N_3897,N_3666,N_3794);
and U3898 (N_3898,N_3670,N_3605);
nand U3899 (N_3899,N_3783,N_3735);
nor U3900 (N_3900,N_3787,N_3691);
nand U3901 (N_3901,N_3664,N_3600);
xor U3902 (N_3902,N_3749,N_3628);
nand U3903 (N_3903,N_3766,N_3619);
nand U3904 (N_3904,N_3742,N_3649);
xnor U3905 (N_3905,N_3749,N_3706);
or U3906 (N_3906,N_3629,N_3754);
and U3907 (N_3907,N_3681,N_3616);
or U3908 (N_3908,N_3768,N_3797);
and U3909 (N_3909,N_3715,N_3731);
or U3910 (N_3910,N_3765,N_3630);
or U3911 (N_3911,N_3785,N_3767);
nor U3912 (N_3912,N_3653,N_3766);
nor U3913 (N_3913,N_3655,N_3661);
xor U3914 (N_3914,N_3796,N_3611);
nor U3915 (N_3915,N_3671,N_3628);
xnor U3916 (N_3916,N_3684,N_3685);
or U3917 (N_3917,N_3668,N_3739);
and U3918 (N_3918,N_3663,N_3669);
nor U3919 (N_3919,N_3750,N_3785);
xnor U3920 (N_3920,N_3702,N_3660);
nor U3921 (N_3921,N_3794,N_3656);
or U3922 (N_3922,N_3624,N_3609);
nand U3923 (N_3923,N_3750,N_3766);
and U3924 (N_3924,N_3614,N_3663);
xor U3925 (N_3925,N_3696,N_3652);
nor U3926 (N_3926,N_3716,N_3715);
xnor U3927 (N_3927,N_3783,N_3640);
nor U3928 (N_3928,N_3710,N_3770);
xor U3929 (N_3929,N_3739,N_3610);
nand U3930 (N_3930,N_3790,N_3649);
nor U3931 (N_3931,N_3732,N_3663);
xnor U3932 (N_3932,N_3687,N_3737);
nand U3933 (N_3933,N_3733,N_3772);
and U3934 (N_3934,N_3728,N_3758);
nor U3935 (N_3935,N_3668,N_3717);
xnor U3936 (N_3936,N_3792,N_3715);
xor U3937 (N_3937,N_3642,N_3762);
and U3938 (N_3938,N_3744,N_3763);
nand U3939 (N_3939,N_3755,N_3633);
nor U3940 (N_3940,N_3767,N_3777);
nor U3941 (N_3941,N_3702,N_3654);
nor U3942 (N_3942,N_3639,N_3784);
nand U3943 (N_3943,N_3693,N_3782);
nor U3944 (N_3944,N_3749,N_3758);
and U3945 (N_3945,N_3672,N_3761);
and U3946 (N_3946,N_3660,N_3641);
nand U3947 (N_3947,N_3660,N_3652);
nor U3948 (N_3948,N_3724,N_3688);
nand U3949 (N_3949,N_3601,N_3720);
nor U3950 (N_3950,N_3719,N_3613);
xnor U3951 (N_3951,N_3627,N_3640);
and U3952 (N_3952,N_3794,N_3734);
or U3953 (N_3953,N_3734,N_3714);
xor U3954 (N_3954,N_3765,N_3600);
or U3955 (N_3955,N_3703,N_3673);
and U3956 (N_3956,N_3759,N_3639);
nand U3957 (N_3957,N_3601,N_3678);
xor U3958 (N_3958,N_3653,N_3793);
and U3959 (N_3959,N_3791,N_3629);
nand U3960 (N_3960,N_3689,N_3667);
and U3961 (N_3961,N_3605,N_3608);
and U3962 (N_3962,N_3660,N_3657);
and U3963 (N_3963,N_3612,N_3602);
or U3964 (N_3964,N_3758,N_3734);
nand U3965 (N_3965,N_3714,N_3712);
nand U3966 (N_3966,N_3796,N_3718);
nor U3967 (N_3967,N_3743,N_3739);
nand U3968 (N_3968,N_3783,N_3758);
or U3969 (N_3969,N_3669,N_3793);
and U3970 (N_3970,N_3792,N_3725);
xnor U3971 (N_3971,N_3696,N_3754);
nand U3972 (N_3972,N_3689,N_3610);
or U3973 (N_3973,N_3782,N_3643);
xnor U3974 (N_3974,N_3731,N_3642);
nand U3975 (N_3975,N_3604,N_3770);
nand U3976 (N_3976,N_3632,N_3677);
nand U3977 (N_3977,N_3607,N_3634);
or U3978 (N_3978,N_3621,N_3635);
nand U3979 (N_3979,N_3753,N_3799);
and U3980 (N_3980,N_3737,N_3613);
xor U3981 (N_3981,N_3690,N_3778);
nand U3982 (N_3982,N_3709,N_3731);
or U3983 (N_3983,N_3763,N_3659);
nand U3984 (N_3984,N_3779,N_3704);
xnor U3985 (N_3985,N_3659,N_3644);
and U3986 (N_3986,N_3663,N_3694);
xnor U3987 (N_3987,N_3697,N_3722);
and U3988 (N_3988,N_3715,N_3603);
and U3989 (N_3989,N_3675,N_3668);
and U3990 (N_3990,N_3692,N_3629);
nand U3991 (N_3991,N_3603,N_3787);
nand U3992 (N_3992,N_3671,N_3790);
xnor U3993 (N_3993,N_3653,N_3784);
nand U3994 (N_3994,N_3698,N_3723);
or U3995 (N_3995,N_3622,N_3795);
and U3996 (N_3996,N_3673,N_3792);
nand U3997 (N_3997,N_3657,N_3614);
nor U3998 (N_3998,N_3780,N_3628);
or U3999 (N_3999,N_3656,N_3748);
nand U4000 (N_4000,N_3839,N_3858);
nor U4001 (N_4001,N_3854,N_3926);
or U4002 (N_4002,N_3985,N_3977);
or U4003 (N_4003,N_3894,N_3984);
nor U4004 (N_4004,N_3893,N_3986);
and U4005 (N_4005,N_3993,N_3825);
or U4006 (N_4006,N_3980,N_3949);
or U4007 (N_4007,N_3955,N_3807);
xnor U4008 (N_4008,N_3939,N_3982);
or U4009 (N_4009,N_3874,N_3851);
or U4010 (N_4010,N_3952,N_3948);
xor U4011 (N_4011,N_3898,N_3885);
nor U4012 (N_4012,N_3959,N_3826);
or U4013 (N_4013,N_3829,N_3996);
or U4014 (N_4014,N_3922,N_3877);
nor U4015 (N_4015,N_3816,N_3916);
xor U4016 (N_4016,N_3850,N_3962);
or U4017 (N_4017,N_3995,N_3805);
nand U4018 (N_4018,N_3950,N_3987);
xor U4019 (N_4019,N_3815,N_3974);
nor U4020 (N_4020,N_3803,N_3998);
xnor U4021 (N_4021,N_3923,N_3904);
nor U4022 (N_4022,N_3873,N_3837);
xor U4023 (N_4023,N_3888,N_3835);
nor U4024 (N_4024,N_3940,N_3981);
xor U4025 (N_4025,N_3957,N_3883);
nor U4026 (N_4026,N_3832,N_3869);
nand U4027 (N_4027,N_3802,N_3897);
or U4028 (N_4028,N_3817,N_3820);
xnor U4029 (N_4029,N_3983,N_3831);
nand U4030 (N_4030,N_3862,N_3936);
nand U4031 (N_4031,N_3878,N_3863);
and U4032 (N_4032,N_3935,N_3997);
and U4033 (N_4033,N_3823,N_3901);
xnor U4034 (N_4034,N_3961,N_3965);
and U4035 (N_4035,N_3818,N_3887);
nor U4036 (N_4036,N_3973,N_3937);
and U4037 (N_4037,N_3848,N_3830);
or U4038 (N_4038,N_3907,N_3975);
nand U4039 (N_4039,N_3889,N_3976);
or U4040 (N_4040,N_3913,N_3842);
xor U4041 (N_4041,N_3972,N_3882);
xor U4042 (N_4042,N_3969,N_3932);
nand U4043 (N_4043,N_3819,N_3876);
and U4044 (N_4044,N_3903,N_3872);
xnor U4045 (N_4045,N_3956,N_3895);
nor U4046 (N_4046,N_3875,N_3960);
or U4047 (N_4047,N_3989,N_3917);
or U4048 (N_4048,N_3990,N_3945);
nor U4049 (N_4049,N_3841,N_3967);
nand U4050 (N_4050,N_3920,N_3924);
nor U4051 (N_4051,N_3906,N_3810);
or U4052 (N_4052,N_3951,N_3812);
or U4053 (N_4053,N_3813,N_3840);
xor U4054 (N_4054,N_3827,N_3927);
or U4055 (N_4055,N_3910,N_3800);
or U4056 (N_4056,N_3919,N_3908);
xnor U4057 (N_4057,N_3915,N_3867);
xnor U4058 (N_4058,N_3892,N_3999);
xor U4059 (N_4059,N_3931,N_3943);
nor U4060 (N_4060,N_3804,N_3970);
nor U4061 (N_4061,N_3861,N_3966);
nor U4062 (N_4062,N_3806,N_3994);
nand U4063 (N_4063,N_3822,N_3871);
nand U4064 (N_4064,N_3844,N_3953);
and U4065 (N_4065,N_3857,N_3947);
nand U4066 (N_4066,N_3801,N_3828);
xor U4067 (N_4067,N_3902,N_3941);
nand U4068 (N_4068,N_3944,N_3880);
xnor U4069 (N_4069,N_3836,N_3847);
nor U4070 (N_4070,N_3925,N_3938);
nand U4071 (N_4071,N_3864,N_3954);
xnor U4072 (N_4072,N_3853,N_3881);
nor U4073 (N_4073,N_3934,N_3884);
or U4074 (N_4074,N_3933,N_3814);
and U4075 (N_4075,N_3890,N_3905);
nand U4076 (N_4076,N_3870,N_3866);
xnor U4077 (N_4077,N_3988,N_3891);
xnor U4078 (N_4078,N_3886,N_3843);
and U4079 (N_4079,N_3809,N_3968);
nor U4080 (N_4080,N_3911,N_3921);
and U4081 (N_4081,N_3868,N_3942);
and U4082 (N_4082,N_3821,N_3852);
nand U4083 (N_4083,N_3811,N_3963);
nand U4084 (N_4084,N_3846,N_3855);
xor U4085 (N_4085,N_3879,N_3958);
nor U4086 (N_4086,N_3838,N_3964);
nand U4087 (N_4087,N_3896,N_3845);
or U4088 (N_4088,N_3978,N_3930);
or U4089 (N_4089,N_3900,N_3991);
xnor U4090 (N_4090,N_3859,N_3824);
or U4091 (N_4091,N_3914,N_3979);
xor U4092 (N_4092,N_3992,N_3899);
and U4093 (N_4093,N_3849,N_3909);
or U4094 (N_4094,N_3912,N_3971);
nor U4095 (N_4095,N_3928,N_3918);
or U4096 (N_4096,N_3856,N_3808);
and U4097 (N_4097,N_3946,N_3929);
xor U4098 (N_4098,N_3865,N_3833);
xor U4099 (N_4099,N_3860,N_3834);
nand U4100 (N_4100,N_3992,N_3999);
nor U4101 (N_4101,N_3822,N_3898);
nor U4102 (N_4102,N_3961,N_3833);
or U4103 (N_4103,N_3804,N_3820);
xor U4104 (N_4104,N_3856,N_3927);
xor U4105 (N_4105,N_3918,N_3854);
xor U4106 (N_4106,N_3995,N_3804);
or U4107 (N_4107,N_3953,N_3819);
or U4108 (N_4108,N_3977,N_3839);
nand U4109 (N_4109,N_3836,N_3864);
nor U4110 (N_4110,N_3860,N_3845);
nand U4111 (N_4111,N_3953,N_3962);
nand U4112 (N_4112,N_3982,N_3947);
nand U4113 (N_4113,N_3945,N_3940);
nand U4114 (N_4114,N_3966,N_3894);
nand U4115 (N_4115,N_3976,N_3967);
nor U4116 (N_4116,N_3955,N_3881);
or U4117 (N_4117,N_3938,N_3986);
or U4118 (N_4118,N_3937,N_3899);
or U4119 (N_4119,N_3936,N_3996);
nand U4120 (N_4120,N_3943,N_3894);
xnor U4121 (N_4121,N_3807,N_3938);
and U4122 (N_4122,N_3818,N_3815);
xor U4123 (N_4123,N_3813,N_3966);
and U4124 (N_4124,N_3975,N_3916);
nand U4125 (N_4125,N_3966,N_3993);
nor U4126 (N_4126,N_3957,N_3958);
nand U4127 (N_4127,N_3819,N_3917);
nand U4128 (N_4128,N_3970,N_3876);
and U4129 (N_4129,N_3910,N_3992);
xnor U4130 (N_4130,N_3971,N_3834);
or U4131 (N_4131,N_3813,N_3924);
nor U4132 (N_4132,N_3857,N_3894);
nand U4133 (N_4133,N_3864,N_3802);
nor U4134 (N_4134,N_3904,N_3983);
nor U4135 (N_4135,N_3963,N_3955);
and U4136 (N_4136,N_3870,N_3876);
and U4137 (N_4137,N_3810,N_3872);
nor U4138 (N_4138,N_3856,N_3969);
nor U4139 (N_4139,N_3934,N_3903);
nand U4140 (N_4140,N_3926,N_3800);
nand U4141 (N_4141,N_3826,N_3901);
and U4142 (N_4142,N_3878,N_3921);
and U4143 (N_4143,N_3918,N_3991);
nand U4144 (N_4144,N_3957,N_3898);
and U4145 (N_4145,N_3919,N_3822);
nor U4146 (N_4146,N_3808,N_3876);
or U4147 (N_4147,N_3833,N_3847);
or U4148 (N_4148,N_3924,N_3922);
nand U4149 (N_4149,N_3948,N_3880);
or U4150 (N_4150,N_3903,N_3988);
xnor U4151 (N_4151,N_3907,N_3993);
nand U4152 (N_4152,N_3969,N_3972);
and U4153 (N_4153,N_3993,N_3863);
xor U4154 (N_4154,N_3886,N_3988);
nor U4155 (N_4155,N_3893,N_3814);
xnor U4156 (N_4156,N_3821,N_3979);
and U4157 (N_4157,N_3866,N_3972);
xor U4158 (N_4158,N_3866,N_3973);
nand U4159 (N_4159,N_3828,N_3804);
and U4160 (N_4160,N_3966,N_3906);
xor U4161 (N_4161,N_3850,N_3873);
nor U4162 (N_4162,N_3942,N_3925);
or U4163 (N_4163,N_3933,N_3905);
xnor U4164 (N_4164,N_3830,N_3800);
nand U4165 (N_4165,N_3975,N_3998);
and U4166 (N_4166,N_3915,N_3870);
and U4167 (N_4167,N_3979,N_3927);
xor U4168 (N_4168,N_3942,N_3860);
or U4169 (N_4169,N_3820,N_3877);
nor U4170 (N_4170,N_3858,N_3962);
and U4171 (N_4171,N_3962,N_3802);
or U4172 (N_4172,N_3901,N_3843);
nor U4173 (N_4173,N_3930,N_3865);
nor U4174 (N_4174,N_3861,N_3896);
xnor U4175 (N_4175,N_3963,N_3977);
nand U4176 (N_4176,N_3821,N_3819);
nand U4177 (N_4177,N_3910,N_3977);
xor U4178 (N_4178,N_3863,N_3897);
xor U4179 (N_4179,N_3992,N_3857);
and U4180 (N_4180,N_3847,N_3809);
nand U4181 (N_4181,N_3878,N_3956);
nor U4182 (N_4182,N_3936,N_3938);
nand U4183 (N_4183,N_3970,N_3801);
and U4184 (N_4184,N_3909,N_3809);
xor U4185 (N_4185,N_3945,N_3881);
xnor U4186 (N_4186,N_3947,N_3820);
or U4187 (N_4187,N_3948,N_3801);
or U4188 (N_4188,N_3958,N_3962);
or U4189 (N_4189,N_3861,N_3822);
or U4190 (N_4190,N_3984,N_3937);
or U4191 (N_4191,N_3924,N_3976);
xor U4192 (N_4192,N_3882,N_3804);
xnor U4193 (N_4193,N_3899,N_3864);
xnor U4194 (N_4194,N_3995,N_3910);
nand U4195 (N_4195,N_3874,N_3899);
nor U4196 (N_4196,N_3806,N_3824);
or U4197 (N_4197,N_3942,N_3940);
nor U4198 (N_4198,N_3971,N_3988);
nand U4199 (N_4199,N_3957,N_3806);
or U4200 (N_4200,N_4194,N_4017);
xnor U4201 (N_4201,N_4129,N_4006);
and U4202 (N_4202,N_4057,N_4103);
nor U4203 (N_4203,N_4077,N_4113);
and U4204 (N_4204,N_4065,N_4169);
xnor U4205 (N_4205,N_4097,N_4162);
nand U4206 (N_4206,N_4196,N_4166);
nand U4207 (N_4207,N_4193,N_4188);
nor U4208 (N_4208,N_4107,N_4036);
or U4209 (N_4209,N_4091,N_4032);
xor U4210 (N_4210,N_4068,N_4198);
nor U4211 (N_4211,N_4058,N_4126);
or U4212 (N_4212,N_4012,N_4165);
nor U4213 (N_4213,N_4007,N_4128);
nand U4214 (N_4214,N_4172,N_4079);
xnor U4215 (N_4215,N_4029,N_4019);
xnor U4216 (N_4216,N_4054,N_4038);
or U4217 (N_4217,N_4050,N_4021);
or U4218 (N_4218,N_4060,N_4144);
and U4219 (N_4219,N_4010,N_4122);
or U4220 (N_4220,N_4150,N_4000);
xnor U4221 (N_4221,N_4022,N_4143);
xor U4222 (N_4222,N_4084,N_4180);
nor U4223 (N_4223,N_4158,N_4127);
xnor U4224 (N_4224,N_4072,N_4189);
or U4225 (N_4225,N_4136,N_4089);
nand U4226 (N_4226,N_4164,N_4004);
xor U4227 (N_4227,N_4159,N_4005);
or U4228 (N_4228,N_4098,N_4132);
or U4229 (N_4229,N_4121,N_4048);
nand U4230 (N_4230,N_4120,N_4197);
nor U4231 (N_4231,N_4140,N_4085);
xnor U4232 (N_4232,N_4053,N_4177);
or U4233 (N_4233,N_4183,N_4145);
xnor U4234 (N_4234,N_4192,N_4039);
and U4235 (N_4235,N_4047,N_4033);
xor U4236 (N_4236,N_4106,N_4093);
nor U4237 (N_4237,N_4049,N_4104);
or U4238 (N_4238,N_4149,N_4185);
and U4239 (N_4239,N_4034,N_4105);
nor U4240 (N_4240,N_4073,N_4024);
nand U4241 (N_4241,N_4176,N_4043);
and U4242 (N_4242,N_4152,N_4002);
or U4243 (N_4243,N_4088,N_4195);
and U4244 (N_4244,N_4118,N_4109);
nor U4245 (N_4245,N_4061,N_4167);
or U4246 (N_4246,N_4171,N_4100);
and U4247 (N_4247,N_4044,N_4151);
xnor U4248 (N_4248,N_4134,N_4018);
and U4249 (N_4249,N_4069,N_4090);
and U4250 (N_4250,N_4011,N_4020);
xnor U4251 (N_4251,N_4092,N_4028);
and U4252 (N_4252,N_4131,N_4087);
and U4253 (N_4253,N_4045,N_4095);
nand U4254 (N_4254,N_4133,N_4147);
or U4255 (N_4255,N_4070,N_4081);
and U4256 (N_4256,N_4067,N_4124);
nor U4257 (N_4257,N_4137,N_4052);
nor U4258 (N_4258,N_4080,N_4064);
nor U4259 (N_4259,N_4001,N_4123);
or U4260 (N_4260,N_4117,N_4157);
nand U4261 (N_4261,N_4115,N_4026);
nand U4262 (N_4262,N_4178,N_4191);
nor U4263 (N_4263,N_4186,N_4146);
and U4264 (N_4264,N_4108,N_4155);
or U4265 (N_4265,N_4040,N_4173);
and U4266 (N_4266,N_4030,N_4111);
xor U4267 (N_4267,N_4078,N_4014);
nand U4268 (N_4268,N_4042,N_4076);
and U4269 (N_4269,N_4125,N_4035);
nand U4270 (N_4270,N_4056,N_4016);
and U4271 (N_4271,N_4175,N_4025);
or U4272 (N_4272,N_4156,N_4160);
xor U4273 (N_4273,N_4199,N_4153);
or U4274 (N_4274,N_4094,N_4142);
xnor U4275 (N_4275,N_4139,N_4101);
or U4276 (N_4276,N_4027,N_4074);
nand U4277 (N_4277,N_4059,N_4135);
and U4278 (N_4278,N_4130,N_4003);
or U4279 (N_4279,N_4179,N_4114);
nand U4280 (N_4280,N_4184,N_4141);
or U4281 (N_4281,N_4083,N_4041);
nand U4282 (N_4282,N_4009,N_4046);
and U4283 (N_4283,N_4008,N_4096);
or U4284 (N_4284,N_4082,N_4110);
xor U4285 (N_4285,N_4023,N_4174);
nand U4286 (N_4286,N_4037,N_4161);
xor U4287 (N_4287,N_4154,N_4031);
or U4288 (N_4288,N_4190,N_4119);
nand U4289 (N_4289,N_4015,N_4112);
nor U4290 (N_4290,N_4102,N_4187);
nor U4291 (N_4291,N_4181,N_4138);
xor U4292 (N_4292,N_4075,N_4063);
nand U4293 (N_4293,N_4170,N_4013);
and U4294 (N_4294,N_4071,N_4168);
nand U4295 (N_4295,N_4148,N_4163);
and U4296 (N_4296,N_4086,N_4051);
and U4297 (N_4297,N_4062,N_4055);
xnor U4298 (N_4298,N_4116,N_4182);
nand U4299 (N_4299,N_4066,N_4099);
nand U4300 (N_4300,N_4038,N_4165);
or U4301 (N_4301,N_4105,N_4122);
xnor U4302 (N_4302,N_4149,N_4027);
and U4303 (N_4303,N_4139,N_4013);
nand U4304 (N_4304,N_4055,N_4079);
and U4305 (N_4305,N_4066,N_4121);
and U4306 (N_4306,N_4116,N_4138);
nand U4307 (N_4307,N_4007,N_4131);
nor U4308 (N_4308,N_4063,N_4124);
nor U4309 (N_4309,N_4021,N_4009);
or U4310 (N_4310,N_4057,N_4155);
or U4311 (N_4311,N_4040,N_4079);
xor U4312 (N_4312,N_4036,N_4185);
nor U4313 (N_4313,N_4108,N_4111);
or U4314 (N_4314,N_4097,N_4125);
and U4315 (N_4315,N_4052,N_4106);
xnor U4316 (N_4316,N_4036,N_4159);
nand U4317 (N_4317,N_4115,N_4056);
and U4318 (N_4318,N_4137,N_4130);
or U4319 (N_4319,N_4159,N_4107);
nand U4320 (N_4320,N_4005,N_4104);
or U4321 (N_4321,N_4147,N_4004);
and U4322 (N_4322,N_4050,N_4037);
or U4323 (N_4323,N_4007,N_4021);
or U4324 (N_4324,N_4097,N_4164);
xnor U4325 (N_4325,N_4187,N_4182);
nand U4326 (N_4326,N_4022,N_4109);
nor U4327 (N_4327,N_4019,N_4009);
nor U4328 (N_4328,N_4114,N_4001);
nor U4329 (N_4329,N_4004,N_4115);
nor U4330 (N_4330,N_4031,N_4071);
xor U4331 (N_4331,N_4025,N_4019);
nand U4332 (N_4332,N_4095,N_4030);
or U4333 (N_4333,N_4036,N_4180);
nand U4334 (N_4334,N_4035,N_4189);
nand U4335 (N_4335,N_4130,N_4033);
or U4336 (N_4336,N_4122,N_4197);
or U4337 (N_4337,N_4139,N_4069);
xor U4338 (N_4338,N_4170,N_4182);
or U4339 (N_4339,N_4022,N_4014);
nor U4340 (N_4340,N_4010,N_4054);
and U4341 (N_4341,N_4176,N_4001);
and U4342 (N_4342,N_4002,N_4108);
and U4343 (N_4343,N_4019,N_4124);
and U4344 (N_4344,N_4168,N_4017);
or U4345 (N_4345,N_4013,N_4098);
nor U4346 (N_4346,N_4054,N_4011);
or U4347 (N_4347,N_4142,N_4062);
nand U4348 (N_4348,N_4109,N_4111);
and U4349 (N_4349,N_4133,N_4176);
and U4350 (N_4350,N_4123,N_4052);
or U4351 (N_4351,N_4121,N_4109);
or U4352 (N_4352,N_4165,N_4158);
nor U4353 (N_4353,N_4075,N_4153);
nor U4354 (N_4354,N_4088,N_4021);
or U4355 (N_4355,N_4048,N_4195);
nand U4356 (N_4356,N_4150,N_4197);
nand U4357 (N_4357,N_4141,N_4097);
nor U4358 (N_4358,N_4051,N_4188);
nand U4359 (N_4359,N_4083,N_4090);
or U4360 (N_4360,N_4173,N_4000);
or U4361 (N_4361,N_4010,N_4084);
nand U4362 (N_4362,N_4109,N_4197);
nand U4363 (N_4363,N_4021,N_4144);
or U4364 (N_4364,N_4139,N_4067);
nor U4365 (N_4365,N_4010,N_4069);
nor U4366 (N_4366,N_4177,N_4160);
nand U4367 (N_4367,N_4022,N_4035);
or U4368 (N_4368,N_4000,N_4064);
xor U4369 (N_4369,N_4173,N_4033);
or U4370 (N_4370,N_4159,N_4034);
nor U4371 (N_4371,N_4071,N_4029);
xor U4372 (N_4372,N_4193,N_4125);
xor U4373 (N_4373,N_4168,N_4077);
xnor U4374 (N_4374,N_4189,N_4148);
nand U4375 (N_4375,N_4070,N_4034);
nor U4376 (N_4376,N_4116,N_4068);
or U4377 (N_4377,N_4129,N_4039);
xnor U4378 (N_4378,N_4174,N_4182);
or U4379 (N_4379,N_4012,N_4059);
or U4380 (N_4380,N_4150,N_4102);
or U4381 (N_4381,N_4176,N_4029);
or U4382 (N_4382,N_4055,N_4117);
or U4383 (N_4383,N_4158,N_4191);
nand U4384 (N_4384,N_4131,N_4097);
and U4385 (N_4385,N_4177,N_4048);
or U4386 (N_4386,N_4090,N_4183);
nand U4387 (N_4387,N_4138,N_4197);
nand U4388 (N_4388,N_4171,N_4136);
nor U4389 (N_4389,N_4025,N_4036);
nand U4390 (N_4390,N_4193,N_4028);
nor U4391 (N_4391,N_4077,N_4102);
or U4392 (N_4392,N_4052,N_4186);
or U4393 (N_4393,N_4120,N_4178);
xnor U4394 (N_4394,N_4031,N_4148);
and U4395 (N_4395,N_4187,N_4115);
xnor U4396 (N_4396,N_4009,N_4181);
nor U4397 (N_4397,N_4057,N_4030);
and U4398 (N_4398,N_4068,N_4006);
xor U4399 (N_4399,N_4186,N_4079);
nor U4400 (N_4400,N_4330,N_4314);
xnor U4401 (N_4401,N_4393,N_4390);
or U4402 (N_4402,N_4354,N_4395);
or U4403 (N_4403,N_4289,N_4215);
nand U4404 (N_4404,N_4300,N_4341);
or U4405 (N_4405,N_4281,N_4368);
nand U4406 (N_4406,N_4373,N_4356);
xor U4407 (N_4407,N_4298,N_4308);
xor U4408 (N_4408,N_4374,N_4222);
nor U4409 (N_4409,N_4353,N_4247);
nand U4410 (N_4410,N_4325,N_4227);
nand U4411 (N_4411,N_4349,N_4223);
nor U4412 (N_4412,N_4217,N_4329);
nor U4413 (N_4413,N_4305,N_4299);
or U4414 (N_4414,N_4372,N_4363);
nor U4415 (N_4415,N_4271,N_4234);
nor U4416 (N_4416,N_4243,N_4250);
nor U4417 (N_4417,N_4273,N_4352);
or U4418 (N_4418,N_4318,N_4362);
or U4419 (N_4419,N_4361,N_4360);
and U4420 (N_4420,N_4212,N_4224);
xnor U4421 (N_4421,N_4201,N_4328);
nand U4422 (N_4422,N_4336,N_4275);
nor U4423 (N_4423,N_4254,N_4256);
nand U4424 (N_4424,N_4295,N_4345);
nor U4425 (N_4425,N_4204,N_4249);
nor U4426 (N_4426,N_4294,N_4214);
and U4427 (N_4427,N_4288,N_4303);
and U4428 (N_4428,N_4225,N_4241);
and U4429 (N_4429,N_4283,N_4244);
xnor U4430 (N_4430,N_4348,N_4280);
nand U4431 (N_4431,N_4231,N_4350);
nand U4432 (N_4432,N_4268,N_4251);
xnor U4433 (N_4433,N_4310,N_4388);
or U4434 (N_4434,N_4376,N_4226);
or U4435 (N_4435,N_4302,N_4365);
xor U4436 (N_4436,N_4324,N_4320);
xor U4437 (N_4437,N_4357,N_4316);
nor U4438 (N_4438,N_4384,N_4342);
or U4439 (N_4439,N_4210,N_4291);
and U4440 (N_4440,N_4208,N_4367);
or U4441 (N_4441,N_4257,N_4380);
nor U4442 (N_4442,N_4202,N_4266);
and U4443 (N_4443,N_4397,N_4209);
nor U4444 (N_4444,N_4386,N_4265);
nor U4445 (N_4445,N_4293,N_4383);
xor U4446 (N_4446,N_4355,N_4205);
xor U4447 (N_4447,N_4274,N_4370);
nor U4448 (N_4448,N_4375,N_4272);
or U4449 (N_4449,N_4358,N_4239);
xor U4450 (N_4450,N_4396,N_4344);
xnor U4451 (N_4451,N_4269,N_4304);
and U4452 (N_4452,N_4259,N_4220);
and U4453 (N_4453,N_4366,N_4240);
xnor U4454 (N_4454,N_4238,N_4385);
nor U4455 (N_4455,N_4399,N_4253);
or U4456 (N_4456,N_4233,N_4230);
or U4457 (N_4457,N_4279,N_4287);
xor U4458 (N_4458,N_4282,N_4377);
xor U4459 (N_4459,N_4301,N_4260);
nand U4460 (N_4460,N_4292,N_4248);
xor U4461 (N_4461,N_4270,N_4319);
and U4462 (N_4462,N_4277,N_4252);
and U4463 (N_4463,N_4242,N_4246);
and U4464 (N_4464,N_4317,N_4286);
nor U4465 (N_4465,N_4284,N_4331);
and U4466 (N_4466,N_4258,N_4381);
nor U4467 (N_4467,N_4387,N_4369);
nor U4468 (N_4468,N_4236,N_4335);
and U4469 (N_4469,N_4309,N_4321);
nand U4470 (N_4470,N_4327,N_4211);
nand U4471 (N_4471,N_4340,N_4263);
and U4472 (N_4472,N_4219,N_4262);
or U4473 (N_4473,N_4255,N_4326);
nand U4474 (N_4474,N_4228,N_4278);
and U4475 (N_4475,N_4245,N_4359);
xnor U4476 (N_4476,N_4285,N_4261);
nand U4477 (N_4477,N_4206,N_4313);
nand U4478 (N_4478,N_4267,N_4237);
and U4479 (N_4479,N_4391,N_4351);
or U4480 (N_4480,N_4323,N_4276);
nand U4481 (N_4481,N_4218,N_4382);
nand U4482 (N_4482,N_4296,N_4394);
and U4483 (N_4483,N_4312,N_4297);
nand U4484 (N_4484,N_4378,N_4334);
xnor U4485 (N_4485,N_4307,N_4371);
nor U4486 (N_4486,N_4290,N_4339);
nor U4487 (N_4487,N_4200,N_4392);
or U4488 (N_4488,N_4364,N_4338);
nand U4489 (N_4489,N_4221,N_4332);
or U4490 (N_4490,N_4235,N_4337);
xnor U4491 (N_4491,N_4229,N_4347);
xor U4492 (N_4492,N_4216,N_4232);
or U4493 (N_4493,N_4346,N_4306);
or U4494 (N_4494,N_4203,N_4207);
and U4495 (N_4495,N_4213,N_4322);
nand U4496 (N_4496,N_4389,N_4343);
nand U4497 (N_4497,N_4379,N_4311);
xor U4498 (N_4498,N_4398,N_4333);
and U4499 (N_4499,N_4315,N_4264);
nor U4500 (N_4500,N_4357,N_4245);
or U4501 (N_4501,N_4315,N_4342);
xnor U4502 (N_4502,N_4249,N_4329);
nand U4503 (N_4503,N_4273,N_4303);
nand U4504 (N_4504,N_4251,N_4293);
or U4505 (N_4505,N_4259,N_4209);
nor U4506 (N_4506,N_4370,N_4368);
or U4507 (N_4507,N_4333,N_4275);
nor U4508 (N_4508,N_4253,N_4286);
xnor U4509 (N_4509,N_4276,N_4397);
or U4510 (N_4510,N_4205,N_4399);
nand U4511 (N_4511,N_4272,N_4234);
xor U4512 (N_4512,N_4242,N_4219);
and U4513 (N_4513,N_4288,N_4276);
xnor U4514 (N_4514,N_4318,N_4245);
and U4515 (N_4515,N_4300,N_4291);
or U4516 (N_4516,N_4333,N_4387);
nor U4517 (N_4517,N_4380,N_4276);
or U4518 (N_4518,N_4322,N_4382);
or U4519 (N_4519,N_4298,N_4225);
or U4520 (N_4520,N_4330,N_4297);
nand U4521 (N_4521,N_4319,N_4399);
xnor U4522 (N_4522,N_4334,N_4391);
or U4523 (N_4523,N_4216,N_4214);
nor U4524 (N_4524,N_4379,N_4393);
nor U4525 (N_4525,N_4250,N_4315);
or U4526 (N_4526,N_4222,N_4221);
nor U4527 (N_4527,N_4241,N_4331);
nor U4528 (N_4528,N_4330,N_4265);
or U4529 (N_4529,N_4285,N_4394);
and U4530 (N_4530,N_4227,N_4335);
xor U4531 (N_4531,N_4332,N_4275);
nand U4532 (N_4532,N_4247,N_4334);
nand U4533 (N_4533,N_4393,N_4267);
or U4534 (N_4534,N_4223,N_4367);
nand U4535 (N_4535,N_4333,N_4223);
nor U4536 (N_4536,N_4331,N_4210);
and U4537 (N_4537,N_4246,N_4397);
xor U4538 (N_4538,N_4344,N_4265);
nor U4539 (N_4539,N_4319,N_4214);
and U4540 (N_4540,N_4369,N_4320);
xor U4541 (N_4541,N_4222,N_4216);
nand U4542 (N_4542,N_4381,N_4262);
or U4543 (N_4543,N_4377,N_4207);
xnor U4544 (N_4544,N_4220,N_4315);
or U4545 (N_4545,N_4399,N_4339);
and U4546 (N_4546,N_4245,N_4356);
nand U4547 (N_4547,N_4338,N_4358);
nor U4548 (N_4548,N_4329,N_4283);
nor U4549 (N_4549,N_4246,N_4374);
nand U4550 (N_4550,N_4254,N_4225);
and U4551 (N_4551,N_4390,N_4269);
nand U4552 (N_4552,N_4304,N_4396);
nand U4553 (N_4553,N_4398,N_4304);
xor U4554 (N_4554,N_4256,N_4357);
xnor U4555 (N_4555,N_4304,N_4252);
xor U4556 (N_4556,N_4293,N_4394);
or U4557 (N_4557,N_4334,N_4288);
and U4558 (N_4558,N_4376,N_4273);
nor U4559 (N_4559,N_4315,N_4278);
nand U4560 (N_4560,N_4227,N_4210);
xnor U4561 (N_4561,N_4385,N_4381);
or U4562 (N_4562,N_4224,N_4253);
nand U4563 (N_4563,N_4359,N_4303);
nand U4564 (N_4564,N_4379,N_4396);
nor U4565 (N_4565,N_4248,N_4234);
xnor U4566 (N_4566,N_4394,N_4248);
and U4567 (N_4567,N_4294,N_4228);
or U4568 (N_4568,N_4341,N_4278);
nor U4569 (N_4569,N_4345,N_4206);
xor U4570 (N_4570,N_4307,N_4207);
and U4571 (N_4571,N_4274,N_4385);
nor U4572 (N_4572,N_4328,N_4220);
nand U4573 (N_4573,N_4200,N_4279);
or U4574 (N_4574,N_4237,N_4220);
or U4575 (N_4575,N_4323,N_4259);
xor U4576 (N_4576,N_4393,N_4332);
and U4577 (N_4577,N_4348,N_4342);
nor U4578 (N_4578,N_4380,N_4215);
and U4579 (N_4579,N_4354,N_4290);
xnor U4580 (N_4580,N_4357,N_4215);
nor U4581 (N_4581,N_4278,N_4208);
nand U4582 (N_4582,N_4390,N_4377);
and U4583 (N_4583,N_4318,N_4214);
xor U4584 (N_4584,N_4388,N_4317);
or U4585 (N_4585,N_4378,N_4357);
xor U4586 (N_4586,N_4245,N_4378);
nor U4587 (N_4587,N_4207,N_4290);
or U4588 (N_4588,N_4247,N_4208);
nor U4589 (N_4589,N_4376,N_4224);
or U4590 (N_4590,N_4259,N_4288);
and U4591 (N_4591,N_4323,N_4395);
or U4592 (N_4592,N_4201,N_4250);
nor U4593 (N_4593,N_4262,N_4225);
and U4594 (N_4594,N_4324,N_4264);
nor U4595 (N_4595,N_4286,N_4393);
or U4596 (N_4596,N_4234,N_4209);
nor U4597 (N_4597,N_4325,N_4308);
nor U4598 (N_4598,N_4258,N_4296);
nor U4599 (N_4599,N_4364,N_4359);
and U4600 (N_4600,N_4516,N_4560);
xnor U4601 (N_4601,N_4475,N_4499);
xnor U4602 (N_4602,N_4425,N_4507);
or U4603 (N_4603,N_4583,N_4474);
nand U4604 (N_4604,N_4437,N_4549);
nor U4605 (N_4605,N_4594,N_4568);
xor U4606 (N_4606,N_4466,N_4447);
or U4607 (N_4607,N_4543,N_4426);
nor U4608 (N_4608,N_4409,N_4461);
xnor U4609 (N_4609,N_4443,N_4451);
and U4610 (N_4610,N_4439,N_4541);
xor U4611 (N_4611,N_4411,N_4533);
xnor U4612 (N_4612,N_4542,N_4529);
and U4613 (N_4613,N_4492,N_4571);
nand U4614 (N_4614,N_4478,N_4458);
or U4615 (N_4615,N_4579,N_4525);
or U4616 (N_4616,N_4471,N_4555);
xnor U4617 (N_4617,N_4495,N_4587);
or U4618 (N_4618,N_4422,N_4586);
xnor U4619 (N_4619,N_4420,N_4427);
xnor U4620 (N_4620,N_4459,N_4527);
nand U4621 (N_4621,N_4538,N_4450);
or U4622 (N_4622,N_4554,N_4530);
or U4623 (N_4623,N_4517,N_4493);
or U4624 (N_4624,N_4569,N_4465);
or U4625 (N_4625,N_4536,N_4598);
xor U4626 (N_4626,N_4490,N_4468);
xnor U4627 (N_4627,N_4513,N_4452);
or U4628 (N_4628,N_4562,N_4593);
xor U4629 (N_4629,N_4528,N_4585);
xnor U4630 (N_4630,N_4547,N_4537);
nor U4631 (N_4631,N_4556,N_4494);
nor U4632 (N_4632,N_4462,N_4557);
nand U4633 (N_4633,N_4421,N_4472);
nand U4634 (N_4634,N_4417,N_4401);
nand U4635 (N_4635,N_4581,N_4481);
nor U4636 (N_4636,N_4505,N_4546);
nor U4637 (N_4637,N_4564,N_4498);
and U4638 (N_4638,N_4503,N_4436);
nand U4639 (N_4639,N_4489,N_4567);
nand U4640 (N_4640,N_4403,N_4497);
nor U4641 (N_4641,N_4442,N_4559);
and U4642 (N_4642,N_4438,N_4519);
nand U4643 (N_4643,N_4446,N_4590);
xor U4644 (N_4644,N_4469,N_4434);
nand U4645 (N_4645,N_4432,N_4576);
or U4646 (N_4646,N_4402,N_4539);
nand U4647 (N_4647,N_4400,N_4405);
nand U4648 (N_4648,N_4440,N_4512);
nand U4649 (N_4649,N_4552,N_4535);
and U4650 (N_4650,N_4476,N_4496);
or U4651 (N_4651,N_4532,N_4514);
and U4652 (N_4652,N_4448,N_4534);
and U4653 (N_4653,N_4423,N_4435);
nor U4654 (N_4654,N_4577,N_4418);
nand U4655 (N_4655,N_4470,N_4483);
nand U4656 (N_4656,N_4460,N_4433);
or U4657 (N_4657,N_4561,N_4485);
nor U4658 (N_4658,N_4410,N_4551);
or U4659 (N_4659,N_4502,N_4595);
and U4660 (N_4660,N_4416,N_4566);
xor U4661 (N_4661,N_4415,N_4531);
xor U4662 (N_4662,N_4526,N_4412);
or U4663 (N_4663,N_4563,N_4570);
or U4664 (N_4664,N_4413,N_4456);
nand U4665 (N_4665,N_4597,N_4599);
nor U4666 (N_4666,N_4467,N_4473);
nor U4667 (N_4667,N_4484,N_4584);
or U4668 (N_4668,N_4540,N_4449);
nand U4669 (N_4669,N_4588,N_4444);
or U4670 (N_4670,N_4515,N_4408);
or U4671 (N_4671,N_4574,N_4510);
or U4672 (N_4672,N_4550,N_4428);
nand U4673 (N_4673,N_4548,N_4463);
or U4674 (N_4674,N_4582,N_4487);
or U4675 (N_4675,N_4580,N_4407);
and U4676 (N_4676,N_4477,N_4575);
nor U4677 (N_4677,N_4431,N_4455);
xnor U4678 (N_4678,N_4565,N_4501);
nand U4679 (N_4679,N_4509,N_4491);
and U4680 (N_4680,N_4482,N_4419);
or U4681 (N_4681,N_4592,N_4480);
or U4682 (N_4682,N_4479,N_4404);
and U4683 (N_4683,N_4596,N_4520);
or U4684 (N_4684,N_4518,N_4572);
and U4685 (N_4685,N_4553,N_4430);
and U4686 (N_4686,N_4591,N_4521);
xnor U4687 (N_4687,N_4544,N_4523);
nand U4688 (N_4688,N_4486,N_4508);
and U4689 (N_4689,N_4414,N_4545);
nand U4690 (N_4690,N_4500,N_4457);
xor U4691 (N_4691,N_4589,N_4406);
and U4692 (N_4692,N_4429,N_4524);
nand U4693 (N_4693,N_4506,N_4464);
xor U4694 (N_4694,N_4558,N_4488);
nand U4695 (N_4695,N_4578,N_4453);
nor U4696 (N_4696,N_4424,N_4441);
and U4697 (N_4697,N_4454,N_4573);
and U4698 (N_4698,N_4522,N_4445);
xor U4699 (N_4699,N_4511,N_4504);
xnor U4700 (N_4700,N_4575,N_4537);
nor U4701 (N_4701,N_4463,N_4593);
or U4702 (N_4702,N_4505,N_4453);
xor U4703 (N_4703,N_4474,N_4476);
and U4704 (N_4704,N_4512,N_4422);
and U4705 (N_4705,N_4567,N_4470);
nor U4706 (N_4706,N_4474,N_4415);
nor U4707 (N_4707,N_4442,N_4434);
or U4708 (N_4708,N_4544,N_4413);
nand U4709 (N_4709,N_4555,N_4566);
xnor U4710 (N_4710,N_4595,N_4590);
or U4711 (N_4711,N_4411,N_4595);
nand U4712 (N_4712,N_4509,N_4472);
nand U4713 (N_4713,N_4456,N_4447);
nand U4714 (N_4714,N_4401,N_4535);
nor U4715 (N_4715,N_4533,N_4442);
nand U4716 (N_4716,N_4567,N_4518);
nor U4717 (N_4717,N_4599,N_4400);
nor U4718 (N_4718,N_4416,N_4579);
xnor U4719 (N_4719,N_4438,N_4454);
or U4720 (N_4720,N_4434,N_4536);
and U4721 (N_4721,N_4517,N_4452);
or U4722 (N_4722,N_4409,N_4424);
nor U4723 (N_4723,N_4469,N_4560);
xnor U4724 (N_4724,N_4476,N_4482);
or U4725 (N_4725,N_4462,N_4417);
nor U4726 (N_4726,N_4530,N_4591);
and U4727 (N_4727,N_4509,N_4429);
and U4728 (N_4728,N_4583,N_4569);
or U4729 (N_4729,N_4590,N_4484);
or U4730 (N_4730,N_4504,N_4484);
nor U4731 (N_4731,N_4532,N_4585);
and U4732 (N_4732,N_4435,N_4418);
nor U4733 (N_4733,N_4482,N_4582);
xor U4734 (N_4734,N_4411,N_4544);
xnor U4735 (N_4735,N_4449,N_4413);
nor U4736 (N_4736,N_4461,N_4557);
nor U4737 (N_4737,N_4504,N_4475);
xnor U4738 (N_4738,N_4472,N_4406);
xnor U4739 (N_4739,N_4401,N_4522);
nor U4740 (N_4740,N_4480,N_4504);
xor U4741 (N_4741,N_4591,N_4422);
or U4742 (N_4742,N_4486,N_4589);
nand U4743 (N_4743,N_4440,N_4470);
xnor U4744 (N_4744,N_4403,N_4520);
nor U4745 (N_4745,N_4420,N_4509);
nor U4746 (N_4746,N_4471,N_4502);
xnor U4747 (N_4747,N_4490,N_4421);
nor U4748 (N_4748,N_4589,N_4447);
nand U4749 (N_4749,N_4469,N_4473);
nand U4750 (N_4750,N_4499,N_4595);
and U4751 (N_4751,N_4525,N_4547);
nor U4752 (N_4752,N_4563,N_4546);
xnor U4753 (N_4753,N_4508,N_4547);
xor U4754 (N_4754,N_4464,N_4517);
and U4755 (N_4755,N_4450,N_4471);
and U4756 (N_4756,N_4479,N_4595);
and U4757 (N_4757,N_4424,N_4522);
nand U4758 (N_4758,N_4496,N_4502);
nor U4759 (N_4759,N_4530,N_4482);
nor U4760 (N_4760,N_4596,N_4467);
nand U4761 (N_4761,N_4538,N_4568);
nand U4762 (N_4762,N_4484,N_4511);
nor U4763 (N_4763,N_4455,N_4404);
and U4764 (N_4764,N_4414,N_4510);
and U4765 (N_4765,N_4458,N_4450);
or U4766 (N_4766,N_4482,N_4510);
xor U4767 (N_4767,N_4461,N_4582);
or U4768 (N_4768,N_4526,N_4538);
nor U4769 (N_4769,N_4405,N_4539);
nor U4770 (N_4770,N_4597,N_4506);
nand U4771 (N_4771,N_4562,N_4455);
xor U4772 (N_4772,N_4424,N_4586);
xor U4773 (N_4773,N_4558,N_4536);
and U4774 (N_4774,N_4560,N_4414);
nor U4775 (N_4775,N_4400,N_4518);
nor U4776 (N_4776,N_4424,N_4489);
xnor U4777 (N_4777,N_4594,N_4467);
or U4778 (N_4778,N_4566,N_4453);
or U4779 (N_4779,N_4476,N_4418);
nor U4780 (N_4780,N_4585,N_4445);
and U4781 (N_4781,N_4575,N_4597);
and U4782 (N_4782,N_4498,N_4460);
and U4783 (N_4783,N_4456,N_4503);
and U4784 (N_4784,N_4533,N_4458);
xnor U4785 (N_4785,N_4440,N_4467);
and U4786 (N_4786,N_4520,N_4427);
and U4787 (N_4787,N_4547,N_4553);
nand U4788 (N_4788,N_4575,N_4503);
nor U4789 (N_4789,N_4492,N_4517);
and U4790 (N_4790,N_4529,N_4458);
or U4791 (N_4791,N_4413,N_4586);
or U4792 (N_4792,N_4544,N_4451);
nand U4793 (N_4793,N_4407,N_4421);
or U4794 (N_4794,N_4402,N_4548);
nor U4795 (N_4795,N_4501,N_4522);
xor U4796 (N_4796,N_4536,N_4465);
nor U4797 (N_4797,N_4550,N_4409);
xnor U4798 (N_4798,N_4580,N_4510);
nand U4799 (N_4799,N_4563,N_4450);
xor U4800 (N_4800,N_4715,N_4699);
and U4801 (N_4801,N_4700,N_4749);
xnor U4802 (N_4802,N_4775,N_4799);
or U4803 (N_4803,N_4671,N_4609);
nor U4804 (N_4804,N_4790,N_4618);
nand U4805 (N_4805,N_4777,N_4630);
nor U4806 (N_4806,N_4631,N_4744);
xnor U4807 (N_4807,N_4607,N_4642);
or U4808 (N_4808,N_4745,N_4623);
and U4809 (N_4809,N_4622,N_4606);
nor U4810 (N_4810,N_4646,N_4663);
nor U4811 (N_4811,N_4698,N_4774);
nor U4812 (N_4812,N_4685,N_4641);
nand U4813 (N_4813,N_4769,N_4668);
nor U4814 (N_4814,N_4713,N_4649);
nand U4815 (N_4815,N_4677,N_4759);
nand U4816 (N_4816,N_4683,N_4706);
nor U4817 (N_4817,N_4637,N_4746);
and U4818 (N_4818,N_4751,N_4690);
nor U4819 (N_4819,N_4718,N_4738);
nand U4820 (N_4820,N_4610,N_4714);
nand U4821 (N_4821,N_4648,N_4757);
or U4822 (N_4822,N_4786,N_4734);
and U4823 (N_4823,N_4693,N_4779);
xor U4824 (N_4824,N_4628,N_4695);
nand U4825 (N_4825,N_4652,N_4662);
or U4826 (N_4826,N_4711,N_4621);
nor U4827 (N_4827,N_4608,N_4666);
nor U4828 (N_4828,N_4735,N_4710);
xor U4829 (N_4829,N_4686,N_4747);
or U4830 (N_4830,N_4627,N_4721);
or U4831 (N_4831,N_4616,N_4673);
xnor U4832 (N_4832,N_4687,N_4697);
and U4833 (N_4833,N_4667,N_4740);
xor U4834 (N_4834,N_4764,N_4602);
or U4835 (N_4835,N_4682,N_4741);
xor U4836 (N_4836,N_4678,N_4692);
xor U4837 (N_4837,N_4771,N_4742);
xnor U4838 (N_4838,N_4674,N_4719);
nand U4839 (N_4839,N_4708,N_4725);
or U4840 (N_4840,N_4696,N_4679);
nor U4841 (N_4841,N_4644,N_4676);
or U4842 (N_4842,N_4611,N_4773);
xor U4843 (N_4843,N_4636,N_4617);
xnor U4844 (N_4844,N_4707,N_4785);
nor U4845 (N_4845,N_4780,N_4643);
nor U4846 (N_4846,N_4659,N_4615);
xnor U4847 (N_4847,N_4796,N_4728);
or U4848 (N_4848,N_4655,N_4691);
nand U4849 (N_4849,N_4654,N_4603);
nand U4850 (N_4850,N_4752,N_4704);
nand U4851 (N_4851,N_4753,N_4722);
or U4852 (N_4852,N_4781,N_4614);
xor U4853 (N_4853,N_4772,N_4716);
or U4854 (N_4854,N_4689,N_4723);
and U4855 (N_4855,N_4684,N_4656);
nor U4856 (N_4856,N_4776,N_4768);
or U4857 (N_4857,N_4797,N_4794);
and U4858 (N_4858,N_4755,N_4733);
and U4859 (N_4859,N_4795,N_4660);
or U4860 (N_4860,N_4680,N_4743);
and U4861 (N_4861,N_4625,N_4653);
nand U4862 (N_4862,N_4760,N_4657);
nand U4863 (N_4863,N_4635,N_4709);
and U4864 (N_4864,N_4729,N_4737);
xor U4865 (N_4865,N_4720,N_4748);
or U4866 (N_4866,N_4633,N_4758);
and U4867 (N_4867,N_4702,N_4640);
nand U4868 (N_4868,N_4754,N_4750);
xnor U4869 (N_4869,N_4767,N_4626);
nor U4870 (N_4870,N_4634,N_4600);
nor U4871 (N_4871,N_4647,N_4724);
nand U4872 (N_4872,N_4792,N_4661);
and U4873 (N_4873,N_4739,N_4778);
and U4874 (N_4874,N_4620,N_4730);
or U4875 (N_4875,N_4761,N_4782);
and U4876 (N_4876,N_4613,N_4669);
nor U4877 (N_4877,N_4784,N_4670);
nor U4878 (N_4878,N_4766,N_4675);
nand U4879 (N_4879,N_4701,N_4732);
nor U4880 (N_4880,N_4639,N_4717);
or U4881 (N_4881,N_4601,N_4705);
nand U4882 (N_4882,N_4756,N_4783);
xnor U4883 (N_4883,N_4694,N_4665);
or U4884 (N_4884,N_4798,N_4651);
or U4885 (N_4885,N_4789,N_4672);
xor U4886 (N_4886,N_4765,N_4787);
or U4887 (N_4887,N_4650,N_4726);
and U4888 (N_4888,N_4791,N_4612);
xor U4889 (N_4889,N_4762,N_4664);
nand U4890 (N_4890,N_4731,N_4703);
nor U4891 (N_4891,N_4788,N_4605);
or U4892 (N_4892,N_4770,N_4619);
and U4893 (N_4893,N_4624,N_4793);
or U4894 (N_4894,N_4712,N_4604);
xnor U4895 (N_4895,N_4629,N_4763);
and U4896 (N_4896,N_4658,N_4638);
xor U4897 (N_4897,N_4632,N_4688);
nor U4898 (N_4898,N_4727,N_4736);
or U4899 (N_4899,N_4645,N_4681);
nand U4900 (N_4900,N_4739,N_4630);
nor U4901 (N_4901,N_4733,N_4667);
and U4902 (N_4902,N_4637,N_4620);
nor U4903 (N_4903,N_4765,N_4614);
nand U4904 (N_4904,N_4689,N_4725);
xor U4905 (N_4905,N_4700,N_4710);
or U4906 (N_4906,N_4632,N_4796);
nand U4907 (N_4907,N_4753,N_4621);
xnor U4908 (N_4908,N_4601,N_4790);
nor U4909 (N_4909,N_4768,N_4710);
xnor U4910 (N_4910,N_4749,N_4649);
or U4911 (N_4911,N_4684,N_4615);
nand U4912 (N_4912,N_4722,N_4735);
and U4913 (N_4913,N_4659,N_4694);
or U4914 (N_4914,N_4708,N_4731);
and U4915 (N_4915,N_4762,N_4680);
and U4916 (N_4916,N_4778,N_4771);
xor U4917 (N_4917,N_4737,N_4777);
xnor U4918 (N_4918,N_4692,N_4774);
nand U4919 (N_4919,N_4745,N_4614);
nand U4920 (N_4920,N_4685,N_4767);
nor U4921 (N_4921,N_4723,N_4753);
and U4922 (N_4922,N_4737,N_4683);
and U4923 (N_4923,N_4653,N_4795);
nand U4924 (N_4924,N_4756,N_4675);
nand U4925 (N_4925,N_4681,N_4677);
xnor U4926 (N_4926,N_4713,N_4651);
or U4927 (N_4927,N_4727,N_4753);
or U4928 (N_4928,N_4701,N_4673);
and U4929 (N_4929,N_4738,N_4657);
or U4930 (N_4930,N_4602,N_4715);
nor U4931 (N_4931,N_4715,N_4773);
xnor U4932 (N_4932,N_4639,N_4741);
nand U4933 (N_4933,N_4688,N_4692);
xor U4934 (N_4934,N_4787,N_4683);
and U4935 (N_4935,N_4605,N_4674);
xnor U4936 (N_4936,N_4659,N_4628);
and U4937 (N_4937,N_4643,N_4700);
and U4938 (N_4938,N_4763,N_4694);
nand U4939 (N_4939,N_4672,N_4702);
and U4940 (N_4940,N_4784,N_4723);
xor U4941 (N_4941,N_4763,N_4744);
nor U4942 (N_4942,N_4764,N_4672);
nor U4943 (N_4943,N_4706,N_4714);
nor U4944 (N_4944,N_4767,N_4707);
and U4945 (N_4945,N_4777,N_4680);
nor U4946 (N_4946,N_4620,N_4756);
or U4947 (N_4947,N_4630,N_4652);
and U4948 (N_4948,N_4645,N_4659);
nor U4949 (N_4949,N_4690,N_4695);
and U4950 (N_4950,N_4786,N_4735);
and U4951 (N_4951,N_4606,N_4779);
nor U4952 (N_4952,N_4788,N_4713);
or U4953 (N_4953,N_4795,N_4610);
and U4954 (N_4954,N_4713,N_4766);
xnor U4955 (N_4955,N_4714,N_4717);
and U4956 (N_4956,N_4682,N_4774);
nor U4957 (N_4957,N_4601,N_4637);
nand U4958 (N_4958,N_4765,N_4677);
and U4959 (N_4959,N_4627,N_4667);
nand U4960 (N_4960,N_4639,N_4703);
nor U4961 (N_4961,N_4702,N_4696);
nand U4962 (N_4962,N_4763,N_4716);
nand U4963 (N_4963,N_4632,N_4690);
and U4964 (N_4964,N_4680,N_4706);
nor U4965 (N_4965,N_4749,N_4763);
or U4966 (N_4966,N_4681,N_4769);
xnor U4967 (N_4967,N_4768,N_4753);
xor U4968 (N_4968,N_4678,N_4677);
xnor U4969 (N_4969,N_4717,N_4675);
nor U4970 (N_4970,N_4700,N_4673);
or U4971 (N_4971,N_4705,N_4783);
and U4972 (N_4972,N_4699,N_4793);
and U4973 (N_4973,N_4606,N_4623);
or U4974 (N_4974,N_4636,N_4698);
or U4975 (N_4975,N_4635,N_4726);
nand U4976 (N_4976,N_4707,N_4730);
nor U4977 (N_4977,N_4782,N_4723);
and U4978 (N_4978,N_4648,N_4786);
xnor U4979 (N_4979,N_4652,N_4685);
nand U4980 (N_4980,N_4767,N_4637);
or U4981 (N_4981,N_4773,N_4628);
or U4982 (N_4982,N_4741,N_4758);
nor U4983 (N_4983,N_4706,N_4684);
or U4984 (N_4984,N_4689,N_4691);
nand U4985 (N_4985,N_4769,N_4658);
nand U4986 (N_4986,N_4659,N_4795);
nand U4987 (N_4987,N_4754,N_4622);
and U4988 (N_4988,N_4771,N_4748);
or U4989 (N_4989,N_4678,N_4606);
nand U4990 (N_4990,N_4797,N_4793);
and U4991 (N_4991,N_4735,N_4720);
or U4992 (N_4992,N_4710,N_4704);
and U4993 (N_4993,N_4787,N_4646);
and U4994 (N_4994,N_4749,N_4778);
and U4995 (N_4995,N_4720,N_4728);
nand U4996 (N_4996,N_4683,N_4752);
nand U4997 (N_4997,N_4693,N_4704);
nor U4998 (N_4998,N_4716,N_4646);
or U4999 (N_4999,N_4734,N_4685);
xnor U5000 (N_5000,N_4861,N_4964);
xnor U5001 (N_5001,N_4983,N_4841);
or U5002 (N_5002,N_4806,N_4801);
nand U5003 (N_5003,N_4954,N_4869);
xnor U5004 (N_5004,N_4895,N_4957);
or U5005 (N_5005,N_4909,N_4887);
or U5006 (N_5006,N_4831,N_4902);
and U5007 (N_5007,N_4838,N_4808);
or U5008 (N_5008,N_4811,N_4935);
and U5009 (N_5009,N_4839,N_4804);
xnor U5010 (N_5010,N_4810,N_4953);
xnor U5011 (N_5011,N_4986,N_4949);
and U5012 (N_5012,N_4980,N_4930);
or U5013 (N_5013,N_4842,N_4919);
nor U5014 (N_5014,N_4928,N_4982);
nand U5015 (N_5015,N_4945,N_4950);
xor U5016 (N_5016,N_4884,N_4888);
or U5017 (N_5017,N_4819,N_4933);
and U5018 (N_5018,N_4815,N_4875);
xnor U5019 (N_5019,N_4860,N_4901);
xor U5020 (N_5020,N_4961,N_4971);
nor U5021 (N_5021,N_4824,N_4833);
nor U5022 (N_5022,N_4886,N_4959);
xor U5023 (N_5023,N_4891,N_4898);
nor U5024 (N_5024,N_4848,N_4876);
nand U5025 (N_5025,N_4904,N_4962);
xor U5026 (N_5026,N_4994,N_4881);
nand U5027 (N_5027,N_4927,N_4958);
nor U5028 (N_5028,N_4979,N_4821);
or U5029 (N_5029,N_4925,N_4834);
nand U5030 (N_5030,N_4952,N_4846);
xor U5031 (N_5031,N_4936,N_4939);
nand U5032 (N_5032,N_4974,N_4987);
nor U5033 (N_5033,N_4870,N_4803);
or U5034 (N_5034,N_4931,N_4865);
or U5035 (N_5035,N_4911,N_4934);
or U5036 (N_5036,N_4910,N_4960);
nor U5037 (N_5037,N_4997,N_4890);
xor U5038 (N_5038,N_4867,N_4868);
and U5039 (N_5039,N_4857,N_4832);
xor U5040 (N_5040,N_4844,N_4991);
nor U5041 (N_5041,N_4829,N_4995);
nand U5042 (N_5042,N_4929,N_4955);
nand U5043 (N_5043,N_4851,N_4858);
xor U5044 (N_5044,N_4800,N_4866);
and U5045 (N_5045,N_4988,N_4826);
or U5046 (N_5046,N_4940,N_4921);
and U5047 (N_5047,N_4996,N_4863);
and U5048 (N_5048,N_4873,N_4981);
nor U5049 (N_5049,N_4847,N_4913);
nor U5050 (N_5050,N_4918,N_4874);
nand U5051 (N_5051,N_4802,N_4809);
or U5052 (N_5052,N_4830,N_4855);
or U5053 (N_5053,N_4947,N_4926);
or U5054 (N_5054,N_4879,N_4906);
xor U5055 (N_5055,N_4818,N_4938);
nand U5056 (N_5056,N_4896,N_4862);
nand U5057 (N_5057,N_4893,N_4812);
and U5058 (N_5058,N_4871,N_4817);
nor U5059 (N_5059,N_4880,N_4963);
and U5060 (N_5060,N_4970,N_4903);
and U5061 (N_5061,N_4859,N_4828);
and U5062 (N_5062,N_4977,N_4998);
nand U5063 (N_5063,N_4942,N_4882);
nand U5064 (N_5064,N_4856,N_4992);
nor U5065 (N_5065,N_4976,N_4984);
nand U5066 (N_5066,N_4816,N_4968);
nor U5067 (N_5067,N_4972,N_4840);
nand U5068 (N_5068,N_4822,N_4897);
and U5069 (N_5069,N_4877,N_4924);
nor U5070 (N_5070,N_4907,N_4892);
nand U5071 (N_5071,N_4985,N_4894);
nor U5072 (N_5072,N_4989,N_4843);
and U5073 (N_5073,N_4975,N_4872);
nor U5074 (N_5074,N_4946,N_4937);
and U5075 (N_5075,N_4845,N_4864);
nand U5076 (N_5076,N_4827,N_4967);
and U5077 (N_5077,N_4965,N_4923);
xor U5078 (N_5078,N_4823,N_4966);
nor U5079 (N_5079,N_4993,N_4956);
or U5080 (N_5080,N_4999,N_4948);
or U5081 (N_5081,N_4969,N_4820);
xnor U5082 (N_5082,N_4978,N_4932);
xnor U5083 (N_5083,N_4922,N_4912);
nor U5084 (N_5084,N_4900,N_4916);
xnor U5085 (N_5085,N_4805,N_4990);
nand U5086 (N_5086,N_4853,N_4889);
nor U5087 (N_5087,N_4849,N_4899);
or U5088 (N_5088,N_4941,N_4883);
xnor U5089 (N_5089,N_4825,N_4973);
xnor U5090 (N_5090,N_4908,N_4944);
and U5091 (N_5091,N_4854,N_4905);
nor U5092 (N_5092,N_4878,N_4885);
and U5093 (N_5093,N_4813,N_4836);
nand U5094 (N_5094,N_4915,N_4814);
nor U5095 (N_5095,N_4835,N_4951);
nor U5096 (N_5096,N_4852,N_4807);
or U5097 (N_5097,N_4943,N_4850);
or U5098 (N_5098,N_4837,N_4920);
or U5099 (N_5099,N_4917,N_4914);
nand U5100 (N_5100,N_4825,N_4832);
nor U5101 (N_5101,N_4941,N_4828);
nand U5102 (N_5102,N_4926,N_4934);
and U5103 (N_5103,N_4942,N_4940);
or U5104 (N_5104,N_4895,N_4874);
nand U5105 (N_5105,N_4968,N_4830);
or U5106 (N_5106,N_4895,N_4850);
nor U5107 (N_5107,N_4866,N_4849);
nand U5108 (N_5108,N_4890,N_4906);
nand U5109 (N_5109,N_4998,N_4941);
xor U5110 (N_5110,N_4877,N_4839);
nor U5111 (N_5111,N_4806,N_4892);
xor U5112 (N_5112,N_4873,N_4953);
xnor U5113 (N_5113,N_4908,N_4886);
and U5114 (N_5114,N_4960,N_4984);
and U5115 (N_5115,N_4951,N_4984);
or U5116 (N_5116,N_4807,N_4883);
nor U5117 (N_5117,N_4894,N_4810);
nor U5118 (N_5118,N_4949,N_4859);
or U5119 (N_5119,N_4944,N_4927);
nand U5120 (N_5120,N_4996,N_4978);
xor U5121 (N_5121,N_4890,N_4935);
nor U5122 (N_5122,N_4893,N_4843);
and U5123 (N_5123,N_4955,N_4961);
nand U5124 (N_5124,N_4930,N_4904);
xnor U5125 (N_5125,N_4809,N_4999);
xnor U5126 (N_5126,N_4964,N_4889);
nand U5127 (N_5127,N_4970,N_4929);
or U5128 (N_5128,N_4991,N_4921);
and U5129 (N_5129,N_4861,N_4852);
nand U5130 (N_5130,N_4817,N_4835);
and U5131 (N_5131,N_4994,N_4900);
or U5132 (N_5132,N_4873,N_4995);
and U5133 (N_5133,N_4896,N_4844);
nand U5134 (N_5134,N_4974,N_4983);
nor U5135 (N_5135,N_4857,N_4843);
nor U5136 (N_5136,N_4947,N_4839);
and U5137 (N_5137,N_4883,N_4993);
xor U5138 (N_5138,N_4919,N_4848);
and U5139 (N_5139,N_4906,N_4976);
xnor U5140 (N_5140,N_4856,N_4803);
xnor U5141 (N_5141,N_4967,N_4940);
or U5142 (N_5142,N_4985,N_4976);
and U5143 (N_5143,N_4892,N_4983);
nand U5144 (N_5144,N_4937,N_4868);
xnor U5145 (N_5145,N_4942,N_4845);
xor U5146 (N_5146,N_4920,N_4927);
nor U5147 (N_5147,N_4885,N_4981);
nand U5148 (N_5148,N_4994,N_4879);
and U5149 (N_5149,N_4904,N_4809);
or U5150 (N_5150,N_4832,N_4978);
nor U5151 (N_5151,N_4859,N_4838);
and U5152 (N_5152,N_4854,N_4829);
and U5153 (N_5153,N_4857,N_4825);
and U5154 (N_5154,N_4867,N_4936);
or U5155 (N_5155,N_4970,N_4947);
nor U5156 (N_5156,N_4807,N_4967);
nand U5157 (N_5157,N_4938,N_4957);
and U5158 (N_5158,N_4964,N_4973);
and U5159 (N_5159,N_4914,N_4987);
nor U5160 (N_5160,N_4913,N_4959);
or U5161 (N_5161,N_4930,N_4822);
nand U5162 (N_5162,N_4896,N_4929);
and U5163 (N_5163,N_4941,N_4970);
and U5164 (N_5164,N_4923,N_4832);
nand U5165 (N_5165,N_4973,N_4829);
and U5166 (N_5166,N_4967,N_4981);
or U5167 (N_5167,N_4868,N_4825);
nand U5168 (N_5168,N_4801,N_4920);
nand U5169 (N_5169,N_4900,N_4847);
and U5170 (N_5170,N_4834,N_4990);
nand U5171 (N_5171,N_4987,N_4860);
nand U5172 (N_5172,N_4840,N_4977);
or U5173 (N_5173,N_4981,N_4827);
and U5174 (N_5174,N_4919,N_4840);
nand U5175 (N_5175,N_4977,N_4963);
nor U5176 (N_5176,N_4892,N_4901);
nand U5177 (N_5177,N_4931,N_4886);
nor U5178 (N_5178,N_4892,N_4838);
nand U5179 (N_5179,N_4951,N_4973);
nor U5180 (N_5180,N_4984,N_4892);
and U5181 (N_5181,N_4803,N_4836);
nand U5182 (N_5182,N_4909,N_4936);
nor U5183 (N_5183,N_4933,N_4861);
and U5184 (N_5184,N_4940,N_4891);
nand U5185 (N_5185,N_4996,N_4909);
and U5186 (N_5186,N_4850,N_4852);
xnor U5187 (N_5187,N_4819,N_4910);
nor U5188 (N_5188,N_4957,N_4986);
or U5189 (N_5189,N_4812,N_4835);
nor U5190 (N_5190,N_4995,N_4973);
xnor U5191 (N_5191,N_4901,N_4999);
nor U5192 (N_5192,N_4855,N_4895);
nor U5193 (N_5193,N_4936,N_4833);
xor U5194 (N_5194,N_4894,N_4893);
and U5195 (N_5195,N_4952,N_4975);
xor U5196 (N_5196,N_4859,N_4879);
nor U5197 (N_5197,N_4901,N_4977);
or U5198 (N_5198,N_4938,N_4817);
and U5199 (N_5199,N_4955,N_4952);
or U5200 (N_5200,N_5066,N_5161);
nand U5201 (N_5201,N_5186,N_5012);
and U5202 (N_5202,N_5144,N_5058);
or U5203 (N_5203,N_5117,N_5104);
or U5204 (N_5204,N_5131,N_5015);
or U5205 (N_5205,N_5160,N_5102);
and U5206 (N_5206,N_5106,N_5087);
xnor U5207 (N_5207,N_5014,N_5162);
or U5208 (N_5208,N_5021,N_5056);
and U5209 (N_5209,N_5115,N_5006);
xnor U5210 (N_5210,N_5134,N_5199);
nand U5211 (N_5211,N_5107,N_5089);
or U5212 (N_5212,N_5183,N_5072);
nor U5213 (N_5213,N_5110,N_5039);
and U5214 (N_5214,N_5195,N_5132);
or U5215 (N_5215,N_5119,N_5020);
nand U5216 (N_5216,N_5022,N_5185);
and U5217 (N_5217,N_5179,N_5143);
xnor U5218 (N_5218,N_5044,N_5198);
nor U5219 (N_5219,N_5111,N_5060);
and U5220 (N_5220,N_5136,N_5083);
nor U5221 (N_5221,N_5177,N_5197);
nand U5222 (N_5222,N_5135,N_5045);
nor U5223 (N_5223,N_5137,N_5000);
and U5224 (N_5224,N_5148,N_5105);
nand U5225 (N_5225,N_5079,N_5092);
nor U5226 (N_5226,N_5168,N_5149);
and U5227 (N_5227,N_5171,N_5080);
and U5228 (N_5228,N_5170,N_5184);
nor U5229 (N_5229,N_5049,N_5057);
and U5230 (N_5230,N_5167,N_5155);
and U5231 (N_5231,N_5016,N_5047);
xor U5232 (N_5232,N_5188,N_5126);
nor U5233 (N_5233,N_5048,N_5076);
xnor U5234 (N_5234,N_5031,N_5069);
and U5235 (N_5235,N_5001,N_5068);
nand U5236 (N_5236,N_5026,N_5100);
nand U5237 (N_5237,N_5173,N_5112);
nand U5238 (N_5238,N_5038,N_5011);
or U5239 (N_5239,N_5037,N_5147);
xnor U5240 (N_5240,N_5190,N_5040);
nand U5241 (N_5241,N_5120,N_5055);
or U5242 (N_5242,N_5182,N_5067);
xnor U5243 (N_5243,N_5164,N_5003);
or U5244 (N_5244,N_5029,N_5093);
and U5245 (N_5245,N_5123,N_5024);
nand U5246 (N_5246,N_5151,N_5059);
xnor U5247 (N_5247,N_5146,N_5073);
nor U5248 (N_5248,N_5050,N_5193);
nor U5249 (N_5249,N_5108,N_5007);
xor U5250 (N_5250,N_5094,N_5121);
nor U5251 (N_5251,N_5139,N_5042);
xor U5252 (N_5252,N_5169,N_5172);
nand U5253 (N_5253,N_5174,N_5078);
nand U5254 (N_5254,N_5129,N_5189);
xor U5255 (N_5255,N_5157,N_5036);
and U5256 (N_5256,N_5019,N_5033);
nand U5257 (N_5257,N_5165,N_5192);
nand U5258 (N_5258,N_5158,N_5175);
nand U5259 (N_5259,N_5109,N_5034);
or U5260 (N_5260,N_5181,N_5085);
and U5261 (N_5261,N_5013,N_5023);
or U5262 (N_5262,N_5098,N_5004);
nand U5263 (N_5263,N_5065,N_5027);
or U5264 (N_5264,N_5116,N_5043);
and U5265 (N_5265,N_5070,N_5075);
nor U5266 (N_5266,N_5035,N_5061);
nor U5267 (N_5267,N_5010,N_5051);
nor U5268 (N_5268,N_5071,N_5113);
xnor U5269 (N_5269,N_5009,N_5159);
and U5270 (N_5270,N_5156,N_5145);
and U5271 (N_5271,N_5127,N_5090);
or U5272 (N_5272,N_5088,N_5063);
and U5273 (N_5273,N_5150,N_5142);
nor U5274 (N_5274,N_5082,N_5028);
xor U5275 (N_5275,N_5054,N_5002);
or U5276 (N_5276,N_5141,N_5086);
or U5277 (N_5277,N_5128,N_5095);
and U5278 (N_5278,N_5008,N_5052);
xnor U5279 (N_5279,N_5041,N_5196);
and U5280 (N_5280,N_5018,N_5152);
xor U5281 (N_5281,N_5138,N_5194);
and U5282 (N_5282,N_5084,N_5191);
and U5283 (N_5283,N_5114,N_5091);
or U5284 (N_5284,N_5180,N_5046);
and U5285 (N_5285,N_5154,N_5163);
nand U5286 (N_5286,N_5140,N_5118);
nor U5287 (N_5287,N_5096,N_5005);
nand U5288 (N_5288,N_5166,N_5030);
or U5289 (N_5289,N_5099,N_5178);
nor U5290 (N_5290,N_5017,N_5077);
nor U5291 (N_5291,N_5025,N_5187);
xor U5292 (N_5292,N_5122,N_5130);
nor U5293 (N_5293,N_5062,N_5074);
xnor U5294 (N_5294,N_5125,N_5101);
xnor U5295 (N_5295,N_5133,N_5103);
and U5296 (N_5296,N_5081,N_5032);
nor U5297 (N_5297,N_5053,N_5176);
nand U5298 (N_5298,N_5064,N_5153);
nor U5299 (N_5299,N_5124,N_5097);
xnor U5300 (N_5300,N_5131,N_5036);
or U5301 (N_5301,N_5191,N_5028);
nor U5302 (N_5302,N_5182,N_5119);
and U5303 (N_5303,N_5084,N_5193);
or U5304 (N_5304,N_5003,N_5192);
nor U5305 (N_5305,N_5038,N_5051);
nor U5306 (N_5306,N_5141,N_5188);
and U5307 (N_5307,N_5158,N_5190);
xor U5308 (N_5308,N_5012,N_5018);
and U5309 (N_5309,N_5182,N_5085);
xnor U5310 (N_5310,N_5141,N_5177);
or U5311 (N_5311,N_5162,N_5086);
and U5312 (N_5312,N_5024,N_5001);
nor U5313 (N_5313,N_5000,N_5166);
and U5314 (N_5314,N_5199,N_5077);
nand U5315 (N_5315,N_5011,N_5014);
xor U5316 (N_5316,N_5199,N_5078);
nor U5317 (N_5317,N_5195,N_5147);
nand U5318 (N_5318,N_5004,N_5184);
xor U5319 (N_5319,N_5170,N_5056);
nor U5320 (N_5320,N_5152,N_5134);
xnor U5321 (N_5321,N_5181,N_5186);
nand U5322 (N_5322,N_5157,N_5016);
xnor U5323 (N_5323,N_5032,N_5106);
or U5324 (N_5324,N_5119,N_5011);
nand U5325 (N_5325,N_5031,N_5178);
nand U5326 (N_5326,N_5185,N_5152);
xor U5327 (N_5327,N_5175,N_5039);
nand U5328 (N_5328,N_5041,N_5111);
nand U5329 (N_5329,N_5053,N_5115);
nor U5330 (N_5330,N_5129,N_5086);
xnor U5331 (N_5331,N_5060,N_5134);
or U5332 (N_5332,N_5008,N_5060);
nand U5333 (N_5333,N_5109,N_5166);
nand U5334 (N_5334,N_5173,N_5066);
nand U5335 (N_5335,N_5032,N_5003);
nand U5336 (N_5336,N_5042,N_5120);
xor U5337 (N_5337,N_5085,N_5195);
nor U5338 (N_5338,N_5111,N_5148);
xor U5339 (N_5339,N_5111,N_5153);
and U5340 (N_5340,N_5031,N_5171);
nor U5341 (N_5341,N_5027,N_5139);
nor U5342 (N_5342,N_5119,N_5077);
nor U5343 (N_5343,N_5114,N_5152);
nor U5344 (N_5344,N_5112,N_5122);
or U5345 (N_5345,N_5167,N_5139);
nor U5346 (N_5346,N_5135,N_5008);
nand U5347 (N_5347,N_5076,N_5038);
or U5348 (N_5348,N_5141,N_5139);
and U5349 (N_5349,N_5137,N_5106);
nand U5350 (N_5350,N_5031,N_5043);
nor U5351 (N_5351,N_5157,N_5139);
and U5352 (N_5352,N_5115,N_5122);
xor U5353 (N_5353,N_5199,N_5094);
nor U5354 (N_5354,N_5012,N_5196);
xnor U5355 (N_5355,N_5144,N_5034);
nand U5356 (N_5356,N_5159,N_5095);
or U5357 (N_5357,N_5141,N_5010);
nor U5358 (N_5358,N_5169,N_5001);
nor U5359 (N_5359,N_5068,N_5147);
and U5360 (N_5360,N_5153,N_5184);
xor U5361 (N_5361,N_5083,N_5039);
nor U5362 (N_5362,N_5113,N_5027);
xnor U5363 (N_5363,N_5042,N_5059);
or U5364 (N_5364,N_5042,N_5005);
xnor U5365 (N_5365,N_5072,N_5121);
nor U5366 (N_5366,N_5146,N_5080);
nand U5367 (N_5367,N_5016,N_5051);
nand U5368 (N_5368,N_5042,N_5024);
nor U5369 (N_5369,N_5100,N_5086);
and U5370 (N_5370,N_5044,N_5132);
or U5371 (N_5371,N_5076,N_5062);
nor U5372 (N_5372,N_5051,N_5059);
or U5373 (N_5373,N_5016,N_5111);
xnor U5374 (N_5374,N_5186,N_5083);
nand U5375 (N_5375,N_5057,N_5031);
nand U5376 (N_5376,N_5155,N_5112);
xnor U5377 (N_5377,N_5161,N_5117);
nand U5378 (N_5378,N_5139,N_5030);
and U5379 (N_5379,N_5165,N_5084);
nand U5380 (N_5380,N_5083,N_5161);
and U5381 (N_5381,N_5001,N_5192);
and U5382 (N_5382,N_5175,N_5194);
or U5383 (N_5383,N_5066,N_5152);
and U5384 (N_5384,N_5007,N_5097);
nand U5385 (N_5385,N_5142,N_5002);
nand U5386 (N_5386,N_5144,N_5101);
or U5387 (N_5387,N_5096,N_5028);
nand U5388 (N_5388,N_5019,N_5096);
xor U5389 (N_5389,N_5079,N_5117);
xnor U5390 (N_5390,N_5152,N_5051);
nand U5391 (N_5391,N_5111,N_5094);
or U5392 (N_5392,N_5004,N_5116);
or U5393 (N_5393,N_5163,N_5096);
nand U5394 (N_5394,N_5020,N_5062);
or U5395 (N_5395,N_5037,N_5041);
nand U5396 (N_5396,N_5131,N_5080);
xor U5397 (N_5397,N_5073,N_5066);
or U5398 (N_5398,N_5123,N_5045);
xor U5399 (N_5399,N_5046,N_5170);
nand U5400 (N_5400,N_5292,N_5305);
and U5401 (N_5401,N_5299,N_5208);
nand U5402 (N_5402,N_5355,N_5265);
xor U5403 (N_5403,N_5308,N_5363);
nand U5404 (N_5404,N_5329,N_5200);
nor U5405 (N_5405,N_5237,N_5354);
xnor U5406 (N_5406,N_5277,N_5294);
xnor U5407 (N_5407,N_5370,N_5297);
or U5408 (N_5408,N_5357,N_5252);
xor U5409 (N_5409,N_5359,N_5256);
xnor U5410 (N_5410,N_5219,N_5241);
or U5411 (N_5411,N_5301,N_5242);
nor U5412 (N_5412,N_5215,N_5295);
nor U5413 (N_5413,N_5386,N_5320);
xnor U5414 (N_5414,N_5323,N_5396);
nand U5415 (N_5415,N_5239,N_5206);
nand U5416 (N_5416,N_5293,N_5374);
xnor U5417 (N_5417,N_5300,N_5368);
xnor U5418 (N_5418,N_5321,N_5273);
and U5419 (N_5419,N_5360,N_5207);
nand U5420 (N_5420,N_5254,N_5231);
nand U5421 (N_5421,N_5384,N_5358);
or U5422 (N_5422,N_5266,N_5213);
nand U5423 (N_5423,N_5344,N_5341);
and U5424 (N_5424,N_5204,N_5324);
nand U5425 (N_5425,N_5263,N_5312);
or U5426 (N_5426,N_5269,N_5334);
and U5427 (N_5427,N_5361,N_5303);
xor U5428 (N_5428,N_5391,N_5210);
or U5429 (N_5429,N_5282,N_5283);
xor U5430 (N_5430,N_5365,N_5238);
xnor U5431 (N_5431,N_5319,N_5209);
nor U5432 (N_5432,N_5378,N_5275);
nor U5433 (N_5433,N_5298,N_5349);
xor U5434 (N_5434,N_5388,N_5232);
xnor U5435 (N_5435,N_5271,N_5247);
or U5436 (N_5436,N_5214,N_5398);
nor U5437 (N_5437,N_5267,N_5202);
nand U5438 (N_5438,N_5274,N_5278);
or U5439 (N_5439,N_5333,N_5351);
nor U5440 (N_5440,N_5394,N_5253);
nand U5441 (N_5441,N_5399,N_5234);
and U5442 (N_5442,N_5325,N_5326);
or U5443 (N_5443,N_5330,N_5339);
or U5444 (N_5444,N_5311,N_5211);
or U5445 (N_5445,N_5364,N_5317);
and U5446 (N_5446,N_5286,N_5250);
or U5447 (N_5447,N_5327,N_5217);
nand U5448 (N_5448,N_5362,N_5243);
xnor U5449 (N_5449,N_5379,N_5348);
xor U5450 (N_5450,N_5316,N_5233);
xnor U5451 (N_5451,N_5260,N_5347);
and U5452 (N_5452,N_5350,N_5377);
and U5453 (N_5453,N_5255,N_5389);
or U5454 (N_5454,N_5246,N_5236);
xnor U5455 (N_5455,N_5335,N_5338);
nor U5456 (N_5456,N_5343,N_5262);
xor U5457 (N_5457,N_5235,N_5291);
or U5458 (N_5458,N_5390,N_5385);
xor U5459 (N_5459,N_5284,N_5230);
nor U5460 (N_5460,N_5203,N_5318);
nor U5461 (N_5461,N_5369,N_5337);
nor U5462 (N_5462,N_5220,N_5240);
nand U5463 (N_5463,N_5251,N_5397);
nor U5464 (N_5464,N_5258,N_5395);
xnor U5465 (N_5465,N_5322,N_5229);
nand U5466 (N_5466,N_5222,N_5356);
nor U5467 (N_5467,N_5328,N_5393);
and U5468 (N_5468,N_5218,N_5366);
xnor U5469 (N_5469,N_5310,N_5345);
nor U5470 (N_5470,N_5261,N_5280);
nand U5471 (N_5471,N_5268,N_5287);
nor U5472 (N_5472,N_5221,N_5245);
and U5473 (N_5473,N_5290,N_5281);
and U5474 (N_5474,N_5342,N_5257);
and U5475 (N_5475,N_5307,N_5313);
nor U5476 (N_5476,N_5387,N_5352);
nand U5477 (N_5477,N_5332,N_5340);
nor U5478 (N_5478,N_5372,N_5201);
and U5479 (N_5479,N_5226,N_5383);
or U5480 (N_5480,N_5373,N_5382);
xor U5481 (N_5481,N_5224,N_5270);
xor U5482 (N_5482,N_5248,N_5259);
nand U5483 (N_5483,N_5304,N_5376);
xor U5484 (N_5484,N_5249,N_5288);
and U5485 (N_5485,N_5279,N_5276);
xor U5486 (N_5486,N_5336,N_5392);
nor U5487 (N_5487,N_5380,N_5228);
and U5488 (N_5488,N_5371,N_5272);
and U5489 (N_5489,N_5315,N_5227);
xnor U5490 (N_5490,N_5302,N_5367);
and U5491 (N_5491,N_5212,N_5309);
nand U5492 (N_5492,N_5381,N_5285);
nor U5493 (N_5493,N_5375,N_5346);
and U5494 (N_5494,N_5289,N_5296);
nor U5495 (N_5495,N_5216,N_5225);
and U5496 (N_5496,N_5223,N_5353);
nor U5497 (N_5497,N_5314,N_5244);
and U5498 (N_5498,N_5306,N_5264);
nand U5499 (N_5499,N_5205,N_5331);
nand U5500 (N_5500,N_5393,N_5200);
xnor U5501 (N_5501,N_5300,N_5372);
nand U5502 (N_5502,N_5323,N_5255);
nand U5503 (N_5503,N_5278,N_5201);
nand U5504 (N_5504,N_5294,N_5327);
or U5505 (N_5505,N_5358,N_5372);
xnor U5506 (N_5506,N_5219,N_5295);
or U5507 (N_5507,N_5221,N_5386);
nand U5508 (N_5508,N_5366,N_5318);
or U5509 (N_5509,N_5264,N_5389);
xnor U5510 (N_5510,N_5335,N_5354);
or U5511 (N_5511,N_5216,N_5349);
nor U5512 (N_5512,N_5352,N_5274);
xnor U5513 (N_5513,N_5284,N_5225);
xnor U5514 (N_5514,N_5359,N_5259);
or U5515 (N_5515,N_5234,N_5319);
or U5516 (N_5516,N_5367,N_5245);
nand U5517 (N_5517,N_5263,N_5227);
nand U5518 (N_5518,N_5310,N_5247);
xor U5519 (N_5519,N_5235,N_5224);
xor U5520 (N_5520,N_5253,N_5219);
nor U5521 (N_5521,N_5229,N_5386);
nand U5522 (N_5522,N_5210,N_5340);
nor U5523 (N_5523,N_5208,N_5394);
nor U5524 (N_5524,N_5375,N_5366);
nor U5525 (N_5525,N_5361,N_5201);
and U5526 (N_5526,N_5347,N_5350);
and U5527 (N_5527,N_5397,N_5214);
nor U5528 (N_5528,N_5240,N_5239);
or U5529 (N_5529,N_5366,N_5225);
nor U5530 (N_5530,N_5223,N_5273);
nor U5531 (N_5531,N_5258,N_5376);
nor U5532 (N_5532,N_5211,N_5235);
nand U5533 (N_5533,N_5243,N_5227);
nor U5534 (N_5534,N_5212,N_5396);
nand U5535 (N_5535,N_5222,N_5286);
and U5536 (N_5536,N_5230,N_5256);
nor U5537 (N_5537,N_5305,N_5219);
nand U5538 (N_5538,N_5210,N_5347);
nand U5539 (N_5539,N_5243,N_5387);
and U5540 (N_5540,N_5302,N_5343);
nor U5541 (N_5541,N_5333,N_5379);
and U5542 (N_5542,N_5397,N_5330);
nor U5543 (N_5543,N_5273,N_5360);
xnor U5544 (N_5544,N_5231,N_5380);
nor U5545 (N_5545,N_5325,N_5261);
nor U5546 (N_5546,N_5250,N_5393);
and U5547 (N_5547,N_5217,N_5213);
nand U5548 (N_5548,N_5357,N_5340);
nor U5549 (N_5549,N_5379,N_5294);
nand U5550 (N_5550,N_5347,N_5399);
nand U5551 (N_5551,N_5377,N_5223);
or U5552 (N_5552,N_5312,N_5335);
xnor U5553 (N_5553,N_5243,N_5377);
xnor U5554 (N_5554,N_5318,N_5300);
or U5555 (N_5555,N_5203,N_5347);
nand U5556 (N_5556,N_5270,N_5380);
or U5557 (N_5557,N_5327,N_5277);
nand U5558 (N_5558,N_5320,N_5271);
nor U5559 (N_5559,N_5237,N_5317);
xor U5560 (N_5560,N_5285,N_5360);
xor U5561 (N_5561,N_5357,N_5286);
and U5562 (N_5562,N_5245,N_5388);
and U5563 (N_5563,N_5392,N_5356);
and U5564 (N_5564,N_5216,N_5306);
xnor U5565 (N_5565,N_5394,N_5215);
and U5566 (N_5566,N_5396,N_5306);
xnor U5567 (N_5567,N_5334,N_5389);
or U5568 (N_5568,N_5357,N_5389);
and U5569 (N_5569,N_5324,N_5353);
xnor U5570 (N_5570,N_5303,N_5216);
nand U5571 (N_5571,N_5324,N_5350);
nand U5572 (N_5572,N_5291,N_5278);
nor U5573 (N_5573,N_5287,N_5333);
and U5574 (N_5574,N_5242,N_5336);
nor U5575 (N_5575,N_5333,N_5312);
and U5576 (N_5576,N_5291,N_5362);
nand U5577 (N_5577,N_5329,N_5272);
xnor U5578 (N_5578,N_5214,N_5296);
xor U5579 (N_5579,N_5396,N_5357);
or U5580 (N_5580,N_5238,N_5352);
nand U5581 (N_5581,N_5331,N_5235);
or U5582 (N_5582,N_5351,N_5361);
and U5583 (N_5583,N_5276,N_5278);
or U5584 (N_5584,N_5227,N_5292);
and U5585 (N_5585,N_5369,N_5344);
nor U5586 (N_5586,N_5213,N_5303);
xnor U5587 (N_5587,N_5313,N_5245);
nand U5588 (N_5588,N_5371,N_5233);
nand U5589 (N_5589,N_5322,N_5205);
and U5590 (N_5590,N_5338,N_5200);
nand U5591 (N_5591,N_5235,N_5288);
and U5592 (N_5592,N_5240,N_5345);
or U5593 (N_5593,N_5278,N_5244);
or U5594 (N_5594,N_5359,N_5211);
and U5595 (N_5595,N_5313,N_5239);
nor U5596 (N_5596,N_5346,N_5223);
nor U5597 (N_5597,N_5268,N_5206);
nand U5598 (N_5598,N_5242,N_5200);
nor U5599 (N_5599,N_5337,N_5256);
nand U5600 (N_5600,N_5549,N_5545);
nor U5601 (N_5601,N_5487,N_5574);
nand U5602 (N_5602,N_5445,N_5468);
xor U5603 (N_5603,N_5558,N_5486);
and U5604 (N_5604,N_5570,N_5471);
nor U5605 (N_5605,N_5449,N_5564);
and U5606 (N_5606,N_5478,N_5470);
or U5607 (N_5607,N_5527,N_5506);
nor U5608 (N_5608,N_5481,N_5571);
nor U5609 (N_5609,N_5442,N_5461);
and U5610 (N_5610,N_5436,N_5451);
or U5611 (N_5611,N_5554,N_5524);
nor U5612 (N_5612,N_5443,N_5579);
and U5613 (N_5613,N_5525,N_5419);
or U5614 (N_5614,N_5508,N_5563);
and U5615 (N_5615,N_5575,N_5535);
nor U5616 (N_5616,N_5592,N_5569);
nor U5617 (N_5617,N_5441,N_5502);
nand U5618 (N_5618,N_5400,N_5537);
nor U5619 (N_5619,N_5418,N_5446);
nand U5620 (N_5620,N_5505,N_5476);
and U5621 (N_5621,N_5496,N_5405);
and U5622 (N_5622,N_5521,N_5447);
xor U5623 (N_5623,N_5433,N_5407);
nand U5624 (N_5624,N_5431,N_5528);
xnor U5625 (N_5625,N_5504,N_5541);
or U5626 (N_5626,N_5596,N_5529);
or U5627 (N_5627,N_5517,N_5588);
nand U5628 (N_5628,N_5411,N_5475);
xor U5629 (N_5629,N_5429,N_5493);
and U5630 (N_5630,N_5582,N_5538);
nor U5631 (N_5631,N_5587,N_5408);
or U5632 (N_5632,N_5484,N_5498);
or U5633 (N_5633,N_5514,N_5415);
nand U5634 (N_5634,N_5477,N_5583);
nand U5635 (N_5635,N_5499,N_5580);
nor U5636 (N_5636,N_5594,N_5520);
xor U5637 (N_5637,N_5577,N_5483);
nand U5638 (N_5638,N_5553,N_5454);
xnor U5639 (N_5639,N_5550,N_5465);
xnor U5640 (N_5640,N_5503,N_5507);
nand U5641 (N_5641,N_5469,N_5425);
and U5642 (N_5642,N_5539,N_5547);
nor U5643 (N_5643,N_5556,N_5559);
nand U5644 (N_5644,N_5572,N_5457);
nand U5645 (N_5645,N_5435,N_5422);
and U5646 (N_5646,N_5573,N_5552);
nand U5647 (N_5647,N_5568,N_5463);
nor U5648 (N_5648,N_5488,N_5462);
xor U5649 (N_5649,N_5453,N_5585);
and U5650 (N_5650,N_5417,N_5432);
nor U5651 (N_5651,N_5450,N_5590);
xnor U5652 (N_5652,N_5599,N_5515);
and U5653 (N_5653,N_5482,N_5567);
nor U5654 (N_5654,N_5536,N_5557);
nor U5655 (N_5655,N_5455,N_5413);
nand U5656 (N_5656,N_5452,N_5533);
xnor U5657 (N_5657,N_5509,N_5561);
nand U5658 (N_5658,N_5566,N_5512);
nor U5659 (N_5659,N_5458,N_5534);
or U5660 (N_5660,N_5479,N_5522);
nor U5661 (N_5661,N_5430,N_5597);
and U5662 (N_5662,N_5519,N_5409);
and U5663 (N_5663,N_5560,N_5420);
and U5664 (N_5664,N_5490,N_5555);
xor U5665 (N_5665,N_5434,N_5516);
xnor U5666 (N_5666,N_5466,N_5510);
nand U5667 (N_5667,N_5591,N_5460);
or U5668 (N_5668,N_5403,N_5439);
nor U5669 (N_5669,N_5531,N_5489);
and U5670 (N_5670,N_5424,N_5428);
xor U5671 (N_5671,N_5495,N_5523);
nor U5672 (N_5672,N_5438,N_5401);
xor U5673 (N_5673,N_5480,N_5578);
nor U5674 (N_5674,N_5513,N_5426);
nor U5675 (N_5675,N_5404,N_5402);
nor U5676 (N_5676,N_5530,N_5584);
xnor U5677 (N_5677,N_5542,N_5593);
or U5678 (N_5678,N_5459,N_5444);
or U5679 (N_5679,N_5544,N_5501);
xor U5680 (N_5680,N_5440,N_5456);
or U5681 (N_5681,N_5474,N_5532);
and U5682 (N_5682,N_5586,N_5448);
nand U5683 (N_5683,N_5562,N_5467);
or U5684 (N_5684,N_5497,N_5526);
xor U5685 (N_5685,N_5576,N_5421);
and U5686 (N_5686,N_5473,N_5518);
nand U5687 (N_5687,N_5410,N_5548);
or U5688 (N_5688,N_5427,N_5589);
and U5689 (N_5689,N_5406,N_5412);
or U5690 (N_5690,N_5414,N_5494);
and U5691 (N_5691,N_5492,N_5546);
and U5692 (N_5692,N_5543,N_5472);
or U5693 (N_5693,N_5437,N_5464);
xnor U5694 (N_5694,N_5485,N_5565);
xor U5695 (N_5695,N_5500,N_5423);
xor U5696 (N_5696,N_5598,N_5581);
and U5697 (N_5697,N_5511,N_5491);
nor U5698 (N_5698,N_5595,N_5551);
xor U5699 (N_5699,N_5416,N_5540);
nand U5700 (N_5700,N_5431,N_5582);
nor U5701 (N_5701,N_5528,N_5589);
nor U5702 (N_5702,N_5586,N_5580);
or U5703 (N_5703,N_5565,N_5529);
nor U5704 (N_5704,N_5484,N_5591);
nand U5705 (N_5705,N_5589,N_5548);
and U5706 (N_5706,N_5547,N_5423);
nand U5707 (N_5707,N_5407,N_5453);
xnor U5708 (N_5708,N_5509,N_5422);
or U5709 (N_5709,N_5537,N_5511);
xor U5710 (N_5710,N_5524,N_5400);
and U5711 (N_5711,N_5514,N_5444);
and U5712 (N_5712,N_5404,N_5531);
nand U5713 (N_5713,N_5413,N_5591);
or U5714 (N_5714,N_5441,N_5545);
or U5715 (N_5715,N_5476,N_5562);
xnor U5716 (N_5716,N_5503,N_5560);
xor U5717 (N_5717,N_5418,N_5442);
xor U5718 (N_5718,N_5517,N_5521);
or U5719 (N_5719,N_5596,N_5535);
or U5720 (N_5720,N_5560,N_5483);
xnor U5721 (N_5721,N_5585,N_5423);
or U5722 (N_5722,N_5578,N_5586);
nor U5723 (N_5723,N_5559,N_5561);
and U5724 (N_5724,N_5405,N_5418);
nand U5725 (N_5725,N_5515,N_5591);
nand U5726 (N_5726,N_5599,N_5455);
xor U5727 (N_5727,N_5410,N_5505);
nand U5728 (N_5728,N_5489,N_5419);
or U5729 (N_5729,N_5429,N_5489);
nor U5730 (N_5730,N_5476,N_5441);
xnor U5731 (N_5731,N_5432,N_5550);
nand U5732 (N_5732,N_5589,N_5431);
xor U5733 (N_5733,N_5418,N_5500);
xnor U5734 (N_5734,N_5553,N_5572);
xnor U5735 (N_5735,N_5420,N_5462);
and U5736 (N_5736,N_5412,N_5574);
and U5737 (N_5737,N_5592,N_5531);
or U5738 (N_5738,N_5503,N_5584);
or U5739 (N_5739,N_5516,N_5421);
xnor U5740 (N_5740,N_5532,N_5445);
and U5741 (N_5741,N_5578,N_5556);
nand U5742 (N_5742,N_5408,N_5540);
xnor U5743 (N_5743,N_5591,N_5595);
xor U5744 (N_5744,N_5545,N_5440);
or U5745 (N_5745,N_5479,N_5461);
nor U5746 (N_5746,N_5512,N_5519);
xnor U5747 (N_5747,N_5467,N_5533);
and U5748 (N_5748,N_5439,N_5565);
and U5749 (N_5749,N_5513,N_5494);
nand U5750 (N_5750,N_5406,N_5589);
nor U5751 (N_5751,N_5481,N_5400);
and U5752 (N_5752,N_5556,N_5414);
nor U5753 (N_5753,N_5442,N_5464);
xor U5754 (N_5754,N_5559,N_5596);
nand U5755 (N_5755,N_5570,N_5558);
or U5756 (N_5756,N_5479,N_5557);
xnor U5757 (N_5757,N_5532,N_5564);
or U5758 (N_5758,N_5534,N_5440);
nand U5759 (N_5759,N_5518,N_5545);
xnor U5760 (N_5760,N_5439,N_5487);
nand U5761 (N_5761,N_5569,N_5542);
nand U5762 (N_5762,N_5518,N_5575);
or U5763 (N_5763,N_5536,N_5528);
xor U5764 (N_5764,N_5403,N_5547);
xor U5765 (N_5765,N_5520,N_5422);
nand U5766 (N_5766,N_5520,N_5473);
and U5767 (N_5767,N_5416,N_5553);
xnor U5768 (N_5768,N_5502,N_5454);
xor U5769 (N_5769,N_5573,N_5449);
nor U5770 (N_5770,N_5458,N_5426);
nand U5771 (N_5771,N_5407,N_5590);
and U5772 (N_5772,N_5490,N_5405);
nor U5773 (N_5773,N_5546,N_5477);
and U5774 (N_5774,N_5501,N_5588);
xnor U5775 (N_5775,N_5441,N_5429);
nor U5776 (N_5776,N_5448,N_5442);
or U5777 (N_5777,N_5494,N_5476);
or U5778 (N_5778,N_5592,N_5410);
or U5779 (N_5779,N_5478,N_5444);
and U5780 (N_5780,N_5443,N_5520);
nor U5781 (N_5781,N_5457,N_5574);
xor U5782 (N_5782,N_5434,N_5433);
or U5783 (N_5783,N_5453,N_5422);
and U5784 (N_5784,N_5591,N_5457);
and U5785 (N_5785,N_5530,N_5462);
and U5786 (N_5786,N_5562,N_5528);
nand U5787 (N_5787,N_5435,N_5481);
nand U5788 (N_5788,N_5435,N_5412);
or U5789 (N_5789,N_5501,N_5556);
or U5790 (N_5790,N_5420,N_5489);
or U5791 (N_5791,N_5446,N_5428);
or U5792 (N_5792,N_5583,N_5530);
or U5793 (N_5793,N_5476,N_5447);
or U5794 (N_5794,N_5512,N_5549);
and U5795 (N_5795,N_5564,N_5417);
or U5796 (N_5796,N_5415,N_5550);
nand U5797 (N_5797,N_5513,N_5499);
nor U5798 (N_5798,N_5563,N_5469);
or U5799 (N_5799,N_5512,N_5467);
and U5800 (N_5800,N_5730,N_5682);
nand U5801 (N_5801,N_5789,N_5669);
or U5802 (N_5802,N_5672,N_5668);
nand U5803 (N_5803,N_5770,N_5633);
and U5804 (N_5804,N_5641,N_5745);
nor U5805 (N_5805,N_5796,N_5675);
nand U5806 (N_5806,N_5613,N_5687);
nor U5807 (N_5807,N_5747,N_5765);
nor U5808 (N_5808,N_5772,N_5715);
xor U5809 (N_5809,N_5681,N_5686);
and U5810 (N_5810,N_5695,N_5670);
xnor U5811 (N_5811,N_5746,N_5794);
nand U5812 (N_5812,N_5754,N_5767);
and U5813 (N_5813,N_5766,N_5733);
xnor U5814 (N_5814,N_5724,N_5647);
nor U5815 (N_5815,N_5702,N_5786);
nand U5816 (N_5816,N_5755,N_5777);
nand U5817 (N_5817,N_5607,N_5790);
or U5818 (N_5818,N_5758,N_5763);
or U5819 (N_5819,N_5627,N_5660);
nand U5820 (N_5820,N_5787,N_5707);
nor U5821 (N_5821,N_5750,N_5698);
nor U5822 (N_5822,N_5743,N_5760);
nand U5823 (N_5823,N_5637,N_5601);
and U5824 (N_5824,N_5725,N_5652);
nand U5825 (N_5825,N_5769,N_5700);
nor U5826 (N_5826,N_5634,N_5640);
and U5827 (N_5827,N_5720,N_5781);
nor U5828 (N_5828,N_5731,N_5716);
nand U5829 (N_5829,N_5629,N_5723);
or U5830 (N_5830,N_5775,N_5639);
nand U5831 (N_5831,N_5677,N_5791);
xnor U5832 (N_5832,N_5734,N_5752);
nand U5833 (N_5833,N_5691,N_5737);
nor U5834 (N_5834,N_5728,N_5608);
or U5835 (N_5835,N_5784,N_5751);
xnor U5836 (N_5836,N_5671,N_5719);
and U5837 (N_5837,N_5600,N_5711);
xnor U5838 (N_5838,N_5776,N_5705);
xor U5839 (N_5839,N_5646,N_5757);
xnor U5840 (N_5840,N_5657,N_5604);
and U5841 (N_5841,N_5628,N_5643);
and U5842 (N_5842,N_5611,N_5764);
nand U5843 (N_5843,N_5683,N_5762);
and U5844 (N_5844,N_5727,N_5736);
nand U5845 (N_5845,N_5697,N_5780);
nand U5846 (N_5846,N_5740,N_5678);
or U5847 (N_5847,N_5653,N_5708);
xnor U5848 (N_5848,N_5706,N_5609);
or U5849 (N_5849,N_5696,N_5620);
nand U5850 (N_5850,N_5779,N_5621);
nand U5851 (N_5851,N_5645,N_5717);
nand U5852 (N_5852,N_5605,N_5674);
nand U5853 (N_5853,N_5616,N_5744);
or U5854 (N_5854,N_5713,N_5648);
nor U5855 (N_5855,N_5785,N_5739);
nor U5856 (N_5856,N_5676,N_5666);
nor U5857 (N_5857,N_5735,N_5714);
or U5858 (N_5858,N_5649,N_5632);
nand U5859 (N_5859,N_5679,N_5651);
or U5860 (N_5860,N_5729,N_5658);
and U5861 (N_5861,N_5721,N_5662);
nand U5862 (N_5862,N_5655,N_5704);
nand U5863 (N_5863,N_5756,N_5782);
nor U5864 (N_5864,N_5688,N_5602);
and U5865 (N_5865,N_5783,N_5685);
and U5866 (N_5866,N_5771,N_5699);
nand U5867 (N_5867,N_5689,N_5664);
xor U5868 (N_5868,N_5603,N_5615);
nand U5869 (N_5869,N_5788,N_5774);
or U5870 (N_5870,N_5793,N_5659);
or U5871 (N_5871,N_5654,N_5741);
xor U5872 (N_5872,N_5690,N_5606);
or U5873 (N_5873,N_5625,N_5644);
xor U5874 (N_5874,N_5738,N_5693);
nand U5875 (N_5875,N_5798,N_5619);
nand U5876 (N_5876,N_5701,N_5624);
xnor U5877 (N_5877,N_5795,N_5748);
and U5878 (N_5878,N_5742,N_5692);
xor U5879 (N_5879,N_5665,N_5663);
and U5880 (N_5880,N_5749,N_5631);
nor U5881 (N_5881,N_5710,N_5703);
nand U5882 (N_5882,N_5661,N_5650);
nand U5883 (N_5883,N_5759,N_5684);
nand U5884 (N_5884,N_5726,N_5622);
xor U5885 (N_5885,N_5712,N_5623);
nor U5886 (N_5886,N_5753,N_5638);
or U5887 (N_5887,N_5667,N_5642);
xnor U5888 (N_5888,N_5709,N_5792);
or U5889 (N_5889,N_5732,N_5614);
and U5890 (N_5890,N_5694,N_5618);
nand U5891 (N_5891,N_5656,N_5722);
and U5892 (N_5892,N_5718,N_5761);
nor U5893 (N_5893,N_5680,N_5799);
or U5894 (N_5894,N_5630,N_5635);
or U5895 (N_5895,N_5797,N_5612);
nor U5896 (N_5896,N_5626,N_5773);
nand U5897 (N_5897,N_5610,N_5778);
nand U5898 (N_5898,N_5673,N_5768);
or U5899 (N_5899,N_5636,N_5617);
or U5900 (N_5900,N_5654,N_5642);
nand U5901 (N_5901,N_5784,N_5755);
and U5902 (N_5902,N_5757,N_5611);
nand U5903 (N_5903,N_5657,N_5788);
or U5904 (N_5904,N_5789,N_5622);
nand U5905 (N_5905,N_5689,N_5637);
xor U5906 (N_5906,N_5719,N_5746);
xor U5907 (N_5907,N_5644,N_5613);
xnor U5908 (N_5908,N_5724,N_5783);
xnor U5909 (N_5909,N_5662,N_5794);
nand U5910 (N_5910,N_5722,N_5774);
and U5911 (N_5911,N_5778,N_5740);
xor U5912 (N_5912,N_5684,N_5647);
and U5913 (N_5913,N_5789,N_5627);
and U5914 (N_5914,N_5731,N_5733);
and U5915 (N_5915,N_5677,N_5709);
and U5916 (N_5916,N_5666,N_5689);
and U5917 (N_5917,N_5639,N_5637);
and U5918 (N_5918,N_5773,N_5715);
or U5919 (N_5919,N_5675,N_5779);
xnor U5920 (N_5920,N_5749,N_5767);
nor U5921 (N_5921,N_5632,N_5767);
xnor U5922 (N_5922,N_5743,N_5663);
xor U5923 (N_5923,N_5776,N_5707);
nor U5924 (N_5924,N_5764,N_5695);
or U5925 (N_5925,N_5763,N_5717);
and U5926 (N_5926,N_5642,N_5726);
nand U5927 (N_5927,N_5729,N_5694);
or U5928 (N_5928,N_5702,N_5731);
nor U5929 (N_5929,N_5724,N_5728);
or U5930 (N_5930,N_5655,N_5781);
nor U5931 (N_5931,N_5616,N_5705);
xnor U5932 (N_5932,N_5723,N_5732);
or U5933 (N_5933,N_5709,N_5796);
or U5934 (N_5934,N_5612,N_5684);
and U5935 (N_5935,N_5626,N_5739);
or U5936 (N_5936,N_5695,N_5618);
nor U5937 (N_5937,N_5744,N_5628);
or U5938 (N_5938,N_5773,N_5789);
nand U5939 (N_5939,N_5727,N_5614);
and U5940 (N_5940,N_5618,N_5675);
nand U5941 (N_5941,N_5736,N_5608);
and U5942 (N_5942,N_5795,N_5775);
or U5943 (N_5943,N_5775,N_5671);
nor U5944 (N_5944,N_5606,N_5687);
xor U5945 (N_5945,N_5629,N_5717);
xnor U5946 (N_5946,N_5678,N_5684);
and U5947 (N_5947,N_5732,N_5790);
nand U5948 (N_5948,N_5617,N_5643);
nor U5949 (N_5949,N_5613,N_5641);
nor U5950 (N_5950,N_5702,N_5631);
nor U5951 (N_5951,N_5681,N_5639);
and U5952 (N_5952,N_5782,N_5709);
or U5953 (N_5953,N_5718,N_5778);
nand U5954 (N_5954,N_5766,N_5763);
nor U5955 (N_5955,N_5608,N_5630);
nor U5956 (N_5956,N_5624,N_5667);
nor U5957 (N_5957,N_5602,N_5668);
nand U5958 (N_5958,N_5622,N_5681);
and U5959 (N_5959,N_5715,N_5730);
nor U5960 (N_5960,N_5628,N_5733);
nand U5961 (N_5961,N_5621,N_5774);
nand U5962 (N_5962,N_5678,N_5669);
nand U5963 (N_5963,N_5747,N_5621);
and U5964 (N_5964,N_5668,N_5604);
xor U5965 (N_5965,N_5610,N_5623);
xor U5966 (N_5966,N_5679,N_5615);
xor U5967 (N_5967,N_5760,N_5714);
nand U5968 (N_5968,N_5689,N_5658);
and U5969 (N_5969,N_5790,N_5766);
nor U5970 (N_5970,N_5670,N_5715);
nor U5971 (N_5971,N_5671,N_5777);
xor U5972 (N_5972,N_5771,N_5647);
and U5973 (N_5973,N_5657,N_5760);
xor U5974 (N_5974,N_5689,N_5746);
and U5975 (N_5975,N_5620,N_5643);
and U5976 (N_5976,N_5776,N_5759);
nand U5977 (N_5977,N_5700,N_5777);
or U5978 (N_5978,N_5677,N_5765);
xnor U5979 (N_5979,N_5725,N_5788);
xnor U5980 (N_5980,N_5671,N_5752);
xnor U5981 (N_5981,N_5665,N_5750);
xnor U5982 (N_5982,N_5680,N_5678);
nand U5983 (N_5983,N_5639,N_5755);
nor U5984 (N_5984,N_5677,N_5796);
nand U5985 (N_5985,N_5701,N_5674);
and U5986 (N_5986,N_5770,N_5781);
xnor U5987 (N_5987,N_5716,N_5666);
nand U5988 (N_5988,N_5608,N_5786);
xor U5989 (N_5989,N_5785,N_5618);
nor U5990 (N_5990,N_5667,N_5725);
or U5991 (N_5991,N_5693,N_5620);
xor U5992 (N_5992,N_5791,N_5724);
xor U5993 (N_5993,N_5742,N_5683);
xor U5994 (N_5994,N_5664,N_5785);
or U5995 (N_5995,N_5752,N_5645);
or U5996 (N_5996,N_5664,N_5609);
nor U5997 (N_5997,N_5740,N_5702);
nand U5998 (N_5998,N_5749,N_5751);
nand U5999 (N_5999,N_5666,N_5745);
nand U6000 (N_6000,N_5811,N_5832);
or U6001 (N_6001,N_5884,N_5962);
nand U6002 (N_6002,N_5886,N_5843);
and U6003 (N_6003,N_5831,N_5813);
or U6004 (N_6004,N_5940,N_5863);
nand U6005 (N_6005,N_5878,N_5806);
nand U6006 (N_6006,N_5824,N_5812);
nand U6007 (N_6007,N_5897,N_5972);
xor U6008 (N_6008,N_5872,N_5816);
and U6009 (N_6009,N_5985,N_5921);
nor U6010 (N_6010,N_5866,N_5916);
or U6011 (N_6011,N_5987,N_5818);
and U6012 (N_6012,N_5966,N_5926);
or U6013 (N_6013,N_5906,N_5857);
xor U6014 (N_6014,N_5901,N_5943);
and U6015 (N_6015,N_5977,N_5929);
nand U6016 (N_6016,N_5837,N_5822);
nand U6017 (N_6017,N_5984,N_5991);
nand U6018 (N_6018,N_5868,N_5877);
xor U6019 (N_6019,N_5882,N_5983);
xor U6020 (N_6020,N_5900,N_5969);
and U6021 (N_6021,N_5920,N_5963);
nor U6022 (N_6022,N_5802,N_5941);
xnor U6023 (N_6023,N_5856,N_5980);
xor U6024 (N_6024,N_5883,N_5865);
nand U6025 (N_6025,N_5930,N_5800);
nand U6026 (N_6026,N_5880,N_5989);
nor U6027 (N_6027,N_5892,N_5875);
or U6028 (N_6028,N_5820,N_5905);
or U6029 (N_6029,N_5844,N_5842);
and U6030 (N_6030,N_5952,N_5879);
and U6031 (N_6031,N_5808,N_5815);
and U6032 (N_6032,N_5833,N_5978);
xor U6033 (N_6033,N_5846,N_5829);
nor U6034 (N_6034,N_5814,N_5853);
nand U6035 (N_6035,N_5973,N_5953);
or U6036 (N_6036,N_5986,N_5828);
nand U6037 (N_6037,N_5970,N_5994);
or U6038 (N_6038,N_5888,N_5827);
and U6039 (N_6039,N_5993,N_5890);
and U6040 (N_6040,N_5917,N_5944);
and U6041 (N_6041,N_5976,N_5936);
and U6042 (N_6042,N_5847,N_5912);
or U6043 (N_6043,N_5830,N_5927);
xnor U6044 (N_6044,N_5909,N_5841);
nand U6045 (N_6045,N_5959,N_5988);
nand U6046 (N_6046,N_5967,N_5965);
nand U6047 (N_6047,N_5981,N_5859);
xor U6048 (N_6048,N_5998,N_5861);
xor U6049 (N_6049,N_5975,N_5925);
and U6050 (N_6050,N_5979,N_5948);
nand U6051 (N_6051,N_5937,N_5821);
nor U6052 (N_6052,N_5947,N_5896);
and U6053 (N_6053,N_5955,N_5950);
or U6054 (N_6054,N_5903,N_5982);
nand U6055 (N_6055,N_5838,N_5845);
or U6056 (N_6056,N_5858,N_5922);
or U6057 (N_6057,N_5935,N_5898);
or U6058 (N_6058,N_5915,N_5911);
nand U6059 (N_6059,N_5819,N_5889);
and U6060 (N_6060,N_5893,N_5839);
nor U6061 (N_6061,N_5913,N_5864);
nor U6062 (N_6062,N_5942,N_5971);
and U6063 (N_6063,N_5876,N_5992);
or U6064 (N_6064,N_5885,N_5804);
nand U6065 (N_6065,N_5990,N_5840);
nand U6066 (N_6066,N_5874,N_5958);
nand U6067 (N_6067,N_5891,N_5836);
nand U6068 (N_6068,N_5968,N_5894);
or U6069 (N_6069,N_5803,N_5809);
nor U6070 (N_6070,N_5849,N_5862);
xnor U6071 (N_6071,N_5933,N_5945);
xnor U6072 (N_6072,N_5995,N_5850);
xor U6073 (N_6073,N_5996,N_5873);
nor U6074 (N_6074,N_5960,N_5907);
and U6075 (N_6075,N_5902,N_5825);
and U6076 (N_6076,N_5810,N_5817);
xnor U6077 (N_6077,N_5928,N_5908);
xor U6078 (N_6078,N_5848,N_5854);
or U6079 (N_6079,N_5835,N_5931);
nand U6080 (N_6080,N_5974,N_5910);
nand U6081 (N_6081,N_5881,N_5860);
or U6082 (N_6082,N_5869,N_5914);
nor U6083 (N_6083,N_5855,N_5918);
nand U6084 (N_6084,N_5870,N_5895);
and U6085 (N_6085,N_5919,N_5807);
and U6086 (N_6086,N_5904,N_5934);
nor U6087 (N_6087,N_5887,N_5867);
or U6088 (N_6088,N_5826,N_5946);
or U6089 (N_6089,N_5999,N_5851);
or U6090 (N_6090,N_5852,N_5997);
nor U6091 (N_6091,N_5938,N_5805);
and U6092 (N_6092,N_5871,N_5923);
xor U6093 (N_6093,N_5932,N_5801);
nor U6094 (N_6094,N_5924,N_5951);
and U6095 (N_6095,N_5957,N_5949);
nand U6096 (N_6096,N_5823,N_5961);
xor U6097 (N_6097,N_5939,N_5899);
and U6098 (N_6098,N_5964,N_5834);
nand U6099 (N_6099,N_5956,N_5954);
or U6100 (N_6100,N_5863,N_5999);
nand U6101 (N_6101,N_5872,N_5813);
nor U6102 (N_6102,N_5816,N_5937);
and U6103 (N_6103,N_5874,N_5896);
nand U6104 (N_6104,N_5952,N_5857);
nand U6105 (N_6105,N_5879,N_5805);
and U6106 (N_6106,N_5894,N_5908);
or U6107 (N_6107,N_5956,N_5998);
or U6108 (N_6108,N_5845,N_5977);
xor U6109 (N_6109,N_5886,N_5971);
nor U6110 (N_6110,N_5851,N_5876);
and U6111 (N_6111,N_5952,N_5947);
nand U6112 (N_6112,N_5890,N_5847);
xor U6113 (N_6113,N_5826,N_5889);
nor U6114 (N_6114,N_5933,N_5859);
or U6115 (N_6115,N_5957,N_5940);
xnor U6116 (N_6116,N_5800,N_5948);
xnor U6117 (N_6117,N_5905,N_5936);
or U6118 (N_6118,N_5835,N_5888);
and U6119 (N_6119,N_5864,N_5855);
nor U6120 (N_6120,N_5823,N_5956);
nand U6121 (N_6121,N_5903,N_5964);
and U6122 (N_6122,N_5933,N_5820);
or U6123 (N_6123,N_5860,N_5883);
xnor U6124 (N_6124,N_5850,N_5973);
xnor U6125 (N_6125,N_5982,N_5808);
and U6126 (N_6126,N_5909,N_5961);
nor U6127 (N_6127,N_5959,N_5830);
xor U6128 (N_6128,N_5948,N_5874);
or U6129 (N_6129,N_5923,N_5867);
nand U6130 (N_6130,N_5879,N_5854);
or U6131 (N_6131,N_5928,N_5986);
nor U6132 (N_6132,N_5812,N_5811);
nand U6133 (N_6133,N_5956,N_5900);
or U6134 (N_6134,N_5937,N_5930);
nand U6135 (N_6135,N_5920,N_5880);
nand U6136 (N_6136,N_5834,N_5978);
nand U6137 (N_6137,N_5967,N_5948);
nor U6138 (N_6138,N_5816,N_5925);
and U6139 (N_6139,N_5992,N_5805);
and U6140 (N_6140,N_5892,N_5837);
and U6141 (N_6141,N_5958,N_5844);
nor U6142 (N_6142,N_5889,N_5887);
nor U6143 (N_6143,N_5996,N_5983);
nand U6144 (N_6144,N_5941,N_5803);
xnor U6145 (N_6145,N_5920,N_5820);
nor U6146 (N_6146,N_5919,N_5897);
and U6147 (N_6147,N_5890,N_5820);
nor U6148 (N_6148,N_5862,N_5994);
nand U6149 (N_6149,N_5948,N_5908);
or U6150 (N_6150,N_5909,N_5853);
nor U6151 (N_6151,N_5922,N_5966);
xor U6152 (N_6152,N_5900,N_5809);
or U6153 (N_6153,N_5997,N_5891);
or U6154 (N_6154,N_5982,N_5809);
nor U6155 (N_6155,N_5942,N_5966);
nor U6156 (N_6156,N_5912,N_5988);
nor U6157 (N_6157,N_5850,N_5998);
nor U6158 (N_6158,N_5939,N_5968);
nand U6159 (N_6159,N_5908,N_5851);
nand U6160 (N_6160,N_5866,N_5980);
and U6161 (N_6161,N_5897,N_5827);
or U6162 (N_6162,N_5901,N_5865);
xnor U6163 (N_6163,N_5984,N_5986);
and U6164 (N_6164,N_5969,N_5979);
or U6165 (N_6165,N_5954,N_5828);
xnor U6166 (N_6166,N_5804,N_5830);
xnor U6167 (N_6167,N_5912,N_5977);
or U6168 (N_6168,N_5902,N_5999);
xor U6169 (N_6169,N_5930,N_5811);
nand U6170 (N_6170,N_5857,N_5955);
and U6171 (N_6171,N_5925,N_5924);
nor U6172 (N_6172,N_5832,N_5994);
nor U6173 (N_6173,N_5932,N_5817);
xor U6174 (N_6174,N_5885,N_5957);
nor U6175 (N_6175,N_5850,N_5859);
nand U6176 (N_6176,N_5868,N_5824);
nand U6177 (N_6177,N_5995,N_5820);
nand U6178 (N_6178,N_5813,N_5838);
nand U6179 (N_6179,N_5893,N_5967);
xor U6180 (N_6180,N_5863,N_5847);
and U6181 (N_6181,N_5942,N_5844);
xor U6182 (N_6182,N_5817,N_5966);
nand U6183 (N_6183,N_5994,N_5958);
or U6184 (N_6184,N_5830,N_5982);
nor U6185 (N_6185,N_5851,N_5930);
nand U6186 (N_6186,N_5814,N_5981);
nor U6187 (N_6187,N_5894,N_5981);
nor U6188 (N_6188,N_5811,N_5940);
nor U6189 (N_6189,N_5943,N_5914);
xor U6190 (N_6190,N_5953,N_5801);
or U6191 (N_6191,N_5896,N_5956);
and U6192 (N_6192,N_5881,N_5995);
and U6193 (N_6193,N_5963,N_5889);
and U6194 (N_6194,N_5920,N_5918);
and U6195 (N_6195,N_5978,N_5943);
xor U6196 (N_6196,N_5932,N_5858);
xor U6197 (N_6197,N_5842,N_5995);
nor U6198 (N_6198,N_5933,N_5973);
nand U6199 (N_6199,N_5957,N_5934);
and U6200 (N_6200,N_6025,N_6144);
xor U6201 (N_6201,N_6009,N_6052);
xor U6202 (N_6202,N_6157,N_6090);
and U6203 (N_6203,N_6000,N_6104);
or U6204 (N_6204,N_6139,N_6198);
xnor U6205 (N_6205,N_6190,N_6124);
nor U6206 (N_6206,N_6047,N_6061);
nand U6207 (N_6207,N_6016,N_6014);
and U6208 (N_6208,N_6103,N_6017);
nand U6209 (N_6209,N_6121,N_6147);
xor U6210 (N_6210,N_6087,N_6132);
nor U6211 (N_6211,N_6065,N_6027);
nand U6212 (N_6212,N_6141,N_6182);
or U6213 (N_6213,N_6019,N_6118);
or U6214 (N_6214,N_6033,N_6093);
xor U6215 (N_6215,N_6167,N_6142);
and U6216 (N_6216,N_6015,N_6148);
or U6217 (N_6217,N_6077,N_6078);
or U6218 (N_6218,N_6028,N_6038);
nor U6219 (N_6219,N_6039,N_6161);
nand U6220 (N_6220,N_6174,N_6002);
or U6221 (N_6221,N_6081,N_6140);
xnor U6222 (N_6222,N_6022,N_6136);
xor U6223 (N_6223,N_6099,N_6199);
nand U6224 (N_6224,N_6073,N_6040);
nand U6225 (N_6225,N_6029,N_6131);
xnor U6226 (N_6226,N_6170,N_6079);
xor U6227 (N_6227,N_6057,N_6066);
nor U6228 (N_6228,N_6153,N_6169);
xor U6229 (N_6229,N_6159,N_6069);
nor U6230 (N_6230,N_6089,N_6092);
xnor U6231 (N_6231,N_6171,N_6107);
nand U6232 (N_6232,N_6063,N_6135);
and U6233 (N_6233,N_6080,N_6185);
nand U6234 (N_6234,N_6082,N_6195);
or U6235 (N_6235,N_6156,N_6095);
xor U6236 (N_6236,N_6058,N_6133);
nor U6237 (N_6237,N_6055,N_6129);
xor U6238 (N_6238,N_6197,N_6074);
nor U6239 (N_6239,N_6101,N_6184);
nand U6240 (N_6240,N_6173,N_6031);
xor U6241 (N_6241,N_6044,N_6163);
or U6242 (N_6242,N_6168,N_6162);
or U6243 (N_6243,N_6021,N_6100);
nand U6244 (N_6244,N_6037,N_6030);
nor U6245 (N_6245,N_6186,N_6084);
xnor U6246 (N_6246,N_6102,N_6166);
nand U6247 (N_6247,N_6032,N_6117);
and U6248 (N_6248,N_6149,N_6194);
nand U6249 (N_6249,N_6013,N_6006);
or U6250 (N_6250,N_6043,N_6172);
nand U6251 (N_6251,N_6164,N_6126);
or U6252 (N_6252,N_6108,N_6076);
and U6253 (N_6253,N_6110,N_6008);
xnor U6254 (N_6254,N_6051,N_6054);
xor U6255 (N_6255,N_6094,N_6062);
and U6256 (N_6256,N_6127,N_6111);
nor U6257 (N_6257,N_6049,N_6130);
and U6258 (N_6258,N_6070,N_6120);
and U6259 (N_6259,N_6085,N_6024);
and U6260 (N_6260,N_6088,N_6020);
nor U6261 (N_6261,N_6138,N_6083);
or U6262 (N_6262,N_6113,N_6096);
or U6263 (N_6263,N_6177,N_6145);
and U6264 (N_6264,N_6045,N_6183);
and U6265 (N_6265,N_6137,N_6067);
xnor U6266 (N_6266,N_6114,N_6011);
nand U6267 (N_6267,N_6181,N_6165);
nor U6268 (N_6268,N_6155,N_6046);
and U6269 (N_6269,N_6123,N_6018);
nand U6270 (N_6270,N_6176,N_6041);
xor U6271 (N_6271,N_6036,N_6086);
nor U6272 (N_6272,N_6026,N_6158);
nand U6273 (N_6273,N_6034,N_6003);
or U6274 (N_6274,N_6035,N_6134);
or U6275 (N_6275,N_6042,N_6189);
and U6276 (N_6276,N_6056,N_6109);
nand U6277 (N_6277,N_6115,N_6059);
or U6278 (N_6278,N_6071,N_6188);
nand U6279 (N_6279,N_6146,N_6119);
xor U6280 (N_6280,N_6023,N_6143);
xnor U6281 (N_6281,N_6001,N_6178);
xor U6282 (N_6282,N_6154,N_6004);
nand U6283 (N_6283,N_6060,N_6125);
nor U6284 (N_6284,N_6064,N_6112);
and U6285 (N_6285,N_6106,N_6075);
and U6286 (N_6286,N_6105,N_6050);
or U6287 (N_6287,N_6007,N_6005);
xnor U6288 (N_6288,N_6012,N_6091);
xnor U6289 (N_6289,N_6152,N_6151);
xor U6290 (N_6290,N_6191,N_6010);
and U6291 (N_6291,N_6160,N_6053);
nor U6292 (N_6292,N_6116,N_6150);
and U6293 (N_6293,N_6128,N_6097);
nor U6294 (N_6294,N_6196,N_6072);
and U6295 (N_6295,N_6187,N_6193);
and U6296 (N_6296,N_6122,N_6180);
or U6297 (N_6297,N_6175,N_6068);
nand U6298 (N_6298,N_6098,N_6192);
or U6299 (N_6299,N_6179,N_6048);
or U6300 (N_6300,N_6143,N_6080);
xnor U6301 (N_6301,N_6131,N_6167);
xor U6302 (N_6302,N_6119,N_6192);
xnor U6303 (N_6303,N_6027,N_6091);
nand U6304 (N_6304,N_6077,N_6065);
and U6305 (N_6305,N_6031,N_6129);
nor U6306 (N_6306,N_6098,N_6158);
nor U6307 (N_6307,N_6042,N_6094);
or U6308 (N_6308,N_6000,N_6043);
or U6309 (N_6309,N_6025,N_6198);
xnor U6310 (N_6310,N_6147,N_6096);
or U6311 (N_6311,N_6052,N_6140);
nor U6312 (N_6312,N_6119,N_6090);
nand U6313 (N_6313,N_6195,N_6104);
nand U6314 (N_6314,N_6064,N_6110);
nor U6315 (N_6315,N_6197,N_6162);
nor U6316 (N_6316,N_6124,N_6185);
nand U6317 (N_6317,N_6183,N_6072);
nor U6318 (N_6318,N_6177,N_6076);
or U6319 (N_6319,N_6007,N_6107);
and U6320 (N_6320,N_6142,N_6112);
or U6321 (N_6321,N_6158,N_6017);
and U6322 (N_6322,N_6152,N_6002);
xor U6323 (N_6323,N_6066,N_6139);
and U6324 (N_6324,N_6154,N_6121);
nand U6325 (N_6325,N_6129,N_6112);
or U6326 (N_6326,N_6005,N_6151);
nor U6327 (N_6327,N_6076,N_6007);
xor U6328 (N_6328,N_6148,N_6132);
nor U6329 (N_6329,N_6093,N_6095);
or U6330 (N_6330,N_6017,N_6002);
nor U6331 (N_6331,N_6049,N_6070);
and U6332 (N_6332,N_6182,N_6113);
or U6333 (N_6333,N_6166,N_6144);
nor U6334 (N_6334,N_6035,N_6010);
or U6335 (N_6335,N_6105,N_6154);
nor U6336 (N_6336,N_6047,N_6035);
nand U6337 (N_6337,N_6058,N_6028);
or U6338 (N_6338,N_6130,N_6032);
or U6339 (N_6339,N_6084,N_6089);
or U6340 (N_6340,N_6099,N_6113);
and U6341 (N_6341,N_6044,N_6067);
xor U6342 (N_6342,N_6138,N_6086);
nor U6343 (N_6343,N_6167,N_6174);
nand U6344 (N_6344,N_6096,N_6135);
nand U6345 (N_6345,N_6146,N_6124);
xnor U6346 (N_6346,N_6061,N_6177);
xnor U6347 (N_6347,N_6098,N_6109);
xnor U6348 (N_6348,N_6133,N_6156);
or U6349 (N_6349,N_6194,N_6036);
xor U6350 (N_6350,N_6170,N_6194);
nand U6351 (N_6351,N_6041,N_6066);
nand U6352 (N_6352,N_6192,N_6139);
or U6353 (N_6353,N_6197,N_6180);
xor U6354 (N_6354,N_6148,N_6040);
nand U6355 (N_6355,N_6043,N_6008);
nor U6356 (N_6356,N_6083,N_6124);
xnor U6357 (N_6357,N_6137,N_6132);
xnor U6358 (N_6358,N_6163,N_6004);
xnor U6359 (N_6359,N_6115,N_6019);
or U6360 (N_6360,N_6105,N_6010);
nand U6361 (N_6361,N_6149,N_6119);
nand U6362 (N_6362,N_6129,N_6068);
xnor U6363 (N_6363,N_6079,N_6187);
and U6364 (N_6364,N_6121,N_6169);
nand U6365 (N_6365,N_6104,N_6126);
xor U6366 (N_6366,N_6082,N_6058);
and U6367 (N_6367,N_6148,N_6192);
and U6368 (N_6368,N_6153,N_6151);
nor U6369 (N_6369,N_6196,N_6173);
nor U6370 (N_6370,N_6071,N_6179);
nor U6371 (N_6371,N_6199,N_6165);
xnor U6372 (N_6372,N_6158,N_6137);
xor U6373 (N_6373,N_6166,N_6002);
xor U6374 (N_6374,N_6154,N_6065);
and U6375 (N_6375,N_6117,N_6042);
xnor U6376 (N_6376,N_6037,N_6044);
and U6377 (N_6377,N_6099,N_6186);
nor U6378 (N_6378,N_6067,N_6128);
nand U6379 (N_6379,N_6127,N_6178);
xor U6380 (N_6380,N_6085,N_6165);
and U6381 (N_6381,N_6167,N_6026);
nand U6382 (N_6382,N_6156,N_6045);
nor U6383 (N_6383,N_6031,N_6113);
or U6384 (N_6384,N_6125,N_6038);
nand U6385 (N_6385,N_6014,N_6169);
and U6386 (N_6386,N_6152,N_6091);
nand U6387 (N_6387,N_6045,N_6186);
or U6388 (N_6388,N_6134,N_6069);
or U6389 (N_6389,N_6024,N_6018);
nor U6390 (N_6390,N_6029,N_6096);
or U6391 (N_6391,N_6064,N_6024);
nor U6392 (N_6392,N_6039,N_6114);
nor U6393 (N_6393,N_6026,N_6148);
nand U6394 (N_6394,N_6020,N_6173);
nor U6395 (N_6395,N_6051,N_6018);
xor U6396 (N_6396,N_6057,N_6067);
nand U6397 (N_6397,N_6026,N_6129);
or U6398 (N_6398,N_6015,N_6075);
and U6399 (N_6399,N_6015,N_6092);
nand U6400 (N_6400,N_6389,N_6388);
nor U6401 (N_6401,N_6225,N_6373);
and U6402 (N_6402,N_6312,N_6292);
nand U6403 (N_6403,N_6380,N_6239);
and U6404 (N_6404,N_6356,N_6332);
nand U6405 (N_6405,N_6208,N_6290);
nand U6406 (N_6406,N_6237,N_6258);
nand U6407 (N_6407,N_6355,N_6251);
and U6408 (N_6408,N_6393,N_6291);
nor U6409 (N_6409,N_6215,N_6320);
nand U6410 (N_6410,N_6204,N_6232);
nand U6411 (N_6411,N_6354,N_6299);
and U6412 (N_6412,N_6288,N_6358);
nor U6413 (N_6413,N_6305,N_6347);
and U6414 (N_6414,N_6316,N_6360);
or U6415 (N_6415,N_6362,N_6370);
xor U6416 (N_6416,N_6308,N_6313);
nor U6417 (N_6417,N_6272,N_6333);
or U6418 (N_6418,N_6218,N_6234);
nor U6419 (N_6419,N_6350,N_6298);
and U6420 (N_6420,N_6341,N_6260);
nand U6421 (N_6421,N_6229,N_6274);
nand U6422 (N_6422,N_6357,N_6361);
xor U6423 (N_6423,N_6322,N_6226);
or U6424 (N_6424,N_6331,N_6275);
nor U6425 (N_6425,N_6295,N_6217);
nand U6426 (N_6426,N_6265,N_6256);
nand U6427 (N_6427,N_6236,N_6387);
nor U6428 (N_6428,N_6335,N_6321);
xnor U6429 (N_6429,N_6203,N_6318);
xnor U6430 (N_6430,N_6398,N_6276);
nand U6431 (N_6431,N_6392,N_6264);
xor U6432 (N_6432,N_6268,N_6329);
xor U6433 (N_6433,N_6270,N_6222);
nand U6434 (N_6434,N_6255,N_6266);
or U6435 (N_6435,N_6301,N_6365);
nor U6436 (N_6436,N_6330,N_6382);
and U6437 (N_6437,N_6383,N_6348);
nor U6438 (N_6438,N_6212,N_6249);
nand U6439 (N_6439,N_6248,N_6206);
nor U6440 (N_6440,N_6394,N_6257);
xnor U6441 (N_6441,N_6364,N_6377);
xor U6442 (N_6442,N_6381,N_6340);
and U6443 (N_6443,N_6384,N_6244);
and U6444 (N_6444,N_6343,N_6303);
or U6445 (N_6445,N_6349,N_6317);
xnor U6446 (N_6446,N_6363,N_6399);
or U6447 (N_6447,N_6294,N_6259);
nand U6448 (N_6448,N_6241,N_6211);
or U6449 (N_6449,N_6284,N_6385);
nor U6450 (N_6450,N_6325,N_6280);
nand U6451 (N_6451,N_6337,N_6221);
or U6452 (N_6452,N_6334,N_6353);
or U6453 (N_6453,N_6202,N_6395);
and U6454 (N_6454,N_6319,N_6216);
nand U6455 (N_6455,N_6231,N_6367);
nand U6456 (N_6456,N_6324,N_6397);
nand U6457 (N_6457,N_6338,N_6224);
nand U6458 (N_6458,N_6315,N_6201);
xor U6459 (N_6459,N_6366,N_6287);
nand U6460 (N_6460,N_6371,N_6228);
nand U6461 (N_6461,N_6327,N_6261);
nand U6462 (N_6462,N_6219,N_6336);
nor U6463 (N_6463,N_6283,N_6304);
nand U6464 (N_6464,N_6247,N_6390);
nand U6465 (N_6465,N_6378,N_6375);
and U6466 (N_6466,N_6372,N_6230);
and U6467 (N_6467,N_6220,N_6253);
nor U6468 (N_6468,N_6296,N_6242);
nor U6469 (N_6469,N_6200,N_6233);
xor U6470 (N_6470,N_6302,N_6345);
xnor U6471 (N_6471,N_6289,N_6271);
or U6472 (N_6472,N_6269,N_6267);
xnor U6473 (N_6473,N_6376,N_6246);
and U6474 (N_6474,N_6245,N_6278);
xor U6475 (N_6475,N_6374,N_6310);
nor U6476 (N_6476,N_6368,N_6396);
nor U6477 (N_6477,N_6352,N_6293);
nor U6478 (N_6478,N_6207,N_6300);
and U6479 (N_6479,N_6227,N_6277);
nand U6480 (N_6480,N_6344,N_6235);
or U6481 (N_6481,N_6223,N_6307);
nand U6482 (N_6482,N_6213,N_6282);
xnor U6483 (N_6483,N_6311,N_6309);
or U6484 (N_6484,N_6243,N_6286);
and U6485 (N_6485,N_6339,N_6369);
and U6486 (N_6486,N_6214,N_6250);
and U6487 (N_6487,N_6205,N_6254);
or U6488 (N_6488,N_6351,N_6314);
nand U6489 (N_6489,N_6263,N_6306);
xnor U6490 (N_6490,N_6346,N_6359);
nor U6491 (N_6491,N_6279,N_6297);
nor U6492 (N_6492,N_6238,N_6285);
xor U6493 (N_6493,N_6391,N_6240);
xor U6494 (N_6494,N_6326,N_6342);
and U6495 (N_6495,N_6328,N_6209);
nand U6496 (N_6496,N_6386,N_6252);
xor U6497 (N_6497,N_6262,N_6210);
nor U6498 (N_6498,N_6379,N_6273);
nor U6499 (N_6499,N_6281,N_6323);
or U6500 (N_6500,N_6298,N_6335);
and U6501 (N_6501,N_6343,N_6363);
and U6502 (N_6502,N_6294,N_6284);
or U6503 (N_6503,N_6299,N_6393);
or U6504 (N_6504,N_6246,N_6235);
nor U6505 (N_6505,N_6359,N_6363);
or U6506 (N_6506,N_6223,N_6277);
nand U6507 (N_6507,N_6373,N_6343);
xnor U6508 (N_6508,N_6271,N_6346);
nor U6509 (N_6509,N_6261,N_6227);
nand U6510 (N_6510,N_6230,N_6262);
xnor U6511 (N_6511,N_6365,N_6387);
nor U6512 (N_6512,N_6303,N_6250);
nand U6513 (N_6513,N_6203,N_6353);
xnor U6514 (N_6514,N_6211,N_6336);
and U6515 (N_6515,N_6294,N_6361);
nor U6516 (N_6516,N_6284,N_6208);
and U6517 (N_6517,N_6273,N_6322);
and U6518 (N_6518,N_6208,N_6308);
xor U6519 (N_6519,N_6241,N_6270);
nand U6520 (N_6520,N_6342,N_6219);
nor U6521 (N_6521,N_6234,N_6382);
xor U6522 (N_6522,N_6280,N_6235);
xor U6523 (N_6523,N_6386,N_6328);
nand U6524 (N_6524,N_6313,N_6223);
and U6525 (N_6525,N_6317,N_6253);
and U6526 (N_6526,N_6205,N_6237);
nand U6527 (N_6527,N_6212,N_6229);
or U6528 (N_6528,N_6374,N_6370);
or U6529 (N_6529,N_6241,N_6264);
or U6530 (N_6530,N_6224,N_6252);
or U6531 (N_6531,N_6307,N_6321);
or U6532 (N_6532,N_6265,N_6372);
xor U6533 (N_6533,N_6360,N_6210);
and U6534 (N_6534,N_6268,N_6242);
and U6535 (N_6535,N_6348,N_6289);
and U6536 (N_6536,N_6324,N_6238);
and U6537 (N_6537,N_6234,N_6216);
and U6538 (N_6538,N_6239,N_6237);
nand U6539 (N_6539,N_6344,N_6328);
and U6540 (N_6540,N_6311,N_6373);
xnor U6541 (N_6541,N_6274,N_6321);
nand U6542 (N_6542,N_6389,N_6207);
and U6543 (N_6543,N_6285,N_6329);
and U6544 (N_6544,N_6280,N_6399);
and U6545 (N_6545,N_6355,N_6267);
or U6546 (N_6546,N_6327,N_6395);
nand U6547 (N_6547,N_6351,N_6306);
and U6548 (N_6548,N_6376,N_6252);
and U6549 (N_6549,N_6206,N_6371);
xnor U6550 (N_6550,N_6201,N_6204);
nand U6551 (N_6551,N_6247,N_6346);
or U6552 (N_6552,N_6379,N_6377);
and U6553 (N_6553,N_6234,N_6340);
nand U6554 (N_6554,N_6309,N_6344);
nor U6555 (N_6555,N_6203,N_6341);
nor U6556 (N_6556,N_6377,N_6358);
nor U6557 (N_6557,N_6296,N_6354);
or U6558 (N_6558,N_6209,N_6391);
and U6559 (N_6559,N_6346,N_6263);
nor U6560 (N_6560,N_6323,N_6290);
xor U6561 (N_6561,N_6325,N_6377);
and U6562 (N_6562,N_6349,N_6370);
or U6563 (N_6563,N_6227,N_6390);
nand U6564 (N_6564,N_6308,N_6300);
nand U6565 (N_6565,N_6362,N_6327);
or U6566 (N_6566,N_6227,N_6266);
and U6567 (N_6567,N_6218,N_6381);
or U6568 (N_6568,N_6397,N_6388);
nand U6569 (N_6569,N_6247,N_6282);
xnor U6570 (N_6570,N_6297,N_6344);
and U6571 (N_6571,N_6202,N_6287);
xnor U6572 (N_6572,N_6368,N_6394);
nor U6573 (N_6573,N_6231,N_6260);
and U6574 (N_6574,N_6379,N_6325);
xor U6575 (N_6575,N_6279,N_6350);
nor U6576 (N_6576,N_6379,N_6208);
or U6577 (N_6577,N_6238,N_6320);
nor U6578 (N_6578,N_6262,N_6357);
and U6579 (N_6579,N_6366,N_6258);
nand U6580 (N_6580,N_6308,N_6330);
nor U6581 (N_6581,N_6319,N_6298);
nand U6582 (N_6582,N_6397,N_6229);
or U6583 (N_6583,N_6219,N_6373);
or U6584 (N_6584,N_6393,N_6251);
and U6585 (N_6585,N_6316,N_6282);
xnor U6586 (N_6586,N_6314,N_6336);
nor U6587 (N_6587,N_6304,N_6294);
and U6588 (N_6588,N_6320,N_6280);
xnor U6589 (N_6589,N_6280,N_6343);
or U6590 (N_6590,N_6275,N_6278);
and U6591 (N_6591,N_6224,N_6298);
nor U6592 (N_6592,N_6228,N_6255);
nor U6593 (N_6593,N_6351,N_6260);
nand U6594 (N_6594,N_6231,N_6256);
or U6595 (N_6595,N_6292,N_6241);
nor U6596 (N_6596,N_6300,N_6225);
nor U6597 (N_6597,N_6209,N_6386);
nand U6598 (N_6598,N_6218,N_6216);
and U6599 (N_6599,N_6238,N_6365);
nor U6600 (N_6600,N_6464,N_6501);
nor U6601 (N_6601,N_6412,N_6436);
nor U6602 (N_6602,N_6551,N_6478);
nor U6603 (N_6603,N_6535,N_6404);
or U6604 (N_6604,N_6511,N_6423);
nor U6605 (N_6605,N_6562,N_6589);
xor U6606 (N_6606,N_6523,N_6492);
xnor U6607 (N_6607,N_6487,N_6587);
and U6608 (N_6608,N_6543,N_6597);
nand U6609 (N_6609,N_6515,N_6495);
nor U6610 (N_6610,N_6552,N_6559);
and U6611 (N_6611,N_6558,N_6516);
nor U6612 (N_6612,N_6406,N_6434);
nor U6613 (N_6613,N_6514,N_6496);
or U6614 (N_6614,N_6534,N_6456);
nand U6615 (N_6615,N_6498,N_6599);
or U6616 (N_6616,N_6556,N_6424);
or U6617 (N_6617,N_6444,N_6462);
nor U6618 (N_6618,N_6421,N_6526);
nor U6619 (N_6619,N_6438,N_6585);
nand U6620 (N_6620,N_6544,N_6477);
and U6621 (N_6621,N_6512,N_6454);
nor U6622 (N_6622,N_6417,N_6595);
and U6623 (N_6623,N_6431,N_6486);
xor U6624 (N_6624,N_6504,N_6485);
or U6625 (N_6625,N_6531,N_6400);
and U6626 (N_6626,N_6576,N_6508);
and U6627 (N_6627,N_6510,N_6458);
xor U6628 (N_6628,N_6560,N_6468);
nor U6629 (N_6629,N_6432,N_6461);
or U6630 (N_6630,N_6455,N_6569);
xnor U6631 (N_6631,N_6577,N_6440);
and U6632 (N_6632,N_6573,N_6443);
or U6633 (N_6633,N_6401,N_6415);
xor U6634 (N_6634,N_6584,N_6507);
nand U6635 (N_6635,N_6442,N_6546);
or U6636 (N_6636,N_6448,N_6525);
xnor U6637 (N_6637,N_6418,N_6593);
xnor U6638 (N_6638,N_6467,N_6583);
and U6639 (N_6639,N_6446,N_6567);
nor U6640 (N_6640,N_6413,N_6465);
and U6641 (N_6641,N_6565,N_6489);
nand U6642 (N_6642,N_6453,N_6591);
xnor U6643 (N_6643,N_6503,N_6528);
nor U6644 (N_6644,N_6532,N_6491);
or U6645 (N_6645,N_6469,N_6476);
nor U6646 (N_6646,N_6439,N_6422);
xor U6647 (N_6647,N_6407,N_6445);
and U6648 (N_6648,N_6426,N_6568);
nor U6649 (N_6649,N_6564,N_6509);
nand U6650 (N_6650,N_6410,N_6566);
and U6651 (N_6651,N_6493,N_6527);
nand U6652 (N_6652,N_6450,N_6409);
or U6653 (N_6653,N_6484,N_6538);
nand U6654 (N_6654,N_6460,N_6433);
xnor U6655 (N_6655,N_6557,N_6449);
or U6656 (N_6656,N_6517,N_6437);
and U6657 (N_6657,N_6466,N_6518);
xor U6658 (N_6658,N_6579,N_6554);
nor U6659 (N_6659,N_6561,N_6420);
and U6660 (N_6660,N_6419,N_6494);
nor U6661 (N_6661,N_6403,N_6540);
and U6662 (N_6662,N_6483,N_6529);
nand U6663 (N_6663,N_6451,N_6513);
nand U6664 (N_6664,N_6479,N_6574);
nand U6665 (N_6665,N_6429,N_6598);
nand U6666 (N_6666,N_6572,N_6482);
and U6667 (N_6667,N_6472,N_6530);
and U6668 (N_6668,N_6555,N_6505);
nor U6669 (N_6669,N_6571,N_6553);
nor U6670 (N_6670,N_6549,N_6402);
nor U6671 (N_6671,N_6473,N_6457);
nand U6672 (N_6672,N_6547,N_6480);
or U6673 (N_6673,N_6506,N_6519);
xor U6674 (N_6674,N_6490,N_6575);
nor U6675 (N_6675,N_6435,N_6548);
or U6676 (N_6676,N_6563,N_6416);
and U6677 (N_6677,N_6475,N_6578);
xor U6678 (N_6678,N_6545,N_6592);
xnor U6679 (N_6679,N_6536,N_6539);
nor U6680 (N_6680,N_6537,N_6428);
xnor U6681 (N_6681,N_6550,N_6580);
or U6682 (N_6682,N_6541,N_6414);
or U6683 (N_6683,N_6521,N_6471);
nor U6684 (N_6684,N_6542,N_6499);
and U6685 (N_6685,N_6586,N_6441);
or U6686 (N_6686,N_6520,N_6596);
xor U6687 (N_6687,N_6463,N_6427);
xnor U6688 (N_6688,N_6405,N_6590);
and U6689 (N_6689,N_6459,N_6581);
xnor U6690 (N_6690,N_6481,N_6588);
nor U6691 (N_6691,N_6408,N_6470);
or U6692 (N_6692,N_6430,N_6452);
nand U6693 (N_6693,N_6488,N_6522);
nand U6694 (N_6694,N_6447,N_6502);
nand U6695 (N_6695,N_6524,N_6570);
and U6696 (N_6696,N_6533,N_6497);
nand U6697 (N_6697,N_6500,N_6425);
and U6698 (N_6698,N_6474,N_6594);
or U6699 (N_6699,N_6411,N_6582);
or U6700 (N_6700,N_6459,N_6572);
nor U6701 (N_6701,N_6430,N_6567);
xnor U6702 (N_6702,N_6457,N_6529);
nand U6703 (N_6703,N_6534,N_6402);
nand U6704 (N_6704,N_6511,N_6591);
nor U6705 (N_6705,N_6420,N_6584);
nor U6706 (N_6706,N_6455,N_6491);
nand U6707 (N_6707,N_6519,N_6408);
xnor U6708 (N_6708,N_6560,N_6403);
nor U6709 (N_6709,N_6430,N_6411);
xor U6710 (N_6710,N_6538,N_6483);
and U6711 (N_6711,N_6565,N_6445);
and U6712 (N_6712,N_6577,N_6597);
and U6713 (N_6713,N_6494,N_6483);
and U6714 (N_6714,N_6596,N_6466);
and U6715 (N_6715,N_6556,N_6420);
or U6716 (N_6716,N_6583,N_6569);
xor U6717 (N_6717,N_6417,N_6533);
or U6718 (N_6718,N_6583,N_6494);
and U6719 (N_6719,N_6544,N_6453);
nand U6720 (N_6720,N_6523,N_6585);
or U6721 (N_6721,N_6432,N_6597);
xor U6722 (N_6722,N_6511,N_6556);
nor U6723 (N_6723,N_6591,N_6596);
xor U6724 (N_6724,N_6401,N_6443);
nand U6725 (N_6725,N_6440,N_6456);
nand U6726 (N_6726,N_6461,N_6463);
and U6727 (N_6727,N_6599,N_6580);
xor U6728 (N_6728,N_6451,N_6455);
nor U6729 (N_6729,N_6427,N_6445);
or U6730 (N_6730,N_6431,N_6497);
or U6731 (N_6731,N_6553,N_6461);
and U6732 (N_6732,N_6436,N_6469);
xnor U6733 (N_6733,N_6526,N_6403);
and U6734 (N_6734,N_6405,N_6507);
nor U6735 (N_6735,N_6448,N_6580);
nand U6736 (N_6736,N_6558,N_6443);
and U6737 (N_6737,N_6449,N_6565);
or U6738 (N_6738,N_6527,N_6465);
or U6739 (N_6739,N_6588,N_6448);
nand U6740 (N_6740,N_6523,N_6453);
or U6741 (N_6741,N_6527,N_6473);
nand U6742 (N_6742,N_6530,N_6521);
and U6743 (N_6743,N_6410,N_6533);
nand U6744 (N_6744,N_6433,N_6599);
and U6745 (N_6745,N_6403,N_6467);
nand U6746 (N_6746,N_6535,N_6537);
and U6747 (N_6747,N_6539,N_6579);
nor U6748 (N_6748,N_6418,N_6458);
and U6749 (N_6749,N_6556,N_6546);
nand U6750 (N_6750,N_6436,N_6431);
nor U6751 (N_6751,N_6550,N_6436);
nand U6752 (N_6752,N_6499,N_6462);
or U6753 (N_6753,N_6508,N_6548);
nand U6754 (N_6754,N_6551,N_6555);
nand U6755 (N_6755,N_6448,N_6592);
xnor U6756 (N_6756,N_6538,N_6424);
or U6757 (N_6757,N_6579,N_6446);
and U6758 (N_6758,N_6512,N_6532);
and U6759 (N_6759,N_6587,N_6411);
nand U6760 (N_6760,N_6587,N_6524);
or U6761 (N_6761,N_6488,N_6425);
or U6762 (N_6762,N_6424,N_6471);
nor U6763 (N_6763,N_6425,N_6411);
nand U6764 (N_6764,N_6514,N_6465);
xnor U6765 (N_6765,N_6570,N_6460);
nand U6766 (N_6766,N_6548,N_6443);
and U6767 (N_6767,N_6452,N_6584);
or U6768 (N_6768,N_6450,N_6452);
or U6769 (N_6769,N_6597,N_6406);
and U6770 (N_6770,N_6471,N_6564);
nand U6771 (N_6771,N_6504,N_6524);
or U6772 (N_6772,N_6440,N_6410);
xnor U6773 (N_6773,N_6555,N_6520);
xor U6774 (N_6774,N_6550,N_6413);
and U6775 (N_6775,N_6465,N_6576);
nor U6776 (N_6776,N_6467,N_6590);
xnor U6777 (N_6777,N_6492,N_6566);
nand U6778 (N_6778,N_6577,N_6403);
or U6779 (N_6779,N_6450,N_6469);
and U6780 (N_6780,N_6586,N_6426);
nor U6781 (N_6781,N_6531,N_6494);
xnor U6782 (N_6782,N_6526,N_6558);
or U6783 (N_6783,N_6427,N_6536);
or U6784 (N_6784,N_6422,N_6539);
and U6785 (N_6785,N_6405,N_6521);
and U6786 (N_6786,N_6471,N_6419);
nor U6787 (N_6787,N_6588,N_6573);
nor U6788 (N_6788,N_6553,N_6556);
and U6789 (N_6789,N_6570,N_6428);
nand U6790 (N_6790,N_6469,N_6553);
or U6791 (N_6791,N_6420,N_6582);
nand U6792 (N_6792,N_6598,N_6545);
xnor U6793 (N_6793,N_6434,N_6595);
nor U6794 (N_6794,N_6480,N_6594);
and U6795 (N_6795,N_6514,N_6540);
xnor U6796 (N_6796,N_6403,N_6525);
xnor U6797 (N_6797,N_6429,N_6525);
or U6798 (N_6798,N_6559,N_6445);
xor U6799 (N_6799,N_6559,N_6495);
nor U6800 (N_6800,N_6710,N_6748);
xor U6801 (N_6801,N_6696,N_6611);
xnor U6802 (N_6802,N_6691,N_6772);
and U6803 (N_6803,N_6700,N_6787);
and U6804 (N_6804,N_6750,N_6646);
nand U6805 (N_6805,N_6686,N_6753);
nand U6806 (N_6806,N_6645,N_6720);
and U6807 (N_6807,N_6746,N_6707);
nor U6808 (N_6808,N_6791,N_6647);
or U6809 (N_6809,N_6784,N_6719);
nand U6810 (N_6810,N_6766,N_6642);
xor U6811 (N_6811,N_6758,N_6716);
xor U6812 (N_6812,N_6644,N_6683);
nand U6813 (N_6813,N_6681,N_6737);
or U6814 (N_6814,N_6775,N_6661);
or U6815 (N_6815,N_6634,N_6636);
nor U6816 (N_6816,N_6643,N_6672);
nor U6817 (N_6817,N_6630,N_6654);
nand U6818 (N_6818,N_6713,N_6679);
and U6819 (N_6819,N_6781,N_6722);
nand U6820 (N_6820,N_6721,N_6633);
nor U6821 (N_6821,N_6733,N_6675);
xnor U6822 (N_6822,N_6715,N_6616);
nor U6823 (N_6823,N_6635,N_6751);
and U6824 (N_6824,N_6756,N_6745);
or U6825 (N_6825,N_6712,N_6651);
and U6826 (N_6826,N_6671,N_6740);
nand U6827 (N_6827,N_6778,N_6797);
nor U6828 (N_6828,N_6793,N_6706);
xor U6829 (N_6829,N_6732,N_6620);
nor U6830 (N_6830,N_6762,N_6780);
or U6831 (N_6831,N_6689,N_6729);
xnor U6832 (N_6832,N_6697,N_6698);
or U6833 (N_6833,N_6747,N_6627);
nor U6834 (N_6834,N_6763,N_6769);
nor U6835 (N_6835,N_6779,N_6743);
xnor U6836 (N_6836,N_6760,N_6704);
or U6837 (N_6837,N_6711,N_6687);
nand U6838 (N_6838,N_6602,N_6776);
or U6839 (N_6839,N_6640,N_6610);
and U6840 (N_6840,N_6741,N_6673);
and U6841 (N_6841,N_6629,N_6755);
nor U6842 (N_6842,N_6724,N_6608);
nor U6843 (N_6843,N_6718,N_6670);
and U6844 (N_6844,N_6663,N_6702);
xor U6845 (N_6845,N_6777,N_6761);
nor U6846 (N_6846,N_6767,N_6768);
and U6847 (N_6847,N_6674,N_6714);
xnor U6848 (N_6848,N_6625,N_6662);
xor U6849 (N_6849,N_6790,N_6771);
xnor U6850 (N_6850,N_6744,N_6639);
and U6851 (N_6851,N_6600,N_6786);
and U6852 (N_6852,N_6624,N_6655);
nand U6853 (N_6853,N_6676,N_6641);
xor U6854 (N_6854,N_6736,N_6626);
nand U6855 (N_6855,N_6660,N_6703);
nor U6856 (N_6856,N_6694,N_6795);
and U6857 (N_6857,N_6618,N_6613);
nor U6858 (N_6858,N_6604,N_6677);
and U6859 (N_6859,N_6765,N_6690);
or U6860 (N_6860,N_6658,N_6606);
nor U6861 (N_6861,N_6603,N_6725);
and U6862 (N_6862,N_6742,N_6664);
or U6863 (N_6863,N_6609,N_6623);
nor U6864 (N_6864,N_6785,N_6705);
nand U6865 (N_6865,N_6678,N_6657);
and U6866 (N_6866,N_6788,N_6631);
xnor U6867 (N_6867,N_6666,N_6726);
nor U6868 (N_6868,N_6653,N_6773);
and U6869 (N_6869,N_6628,N_6692);
nor U6870 (N_6870,N_6728,N_6648);
nand U6871 (N_6871,N_6649,N_6796);
or U6872 (N_6872,N_6738,N_6799);
or U6873 (N_6873,N_6665,N_6637);
or U6874 (N_6874,N_6684,N_6759);
or U6875 (N_6875,N_6727,N_6695);
xor U6876 (N_6876,N_6764,N_6617);
nand U6877 (N_6877,N_6717,N_6621);
and U6878 (N_6878,N_6622,N_6693);
and U6879 (N_6879,N_6783,N_6730);
or U6880 (N_6880,N_6774,N_6770);
xnor U6881 (N_6881,N_6656,N_6699);
xor U6882 (N_6882,N_6638,N_6659);
nand U6883 (N_6883,N_6735,N_6792);
and U6884 (N_6884,N_6731,N_6601);
nand U6885 (N_6885,N_6685,N_6734);
xnor U6886 (N_6886,N_6723,N_6632);
nor U6887 (N_6887,N_6754,N_6612);
nor U6888 (N_6888,N_6619,N_6798);
xnor U6889 (N_6889,N_6668,N_6667);
and U6890 (N_6890,N_6709,N_6701);
nor U6891 (N_6891,N_6749,N_6688);
nand U6892 (N_6892,N_6669,N_6682);
nor U6893 (N_6893,N_6652,N_6794);
nor U6894 (N_6894,N_6615,N_6650);
and U6895 (N_6895,N_6752,N_6680);
and U6896 (N_6896,N_6789,N_6607);
xor U6897 (N_6897,N_6757,N_6605);
or U6898 (N_6898,N_6782,N_6739);
or U6899 (N_6899,N_6614,N_6708);
and U6900 (N_6900,N_6763,N_6706);
nor U6901 (N_6901,N_6754,N_6601);
and U6902 (N_6902,N_6757,N_6744);
and U6903 (N_6903,N_6715,N_6719);
or U6904 (N_6904,N_6799,N_6630);
xnor U6905 (N_6905,N_6669,N_6695);
nor U6906 (N_6906,N_6743,N_6775);
or U6907 (N_6907,N_6689,N_6786);
and U6908 (N_6908,N_6621,N_6688);
or U6909 (N_6909,N_6748,N_6767);
nand U6910 (N_6910,N_6638,N_6642);
or U6911 (N_6911,N_6760,N_6699);
and U6912 (N_6912,N_6648,N_6783);
xnor U6913 (N_6913,N_6619,N_6749);
and U6914 (N_6914,N_6683,N_6676);
and U6915 (N_6915,N_6618,N_6714);
nor U6916 (N_6916,N_6645,N_6629);
xor U6917 (N_6917,N_6619,N_6724);
or U6918 (N_6918,N_6625,N_6704);
nand U6919 (N_6919,N_6604,N_6706);
xor U6920 (N_6920,N_6661,N_6754);
nand U6921 (N_6921,N_6762,N_6638);
and U6922 (N_6922,N_6683,N_6744);
xnor U6923 (N_6923,N_6746,N_6789);
or U6924 (N_6924,N_6763,N_6602);
nor U6925 (N_6925,N_6618,N_6640);
nor U6926 (N_6926,N_6624,N_6653);
and U6927 (N_6927,N_6704,N_6749);
or U6928 (N_6928,N_6607,N_6627);
or U6929 (N_6929,N_6790,N_6772);
nor U6930 (N_6930,N_6637,N_6755);
nand U6931 (N_6931,N_6799,N_6790);
and U6932 (N_6932,N_6783,N_6670);
xnor U6933 (N_6933,N_6651,N_6689);
xor U6934 (N_6934,N_6778,N_6698);
nand U6935 (N_6935,N_6765,N_6749);
and U6936 (N_6936,N_6784,N_6707);
or U6937 (N_6937,N_6783,N_6656);
xor U6938 (N_6938,N_6631,N_6626);
or U6939 (N_6939,N_6764,N_6644);
nand U6940 (N_6940,N_6797,N_6623);
and U6941 (N_6941,N_6664,N_6685);
nand U6942 (N_6942,N_6705,N_6767);
and U6943 (N_6943,N_6658,N_6780);
and U6944 (N_6944,N_6763,N_6624);
nor U6945 (N_6945,N_6660,N_6748);
nand U6946 (N_6946,N_6755,N_6612);
and U6947 (N_6947,N_6615,N_6671);
xnor U6948 (N_6948,N_6778,N_6600);
nand U6949 (N_6949,N_6767,N_6636);
and U6950 (N_6950,N_6733,N_6775);
xor U6951 (N_6951,N_6731,N_6631);
nor U6952 (N_6952,N_6612,N_6609);
or U6953 (N_6953,N_6752,N_6663);
and U6954 (N_6954,N_6660,N_6704);
nand U6955 (N_6955,N_6743,N_6618);
and U6956 (N_6956,N_6723,N_6759);
or U6957 (N_6957,N_6651,N_6601);
xor U6958 (N_6958,N_6755,N_6618);
and U6959 (N_6959,N_6705,N_6656);
xnor U6960 (N_6960,N_6776,N_6629);
and U6961 (N_6961,N_6625,N_6766);
nor U6962 (N_6962,N_6797,N_6616);
and U6963 (N_6963,N_6721,N_6718);
nand U6964 (N_6964,N_6733,N_6638);
and U6965 (N_6965,N_6770,N_6700);
or U6966 (N_6966,N_6626,N_6606);
and U6967 (N_6967,N_6765,N_6670);
nor U6968 (N_6968,N_6745,N_6671);
nor U6969 (N_6969,N_6688,N_6760);
nor U6970 (N_6970,N_6780,N_6662);
nor U6971 (N_6971,N_6687,N_6766);
nor U6972 (N_6972,N_6662,N_6681);
or U6973 (N_6973,N_6635,N_6768);
or U6974 (N_6974,N_6737,N_6787);
and U6975 (N_6975,N_6764,N_6746);
nand U6976 (N_6976,N_6782,N_6722);
and U6977 (N_6977,N_6652,N_6731);
or U6978 (N_6978,N_6786,N_6697);
nand U6979 (N_6979,N_6756,N_6686);
nand U6980 (N_6980,N_6641,N_6730);
xor U6981 (N_6981,N_6791,N_6717);
nor U6982 (N_6982,N_6677,N_6790);
nor U6983 (N_6983,N_6695,N_6697);
xor U6984 (N_6984,N_6747,N_6703);
or U6985 (N_6985,N_6604,N_6703);
and U6986 (N_6986,N_6644,N_6786);
nor U6987 (N_6987,N_6639,N_6656);
and U6988 (N_6988,N_6652,N_6711);
nand U6989 (N_6989,N_6720,N_6774);
nand U6990 (N_6990,N_6722,N_6718);
nor U6991 (N_6991,N_6709,N_6781);
or U6992 (N_6992,N_6608,N_6726);
or U6993 (N_6993,N_6656,N_6671);
or U6994 (N_6994,N_6621,N_6648);
or U6995 (N_6995,N_6706,N_6665);
nand U6996 (N_6996,N_6670,N_6757);
nor U6997 (N_6997,N_6636,N_6712);
xor U6998 (N_6998,N_6644,N_6738);
or U6999 (N_6999,N_6757,N_6700);
nor U7000 (N_7000,N_6895,N_6859);
nor U7001 (N_7001,N_6872,N_6876);
and U7002 (N_7002,N_6953,N_6816);
or U7003 (N_7003,N_6873,N_6866);
nor U7004 (N_7004,N_6985,N_6824);
nor U7005 (N_7005,N_6913,N_6814);
nor U7006 (N_7006,N_6957,N_6904);
nand U7007 (N_7007,N_6834,N_6871);
nand U7008 (N_7008,N_6813,N_6833);
xor U7009 (N_7009,N_6979,N_6861);
or U7010 (N_7010,N_6903,N_6900);
and U7011 (N_7011,N_6839,N_6853);
and U7012 (N_7012,N_6973,N_6880);
and U7013 (N_7013,N_6998,N_6817);
xnor U7014 (N_7014,N_6920,N_6825);
nor U7015 (N_7015,N_6863,N_6815);
or U7016 (N_7016,N_6927,N_6980);
and U7017 (N_7017,N_6965,N_6902);
xor U7018 (N_7018,N_6964,N_6906);
nand U7019 (N_7019,N_6974,N_6832);
and U7020 (N_7020,N_6898,N_6990);
or U7021 (N_7021,N_6919,N_6981);
and U7022 (N_7022,N_6933,N_6955);
nand U7023 (N_7023,N_6970,N_6862);
xnor U7024 (N_7024,N_6810,N_6860);
xor U7025 (N_7025,N_6851,N_6910);
nor U7026 (N_7026,N_6847,N_6867);
nand U7027 (N_7027,N_6891,N_6864);
and U7028 (N_7028,N_6940,N_6812);
nand U7029 (N_7029,N_6943,N_6885);
nor U7030 (N_7030,N_6941,N_6952);
xor U7031 (N_7031,N_6987,N_6956);
or U7032 (N_7032,N_6869,N_6884);
and U7033 (N_7033,N_6944,N_6971);
or U7034 (N_7034,N_6950,N_6909);
xnor U7035 (N_7035,N_6858,N_6951);
nor U7036 (N_7036,N_6838,N_6837);
or U7037 (N_7037,N_6842,N_6830);
xnor U7038 (N_7038,N_6854,N_6845);
and U7039 (N_7039,N_6959,N_6829);
or U7040 (N_7040,N_6921,N_6881);
nor U7041 (N_7041,N_6984,N_6879);
xnor U7042 (N_7042,N_6882,N_6823);
xor U7043 (N_7043,N_6877,N_6992);
and U7044 (N_7044,N_6975,N_6938);
xnor U7045 (N_7045,N_6945,N_6937);
xnor U7046 (N_7046,N_6896,N_6994);
nand U7047 (N_7047,N_6855,N_6849);
and U7048 (N_7048,N_6907,N_6978);
or U7049 (N_7049,N_6991,N_6905);
xor U7050 (N_7050,N_6948,N_6843);
or U7051 (N_7051,N_6966,N_6846);
nand U7052 (N_7052,N_6878,N_6960);
and U7053 (N_7053,N_6865,N_6932);
and U7054 (N_7054,N_6894,N_6897);
nor U7055 (N_7055,N_6831,N_6806);
or U7056 (N_7056,N_6803,N_6982);
nor U7057 (N_7057,N_6805,N_6883);
and U7058 (N_7058,N_6874,N_6804);
and U7059 (N_7059,N_6848,N_6931);
xnor U7060 (N_7060,N_6901,N_6995);
nand U7061 (N_7061,N_6929,N_6809);
and U7062 (N_7062,N_6989,N_6999);
nand U7063 (N_7063,N_6870,N_6852);
nor U7064 (N_7064,N_6801,N_6886);
nor U7065 (N_7065,N_6868,N_6947);
nor U7066 (N_7066,N_6908,N_6841);
xnor U7067 (N_7067,N_6976,N_6887);
and U7068 (N_7068,N_6961,N_6915);
nor U7069 (N_7069,N_6856,N_6923);
and U7070 (N_7070,N_6818,N_6821);
nand U7071 (N_7071,N_6912,N_6958);
or U7072 (N_7072,N_6967,N_6917);
and U7073 (N_7073,N_6936,N_6836);
nand U7074 (N_7074,N_6934,N_6889);
nand U7075 (N_7075,N_6827,N_6914);
or U7076 (N_7076,N_6969,N_6993);
and U7077 (N_7077,N_6850,N_6963);
nand U7078 (N_7078,N_6949,N_6888);
nor U7079 (N_7079,N_6835,N_6997);
nor U7080 (N_7080,N_6922,N_6928);
or U7081 (N_7081,N_6946,N_6996);
xor U7082 (N_7082,N_6962,N_6802);
xor U7083 (N_7083,N_6939,N_6828);
nor U7084 (N_7084,N_6972,N_6800);
nand U7085 (N_7085,N_6935,N_6840);
and U7086 (N_7086,N_6924,N_6986);
nor U7087 (N_7087,N_6918,N_6988);
and U7088 (N_7088,N_6892,N_6930);
nor U7089 (N_7089,N_6890,N_6811);
nand U7090 (N_7090,N_6857,N_6820);
nand U7091 (N_7091,N_6911,N_6954);
and U7092 (N_7092,N_6844,N_6899);
xnor U7093 (N_7093,N_6968,N_6893);
nor U7094 (N_7094,N_6819,N_6926);
and U7095 (N_7095,N_6826,N_6808);
or U7096 (N_7096,N_6916,N_6822);
or U7097 (N_7097,N_6925,N_6807);
nor U7098 (N_7098,N_6875,N_6942);
xnor U7099 (N_7099,N_6983,N_6977);
nand U7100 (N_7100,N_6940,N_6891);
and U7101 (N_7101,N_6987,N_6995);
nand U7102 (N_7102,N_6863,N_6922);
nand U7103 (N_7103,N_6948,N_6842);
and U7104 (N_7104,N_6836,N_6904);
nor U7105 (N_7105,N_6902,N_6807);
nand U7106 (N_7106,N_6803,N_6845);
xor U7107 (N_7107,N_6841,N_6931);
and U7108 (N_7108,N_6845,N_6827);
xor U7109 (N_7109,N_6883,N_6809);
nand U7110 (N_7110,N_6996,N_6884);
xor U7111 (N_7111,N_6845,N_6921);
or U7112 (N_7112,N_6848,N_6985);
xnor U7113 (N_7113,N_6821,N_6917);
nand U7114 (N_7114,N_6856,N_6815);
or U7115 (N_7115,N_6930,N_6905);
nor U7116 (N_7116,N_6833,N_6950);
nor U7117 (N_7117,N_6859,N_6957);
xnor U7118 (N_7118,N_6867,N_6891);
nand U7119 (N_7119,N_6981,N_6992);
and U7120 (N_7120,N_6980,N_6928);
xnor U7121 (N_7121,N_6873,N_6967);
xor U7122 (N_7122,N_6982,N_6840);
xor U7123 (N_7123,N_6824,N_6980);
nor U7124 (N_7124,N_6849,N_6973);
xnor U7125 (N_7125,N_6882,N_6984);
or U7126 (N_7126,N_6972,N_6968);
nor U7127 (N_7127,N_6855,N_6898);
nor U7128 (N_7128,N_6853,N_6828);
nand U7129 (N_7129,N_6962,N_6985);
or U7130 (N_7130,N_6935,N_6942);
xor U7131 (N_7131,N_6901,N_6884);
nand U7132 (N_7132,N_6931,N_6866);
xnor U7133 (N_7133,N_6809,N_6977);
or U7134 (N_7134,N_6870,N_6807);
and U7135 (N_7135,N_6869,N_6881);
or U7136 (N_7136,N_6885,N_6912);
xor U7137 (N_7137,N_6947,N_6970);
xor U7138 (N_7138,N_6850,N_6830);
or U7139 (N_7139,N_6823,N_6858);
xnor U7140 (N_7140,N_6920,N_6865);
and U7141 (N_7141,N_6801,N_6969);
xnor U7142 (N_7142,N_6808,N_6985);
and U7143 (N_7143,N_6937,N_6925);
nand U7144 (N_7144,N_6961,N_6981);
nor U7145 (N_7145,N_6950,N_6938);
or U7146 (N_7146,N_6974,N_6929);
nand U7147 (N_7147,N_6832,N_6912);
nor U7148 (N_7148,N_6889,N_6829);
xnor U7149 (N_7149,N_6883,N_6974);
nor U7150 (N_7150,N_6882,N_6968);
nand U7151 (N_7151,N_6896,N_6856);
or U7152 (N_7152,N_6897,N_6921);
nand U7153 (N_7153,N_6920,N_6851);
and U7154 (N_7154,N_6876,N_6887);
nand U7155 (N_7155,N_6936,N_6875);
nor U7156 (N_7156,N_6981,N_6990);
nor U7157 (N_7157,N_6941,N_6876);
nand U7158 (N_7158,N_6894,N_6961);
xor U7159 (N_7159,N_6937,N_6889);
xnor U7160 (N_7160,N_6987,N_6817);
or U7161 (N_7161,N_6841,N_6998);
xor U7162 (N_7162,N_6998,N_6908);
and U7163 (N_7163,N_6992,N_6998);
nor U7164 (N_7164,N_6880,N_6836);
nor U7165 (N_7165,N_6838,N_6812);
and U7166 (N_7166,N_6869,N_6821);
and U7167 (N_7167,N_6850,N_6926);
nand U7168 (N_7168,N_6999,N_6869);
xnor U7169 (N_7169,N_6900,N_6833);
or U7170 (N_7170,N_6848,N_6849);
nand U7171 (N_7171,N_6974,N_6980);
nand U7172 (N_7172,N_6849,N_6865);
nand U7173 (N_7173,N_6836,N_6959);
or U7174 (N_7174,N_6813,N_6872);
or U7175 (N_7175,N_6824,N_6987);
nand U7176 (N_7176,N_6986,N_6845);
xnor U7177 (N_7177,N_6898,N_6860);
xnor U7178 (N_7178,N_6969,N_6831);
or U7179 (N_7179,N_6874,N_6948);
or U7180 (N_7180,N_6930,N_6870);
or U7181 (N_7181,N_6893,N_6911);
nand U7182 (N_7182,N_6828,N_6867);
xor U7183 (N_7183,N_6979,N_6838);
or U7184 (N_7184,N_6858,N_6845);
and U7185 (N_7185,N_6863,N_6800);
and U7186 (N_7186,N_6919,N_6947);
nand U7187 (N_7187,N_6924,N_6816);
and U7188 (N_7188,N_6904,N_6994);
xnor U7189 (N_7189,N_6855,N_6990);
nor U7190 (N_7190,N_6893,N_6903);
or U7191 (N_7191,N_6806,N_6913);
and U7192 (N_7192,N_6988,N_6872);
nor U7193 (N_7193,N_6916,N_6991);
nand U7194 (N_7194,N_6912,N_6948);
or U7195 (N_7195,N_6845,N_6897);
nand U7196 (N_7196,N_6919,N_6963);
nor U7197 (N_7197,N_6888,N_6962);
or U7198 (N_7198,N_6819,N_6994);
and U7199 (N_7199,N_6945,N_6821);
and U7200 (N_7200,N_7174,N_7103);
xnor U7201 (N_7201,N_7069,N_7167);
xor U7202 (N_7202,N_7175,N_7128);
or U7203 (N_7203,N_7044,N_7171);
or U7204 (N_7204,N_7155,N_7054);
xor U7205 (N_7205,N_7085,N_7192);
nor U7206 (N_7206,N_7023,N_7066);
nor U7207 (N_7207,N_7083,N_7132);
or U7208 (N_7208,N_7135,N_7159);
xnor U7209 (N_7209,N_7068,N_7150);
or U7210 (N_7210,N_7084,N_7047);
nor U7211 (N_7211,N_7163,N_7017);
nand U7212 (N_7212,N_7067,N_7111);
xnor U7213 (N_7213,N_7016,N_7166);
xnor U7214 (N_7214,N_7057,N_7036);
or U7215 (N_7215,N_7061,N_7152);
xor U7216 (N_7216,N_7194,N_7091);
xnor U7217 (N_7217,N_7088,N_7018);
and U7218 (N_7218,N_7006,N_7026);
xor U7219 (N_7219,N_7079,N_7186);
xor U7220 (N_7220,N_7092,N_7131);
and U7221 (N_7221,N_7191,N_7099);
and U7222 (N_7222,N_7060,N_7119);
or U7223 (N_7223,N_7185,N_7056);
nor U7224 (N_7224,N_7145,N_7179);
and U7225 (N_7225,N_7102,N_7130);
xor U7226 (N_7226,N_7143,N_7096);
and U7227 (N_7227,N_7183,N_7195);
nor U7228 (N_7228,N_7029,N_7072);
nand U7229 (N_7229,N_7107,N_7041);
or U7230 (N_7230,N_7073,N_7090);
and U7231 (N_7231,N_7037,N_7021);
xor U7232 (N_7232,N_7173,N_7100);
and U7233 (N_7233,N_7011,N_7022);
nand U7234 (N_7234,N_7063,N_7129);
nand U7235 (N_7235,N_7162,N_7013);
or U7236 (N_7236,N_7080,N_7115);
or U7237 (N_7237,N_7113,N_7187);
and U7238 (N_7238,N_7008,N_7127);
nand U7239 (N_7239,N_7114,N_7108);
nor U7240 (N_7240,N_7146,N_7116);
nand U7241 (N_7241,N_7025,N_7141);
and U7242 (N_7242,N_7045,N_7078);
nand U7243 (N_7243,N_7059,N_7032);
and U7244 (N_7244,N_7055,N_7065);
xor U7245 (N_7245,N_7147,N_7176);
nor U7246 (N_7246,N_7051,N_7058);
nor U7247 (N_7247,N_7052,N_7198);
xnor U7248 (N_7248,N_7024,N_7199);
nor U7249 (N_7249,N_7031,N_7089);
nor U7250 (N_7250,N_7180,N_7181);
xor U7251 (N_7251,N_7039,N_7140);
nor U7252 (N_7252,N_7124,N_7144);
or U7253 (N_7253,N_7014,N_7064);
xor U7254 (N_7254,N_7189,N_7000);
or U7255 (N_7255,N_7075,N_7093);
or U7256 (N_7256,N_7133,N_7053);
or U7257 (N_7257,N_7003,N_7138);
and U7258 (N_7258,N_7038,N_7027);
xor U7259 (N_7259,N_7010,N_7034);
nand U7260 (N_7260,N_7196,N_7046);
and U7261 (N_7261,N_7148,N_7033);
and U7262 (N_7262,N_7012,N_7197);
or U7263 (N_7263,N_7050,N_7042);
nand U7264 (N_7264,N_7164,N_7048);
nand U7265 (N_7265,N_7007,N_7104);
nand U7266 (N_7266,N_7178,N_7110);
nand U7267 (N_7267,N_7154,N_7184);
and U7268 (N_7268,N_7005,N_7004);
xnor U7269 (N_7269,N_7120,N_7095);
and U7270 (N_7270,N_7071,N_7160);
and U7271 (N_7271,N_7123,N_7121);
or U7272 (N_7272,N_7074,N_7168);
xor U7273 (N_7273,N_7142,N_7112);
and U7274 (N_7274,N_7082,N_7137);
nand U7275 (N_7275,N_7169,N_7028);
or U7276 (N_7276,N_7001,N_7076);
nand U7277 (N_7277,N_7101,N_7020);
and U7278 (N_7278,N_7134,N_7081);
nand U7279 (N_7279,N_7158,N_7040);
nor U7280 (N_7280,N_7106,N_7151);
or U7281 (N_7281,N_7002,N_7009);
xnor U7282 (N_7282,N_7190,N_7153);
xnor U7283 (N_7283,N_7043,N_7139);
or U7284 (N_7284,N_7149,N_7109);
nor U7285 (N_7285,N_7193,N_7035);
or U7286 (N_7286,N_7077,N_7019);
xor U7287 (N_7287,N_7126,N_7097);
or U7288 (N_7288,N_7062,N_7049);
nor U7289 (N_7289,N_7117,N_7170);
and U7290 (N_7290,N_7188,N_7177);
and U7291 (N_7291,N_7094,N_7125);
nor U7292 (N_7292,N_7165,N_7030);
or U7293 (N_7293,N_7118,N_7087);
xor U7294 (N_7294,N_7105,N_7157);
and U7295 (N_7295,N_7015,N_7182);
or U7296 (N_7296,N_7070,N_7098);
or U7297 (N_7297,N_7156,N_7161);
and U7298 (N_7298,N_7122,N_7086);
xnor U7299 (N_7299,N_7136,N_7172);
nand U7300 (N_7300,N_7068,N_7031);
xor U7301 (N_7301,N_7170,N_7010);
or U7302 (N_7302,N_7072,N_7076);
nand U7303 (N_7303,N_7130,N_7026);
nand U7304 (N_7304,N_7109,N_7022);
or U7305 (N_7305,N_7030,N_7088);
or U7306 (N_7306,N_7134,N_7099);
and U7307 (N_7307,N_7121,N_7152);
or U7308 (N_7308,N_7142,N_7015);
xor U7309 (N_7309,N_7194,N_7198);
xor U7310 (N_7310,N_7048,N_7180);
nand U7311 (N_7311,N_7109,N_7091);
nor U7312 (N_7312,N_7069,N_7102);
or U7313 (N_7313,N_7175,N_7164);
nor U7314 (N_7314,N_7154,N_7159);
nor U7315 (N_7315,N_7059,N_7066);
or U7316 (N_7316,N_7140,N_7102);
nor U7317 (N_7317,N_7040,N_7154);
xnor U7318 (N_7318,N_7081,N_7069);
or U7319 (N_7319,N_7094,N_7066);
and U7320 (N_7320,N_7159,N_7146);
nand U7321 (N_7321,N_7008,N_7099);
nor U7322 (N_7322,N_7035,N_7062);
nand U7323 (N_7323,N_7028,N_7145);
and U7324 (N_7324,N_7107,N_7192);
nand U7325 (N_7325,N_7167,N_7008);
and U7326 (N_7326,N_7077,N_7022);
nand U7327 (N_7327,N_7120,N_7103);
or U7328 (N_7328,N_7127,N_7149);
xnor U7329 (N_7329,N_7037,N_7147);
nand U7330 (N_7330,N_7022,N_7179);
nand U7331 (N_7331,N_7001,N_7075);
nand U7332 (N_7332,N_7088,N_7199);
nand U7333 (N_7333,N_7119,N_7141);
xor U7334 (N_7334,N_7035,N_7033);
nand U7335 (N_7335,N_7057,N_7198);
and U7336 (N_7336,N_7064,N_7051);
nor U7337 (N_7337,N_7014,N_7139);
xor U7338 (N_7338,N_7113,N_7080);
xor U7339 (N_7339,N_7020,N_7185);
nor U7340 (N_7340,N_7116,N_7119);
or U7341 (N_7341,N_7038,N_7015);
nor U7342 (N_7342,N_7177,N_7027);
xnor U7343 (N_7343,N_7045,N_7166);
xor U7344 (N_7344,N_7158,N_7061);
nor U7345 (N_7345,N_7197,N_7148);
or U7346 (N_7346,N_7127,N_7181);
nand U7347 (N_7347,N_7024,N_7033);
xor U7348 (N_7348,N_7116,N_7192);
or U7349 (N_7349,N_7059,N_7013);
and U7350 (N_7350,N_7075,N_7124);
or U7351 (N_7351,N_7128,N_7025);
and U7352 (N_7352,N_7009,N_7131);
and U7353 (N_7353,N_7114,N_7034);
nor U7354 (N_7354,N_7147,N_7124);
and U7355 (N_7355,N_7081,N_7090);
and U7356 (N_7356,N_7138,N_7130);
or U7357 (N_7357,N_7028,N_7024);
xor U7358 (N_7358,N_7139,N_7167);
and U7359 (N_7359,N_7035,N_7006);
xor U7360 (N_7360,N_7003,N_7136);
xor U7361 (N_7361,N_7008,N_7198);
or U7362 (N_7362,N_7152,N_7067);
nand U7363 (N_7363,N_7040,N_7001);
xor U7364 (N_7364,N_7195,N_7120);
nor U7365 (N_7365,N_7056,N_7072);
xor U7366 (N_7366,N_7166,N_7012);
and U7367 (N_7367,N_7101,N_7062);
or U7368 (N_7368,N_7144,N_7080);
or U7369 (N_7369,N_7067,N_7098);
nand U7370 (N_7370,N_7008,N_7012);
nor U7371 (N_7371,N_7086,N_7167);
nand U7372 (N_7372,N_7074,N_7106);
and U7373 (N_7373,N_7184,N_7119);
xnor U7374 (N_7374,N_7082,N_7099);
and U7375 (N_7375,N_7177,N_7169);
or U7376 (N_7376,N_7184,N_7127);
nand U7377 (N_7377,N_7185,N_7145);
xor U7378 (N_7378,N_7039,N_7068);
nand U7379 (N_7379,N_7176,N_7099);
or U7380 (N_7380,N_7186,N_7008);
or U7381 (N_7381,N_7033,N_7072);
or U7382 (N_7382,N_7127,N_7002);
or U7383 (N_7383,N_7199,N_7152);
nor U7384 (N_7384,N_7060,N_7071);
nor U7385 (N_7385,N_7055,N_7177);
xnor U7386 (N_7386,N_7150,N_7048);
nor U7387 (N_7387,N_7059,N_7121);
xnor U7388 (N_7388,N_7188,N_7019);
or U7389 (N_7389,N_7044,N_7038);
and U7390 (N_7390,N_7052,N_7105);
and U7391 (N_7391,N_7124,N_7038);
or U7392 (N_7392,N_7144,N_7074);
xnor U7393 (N_7393,N_7005,N_7060);
nor U7394 (N_7394,N_7178,N_7150);
and U7395 (N_7395,N_7067,N_7144);
xor U7396 (N_7396,N_7126,N_7066);
and U7397 (N_7397,N_7005,N_7155);
and U7398 (N_7398,N_7130,N_7199);
or U7399 (N_7399,N_7004,N_7150);
xnor U7400 (N_7400,N_7281,N_7306);
nand U7401 (N_7401,N_7216,N_7270);
and U7402 (N_7402,N_7315,N_7239);
xnor U7403 (N_7403,N_7250,N_7334);
nand U7404 (N_7404,N_7246,N_7266);
or U7405 (N_7405,N_7273,N_7272);
and U7406 (N_7406,N_7206,N_7292);
nor U7407 (N_7407,N_7257,N_7202);
or U7408 (N_7408,N_7370,N_7307);
or U7409 (N_7409,N_7319,N_7209);
nand U7410 (N_7410,N_7230,N_7219);
nand U7411 (N_7411,N_7335,N_7236);
xor U7412 (N_7412,N_7278,N_7240);
nand U7413 (N_7413,N_7215,N_7291);
xnor U7414 (N_7414,N_7271,N_7325);
nor U7415 (N_7415,N_7374,N_7204);
xor U7416 (N_7416,N_7386,N_7346);
nor U7417 (N_7417,N_7352,N_7289);
nor U7418 (N_7418,N_7213,N_7262);
nand U7419 (N_7419,N_7380,N_7345);
nor U7420 (N_7420,N_7222,N_7221);
or U7421 (N_7421,N_7212,N_7310);
xor U7422 (N_7422,N_7354,N_7260);
xnor U7423 (N_7423,N_7338,N_7397);
and U7424 (N_7424,N_7234,N_7360);
nand U7425 (N_7425,N_7347,N_7376);
nor U7426 (N_7426,N_7332,N_7235);
nand U7427 (N_7427,N_7339,N_7369);
or U7428 (N_7428,N_7264,N_7207);
or U7429 (N_7429,N_7241,N_7217);
and U7430 (N_7430,N_7284,N_7329);
nand U7431 (N_7431,N_7205,N_7247);
and U7432 (N_7432,N_7224,N_7201);
xnor U7433 (N_7433,N_7259,N_7277);
xnor U7434 (N_7434,N_7309,N_7210);
nor U7435 (N_7435,N_7223,N_7242);
nor U7436 (N_7436,N_7320,N_7237);
or U7437 (N_7437,N_7378,N_7274);
nand U7438 (N_7438,N_7389,N_7294);
nor U7439 (N_7439,N_7233,N_7293);
and U7440 (N_7440,N_7313,N_7364);
nor U7441 (N_7441,N_7256,N_7381);
nor U7442 (N_7442,N_7371,N_7361);
or U7443 (N_7443,N_7318,N_7349);
xor U7444 (N_7444,N_7363,N_7341);
and U7445 (N_7445,N_7392,N_7308);
nand U7446 (N_7446,N_7228,N_7254);
and U7447 (N_7447,N_7220,N_7385);
nand U7448 (N_7448,N_7387,N_7323);
and U7449 (N_7449,N_7253,N_7322);
nor U7450 (N_7450,N_7314,N_7229);
or U7451 (N_7451,N_7303,N_7261);
and U7452 (N_7452,N_7214,N_7382);
and U7453 (N_7453,N_7280,N_7298);
xor U7454 (N_7454,N_7267,N_7227);
nand U7455 (N_7455,N_7342,N_7357);
nand U7456 (N_7456,N_7203,N_7226);
nand U7457 (N_7457,N_7299,N_7359);
xnor U7458 (N_7458,N_7383,N_7248);
or U7459 (N_7459,N_7343,N_7321);
and U7460 (N_7460,N_7398,N_7288);
xnor U7461 (N_7461,N_7311,N_7328);
xnor U7462 (N_7462,N_7336,N_7379);
xor U7463 (N_7463,N_7393,N_7396);
xnor U7464 (N_7464,N_7208,N_7218);
or U7465 (N_7465,N_7367,N_7331);
nand U7466 (N_7466,N_7375,N_7252);
nand U7467 (N_7467,N_7211,N_7305);
or U7468 (N_7468,N_7317,N_7324);
or U7469 (N_7469,N_7268,N_7388);
nand U7470 (N_7470,N_7290,N_7344);
nand U7471 (N_7471,N_7285,N_7337);
nor U7472 (N_7472,N_7368,N_7304);
or U7473 (N_7473,N_7394,N_7286);
and U7474 (N_7474,N_7263,N_7300);
xor U7475 (N_7475,N_7244,N_7238);
or U7476 (N_7476,N_7316,N_7312);
or U7477 (N_7477,N_7279,N_7399);
or U7478 (N_7478,N_7333,N_7355);
and U7479 (N_7479,N_7348,N_7326);
xor U7480 (N_7480,N_7255,N_7231);
xnor U7481 (N_7481,N_7225,N_7296);
nand U7482 (N_7482,N_7249,N_7391);
xnor U7483 (N_7483,N_7362,N_7275);
nor U7484 (N_7484,N_7356,N_7340);
nand U7485 (N_7485,N_7365,N_7327);
nor U7486 (N_7486,N_7350,N_7390);
or U7487 (N_7487,N_7297,N_7377);
nand U7488 (N_7488,N_7200,N_7373);
and U7489 (N_7489,N_7302,N_7351);
nand U7490 (N_7490,N_7245,N_7384);
nand U7491 (N_7491,N_7243,N_7372);
nor U7492 (N_7492,N_7287,N_7276);
nand U7493 (N_7493,N_7258,N_7282);
and U7494 (N_7494,N_7358,N_7353);
xnor U7495 (N_7495,N_7330,N_7366);
xor U7496 (N_7496,N_7269,N_7301);
nor U7497 (N_7497,N_7283,N_7395);
nand U7498 (N_7498,N_7295,N_7265);
xor U7499 (N_7499,N_7251,N_7232);
and U7500 (N_7500,N_7324,N_7350);
nor U7501 (N_7501,N_7374,N_7227);
nand U7502 (N_7502,N_7360,N_7313);
or U7503 (N_7503,N_7297,N_7318);
nand U7504 (N_7504,N_7205,N_7312);
nor U7505 (N_7505,N_7226,N_7375);
or U7506 (N_7506,N_7301,N_7289);
xnor U7507 (N_7507,N_7398,N_7232);
or U7508 (N_7508,N_7389,N_7346);
and U7509 (N_7509,N_7294,N_7267);
and U7510 (N_7510,N_7246,N_7260);
xor U7511 (N_7511,N_7353,N_7360);
and U7512 (N_7512,N_7250,N_7399);
and U7513 (N_7513,N_7284,N_7389);
xnor U7514 (N_7514,N_7238,N_7360);
xor U7515 (N_7515,N_7354,N_7317);
and U7516 (N_7516,N_7379,N_7343);
nand U7517 (N_7517,N_7201,N_7362);
nor U7518 (N_7518,N_7362,N_7237);
xor U7519 (N_7519,N_7365,N_7299);
or U7520 (N_7520,N_7231,N_7284);
nor U7521 (N_7521,N_7233,N_7336);
nand U7522 (N_7522,N_7251,N_7358);
xor U7523 (N_7523,N_7227,N_7213);
nor U7524 (N_7524,N_7221,N_7299);
and U7525 (N_7525,N_7367,N_7229);
xnor U7526 (N_7526,N_7261,N_7256);
nand U7527 (N_7527,N_7382,N_7393);
nor U7528 (N_7528,N_7281,N_7283);
nand U7529 (N_7529,N_7208,N_7205);
nor U7530 (N_7530,N_7366,N_7328);
nor U7531 (N_7531,N_7248,N_7381);
or U7532 (N_7532,N_7217,N_7254);
xnor U7533 (N_7533,N_7337,N_7251);
xor U7534 (N_7534,N_7203,N_7247);
or U7535 (N_7535,N_7300,N_7200);
nor U7536 (N_7536,N_7328,N_7279);
and U7537 (N_7537,N_7283,N_7230);
or U7538 (N_7538,N_7267,N_7218);
or U7539 (N_7539,N_7376,N_7334);
nand U7540 (N_7540,N_7265,N_7387);
or U7541 (N_7541,N_7231,N_7317);
and U7542 (N_7542,N_7290,N_7203);
nand U7543 (N_7543,N_7240,N_7312);
and U7544 (N_7544,N_7326,N_7276);
or U7545 (N_7545,N_7330,N_7211);
xnor U7546 (N_7546,N_7232,N_7378);
nor U7547 (N_7547,N_7231,N_7271);
nor U7548 (N_7548,N_7282,N_7370);
xor U7549 (N_7549,N_7369,N_7310);
or U7550 (N_7550,N_7331,N_7373);
nor U7551 (N_7551,N_7365,N_7210);
xor U7552 (N_7552,N_7246,N_7273);
or U7553 (N_7553,N_7284,N_7383);
or U7554 (N_7554,N_7352,N_7346);
and U7555 (N_7555,N_7237,N_7202);
and U7556 (N_7556,N_7283,N_7305);
xnor U7557 (N_7557,N_7389,N_7373);
nand U7558 (N_7558,N_7333,N_7294);
nor U7559 (N_7559,N_7353,N_7248);
xor U7560 (N_7560,N_7240,N_7230);
nor U7561 (N_7561,N_7281,N_7222);
and U7562 (N_7562,N_7326,N_7287);
xnor U7563 (N_7563,N_7375,N_7330);
xor U7564 (N_7564,N_7269,N_7386);
nor U7565 (N_7565,N_7224,N_7295);
nand U7566 (N_7566,N_7375,N_7249);
and U7567 (N_7567,N_7304,N_7339);
or U7568 (N_7568,N_7364,N_7281);
xnor U7569 (N_7569,N_7368,N_7310);
xor U7570 (N_7570,N_7236,N_7215);
xnor U7571 (N_7571,N_7340,N_7302);
xnor U7572 (N_7572,N_7364,N_7262);
xnor U7573 (N_7573,N_7266,N_7249);
xnor U7574 (N_7574,N_7296,N_7286);
nor U7575 (N_7575,N_7200,N_7397);
nor U7576 (N_7576,N_7388,N_7298);
or U7577 (N_7577,N_7322,N_7288);
nor U7578 (N_7578,N_7328,N_7363);
nor U7579 (N_7579,N_7293,N_7343);
and U7580 (N_7580,N_7362,N_7329);
nand U7581 (N_7581,N_7308,N_7293);
xor U7582 (N_7582,N_7343,N_7353);
xnor U7583 (N_7583,N_7207,N_7321);
and U7584 (N_7584,N_7336,N_7337);
nor U7585 (N_7585,N_7311,N_7312);
or U7586 (N_7586,N_7223,N_7299);
nor U7587 (N_7587,N_7230,N_7326);
xor U7588 (N_7588,N_7392,N_7312);
nor U7589 (N_7589,N_7219,N_7257);
nor U7590 (N_7590,N_7226,N_7362);
nand U7591 (N_7591,N_7381,N_7209);
and U7592 (N_7592,N_7276,N_7333);
xnor U7593 (N_7593,N_7286,N_7259);
xor U7594 (N_7594,N_7250,N_7313);
xnor U7595 (N_7595,N_7358,N_7226);
and U7596 (N_7596,N_7243,N_7205);
nand U7597 (N_7597,N_7258,N_7222);
and U7598 (N_7598,N_7232,N_7327);
or U7599 (N_7599,N_7383,N_7217);
and U7600 (N_7600,N_7566,N_7457);
xnor U7601 (N_7601,N_7431,N_7515);
or U7602 (N_7602,N_7425,N_7408);
and U7603 (N_7603,N_7534,N_7502);
nor U7604 (N_7604,N_7568,N_7477);
xor U7605 (N_7605,N_7591,N_7407);
nand U7606 (N_7606,N_7553,N_7433);
or U7607 (N_7607,N_7449,N_7590);
nor U7608 (N_7608,N_7558,N_7466);
nor U7609 (N_7609,N_7528,N_7594);
xor U7610 (N_7610,N_7579,N_7587);
and U7611 (N_7611,N_7450,N_7514);
nor U7612 (N_7612,N_7415,N_7420);
xor U7613 (N_7613,N_7578,N_7496);
or U7614 (N_7614,N_7435,N_7512);
and U7615 (N_7615,N_7479,N_7539);
xnor U7616 (N_7616,N_7423,N_7405);
nand U7617 (N_7617,N_7453,N_7441);
and U7618 (N_7618,N_7552,N_7540);
and U7619 (N_7619,N_7555,N_7464);
or U7620 (N_7620,N_7560,N_7535);
and U7621 (N_7621,N_7537,N_7510);
nand U7622 (N_7622,N_7522,N_7509);
nand U7623 (N_7623,N_7513,N_7478);
xor U7624 (N_7624,N_7440,N_7419);
and U7625 (N_7625,N_7462,N_7572);
xnor U7626 (N_7626,N_7442,N_7546);
or U7627 (N_7627,N_7593,N_7575);
nand U7628 (N_7628,N_7417,N_7573);
nand U7629 (N_7629,N_7469,N_7526);
nand U7630 (N_7630,N_7421,N_7556);
xor U7631 (N_7631,N_7564,N_7549);
and U7632 (N_7632,N_7489,N_7503);
nor U7633 (N_7633,N_7404,N_7411);
and U7634 (N_7634,N_7451,N_7460);
or U7635 (N_7635,N_7544,N_7493);
nand U7636 (N_7636,N_7530,N_7481);
nor U7637 (N_7637,N_7531,N_7452);
nor U7638 (N_7638,N_7585,N_7444);
nand U7639 (N_7639,N_7467,N_7589);
and U7640 (N_7640,N_7427,N_7559);
or U7641 (N_7641,N_7519,N_7429);
xor U7642 (N_7642,N_7500,N_7548);
nor U7643 (N_7643,N_7584,N_7463);
nand U7644 (N_7644,N_7545,N_7508);
xor U7645 (N_7645,N_7538,N_7474);
or U7646 (N_7646,N_7565,N_7482);
nand U7647 (N_7647,N_7426,N_7468);
xnor U7648 (N_7648,N_7569,N_7438);
xor U7649 (N_7649,N_7458,N_7413);
or U7650 (N_7650,N_7432,N_7434);
or U7651 (N_7651,N_7486,N_7582);
xnor U7652 (N_7652,N_7583,N_7504);
or U7653 (N_7653,N_7542,N_7445);
and U7654 (N_7654,N_7588,N_7473);
and U7655 (N_7655,N_7499,N_7595);
and U7656 (N_7656,N_7581,N_7492);
nor U7657 (N_7657,N_7495,N_7505);
or U7658 (N_7658,N_7485,N_7401);
or U7659 (N_7659,N_7497,N_7580);
and U7660 (N_7660,N_7567,N_7576);
and U7661 (N_7661,N_7570,N_7416);
and U7662 (N_7662,N_7527,N_7557);
nand U7663 (N_7663,N_7574,N_7409);
and U7664 (N_7664,N_7472,N_7551);
nor U7665 (N_7665,N_7403,N_7506);
nor U7666 (N_7666,N_7488,N_7471);
and U7667 (N_7667,N_7533,N_7521);
and U7668 (N_7668,N_7571,N_7597);
nand U7669 (N_7669,N_7418,N_7428);
xor U7670 (N_7670,N_7524,N_7443);
and U7671 (N_7671,N_7554,N_7596);
nor U7672 (N_7672,N_7518,N_7547);
or U7673 (N_7673,N_7446,N_7586);
or U7674 (N_7674,N_7498,N_7599);
nor U7675 (N_7675,N_7541,N_7454);
nand U7676 (N_7676,N_7465,N_7563);
nor U7677 (N_7677,N_7414,N_7523);
nand U7678 (N_7678,N_7550,N_7592);
nand U7679 (N_7679,N_7529,N_7536);
or U7680 (N_7680,N_7475,N_7484);
xnor U7681 (N_7681,N_7410,N_7470);
xor U7682 (N_7682,N_7487,N_7491);
xnor U7683 (N_7683,N_7422,N_7447);
nor U7684 (N_7684,N_7439,N_7412);
xor U7685 (N_7685,N_7437,N_7402);
xor U7686 (N_7686,N_7461,N_7455);
or U7687 (N_7687,N_7490,N_7483);
xor U7688 (N_7688,N_7476,N_7562);
nor U7689 (N_7689,N_7480,N_7516);
and U7690 (N_7690,N_7511,N_7501);
nor U7691 (N_7691,N_7424,N_7436);
nand U7692 (N_7692,N_7532,N_7543);
nor U7693 (N_7693,N_7525,N_7456);
nand U7694 (N_7694,N_7507,N_7561);
nor U7695 (N_7695,N_7406,N_7459);
nand U7696 (N_7696,N_7598,N_7430);
nor U7697 (N_7697,N_7494,N_7577);
or U7698 (N_7698,N_7517,N_7448);
nand U7699 (N_7699,N_7520,N_7400);
and U7700 (N_7700,N_7456,N_7533);
and U7701 (N_7701,N_7414,N_7446);
and U7702 (N_7702,N_7433,N_7496);
xnor U7703 (N_7703,N_7589,N_7478);
nand U7704 (N_7704,N_7478,N_7476);
nor U7705 (N_7705,N_7482,N_7517);
nand U7706 (N_7706,N_7527,N_7526);
nor U7707 (N_7707,N_7521,N_7558);
and U7708 (N_7708,N_7579,N_7462);
xnor U7709 (N_7709,N_7420,N_7468);
nor U7710 (N_7710,N_7533,N_7539);
nor U7711 (N_7711,N_7533,N_7422);
nand U7712 (N_7712,N_7493,N_7462);
or U7713 (N_7713,N_7460,N_7497);
xnor U7714 (N_7714,N_7505,N_7509);
or U7715 (N_7715,N_7406,N_7446);
or U7716 (N_7716,N_7430,N_7431);
and U7717 (N_7717,N_7415,N_7583);
xnor U7718 (N_7718,N_7554,N_7520);
and U7719 (N_7719,N_7518,N_7400);
nand U7720 (N_7720,N_7491,N_7471);
nor U7721 (N_7721,N_7472,N_7524);
nand U7722 (N_7722,N_7557,N_7453);
nand U7723 (N_7723,N_7404,N_7560);
and U7724 (N_7724,N_7588,N_7433);
or U7725 (N_7725,N_7409,N_7515);
or U7726 (N_7726,N_7416,N_7491);
nand U7727 (N_7727,N_7457,N_7407);
nand U7728 (N_7728,N_7513,N_7520);
nor U7729 (N_7729,N_7512,N_7514);
and U7730 (N_7730,N_7588,N_7549);
nor U7731 (N_7731,N_7439,N_7565);
or U7732 (N_7732,N_7529,N_7532);
xor U7733 (N_7733,N_7410,N_7506);
and U7734 (N_7734,N_7531,N_7516);
or U7735 (N_7735,N_7559,N_7527);
nor U7736 (N_7736,N_7527,N_7502);
or U7737 (N_7737,N_7435,N_7565);
nand U7738 (N_7738,N_7516,N_7574);
or U7739 (N_7739,N_7448,N_7555);
and U7740 (N_7740,N_7436,N_7592);
xnor U7741 (N_7741,N_7496,N_7509);
nor U7742 (N_7742,N_7454,N_7590);
nand U7743 (N_7743,N_7523,N_7424);
nand U7744 (N_7744,N_7438,N_7419);
or U7745 (N_7745,N_7587,N_7454);
nand U7746 (N_7746,N_7404,N_7403);
nand U7747 (N_7747,N_7528,N_7549);
nor U7748 (N_7748,N_7449,N_7531);
xor U7749 (N_7749,N_7527,N_7588);
nand U7750 (N_7750,N_7536,N_7426);
nand U7751 (N_7751,N_7415,N_7435);
nand U7752 (N_7752,N_7484,N_7511);
xor U7753 (N_7753,N_7415,N_7566);
and U7754 (N_7754,N_7453,N_7569);
or U7755 (N_7755,N_7580,N_7465);
nand U7756 (N_7756,N_7490,N_7512);
and U7757 (N_7757,N_7496,N_7591);
xor U7758 (N_7758,N_7543,N_7509);
and U7759 (N_7759,N_7464,N_7419);
and U7760 (N_7760,N_7423,N_7564);
nand U7761 (N_7761,N_7405,N_7594);
nor U7762 (N_7762,N_7431,N_7448);
nand U7763 (N_7763,N_7427,N_7488);
nand U7764 (N_7764,N_7511,N_7571);
nand U7765 (N_7765,N_7416,N_7544);
nor U7766 (N_7766,N_7450,N_7478);
nand U7767 (N_7767,N_7530,N_7570);
or U7768 (N_7768,N_7463,N_7595);
nand U7769 (N_7769,N_7427,N_7447);
nor U7770 (N_7770,N_7451,N_7569);
and U7771 (N_7771,N_7433,N_7481);
and U7772 (N_7772,N_7494,N_7454);
and U7773 (N_7773,N_7580,N_7529);
xor U7774 (N_7774,N_7455,N_7597);
xnor U7775 (N_7775,N_7444,N_7513);
and U7776 (N_7776,N_7577,N_7497);
nor U7777 (N_7777,N_7530,N_7541);
xnor U7778 (N_7778,N_7449,N_7527);
or U7779 (N_7779,N_7550,N_7533);
and U7780 (N_7780,N_7463,N_7494);
nand U7781 (N_7781,N_7475,N_7538);
nand U7782 (N_7782,N_7409,N_7422);
nor U7783 (N_7783,N_7400,N_7579);
xor U7784 (N_7784,N_7550,N_7598);
xor U7785 (N_7785,N_7421,N_7474);
nand U7786 (N_7786,N_7533,N_7491);
and U7787 (N_7787,N_7505,N_7511);
nor U7788 (N_7788,N_7407,N_7581);
and U7789 (N_7789,N_7502,N_7500);
and U7790 (N_7790,N_7443,N_7578);
or U7791 (N_7791,N_7581,N_7470);
nand U7792 (N_7792,N_7547,N_7466);
nor U7793 (N_7793,N_7560,N_7409);
xnor U7794 (N_7794,N_7583,N_7461);
or U7795 (N_7795,N_7544,N_7506);
xnor U7796 (N_7796,N_7530,N_7473);
nand U7797 (N_7797,N_7472,N_7447);
or U7798 (N_7798,N_7529,N_7478);
nand U7799 (N_7799,N_7533,N_7408);
nor U7800 (N_7800,N_7733,N_7724);
or U7801 (N_7801,N_7760,N_7775);
nor U7802 (N_7802,N_7672,N_7648);
or U7803 (N_7803,N_7638,N_7719);
nor U7804 (N_7804,N_7717,N_7683);
and U7805 (N_7805,N_7787,N_7766);
nor U7806 (N_7806,N_7780,N_7710);
or U7807 (N_7807,N_7688,N_7612);
xnor U7808 (N_7808,N_7636,N_7729);
or U7809 (N_7809,N_7685,N_7742);
and U7810 (N_7810,N_7791,N_7681);
nand U7811 (N_7811,N_7745,N_7796);
and U7812 (N_7812,N_7749,N_7650);
nor U7813 (N_7813,N_7605,N_7631);
nand U7814 (N_7814,N_7794,N_7664);
and U7815 (N_7815,N_7644,N_7614);
nor U7816 (N_7816,N_7726,N_7739);
or U7817 (N_7817,N_7759,N_7736);
xor U7818 (N_7818,N_7767,N_7645);
and U7819 (N_7819,N_7675,N_7676);
nand U7820 (N_7820,N_7769,N_7666);
xor U7821 (N_7821,N_7763,N_7626);
nand U7822 (N_7822,N_7738,N_7754);
nand U7823 (N_7823,N_7623,N_7607);
and U7824 (N_7824,N_7609,N_7669);
or U7825 (N_7825,N_7750,N_7707);
xnor U7826 (N_7826,N_7720,N_7620);
or U7827 (N_7827,N_7723,N_7694);
xor U7828 (N_7828,N_7686,N_7728);
xor U7829 (N_7829,N_7776,N_7658);
and U7830 (N_7830,N_7630,N_7722);
nor U7831 (N_7831,N_7799,N_7655);
nor U7832 (N_7832,N_7735,N_7684);
nand U7833 (N_7833,N_7632,N_7677);
and U7834 (N_7834,N_7639,N_7654);
or U7835 (N_7835,N_7687,N_7696);
nor U7836 (N_7836,N_7792,N_7680);
nand U7837 (N_7837,N_7613,N_7715);
and U7838 (N_7838,N_7627,N_7635);
xor U7839 (N_7839,N_7732,N_7641);
nand U7840 (N_7840,N_7611,N_7712);
xnor U7841 (N_7841,N_7706,N_7716);
nor U7842 (N_7842,N_7662,N_7689);
and U7843 (N_7843,N_7700,N_7621);
nand U7844 (N_7844,N_7744,N_7606);
or U7845 (N_7845,N_7610,N_7771);
nor U7846 (N_7846,N_7778,N_7755);
or U7847 (N_7847,N_7779,N_7603);
nor U7848 (N_7848,N_7757,N_7708);
and U7849 (N_7849,N_7659,N_7622);
or U7850 (N_7850,N_7682,N_7668);
or U7851 (N_7851,N_7774,N_7727);
nor U7852 (N_7852,N_7737,N_7753);
and U7853 (N_7853,N_7643,N_7629);
xor U7854 (N_7854,N_7633,N_7797);
xor U7855 (N_7855,N_7784,N_7725);
xor U7856 (N_7856,N_7673,N_7702);
nand U7857 (N_7857,N_7657,N_7697);
nor U7858 (N_7858,N_7795,N_7785);
xor U7859 (N_7859,N_7798,N_7670);
xor U7860 (N_7860,N_7615,N_7600);
nor U7861 (N_7861,N_7756,N_7768);
nor U7862 (N_7862,N_7730,N_7663);
nor U7863 (N_7863,N_7665,N_7713);
xor U7864 (N_7864,N_7781,N_7741);
and U7865 (N_7865,N_7705,N_7652);
nor U7866 (N_7866,N_7709,N_7698);
xnor U7867 (N_7867,N_7770,N_7695);
nor U7868 (N_7868,N_7762,N_7651);
nor U7869 (N_7869,N_7667,N_7786);
and U7870 (N_7870,N_7616,N_7637);
xor U7871 (N_7871,N_7788,N_7691);
or U7872 (N_7872,N_7747,N_7721);
nor U7873 (N_7873,N_7634,N_7783);
nor U7874 (N_7874,N_7671,N_7625);
xor U7875 (N_7875,N_7758,N_7743);
or U7876 (N_7876,N_7793,N_7678);
and U7877 (N_7877,N_7690,N_7692);
xor U7878 (N_7878,N_7777,N_7772);
nor U7879 (N_7879,N_7602,N_7714);
nor U7880 (N_7880,N_7679,N_7718);
nor U7881 (N_7881,N_7604,N_7765);
or U7882 (N_7882,N_7674,N_7656);
xnor U7883 (N_7883,N_7649,N_7764);
xor U7884 (N_7884,N_7661,N_7618);
xor U7885 (N_7885,N_7731,N_7782);
or U7886 (N_7886,N_7624,N_7790);
xor U7887 (N_7887,N_7711,N_7619);
nor U7888 (N_7888,N_7693,N_7761);
nor U7889 (N_7889,N_7628,N_7746);
and U7890 (N_7890,N_7646,N_7647);
nand U7891 (N_7891,N_7703,N_7617);
xnor U7892 (N_7892,N_7752,N_7701);
and U7893 (N_7893,N_7640,N_7642);
xnor U7894 (N_7894,N_7608,N_7789);
and U7895 (N_7895,N_7653,N_7601);
nor U7896 (N_7896,N_7751,N_7748);
xnor U7897 (N_7897,N_7734,N_7704);
or U7898 (N_7898,N_7740,N_7773);
or U7899 (N_7899,N_7660,N_7699);
nand U7900 (N_7900,N_7661,N_7779);
xnor U7901 (N_7901,N_7720,N_7699);
and U7902 (N_7902,N_7780,N_7770);
or U7903 (N_7903,N_7602,N_7686);
xnor U7904 (N_7904,N_7717,N_7646);
nand U7905 (N_7905,N_7606,N_7605);
and U7906 (N_7906,N_7621,N_7720);
and U7907 (N_7907,N_7794,N_7722);
nand U7908 (N_7908,N_7762,N_7604);
or U7909 (N_7909,N_7641,N_7623);
xnor U7910 (N_7910,N_7700,N_7602);
nor U7911 (N_7911,N_7630,N_7749);
or U7912 (N_7912,N_7710,N_7754);
xor U7913 (N_7913,N_7762,N_7731);
and U7914 (N_7914,N_7670,N_7714);
nand U7915 (N_7915,N_7757,N_7672);
nor U7916 (N_7916,N_7775,N_7764);
nand U7917 (N_7917,N_7675,N_7672);
and U7918 (N_7918,N_7608,N_7743);
xor U7919 (N_7919,N_7674,N_7679);
xnor U7920 (N_7920,N_7769,N_7799);
xnor U7921 (N_7921,N_7727,N_7683);
or U7922 (N_7922,N_7764,N_7663);
or U7923 (N_7923,N_7636,N_7748);
xor U7924 (N_7924,N_7782,N_7675);
or U7925 (N_7925,N_7676,N_7683);
nand U7926 (N_7926,N_7665,N_7641);
or U7927 (N_7927,N_7779,N_7728);
and U7928 (N_7928,N_7753,N_7730);
xnor U7929 (N_7929,N_7797,N_7663);
nand U7930 (N_7930,N_7681,N_7734);
and U7931 (N_7931,N_7777,N_7714);
nor U7932 (N_7932,N_7782,N_7691);
xor U7933 (N_7933,N_7778,N_7767);
and U7934 (N_7934,N_7711,N_7771);
xor U7935 (N_7935,N_7738,N_7669);
nor U7936 (N_7936,N_7614,N_7754);
nand U7937 (N_7937,N_7629,N_7625);
or U7938 (N_7938,N_7798,N_7690);
and U7939 (N_7939,N_7763,N_7620);
nand U7940 (N_7940,N_7674,N_7665);
and U7941 (N_7941,N_7706,N_7777);
nand U7942 (N_7942,N_7712,N_7603);
or U7943 (N_7943,N_7630,N_7606);
or U7944 (N_7944,N_7763,N_7651);
nand U7945 (N_7945,N_7699,N_7662);
or U7946 (N_7946,N_7754,N_7721);
nand U7947 (N_7947,N_7668,N_7735);
nor U7948 (N_7948,N_7766,N_7778);
and U7949 (N_7949,N_7759,N_7782);
nand U7950 (N_7950,N_7659,N_7626);
xor U7951 (N_7951,N_7778,N_7614);
or U7952 (N_7952,N_7619,N_7698);
or U7953 (N_7953,N_7720,N_7765);
nor U7954 (N_7954,N_7605,N_7718);
and U7955 (N_7955,N_7634,N_7636);
or U7956 (N_7956,N_7743,N_7654);
nor U7957 (N_7957,N_7708,N_7733);
and U7958 (N_7958,N_7657,N_7654);
and U7959 (N_7959,N_7610,N_7667);
xnor U7960 (N_7960,N_7683,N_7768);
nor U7961 (N_7961,N_7691,N_7771);
nor U7962 (N_7962,N_7751,N_7722);
xnor U7963 (N_7963,N_7685,N_7773);
and U7964 (N_7964,N_7633,N_7613);
or U7965 (N_7965,N_7667,N_7724);
xor U7966 (N_7966,N_7613,N_7658);
and U7967 (N_7967,N_7612,N_7756);
nor U7968 (N_7968,N_7762,N_7707);
nor U7969 (N_7969,N_7736,N_7761);
xor U7970 (N_7970,N_7699,N_7763);
nor U7971 (N_7971,N_7652,N_7781);
nor U7972 (N_7972,N_7625,N_7637);
and U7973 (N_7973,N_7724,N_7606);
nand U7974 (N_7974,N_7765,N_7775);
nand U7975 (N_7975,N_7707,N_7781);
nand U7976 (N_7976,N_7616,N_7624);
and U7977 (N_7977,N_7702,N_7649);
xnor U7978 (N_7978,N_7695,N_7701);
and U7979 (N_7979,N_7729,N_7639);
and U7980 (N_7980,N_7697,N_7794);
nand U7981 (N_7981,N_7700,N_7687);
and U7982 (N_7982,N_7635,N_7617);
nand U7983 (N_7983,N_7680,N_7668);
nor U7984 (N_7984,N_7645,N_7644);
nor U7985 (N_7985,N_7720,N_7791);
or U7986 (N_7986,N_7703,N_7797);
or U7987 (N_7987,N_7720,N_7647);
xnor U7988 (N_7988,N_7790,N_7747);
nor U7989 (N_7989,N_7645,N_7623);
and U7990 (N_7990,N_7797,N_7679);
nand U7991 (N_7991,N_7640,N_7725);
nor U7992 (N_7992,N_7776,N_7641);
nand U7993 (N_7993,N_7780,N_7705);
xor U7994 (N_7994,N_7772,N_7658);
and U7995 (N_7995,N_7619,N_7640);
nand U7996 (N_7996,N_7675,N_7744);
and U7997 (N_7997,N_7608,N_7700);
or U7998 (N_7998,N_7735,N_7651);
nor U7999 (N_7999,N_7714,N_7746);
nand U8000 (N_8000,N_7888,N_7881);
nor U8001 (N_8001,N_7963,N_7821);
xor U8002 (N_8002,N_7875,N_7907);
nand U8003 (N_8003,N_7988,N_7996);
nand U8004 (N_8004,N_7912,N_7987);
or U8005 (N_8005,N_7946,N_7871);
xnor U8006 (N_8006,N_7842,N_7853);
or U8007 (N_8007,N_7936,N_7860);
nor U8008 (N_8008,N_7990,N_7953);
xor U8009 (N_8009,N_7819,N_7964);
and U8010 (N_8010,N_7920,N_7803);
or U8011 (N_8011,N_7890,N_7976);
nor U8012 (N_8012,N_7802,N_7922);
and U8013 (N_8013,N_7828,N_7816);
nor U8014 (N_8014,N_7809,N_7966);
or U8015 (N_8015,N_7844,N_7868);
nand U8016 (N_8016,N_7902,N_7841);
nand U8017 (N_8017,N_7931,N_7975);
nand U8018 (N_8018,N_7847,N_7956);
nor U8019 (N_8019,N_7858,N_7991);
and U8020 (N_8020,N_7850,N_7983);
nor U8021 (N_8021,N_7883,N_7910);
nor U8022 (N_8022,N_7834,N_7932);
and U8023 (N_8023,N_7807,N_7814);
and U8024 (N_8024,N_7820,N_7977);
nand U8025 (N_8025,N_7954,N_7800);
nor U8026 (N_8026,N_7856,N_7859);
or U8027 (N_8027,N_7862,N_7974);
xnor U8028 (N_8028,N_7864,N_7944);
xor U8029 (N_8029,N_7906,N_7805);
nand U8030 (N_8030,N_7969,N_7855);
nand U8031 (N_8031,N_7827,N_7957);
or U8032 (N_8032,N_7877,N_7926);
nand U8033 (N_8033,N_7942,N_7825);
nor U8034 (N_8034,N_7979,N_7836);
nand U8035 (N_8035,N_7960,N_7846);
xnor U8036 (N_8036,N_7882,N_7921);
and U8037 (N_8037,N_7849,N_7985);
xor U8038 (N_8038,N_7848,N_7812);
or U8039 (N_8039,N_7952,N_7925);
xnor U8040 (N_8040,N_7845,N_7945);
nand U8041 (N_8041,N_7923,N_7895);
nor U8042 (N_8042,N_7880,N_7886);
or U8043 (N_8043,N_7872,N_7801);
nor U8044 (N_8044,N_7951,N_7980);
nor U8045 (N_8045,N_7904,N_7824);
nor U8046 (N_8046,N_7937,N_7822);
nand U8047 (N_8047,N_7998,N_7941);
nand U8048 (N_8048,N_7982,N_7893);
and U8049 (N_8049,N_7823,N_7870);
nand U8050 (N_8050,N_7999,N_7949);
or U8051 (N_8051,N_7894,N_7914);
or U8052 (N_8052,N_7948,N_7815);
nor U8053 (N_8053,N_7986,N_7924);
nand U8054 (N_8054,N_7934,N_7843);
nor U8055 (N_8055,N_7808,N_7971);
or U8056 (N_8056,N_7885,N_7903);
or U8057 (N_8057,N_7935,N_7879);
and U8058 (N_8058,N_7818,N_7909);
xnor U8059 (N_8059,N_7992,N_7826);
nand U8060 (N_8060,N_7984,N_7857);
xnor U8061 (N_8061,N_7835,N_7892);
xnor U8062 (N_8062,N_7867,N_7940);
nor U8063 (N_8063,N_7861,N_7866);
or U8064 (N_8064,N_7968,N_7878);
nand U8065 (N_8065,N_7905,N_7897);
or U8066 (N_8066,N_7947,N_7938);
nand U8067 (N_8067,N_7851,N_7813);
or U8068 (N_8068,N_7967,N_7919);
nor U8069 (N_8069,N_7865,N_7959);
nand U8070 (N_8070,N_7943,N_7831);
nor U8071 (N_8071,N_7874,N_7939);
nor U8072 (N_8072,N_7927,N_7928);
xnor U8073 (N_8073,N_7899,N_7917);
nand U8074 (N_8074,N_7840,N_7911);
nand U8075 (N_8075,N_7804,N_7854);
and U8076 (N_8076,N_7933,N_7833);
nand U8077 (N_8077,N_7981,N_7852);
or U8078 (N_8078,N_7916,N_7901);
nand U8079 (N_8079,N_7989,N_7950);
nand U8080 (N_8080,N_7973,N_7955);
xnor U8081 (N_8081,N_7900,N_7806);
xnor U8082 (N_8082,N_7930,N_7962);
or U8083 (N_8083,N_7863,N_7997);
xnor U8084 (N_8084,N_7972,N_7913);
xor U8085 (N_8085,N_7993,N_7958);
and U8086 (N_8086,N_7811,N_7994);
xor U8087 (N_8087,N_7965,N_7832);
nand U8088 (N_8088,N_7891,N_7838);
xnor U8089 (N_8089,N_7837,N_7978);
or U8090 (N_8090,N_7908,N_7961);
nand U8091 (N_8091,N_7876,N_7810);
or U8092 (N_8092,N_7839,N_7929);
and U8093 (N_8093,N_7830,N_7887);
nand U8094 (N_8094,N_7896,N_7995);
or U8095 (N_8095,N_7970,N_7869);
and U8096 (N_8096,N_7898,N_7915);
or U8097 (N_8097,N_7817,N_7884);
nand U8098 (N_8098,N_7873,N_7889);
and U8099 (N_8099,N_7918,N_7829);
and U8100 (N_8100,N_7887,N_7969);
xor U8101 (N_8101,N_7842,N_7890);
nand U8102 (N_8102,N_7917,N_7862);
nand U8103 (N_8103,N_7940,N_7844);
and U8104 (N_8104,N_7802,N_7844);
nand U8105 (N_8105,N_7872,N_7843);
nand U8106 (N_8106,N_7857,N_7963);
xor U8107 (N_8107,N_7800,N_7920);
nand U8108 (N_8108,N_7860,N_7888);
or U8109 (N_8109,N_7912,N_7902);
xor U8110 (N_8110,N_7846,N_7999);
nor U8111 (N_8111,N_7935,N_7936);
or U8112 (N_8112,N_7998,N_7873);
nor U8113 (N_8113,N_7919,N_7957);
nand U8114 (N_8114,N_7856,N_7871);
or U8115 (N_8115,N_7977,N_7837);
nor U8116 (N_8116,N_7834,N_7929);
nand U8117 (N_8117,N_7859,N_7945);
or U8118 (N_8118,N_7947,N_7880);
xor U8119 (N_8119,N_7908,N_7948);
or U8120 (N_8120,N_7868,N_7869);
nand U8121 (N_8121,N_7838,N_7839);
xnor U8122 (N_8122,N_7958,N_7851);
or U8123 (N_8123,N_7907,N_7886);
nand U8124 (N_8124,N_7946,N_7992);
xnor U8125 (N_8125,N_7919,N_7864);
nand U8126 (N_8126,N_7823,N_7814);
or U8127 (N_8127,N_7820,N_7877);
xnor U8128 (N_8128,N_7924,N_7823);
nor U8129 (N_8129,N_7929,N_7873);
and U8130 (N_8130,N_7826,N_7943);
and U8131 (N_8131,N_7935,N_7919);
xor U8132 (N_8132,N_7890,N_7872);
or U8133 (N_8133,N_7884,N_7818);
nand U8134 (N_8134,N_7924,N_7999);
nor U8135 (N_8135,N_7828,N_7946);
nor U8136 (N_8136,N_7844,N_7893);
or U8137 (N_8137,N_7840,N_7927);
or U8138 (N_8138,N_7939,N_7818);
and U8139 (N_8139,N_7971,N_7953);
nand U8140 (N_8140,N_7906,N_7900);
nand U8141 (N_8141,N_7934,N_7885);
or U8142 (N_8142,N_7996,N_7911);
and U8143 (N_8143,N_7822,N_7847);
nand U8144 (N_8144,N_7888,N_7935);
or U8145 (N_8145,N_7938,N_7863);
xor U8146 (N_8146,N_7924,N_7852);
nand U8147 (N_8147,N_7965,N_7942);
and U8148 (N_8148,N_7806,N_7846);
nand U8149 (N_8149,N_7923,N_7869);
and U8150 (N_8150,N_7883,N_7929);
xor U8151 (N_8151,N_7920,N_7991);
nor U8152 (N_8152,N_7966,N_7978);
nor U8153 (N_8153,N_7974,N_7904);
or U8154 (N_8154,N_7816,N_7893);
and U8155 (N_8155,N_7804,N_7957);
nand U8156 (N_8156,N_7916,N_7937);
nand U8157 (N_8157,N_7906,N_7859);
nand U8158 (N_8158,N_7858,N_7854);
or U8159 (N_8159,N_7937,N_7876);
xor U8160 (N_8160,N_7975,N_7986);
nor U8161 (N_8161,N_7952,N_7802);
and U8162 (N_8162,N_7923,N_7976);
and U8163 (N_8163,N_7852,N_7891);
nor U8164 (N_8164,N_7950,N_7895);
or U8165 (N_8165,N_7806,N_7885);
nor U8166 (N_8166,N_7844,N_7815);
nor U8167 (N_8167,N_7894,N_7801);
or U8168 (N_8168,N_7901,N_7969);
and U8169 (N_8169,N_7835,N_7802);
or U8170 (N_8170,N_7969,N_7937);
nand U8171 (N_8171,N_7955,N_7964);
nand U8172 (N_8172,N_7829,N_7894);
or U8173 (N_8173,N_7984,N_7825);
or U8174 (N_8174,N_7949,N_7954);
nand U8175 (N_8175,N_7880,N_7998);
xnor U8176 (N_8176,N_7866,N_7813);
nor U8177 (N_8177,N_7911,N_7922);
xnor U8178 (N_8178,N_7930,N_7959);
and U8179 (N_8179,N_7980,N_7913);
or U8180 (N_8180,N_7936,N_7908);
nor U8181 (N_8181,N_7918,N_7827);
nor U8182 (N_8182,N_7944,N_7827);
nand U8183 (N_8183,N_7903,N_7859);
xnor U8184 (N_8184,N_7922,N_7847);
nor U8185 (N_8185,N_7930,N_7949);
nor U8186 (N_8186,N_7813,N_7903);
or U8187 (N_8187,N_7852,N_7953);
and U8188 (N_8188,N_7823,N_7819);
nor U8189 (N_8189,N_7827,N_7946);
and U8190 (N_8190,N_7844,N_7816);
xnor U8191 (N_8191,N_7950,N_7977);
nand U8192 (N_8192,N_7961,N_7946);
and U8193 (N_8193,N_7870,N_7918);
xnor U8194 (N_8194,N_7944,N_7852);
nor U8195 (N_8195,N_7900,N_7922);
nor U8196 (N_8196,N_7968,N_7930);
xnor U8197 (N_8197,N_7944,N_7871);
and U8198 (N_8198,N_7884,N_7935);
nand U8199 (N_8199,N_7960,N_7955);
nand U8200 (N_8200,N_8096,N_8026);
or U8201 (N_8201,N_8065,N_8048);
nor U8202 (N_8202,N_8138,N_8010);
and U8203 (N_8203,N_8066,N_8140);
nand U8204 (N_8204,N_8106,N_8193);
xor U8205 (N_8205,N_8086,N_8017);
and U8206 (N_8206,N_8003,N_8141);
xnor U8207 (N_8207,N_8186,N_8071);
xor U8208 (N_8208,N_8197,N_8150);
nor U8209 (N_8209,N_8101,N_8185);
and U8210 (N_8210,N_8155,N_8161);
nand U8211 (N_8211,N_8131,N_8002);
xor U8212 (N_8212,N_8173,N_8180);
nor U8213 (N_8213,N_8135,N_8073);
or U8214 (N_8214,N_8108,N_8023);
nand U8215 (N_8215,N_8132,N_8170);
and U8216 (N_8216,N_8184,N_8178);
or U8217 (N_8217,N_8063,N_8092);
or U8218 (N_8218,N_8115,N_8041);
and U8219 (N_8219,N_8129,N_8085);
nand U8220 (N_8220,N_8008,N_8105);
or U8221 (N_8221,N_8147,N_8035);
nor U8222 (N_8222,N_8036,N_8179);
and U8223 (N_8223,N_8011,N_8081);
or U8224 (N_8224,N_8089,N_8118);
xnor U8225 (N_8225,N_8083,N_8004);
and U8226 (N_8226,N_8014,N_8049);
and U8227 (N_8227,N_8075,N_8022);
and U8228 (N_8228,N_8149,N_8121);
xnor U8229 (N_8229,N_8055,N_8152);
nor U8230 (N_8230,N_8124,N_8039);
nor U8231 (N_8231,N_8166,N_8056);
nor U8232 (N_8232,N_8126,N_8069);
nor U8233 (N_8233,N_8006,N_8163);
and U8234 (N_8234,N_8146,N_8079);
or U8235 (N_8235,N_8028,N_8052);
nand U8236 (N_8236,N_8188,N_8187);
xor U8237 (N_8237,N_8076,N_8154);
nor U8238 (N_8238,N_8169,N_8198);
or U8239 (N_8239,N_8134,N_8088);
nor U8240 (N_8240,N_8156,N_8040);
nor U8241 (N_8241,N_8189,N_8122);
or U8242 (N_8242,N_8031,N_8057);
and U8243 (N_8243,N_8018,N_8177);
or U8244 (N_8244,N_8133,N_8125);
nor U8245 (N_8245,N_8142,N_8045);
or U8246 (N_8246,N_8044,N_8060);
nor U8247 (N_8247,N_8171,N_8194);
nor U8248 (N_8248,N_8054,N_8084);
nor U8249 (N_8249,N_8007,N_8047);
nand U8250 (N_8250,N_8061,N_8137);
xor U8251 (N_8251,N_8144,N_8151);
nand U8252 (N_8252,N_8001,N_8119);
nand U8253 (N_8253,N_8013,N_8114);
xor U8254 (N_8254,N_8080,N_8168);
xor U8255 (N_8255,N_8158,N_8067);
and U8256 (N_8256,N_8062,N_8019);
nand U8257 (N_8257,N_8025,N_8099);
nand U8258 (N_8258,N_8005,N_8127);
nor U8259 (N_8259,N_8094,N_8190);
nand U8260 (N_8260,N_8000,N_8109);
nand U8261 (N_8261,N_8037,N_8090);
nor U8262 (N_8262,N_8033,N_8183);
xnor U8263 (N_8263,N_8059,N_8139);
xnor U8264 (N_8264,N_8091,N_8136);
and U8265 (N_8265,N_8123,N_8087);
or U8266 (N_8266,N_8078,N_8100);
and U8267 (N_8267,N_8012,N_8107);
nand U8268 (N_8268,N_8165,N_8145);
nand U8269 (N_8269,N_8016,N_8064);
nor U8270 (N_8270,N_8191,N_8176);
and U8271 (N_8271,N_8110,N_8162);
or U8272 (N_8272,N_8120,N_8070);
xor U8273 (N_8273,N_8172,N_8074);
xnor U8274 (N_8274,N_8116,N_8153);
xnor U8275 (N_8275,N_8046,N_8042);
or U8276 (N_8276,N_8093,N_8103);
and U8277 (N_8277,N_8192,N_8164);
nand U8278 (N_8278,N_8098,N_8104);
or U8279 (N_8279,N_8175,N_8029);
or U8280 (N_8280,N_8195,N_8053);
nor U8281 (N_8281,N_8182,N_8058);
nor U8282 (N_8282,N_8095,N_8160);
nor U8283 (N_8283,N_8181,N_8097);
or U8284 (N_8284,N_8043,N_8020);
and U8285 (N_8285,N_8174,N_8117);
and U8286 (N_8286,N_8024,N_8112);
and U8287 (N_8287,N_8034,N_8038);
nor U8288 (N_8288,N_8027,N_8015);
or U8289 (N_8289,N_8111,N_8009);
nor U8290 (N_8290,N_8113,N_8032);
nand U8291 (N_8291,N_8030,N_8077);
and U8292 (N_8292,N_8157,N_8050);
xor U8293 (N_8293,N_8159,N_8082);
xor U8294 (N_8294,N_8130,N_8051);
nand U8295 (N_8295,N_8167,N_8196);
nor U8296 (N_8296,N_8143,N_8021);
nor U8297 (N_8297,N_8199,N_8128);
and U8298 (N_8298,N_8148,N_8072);
and U8299 (N_8299,N_8102,N_8068);
xnor U8300 (N_8300,N_8062,N_8045);
nor U8301 (N_8301,N_8069,N_8170);
or U8302 (N_8302,N_8188,N_8143);
xnor U8303 (N_8303,N_8197,N_8098);
or U8304 (N_8304,N_8081,N_8196);
or U8305 (N_8305,N_8062,N_8178);
nor U8306 (N_8306,N_8155,N_8010);
or U8307 (N_8307,N_8174,N_8088);
nor U8308 (N_8308,N_8058,N_8130);
or U8309 (N_8309,N_8076,N_8192);
or U8310 (N_8310,N_8040,N_8139);
nor U8311 (N_8311,N_8176,N_8013);
nor U8312 (N_8312,N_8172,N_8110);
and U8313 (N_8313,N_8070,N_8118);
nor U8314 (N_8314,N_8000,N_8124);
and U8315 (N_8315,N_8108,N_8113);
nand U8316 (N_8316,N_8116,N_8109);
or U8317 (N_8317,N_8151,N_8022);
nand U8318 (N_8318,N_8106,N_8151);
or U8319 (N_8319,N_8134,N_8196);
or U8320 (N_8320,N_8182,N_8012);
nor U8321 (N_8321,N_8040,N_8194);
and U8322 (N_8322,N_8180,N_8135);
and U8323 (N_8323,N_8095,N_8097);
xor U8324 (N_8324,N_8092,N_8081);
xnor U8325 (N_8325,N_8138,N_8127);
and U8326 (N_8326,N_8175,N_8188);
nand U8327 (N_8327,N_8165,N_8060);
xnor U8328 (N_8328,N_8118,N_8021);
nor U8329 (N_8329,N_8060,N_8094);
nor U8330 (N_8330,N_8081,N_8137);
nor U8331 (N_8331,N_8181,N_8160);
or U8332 (N_8332,N_8154,N_8031);
or U8333 (N_8333,N_8017,N_8030);
and U8334 (N_8334,N_8047,N_8144);
nor U8335 (N_8335,N_8018,N_8054);
xor U8336 (N_8336,N_8153,N_8134);
or U8337 (N_8337,N_8130,N_8158);
or U8338 (N_8338,N_8154,N_8088);
xor U8339 (N_8339,N_8004,N_8191);
nor U8340 (N_8340,N_8006,N_8085);
or U8341 (N_8341,N_8024,N_8051);
nor U8342 (N_8342,N_8184,N_8052);
nand U8343 (N_8343,N_8182,N_8151);
and U8344 (N_8344,N_8101,N_8110);
or U8345 (N_8345,N_8176,N_8136);
xnor U8346 (N_8346,N_8020,N_8079);
nand U8347 (N_8347,N_8097,N_8023);
or U8348 (N_8348,N_8020,N_8069);
nand U8349 (N_8349,N_8142,N_8166);
xor U8350 (N_8350,N_8151,N_8143);
or U8351 (N_8351,N_8076,N_8075);
nor U8352 (N_8352,N_8045,N_8133);
and U8353 (N_8353,N_8017,N_8054);
xor U8354 (N_8354,N_8170,N_8061);
or U8355 (N_8355,N_8127,N_8166);
nand U8356 (N_8356,N_8072,N_8016);
xor U8357 (N_8357,N_8001,N_8016);
xor U8358 (N_8358,N_8117,N_8148);
or U8359 (N_8359,N_8084,N_8148);
nand U8360 (N_8360,N_8194,N_8114);
xor U8361 (N_8361,N_8160,N_8012);
nand U8362 (N_8362,N_8058,N_8029);
nor U8363 (N_8363,N_8191,N_8103);
xor U8364 (N_8364,N_8149,N_8092);
or U8365 (N_8365,N_8128,N_8134);
xnor U8366 (N_8366,N_8002,N_8197);
xnor U8367 (N_8367,N_8026,N_8156);
nand U8368 (N_8368,N_8169,N_8164);
xor U8369 (N_8369,N_8084,N_8064);
nand U8370 (N_8370,N_8045,N_8000);
xnor U8371 (N_8371,N_8138,N_8094);
nand U8372 (N_8372,N_8191,N_8139);
nand U8373 (N_8373,N_8008,N_8130);
or U8374 (N_8374,N_8067,N_8177);
and U8375 (N_8375,N_8026,N_8020);
nor U8376 (N_8376,N_8044,N_8013);
or U8377 (N_8377,N_8037,N_8038);
nor U8378 (N_8378,N_8052,N_8015);
nand U8379 (N_8379,N_8048,N_8171);
and U8380 (N_8380,N_8079,N_8157);
nand U8381 (N_8381,N_8153,N_8082);
nand U8382 (N_8382,N_8113,N_8105);
nor U8383 (N_8383,N_8041,N_8031);
nor U8384 (N_8384,N_8089,N_8183);
nor U8385 (N_8385,N_8042,N_8081);
nand U8386 (N_8386,N_8121,N_8196);
and U8387 (N_8387,N_8033,N_8072);
and U8388 (N_8388,N_8149,N_8091);
and U8389 (N_8389,N_8003,N_8006);
and U8390 (N_8390,N_8142,N_8008);
or U8391 (N_8391,N_8023,N_8094);
nor U8392 (N_8392,N_8053,N_8018);
and U8393 (N_8393,N_8029,N_8127);
and U8394 (N_8394,N_8097,N_8153);
and U8395 (N_8395,N_8029,N_8044);
nor U8396 (N_8396,N_8147,N_8170);
nand U8397 (N_8397,N_8090,N_8039);
xnor U8398 (N_8398,N_8176,N_8075);
nand U8399 (N_8399,N_8191,N_8040);
nor U8400 (N_8400,N_8325,N_8238);
nand U8401 (N_8401,N_8387,N_8237);
and U8402 (N_8402,N_8383,N_8294);
or U8403 (N_8403,N_8345,N_8394);
xor U8404 (N_8404,N_8267,N_8228);
xor U8405 (N_8405,N_8232,N_8365);
or U8406 (N_8406,N_8210,N_8209);
nor U8407 (N_8407,N_8310,N_8396);
nand U8408 (N_8408,N_8219,N_8262);
nor U8409 (N_8409,N_8206,N_8271);
or U8410 (N_8410,N_8280,N_8348);
and U8411 (N_8411,N_8249,N_8245);
nor U8412 (N_8412,N_8288,N_8257);
nor U8413 (N_8413,N_8269,N_8374);
and U8414 (N_8414,N_8241,N_8347);
nand U8415 (N_8415,N_8266,N_8373);
and U8416 (N_8416,N_8247,N_8342);
and U8417 (N_8417,N_8334,N_8320);
and U8418 (N_8418,N_8371,N_8358);
nor U8419 (N_8419,N_8290,N_8344);
xor U8420 (N_8420,N_8351,N_8366);
or U8421 (N_8421,N_8355,N_8313);
xnor U8422 (N_8422,N_8328,N_8382);
xor U8423 (N_8423,N_8251,N_8226);
and U8424 (N_8424,N_8263,N_8367);
and U8425 (N_8425,N_8331,N_8312);
nand U8426 (N_8426,N_8399,N_8332);
nor U8427 (N_8427,N_8272,N_8319);
and U8428 (N_8428,N_8281,N_8346);
and U8429 (N_8429,N_8391,N_8393);
and U8430 (N_8430,N_8315,N_8274);
nand U8431 (N_8431,N_8317,N_8341);
or U8432 (N_8432,N_8316,N_8250);
nand U8433 (N_8433,N_8352,N_8392);
and U8434 (N_8434,N_8208,N_8284);
xnor U8435 (N_8435,N_8283,N_8368);
and U8436 (N_8436,N_8212,N_8304);
nand U8437 (N_8437,N_8329,N_8282);
nand U8438 (N_8438,N_8398,N_8216);
and U8439 (N_8439,N_8207,N_8385);
or U8440 (N_8440,N_8203,N_8381);
and U8441 (N_8441,N_8264,N_8268);
and U8442 (N_8442,N_8229,N_8278);
xor U8443 (N_8443,N_8379,N_8301);
nor U8444 (N_8444,N_8397,N_8361);
nor U8445 (N_8445,N_8225,N_8293);
or U8446 (N_8446,N_8298,N_8255);
xor U8447 (N_8447,N_8338,N_8235);
or U8448 (N_8448,N_8380,N_8236);
or U8449 (N_8449,N_8340,N_8299);
and U8450 (N_8450,N_8211,N_8221);
nand U8451 (N_8451,N_8386,N_8200);
and U8452 (N_8452,N_8217,N_8395);
nor U8453 (N_8453,N_8214,N_8307);
xor U8454 (N_8454,N_8343,N_8376);
or U8455 (N_8455,N_8349,N_8285);
or U8456 (N_8456,N_8318,N_8233);
xor U8457 (N_8457,N_8324,N_8305);
or U8458 (N_8458,N_8254,N_8270);
nand U8459 (N_8459,N_8296,N_8370);
and U8460 (N_8460,N_8289,N_8350);
xor U8461 (N_8461,N_8356,N_8357);
nand U8462 (N_8462,N_8260,N_8378);
and U8463 (N_8463,N_8390,N_8323);
nor U8464 (N_8464,N_8248,N_8220);
nand U8465 (N_8465,N_8333,N_8353);
nand U8466 (N_8466,N_8253,N_8375);
and U8467 (N_8467,N_8306,N_8201);
or U8468 (N_8468,N_8292,N_8384);
nor U8469 (N_8469,N_8234,N_8321);
nor U8470 (N_8470,N_8314,N_8388);
xor U8471 (N_8471,N_8279,N_8336);
or U8472 (N_8472,N_8308,N_8327);
xnor U8473 (N_8473,N_8354,N_8243);
and U8474 (N_8474,N_8363,N_8204);
or U8475 (N_8475,N_8256,N_8205);
xnor U8476 (N_8476,N_8300,N_8261);
nor U8477 (N_8477,N_8275,N_8218);
and U8478 (N_8478,N_8252,N_8240);
nor U8479 (N_8479,N_8223,N_8202);
nor U8480 (N_8480,N_8311,N_8227);
xnor U8481 (N_8481,N_8291,N_8295);
or U8482 (N_8482,N_8309,N_8359);
nor U8483 (N_8483,N_8389,N_8360);
and U8484 (N_8484,N_8239,N_8215);
nor U8485 (N_8485,N_8362,N_8246);
xor U8486 (N_8486,N_8302,N_8372);
nand U8487 (N_8487,N_8222,N_8224);
nand U8488 (N_8488,N_8213,N_8322);
nand U8489 (N_8489,N_8258,N_8244);
or U8490 (N_8490,N_8377,N_8330);
or U8491 (N_8491,N_8287,N_8242);
xnor U8492 (N_8492,N_8231,N_8277);
or U8493 (N_8493,N_8335,N_8337);
nand U8494 (N_8494,N_8265,N_8259);
nand U8495 (N_8495,N_8276,N_8364);
or U8496 (N_8496,N_8273,N_8339);
nor U8497 (N_8497,N_8297,N_8369);
or U8498 (N_8498,N_8286,N_8230);
nor U8499 (N_8499,N_8303,N_8326);
xor U8500 (N_8500,N_8306,N_8363);
or U8501 (N_8501,N_8277,N_8366);
xnor U8502 (N_8502,N_8353,N_8298);
and U8503 (N_8503,N_8228,N_8277);
or U8504 (N_8504,N_8361,N_8216);
nand U8505 (N_8505,N_8233,N_8365);
xnor U8506 (N_8506,N_8314,N_8210);
or U8507 (N_8507,N_8277,N_8203);
xnor U8508 (N_8508,N_8321,N_8327);
or U8509 (N_8509,N_8345,N_8277);
xor U8510 (N_8510,N_8378,N_8311);
nor U8511 (N_8511,N_8351,N_8278);
nor U8512 (N_8512,N_8219,N_8384);
or U8513 (N_8513,N_8250,N_8345);
and U8514 (N_8514,N_8272,N_8396);
xor U8515 (N_8515,N_8215,N_8331);
nor U8516 (N_8516,N_8351,N_8232);
nor U8517 (N_8517,N_8382,N_8323);
and U8518 (N_8518,N_8254,N_8383);
or U8519 (N_8519,N_8296,N_8364);
or U8520 (N_8520,N_8233,N_8283);
xnor U8521 (N_8521,N_8382,N_8229);
and U8522 (N_8522,N_8379,N_8382);
nand U8523 (N_8523,N_8307,N_8264);
or U8524 (N_8524,N_8296,N_8315);
xor U8525 (N_8525,N_8238,N_8320);
xor U8526 (N_8526,N_8303,N_8353);
nor U8527 (N_8527,N_8214,N_8388);
xnor U8528 (N_8528,N_8354,N_8245);
nor U8529 (N_8529,N_8395,N_8246);
nor U8530 (N_8530,N_8313,N_8340);
xor U8531 (N_8531,N_8292,N_8319);
nand U8532 (N_8532,N_8266,N_8223);
and U8533 (N_8533,N_8327,N_8239);
nor U8534 (N_8534,N_8393,N_8310);
nand U8535 (N_8535,N_8378,N_8327);
nand U8536 (N_8536,N_8210,N_8276);
nand U8537 (N_8537,N_8373,N_8242);
xor U8538 (N_8538,N_8208,N_8322);
or U8539 (N_8539,N_8259,N_8207);
nor U8540 (N_8540,N_8324,N_8286);
xor U8541 (N_8541,N_8321,N_8367);
nor U8542 (N_8542,N_8282,N_8249);
xor U8543 (N_8543,N_8390,N_8279);
and U8544 (N_8544,N_8372,N_8390);
or U8545 (N_8545,N_8280,N_8271);
and U8546 (N_8546,N_8364,N_8235);
xor U8547 (N_8547,N_8340,N_8253);
or U8548 (N_8548,N_8242,N_8255);
or U8549 (N_8549,N_8237,N_8244);
or U8550 (N_8550,N_8307,N_8219);
nand U8551 (N_8551,N_8289,N_8278);
and U8552 (N_8552,N_8344,N_8308);
or U8553 (N_8553,N_8349,N_8321);
and U8554 (N_8554,N_8213,N_8286);
and U8555 (N_8555,N_8375,N_8343);
nand U8556 (N_8556,N_8310,N_8225);
and U8557 (N_8557,N_8301,N_8313);
nor U8558 (N_8558,N_8334,N_8223);
and U8559 (N_8559,N_8330,N_8320);
xor U8560 (N_8560,N_8391,N_8305);
or U8561 (N_8561,N_8346,N_8290);
xnor U8562 (N_8562,N_8202,N_8218);
nand U8563 (N_8563,N_8270,N_8395);
nor U8564 (N_8564,N_8393,N_8221);
xor U8565 (N_8565,N_8333,N_8268);
nand U8566 (N_8566,N_8247,N_8261);
and U8567 (N_8567,N_8396,N_8325);
xor U8568 (N_8568,N_8292,N_8287);
nand U8569 (N_8569,N_8329,N_8253);
nor U8570 (N_8570,N_8239,N_8234);
nor U8571 (N_8571,N_8303,N_8294);
nand U8572 (N_8572,N_8265,N_8205);
nor U8573 (N_8573,N_8377,N_8301);
nor U8574 (N_8574,N_8261,N_8208);
xor U8575 (N_8575,N_8344,N_8352);
nand U8576 (N_8576,N_8233,N_8353);
or U8577 (N_8577,N_8214,N_8226);
xnor U8578 (N_8578,N_8294,N_8262);
and U8579 (N_8579,N_8318,N_8386);
nand U8580 (N_8580,N_8246,N_8217);
or U8581 (N_8581,N_8272,N_8245);
and U8582 (N_8582,N_8257,N_8221);
nand U8583 (N_8583,N_8397,N_8318);
nand U8584 (N_8584,N_8353,N_8366);
or U8585 (N_8585,N_8394,N_8259);
xnor U8586 (N_8586,N_8393,N_8213);
and U8587 (N_8587,N_8352,N_8324);
and U8588 (N_8588,N_8380,N_8210);
xor U8589 (N_8589,N_8349,N_8367);
xor U8590 (N_8590,N_8351,N_8330);
nor U8591 (N_8591,N_8322,N_8391);
nand U8592 (N_8592,N_8242,N_8203);
xor U8593 (N_8593,N_8240,N_8292);
or U8594 (N_8594,N_8369,N_8292);
xnor U8595 (N_8595,N_8375,N_8370);
xor U8596 (N_8596,N_8369,N_8294);
nand U8597 (N_8597,N_8360,N_8399);
nand U8598 (N_8598,N_8289,N_8218);
nand U8599 (N_8599,N_8205,N_8315);
or U8600 (N_8600,N_8461,N_8589);
nor U8601 (N_8601,N_8582,N_8544);
nor U8602 (N_8602,N_8476,N_8592);
or U8603 (N_8603,N_8401,N_8446);
xnor U8604 (N_8604,N_8411,N_8400);
nand U8605 (N_8605,N_8478,N_8410);
xor U8606 (N_8606,N_8509,N_8429);
nor U8607 (N_8607,N_8523,N_8578);
nand U8608 (N_8608,N_8414,N_8541);
nand U8609 (N_8609,N_8466,N_8535);
or U8610 (N_8610,N_8454,N_8562);
xnor U8611 (N_8611,N_8568,N_8539);
and U8612 (N_8612,N_8576,N_8444);
xnor U8613 (N_8613,N_8525,N_8452);
or U8614 (N_8614,N_8565,N_8448);
xor U8615 (N_8615,N_8551,N_8538);
nand U8616 (N_8616,N_8472,N_8459);
or U8617 (N_8617,N_8458,N_8487);
nor U8618 (N_8618,N_8587,N_8548);
or U8619 (N_8619,N_8475,N_8520);
and U8620 (N_8620,N_8591,N_8517);
nor U8621 (N_8621,N_8464,N_8491);
or U8622 (N_8622,N_8500,N_8564);
or U8623 (N_8623,N_8511,N_8413);
and U8624 (N_8624,N_8490,N_8431);
xnor U8625 (N_8625,N_8501,N_8415);
or U8626 (N_8626,N_8516,N_8424);
and U8627 (N_8627,N_8499,N_8486);
nand U8628 (N_8628,N_8596,N_8566);
xor U8629 (N_8629,N_8572,N_8418);
nor U8630 (N_8630,N_8599,N_8470);
and U8631 (N_8631,N_8494,N_8594);
nand U8632 (N_8632,N_8460,N_8546);
nand U8633 (N_8633,N_8557,N_8412);
nor U8634 (N_8634,N_8570,N_8545);
xor U8635 (N_8635,N_8531,N_8480);
nand U8636 (N_8636,N_8574,N_8498);
nor U8637 (N_8637,N_8507,N_8532);
nor U8638 (N_8638,N_8456,N_8423);
and U8639 (N_8639,N_8484,N_8425);
and U8640 (N_8640,N_8407,N_8518);
nand U8641 (N_8641,N_8477,N_8502);
or U8642 (N_8642,N_8434,N_8467);
xor U8643 (N_8643,N_8543,N_8519);
or U8644 (N_8644,N_8471,N_8584);
nand U8645 (N_8645,N_8438,N_8482);
xnor U8646 (N_8646,N_8526,N_8527);
nand U8647 (N_8647,N_8469,N_8553);
or U8648 (N_8648,N_8581,N_8528);
xor U8649 (N_8649,N_8559,N_8445);
nor U8650 (N_8650,N_8536,N_8510);
xor U8651 (N_8651,N_8497,N_8583);
or U8652 (N_8652,N_8416,N_8503);
nand U8653 (N_8653,N_8549,N_8409);
and U8654 (N_8654,N_8505,N_8512);
xnor U8655 (N_8655,N_8421,N_8463);
or U8656 (N_8656,N_8436,N_8521);
nand U8657 (N_8657,N_8455,N_8428);
nand U8658 (N_8658,N_8427,N_8437);
or U8659 (N_8659,N_8481,N_8558);
or U8660 (N_8660,N_8529,N_8561);
xnor U8661 (N_8661,N_8417,N_8440);
xor U8662 (N_8662,N_8408,N_8493);
nand U8663 (N_8663,N_8524,N_8441);
and U8664 (N_8664,N_8598,N_8547);
xnor U8665 (N_8665,N_8593,N_8595);
nand U8666 (N_8666,N_8406,N_8567);
nand U8667 (N_8667,N_8462,N_8485);
nor U8668 (N_8668,N_8571,N_8468);
nand U8669 (N_8669,N_8569,N_8560);
nor U8670 (N_8670,N_8451,N_8435);
nor U8671 (N_8671,N_8432,N_8439);
nand U8672 (N_8672,N_8530,N_8483);
or U8673 (N_8673,N_8573,N_8496);
nand U8674 (N_8674,N_8449,N_8443);
and U8675 (N_8675,N_8514,N_8474);
or U8676 (N_8676,N_8504,N_8597);
nand U8677 (N_8677,N_8492,N_8508);
xor U8678 (N_8678,N_8457,N_8540);
nor U8679 (N_8679,N_8522,N_8542);
or U8680 (N_8680,N_8402,N_8556);
nand U8681 (N_8681,N_8404,N_8506);
and U8682 (N_8682,N_8495,N_8585);
and U8683 (N_8683,N_8575,N_8554);
nand U8684 (N_8684,N_8513,N_8580);
and U8685 (N_8685,N_8555,N_8420);
nand U8686 (N_8686,N_8405,N_8453);
nand U8687 (N_8687,N_8465,N_8489);
nor U8688 (N_8688,N_8550,N_8426);
xnor U8689 (N_8689,N_8419,N_8515);
xnor U8690 (N_8690,N_8422,N_8590);
nor U8691 (N_8691,N_8473,N_8433);
xor U8692 (N_8692,N_8577,N_8534);
and U8693 (N_8693,N_8447,N_8442);
nand U8694 (N_8694,N_8579,N_8586);
xnor U8695 (N_8695,N_8450,N_8430);
nor U8696 (N_8696,N_8488,N_8588);
nor U8697 (N_8697,N_8537,N_8563);
nand U8698 (N_8698,N_8533,N_8403);
nor U8699 (N_8699,N_8479,N_8552);
xor U8700 (N_8700,N_8546,N_8513);
nand U8701 (N_8701,N_8514,N_8576);
and U8702 (N_8702,N_8533,N_8529);
nor U8703 (N_8703,N_8544,N_8400);
xor U8704 (N_8704,N_8420,N_8463);
and U8705 (N_8705,N_8572,N_8554);
nand U8706 (N_8706,N_8530,N_8516);
nor U8707 (N_8707,N_8467,N_8497);
xor U8708 (N_8708,N_8490,N_8472);
nand U8709 (N_8709,N_8489,N_8477);
and U8710 (N_8710,N_8433,N_8471);
nor U8711 (N_8711,N_8576,N_8529);
xor U8712 (N_8712,N_8472,N_8406);
xor U8713 (N_8713,N_8406,N_8461);
nor U8714 (N_8714,N_8529,N_8596);
and U8715 (N_8715,N_8492,N_8498);
nand U8716 (N_8716,N_8490,N_8476);
and U8717 (N_8717,N_8584,N_8535);
or U8718 (N_8718,N_8559,N_8533);
and U8719 (N_8719,N_8569,N_8406);
or U8720 (N_8720,N_8458,N_8461);
or U8721 (N_8721,N_8570,N_8440);
xor U8722 (N_8722,N_8515,N_8433);
or U8723 (N_8723,N_8426,N_8575);
nand U8724 (N_8724,N_8492,N_8519);
nor U8725 (N_8725,N_8583,N_8526);
nand U8726 (N_8726,N_8434,N_8465);
and U8727 (N_8727,N_8503,N_8442);
nor U8728 (N_8728,N_8527,N_8572);
or U8729 (N_8729,N_8533,N_8589);
xor U8730 (N_8730,N_8441,N_8548);
xnor U8731 (N_8731,N_8514,N_8594);
or U8732 (N_8732,N_8554,N_8574);
xnor U8733 (N_8733,N_8503,N_8412);
xor U8734 (N_8734,N_8422,N_8476);
or U8735 (N_8735,N_8500,N_8506);
and U8736 (N_8736,N_8519,N_8448);
nor U8737 (N_8737,N_8412,N_8421);
or U8738 (N_8738,N_8462,N_8529);
or U8739 (N_8739,N_8582,N_8459);
xnor U8740 (N_8740,N_8432,N_8427);
nor U8741 (N_8741,N_8556,N_8522);
nor U8742 (N_8742,N_8454,N_8501);
or U8743 (N_8743,N_8409,N_8435);
nand U8744 (N_8744,N_8549,N_8555);
xor U8745 (N_8745,N_8566,N_8449);
xor U8746 (N_8746,N_8415,N_8421);
nand U8747 (N_8747,N_8436,N_8493);
nor U8748 (N_8748,N_8492,N_8437);
nor U8749 (N_8749,N_8463,N_8558);
or U8750 (N_8750,N_8547,N_8426);
or U8751 (N_8751,N_8449,N_8541);
nor U8752 (N_8752,N_8417,N_8564);
nand U8753 (N_8753,N_8572,N_8510);
nand U8754 (N_8754,N_8533,N_8495);
or U8755 (N_8755,N_8566,N_8458);
nor U8756 (N_8756,N_8508,N_8514);
or U8757 (N_8757,N_8490,N_8477);
and U8758 (N_8758,N_8443,N_8464);
or U8759 (N_8759,N_8587,N_8454);
and U8760 (N_8760,N_8540,N_8572);
nand U8761 (N_8761,N_8456,N_8411);
and U8762 (N_8762,N_8588,N_8411);
xor U8763 (N_8763,N_8516,N_8418);
xnor U8764 (N_8764,N_8457,N_8404);
nor U8765 (N_8765,N_8576,N_8441);
or U8766 (N_8766,N_8560,N_8426);
nand U8767 (N_8767,N_8566,N_8436);
and U8768 (N_8768,N_8511,N_8577);
nand U8769 (N_8769,N_8551,N_8581);
nand U8770 (N_8770,N_8562,N_8447);
or U8771 (N_8771,N_8529,N_8487);
or U8772 (N_8772,N_8496,N_8449);
xnor U8773 (N_8773,N_8539,N_8476);
and U8774 (N_8774,N_8526,N_8487);
nor U8775 (N_8775,N_8470,N_8476);
nor U8776 (N_8776,N_8557,N_8460);
xor U8777 (N_8777,N_8464,N_8561);
or U8778 (N_8778,N_8443,N_8586);
and U8779 (N_8779,N_8445,N_8410);
and U8780 (N_8780,N_8489,N_8490);
nand U8781 (N_8781,N_8562,N_8509);
nor U8782 (N_8782,N_8595,N_8463);
and U8783 (N_8783,N_8587,N_8475);
and U8784 (N_8784,N_8477,N_8545);
or U8785 (N_8785,N_8523,N_8571);
nor U8786 (N_8786,N_8468,N_8428);
nor U8787 (N_8787,N_8563,N_8455);
or U8788 (N_8788,N_8558,N_8544);
xor U8789 (N_8789,N_8499,N_8521);
or U8790 (N_8790,N_8511,N_8568);
xor U8791 (N_8791,N_8562,N_8495);
and U8792 (N_8792,N_8555,N_8482);
xor U8793 (N_8793,N_8465,N_8591);
xor U8794 (N_8794,N_8591,N_8487);
or U8795 (N_8795,N_8489,N_8515);
nor U8796 (N_8796,N_8558,N_8527);
and U8797 (N_8797,N_8491,N_8537);
and U8798 (N_8798,N_8597,N_8423);
or U8799 (N_8799,N_8539,N_8546);
or U8800 (N_8800,N_8694,N_8655);
nor U8801 (N_8801,N_8781,N_8798);
or U8802 (N_8802,N_8662,N_8706);
or U8803 (N_8803,N_8600,N_8714);
and U8804 (N_8804,N_8792,N_8693);
nand U8805 (N_8805,N_8719,N_8661);
and U8806 (N_8806,N_8635,N_8616);
nor U8807 (N_8807,N_8627,N_8771);
xnor U8808 (N_8808,N_8684,N_8794);
nor U8809 (N_8809,N_8663,N_8727);
or U8810 (N_8810,N_8678,N_8692);
xnor U8811 (N_8811,N_8707,N_8749);
nor U8812 (N_8812,N_8746,N_8710);
and U8813 (N_8813,N_8711,N_8695);
nor U8814 (N_8814,N_8708,N_8732);
xor U8815 (N_8815,N_8772,N_8704);
nand U8816 (N_8816,N_8631,N_8786);
or U8817 (N_8817,N_8670,N_8783);
xor U8818 (N_8818,N_8736,N_8745);
and U8819 (N_8819,N_8741,N_8701);
xor U8820 (N_8820,N_8784,N_8716);
or U8821 (N_8821,N_8766,N_8666);
nand U8822 (N_8822,N_8776,N_8756);
nor U8823 (N_8823,N_8624,N_8737);
or U8824 (N_8824,N_8712,N_8677);
nor U8825 (N_8825,N_8683,N_8744);
or U8826 (N_8826,N_8622,N_8752);
and U8827 (N_8827,N_8601,N_8775);
nand U8828 (N_8828,N_8690,N_8691);
and U8829 (N_8829,N_8636,N_8721);
and U8830 (N_8830,N_8617,N_8672);
nor U8831 (N_8831,N_8671,N_8674);
xnor U8832 (N_8832,N_8688,N_8620);
nand U8833 (N_8833,N_8668,N_8682);
and U8834 (N_8834,N_8687,N_8720);
nand U8835 (N_8835,N_8667,N_8726);
nand U8836 (N_8836,N_8748,N_8757);
nor U8837 (N_8837,N_8614,N_8760);
nand U8838 (N_8838,N_8651,N_8603);
or U8839 (N_8839,N_8669,N_8633);
or U8840 (N_8840,N_8619,N_8640);
or U8841 (N_8841,N_8626,N_8612);
and U8842 (N_8842,N_8686,N_8761);
and U8843 (N_8843,N_8739,N_8785);
or U8844 (N_8844,N_8689,N_8762);
nand U8845 (N_8845,N_8729,N_8625);
or U8846 (N_8846,N_8656,N_8724);
xor U8847 (N_8847,N_8657,N_8638);
xor U8848 (N_8848,N_8782,N_8650);
and U8849 (N_8849,N_8604,N_8702);
and U8850 (N_8850,N_8780,N_8796);
xnor U8851 (N_8851,N_8623,N_8709);
or U8852 (N_8852,N_8607,N_8703);
nor U8853 (N_8853,N_8643,N_8791);
or U8854 (N_8854,N_8725,N_8779);
or U8855 (N_8855,N_8755,N_8613);
nor U8856 (N_8856,N_8773,N_8658);
and U8857 (N_8857,N_8675,N_8673);
and U8858 (N_8858,N_8734,N_8769);
nor U8859 (N_8859,N_8767,N_8676);
xnor U8860 (N_8860,N_8700,N_8774);
xnor U8861 (N_8861,N_8759,N_8758);
nor U8862 (N_8862,N_8634,N_8718);
nand U8863 (N_8863,N_8610,N_8679);
xnor U8864 (N_8864,N_8728,N_8723);
and U8865 (N_8865,N_8750,N_8681);
nand U8866 (N_8866,N_8685,N_8680);
nand U8867 (N_8867,N_8653,N_8713);
xor U8868 (N_8868,N_8615,N_8611);
and U8869 (N_8869,N_8699,N_8664);
nor U8870 (N_8870,N_8799,N_8641);
nor U8871 (N_8871,N_8742,N_8722);
or U8872 (N_8872,N_8637,N_8705);
xor U8873 (N_8873,N_8731,N_8659);
xnor U8874 (N_8874,N_8777,N_8645);
nor U8875 (N_8875,N_8764,N_8618);
nor U8876 (N_8876,N_8738,N_8795);
nor U8877 (N_8877,N_8751,N_8608);
xor U8878 (N_8878,N_8647,N_8628);
nand U8879 (N_8879,N_8793,N_8717);
nand U8880 (N_8880,N_8609,N_8763);
or U8881 (N_8881,N_8765,N_8754);
xnor U8882 (N_8882,N_8629,N_8648);
or U8883 (N_8883,N_8778,N_8715);
or U8884 (N_8884,N_8654,N_8770);
nor U8885 (N_8885,N_8632,N_8698);
and U8886 (N_8886,N_8753,N_8644);
and U8887 (N_8887,N_8660,N_8652);
nor U8888 (N_8888,N_8735,N_8747);
nand U8889 (N_8889,N_8605,N_8768);
xnor U8890 (N_8890,N_8606,N_8642);
and U8891 (N_8891,N_8665,N_8730);
or U8892 (N_8892,N_8788,N_8733);
xnor U8893 (N_8893,N_8787,N_8790);
or U8894 (N_8894,N_8639,N_8797);
xnor U8895 (N_8895,N_8602,N_8789);
xor U8896 (N_8896,N_8743,N_8646);
and U8897 (N_8897,N_8630,N_8621);
or U8898 (N_8898,N_8740,N_8649);
xnor U8899 (N_8899,N_8697,N_8696);
or U8900 (N_8900,N_8647,N_8638);
nor U8901 (N_8901,N_8662,N_8623);
nand U8902 (N_8902,N_8707,N_8735);
and U8903 (N_8903,N_8722,N_8658);
nand U8904 (N_8904,N_8687,N_8729);
and U8905 (N_8905,N_8726,N_8685);
or U8906 (N_8906,N_8656,N_8649);
xor U8907 (N_8907,N_8719,N_8669);
xor U8908 (N_8908,N_8799,N_8789);
nand U8909 (N_8909,N_8778,N_8719);
and U8910 (N_8910,N_8674,N_8639);
or U8911 (N_8911,N_8687,N_8794);
nand U8912 (N_8912,N_8773,N_8713);
nand U8913 (N_8913,N_8724,N_8737);
nor U8914 (N_8914,N_8626,N_8668);
or U8915 (N_8915,N_8771,N_8739);
nor U8916 (N_8916,N_8687,N_8694);
xor U8917 (N_8917,N_8631,N_8688);
or U8918 (N_8918,N_8646,N_8688);
nor U8919 (N_8919,N_8686,N_8715);
or U8920 (N_8920,N_8693,N_8766);
nor U8921 (N_8921,N_8726,N_8724);
nand U8922 (N_8922,N_8683,N_8757);
nand U8923 (N_8923,N_8763,N_8623);
nand U8924 (N_8924,N_8699,N_8771);
and U8925 (N_8925,N_8664,N_8663);
xor U8926 (N_8926,N_8749,N_8627);
and U8927 (N_8927,N_8659,N_8686);
or U8928 (N_8928,N_8659,N_8746);
or U8929 (N_8929,N_8787,N_8641);
and U8930 (N_8930,N_8647,N_8646);
xor U8931 (N_8931,N_8622,N_8692);
and U8932 (N_8932,N_8601,N_8742);
nor U8933 (N_8933,N_8785,N_8764);
xnor U8934 (N_8934,N_8773,N_8739);
nand U8935 (N_8935,N_8754,N_8707);
and U8936 (N_8936,N_8777,N_8706);
xnor U8937 (N_8937,N_8740,N_8689);
or U8938 (N_8938,N_8740,N_8640);
or U8939 (N_8939,N_8726,N_8722);
or U8940 (N_8940,N_8730,N_8602);
nand U8941 (N_8941,N_8690,N_8761);
and U8942 (N_8942,N_8649,N_8688);
nor U8943 (N_8943,N_8742,N_8752);
nand U8944 (N_8944,N_8637,N_8753);
nand U8945 (N_8945,N_8715,N_8796);
xor U8946 (N_8946,N_8736,N_8617);
nand U8947 (N_8947,N_8620,N_8760);
nand U8948 (N_8948,N_8609,N_8672);
and U8949 (N_8949,N_8670,N_8715);
and U8950 (N_8950,N_8682,N_8681);
nor U8951 (N_8951,N_8768,N_8662);
and U8952 (N_8952,N_8693,N_8774);
and U8953 (N_8953,N_8745,N_8781);
xor U8954 (N_8954,N_8645,N_8787);
nor U8955 (N_8955,N_8613,N_8790);
or U8956 (N_8956,N_8683,N_8652);
nand U8957 (N_8957,N_8737,N_8761);
or U8958 (N_8958,N_8792,N_8692);
nor U8959 (N_8959,N_8656,N_8796);
xor U8960 (N_8960,N_8708,N_8794);
nor U8961 (N_8961,N_8692,N_8713);
or U8962 (N_8962,N_8674,N_8613);
nand U8963 (N_8963,N_8651,N_8792);
xnor U8964 (N_8964,N_8662,N_8712);
and U8965 (N_8965,N_8661,N_8757);
nor U8966 (N_8966,N_8601,N_8735);
and U8967 (N_8967,N_8638,N_8736);
nor U8968 (N_8968,N_8691,N_8631);
or U8969 (N_8969,N_8698,N_8768);
nor U8970 (N_8970,N_8783,N_8781);
xnor U8971 (N_8971,N_8659,N_8735);
and U8972 (N_8972,N_8635,N_8753);
nand U8973 (N_8973,N_8795,N_8735);
xnor U8974 (N_8974,N_8788,N_8651);
nand U8975 (N_8975,N_8784,N_8673);
nor U8976 (N_8976,N_8721,N_8744);
nand U8977 (N_8977,N_8670,N_8768);
nor U8978 (N_8978,N_8664,N_8733);
or U8979 (N_8979,N_8655,N_8647);
and U8980 (N_8980,N_8686,N_8702);
nand U8981 (N_8981,N_8609,N_8762);
xnor U8982 (N_8982,N_8755,N_8728);
or U8983 (N_8983,N_8765,N_8629);
or U8984 (N_8984,N_8675,N_8637);
nand U8985 (N_8985,N_8699,N_8735);
or U8986 (N_8986,N_8702,N_8799);
and U8987 (N_8987,N_8746,N_8669);
or U8988 (N_8988,N_8674,N_8716);
and U8989 (N_8989,N_8740,N_8759);
or U8990 (N_8990,N_8619,N_8708);
or U8991 (N_8991,N_8736,N_8623);
nand U8992 (N_8992,N_8702,N_8770);
nand U8993 (N_8993,N_8720,N_8790);
or U8994 (N_8994,N_8705,N_8787);
or U8995 (N_8995,N_8776,N_8728);
xnor U8996 (N_8996,N_8687,N_8664);
nand U8997 (N_8997,N_8798,N_8720);
or U8998 (N_8998,N_8753,N_8671);
nor U8999 (N_8999,N_8662,N_8718);
nor U9000 (N_9000,N_8816,N_8833);
nor U9001 (N_9001,N_8903,N_8807);
nand U9002 (N_9002,N_8978,N_8943);
or U9003 (N_9003,N_8983,N_8990);
nor U9004 (N_9004,N_8805,N_8898);
nor U9005 (N_9005,N_8991,N_8806);
nand U9006 (N_9006,N_8875,N_8956);
nor U9007 (N_9007,N_8947,N_8800);
and U9008 (N_9008,N_8942,N_8926);
or U9009 (N_9009,N_8963,N_8837);
nor U9010 (N_9010,N_8829,N_8873);
nand U9011 (N_9011,N_8899,N_8891);
xor U9012 (N_9012,N_8999,N_8987);
xor U9013 (N_9013,N_8950,N_8901);
or U9014 (N_9014,N_8844,N_8876);
and U9015 (N_9015,N_8962,N_8867);
nor U9016 (N_9016,N_8986,N_8856);
or U9017 (N_9017,N_8985,N_8890);
nor U9018 (N_9018,N_8839,N_8830);
nand U9019 (N_9019,N_8883,N_8984);
nand U9020 (N_9020,N_8927,N_8848);
nor U9021 (N_9021,N_8946,N_8850);
nor U9022 (N_9022,N_8981,N_8923);
xnor U9023 (N_9023,N_8964,N_8851);
nand U9024 (N_9024,N_8976,N_8825);
nand U9025 (N_9025,N_8847,N_8917);
or U9026 (N_9026,N_8842,N_8953);
and U9027 (N_9027,N_8884,N_8911);
nand U9028 (N_9028,N_8860,N_8827);
nand U9029 (N_9029,N_8905,N_8932);
or U9030 (N_9030,N_8886,N_8998);
or U9031 (N_9031,N_8809,N_8889);
xnor U9032 (N_9032,N_8820,N_8938);
and U9033 (N_9033,N_8902,N_8931);
xnor U9034 (N_9034,N_8933,N_8811);
nor U9035 (N_9035,N_8841,N_8817);
and U9036 (N_9036,N_8865,N_8840);
and U9037 (N_9037,N_8893,N_8862);
nand U9038 (N_9038,N_8966,N_8802);
nand U9039 (N_9039,N_8977,N_8913);
nand U9040 (N_9040,N_8975,N_8834);
and U9041 (N_9041,N_8992,N_8871);
xnor U9042 (N_9042,N_8882,N_8852);
nor U9043 (N_9043,N_8965,N_8944);
or U9044 (N_9044,N_8972,N_8878);
or U9045 (N_9045,N_8821,N_8967);
nand U9046 (N_9046,N_8988,N_8995);
xor U9047 (N_9047,N_8858,N_8813);
nand U9048 (N_9048,N_8803,N_8814);
and U9049 (N_9049,N_8912,N_8952);
xnor U9050 (N_9050,N_8900,N_8866);
or U9051 (N_9051,N_8870,N_8974);
nand U9052 (N_9052,N_8872,N_8994);
nand U9053 (N_9053,N_8928,N_8846);
and U9054 (N_9054,N_8887,N_8838);
nand U9055 (N_9055,N_8874,N_8941);
nand U9056 (N_9056,N_8954,N_8973);
nand U9057 (N_9057,N_8831,N_8859);
and U9058 (N_9058,N_8935,N_8969);
nand U9059 (N_9059,N_8921,N_8922);
nand U9060 (N_9060,N_8989,N_8808);
nand U9061 (N_9061,N_8823,N_8864);
and U9062 (N_9062,N_8924,N_8930);
or U9063 (N_9063,N_8957,N_8920);
or U9064 (N_9064,N_8925,N_8949);
nor U9065 (N_9065,N_8877,N_8822);
nand U9066 (N_9066,N_8904,N_8896);
or U9067 (N_9067,N_8948,N_8937);
and U9068 (N_9068,N_8939,N_8940);
nand U9069 (N_9069,N_8951,N_8826);
or U9070 (N_9070,N_8828,N_8916);
and U9071 (N_9071,N_8863,N_8892);
nor U9072 (N_9072,N_8845,N_8919);
nand U9073 (N_9073,N_8910,N_8855);
and U9074 (N_9074,N_8861,N_8979);
nor U9075 (N_9075,N_8958,N_8936);
and U9076 (N_9076,N_8929,N_8895);
nand U9077 (N_9077,N_8824,N_8908);
nand U9078 (N_9078,N_8971,N_8818);
nor U9079 (N_9079,N_8835,N_8996);
nor U9080 (N_9080,N_8868,N_8857);
nor U9081 (N_9081,N_8853,N_8915);
or U9082 (N_9082,N_8812,N_8810);
or U9083 (N_9083,N_8880,N_8909);
nand U9084 (N_9084,N_8854,N_8961);
and U9085 (N_9085,N_8918,N_8934);
nor U9086 (N_9086,N_8869,N_8885);
xnor U9087 (N_9087,N_8914,N_8819);
or U9088 (N_9088,N_8945,N_8815);
or U9089 (N_9089,N_8907,N_8836);
nor U9090 (N_9090,N_8982,N_8804);
or U9091 (N_9091,N_8997,N_8832);
and U9092 (N_9092,N_8894,N_8888);
nand U9093 (N_9093,N_8897,N_8955);
or U9094 (N_9094,N_8801,N_8879);
nand U9095 (N_9095,N_8968,N_8843);
nand U9096 (N_9096,N_8959,N_8849);
nor U9097 (N_9097,N_8993,N_8970);
nor U9098 (N_9098,N_8906,N_8881);
xnor U9099 (N_9099,N_8960,N_8980);
or U9100 (N_9100,N_8821,N_8889);
and U9101 (N_9101,N_8966,N_8852);
xor U9102 (N_9102,N_8832,N_8926);
xnor U9103 (N_9103,N_8802,N_8893);
or U9104 (N_9104,N_8840,N_8886);
nand U9105 (N_9105,N_8966,N_8867);
nor U9106 (N_9106,N_8903,N_8887);
nand U9107 (N_9107,N_8972,N_8822);
and U9108 (N_9108,N_8886,N_8992);
xnor U9109 (N_9109,N_8935,N_8859);
or U9110 (N_9110,N_8900,N_8908);
nor U9111 (N_9111,N_8942,N_8981);
or U9112 (N_9112,N_8840,N_8908);
or U9113 (N_9113,N_8905,N_8832);
and U9114 (N_9114,N_8853,N_8838);
nor U9115 (N_9115,N_8850,N_8891);
or U9116 (N_9116,N_8843,N_8894);
nor U9117 (N_9117,N_8956,N_8836);
and U9118 (N_9118,N_8870,N_8910);
nand U9119 (N_9119,N_8868,N_8930);
xnor U9120 (N_9120,N_8998,N_8831);
nor U9121 (N_9121,N_8904,N_8800);
nand U9122 (N_9122,N_8895,N_8830);
nor U9123 (N_9123,N_8891,N_8849);
xor U9124 (N_9124,N_8803,N_8866);
or U9125 (N_9125,N_8890,N_8824);
nand U9126 (N_9126,N_8987,N_8863);
or U9127 (N_9127,N_8919,N_8950);
nand U9128 (N_9128,N_8968,N_8821);
nand U9129 (N_9129,N_8866,N_8818);
xor U9130 (N_9130,N_8802,N_8860);
or U9131 (N_9131,N_8842,N_8954);
xor U9132 (N_9132,N_8842,N_8828);
nor U9133 (N_9133,N_8877,N_8821);
nor U9134 (N_9134,N_8992,N_8802);
nand U9135 (N_9135,N_8978,N_8953);
xnor U9136 (N_9136,N_8883,N_8896);
and U9137 (N_9137,N_8845,N_8954);
and U9138 (N_9138,N_8801,N_8932);
nor U9139 (N_9139,N_8858,N_8861);
nor U9140 (N_9140,N_8808,N_8979);
or U9141 (N_9141,N_8984,N_8918);
and U9142 (N_9142,N_8873,N_8826);
nor U9143 (N_9143,N_8902,N_8900);
nand U9144 (N_9144,N_8890,N_8878);
and U9145 (N_9145,N_8971,N_8928);
or U9146 (N_9146,N_8829,N_8924);
xnor U9147 (N_9147,N_8881,N_8972);
nand U9148 (N_9148,N_8972,N_8885);
or U9149 (N_9149,N_8858,N_8972);
and U9150 (N_9150,N_8998,N_8877);
or U9151 (N_9151,N_8824,N_8969);
xnor U9152 (N_9152,N_8880,N_8832);
and U9153 (N_9153,N_8887,N_8821);
nor U9154 (N_9154,N_8961,N_8879);
nand U9155 (N_9155,N_8978,N_8984);
nor U9156 (N_9156,N_8913,N_8922);
nor U9157 (N_9157,N_8955,N_8916);
xor U9158 (N_9158,N_8825,N_8857);
or U9159 (N_9159,N_8891,N_8856);
or U9160 (N_9160,N_8979,N_8932);
xor U9161 (N_9161,N_8820,N_8964);
nand U9162 (N_9162,N_8857,N_8833);
nand U9163 (N_9163,N_8826,N_8878);
nand U9164 (N_9164,N_8838,N_8962);
nor U9165 (N_9165,N_8901,N_8877);
or U9166 (N_9166,N_8959,N_8800);
and U9167 (N_9167,N_8890,N_8863);
xnor U9168 (N_9168,N_8937,N_8841);
nand U9169 (N_9169,N_8810,N_8833);
and U9170 (N_9170,N_8965,N_8804);
nor U9171 (N_9171,N_8984,N_8902);
nand U9172 (N_9172,N_8944,N_8988);
nand U9173 (N_9173,N_8894,N_8893);
or U9174 (N_9174,N_8920,N_8899);
or U9175 (N_9175,N_8900,N_8977);
xnor U9176 (N_9176,N_8896,N_8975);
xnor U9177 (N_9177,N_8840,N_8802);
or U9178 (N_9178,N_8808,N_8944);
nand U9179 (N_9179,N_8845,N_8832);
nor U9180 (N_9180,N_8939,N_8985);
and U9181 (N_9181,N_8920,N_8892);
or U9182 (N_9182,N_8928,N_8815);
and U9183 (N_9183,N_8856,N_8872);
or U9184 (N_9184,N_8980,N_8870);
and U9185 (N_9185,N_8937,N_8956);
xor U9186 (N_9186,N_8976,N_8917);
xor U9187 (N_9187,N_8909,N_8953);
xnor U9188 (N_9188,N_8994,N_8815);
nand U9189 (N_9189,N_8859,N_8827);
and U9190 (N_9190,N_8857,N_8806);
nor U9191 (N_9191,N_8984,N_8840);
xnor U9192 (N_9192,N_8876,N_8889);
and U9193 (N_9193,N_8890,N_8983);
and U9194 (N_9194,N_8855,N_8918);
xnor U9195 (N_9195,N_8967,N_8866);
nand U9196 (N_9196,N_8959,N_8928);
or U9197 (N_9197,N_8865,N_8849);
or U9198 (N_9198,N_8911,N_8950);
or U9199 (N_9199,N_8900,N_8884);
or U9200 (N_9200,N_9071,N_9157);
xnor U9201 (N_9201,N_9127,N_9097);
nor U9202 (N_9202,N_9054,N_9155);
xor U9203 (N_9203,N_9088,N_9138);
nor U9204 (N_9204,N_9099,N_9137);
and U9205 (N_9205,N_9096,N_9171);
nor U9206 (N_9206,N_9024,N_9156);
xor U9207 (N_9207,N_9049,N_9067);
xor U9208 (N_9208,N_9149,N_9189);
xor U9209 (N_9209,N_9101,N_9178);
or U9210 (N_9210,N_9044,N_9022);
or U9211 (N_9211,N_9004,N_9046);
nor U9212 (N_9212,N_9115,N_9095);
nor U9213 (N_9213,N_9185,N_9016);
and U9214 (N_9214,N_9057,N_9082);
xor U9215 (N_9215,N_9053,N_9043);
nand U9216 (N_9216,N_9158,N_9011);
xor U9217 (N_9217,N_9060,N_9111);
or U9218 (N_9218,N_9094,N_9102);
xnor U9219 (N_9219,N_9031,N_9196);
xor U9220 (N_9220,N_9062,N_9110);
nand U9221 (N_9221,N_9114,N_9175);
nand U9222 (N_9222,N_9197,N_9128);
or U9223 (N_9223,N_9194,N_9187);
xor U9224 (N_9224,N_9083,N_9012);
xor U9225 (N_9225,N_9008,N_9131);
or U9226 (N_9226,N_9077,N_9005);
and U9227 (N_9227,N_9001,N_9075);
xnor U9228 (N_9228,N_9091,N_9190);
nand U9229 (N_9229,N_9032,N_9074);
or U9230 (N_9230,N_9122,N_9010);
and U9231 (N_9231,N_9141,N_9058);
and U9232 (N_9232,N_9145,N_9052);
and U9233 (N_9233,N_9180,N_9025);
and U9234 (N_9234,N_9160,N_9023);
or U9235 (N_9235,N_9000,N_9090);
nand U9236 (N_9236,N_9105,N_9027);
nor U9237 (N_9237,N_9120,N_9084);
and U9238 (N_9238,N_9037,N_9170);
xor U9239 (N_9239,N_9124,N_9143);
and U9240 (N_9240,N_9148,N_9006);
and U9241 (N_9241,N_9162,N_9179);
or U9242 (N_9242,N_9125,N_9161);
nor U9243 (N_9243,N_9177,N_9165);
nand U9244 (N_9244,N_9139,N_9045);
nor U9245 (N_9245,N_9080,N_9159);
and U9246 (N_9246,N_9142,N_9051);
nor U9247 (N_9247,N_9106,N_9002);
xnor U9248 (N_9248,N_9119,N_9059);
nor U9249 (N_9249,N_9117,N_9041);
or U9250 (N_9250,N_9042,N_9078);
and U9251 (N_9251,N_9169,N_9068);
nor U9252 (N_9252,N_9166,N_9144);
nor U9253 (N_9253,N_9035,N_9118);
nor U9254 (N_9254,N_9168,N_9065);
or U9255 (N_9255,N_9086,N_9007);
and U9256 (N_9256,N_9040,N_9019);
nor U9257 (N_9257,N_9018,N_9164);
xnor U9258 (N_9258,N_9134,N_9104);
nand U9259 (N_9259,N_9017,N_9063);
and U9260 (N_9260,N_9199,N_9009);
nor U9261 (N_9261,N_9123,N_9072);
or U9262 (N_9262,N_9050,N_9092);
xor U9263 (N_9263,N_9147,N_9135);
or U9264 (N_9264,N_9021,N_9188);
xnor U9265 (N_9265,N_9061,N_9140);
xor U9266 (N_9266,N_9081,N_9153);
nor U9267 (N_9267,N_9013,N_9100);
nand U9268 (N_9268,N_9056,N_9047);
and U9269 (N_9269,N_9015,N_9033);
or U9270 (N_9270,N_9183,N_9181);
nor U9271 (N_9271,N_9113,N_9003);
nand U9272 (N_9272,N_9030,N_9020);
nor U9273 (N_9273,N_9186,N_9191);
and U9274 (N_9274,N_9126,N_9163);
nand U9275 (N_9275,N_9089,N_9055);
nand U9276 (N_9276,N_9026,N_9048);
xor U9277 (N_9277,N_9014,N_9085);
xnor U9278 (N_9278,N_9079,N_9193);
nand U9279 (N_9279,N_9073,N_9192);
nand U9280 (N_9280,N_9146,N_9184);
xor U9281 (N_9281,N_9098,N_9093);
nand U9282 (N_9282,N_9076,N_9174);
xor U9283 (N_9283,N_9130,N_9112);
and U9284 (N_9284,N_9132,N_9172);
and U9285 (N_9285,N_9038,N_9121);
nor U9286 (N_9286,N_9167,N_9039);
nand U9287 (N_9287,N_9066,N_9103);
nand U9288 (N_9288,N_9109,N_9133);
and U9289 (N_9289,N_9195,N_9108);
nor U9290 (N_9290,N_9036,N_9150);
and U9291 (N_9291,N_9154,N_9116);
nand U9292 (N_9292,N_9152,N_9176);
or U9293 (N_9293,N_9064,N_9173);
and U9294 (N_9294,N_9034,N_9070);
xor U9295 (N_9295,N_9029,N_9028);
or U9296 (N_9296,N_9198,N_9069);
nor U9297 (N_9297,N_9136,N_9129);
and U9298 (N_9298,N_9182,N_9151);
xor U9299 (N_9299,N_9107,N_9087);
xnor U9300 (N_9300,N_9078,N_9020);
xor U9301 (N_9301,N_9019,N_9171);
nor U9302 (N_9302,N_9189,N_9046);
xor U9303 (N_9303,N_9022,N_9100);
and U9304 (N_9304,N_9125,N_9156);
nand U9305 (N_9305,N_9184,N_9083);
and U9306 (N_9306,N_9175,N_9072);
or U9307 (N_9307,N_9164,N_9012);
or U9308 (N_9308,N_9139,N_9007);
nand U9309 (N_9309,N_9003,N_9114);
nor U9310 (N_9310,N_9156,N_9048);
and U9311 (N_9311,N_9069,N_9084);
nand U9312 (N_9312,N_9007,N_9107);
nand U9313 (N_9313,N_9164,N_9075);
and U9314 (N_9314,N_9030,N_9139);
nand U9315 (N_9315,N_9030,N_9131);
xnor U9316 (N_9316,N_9073,N_9043);
and U9317 (N_9317,N_9057,N_9081);
nand U9318 (N_9318,N_9023,N_9161);
nand U9319 (N_9319,N_9098,N_9002);
xnor U9320 (N_9320,N_9043,N_9183);
xnor U9321 (N_9321,N_9169,N_9152);
or U9322 (N_9322,N_9198,N_9087);
xor U9323 (N_9323,N_9144,N_9075);
nand U9324 (N_9324,N_9119,N_9011);
nand U9325 (N_9325,N_9157,N_9125);
or U9326 (N_9326,N_9068,N_9170);
and U9327 (N_9327,N_9164,N_9024);
nand U9328 (N_9328,N_9195,N_9030);
and U9329 (N_9329,N_9141,N_9006);
or U9330 (N_9330,N_9051,N_9020);
xnor U9331 (N_9331,N_9195,N_9068);
and U9332 (N_9332,N_9088,N_9067);
and U9333 (N_9333,N_9047,N_9082);
xor U9334 (N_9334,N_9013,N_9044);
and U9335 (N_9335,N_9009,N_9197);
or U9336 (N_9336,N_9107,N_9065);
and U9337 (N_9337,N_9071,N_9143);
and U9338 (N_9338,N_9010,N_9092);
nor U9339 (N_9339,N_9034,N_9133);
nand U9340 (N_9340,N_9086,N_9025);
and U9341 (N_9341,N_9102,N_9154);
and U9342 (N_9342,N_9015,N_9072);
nand U9343 (N_9343,N_9138,N_9152);
nand U9344 (N_9344,N_9174,N_9079);
nor U9345 (N_9345,N_9085,N_9030);
nor U9346 (N_9346,N_9010,N_9197);
and U9347 (N_9347,N_9028,N_9047);
nor U9348 (N_9348,N_9144,N_9134);
or U9349 (N_9349,N_9181,N_9056);
nor U9350 (N_9350,N_9010,N_9168);
or U9351 (N_9351,N_9135,N_9050);
or U9352 (N_9352,N_9113,N_9171);
nor U9353 (N_9353,N_9113,N_9119);
nor U9354 (N_9354,N_9008,N_9040);
or U9355 (N_9355,N_9075,N_9047);
and U9356 (N_9356,N_9086,N_9044);
nand U9357 (N_9357,N_9109,N_9088);
nor U9358 (N_9358,N_9157,N_9160);
and U9359 (N_9359,N_9134,N_9083);
xnor U9360 (N_9360,N_9138,N_9151);
or U9361 (N_9361,N_9149,N_9070);
nor U9362 (N_9362,N_9177,N_9132);
xnor U9363 (N_9363,N_9044,N_9101);
and U9364 (N_9364,N_9082,N_9016);
nor U9365 (N_9365,N_9118,N_9191);
and U9366 (N_9366,N_9073,N_9113);
nor U9367 (N_9367,N_9149,N_9009);
nand U9368 (N_9368,N_9123,N_9065);
or U9369 (N_9369,N_9079,N_9084);
nor U9370 (N_9370,N_9159,N_9061);
and U9371 (N_9371,N_9116,N_9198);
xor U9372 (N_9372,N_9119,N_9057);
nor U9373 (N_9373,N_9103,N_9162);
and U9374 (N_9374,N_9007,N_9122);
or U9375 (N_9375,N_9178,N_9088);
and U9376 (N_9376,N_9115,N_9079);
nor U9377 (N_9377,N_9062,N_9028);
and U9378 (N_9378,N_9111,N_9179);
and U9379 (N_9379,N_9078,N_9116);
nand U9380 (N_9380,N_9163,N_9165);
nor U9381 (N_9381,N_9108,N_9092);
nand U9382 (N_9382,N_9113,N_9158);
or U9383 (N_9383,N_9197,N_9063);
and U9384 (N_9384,N_9188,N_9138);
nor U9385 (N_9385,N_9086,N_9019);
nand U9386 (N_9386,N_9188,N_9051);
nor U9387 (N_9387,N_9057,N_9157);
xor U9388 (N_9388,N_9183,N_9190);
and U9389 (N_9389,N_9134,N_9061);
xor U9390 (N_9390,N_9187,N_9141);
nand U9391 (N_9391,N_9129,N_9059);
xor U9392 (N_9392,N_9009,N_9127);
and U9393 (N_9393,N_9131,N_9043);
or U9394 (N_9394,N_9038,N_9035);
or U9395 (N_9395,N_9118,N_9023);
and U9396 (N_9396,N_9155,N_9061);
or U9397 (N_9397,N_9106,N_9063);
or U9398 (N_9398,N_9030,N_9174);
or U9399 (N_9399,N_9102,N_9178);
and U9400 (N_9400,N_9246,N_9392);
or U9401 (N_9401,N_9357,N_9264);
nor U9402 (N_9402,N_9303,N_9225);
or U9403 (N_9403,N_9239,N_9292);
nor U9404 (N_9404,N_9272,N_9300);
or U9405 (N_9405,N_9384,N_9273);
nand U9406 (N_9406,N_9242,N_9332);
nand U9407 (N_9407,N_9388,N_9323);
nor U9408 (N_9408,N_9285,N_9205);
or U9409 (N_9409,N_9256,N_9330);
or U9410 (N_9410,N_9371,N_9209);
nand U9411 (N_9411,N_9350,N_9354);
or U9412 (N_9412,N_9207,N_9312);
and U9413 (N_9413,N_9348,N_9270);
and U9414 (N_9414,N_9324,N_9274);
or U9415 (N_9415,N_9344,N_9253);
xor U9416 (N_9416,N_9373,N_9391);
and U9417 (N_9417,N_9289,N_9299);
and U9418 (N_9418,N_9311,N_9314);
xnor U9419 (N_9419,N_9240,N_9369);
nand U9420 (N_9420,N_9355,N_9293);
or U9421 (N_9421,N_9263,N_9291);
xor U9422 (N_9422,N_9201,N_9203);
nand U9423 (N_9423,N_9275,N_9220);
nor U9424 (N_9424,N_9361,N_9372);
xor U9425 (N_9425,N_9243,N_9356);
and U9426 (N_9426,N_9305,N_9290);
nand U9427 (N_9427,N_9342,N_9304);
and U9428 (N_9428,N_9394,N_9386);
or U9429 (N_9429,N_9395,N_9206);
or U9430 (N_9430,N_9266,N_9267);
xor U9431 (N_9431,N_9250,N_9238);
nor U9432 (N_9432,N_9310,N_9252);
or U9433 (N_9433,N_9212,N_9251);
nor U9434 (N_9434,N_9258,N_9297);
and U9435 (N_9435,N_9200,N_9296);
nor U9436 (N_9436,N_9337,N_9309);
nand U9437 (N_9437,N_9226,N_9237);
nor U9438 (N_9438,N_9399,N_9277);
nand U9439 (N_9439,N_9318,N_9248);
xnor U9440 (N_9440,N_9364,N_9224);
xor U9441 (N_9441,N_9280,N_9294);
or U9442 (N_9442,N_9281,N_9331);
nand U9443 (N_9443,N_9218,N_9315);
nor U9444 (N_9444,N_9368,N_9276);
and U9445 (N_9445,N_9231,N_9327);
xnor U9446 (N_9446,N_9317,N_9223);
xor U9447 (N_9447,N_9329,N_9319);
and U9448 (N_9448,N_9236,N_9255);
nor U9449 (N_9449,N_9396,N_9346);
nor U9450 (N_9450,N_9343,N_9325);
or U9451 (N_9451,N_9326,N_9335);
xnor U9452 (N_9452,N_9385,N_9262);
nand U9453 (N_9453,N_9283,N_9393);
or U9454 (N_9454,N_9316,N_9397);
xnor U9455 (N_9455,N_9338,N_9378);
and U9456 (N_9456,N_9322,N_9282);
or U9457 (N_9457,N_9221,N_9377);
nor U9458 (N_9458,N_9241,N_9210);
nor U9459 (N_9459,N_9284,N_9298);
and U9460 (N_9460,N_9216,N_9219);
xor U9461 (N_9461,N_9366,N_9244);
xor U9462 (N_9462,N_9261,N_9375);
and U9463 (N_9463,N_9271,N_9227);
nand U9464 (N_9464,N_9213,N_9370);
xnor U9465 (N_9465,N_9363,N_9279);
xnor U9466 (N_9466,N_9353,N_9382);
nand U9467 (N_9467,N_9376,N_9398);
nand U9468 (N_9468,N_9230,N_9257);
nor U9469 (N_9469,N_9383,N_9245);
and U9470 (N_9470,N_9217,N_9387);
nand U9471 (N_9471,N_9345,N_9208);
xnor U9472 (N_9472,N_9259,N_9268);
nand U9473 (N_9473,N_9341,N_9249);
nand U9474 (N_9474,N_9214,N_9222);
and U9475 (N_9475,N_9352,N_9358);
and U9476 (N_9476,N_9389,N_9215);
or U9477 (N_9477,N_9265,N_9288);
nand U9478 (N_9478,N_9381,N_9295);
xor U9479 (N_9479,N_9328,N_9320);
and U9480 (N_9480,N_9286,N_9302);
and U9481 (N_9481,N_9362,N_9321);
xnor U9482 (N_9482,N_9367,N_9202);
and U9483 (N_9483,N_9339,N_9269);
nand U9484 (N_9484,N_9260,N_9204);
xor U9485 (N_9485,N_9360,N_9234);
and U9486 (N_9486,N_9235,N_9359);
nor U9487 (N_9487,N_9351,N_9254);
and U9488 (N_9488,N_9301,N_9306);
nand U9489 (N_9489,N_9308,N_9336);
and U9490 (N_9490,N_9340,N_9374);
nand U9491 (N_9491,N_9228,N_9333);
nand U9492 (N_9492,N_9232,N_9307);
and U9493 (N_9493,N_9347,N_9379);
xor U9494 (N_9494,N_9229,N_9233);
nor U9495 (N_9495,N_9334,N_9380);
or U9496 (N_9496,N_9247,N_9365);
nor U9497 (N_9497,N_9211,N_9349);
or U9498 (N_9498,N_9390,N_9278);
nor U9499 (N_9499,N_9287,N_9313);
xor U9500 (N_9500,N_9295,N_9201);
and U9501 (N_9501,N_9256,N_9262);
nor U9502 (N_9502,N_9297,N_9309);
xnor U9503 (N_9503,N_9272,N_9233);
nand U9504 (N_9504,N_9223,N_9260);
nor U9505 (N_9505,N_9254,N_9302);
or U9506 (N_9506,N_9232,N_9265);
or U9507 (N_9507,N_9200,N_9376);
nor U9508 (N_9508,N_9258,N_9243);
and U9509 (N_9509,N_9380,N_9338);
or U9510 (N_9510,N_9386,N_9217);
nor U9511 (N_9511,N_9362,N_9253);
xnor U9512 (N_9512,N_9389,N_9265);
nor U9513 (N_9513,N_9216,N_9363);
or U9514 (N_9514,N_9330,N_9265);
nand U9515 (N_9515,N_9342,N_9348);
or U9516 (N_9516,N_9299,N_9263);
or U9517 (N_9517,N_9330,N_9360);
nor U9518 (N_9518,N_9312,N_9333);
nor U9519 (N_9519,N_9313,N_9257);
nor U9520 (N_9520,N_9289,N_9380);
and U9521 (N_9521,N_9341,N_9269);
and U9522 (N_9522,N_9317,N_9206);
nor U9523 (N_9523,N_9257,N_9335);
xnor U9524 (N_9524,N_9397,N_9373);
xor U9525 (N_9525,N_9339,N_9377);
nor U9526 (N_9526,N_9272,N_9231);
and U9527 (N_9527,N_9245,N_9314);
xnor U9528 (N_9528,N_9356,N_9388);
or U9529 (N_9529,N_9275,N_9204);
nor U9530 (N_9530,N_9285,N_9213);
nor U9531 (N_9531,N_9342,N_9299);
or U9532 (N_9532,N_9260,N_9384);
nand U9533 (N_9533,N_9216,N_9212);
xor U9534 (N_9534,N_9271,N_9333);
and U9535 (N_9535,N_9333,N_9269);
or U9536 (N_9536,N_9361,N_9351);
nor U9537 (N_9537,N_9267,N_9217);
nor U9538 (N_9538,N_9240,N_9216);
and U9539 (N_9539,N_9207,N_9267);
xor U9540 (N_9540,N_9202,N_9331);
xnor U9541 (N_9541,N_9302,N_9210);
nor U9542 (N_9542,N_9291,N_9395);
nor U9543 (N_9543,N_9362,N_9271);
xnor U9544 (N_9544,N_9383,N_9377);
nand U9545 (N_9545,N_9301,N_9290);
or U9546 (N_9546,N_9332,N_9239);
nand U9547 (N_9547,N_9393,N_9397);
nand U9548 (N_9548,N_9332,N_9201);
nor U9549 (N_9549,N_9243,N_9304);
nand U9550 (N_9550,N_9361,N_9259);
nand U9551 (N_9551,N_9318,N_9346);
or U9552 (N_9552,N_9337,N_9274);
xor U9553 (N_9553,N_9238,N_9316);
and U9554 (N_9554,N_9373,N_9308);
xor U9555 (N_9555,N_9301,N_9324);
xnor U9556 (N_9556,N_9299,N_9284);
and U9557 (N_9557,N_9229,N_9266);
nor U9558 (N_9558,N_9389,N_9253);
xnor U9559 (N_9559,N_9282,N_9234);
nor U9560 (N_9560,N_9239,N_9267);
nand U9561 (N_9561,N_9318,N_9322);
nor U9562 (N_9562,N_9232,N_9231);
and U9563 (N_9563,N_9256,N_9394);
xor U9564 (N_9564,N_9325,N_9396);
nor U9565 (N_9565,N_9224,N_9221);
or U9566 (N_9566,N_9345,N_9232);
xnor U9567 (N_9567,N_9321,N_9393);
and U9568 (N_9568,N_9376,N_9292);
nand U9569 (N_9569,N_9317,N_9344);
and U9570 (N_9570,N_9289,N_9300);
nand U9571 (N_9571,N_9389,N_9234);
nor U9572 (N_9572,N_9259,N_9200);
or U9573 (N_9573,N_9217,N_9201);
xnor U9574 (N_9574,N_9374,N_9368);
or U9575 (N_9575,N_9287,N_9200);
or U9576 (N_9576,N_9369,N_9392);
nand U9577 (N_9577,N_9219,N_9369);
nor U9578 (N_9578,N_9255,N_9312);
xnor U9579 (N_9579,N_9360,N_9210);
nand U9580 (N_9580,N_9235,N_9215);
nor U9581 (N_9581,N_9380,N_9240);
xnor U9582 (N_9582,N_9273,N_9298);
and U9583 (N_9583,N_9383,N_9338);
nand U9584 (N_9584,N_9351,N_9233);
nor U9585 (N_9585,N_9356,N_9327);
nand U9586 (N_9586,N_9372,N_9207);
nor U9587 (N_9587,N_9318,N_9274);
or U9588 (N_9588,N_9390,N_9257);
or U9589 (N_9589,N_9329,N_9223);
xor U9590 (N_9590,N_9283,N_9391);
nor U9591 (N_9591,N_9388,N_9358);
xor U9592 (N_9592,N_9227,N_9379);
or U9593 (N_9593,N_9244,N_9311);
nand U9594 (N_9594,N_9360,N_9277);
or U9595 (N_9595,N_9215,N_9298);
or U9596 (N_9596,N_9392,N_9298);
xnor U9597 (N_9597,N_9200,N_9251);
nand U9598 (N_9598,N_9201,N_9244);
or U9599 (N_9599,N_9230,N_9263);
xnor U9600 (N_9600,N_9473,N_9537);
or U9601 (N_9601,N_9587,N_9573);
and U9602 (N_9602,N_9533,N_9504);
nand U9603 (N_9603,N_9556,N_9497);
xnor U9604 (N_9604,N_9570,N_9430);
or U9605 (N_9605,N_9443,N_9559);
nor U9606 (N_9606,N_9571,N_9458);
and U9607 (N_9607,N_9514,N_9583);
nand U9608 (N_9608,N_9547,N_9588);
and U9609 (N_9609,N_9419,N_9402);
xnor U9610 (N_9610,N_9555,N_9597);
and U9611 (N_9611,N_9535,N_9410);
nand U9612 (N_9612,N_9499,N_9464);
and U9613 (N_9613,N_9538,N_9505);
and U9614 (N_9614,N_9474,N_9426);
xnor U9615 (N_9615,N_9479,N_9433);
xnor U9616 (N_9616,N_9534,N_9503);
and U9617 (N_9617,N_9407,N_9574);
nor U9618 (N_9618,N_9432,N_9521);
nand U9619 (N_9619,N_9586,N_9592);
or U9620 (N_9620,N_9526,N_9468);
nand U9621 (N_9621,N_9506,N_9436);
nand U9622 (N_9622,N_9549,N_9424);
or U9623 (N_9623,N_9470,N_9589);
xor U9624 (N_9624,N_9524,N_9528);
nand U9625 (N_9625,N_9580,N_9544);
nor U9626 (N_9626,N_9400,N_9498);
xor U9627 (N_9627,N_9539,N_9598);
nor U9628 (N_9628,N_9440,N_9569);
and U9629 (N_9629,N_9448,N_9512);
nand U9630 (N_9630,N_9445,N_9449);
nand U9631 (N_9631,N_9591,N_9435);
xor U9632 (N_9632,N_9425,N_9532);
or U9633 (N_9633,N_9416,N_9527);
xnor U9634 (N_9634,N_9542,N_9455);
and U9635 (N_9635,N_9554,N_9561);
or U9636 (N_9636,N_9579,N_9406);
xor U9637 (N_9637,N_9447,N_9516);
or U9638 (N_9638,N_9452,N_9484);
nand U9639 (N_9639,N_9441,N_9476);
and U9640 (N_9640,N_9593,N_9545);
nand U9641 (N_9641,N_9558,N_9482);
and U9642 (N_9642,N_9596,N_9490);
nor U9643 (N_9643,N_9404,N_9408);
and U9644 (N_9644,N_9475,N_9466);
and U9645 (N_9645,N_9502,N_9472);
nor U9646 (N_9646,N_9576,N_9460);
or U9647 (N_9647,N_9531,N_9478);
xnor U9648 (N_9648,N_9513,N_9439);
nand U9649 (N_9649,N_9566,N_9456);
or U9650 (N_9650,N_9438,N_9518);
nand U9651 (N_9651,N_9469,N_9507);
xnor U9652 (N_9652,N_9462,N_9415);
xnor U9653 (N_9653,N_9463,N_9429);
and U9654 (N_9654,N_9495,N_9409);
nor U9655 (N_9655,N_9412,N_9483);
or U9656 (N_9656,N_9508,N_9481);
nor U9657 (N_9657,N_9488,N_9584);
nor U9658 (N_9658,N_9428,N_9489);
nor U9659 (N_9659,N_9465,N_9572);
and U9660 (N_9660,N_9492,N_9459);
or U9661 (N_9661,N_9509,N_9578);
nor U9662 (N_9662,N_9562,N_9461);
or U9663 (N_9663,N_9560,N_9525);
and U9664 (N_9664,N_9413,N_9567);
or U9665 (N_9665,N_9437,N_9417);
nor U9666 (N_9666,N_9444,N_9557);
nor U9667 (N_9667,N_9471,N_9511);
nand U9668 (N_9668,N_9427,N_9553);
and U9669 (N_9669,N_9403,N_9450);
xor U9670 (N_9670,N_9519,N_9480);
nor U9671 (N_9671,N_9563,N_9446);
nand U9672 (N_9672,N_9453,N_9405);
and U9673 (N_9673,N_9494,N_9487);
or U9674 (N_9674,N_9575,N_9510);
and U9675 (N_9675,N_9540,N_9454);
or U9676 (N_9676,N_9414,N_9420);
or U9677 (N_9677,N_9551,N_9529);
nor U9678 (N_9678,N_9530,N_9568);
or U9679 (N_9679,N_9421,N_9590);
or U9680 (N_9680,N_9451,N_9564);
xor U9681 (N_9681,N_9565,N_9501);
nand U9682 (N_9682,N_9418,N_9517);
xnor U9683 (N_9683,N_9577,N_9582);
xor U9684 (N_9684,N_9550,N_9422);
or U9685 (N_9685,N_9541,N_9401);
and U9686 (N_9686,N_9491,N_9585);
and U9687 (N_9687,N_9520,N_9496);
nand U9688 (N_9688,N_9515,N_9467);
and U9689 (N_9689,N_9594,N_9423);
or U9690 (N_9690,N_9411,N_9522);
nor U9691 (N_9691,N_9486,N_9442);
and U9692 (N_9692,N_9523,N_9581);
and U9693 (N_9693,N_9493,N_9434);
nand U9694 (N_9694,N_9548,N_9543);
and U9695 (N_9695,N_9552,N_9431);
nand U9696 (N_9696,N_9485,N_9500);
or U9697 (N_9697,N_9477,N_9536);
or U9698 (N_9698,N_9546,N_9457);
nor U9699 (N_9699,N_9599,N_9595);
and U9700 (N_9700,N_9569,N_9438);
nor U9701 (N_9701,N_9579,N_9445);
or U9702 (N_9702,N_9422,N_9466);
and U9703 (N_9703,N_9484,N_9508);
or U9704 (N_9704,N_9426,N_9573);
xor U9705 (N_9705,N_9552,N_9500);
nand U9706 (N_9706,N_9431,N_9566);
and U9707 (N_9707,N_9569,N_9410);
xnor U9708 (N_9708,N_9509,N_9536);
nor U9709 (N_9709,N_9573,N_9419);
nand U9710 (N_9710,N_9407,N_9539);
or U9711 (N_9711,N_9430,N_9598);
and U9712 (N_9712,N_9553,N_9491);
nor U9713 (N_9713,N_9498,N_9439);
nand U9714 (N_9714,N_9587,N_9540);
or U9715 (N_9715,N_9446,N_9576);
xnor U9716 (N_9716,N_9418,N_9448);
and U9717 (N_9717,N_9479,N_9426);
or U9718 (N_9718,N_9489,N_9443);
and U9719 (N_9719,N_9426,N_9584);
xor U9720 (N_9720,N_9498,N_9418);
nor U9721 (N_9721,N_9589,N_9592);
or U9722 (N_9722,N_9570,N_9499);
or U9723 (N_9723,N_9514,N_9532);
or U9724 (N_9724,N_9557,N_9570);
nor U9725 (N_9725,N_9472,N_9560);
nand U9726 (N_9726,N_9444,N_9513);
and U9727 (N_9727,N_9580,N_9508);
xnor U9728 (N_9728,N_9545,N_9448);
xnor U9729 (N_9729,N_9566,N_9549);
nand U9730 (N_9730,N_9567,N_9469);
nor U9731 (N_9731,N_9531,N_9485);
nand U9732 (N_9732,N_9580,N_9556);
xor U9733 (N_9733,N_9516,N_9460);
nand U9734 (N_9734,N_9574,N_9482);
nor U9735 (N_9735,N_9572,N_9420);
and U9736 (N_9736,N_9569,N_9562);
and U9737 (N_9737,N_9550,N_9542);
and U9738 (N_9738,N_9597,N_9544);
nor U9739 (N_9739,N_9565,N_9463);
xnor U9740 (N_9740,N_9443,N_9492);
and U9741 (N_9741,N_9538,N_9463);
and U9742 (N_9742,N_9585,N_9588);
xnor U9743 (N_9743,N_9555,N_9493);
and U9744 (N_9744,N_9431,N_9435);
xnor U9745 (N_9745,N_9579,N_9546);
or U9746 (N_9746,N_9559,N_9406);
nor U9747 (N_9747,N_9505,N_9418);
nand U9748 (N_9748,N_9511,N_9556);
or U9749 (N_9749,N_9510,N_9422);
and U9750 (N_9750,N_9414,N_9543);
and U9751 (N_9751,N_9580,N_9539);
nand U9752 (N_9752,N_9582,N_9516);
or U9753 (N_9753,N_9568,N_9582);
nand U9754 (N_9754,N_9420,N_9415);
nand U9755 (N_9755,N_9539,N_9487);
xor U9756 (N_9756,N_9553,N_9465);
and U9757 (N_9757,N_9411,N_9440);
nor U9758 (N_9758,N_9542,N_9536);
xnor U9759 (N_9759,N_9517,N_9569);
or U9760 (N_9760,N_9414,N_9547);
or U9761 (N_9761,N_9471,N_9488);
nand U9762 (N_9762,N_9520,N_9522);
xnor U9763 (N_9763,N_9495,N_9469);
nand U9764 (N_9764,N_9440,N_9487);
xor U9765 (N_9765,N_9555,N_9479);
nor U9766 (N_9766,N_9418,N_9482);
nand U9767 (N_9767,N_9472,N_9475);
or U9768 (N_9768,N_9579,N_9468);
and U9769 (N_9769,N_9468,N_9488);
nand U9770 (N_9770,N_9451,N_9520);
nand U9771 (N_9771,N_9440,N_9574);
xnor U9772 (N_9772,N_9423,N_9511);
or U9773 (N_9773,N_9481,N_9555);
or U9774 (N_9774,N_9579,N_9570);
and U9775 (N_9775,N_9555,N_9534);
xor U9776 (N_9776,N_9542,N_9426);
nor U9777 (N_9777,N_9448,N_9474);
nand U9778 (N_9778,N_9550,N_9402);
or U9779 (N_9779,N_9528,N_9426);
nand U9780 (N_9780,N_9509,N_9462);
nand U9781 (N_9781,N_9509,N_9442);
nor U9782 (N_9782,N_9479,N_9594);
or U9783 (N_9783,N_9518,N_9426);
xnor U9784 (N_9784,N_9413,N_9495);
and U9785 (N_9785,N_9467,N_9524);
nand U9786 (N_9786,N_9428,N_9435);
xnor U9787 (N_9787,N_9513,N_9583);
and U9788 (N_9788,N_9433,N_9441);
and U9789 (N_9789,N_9589,N_9548);
xor U9790 (N_9790,N_9593,N_9415);
xor U9791 (N_9791,N_9447,N_9512);
nor U9792 (N_9792,N_9552,N_9516);
nand U9793 (N_9793,N_9416,N_9407);
xor U9794 (N_9794,N_9540,N_9438);
or U9795 (N_9795,N_9591,N_9538);
and U9796 (N_9796,N_9405,N_9538);
xnor U9797 (N_9797,N_9435,N_9525);
nand U9798 (N_9798,N_9505,N_9435);
nor U9799 (N_9799,N_9579,N_9453);
nand U9800 (N_9800,N_9617,N_9680);
and U9801 (N_9801,N_9610,N_9775);
and U9802 (N_9802,N_9671,N_9724);
xnor U9803 (N_9803,N_9607,N_9749);
nor U9804 (N_9804,N_9649,N_9664);
nor U9805 (N_9805,N_9628,N_9714);
nand U9806 (N_9806,N_9631,N_9624);
nor U9807 (N_9807,N_9789,N_9707);
or U9808 (N_9808,N_9634,N_9750);
nand U9809 (N_9809,N_9614,N_9659);
nand U9810 (N_9810,N_9708,N_9786);
nand U9811 (N_9811,N_9788,N_9705);
xor U9812 (N_9812,N_9678,N_9622);
nand U9813 (N_9813,N_9609,N_9641);
nor U9814 (N_9814,N_9650,N_9797);
nor U9815 (N_9815,N_9732,N_9720);
nor U9816 (N_9816,N_9602,N_9765);
and U9817 (N_9817,N_9605,N_9644);
nor U9818 (N_9818,N_9780,N_9698);
and U9819 (N_9819,N_9675,N_9681);
nor U9820 (N_9820,N_9632,N_9737);
nand U9821 (N_9821,N_9767,N_9653);
xor U9822 (N_9822,N_9785,N_9621);
nor U9823 (N_9823,N_9696,N_9616);
xnor U9824 (N_9824,N_9738,N_9691);
nand U9825 (N_9825,N_9783,N_9697);
xnor U9826 (N_9826,N_9763,N_9623);
xor U9827 (N_9827,N_9784,N_9612);
and U9828 (N_9828,N_9673,N_9706);
and U9829 (N_9829,N_9682,N_9625);
and U9830 (N_9830,N_9702,N_9741);
nand U9831 (N_9831,N_9677,N_9759);
or U9832 (N_9832,N_9660,N_9626);
nor U9833 (N_9833,N_9751,N_9651);
and U9834 (N_9834,N_9719,N_9726);
or U9835 (N_9835,N_9661,N_9782);
or U9836 (N_9836,N_9725,N_9755);
xor U9837 (N_9837,N_9655,N_9676);
nand U9838 (N_9838,N_9776,N_9796);
xnor U9839 (N_9839,N_9717,N_9711);
xor U9840 (N_9840,N_9633,N_9667);
nand U9841 (N_9841,N_9638,N_9731);
or U9842 (N_9842,N_9730,N_9608);
nor U9843 (N_9843,N_9700,N_9672);
and U9844 (N_9844,N_9722,N_9777);
nand U9845 (N_9845,N_9668,N_9686);
or U9846 (N_9846,N_9637,N_9630);
xnor U9847 (N_9847,N_9728,N_9640);
and U9848 (N_9848,N_9674,N_9629);
nor U9849 (N_9849,N_9643,N_9773);
xnor U9850 (N_9850,N_9721,N_9606);
and U9851 (N_9851,N_9694,N_9736);
nand U9852 (N_9852,N_9735,N_9727);
nor U9853 (N_9853,N_9740,N_9663);
or U9854 (N_9854,N_9739,N_9613);
or U9855 (N_9855,N_9670,N_9747);
xor U9856 (N_9856,N_9710,N_9748);
nor U9857 (N_9857,N_9648,N_9716);
and U9858 (N_9858,N_9761,N_9757);
xor U9859 (N_9859,N_9699,N_9657);
or U9860 (N_9860,N_9787,N_9669);
nand U9861 (N_9861,N_9723,N_9762);
and U9862 (N_9862,N_9742,N_9662);
nand U9863 (N_9863,N_9770,N_9779);
nand U9864 (N_9864,N_9658,N_9611);
nor U9865 (N_9865,N_9704,N_9746);
or U9866 (N_9866,N_9791,N_9756);
or U9867 (N_9867,N_9693,N_9652);
nand U9868 (N_9868,N_9709,N_9745);
or U9869 (N_9869,N_9620,N_9703);
and U9870 (N_9870,N_9689,N_9795);
nor U9871 (N_9871,N_9683,N_9793);
or U9872 (N_9872,N_9618,N_9772);
xor U9873 (N_9873,N_9774,N_9647);
or U9874 (N_9874,N_9642,N_9687);
nor U9875 (N_9875,N_9656,N_9768);
or U9876 (N_9876,N_9713,N_9619);
nand U9877 (N_9877,N_9604,N_9753);
and U9878 (N_9878,N_9627,N_9679);
xnor U9879 (N_9879,N_9712,N_9790);
and U9880 (N_9880,N_9743,N_9635);
and U9881 (N_9881,N_9636,N_9701);
nand U9882 (N_9882,N_9764,N_9733);
or U9883 (N_9883,N_9754,N_9794);
or U9884 (N_9884,N_9665,N_9666);
and U9885 (N_9885,N_9646,N_9734);
or U9886 (N_9886,N_9685,N_9715);
nand U9887 (N_9887,N_9692,N_9781);
or U9888 (N_9888,N_9729,N_9792);
nor U9889 (N_9889,N_9778,N_9718);
or U9890 (N_9890,N_9639,N_9760);
nor U9891 (N_9891,N_9684,N_9600);
nand U9892 (N_9892,N_9654,N_9695);
or U9893 (N_9893,N_9758,N_9769);
xnor U9894 (N_9894,N_9645,N_9690);
xnor U9895 (N_9895,N_9603,N_9744);
nor U9896 (N_9896,N_9799,N_9601);
or U9897 (N_9897,N_9688,N_9798);
nand U9898 (N_9898,N_9752,N_9771);
and U9899 (N_9899,N_9615,N_9766);
nor U9900 (N_9900,N_9740,N_9793);
nand U9901 (N_9901,N_9656,N_9735);
or U9902 (N_9902,N_9767,N_9659);
and U9903 (N_9903,N_9688,N_9762);
or U9904 (N_9904,N_9672,N_9611);
or U9905 (N_9905,N_9704,N_9612);
and U9906 (N_9906,N_9692,N_9796);
nor U9907 (N_9907,N_9725,N_9724);
xor U9908 (N_9908,N_9740,N_9750);
and U9909 (N_9909,N_9680,N_9761);
xnor U9910 (N_9910,N_9742,N_9792);
and U9911 (N_9911,N_9702,N_9603);
nand U9912 (N_9912,N_9718,N_9700);
and U9913 (N_9913,N_9741,N_9647);
nor U9914 (N_9914,N_9728,N_9797);
or U9915 (N_9915,N_9729,N_9702);
or U9916 (N_9916,N_9781,N_9605);
nand U9917 (N_9917,N_9763,N_9690);
xnor U9918 (N_9918,N_9670,N_9600);
nor U9919 (N_9919,N_9605,N_9705);
nor U9920 (N_9920,N_9740,N_9635);
xor U9921 (N_9921,N_9758,N_9736);
and U9922 (N_9922,N_9646,N_9678);
xnor U9923 (N_9923,N_9749,N_9669);
and U9924 (N_9924,N_9684,N_9655);
xnor U9925 (N_9925,N_9794,N_9785);
nand U9926 (N_9926,N_9799,N_9653);
or U9927 (N_9927,N_9796,N_9779);
and U9928 (N_9928,N_9695,N_9639);
nor U9929 (N_9929,N_9613,N_9755);
nand U9930 (N_9930,N_9723,N_9682);
and U9931 (N_9931,N_9717,N_9601);
or U9932 (N_9932,N_9657,N_9652);
nand U9933 (N_9933,N_9675,N_9730);
xor U9934 (N_9934,N_9777,N_9716);
nor U9935 (N_9935,N_9674,N_9615);
and U9936 (N_9936,N_9604,N_9664);
nand U9937 (N_9937,N_9683,N_9604);
nor U9938 (N_9938,N_9638,N_9724);
xnor U9939 (N_9939,N_9629,N_9776);
nor U9940 (N_9940,N_9653,N_9635);
nand U9941 (N_9941,N_9777,N_9742);
and U9942 (N_9942,N_9708,N_9613);
xnor U9943 (N_9943,N_9762,N_9697);
xor U9944 (N_9944,N_9668,N_9670);
xor U9945 (N_9945,N_9748,N_9724);
nand U9946 (N_9946,N_9618,N_9624);
xnor U9947 (N_9947,N_9714,N_9644);
xor U9948 (N_9948,N_9728,N_9740);
xnor U9949 (N_9949,N_9798,N_9684);
nor U9950 (N_9950,N_9627,N_9729);
xor U9951 (N_9951,N_9619,N_9738);
nand U9952 (N_9952,N_9744,N_9798);
and U9953 (N_9953,N_9620,N_9662);
or U9954 (N_9954,N_9750,N_9725);
and U9955 (N_9955,N_9607,N_9628);
or U9956 (N_9956,N_9664,N_9670);
or U9957 (N_9957,N_9745,N_9770);
and U9958 (N_9958,N_9793,N_9606);
xor U9959 (N_9959,N_9703,N_9636);
xnor U9960 (N_9960,N_9656,N_9728);
xnor U9961 (N_9961,N_9614,N_9603);
or U9962 (N_9962,N_9658,N_9649);
xnor U9963 (N_9963,N_9782,N_9790);
nor U9964 (N_9964,N_9787,N_9763);
and U9965 (N_9965,N_9702,N_9639);
nand U9966 (N_9966,N_9636,N_9761);
nor U9967 (N_9967,N_9631,N_9601);
and U9968 (N_9968,N_9673,N_9613);
or U9969 (N_9969,N_9760,N_9782);
xor U9970 (N_9970,N_9697,N_9664);
and U9971 (N_9971,N_9759,N_9776);
nor U9972 (N_9972,N_9785,N_9641);
xor U9973 (N_9973,N_9722,N_9796);
xnor U9974 (N_9974,N_9746,N_9763);
or U9975 (N_9975,N_9609,N_9719);
nand U9976 (N_9976,N_9693,N_9718);
xnor U9977 (N_9977,N_9724,N_9649);
nand U9978 (N_9978,N_9665,N_9624);
and U9979 (N_9979,N_9729,N_9688);
or U9980 (N_9980,N_9736,N_9792);
nand U9981 (N_9981,N_9731,N_9725);
xnor U9982 (N_9982,N_9665,N_9641);
nand U9983 (N_9983,N_9648,N_9609);
xnor U9984 (N_9984,N_9719,N_9750);
nand U9985 (N_9985,N_9767,N_9747);
xnor U9986 (N_9986,N_9641,N_9695);
nor U9987 (N_9987,N_9721,N_9665);
nand U9988 (N_9988,N_9783,N_9735);
nor U9989 (N_9989,N_9776,N_9676);
nor U9990 (N_9990,N_9708,N_9707);
nand U9991 (N_9991,N_9645,N_9743);
xnor U9992 (N_9992,N_9620,N_9785);
xnor U9993 (N_9993,N_9683,N_9767);
or U9994 (N_9994,N_9784,N_9686);
or U9995 (N_9995,N_9617,N_9783);
nand U9996 (N_9996,N_9764,N_9721);
and U9997 (N_9997,N_9776,N_9784);
or U9998 (N_9998,N_9734,N_9605);
nor U9999 (N_9999,N_9707,N_9751);
xnor U10000 (N_10000,N_9937,N_9852);
nor U10001 (N_10001,N_9979,N_9949);
nand U10002 (N_10002,N_9811,N_9954);
and U10003 (N_10003,N_9923,N_9941);
nor U10004 (N_10004,N_9818,N_9857);
or U10005 (N_10005,N_9877,N_9970);
xor U10006 (N_10006,N_9991,N_9982);
nand U10007 (N_10007,N_9942,N_9875);
or U10008 (N_10008,N_9865,N_9842);
nand U10009 (N_10009,N_9917,N_9878);
nand U10010 (N_10010,N_9934,N_9859);
or U10011 (N_10011,N_9885,N_9994);
and U10012 (N_10012,N_9961,N_9902);
nand U10013 (N_10013,N_9940,N_9884);
and U10014 (N_10014,N_9834,N_9841);
nand U10015 (N_10015,N_9938,N_9922);
nand U10016 (N_10016,N_9847,N_9966);
nor U10017 (N_10017,N_9862,N_9883);
nor U10018 (N_10018,N_9930,N_9825);
or U10019 (N_10019,N_9969,N_9904);
nand U10020 (N_10020,N_9900,N_9879);
xor U10021 (N_10021,N_9999,N_9802);
nor U10022 (N_10022,N_9893,N_9891);
and U10023 (N_10023,N_9898,N_9926);
nor U10024 (N_10024,N_9824,N_9964);
nor U10025 (N_10025,N_9814,N_9952);
and U10026 (N_10026,N_9988,N_9908);
xnor U10027 (N_10027,N_9840,N_9913);
or U10028 (N_10028,N_9861,N_9910);
nor U10029 (N_10029,N_9803,N_9921);
xor U10030 (N_10030,N_9810,N_9983);
nor U10031 (N_10031,N_9989,N_9905);
nand U10032 (N_10032,N_9876,N_9974);
and U10033 (N_10033,N_9909,N_9874);
xnor U10034 (N_10034,N_9820,N_9906);
and U10035 (N_10035,N_9830,N_9967);
xnor U10036 (N_10036,N_9804,N_9960);
and U10037 (N_10037,N_9873,N_9945);
nor U10038 (N_10038,N_9920,N_9837);
nand U10039 (N_10039,N_9843,N_9984);
or U10040 (N_10040,N_9870,N_9950);
xnor U10041 (N_10041,N_9836,N_9943);
or U10042 (N_10042,N_9924,N_9936);
nand U10043 (N_10043,N_9998,N_9899);
xor U10044 (N_10044,N_9946,N_9918);
xnor U10045 (N_10045,N_9866,N_9829);
xnor U10046 (N_10046,N_9897,N_9951);
nor U10047 (N_10047,N_9808,N_9959);
xor U10048 (N_10048,N_9864,N_9911);
nand U10049 (N_10049,N_9932,N_9856);
xor U10050 (N_10050,N_9939,N_9823);
and U10051 (N_10051,N_9848,N_9812);
xor U10052 (N_10052,N_9933,N_9925);
nand U10053 (N_10053,N_9863,N_9963);
nand U10054 (N_10054,N_9809,N_9832);
nand U10055 (N_10055,N_9826,N_9860);
and U10056 (N_10056,N_9929,N_9901);
and U10057 (N_10057,N_9869,N_9995);
nand U10058 (N_10058,N_9935,N_9868);
or U10059 (N_10059,N_9968,N_9928);
nor U10060 (N_10060,N_9962,N_9839);
and U10061 (N_10061,N_9801,N_9976);
and U10062 (N_10062,N_9858,N_9919);
or U10063 (N_10063,N_9944,N_9817);
xor U10064 (N_10064,N_9806,N_9846);
xor U10065 (N_10065,N_9953,N_9957);
nor U10066 (N_10066,N_9977,N_9993);
xnor U10067 (N_10067,N_9854,N_9915);
or U10068 (N_10068,N_9931,N_9822);
nor U10069 (N_10069,N_9831,N_9838);
and U10070 (N_10070,N_9882,N_9971);
and U10071 (N_10071,N_9880,N_9800);
nor U10072 (N_10072,N_9815,N_9805);
and U10073 (N_10073,N_9886,N_9835);
nand U10074 (N_10074,N_9845,N_9907);
nand U10075 (N_10075,N_9986,N_9903);
or U10076 (N_10076,N_9849,N_9914);
or U10077 (N_10077,N_9980,N_9996);
and U10078 (N_10078,N_9985,N_9872);
nor U10079 (N_10079,N_9889,N_9992);
xnor U10080 (N_10080,N_9881,N_9819);
xor U10081 (N_10081,N_9892,N_9844);
or U10082 (N_10082,N_9894,N_9948);
nor U10083 (N_10083,N_9828,N_9947);
nand U10084 (N_10084,N_9821,N_9888);
and U10085 (N_10085,N_9955,N_9816);
and U10086 (N_10086,N_9990,N_9851);
xnor U10087 (N_10087,N_9916,N_9887);
nand U10088 (N_10088,N_9958,N_9827);
and U10089 (N_10089,N_9871,N_9895);
xnor U10090 (N_10090,N_9912,N_9833);
nor U10091 (N_10091,N_9956,N_9972);
or U10092 (N_10092,N_9807,N_9975);
nand U10093 (N_10093,N_9850,N_9890);
nand U10094 (N_10094,N_9853,N_9978);
and U10095 (N_10095,N_9981,N_9987);
nand U10096 (N_10096,N_9867,N_9965);
or U10097 (N_10097,N_9813,N_9997);
or U10098 (N_10098,N_9855,N_9927);
xnor U10099 (N_10099,N_9973,N_9896);
and U10100 (N_10100,N_9809,N_9831);
and U10101 (N_10101,N_9813,N_9820);
and U10102 (N_10102,N_9808,N_9819);
nor U10103 (N_10103,N_9879,N_9881);
nand U10104 (N_10104,N_9869,N_9953);
nor U10105 (N_10105,N_9978,N_9993);
xnor U10106 (N_10106,N_9982,N_9976);
xor U10107 (N_10107,N_9947,N_9907);
xor U10108 (N_10108,N_9931,N_9958);
nand U10109 (N_10109,N_9907,N_9980);
nor U10110 (N_10110,N_9883,N_9880);
and U10111 (N_10111,N_9802,N_9824);
xor U10112 (N_10112,N_9882,N_9897);
and U10113 (N_10113,N_9975,N_9902);
or U10114 (N_10114,N_9851,N_9833);
xor U10115 (N_10115,N_9804,N_9803);
xnor U10116 (N_10116,N_9913,N_9841);
xor U10117 (N_10117,N_9918,N_9935);
and U10118 (N_10118,N_9848,N_9851);
or U10119 (N_10119,N_9943,N_9845);
nor U10120 (N_10120,N_9836,N_9807);
xnor U10121 (N_10121,N_9874,N_9920);
nand U10122 (N_10122,N_9902,N_9969);
nand U10123 (N_10123,N_9879,N_9908);
and U10124 (N_10124,N_9923,N_9991);
or U10125 (N_10125,N_9823,N_9814);
xnor U10126 (N_10126,N_9925,N_9927);
nand U10127 (N_10127,N_9814,N_9815);
xor U10128 (N_10128,N_9857,N_9802);
and U10129 (N_10129,N_9929,N_9966);
or U10130 (N_10130,N_9841,N_9900);
and U10131 (N_10131,N_9806,N_9961);
nor U10132 (N_10132,N_9813,N_9842);
xor U10133 (N_10133,N_9864,N_9822);
and U10134 (N_10134,N_9941,N_9802);
nor U10135 (N_10135,N_9813,N_9831);
xor U10136 (N_10136,N_9925,N_9893);
or U10137 (N_10137,N_9842,N_9832);
nand U10138 (N_10138,N_9949,N_9811);
xor U10139 (N_10139,N_9985,N_9874);
and U10140 (N_10140,N_9855,N_9911);
or U10141 (N_10141,N_9912,N_9867);
nand U10142 (N_10142,N_9930,N_9943);
nand U10143 (N_10143,N_9948,N_9994);
or U10144 (N_10144,N_9884,N_9919);
and U10145 (N_10145,N_9831,N_9899);
and U10146 (N_10146,N_9841,N_9801);
xor U10147 (N_10147,N_9996,N_9955);
and U10148 (N_10148,N_9872,N_9926);
nand U10149 (N_10149,N_9908,N_9987);
xor U10150 (N_10150,N_9827,N_9924);
xnor U10151 (N_10151,N_9871,N_9916);
nor U10152 (N_10152,N_9960,N_9848);
and U10153 (N_10153,N_9964,N_9945);
or U10154 (N_10154,N_9966,N_9838);
and U10155 (N_10155,N_9932,N_9980);
or U10156 (N_10156,N_9802,N_9954);
and U10157 (N_10157,N_9955,N_9944);
or U10158 (N_10158,N_9865,N_9943);
xnor U10159 (N_10159,N_9938,N_9934);
or U10160 (N_10160,N_9853,N_9927);
nor U10161 (N_10161,N_9959,N_9964);
nor U10162 (N_10162,N_9851,N_9819);
or U10163 (N_10163,N_9833,N_9936);
xnor U10164 (N_10164,N_9800,N_9822);
and U10165 (N_10165,N_9958,N_9857);
nand U10166 (N_10166,N_9817,N_9851);
or U10167 (N_10167,N_9865,N_9916);
and U10168 (N_10168,N_9848,N_9920);
nor U10169 (N_10169,N_9832,N_9830);
nand U10170 (N_10170,N_9959,N_9809);
or U10171 (N_10171,N_9835,N_9849);
nor U10172 (N_10172,N_9835,N_9992);
and U10173 (N_10173,N_9847,N_9864);
or U10174 (N_10174,N_9807,N_9919);
nor U10175 (N_10175,N_9860,N_9834);
nor U10176 (N_10176,N_9833,N_9860);
and U10177 (N_10177,N_9816,N_9920);
xor U10178 (N_10178,N_9902,N_9998);
nor U10179 (N_10179,N_9801,N_9954);
xnor U10180 (N_10180,N_9813,N_9949);
and U10181 (N_10181,N_9964,N_9823);
or U10182 (N_10182,N_9802,N_9849);
nor U10183 (N_10183,N_9809,N_9830);
nand U10184 (N_10184,N_9849,N_9996);
nor U10185 (N_10185,N_9810,N_9994);
and U10186 (N_10186,N_9841,N_9907);
or U10187 (N_10187,N_9856,N_9990);
nand U10188 (N_10188,N_9929,N_9923);
xnor U10189 (N_10189,N_9809,N_9915);
and U10190 (N_10190,N_9992,N_9989);
nor U10191 (N_10191,N_9874,N_9870);
xnor U10192 (N_10192,N_9953,N_9980);
and U10193 (N_10193,N_9969,N_9947);
nand U10194 (N_10194,N_9800,N_9977);
or U10195 (N_10195,N_9895,N_9885);
and U10196 (N_10196,N_9860,N_9998);
or U10197 (N_10197,N_9892,N_9894);
nor U10198 (N_10198,N_9851,N_9876);
and U10199 (N_10199,N_9986,N_9987);
nor U10200 (N_10200,N_10153,N_10110);
nand U10201 (N_10201,N_10151,N_10025);
nand U10202 (N_10202,N_10032,N_10036);
nor U10203 (N_10203,N_10106,N_10146);
nand U10204 (N_10204,N_10194,N_10078);
or U10205 (N_10205,N_10026,N_10120);
xor U10206 (N_10206,N_10197,N_10053);
or U10207 (N_10207,N_10126,N_10012);
xnor U10208 (N_10208,N_10062,N_10001);
nand U10209 (N_10209,N_10184,N_10020);
nor U10210 (N_10210,N_10024,N_10190);
xor U10211 (N_10211,N_10162,N_10164);
nand U10212 (N_10212,N_10179,N_10135);
and U10213 (N_10213,N_10176,N_10065);
xnor U10214 (N_10214,N_10009,N_10119);
nand U10215 (N_10215,N_10134,N_10041);
nor U10216 (N_10216,N_10084,N_10122);
nor U10217 (N_10217,N_10014,N_10155);
nand U10218 (N_10218,N_10127,N_10133);
and U10219 (N_10219,N_10035,N_10088);
and U10220 (N_10220,N_10192,N_10031);
xnor U10221 (N_10221,N_10073,N_10067);
and U10222 (N_10222,N_10163,N_10008);
nand U10223 (N_10223,N_10089,N_10158);
or U10224 (N_10224,N_10118,N_10030);
or U10225 (N_10225,N_10125,N_10095);
or U10226 (N_10226,N_10028,N_10047);
xnor U10227 (N_10227,N_10058,N_10108);
or U10228 (N_10228,N_10027,N_10079);
xnor U10229 (N_10229,N_10005,N_10165);
nor U10230 (N_10230,N_10150,N_10191);
nand U10231 (N_10231,N_10104,N_10172);
nand U10232 (N_10232,N_10016,N_10038);
or U10233 (N_10233,N_10050,N_10137);
nor U10234 (N_10234,N_10174,N_10139);
or U10235 (N_10235,N_10037,N_10098);
nand U10236 (N_10236,N_10066,N_10044);
xnor U10237 (N_10237,N_10193,N_10013);
nand U10238 (N_10238,N_10018,N_10010);
or U10239 (N_10239,N_10070,N_10096);
and U10240 (N_10240,N_10007,N_10019);
or U10241 (N_10241,N_10186,N_10034);
and U10242 (N_10242,N_10107,N_10132);
nand U10243 (N_10243,N_10081,N_10130);
or U10244 (N_10244,N_10136,N_10171);
nand U10245 (N_10245,N_10170,N_10011);
xor U10246 (N_10246,N_10188,N_10094);
nand U10247 (N_10247,N_10000,N_10090);
nor U10248 (N_10248,N_10112,N_10195);
nand U10249 (N_10249,N_10059,N_10183);
or U10250 (N_10250,N_10068,N_10128);
xnor U10251 (N_10251,N_10156,N_10131);
nand U10252 (N_10252,N_10141,N_10092);
xor U10253 (N_10253,N_10046,N_10085);
or U10254 (N_10254,N_10033,N_10004);
nand U10255 (N_10255,N_10198,N_10097);
nor U10256 (N_10256,N_10083,N_10076);
nand U10257 (N_10257,N_10178,N_10077);
nand U10258 (N_10258,N_10057,N_10121);
nand U10259 (N_10259,N_10180,N_10091);
xor U10260 (N_10260,N_10093,N_10167);
or U10261 (N_10261,N_10087,N_10111);
nand U10262 (N_10262,N_10115,N_10023);
or U10263 (N_10263,N_10154,N_10143);
nand U10264 (N_10264,N_10051,N_10185);
and U10265 (N_10265,N_10074,N_10075);
nor U10266 (N_10266,N_10022,N_10086);
nor U10267 (N_10267,N_10166,N_10039);
nor U10268 (N_10268,N_10152,N_10103);
or U10269 (N_10269,N_10182,N_10147);
or U10270 (N_10270,N_10105,N_10177);
nand U10271 (N_10271,N_10117,N_10080);
and U10272 (N_10272,N_10049,N_10064);
and U10273 (N_10273,N_10124,N_10144);
nand U10274 (N_10274,N_10148,N_10129);
nand U10275 (N_10275,N_10017,N_10006);
xor U10276 (N_10276,N_10100,N_10056);
nand U10277 (N_10277,N_10045,N_10113);
or U10278 (N_10278,N_10102,N_10189);
or U10279 (N_10279,N_10002,N_10060);
nor U10280 (N_10280,N_10029,N_10175);
or U10281 (N_10281,N_10160,N_10043);
nor U10282 (N_10282,N_10054,N_10161);
nand U10283 (N_10283,N_10003,N_10159);
and U10284 (N_10284,N_10101,N_10199);
xor U10285 (N_10285,N_10116,N_10140);
and U10286 (N_10286,N_10069,N_10055);
nand U10287 (N_10287,N_10149,N_10021);
nor U10288 (N_10288,N_10052,N_10181);
nor U10289 (N_10289,N_10061,N_10048);
xor U10290 (N_10290,N_10173,N_10099);
xnor U10291 (N_10291,N_10082,N_10063);
or U10292 (N_10292,N_10072,N_10109);
and U10293 (N_10293,N_10157,N_10040);
or U10294 (N_10294,N_10169,N_10042);
nand U10295 (N_10295,N_10187,N_10142);
or U10296 (N_10296,N_10015,N_10114);
and U10297 (N_10297,N_10168,N_10138);
nor U10298 (N_10298,N_10071,N_10145);
or U10299 (N_10299,N_10196,N_10123);
xor U10300 (N_10300,N_10067,N_10182);
and U10301 (N_10301,N_10182,N_10025);
nand U10302 (N_10302,N_10095,N_10056);
nand U10303 (N_10303,N_10092,N_10050);
xor U10304 (N_10304,N_10124,N_10130);
or U10305 (N_10305,N_10042,N_10152);
nand U10306 (N_10306,N_10020,N_10069);
xor U10307 (N_10307,N_10043,N_10012);
and U10308 (N_10308,N_10087,N_10157);
or U10309 (N_10309,N_10091,N_10010);
nor U10310 (N_10310,N_10123,N_10095);
nand U10311 (N_10311,N_10059,N_10166);
nand U10312 (N_10312,N_10015,N_10143);
nand U10313 (N_10313,N_10033,N_10118);
xnor U10314 (N_10314,N_10170,N_10148);
nand U10315 (N_10315,N_10158,N_10117);
nor U10316 (N_10316,N_10033,N_10122);
or U10317 (N_10317,N_10072,N_10143);
and U10318 (N_10318,N_10068,N_10171);
nand U10319 (N_10319,N_10150,N_10029);
nor U10320 (N_10320,N_10197,N_10021);
nor U10321 (N_10321,N_10138,N_10114);
or U10322 (N_10322,N_10024,N_10048);
nor U10323 (N_10323,N_10066,N_10088);
nand U10324 (N_10324,N_10064,N_10109);
or U10325 (N_10325,N_10156,N_10128);
nor U10326 (N_10326,N_10011,N_10112);
or U10327 (N_10327,N_10114,N_10198);
nand U10328 (N_10328,N_10012,N_10135);
xnor U10329 (N_10329,N_10148,N_10160);
and U10330 (N_10330,N_10123,N_10126);
nor U10331 (N_10331,N_10163,N_10172);
nand U10332 (N_10332,N_10026,N_10049);
or U10333 (N_10333,N_10136,N_10186);
nor U10334 (N_10334,N_10162,N_10104);
nor U10335 (N_10335,N_10009,N_10167);
or U10336 (N_10336,N_10027,N_10034);
xnor U10337 (N_10337,N_10193,N_10044);
and U10338 (N_10338,N_10183,N_10131);
xor U10339 (N_10339,N_10054,N_10024);
and U10340 (N_10340,N_10160,N_10058);
and U10341 (N_10341,N_10129,N_10136);
xor U10342 (N_10342,N_10193,N_10122);
and U10343 (N_10343,N_10143,N_10023);
nand U10344 (N_10344,N_10192,N_10006);
nand U10345 (N_10345,N_10006,N_10083);
and U10346 (N_10346,N_10185,N_10063);
nand U10347 (N_10347,N_10080,N_10152);
and U10348 (N_10348,N_10014,N_10138);
xor U10349 (N_10349,N_10106,N_10122);
nand U10350 (N_10350,N_10164,N_10116);
xor U10351 (N_10351,N_10180,N_10199);
and U10352 (N_10352,N_10168,N_10180);
nor U10353 (N_10353,N_10055,N_10085);
xor U10354 (N_10354,N_10002,N_10198);
nand U10355 (N_10355,N_10002,N_10122);
and U10356 (N_10356,N_10056,N_10156);
nand U10357 (N_10357,N_10074,N_10064);
nor U10358 (N_10358,N_10150,N_10087);
or U10359 (N_10359,N_10081,N_10082);
or U10360 (N_10360,N_10022,N_10177);
and U10361 (N_10361,N_10182,N_10007);
or U10362 (N_10362,N_10091,N_10120);
nor U10363 (N_10363,N_10065,N_10024);
xnor U10364 (N_10364,N_10086,N_10196);
nand U10365 (N_10365,N_10105,N_10020);
nand U10366 (N_10366,N_10002,N_10026);
and U10367 (N_10367,N_10021,N_10000);
nor U10368 (N_10368,N_10123,N_10102);
xor U10369 (N_10369,N_10140,N_10059);
or U10370 (N_10370,N_10175,N_10155);
nand U10371 (N_10371,N_10053,N_10117);
nand U10372 (N_10372,N_10077,N_10072);
or U10373 (N_10373,N_10030,N_10183);
xor U10374 (N_10374,N_10157,N_10176);
xnor U10375 (N_10375,N_10161,N_10137);
nor U10376 (N_10376,N_10182,N_10145);
nand U10377 (N_10377,N_10024,N_10082);
nor U10378 (N_10378,N_10032,N_10000);
nor U10379 (N_10379,N_10109,N_10014);
nand U10380 (N_10380,N_10000,N_10188);
nand U10381 (N_10381,N_10159,N_10051);
and U10382 (N_10382,N_10042,N_10104);
nor U10383 (N_10383,N_10140,N_10107);
nor U10384 (N_10384,N_10042,N_10044);
nand U10385 (N_10385,N_10195,N_10028);
and U10386 (N_10386,N_10183,N_10054);
and U10387 (N_10387,N_10172,N_10151);
xor U10388 (N_10388,N_10026,N_10156);
or U10389 (N_10389,N_10050,N_10099);
or U10390 (N_10390,N_10195,N_10036);
nor U10391 (N_10391,N_10017,N_10170);
nand U10392 (N_10392,N_10126,N_10169);
or U10393 (N_10393,N_10071,N_10056);
nor U10394 (N_10394,N_10059,N_10066);
or U10395 (N_10395,N_10006,N_10155);
and U10396 (N_10396,N_10058,N_10195);
and U10397 (N_10397,N_10099,N_10199);
nand U10398 (N_10398,N_10136,N_10177);
xor U10399 (N_10399,N_10087,N_10063);
nand U10400 (N_10400,N_10242,N_10204);
nand U10401 (N_10401,N_10208,N_10259);
nand U10402 (N_10402,N_10226,N_10231);
nor U10403 (N_10403,N_10333,N_10292);
xor U10404 (N_10404,N_10367,N_10206);
nor U10405 (N_10405,N_10326,N_10214);
or U10406 (N_10406,N_10249,N_10230);
nand U10407 (N_10407,N_10350,N_10276);
and U10408 (N_10408,N_10235,N_10247);
nor U10409 (N_10409,N_10274,N_10284);
or U10410 (N_10410,N_10312,N_10321);
or U10411 (N_10411,N_10303,N_10228);
and U10412 (N_10412,N_10396,N_10310);
nand U10413 (N_10413,N_10253,N_10278);
nand U10414 (N_10414,N_10239,N_10384);
xnor U10415 (N_10415,N_10313,N_10212);
xnor U10416 (N_10416,N_10366,N_10252);
nor U10417 (N_10417,N_10338,N_10387);
and U10418 (N_10418,N_10322,N_10348);
or U10419 (N_10419,N_10265,N_10325);
and U10420 (N_10420,N_10223,N_10304);
nand U10421 (N_10421,N_10320,N_10262);
and U10422 (N_10422,N_10332,N_10237);
nand U10423 (N_10423,N_10341,N_10364);
nor U10424 (N_10424,N_10275,N_10219);
xnor U10425 (N_10425,N_10296,N_10393);
and U10426 (N_10426,N_10377,N_10391);
xnor U10427 (N_10427,N_10203,N_10392);
xor U10428 (N_10428,N_10314,N_10246);
nor U10429 (N_10429,N_10297,N_10243);
nand U10430 (N_10430,N_10395,N_10373);
or U10431 (N_10431,N_10258,N_10245);
nand U10432 (N_10432,N_10329,N_10376);
nand U10433 (N_10433,N_10291,N_10268);
xor U10434 (N_10434,N_10300,N_10222);
nor U10435 (N_10435,N_10316,N_10397);
nand U10436 (N_10436,N_10398,N_10240);
or U10437 (N_10437,N_10345,N_10357);
xor U10438 (N_10438,N_10279,N_10361);
xor U10439 (N_10439,N_10273,N_10368);
xnor U10440 (N_10440,N_10359,N_10352);
and U10441 (N_10441,N_10374,N_10250);
nand U10442 (N_10442,N_10317,N_10381);
or U10443 (N_10443,N_10379,N_10383);
nand U10444 (N_10444,N_10285,N_10290);
xor U10445 (N_10445,N_10336,N_10389);
nor U10446 (N_10446,N_10347,N_10264);
and U10447 (N_10447,N_10287,N_10318);
nor U10448 (N_10448,N_10390,N_10324);
or U10449 (N_10449,N_10369,N_10309);
or U10450 (N_10450,N_10207,N_10355);
xnor U10451 (N_10451,N_10209,N_10351);
xnor U10452 (N_10452,N_10305,N_10362);
or U10453 (N_10453,N_10319,N_10280);
and U10454 (N_10454,N_10344,N_10202);
xnor U10455 (N_10455,N_10233,N_10220);
xor U10456 (N_10456,N_10328,N_10261);
nand U10457 (N_10457,N_10210,N_10380);
nor U10458 (N_10458,N_10306,N_10358);
nor U10459 (N_10459,N_10386,N_10238);
or U10460 (N_10460,N_10378,N_10311);
and U10461 (N_10461,N_10339,N_10271);
xnor U10462 (N_10462,N_10382,N_10349);
nand U10463 (N_10463,N_10331,N_10283);
nand U10464 (N_10464,N_10353,N_10307);
xnor U10465 (N_10465,N_10255,N_10372);
and U10466 (N_10466,N_10354,N_10236);
nor U10467 (N_10467,N_10330,N_10257);
and U10468 (N_10468,N_10363,N_10327);
xor U10469 (N_10469,N_10360,N_10301);
nor U10470 (N_10470,N_10371,N_10346);
xnor U10471 (N_10471,N_10269,N_10298);
or U10472 (N_10472,N_10343,N_10263);
nor U10473 (N_10473,N_10286,N_10272);
nor U10474 (N_10474,N_10234,N_10248);
or U10475 (N_10475,N_10201,N_10241);
nor U10476 (N_10476,N_10299,N_10356);
nand U10477 (N_10477,N_10337,N_10288);
nor U10478 (N_10478,N_10293,N_10254);
nor U10479 (N_10479,N_10213,N_10244);
or U10480 (N_10480,N_10266,N_10323);
and U10481 (N_10481,N_10281,N_10217);
nand U10482 (N_10482,N_10335,N_10315);
and U10483 (N_10483,N_10218,N_10388);
and U10484 (N_10484,N_10277,N_10308);
nor U10485 (N_10485,N_10251,N_10229);
nand U10486 (N_10486,N_10267,N_10216);
xor U10487 (N_10487,N_10200,N_10375);
nand U10488 (N_10488,N_10256,N_10224);
or U10489 (N_10489,N_10282,N_10225);
or U10490 (N_10490,N_10232,N_10260);
or U10491 (N_10491,N_10295,N_10205);
or U10492 (N_10492,N_10385,N_10394);
xnor U10493 (N_10493,N_10215,N_10399);
nand U10494 (N_10494,N_10227,N_10340);
nor U10495 (N_10495,N_10270,N_10370);
or U10496 (N_10496,N_10289,N_10334);
and U10497 (N_10497,N_10294,N_10365);
and U10498 (N_10498,N_10302,N_10342);
xor U10499 (N_10499,N_10211,N_10221);
nor U10500 (N_10500,N_10315,N_10273);
and U10501 (N_10501,N_10342,N_10316);
xnor U10502 (N_10502,N_10291,N_10334);
nor U10503 (N_10503,N_10342,N_10219);
xnor U10504 (N_10504,N_10393,N_10283);
nand U10505 (N_10505,N_10295,N_10219);
or U10506 (N_10506,N_10375,N_10209);
nand U10507 (N_10507,N_10364,N_10363);
nand U10508 (N_10508,N_10295,N_10264);
nand U10509 (N_10509,N_10349,N_10294);
or U10510 (N_10510,N_10356,N_10221);
xnor U10511 (N_10511,N_10225,N_10363);
or U10512 (N_10512,N_10367,N_10373);
nor U10513 (N_10513,N_10227,N_10324);
or U10514 (N_10514,N_10332,N_10246);
nand U10515 (N_10515,N_10284,N_10300);
xnor U10516 (N_10516,N_10215,N_10201);
nor U10517 (N_10517,N_10229,N_10210);
and U10518 (N_10518,N_10290,N_10215);
nor U10519 (N_10519,N_10334,N_10254);
or U10520 (N_10520,N_10247,N_10297);
xor U10521 (N_10521,N_10392,N_10275);
and U10522 (N_10522,N_10264,N_10282);
nand U10523 (N_10523,N_10280,N_10348);
and U10524 (N_10524,N_10387,N_10221);
or U10525 (N_10525,N_10316,N_10224);
xnor U10526 (N_10526,N_10280,N_10263);
nor U10527 (N_10527,N_10363,N_10319);
nand U10528 (N_10528,N_10358,N_10304);
nor U10529 (N_10529,N_10223,N_10375);
xor U10530 (N_10530,N_10308,N_10361);
nor U10531 (N_10531,N_10337,N_10275);
and U10532 (N_10532,N_10271,N_10285);
nand U10533 (N_10533,N_10206,N_10333);
nor U10534 (N_10534,N_10360,N_10354);
nor U10535 (N_10535,N_10203,N_10394);
xnor U10536 (N_10536,N_10248,N_10299);
or U10537 (N_10537,N_10280,N_10351);
nor U10538 (N_10538,N_10262,N_10325);
and U10539 (N_10539,N_10318,N_10399);
xnor U10540 (N_10540,N_10299,N_10321);
nand U10541 (N_10541,N_10294,N_10314);
and U10542 (N_10542,N_10220,N_10200);
xnor U10543 (N_10543,N_10315,N_10274);
nor U10544 (N_10544,N_10324,N_10278);
and U10545 (N_10545,N_10381,N_10268);
and U10546 (N_10546,N_10317,N_10229);
or U10547 (N_10547,N_10297,N_10369);
nand U10548 (N_10548,N_10205,N_10258);
nor U10549 (N_10549,N_10378,N_10233);
xor U10550 (N_10550,N_10334,N_10210);
nor U10551 (N_10551,N_10283,N_10284);
xor U10552 (N_10552,N_10391,N_10245);
and U10553 (N_10553,N_10319,N_10356);
and U10554 (N_10554,N_10333,N_10353);
nor U10555 (N_10555,N_10343,N_10228);
xnor U10556 (N_10556,N_10273,N_10258);
nand U10557 (N_10557,N_10264,N_10346);
or U10558 (N_10558,N_10276,N_10310);
nor U10559 (N_10559,N_10299,N_10355);
nor U10560 (N_10560,N_10255,N_10264);
and U10561 (N_10561,N_10376,N_10356);
and U10562 (N_10562,N_10204,N_10380);
nor U10563 (N_10563,N_10266,N_10307);
or U10564 (N_10564,N_10264,N_10324);
and U10565 (N_10565,N_10349,N_10223);
and U10566 (N_10566,N_10382,N_10201);
and U10567 (N_10567,N_10218,N_10248);
or U10568 (N_10568,N_10284,N_10390);
or U10569 (N_10569,N_10214,N_10382);
nor U10570 (N_10570,N_10326,N_10246);
or U10571 (N_10571,N_10246,N_10327);
nor U10572 (N_10572,N_10299,N_10288);
or U10573 (N_10573,N_10204,N_10263);
nand U10574 (N_10574,N_10204,N_10327);
nand U10575 (N_10575,N_10318,N_10337);
xor U10576 (N_10576,N_10321,N_10351);
xnor U10577 (N_10577,N_10364,N_10311);
nand U10578 (N_10578,N_10363,N_10305);
and U10579 (N_10579,N_10226,N_10368);
xnor U10580 (N_10580,N_10393,N_10377);
and U10581 (N_10581,N_10399,N_10240);
nor U10582 (N_10582,N_10367,N_10259);
nor U10583 (N_10583,N_10244,N_10264);
and U10584 (N_10584,N_10329,N_10391);
xor U10585 (N_10585,N_10269,N_10225);
xor U10586 (N_10586,N_10223,N_10267);
xnor U10587 (N_10587,N_10289,N_10268);
nand U10588 (N_10588,N_10348,N_10359);
and U10589 (N_10589,N_10225,N_10204);
and U10590 (N_10590,N_10324,N_10218);
nor U10591 (N_10591,N_10329,N_10263);
nand U10592 (N_10592,N_10241,N_10207);
nor U10593 (N_10593,N_10305,N_10285);
and U10594 (N_10594,N_10214,N_10263);
nand U10595 (N_10595,N_10246,N_10224);
or U10596 (N_10596,N_10249,N_10333);
xor U10597 (N_10597,N_10280,N_10246);
and U10598 (N_10598,N_10222,N_10282);
nand U10599 (N_10599,N_10274,N_10312);
and U10600 (N_10600,N_10483,N_10499);
and U10601 (N_10601,N_10440,N_10430);
or U10602 (N_10602,N_10505,N_10422);
nand U10603 (N_10603,N_10509,N_10524);
nand U10604 (N_10604,N_10474,N_10542);
nor U10605 (N_10605,N_10516,N_10508);
xnor U10606 (N_10606,N_10555,N_10530);
nor U10607 (N_10607,N_10460,N_10565);
and U10608 (N_10608,N_10437,N_10598);
and U10609 (N_10609,N_10464,N_10533);
nor U10610 (N_10610,N_10482,N_10506);
and U10611 (N_10611,N_10432,N_10445);
xor U10612 (N_10612,N_10574,N_10449);
and U10613 (N_10613,N_10580,N_10456);
nand U10614 (N_10614,N_10411,N_10402);
nand U10615 (N_10615,N_10450,N_10475);
or U10616 (N_10616,N_10517,N_10541);
xnor U10617 (N_10617,N_10504,N_10590);
and U10618 (N_10618,N_10447,N_10557);
nor U10619 (N_10619,N_10481,N_10407);
and U10620 (N_10620,N_10543,N_10549);
nor U10621 (N_10621,N_10492,N_10438);
and U10622 (N_10622,N_10562,N_10409);
nor U10623 (N_10623,N_10434,N_10412);
and U10624 (N_10624,N_10514,N_10502);
nor U10625 (N_10625,N_10406,N_10540);
xor U10626 (N_10626,N_10489,N_10400);
nor U10627 (N_10627,N_10408,N_10578);
xnor U10628 (N_10628,N_10503,N_10573);
or U10629 (N_10629,N_10446,N_10468);
nor U10630 (N_10630,N_10522,N_10585);
and U10631 (N_10631,N_10419,N_10515);
and U10632 (N_10632,N_10424,N_10576);
nor U10633 (N_10633,N_10403,N_10435);
nor U10634 (N_10634,N_10518,N_10444);
nor U10635 (N_10635,N_10485,N_10563);
or U10636 (N_10636,N_10535,N_10581);
or U10637 (N_10637,N_10548,N_10421);
or U10638 (N_10638,N_10495,N_10560);
xnor U10639 (N_10639,N_10528,N_10554);
nor U10640 (N_10640,N_10488,N_10561);
xnor U10641 (N_10641,N_10582,N_10410);
nand U10642 (N_10642,N_10591,N_10599);
xor U10643 (N_10643,N_10457,N_10583);
or U10644 (N_10644,N_10427,N_10521);
and U10645 (N_10645,N_10507,N_10420);
or U10646 (N_10646,N_10595,N_10458);
nand U10647 (N_10647,N_10428,N_10480);
nor U10648 (N_10648,N_10593,N_10526);
xnor U10649 (N_10649,N_10415,N_10531);
nand U10650 (N_10650,N_10426,N_10550);
xor U10651 (N_10651,N_10529,N_10463);
nand U10652 (N_10652,N_10594,N_10476);
xnor U10653 (N_10653,N_10559,N_10567);
or U10654 (N_10654,N_10575,N_10417);
xnor U10655 (N_10655,N_10493,N_10498);
or U10656 (N_10656,N_10404,N_10461);
or U10657 (N_10657,N_10500,N_10572);
and U10658 (N_10658,N_10441,N_10545);
nand U10659 (N_10659,N_10442,N_10443);
and U10660 (N_10660,N_10587,N_10436);
or U10661 (N_10661,N_10433,N_10484);
nor U10662 (N_10662,N_10425,N_10405);
or U10663 (N_10663,N_10451,N_10538);
or U10664 (N_10664,N_10423,N_10466);
or U10665 (N_10665,N_10553,N_10494);
nor U10666 (N_10666,N_10588,N_10523);
or U10667 (N_10667,N_10592,N_10596);
nor U10668 (N_10668,N_10544,N_10527);
xor U10669 (N_10669,N_10577,N_10497);
nor U10670 (N_10670,N_10501,N_10431);
or U10671 (N_10671,N_10439,N_10534);
or U10672 (N_10672,N_10416,N_10459);
xnor U10673 (N_10673,N_10453,N_10586);
nand U10674 (N_10674,N_10552,N_10584);
nand U10675 (N_10675,N_10547,N_10520);
or U10676 (N_10676,N_10539,N_10566);
nor U10677 (N_10677,N_10571,N_10551);
and U10678 (N_10678,N_10470,N_10569);
xnor U10679 (N_10679,N_10511,N_10487);
or U10680 (N_10680,N_10471,N_10532);
and U10681 (N_10681,N_10589,N_10472);
or U10682 (N_10682,N_10564,N_10414);
and U10683 (N_10683,N_10479,N_10455);
or U10684 (N_10684,N_10452,N_10448);
and U10685 (N_10685,N_10570,N_10469);
or U10686 (N_10686,N_10537,N_10513);
xor U10687 (N_10687,N_10467,N_10536);
and U10688 (N_10688,N_10473,N_10579);
or U10689 (N_10689,N_10546,N_10512);
xnor U10690 (N_10690,N_10429,N_10486);
nor U10691 (N_10691,N_10418,N_10465);
or U10692 (N_10692,N_10556,N_10525);
nor U10693 (N_10693,N_10413,N_10490);
nand U10694 (N_10694,N_10510,N_10519);
and U10695 (N_10695,N_10478,N_10491);
and U10696 (N_10696,N_10558,N_10568);
xnor U10697 (N_10697,N_10597,N_10462);
or U10698 (N_10698,N_10454,N_10477);
or U10699 (N_10699,N_10401,N_10496);
and U10700 (N_10700,N_10502,N_10551);
nor U10701 (N_10701,N_10440,N_10416);
and U10702 (N_10702,N_10429,N_10537);
nand U10703 (N_10703,N_10583,N_10592);
nor U10704 (N_10704,N_10544,N_10506);
xor U10705 (N_10705,N_10415,N_10402);
or U10706 (N_10706,N_10596,N_10496);
and U10707 (N_10707,N_10486,N_10551);
nor U10708 (N_10708,N_10468,N_10438);
and U10709 (N_10709,N_10505,N_10464);
and U10710 (N_10710,N_10423,N_10500);
nand U10711 (N_10711,N_10502,N_10599);
xor U10712 (N_10712,N_10574,N_10563);
xor U10713 (N_10713,N_10580,N_10561);
or U10714 (N_10714,N_10513,N_10463);
nor U10715 (N_10715,N_10558,N_10579);
nor U10716 (N_10716,N_10504,N_10533);
nor U10717 (N_10717,N_10598,N_10475);
nor U10718 (N_10718,N_10496,N_10593);
or U10719 (N_10719,N_10450,N_10500);
nor U10720 (N_10720,N_10485,N_10595);
and U10721 (N_10721,N_10569,N_10418);
xnor U10722 (N_10722,N_10481,N_10419);
or U10723 (N_10723,N_10433,N_10483);
nor U10724 (N_10724,N_10568,N_10419);
or U10725 (N_10725,N_10535,N_10457);
or U10726 (N_10726,N_10595,N_10567);
nor U10727 (N_10727,N_10586,N_10443);
and U10728 (N_10728,N_10460,N_10501);
nand U10729 (N_10729,N_10470,N_10418);
xnor U10730 (N_10730,N_10584,N_10599);
or U10731 (N_10731,N_10523,N_10477);
and U10732 (N_10732,N_10473,N_10537);
nand U10733 (N_10733,N_10510,N_10526);
or U10734 (N_10734,N_10553,N_10509);
xor U10735 (N_10735,N_10562,N_10592);
and U10736 (N_10736,N_10565,N_10498);
nor U10737 (N_10737,N_10475,N_10530);
nand U10738 (N_10738,N_10544,N_10436);
or U10739 (N_10739,N_10426,N_10551);
nand U10740 (N_10740,N_10567,N_10573);
nand U10741 (N_10741,N_10517,N_10468);
nand U10742 (N_10742,N_10590,N_10572);
xor U10743 (N_10743,N_10442,N_10517);
nor U10744 (N_10744,N_10406,N_10439);
xor U10745 (N_10745,N_10417,N_10574);
or U10746 (N_10746,N_10570,N_10540);
nand U10747 (N_10747,N_10537,N_10577);
xor U10748 (N_10748,N_10451,N_10412);
nand U10749 (N_10749,N_10480,N_10417);
xnor U10750 (N_10750,N_10415,N_10547);
nand U10751 (N_10751,N_10554,N_10406);
nand U10752 (N_10752,N_10481,N_10534);
and U10753 (N_10753,N_10535,N_10431);
nor U10754 (N_10754,N_10416,N_10420);
and U10755 (N_10755,N_10526,N_10571);
nand U10756 (N_10756,N_10534,N_10436);
nand U10757 (N_10757,N_10485,N_10400);
nand U10758 (N_10758,N_10482,N_10481);
or U10759 (N_10759,N_10554,N_10459);
xor U10760 (N_10760,N_10414,N_10401);
or U10761 (N_10761,N_10592,N_10440);
and U10762 (N_10762,N_10507,N_10427);
or U10763 (N_10763,N_10569,N_10578);
nor U10764 (N_10764,N_10575,N_10563);
nor U10765 (N_10765,N_10548,N_10474);
nand U10766 (N_10766,N_10593,N_10590);
nor U10767 (N_10767,N_10429,N_10492);
xnor U10768 (N_10768,N_10553,N_10506);
xor U10769 (N_10769,N_10439,N_10468);
nand U10770 (N_10770,N_10499,N_10415);
xor U10771 (N_10771,N_10577,N_10416);
and U10772 (N_10772,N_10573,N_10423);
and U10773 (N_10773,N_10571,N_10461);
or U10774 (N_10774,N_10572,N_10485);
nor U10775 (N_10775,N_10546,N_10574);
xor U10776 (N_10776,N_10479,N_10572);
xnor U10777 (N_10777,N_10578,N_10503);
xor U10778 (N_10778,N_10496,N_10442);
or U10779 (N_10779,N_10543,N_10402);
xor U10780 (N_10780,N_10447,N_10507);
nand U10781 (N_10781,N_10575,N_10404);
nor U10782 (N_10782,N_10403,N_10597);
and U10783 (N_10783,N_10417,N_10558);
nor U10784 (N_10784,N_10587,N_10519);
nand U10785 (N_10785,N_10416,N_10450);
and U10786 (N_10786,N_10474,N_10408);
or U10787 (N_10787,N_10581,N_10477);
or U10788 (N_10788,N_10468,N_10400);
xor U10789 (N_10789,N_10491,N_10506);
nor U10790 (N_10790,N_10460,N_10441);
xor U10791 (N_10791,N_10515,N_10547);
and U10792 (N_10792,N_10469,N_10444);
nor U10793 (N_10793,N_10506,N_10562);
or U10794 (N_10794,N_10519,N_10539);
nand U10795 (N_10795,N_10597,N_10473);
xor U10796 (N_10796,N_10417,N_10569);
or U10797 (N_10797,N_10544,N_10406);
nand U10798 (N_10798,N_10557,N_10555);
or U10799 (N_10799,N_10405,N_10599);
nand U10800 (N_10800,N_10720,N_10600);
and U10801 (N_10801,N_10798,N_10779);
nand U10802 (N_10802,N_10791,N_10755);
xnor U10803 (N_10803,N_10646,N_10612);
nand U10804 (N_10804,N_10776,N_10674);
nor U10805 (N_10805,N_10744,N_10604);
nand U10806 (N_10806,N_10774,N_10635);
nor U10807 (N_10807,N_10777,N_10648);
or U10808 (N_10808,N_10796,N_10641);
and U10809 (N_10809,N_10636,N_10708);
nor U10810 (N_10810,N_10726,N_10675);
and U10811 (N_10811,N_10727,N_10692);
xor U10812 (N_10812,N_10664,N_10799);
nand U10813 (N_10813,N_10792,N_10704);
nor U10814 (N_10814,N_10683,N_10741);
or U10815 (N_10815,N_10676,N_10623);
or U10816 (N_10816,N_10723,N_10733);
nand U10817 (N_10817,N_10647,N_10687);
xor U10818 (N_10818,N_10601,N_10761);
nor U10819 (N_10819,N_10689,N_10719);
xor U10820 (N_10820,N_10637,N_10628);
xnor U10821 (N_10821,N_10681,N_10632);
nor U10822 (N_10822,N_10633,N_10669);
nor U10823 (N_10823,N_10721,N_10619);
nor U10824 (N_10824,N_10668,N_10758);
xnor U10825 (N_10825,N_10609,N_10614);
or U10826 (N_10826,N_10642,N_10728);
or U10827 (N_10827,N_10672,N_10724);
nor U10828 (N_10828,N_10650,N_10762);
nor U10829 (N_10829,N_10731,N_10794);
or U10830 (N_10830,N_10760,N_10662);
xor U10831 (N_10831,N_10678,N_10736);
or U10832 (N_10832,N_10665,N_10702);
nand U10833 (N_10833,N_10691,N_10643);
xnor U10834 (N_10834,N_10603,N_10608);
and U10835 (N_10835,N_10686,N_10706);
and U10836 (N_10836,N_10782,N_10732);
nor U10837 (N_10837,N_10729,N_10640);
nor U10838 (N_10838,N_10751,N_10671);
and U10839 (N_10839,N_10620,N_10673);
nor U10840 (N_10840,N_10630,N_10716);
xnor U10841 (N_10841,N_10784,N_10626);
nor U10842 (N_10842,N_10747,N_10666);
or U10843 (N_10843,N_10622,N_10763);
nand U10844 (N_10844,N_10700,N_10625);
and U10845 (N_10845,N_10655,N_10737);
xor U10846 (N_10846,N_10611,N_10739);
and U10847 (N_10847,N_10746,N_10605);
nand U10848 (N_10848,N_10639,N_10621);
nand U10849 (N_10849,N_10615,N_10772);
or U10850 (N_10850,N_10773,N_10771);
nand U10851 (N_10851,N_10682,N_10734);
nor U10852 (N_10852,N_10789,N_10607);
nor U10853 (N_10853,N_10742,N_10765);
xor U10854 (N_10854,N_10653,N_10712);
nor U10855 (N_10855,N_10645,N_10752);
nor U10856 (N_10856,N_10780,N_10688);
and U10857 (N_10857,N_10748,N_10698);
or U10858 (N_10858,N_10606,N_10616);
xnor U10859 (N_10859,N_10695,N_10663);
nand U10860 (N_10860,N_10667,N_10649);
and U10861 (N_10861,N_10738,N_10694);
nand U10862 (N_10862,N_10631,N_10644);
or U10863 (N_10863,N_10699,N_10617);
xor U10864 (N_10864,N_10743,N_10713);
xor U10865 (N_10865,N_10654,N_10705);
or U10866 (N_10866,N_10679,N_10745);
or U10867 (N_10867,N_10714,N_10753);
or U10868 (N_10868,N_10781,N_10710);
nor U10869 (N_10869,N_10775,N_10627);
or U10870 (N_10870,N_10764,N_10717);
nand U10871 (N_10871,N_10754,N_10759);
xnor U10872 (N_10872,N_10711,N_10749);
nor U10873 (N_10873,N_10680,N_10660);
and U10874 (N_10874,N_10656,N_10659);
and U10875 (N_10875,N_10602,N_10661);
or U10876 (N_10876,N_10652,N_10703);
and U10877 (N_10877,N_10718,N_10657);
nor U10878 (N_10878,N_10767,N_10788);
or U10879 (N_10879,N_10618,N_10707);
nand U10880 (N_10880,N_10786,N_10790);
nand U10881 (N_10881,N_10768,N_10769);
and U10882 (N_10882,N_10709,N_10735);
nor U10883 (N_10883,N_10613,N_10690);
and U10884 (N_10884,N_10685,N_10696);
nor U10885 (N_10885,N_10740,N_10722);
or U10886 (N_10886,N_10670,N_10693);
nor U10887 (N_10887,N_10778,N_10785);
nand U10888 (N_10888,N_10787,N_10795);
or U10889 (N_10889,N_10730,N_10757);
and U10890 (N_10890,N_10715,N_10634);
xor U10891 (N_10891,N_10697,N_10793);
and U10892 (N_10892,N_10770,N_10725);
and U10893 (N_10893,N_10701,N_10624);
or U10894 (N_10894,N_10658,N_10766);
nand U10895 (N_10895,N_10756,N_10629);
xnor U10896 (N_10896,N_10783,N_10750);
nor U10897 (N_10897,N_10684,N_10651);
nand U10898 (N_10898,N_10677,N_10797);
and U10899 (N_10899,N_10638,N_10610);
and U10900 (N_10900,N_10655,N_10617);
or U10901 (N_10901,N_10780,N_10696);
nand U10902 (N_10902,N_10652,N_10654);
and U10903 (N_10903,N_10600,N_10793);
and U10904 (N_10904,N_10666,N_10605);
nor U10905 (N_10905,N_10744,N_10717);
nand U10906 (N_10906,N_10666,N_10640);
nor U10907 (N_10907,N_10742,N_10728);
xor U10908 (N_10908,N_10638,N_10776);
and U10909 (N_10909,N_10686,N_10605);
xor U10910 (N_10910,N_10678,N_10618);
nor U10911 (N_10911,N_10677,N_10766);
nor U10912 (N_10912,N_10681,N_10717);
nor U10913 (N_10913,N_10630,N_10620);
or U10914 (N_10914,N_10726,N_10739);
and U10915 (N_10915,N_10605,N_10770);
and U10916 (N_10916,N_10685,N_10743);
nand U10917 (N_10917,N_10766,N_10725);
and U10918 (N_10918,N_10670,N_10700);
xor U10919 (N_10919,N_10761,N_10707);
xnor U10920 (N_10920,N_10717,N_10723);
and U10921 (N_10921,N_10600,N_10733);
and U10922 (N_10922,N_10663,N_10613);
nor U10923 (N_10923,N_10611,N_10763);
xnor U10924 (N_10924,N_10680,N_10770);
nor U10925 (N_10925,N_10705,N_10768);
nand U10926 (N_10926,N_10601,N_10708);
nor U10927 (N_10927,N_10757,N_10729);
nand U10928 (N_10928,N_10627,N_10739);
nor U10929 (N_10929,N_10666,N_10636);
nand U10930 (N_10930,N_10623,N_10782);
nand U10931 (N_10931,N_10632,N_10746);
and U10932 (N_10932,N_10679,N_10790);
nand U10933 (N_10933,N_10704,N_10603);
or U10934 (N_10934,N_10620,N_10644);
nor U10935 (N_10935,N_10635,N_10728);
and U10936 (N_10936,N_10707,N_10738);
nand U10937 (N_10937,N_10762,N_10707);
and U10938 (N_10938,N_10770,N_10663);
nor U10939 (N_10939,N_10605,N_10732);
or U10940 (N_10940,N_10636,N_10612);
nor U10941 (N_10941,N_10657,N_10649);
xnor U10942 (N_10942,N_10654,N_10740);
nand U10943 (N_10943,N_10764,N_10668);
nand U10944 (N_10944,N_10691,N_10610);
and U10945 (N_10945,N_10627,N_10654);
or U10946 (N_10946,N_10719,N_10627);
nor U10947 (N_10947,N_10657,N_10629);
nand U10948 (N_10948,N_10676,N_10731);
nand U10949 (N_10949,N_10781,N_10602);
xnor U10950 (N_10950,N_10680,N_10656);
nand U10951 (N_10951,N_10614,N_10771);
xnor U10952 (N_10952,N_10787,N_10727);
xor U10953 (N_10953,N_10708,N_10674);
nand U10954 (N_10954,N_10686,N_10792);
or U10955 (N_10955,N_10625,N_10747);
nor U10956 (N_10956,N_10612,N_10639);
nand U10957 (N_10957,N_10658,N_10684);
nor U10958 (N_10958,N_10715,N_10712);
or U10959 (N_10959,N_10786,N_10625);
xnor U10960 (N_10960,N_10692,N_10643);
and U10961 (N_10961,N_10710,N_10716);
or U10962 (N_10962,N_10613,N_10614);
or U10963 (N_10963,N_10707,N_10706);
nand U10964 (N_10964,N_10651,N_10718);
or U10965 (N_10965,N_10678,N_10745);
nand U10966 (N_10966,N_10634,N_10615);
and U10967 (N_10967,N_10777,N_10703);
nand U10968 (N_10968,N_10636,N_10761);
nor U10969 (N_10969,N_10735,N_10661);
or U10970 (N_10970,N_10625,N_10618);
xor U10971 (N_10971,N_10667,N_10630);
or U10972 (N_10972,N_10665,N_10625);
nor U10973 (N_10973,N_10685,N_10716);
nand U10974 (N_10974,N_10639,N_10782);
or U10975 (N_10975,N_10707,N_10741);
or U10976 (N_10976,N_10686,N_10633);
nand U10977 (N_10977,N_10728,N_10750);
nor U10978 (N_10978,N_10655,N_10774);
or U10979 (N_10979,N_10653,N_10754);
nor U10980 (N_10980,N_10724,N_10619);
nand U10981 (N_10981,N_10695,N_10639);
and U10982 (N_10982,N_10799,N_10653);
nor U10983 (N_10983,N_10731,N_10604);
and U10984 (N_10984,N_10678,N_10786);
xnor U10985 (N_10985,N_10764,N_10652);
xor U10986 (N_10986,N_10656,N_10671);
nor U10987 (N_10987,N_10636,N_10627);
or U10988 (N_10988,N_10612,N_10604);
and U10989 (N_10989,N_10619,N_10643);
nor U10990 (N_10990,N_10629,N_10725);
xor U10991 (N_10991,N_10671,N_10774);
nand U10992 (N_10992,N_10634,N_10759);
and U10993 (N_10993,N_10665,N_10658);
nand U10994 (N_10994,N_10740,N_10697);
nand U10995 (N_10995,N_10777,N_10604);
or U10996 (N_10996,N_10762,N_10795);
nand U10997 (N_10997,N_10713,N_10789);
or U10998 (N_10998,N_10617,N_10747);
xor U10999 (N_10999,N_10608,N_10626);
nand U11000 (N_11000,N_10970,N_10941);
or U11001 (N_11001,N_10962,N_10838);
nor U11002 (N_11002,N_10967,N_10948);
or U11003 (N_11003,N_10852,N_10854);
and U11004 (N_11004,N_10861,N_10890);
or U11005 (N_11005,N_10942,N_10969);
xor U11006 (N_11006,N_10824,N_10930);
or U11007 (N_11007,N_10937,N_10829);
and U11008 (N_11008,N_10943,N_10905);
or U11009 (N_11009,N_10806,N_10827);
or U11010 (N_11010,N_10816,N_10856);
xnor U11011 (N_11011,N_10831,N_10834);
xnor U11012 (N_11012,N_10933,N_10884);
nor U11013 (N_11013,N_10862,N_10810);
or U11014 (N_11014,N_10876,N_10888);
nor U11015 (N_11015,N_10853,N_10977);
nor U11016 (N_11016,N_10811,N_10936);
nor U11017 (N_11017,N_10920,N_10898);
xnor U11018 (N_11018,N_10842,N_10953);
and U11019 (N_11019,N_10973,N_10830);
and U11020 (N_11020,N_10966,N_10981);
nor U11021 (N_11021,N_10817,N_10839);
xor U11022 (N_11022,N_10859,N_10877);
or U11023 (N_11023,N_10880,N_10947);
nor U11024 (N_11024,N_10932,N_10922);
or U11025 (N_11025,N_10843,N_10971);
xnor U11026 (N_11026,N_10935,N_10872);
nor U11027 (N_11027,N_10934,N_10865);
nand U11028 (N_11028,N_10945,N_10957);
nor U11029 (N_11029,N_10908,N_10886);
xor U11030 (N_11030,N_10846,N_10864);
xor U11031 (N_11031,N_10983,N_10978);
nor U11032 (N_11032,N_10878,N_10902);
and U11033 (N_11033,N_10927,N_10895);
xnor U11034 (N_11034,N_10801,N_10982);
xor U11035 (N_11035,N_10916,N_10955);
and U11036 (N_11036,N_10950,N_10844);
or U11037 (N_11037,N_10921,N_10813);
nand U11038 (N_11038,N_10826,N_10959);
or U11039 (N_11039,N_10960,N_10989);
xor U11040 (N_11040,N_10938,N_10889);
or U11041 (N_11041,N_10995,N_10993);
nand U11042 (N_11042,N_10828,N_10923);
or U11043 (N_11043,N_10840,N_10911);
or U11044 (N_11044,N_10976,N_10985);
nand U11045 (N_11045,N_10803,N_10894);
nand U11046 (N_11046,N_10928,N_10956);
and U11047 (N_11047,N_10814,N_10847);
nor U11048 (N_11048,N_10899,N_10949);
or U11049 (N_11049,N_10807,N_10964);
or U11050 (N_11050,N_10837,N_10891);
nand U11051 (N_11051,N_10849,N_10907);
nor U11052 (N_11052,N_10841,N_10900);
nor U11053 (N_11053,N_10802,N_10999);
and U11054 (N_11054,N_10820,N_10909);
nor U11055 (N_11055,N_10897,N_10926);
xor U11056 (N_11056,N_10952,N_10991);
or U11057 (N_11057,N_10987,N_10879);
and U11058 (N_11058,N_10883,N_10906);
and U11059 (N_11059,N_10925,N_10954);
nor U11060 (N_11060,N_10994,N_10965);
nor U11061 (N_11061,N_10997,N_10910);
and U11062 (N_11062,N_10975,N_10836);
nand U11063 (N_11063,N_10809,N_10868);
or U11064 (N_11064,N_10961,N_10940);
nor U11065 (N_11065,N_10992,N_10887);
and U11066 (N_11066,N_10924,N_10867);
xnor U11067 (N_11067,N_10804,N_10805);
nor U11068 (N_11068,N_10821,N_10986);
xor U11069 (N_11069,N_10819,N_10939);
nand U11070 (N_11070,N_10896,N_10903);
nor U11071 (N_11071,N_10800,N_10901);
and U11072 (N_11072,N_10913,N_10855);
xor U11073 (N_11073,N_10863,N_10963);
nor U11074 (N_11074,N_10951,N_10968);
or U11075 (N_11075,N_10869,N_10984);
or U11076 (N_11076,N_10866,N_10851);
nand U11077 (N_11077,N_10873,N_10980);
xor U11078 (N_11078,N_10929,N_10919);
xor U11079 (N_11079,N_10835,N_10818);
nor U11080 (N_11080,N_10946,N_10825);
or U11081 (N_11081,N_10988,N_10979);
or U11082 (N_11082,N_10918,N_10931);
and U11083 (N_11083,N_10870,N_10904);
nor U11084 (N_11084,N_10882,N_10857);
or U11085 (N_11085,N_10990,N_10914);
nor U11086 (N_11086,N_10845,N_10881);
xnor U11087 (N_11087,N_10848,N_10885);
or U11088 (N_11088,N_10850,N_10915);
and U11089 (N_11089,N_10808,N_10822);
and U11090 (N_11090,N_10972,N_10892);
nand U11091 (N_11091,N_10833,N_10958);
and U11092 (N_11092,N_10996,N_10871);
nor U11093 (N_11093,N_10823,N_10875);
xnor U11094 (N_11094,N_10858,N_10812);
and U11095 (N_11095,N_10912,N_10998);
nand U11096 (N_11096,N_10893,N_10917);
nand U11097 (N_11097,N_10815,N_10874);
nand U11098 (N_11098,N_10974,N_10832);
or U11099 (N_11099,N_10860,N_10944);
and U11100 (N_11100,N_10813,N_10849);
nand U11101 (N_11101,N_10917,N_10882);
and U11102 (N_11102,N_10862,N_10953);
and U11103 (N_11103,N_10967,N_10963);
or U11104 (N_11104,N_10869,N_10877);
or U11105 (N_11105,N_10904,N_10830);
or U11106 (N_11106,N_10925,N_10813);
nor U11107 (N_11107,N_10871,N_10811);
xnor U11108 (N_11108,N_10972,N_10956);
nand U11109 (N_11109,N_10827,N_10879);
xnor U11110 (N_11110,N_10897,N_10959);
nor U11111 (N_11111,N_10922,N_10903);
xnor U11112 (N_11112,N_10979,N_10989);
xor U11113 (N_11113,N_10960,N_10853);
nand U11114 (N_11114,N_10802,N_10987);
and U11115 (N_11115,N_10883,N_10885);
xor U11116 (N_11116,N_10901,N_10837);
or U11117 (N_11117,N_10885,N_10805);
nor U11118 (N_11118,N_10826,N_10809);
or U11119 (N_11119,N_10917,N_10818);
or U11120 (N_11120,N_10925,N_10931);
nand U11121 (N_11121,N_10900,N_10895);
xor U11122 (N_11122,N_10948,N_10985);
nor U11123 (N_11123,N_10881,N_10933);
nand U11124 (N_11124,N_10814,N_10844);
nor U11125 (N_11125,N_10947,N_10902);
and U11126 (N_11126,N_10950,N_10866);
or U11127 (N_11127,N_10850,N_10805);
xor U11128 (N_11128,N_10904,N_10969);
nand U11129 (N_11129,N_10892,N_10881);
and U11130 (N_11130,N_10901,N_10968);
and U11131 (N_11131,N_10851,N_10838);
or U11132 (N_11132,N_10843,N_10806);
nand U11133 (N_11133,N_10892,N_10828);
nand U11134 (N_11134,N_10822,N_10866);
and U11135 (N_11135,N_10875,N_10906);
nor U11136 (N_11136,N_10800,N_10944);
or U11137 (N_11137,N_10904,N_10869);
and U11138 (N_11138,N_10813,N_10838);
nand U11139 (N_11139,N_10954,N_10801);
or U11140 (N_11140,N_10848,N_10804);
nand U11141 (N_11141,N_10865,N_10987);
xnor U11142 (N_11142,N_10985,N_10979);
nand U11143 (N_11143,N_10826,N_10940);
nor U11144 (N_11144,N_10909,N_10898);
nand U11145 (N_11145,N_10845,N_10922);
and U11146 (N_11146,N_10874,N_10868);
xor U11147 (N_11147,N_10863,N_10865);
and U11148 (N_11148,N_10834,N_10863);
nor U11149 (N_11149,N_10811,N_10938);
nand U11150 (N_11150,N_10800,N_10919);
or U11151 (N_11151,N_10882,N_10811);
or U11152 (N_11152,N_10866,N_10818);
nand U11153 (N_11153,N_10874,N_10803);
or U11154 (N_11154,N_10814,N_10979);
nand U11155 (N_11155,N_10843,N_10954);
nand U11156 (N_11156,N_10975,N_10845);
or U11157 (N_11157,N_10985,N_10810);
xor U11158 (N_11158,N_10802,N_10970);
or U11159 (N_11159,N_10898,N_10998);
or U11160 (N_11160,N_10946,N_10835);
nor U11161 (N_11161,N_10934,N_10922);
xor U11162 (N_11162,N_10883,N_10850);
nor U11163 (N_11163,N_10828,N_10925);
nor U11164 (N_11164,N_10877,N_10865);
and U11165 (N_11165,N_10896,N_10979);
and U11166 (N_11166,N_10983,N_10846);
or U11167 (N_11167,N_10820,N_10953);
nor U11168 (N_11168,N_10933,N_10800);
and U11169 (N_11169,N_10873,N_10819);
or U11170 (N_11170,N_10807,N_10922);
nand U11171 (N_11171,N_10825,N_10894);
nor U11172 (N_11172,N_10812,N_10827);
nor U11173 (N_11173,N_10805,N_10943);
nand U11174 (N_11174,N_10901,N_10882);
and U11175 (N_11175,N_10998,N_10947);
and U11176 (N_11176,N_10801,N_10823);
or U11177 (N_11177,N_10985,N_10918);
xnor U11178 (N_11178,N_10855,N_10950);
nor U11179 (N_11179,N_10984,N_10933);
xor U11180 (N_11180,N_10891,N_10816);
or U11181 (N_11181,N_10868,N_10864);
or U11182 (N_11182,N_10926,N_10932);
nand U11183 (N_11183,N_10998,N_10933);
nand U11184 (N_11184,N_10946,N_10942);
nor U11185 (N_11185,N_10910,N_10923);
or U11186 (N_11186,N_10988,N_10944);
and U11187 (N_11187,N_10909,N_10818);
nand U11188 (N_11188,N_10892,N_10920);
xor U11189 (N_11189,N_10918,N_10815);
nand U11190 (N_11190,N_10892,N_10835);
xor U11191 (N_11191,N_10802,N_10996);
nor U11192 (N_11192,N_10977,N_10868);
and U11193 (N_11193,N_10982,N_10993);
nand U11194 (N_11194,N_10857,N_10904);
and U11195 (N_11195,N_10857,N_10992);
nand U11196 (N_11196,N_10909,N_10829);
nor U11197 (N_11197,N_10853,N_10940);
xnor U11198 (N_11198,N_10887,N_10841);
xor U11199 (N_11199,N_10927,N_10996);
or U11200 (N_11200,N_11091,N_11032);
or U11201 (N_11201,N_11190,N_11176);
nand U11202 (N_11202,N_11074,N_11175);
nor U11203 (N_11203,N_11162,N_11097);
xnor U11204 (N_11204,N_11079,N_11069);
nand U11205 (N_11205,N_11094,N_11167);
nand U11206 (N_11206,N_11105,N_11178);
nand U11207 (N_11207,N_11150,N_11108);
or U11208 (N_11208,N_11125,N_11057);
or U11209 (N_11209,N_11044,N_11071);
or U11210 (N_11210,N_11081,N_11042);
xor U11211 (N_11211,N_11011,N_11188);
xnor U11212 (N_11212,N_11109,N_11124);
nand U11213 (N_11213,N_11120,N_11161);
xnor U11214 (N_11214,N_11163,N_11180);
and U11215 (N_11215,N_11145,N_11060);
and U11216 (N_11216,N_11055,N_11007);
or U11217 (N_11217,N_11054,N_11038);
nand U11218 (N_11218,N_11182,N_11164);
nand U11219 (N_11219,N_11098,N_11148);
or U11220 (N_11220,N_11174,N_11099);
nand U11221 (N_11221,N_11186,N_11039);
nor U11222 (N_11222,N_11119,N_11149);
xnor U11223 (N_11223,N_11113,N_11062);
nand U11224 (N_11224,N_11127,N_11123);
and U11225 (N_11225,N_11107,N_11040);
nor U11226 (N_11226,N_11047,N_11157);
nor U11227 (N_11227,N_11072,N_11014);
and U11228 (N_11228,N_11053,N_11192);
nor U11229 (N_11229,N_11050,N_11096);
nand U11230 (N_11230,N_11139,N_11136);
and U11231 (N_11231,N_11159,N_11179);
nor U11232 (N_11232,N_11025,N_11034);
and U11233 (N_11233,N_11002,N_11144);
nand U11234 (N_11234,N_11198,N_11048);
and U11235 (N_11235,N_11087,N_11064);
and U11236 (N_11236,N_11132,N_11137);
or U11237 (N_11237,N_11067,N_11090);
or U11238 (N_11238,N_11195,N_11005);
nor U11239 (N_11239,N_11029,N_11026);
xor U11240 (N_11240,N_11147,N_11027);
and U11241 (N_11241,N_11017,N_11130);
or U11242 (N_11242,N_11193,N_11103);
and U11243 (N_11243,N_11084,N_11111);
and U11244 (N_11244,N_11022,N_11021);
and U11245 (N_11245,N_11041,N_11122);
nor U11246 (N_11246,N_11000,N_11006);
nand U11247 (N_11247,N_11142,N_11197);
and U11248 (N_11248,N_11092,N_11165);
and U11249 (N_11249,N_11082,N_11128);
nor U11250 (N_11250,N_11115,N_11063);
nand U11251 (N_11251,N_11100,N_11169);
and U11252 (N_11252,N_11199,N_11173);
nor U11253 (N_11253,N_11073,N_11187);
nand U11254 (N_11254,N_11095,N_11101);
and U11255 (N_11255,N_11183,N_11129);
nor U11256 (N_11256,N_11152,N_11166);
or U11257 (N_11257,N_11018,N_11158);
xor U11258 (N_11258,N_11059,N_11177);
and U11259 (N_11259,N_11066,N_11083);
nor U11260 (N_11260,N_11070,N_11110);
nor U11261 (N_11261,N_11019,N_11037);
nor U11262 (N_11262,N_11168,N_11171);
nand U11263 (N_11263,N_11135,N_11146);
nor U11264 (N_11264,N_11134,N_11020);
or U11265 (N_11265,N_11104,N_11030);
nand U11266 (N_11266,N_11024,N_11191);
or U11267 (N_11267,N_11093,N_11194);
xnor U11268 (N_11268,N_11185,N_11051);
or U11269 (N_11269,N_11046,N_11156);
nand U11270 (N_11270,N_11172,N_11118);
or U11271 (N_11271,N_11075,N_11016);
nand U11272 (N_11272,N_11009,N_11045);
nor U11273 (N_11273,N_11056,N_11078);
and U11274 (N_11274,N_11033,N_11116);
and U11275 (N_11275,N_11023,N_11114);
nor U11276 (N_11276,N_11196,N_11102);
or U11277 (N_11277,N_11155,N_11138);
xnor U11278 (N_11278,N_11061,N_11031);
xnor U11279 (N_11279,N_11181,N_11131);
xnor U11280 (N_11280,N_11160,N_11043);
xnor U11281 (N_11281,N_11049,N_11133);
nand U11282 (N_11282,N_11151,N_11012);
and U11283 (N_11283,N_11028,N_11010);
and U11284 (N_11284,N_11126,N_11003);
or U11285 (N_11285,N_11008,N_11184);
or U11286 (N_11286,N_11068,N_11141);
xnor U11287 (N_11287,N_11154,N_11088);
nand U11288 (N_11288,N_11058,N_11170);
nand U11289 (N_11289,N_11153,N_11077);
nand U11290 (N_11290,N_11065,N_11112);
or U11291 (N_11291,N_11080,N_11089);
nor U11292 (N_11292,N_11036,N_11189);
nand U11293 (N_11293,N_11004,N_11140);
xnor U11294 (N_11294,N_11143,N_11086);
nand U11295 (N_11295,N_11106,N_11013);
and U11296 (N_11296,N_11015,N_11001);
or U11297 (N_11297,N_11052,N_11121);
nor U11298 (N_11298,N_11117,N_11076);
xnor U11299 (N_11299,N_11035,N_11085);
and U11300 (N_11300,N_11000,N_11134);
or U11301 (N_11301,N_11035,N_11075);
xnor U11302 (N_11302,N_11001,N_11024);
xnor U11303 (N_11303,N_11039,N_11050);
nor U11304 (N_11304,N_11196,N_11077);
nand U11305 (N_11305,N_11067,N_11011);
nor U11306 (N_11306,N_11089,N_11086);
xor U11307 (N_11307,N_11044,N_11047);
xor U11308 (N_11308,N_11181,N_11154);
or U11309 (N_11309,N_11175,N_11057);
nor U11310 (N_11310,N_11079,N_11192);
or U11311 (N_11311,N_11079,N_11190);
xnor U11312 (N_11312,N_11105,N_11151);
nor U11313 (N_11313,N_11084,N_11188);
nand U11314 (N_11314,N_11065,N_11111);
nor U11315 (N_11315,N_11136,N_11128);
and U11316 (N_11316,N_11030,N_11159);
or U11317 (N_11317,N_11166,N_11191);
or U11318 (N_11318,N_11063,N_11127);
nor U11319 (N_11319,N_11024,N_11184);
nand U11320 (N_11320,N_11018,N_11183);
xor U11321 (N_11321,N_11148,N_11032);
xnor U11322 (N_11322,N_11197,N_11022);
and U11323 (N_11323,N_11112,N_11194);
xor U11324 (N_11324,N_11012,N_11173);
nor U11325 (N_11325,N_11098,N_11011);
xnor U11326 (N_11326,N_11120,N_11007);
and U11327 (N_11327,N_11105,N_11108);
and U11328 (N_11328,N_11086,N_11099);
nor U11329 (N_11329,N_11113,N_11184);
xnor U11330 (N_11330,N_11070,N_11156);
or U11331 (N_11331,N_11053,N_11185);
xnor U11332 (N_11332,N_11013,N_11086);
and U11333 (N_11333,N_11150,N_11001);
and U11334 (N_11334,N_11048,N_11070);
nand U11335 (N_11335,N_11137,N_11192);
nor U11336 (N_11336,N_11001,N_11083);
nand U11337 (N_11337,N_11109,N_11162);
xor U11338 (N_11338,N_11085,N_11032);
or U11339 (N_11339,N_11140,N_11057);
xor U11340 (N_11340,N_11116,N_11122);
and U11341 (N_11341,N_11018,N_11169);
nand U11342 (N_11342,N_11172,N_11017);
xor U11343 (N_11343,N_11139,N_11074);
xor U11344 (N_11344,N_11002,N_11153);
nor U11345 (N_11345,N_11041,N_11049);
nand U11346 (N_11346,N_11181,N_11060);
nor U11347 (N_11347,N_11072,N_11070);
xor U11348 (N_11348,N_11197,N_11143);
or U11349 (N_11349,N_11042,N_11000);
nand U11350 (N_11350,N_11121,N_11045);
xnor U11351 (N_11351,N_11089,N_11176);
or U11352 (N_11352,N_11163,N_11197);
or U11353 (N_11353,N_11074,N_11005);
nor U11354 (N_11354,N_11127,N_11125);
or U11355 (N_11355,N_11191,N_11129);
nand U11356 (N_11356,N_11192,N_11040);
xor U11357 (N_11357,N_11127,N_11118);
xnor U11358 (N_11358,N_11036,N_11155);
xor U11359 (N_11359,N_11137,N_11032);
nor U11360 (N_11360,N_11138,N_11164);
nand U11361 (N_11361,N_11092,N_11061);
nor U11362 (N_11362,N_11013,N_11076);
xnor U11363 (N_11363,N_11033,N_11010);
nand U11364 (N_11364,N_11067,N_11100);
and U11365 (N_11365,N_11010,N_11072);
xnor U11366 (N_11366,N_11182,N_11054);
and U11367 (N_11367,N_11016,N_11181);
xnor U11368 (N_11368,N_11167,N_11149);
xnor U11369 (N_11369,N_11162,N_11196);
xor U11370 (N_11370,N_11071,N_11190);
xor U11371 (N_11371,N_11186,N_11081);
nor U11372 (N_11372,N_11031,N_11132);
xnor U11373 (N_11373,N_11019,N_11174);
nand U11374 (N_11374,N_11086,N_11124);
or U11375 (N_11375,N_11006,N_11065);
nand U11376 (N_11376,N_11033,N_11094);
and U11377 (N_11377,N_11169,N_11099);
nand U11378 (N_11378,N_11020,N_11136);
nor U11379 (N_11379,N_11126,N_11194);
nor U11380 (N_11380,N_11029,N_11174);
nor U11381 (N_11381,N_11196,N_11029);
nand U11382 (N_11382,N_11071,N_11002);
xnor U11383 (N_11383,N_11034,N_11181);
or U11384 (N_11384,N_11167,N_11029);
and U11385 (N_11385,N_11000,N_11113);
xnor U11386 (N_11386,N_11067,N_11184);
and U11387 (N_11387,N_11084,N_11036);
and U11388 (N_11388,N_11171,N_11120);
or U11389 (N_11389,N_11020,N_11192);
nor U11390 (N_11390,N_11015,N_11038);
nor U11391 (N_11391,N_11144,N_11079);
nand U11392 (N_11392,N_11167,N_11023);
or U11393 (N_11393,N_11084,N_11157);
xor U11394 (N_11394,N_11030,N_11162);
xnor U11395 (N_11395,N_11032,N_11000);
or U11396 (N_11396,N_11016,N_11119);
and U11397 (N_11397,N_11065,N_11074);
and U11398 (N_11398,N_11012,N_11031);
xor U11399 (N_11399,N_11089,N_11053);
or U11400 (N_11400,N_11305,N_11353);
nand U11401 (N_11401,N_11396,N_11312);
nand U11402 (N_11402,N_11362,N_11215);
nand U11403 (N_11403,N_11356,N_11339);
xnor U11404 (N_11404,N_11242,N_11207);
and U11405 (N_11405,N_11217,N_11255);
nor U11406 (N_11406,N_11322,N_11277);
and U11407 (N_11407,N_11289,N_11274);
xor U11408 (N_11408,N_11311,N_11320);
xnor U11409 (N_11409,N_11222,N_11397);
nor U11410 (N_11410,N_11286,N_11296);
nor U11411 (N_11411,N_11326,N_11381);
xor U11412 (N_11412,N_11298,N_11342);
nor U11413 (N_11413,N_11398,N_11212);
nand U11414 (N_11414,N_11279,N_11389);
or U11415 (N_11415,N_11351,N_11291);
xnor U11416 (N_11416,N_11294,N_11335);
and U11417 (N_11417,N_11372,N_11243);
or U11418 (N_11418,N_11204,N_11273);
nor U11419 (N_11419,N_11329,N_11369);
nand U11420 (N_11420,N_11364,N_11210);
or U11421 (N_11421,N_11355,N_11350);
and U11422 (N_11422,N_11292,N_11239);
and U11423 (N_11423,N_11205,N_11328);
nand U11424 (N_11424,N_11394,N_11363);
or U11425 (N_11425,N_11283,N_11325);
nand U11426 (N_11426,N_11282,N_11270);
nand U11427 (N_11427,N_11321,N_11391);
nor U11428 (N_11428,N_11280,N_11309);
or U11429 (N_11429,N_11373,N_11330);
nand U11430 (N_11430,N_11357,N_11229);
nor U11431 (N_11431,N_11262,N_11208);
or U11432 (N_11432,N_11201,N_11348);
or U11433 (N_11433,N_11234,N_11246);
and U11434 (N_11434,N_11310,N_11290);
or U11435 (N_11435,N_11316,N_11346);
or U11436 (N_11436,N_11341,N_11386);
xnor U11437 (N_11437,N_11267,N_11380);
or U11438 (N_11438,N_11203,N_11303);
or U11439 (N_11439,N_11314,N_11354);
xor U11440 (N_11440,N_11333,N_11248);
nand U11441 (N_11441,N_11214,N_11327);
nand U11442 (N_11442,N_11281,N_11253);
or U11443 (N_11443,N_11265,N_11340);
or U11444 (N_11444,N_11206,N_11241);
nor U11445 (N_11445,N_11226,N_11285);
nand U11446 (N_11446,N_11221,N_11258);
nor U11447 (N_11447,N_11224,N_11359);
and U11448 (N_11448,N_11399,N_11278);
nand U11449 (N_11449,N_11261,N_11323);
nand U11450 (N_11450,N_11297,N_11284);
nand U11451 (N_11451,N_11266,N_11331);
nand U11452 (N_11452,N_11361,N_11382);
nand U11453 (N_11453,N_11352,N_11299);
nand U11454 (N_11454,N_11384,N_11240);
or U11455 (N_11455,N_11338,N_11378);
nor U11456 (N_11456,N_11371,N_11318);
nand U11457 (N_11457,N_11379,N_11268);
xor U11458 (N_11458,N_11319,N_11202);
and U11459 (N_11459,N_11313,N_11231);
xor U11460 (N_11460,N_11383,N_11332);
nor U11461 (N_11461,N_11232,N_11347);
or U11462 (N_11462,N_11300,N_11235);
nand U11463 (N_11463,N_11307,N_11360);
xnor U11464 (N_11464,N_11392,N_11302);
or U11465 (N_11465,N_11260,N_11367);
nor U11466 (N_11466,N_11276,N_11375);
nor U11467 (N_11467,N_11293,N_11275);
xor U11468 (N_11468,N_11385,N_11209);
nand U11469 (N_11469,N_11349,N_11220);
and U11470 (N_11470,N_11263,N_11388);
nor U11471 (N_11471,N_11344,N_11218);
nor U11472 (N_11472,N_11393,N_11358);
nor U11473 (N_11473,N_11271,N_11236);
xor U11474 (N_11474,N_11254,N_11237);
and U11475 (N_11475,N_11259,N_11230);
xnor U11476 (N_11476,N_11387,N_11317);
and U11477 (N_11477,N_11249,N_11244);
nor U11478 (N_11478,N_11272,N_11223);
nand U11479 (N_11479,N_11227,N_11336);
nand U11480 (N_11480,N_11213,N_11315);
xor U11481 (N_11481,N_11365,N_11264);
xnor U11482 (N_11482,N_11301,N_11245);
nand U11483 (N_11483,N_11343,N_11233);
xnor U11484 (N_11484,N_11252,N_11377);
and U11485 (N_11485,N_11256,N_11366);
nand U11486 (N_11486,N_11304,N_11334);
nand U11487 (N_11487,N_11395,N_11306);
xor U11488 (N_11488,N_11250,N_11238);
or U11489 (N_11489,N_11228,N_11251);
nand U11490 (N_11490,N_11200,N_11216);
xor U11491 (N_11491,N_11368,N_11288);
xnor U11492 (N_11492,N_11211,N_11376);
and U11493 (N_11493,N_11219,N_11257);
and U11494 (N_11494,N_11324,N_11308);
nand U11495 (N_11495,N_11269,N_11295);
nor U11496 (N_11496,N_11390,N_11337);
or U11497 (N_11497,N_11370,N_11345);
nand U11498 (N_11498,N_11247,N_11374);
and U11499 (N_11499,N_11225,N_11287);
nor U11500 (N_11500,N_11249,N_11297);
nor U11501 (N_11501,N_11248,N_11330);
or U11502 (N_11502,N_11297,N_11393);
nor U11503 (N_11503,N_11362,N_11231);
xor U11504 (N_11504,N_11370,N_11210);
nand U11505 (N_11505,N_11319,N_11399);
and U11506 (N_11506,N_11210,N_11205);
or U11507 (N_11507,N_11300,N_11334);
xor U11508 (N_11508,N_11362,N_11361);
xnor U11509 (N_11509,N_11284,N_11310);
nand U11510 (N_11510,N_11389,N_11208);
nand U11511 (N_11511,N_11256,N_11370);
and U11512 (N_11512,N_11250,N_11372);
or U11513 (N_11513,N_11380,N_11207);
nor U11514 (N_11514,N_11310,N_11389);
nor U11515 (N_11515,N_11360,N_11346);
or U11516 (N_11516,N_11220,N_11348);
or U11517 (N_11517,N_11313,N_11290);
xor U11518 (N_11518,N_11358,N_11248);
nor U11519 (N_11519,N_11205,N_11237);
or U11520 (N_11520,N_11314,N_11342);
xor U11521 (N_11521,N_11254,N_11279);
and U11522 (N_11522,N_11306,N_11310);
nor U11523 (N_11523,N_11308,N_11249);
and U11524 (N_11524,N_11387,N_11283);
xor U11525 (N_11525,N_11387,N_11200);
and U11526 (N_11526,N_11334,N_11243);
xnor U11527 (N_11527,N_11352,N_11291);
xnor U11528 (N_11528,N_11292,N_11351);
and U11529 (N_11529,N_11291,N_11325);
and U11530 (N_11530,N_11354,N_11275);
and U11531 (N_11531,N_11262,N_11281);
xor U11532 (N_11532,N_11278,N_11364);
or U11533 (N_11533,N_11387,N_11388);
or U11534 (N_11534,N_11269,N_11394);
xnor U11535 (N_11535,N_11347,N_11340);
nor U11536 (N_11536,N_11311,N_11238);
nor U11537 (N_11537,N_11271,N_11334);
nand U11538 (N_11538,N_11308,N_11326);
and U11539 (N_11539,N_11204,N_11365);
and U11540 (N_11540,N_11311,N_11284);
and U11541 (N_11541,N_11296,N_11232);
or U11542 (N_11542,N_11259,N_11374);
nand U11543 (N_11543,N_11383,N_11251);
and U11544 (N_11544,N_11313,N_11228);
xnor U11545 (N_11545,N_11344,N_11299);
nand U11546 (N_11546,N_11270,N_11257);
and U11547 (N_11547,N_11377,N_11353);
nor U11548 (N_11548,N_11379,N_11270);
nor U11549 (N_11549,N_11394,N_11217);
xnor U11550 (N_11550,N_11365,N_11362);
and U11551 (N_11551,N_11348,N_11362);
or U11552 (N_11552,N_11366,N_11314);
nor U11553 (N_11553,N_11242,N_11225);
or U11554 (N_11554,N_11388,N_11213);
nor U11555 (N_11555,N_11209,N_11361);
or U11556 (N_11556,N_11322,N_11268);
nor U11557 (N_11557,N_11332,N_11328);
and U11558 (N_11558,N_11255,N_11266);
or U11559 (N_11559,N_11317,N_11346);
nand U11560 (N_11560,N_11351,N_11388);
or U11561 (N_11561,N_11266,N_11222);
xnor U11562 (N_11562,N_11352,N_11209);
xor U11563 (N_11563,N_11304,N_11302);
and U11564 (N_11564,N_11391,N_11384);
nand U11565 (N_11565,N_11300,N_11290);
or U11566 (N_11566,N_11344,N_11241);
nor U11567 (N_11567,N_11232,N_11307);
or U11568 (N_11568,N_11275,N_11389);
nor U11569 (N_11569,N_11282,N_11384);
xnor U11570 (N_11570,N_11282,N_11264);
or U11571 (N_11571,N_11394,N_11308);
or U11572 (N_11572,N_11203,N_11244);
and U11573 (N_11573,N_11211,N_11251);
and U11574 (N_11574,N_11398,N_11281);
nand U11575 (N_11575,N_11370,N_11331);
or U11576 (N_11576,N_11275,N_11217);
nand U11577 (N_11577,N_11315,N_11289);
nor U11578 (N_11578,N_11272,N_11386);
or U11579 (N_11579,N_11374,N_11341);
or U11580 (N_11580,N_11318,N_11219);
xnor U11581 (N_11581,N_11347,N_11318);
xnor U11582 (N_11582,N_11378,N_11296);
or U11583 (N_11583,N_11257,N_11205);
nand U11584 (N_11584,N_11306,N_11328);
nor U11585 (N_11585,N_11397,N_11286);
nor U11586 (N_11586,N_11275,N_11211);
and U11587 (N_11587,N_11224,N_11219);
or U11588 (N_11588,N_11271,N_11340);
and U11589 (N_11589,N_11207,N_11241);
nand U11590 (N_11590,N_11280,N_11217);
nor U11591 (N_11591,N_11238,N_11361);
xor U11592 (N_11592,N_11319,N_11318);
nor U11593 (N_11593,N_11245,N_11240);
xor U11594 (N_11594,N_11238,N_11387);
or U11595 (N_11595,N_11292,N_11300);
nor U11596 (N_11596,N_11235,N_11291);
nand U11597 (N_11597,N_11247,N_11361);
or U11598 (N_11598,N_11286,N_11284);
nand U11599 (N_11599,N_11249,N_11215);
nand U11600 (N_11600,N_11466,N_11522);
and U11601 (N_11601,N_11594,N_11531);
nor U11602 (N_11602,N_11517,N_11566);
nand U11603 (N_11603,N_11568,N_11533);
or U11604 (N_11604,N_11450,N_11470);
xor U11605 (N_11605,N_11580,N_11598);
nor U11606 (N_11606,N_11570,N_11595);
nand U11607 (N_11607,N_11519,N_11436);
nand U11608 (N_11608,N_11500,N_11549);
nand U11609 (N_11609,N_11554,N_11557);
and U11610 (N_11610,N_11441,N_11563);
and U11611 (N_11611,N_11488,N_11422);
xnor U11612 (N_11612,N_11419,N_11497);
or U11613 (N_11613,N_11507,N_11477);
nor U11614 (N_11614,N_11532,N_11428);
xnor U11615 (N_11615,N_11453,N_11457);
nor U11616 (N_11616,N_11416,N_11429);
nor U11617 (N_11617,N_11433,N_11505);
xor U11618 (N_11618,N_11430,N_11565);
nor U11619 (N_11619,N_11499,N_11415);
or U11620 (N_11620,N_11410,N_11431);
xor U11621 (N_11621,N_11486,N_11432);
or U11622 (N_11622,N_11485,N_11562);
nand U11623 (N_11623,N_11577,N_11574);
or U11624 (N_11624,N_11455,N_11472);
xor U11625 (N_11625,N_11541,N_11508);
nand U11626 (N_11626,N_11449,N_11534);
nand U11627 (N_11627,N_11439,N_11529);
nand U11628 (N_11628,N_11530,N_11469);
xnor U11629 (N_11629,N_11573,N_11590);
nand U11630 (N_11630,N_11586,N_11403);
nand U11631 (N_11631,N_11588,N_11451);
and U11632 (N_11632,N_11553,N_11467);
nor U11633 (N_11633,N_11448,N_11401);
or U11634 (N_11634,N_11560,N_11561);
and U11635 (N_11635,N_11512,N_11518);
nor U11636 (N_11636,N_11458,N_11504);
nand U11637 (N_11637,N_11539,N_11475);
xnor U11638 (N_11638,N_11482,N_11538);
xor U11639 (N_11639,N_11426,N_11423);
or U11640 (N_11640,N_11589,N_11552);
and U11641 (N_11641,N_11597,N_11537);
and U11642 (N_11642,N_11555,N_11564);
or U11643 (N_11643,N_11514,N_11582);
or U11644 (N_11644,N_11578,N_11461);
nor U11645 (N_11645,N_11459,N_11592);
and U11646 (N_11646,N_11446,N_11525);
xor U11647 (N_11647,N_11526,N_11591);
nand U11648 (N_11648,N_11465,N_11440);
nand U11649 (N_11649,N_11407,N_11575);
nand U11650 (N_11650,N_11442,N_11593);
or U11651 (N_11651,N_11413,N_11583);
nand U11652 (N_11652,N_11543,N_11524);
xnor U11653 (N_11653,N_11444,N_11494);
and U11654 (N_11654,N_11420,N_11464);
nor U11655 (N_11655,N_11409,N_11434);
and U11656 (N_11656,N_11418,N_11468);
nor U11657 (N_11657,N_11547,N_11490);
xnor U11658 (N_11658,N_11585,N_11493);
nor U11659 (N_11659,N_11536,N_11513);
nor U11660 (N_11660,N_11527,N_11454);
xor U11661 (N_11661,N_11491,N_11404);
nor U11662 (N_11662,N_11509,N_11559);
xnor U11663 (N_11663,N_11437,N_11460);
nand U11664 (N_11664,N_11587,N_11596);
xnor U11665 (N_11665,N_11548,N_11584);
and U11666 (N_11666,N_11481,N_11498);
nand U11667 (N_11667,N_11546,N_11506);
and U11668 (N_11668,N_11480,N_11528);
xor U11669 (N_11669,N_11571,N_11540);
nand U11670 (N_11670,N_11414,N_11479);
nor U11671 (N_11671,N_11545,N_11427);
xnor U11672 (N_11672,N_11405,N_11569);
and U11673 (N_11673,N_11447,N_11576);
and U11674 (N_11674,N_11599,N_11474);
or U11675 (N_11675,N_11402,N_11516);
or U11676 (N_11676,N_11424,N_11425);
and U11677 (N_11677,N_11558,N_11544);
and U11678 (N_11678,N_11462,N_11572);
nor U11679 (N_11679,N_11535,N_11408);
nand U11680 (N_11680,N_11471,N_11556);
or U11681 (N_11681,N_11503,N_11581);
nand U11682 (N_11682,N_11452,N_11551);
or U11683 (N_11683,N_11521,N_11445);
nand U11684 (N_11684,N_11443,N_11484);
or U11685 (N_11685,N_11412,N_11483);
nor U11686 (N_11686,N_11456,N_11542);
and U11687 (N_11687,N_11502,N_11515);
xnor U11688 (N_11688,N_11523,N_11496);
or U11689 (N_11689,N_11579,N_11438);
nand U11690 (N_11690,N_11476,N_11435);
nor U11691 (N_11691,N_11489,N_11473);
xnor U11692 (N_11692,N_11510,N_11550);
nor U11693 (N_11693,N_11487,N_11520);
nand U11694 (N_11694,N_11492,N_11400);
and U11695 (N_11695,N_11417,N_11463);
and U11696 (N_11696,N_11511,N_11501);
and U11697 (N_11697,N_11567,N_11411);
and U11698 (N_11698,N_11406,N_11421);
xnor U11699 (N_11699,N_11478,N_11495);
or U11700 (N_11700,N_11538,N_11575);
or U11701 (N_11701,N_11570,N_11517);
nor U11702 (N_11702,N_11418,N_11415);
or U11703 (N_11703,N_11488,N_11410);
and U11704 (N_11704,N_11541,N_11466);
nand U11705 (N_11705,N_11581,N_11542);
nand U11706 (N_11706,N_11561,N_11411);
nand U11707 (N_11707,N_11552,N_11511);
nand U11708 (N_11708,N_11436,N_11506);
nor U11709 (N_11709,N_11444,N_11520);
or U11710 (N_11710,N_11453,N_11576);
nor U11711 (N_11711,N_11479,N_11400);
nand U11712 (N_11712,N_11519,N_11576);
or U11713 (N_11713,N_11546,N_11437);
nand U11714 (N_11714,N_11564,N_11569);
xor U11715 (N_11715,N_11461,N_11588);
or U11716 (N_11716,N_11556,N_11465);
xnor U11717 (N_11717,N_11558,N_11527);
nor U11718 (N_11718,N_11521,N_11587);
nor U11719 (N_11719,N_11586,N_11425);
nand U11720 (N_11720,N_11548,N_11581);
nand U11721 (N_11721,N_11434,N_11478);
or U11722 (N_11722,N_11540,N_11487);
or U11723 (N_11723,N_11499,N_11443);
and U11724 (N_11724,N_11428,N_11424);
xor U11725 (N_11725,N_11498,N_11504);
nor U11726 (N_11726,N_11524,N_11458);
nand U11727 (N_11727,N_11402,N_11526);
and U11728 (N_11728,N_11548,N_11473);
nor U11729 (N_11729,N_11418,N_11528);
or U11730 (N_11730,N_11538,N_11543);
xor U11731 (N_11731,N_11441,N_11410);
and U11732 (N_11732,N_11595,N_11495);
xnor U11733 (N_11733,N_11401,N_11569);
or U11734 (N_11734,N_11411,N_11406);
or U11735 (N_11735,N_11506,N_11421);
and U11736 (N_11736,N_11584,N_11489);
nor U11737 (N_11737,N_11487,N_11510);
xnor U11738 (N_11738,N_11502,N_11593);
nor U11739 (N_11739,N_11484,N_11575);
xnor U11740 (N_11740,N_11498,N_11482);
nand U11741 (N_11741,N_11549,N_11522);
nand U11742 (N_11742,N_11473,N_11488);
nand U11743 (N_11743,N_11563,N_11414);
nor U11744 (N_11744,N_11575,N_11539);
xor U11745 (N_11745,N_11491,N_11524);
and U11746 (N_11746,N_11566,N_11425);
nand U11747 (N_11747,N_11534,N_11571);
and U11748 (N_11748,N_11538,N_11450);
and U11749 (N_11749,N_11419,N_11434);
nor U11750 (N_11750,N_11535,N_11548);
and U11751 (N_11751,N_11413,N_11470);
nand U11752 (N_11752,N_11424,N_11457);
xnor U11753 (N_11753,N_11453,N_11547);
xor U11754 (N_11754,N_11434,N_11422);
and U11755 (N_11755,N_11539,N_11578);
and U11756 (N_11756,N_11569,N_11414);
nor U11757 (N_11757,N_11572,N_11478);
and U11758 (N_11758,N_11470,N_11492);
xnor U11759 (N_11759,N_11422,N_11462);
nor U11760 (N_11760,N_11452,N_11504);
nand U11761 (N_11761,N_11498,N_11546);
nand U11762 (N_11762,N_11528,N_11448);
xor U11763 (N_11763,N_11502,N_11433);
and U11764 (N_11764,N_11526,N_11441);
and U11765 (N_11765,N_11450,N_11569);
and U11766 (N_11766,N_11453,N_11597);
nor U11767 (N_11767,N_11466,N_11588);
nor U11768 (N_11768,N_11433,N_11514);
nor U11769 (N_11769,N_11552,N_11575);
xor U11770 (N_11770,N_11459,N_11572);
or U11771 (N_11771,N_11531,N_11475);
or U11772 (N_11772,N_11441,N_11548);
and U11773 (N_11773,N_11555,N_11443);
nand U11774 (N_11774,N_11494,N_11567);
xnor U11775 (N_11775,N_11522,N_11505);
nor U11776 (N_11776,N_11472,N_11538);
nor U11777 (N_11777,N_11515,N_11417);
or U11778 (N_11778,N_11479,N_11578);
nand U11779 (N_11779,N_11448,N_11454);
nor U11780 (N_11780,N_11596,N_11411);
xnor U11781 (N_11781,N_11589,N_11559);
nor U11782 (N_11782,N_11502,N_11599);
xnor U11783 (N_11783,N_11576,N_11544);
nor U11784 (N_11784,N_11562,N_11431);
nand U11785 (N_11785,N_11411,N_11405);
or U11786 (N_11786,N_11450,N_11409);
nand U11787 (N_11787,N_11453,N_11508);
or U11788 (N_11788,N_11480,N_11558);
nor U11789 (N_11789,N_11530,N_11539);
nand U11790 (N_11790,N_11560,N_11431);
xnor U11791 (N_11791,N_11508,N_11439);
xnor U11792 (N_11792,N_11525,N_11560);
xnor U11793 (N_11793,N_11444,N_11593);
and U11794 (N_11794,N_11411,N_11505);
nand U11795 (N_11795,N_11586,N_11468);
nand U11796 (N_11796,N_11434,N_11463);
or U11797 (N_11797,N_11440,N_11592);
and U11798 (N_11798,N_11567,N_11584);
xnor U11799 (N_11799,N_11466,N_11510);
and U11800 (N_11800,N_11796,N_11655);
xor U11801 (N_11801,N_11619,N_11669);
nand U11802 (N_11802,N_11717,N_11701);
nand U11803 (N_11803,N_11685,N_11670);
nor U11804 (N_11804,N_11654,N_11736);
xnor U11805 (N_11805,N_11767,N_11630);
nand U11806 (N_11806,N_11709,N_11616);
nand U11807 (N_11807,N_11789,N_11686);
nor U11808 (N_11808,N_11641,N_11720);
and U11809 (N_11809,N_11768,N_11611);
nor U11810 (N_11810,N_11741,N_11639);
or U11811 (N_11811,N_11621,N_11673);
nand U11812 (N_11812,N_11704,N_11601);
xnor U11813 (N_11813,N_11700,N_11706);
nor U11814 (N_11814,N_11658,N_11638);
xnor U11815 (N_11815,N_11756,N_11609);
and U11816 (N_11816,N_11691,N_11651);
xor U11817 (N_11817,N_11645,N_11607);
nor U11818 (N_11818,N_11714,N_11681);
nand U11819 (N_11819,N_11780,N_11666);
nor U11820 (N_11820,N_11695,N_11613);
nand U11821 (N_11821,N_11683,N_11699);
xnor U11822 (N_11822,N_11760,N_11791);
nand U11823 (N_11823,N_11786,N_11677);
nor U11824 (N_11824,N_11778,N_11719);
nand U11825 (N_11825,N_11625,N_11674);
nor U11826 (N_11826,N_11637,N_11712);
nand U11827 (N_11827,N_11618,N_11742);
and U11828 (N_11828,N_11600,N_11647);
nand U11829 (N_11829,N_11676,N_11657);
nor U11830 (N_11830,N_11634,N_11765);
nand U11831 (N_11831,N_11708,N_11750);
or U11832 (N_11832,N_11711,N_11693);
nor U11833 (N_11833,N_11675,N_11610);
xnor U11834 (N_11834,N_11792,N_11660);
nand U11835 (N_11835,N_11643,N_11781);
nor U11836 (N_11836,N_11739,N_11662);
or U11837 (N_11837,N_11763,N_11602);
nand U11838 (N_11838,N_11762,N_11731);
or U11839 (N_11839,N_11776,N_11773);
nor U11840 (N_11840,N_11733,N_11748);
xnor U11841 (N_11841,N_11624,N_11653);
nand U11842 (N_11842,N_11735,N_11650);
nand U11843 (N_11843,N_11783,N_11744);
xor U11844 (N_11844,N_11629,N_11603);
nand U11845 (N_11845,N_11617,N_11764);
and U11846 (N_11846,N_11759,N_11646);
and U11847 (N_11847,N_11710,N_11705);
nor U11848 (N_11848,N_11777,N_11730);
or U11849 (N_11849,N_11687,N_11628);
or U11850 (N_11850,N_11732,N_11644);
nand U11851 (N_11851,N_11622,N_11799);
xor U11852 (N_11852,N_11740,N_11788);
or U11853 (N_11853,N_11775,N_11713);
nand U11854 (N_11854,N_11671,N_11614);
nand U11855 (N_11855,N_11604,N_11737);
or U11856 (N_11856,N_11615,N_11631);
xor U11857 (N_11857,N_11702,N_11608);
nand U11858 (N_11858,N_11724,N_11716);
nor U11859 (N_11859,N_11703,N_11769);
xnor U11860 (N_11860,N_11745,N_11652);
xor U11861 (N_11861,N_11640,N_11758);
xnor U11862 (N_11862,N_11635,N_11755);
and U11863 (N_11863,N_11757,N_11667);
nor U11864 (N_11864,N_11746,N_11682);
and U11865 (N_11865,N_11734,N_11656);
and U11866 (N_11866,N_11749,N_11761);
or U11867 (N_11867,N_11689,N_11606);
xor U11868 (N_11868,N_11605,N_11729);
or U11869 (N_11869,N_11770,N_11668);
nand U11870 (N_11870,N_11747,N_11612);
xor U11871 (N_11871,N_11718,N_11627);
or U11872 (N_11872,N_11661,N_11690);
xnor U11873 (N_11873,N_11794,N_11795);
or U11874 (N_11874,N_11680,N_11678);
xnor U11875 (N_11875,N_11692,N_11636);
nor U11876 (N_11876,N_11665,N_11790);
or U11877 (N_11877,N_11620,N_11787);
nand U11878 (N_11878,N_11723,N_11659);
nor U11879 (N_11879,N_11632,N_11688);
or U11880 (N_11880,N_11696,N_11725);
and U11881 (N_11881,N_11779,N_11785);
nand U11882 (N_11882,N_11727,N_11694);
and U11883 (N_11883,N_11772,N_11649);
nand U11884 (N_11884,N_11633,N_11698);
xor U11885 (N_11885,N_11728,N_11707);
nand U11886 (N_11886,N_11782,N_11663);
nor U11887 (N_11887,N_11679,N_11626);
or U11888 (N_11888,N_11623,N_11721);
nor U11889 (N_11889,N_11753,N_11784);
or U11890 (N_11890,N_11684,N_11798);
xnor U11891 (N_11891,N_11715,N_11697);
or U11892 (N_11892,N_11797,N_11751);
xnor U11893 (N_11893,N_11738,N_11743);
or U11894 (N_11894,N_11648,N_11664);
nand U11895 (N_11895,N_11766,N_11726);
nor U11896 (N_11896,N_11793,N_11672);
nor U11897 (N_11897,N_11754,N_11774);
or U11898 (N_11898,N_11642,N_11771);
nand U11899 (N_11899,N_11722,N_11752);
xor U11900 (N_11900,N_11775,N_11699);
and U11901 (N_11901,N_11634,N_11744);
nor U11902 (N_11902,N_11768,N_11789);
nor U11903 (N_11903,N_11654,N_11707);
xnor U11904 (N_11904,N_11613,N_11767);
nand U11905 (N_11905,N_11761,N_11720);
or U11906 (N_11906,N_11689,N_11653);
xor U11907 (N_11907,N_11707,N_11681);
nor U11908 (N_11908,N_11636,N_11666);
or U11909 (N_11909,N_11779,N_11679);
xnor U11910 (N_11910,N_11726,N_11688);
and U11911 (N_11911,N_11762,N_11723);
and U11912 (N_11912,N_11796,N_11648);
nor U11913 (N_11913,N_11618,N_11638);
and U11914 (N_11914,N_11742,N_11757);
or U11915 (N_11915,N_11681,N_11655);
xnor U11916 (N_11916,N_11778,N_11697);
xnor U11917 (N_11917,N_11621,N_11601);
nand U11918 (N_11918,N_11616,N_11637);
xnor U11919 (N_11919,N_11720,N_11772);
and U11920 (N_11920,N_11661,N_11778);
or U11921 (N_11921,N_11651,N_11672);
nor U11922 (N_11922,N_11765,N_11707);
xor U11923 (N_11923,N_11619,N_11747);
xnor U11924 (N_11924,N_11751,N_11670);
nor U11925 (N_11925,N_11626,N_11696);
and U11926 (N_11926,N_11645,N_11796);
nand U11927 (N_11927,N_11648,N_11729);
xor U11928 (N_11928,N_11713,N_11718);
and U11929 (N_11929,N_11628,N_11646);
nor U11930 (N_11930,N_11686,N_11768);
nand U11931 (N_11931,N_11709,N_11728);
nand U11932 (N_11932,N_11694,N_11778);
and U11933 (N_11933,N_11612,N_11650);
or U11934 (N_11934,N_11739,N_11687);
and U11935 (N_11935,N_11736,N_11760);
nor U11936 (N_11936,N_11718,N_11722);
nor U11937 (N_11937,N_11618,N_11678);
xor U11938 (N_11938,N_11751,N_11771);
nand U11939 (N_11939,N_11706,N_11674);
nand U11940 (N_11940,N_11704,N_11647);
nand U11941 (N_11941,N_11731,N_11622);
nor U11942 (N_11942,N_11743,N_11695);
nand U11943 (N_11943,N_11637,N_11670);
nand U11944 (N_11944,N_11765,N_11628);
nor U11945 (N_11945,N_11674,N_11641);
and U11946 (N_11946,N_11693,N_11640);
or U11947 (N_11947,N_11666,N_11674);
xnor U11948 (N_11948,N_11672,N_11769);
and U11949 (N_11949,N_11674,N_11719);
and U11950 (N_11950,N_11786,N_11762);
nor U11951 (N_11951,N_11787,N_11650);
or U11952 (N_11952,N_11609,N_11722);
or U11953 (N_11953,N_11784,N_11640);
xnor U11954 (N_11954,N_11722,N_11622);
xor U11955 (N_11955,N_11654,N_11679);
and U11956 (N_11956,N_11750,N_11782);
nand U11957 (N_11957,N_11699,N_11653);
or U11958 (N_11958,N_11772,N_11692);
and U11959 (N_11959,N_11617,N_11751);
and U11960 (N_11960,N_11796,N_11794);
nor U11961 (N_11961,N_11634,N_11627);
nor U11962 (N_11962,N_11795,N_11646);
or U11963 (N_11963,N_11645,N_11769);
xor U11964 (N_11964,N_11718,N_11755);
nand U11965 (N_11965,N_11721,N_11731);
nand U11966 (N_11966,N_11748,N_11773);
and U11967 (N_11967,N_11618,N_11787);
xnor U11968 (N_11968,N_11646,N_11760);
xnor U11969 (N_11969,N_11601,N_11769);
or U11970 (N_11970,N_11772,N_11647);
nor U11971 (N_11971,N_11745,N_11617);
nand U11972 (N_11972,N_11785,N_11655);
and U11973 (N_11973,N_11774,N_11700);
or U11974 (N_11974,N_11747,N_11683);
or U11975 (N_11975,N_11613,N_11781);
nor U11976 (N_11976,N_11733,N_11606);
or U11977 (N_11977,N_11754,N_11747);
xor U11978 (N_11978,N_11702,N_11662);
xor U11979 (N_11979,N_11674,N_11758);
and U11980 (N_11980,N_11762,N_11772);
or U11981 (N_11981,N_11683,N_11741);
nand U11982 (N_11982,N_11704,N_11777);
nor U11983 (N_11983,N_11663,N_11759);
and U11984 (N_11984,N_11735,N_11700);
or U11985 (N_11985,N_11650,N_11658);
or U11986 (N_11986,N_11734,N_11612);
or U11987 (N_11987,N_11639,N_11755);
nand U11988 (N_11988,N_11737,N_11658);
nor U11989 (N_11989,N_11683,N_11682);
xnor U11990 (N_11990,N_11725,N_11673);
nand U11991 (N_11991,N_11652,N_11794);
nand U11992 (N_11992,N_11778,N_11651);
or U11993 (N_11993,N_11716,N_11698);
nand U11994 (N_11994,N_11647,N_11632);
and U11995 (N_11995,N_11751,N_11762);
nand U11996 (N_11996,N_11652,N_11755);
and U11997 (N_11997,N_11668,N_11702);
nand U11998 (N_11998,N_11786,N_11767);
xnor U11999 (N_11999,N_11759,N_11632);
or U12000 (N_12000,N_11830,N_11816);
and U12001 (N_12001,N_11971,N_11800);
and U12002 (N_12002,N_11872,N_11928);
and U12003 (N_12003,N_11880,N_11992);
nor U12004 (N_12004,N_11814,N_11913);
nor U12005 (N_12005,N_11807,N_11818);
xor U12006 (N_12006,N_11833,N_11918);
nand U12007 (N_12007,N_11850,N_11966);
xnor U12008 (N_12008,N_11988,N_11963);
nor U12009 (N_12009,N_11848,N_11851);
and U12010 (N_12010,N_11859,N_11977);
and U12011 (N_12011,N_11924,N_11939);
and U12012 (N_12012,N_11843,N_11875);
or U12013 (N_12013,N_11975,N_11906);
nor U12014 (N_12014,N_11810,N_11998);
xor U12015 (N_12015,N_11915,N_11813);
nand U12016 (N_12016,N_11925,N_11922);
xnor U12017 (N_12017,N_11914,N_11969);
xor U12018 (N_12018,N_11984,N_11957);
xor U12019 (N_12019,N_11940,N_11888);
nor U12020 (N_12020,N_11997,N_11889);
and U12021 (N_12021,N_11996,N_11912);
or U12022 (N_12022,N_11974,N_11867);
nor U12023 (N_12023,N_11927,N_11802);
nor U12024 (N_12024,N_11943,N_11852);
xor U12025 (N_12025,N_11891,N_11942);
nand U12026 (N_12026,N_11962,N_11999);
nor U12027 (N_12027,N_11834,N_11917);
or U12028 (N_12028,N_11860,N_11865);
or U12029 (N_12029,N_11964,N_11900);
or U12030 (N_12030,N_11911,N_11862);
and U12031 (N_12031,N_11883,N_11908);
and U12032 (N_12032,N_11958,N_11990);
nand U12033 (N_12033,N_11929,N_11920);
nand U12034 (N_12034,N_11973,N_11841);
xnor U12035 (N_12035,N_11948,N_11835);
xnor U12036 (N_12036,N_11854,N_11960);
or U12037 (N_12037,N_11886,N_11968);
xnor U12038 (N_12038,N_11876,N_11897);
nor U12039 (N_12039,N_11882,N_11832);
xnor U12040 (N_12040,N_11831,N_11874);
xor U12041 (N_12041,N_11804,N_11879);
nor U12042 (N_12042,N_11936,N_11801);
and U12043 (N_12043,N_11907,N_11910);
nand U12044 (N_12044,N_11817,N_11961);
and U12045 (N_12045,N_11864,N_11979);
nand U12046 (N_12046,N_11954,N_11965);
nand U12047 (N_12047,N_11902,N_11898);
and U12048 (N_12048,N_11858,N_11950);
or U12049 (N_12049,N_11887,N_11839);
nor U12050 (N_12050,N_11894,N_11982);
or U12051 (N_12051,N_11809,N_11935);
xor U12052 (N_12052,N_11855,N_11993);
or U12053 (N_12053,N_11921,N_11926);
xnor U12054 (N_12054,N_11904,N_11978);
or U12055 (N_12055,N_11892,N_11844);
nor U12056 (N_12056,N_11986,N_11870);
or U12057 (N_12057,N_11947,N_11923);
or U12058 (N_12058,N_11890,N_11896);
nor U12059 (N_12059,N_11949,N_11980);
nand U12060 (N_12060,N_11873,N_11853);
or U12061 (N_12061,N_11951,N_11972);
nor U12062 (N_12062,N_11811,N_11869);
and U12063 (N_12063,N_11885,N_11983);
nor U12064 (N_12064,N_11829,N_11930);
and U12065 (N_12065,N_11823,N_11836);
or U12066 (N_12066,N_11952,N_11955);
or U12067 (N_12067,N_11934,N_11953);
nor U12068 (N_12068,N_11849,N_11846);
or U12069 (N_12069,N_11985,N_11857);
nor U12070 (N_12070,N_11884,N_11893);
xor U12071 (N_12071,N_11822,N_11824);
or U12072 (N_12072,N_11837,N_11805);
nor U12073 (N_12073,N_11877,N_11881);
xor U12074 (N_12074,N_11903,N_11981);
nor U12075 (N_12075,N_11847,N_11899);
nand U12076 (N_12076,N_11991,N_11905);
nand U12077 (N_12077,N_11987,N_11827);
or U12078 (N_12078,N_11863,N_11956);
and U12079 (N_12079,N_11840,N_11819);
nand U12080 (N_12080,N_11916,N_11933);
xnor U12081 (N_12081,N_11861,N_11808);
nor U12082 (N_12082,N_11909,N_11828);
nor U12083 (N_12083,N_11946,N_11941);
or U12084 (N_12084,N_11931,N_11842);
xnor U12085 (N_12085,N_11866,N_11967);
nor U12086 (N_12086,N_11976,N_11838);
nand U12087 (N_12087,N_11821,N_11812);
nand U12088 (N_12088,N_11845,N_11806);
nor U12089 (N_12089,N_11871,N_11959);
xor U12090 (N_12090,N_11938,N_11826);
nand U12091 (N_12091,N_11995,N_11945);
and U12092 (N_12092,N_11815,N_11970);
xor U12093 (N_12093,N_11937,N_11878);
nor U12094 (N_12094,N_11944,N_11825);
nor U12095 (N_12095,N_11856,N_11989);
and U12096 (N_12096,N_11820,N_11895);
or U12097 (N_12097,N_11868,N_11803);
nor U12098 (N_12098,N_11901,N_11932);
xor U12099 (N_12099,N_11994,N_11919);
and U12100 (N_12100,N_11807,N_11947);
or U12101 (N_12101,N_11808,N_11993);
xor U12102 (N_12102,N_11993,N_11848);
and U12103 (N_12103,N_11983,N_11926);
nor U12104 (N_12104,N_11903,N_11806);
xor U12105 (N_12105,N_11953,N_11933);
and U12106 (N_12106,N_11810,N_11911);
and U12107 (N_12107,N_11955,N_11815);
nor U12108 (N_12108,N_11988,N_11977);
nor U12109 (N_12109,N_11994,N_11961);
nand U12110 (N_12110,N_11876,N_11892);
or U12111 (N_12111,N_11879,N_11892);
xor U12112 (N_12112,N_11894,N_11870);
xnor U12113 (N_12113,N_11962,N_11983);
nor U12114 (N_12114,N_11935,N_11984);
nand U12115 (N_12115,N_11892,N_11867);
and U12116 (N_12116,N_11969,N_11878);
xor U12117 (N_12117,N_11897,N_11809);
nand U12118 (N_12118,N_11914,N_11841);
nand U12119 (N_12119,N_11883,N_11808);
xor U12120 (N_12120,N_11886,N_11991);
nor U12121 (N_12121,N_11828,N_11984);
or U12122 (N_12122,N_11842,N_11859);
nor U12123 (N_12123,N_11914,N_11989);
nor U12124 (N_12124,N_11835,N_11816);
nor U12125 (N_12125,N_11839,N_11853);
xnor U12126 (N_12126,N_11996,N_11919);
xor U12127 (N_12127,N_11919,N_11814);
nand U12128 (N_12128,N_11838,N_11991);
xor U12129 (N_12129,N_11851,N_11869);
nand U12130 (N_12130,N_11844,N_11813);
nand U12131 (N_12131,N_11807,N_11855);
nand U12132 (N_12132,N_11984,N_11821);
xor U12133 (N_12133,N_11930,N_11932);
nand U12134 (N_12134,N_11886,N_11964);
nand U12135 (N_12135,N_11823,N_11912);
or U12136 (N_12136,N_11899,N_11858);
xor U12137 (N_12137,N_11880,N_11928);
and U12138 (N_12138,N_11943,N_11960);
nand U12139 (N_12139,N_11873,N_11869);
and U12140 (N_12140,N_11811,N_11816);
nor U12141 (N_12141,N_11930,N_11977);
xor U12142 (N_12142,N_11944,N_11999);
and U12143 (N_12143,N_11804,N_11908);
nor U12144 (N_12144,N_11879,N_11869);
or U12145 (N_12145,N_11963,N_11995);
and U12146 (N_12146,N_11813,N_11832);
or U12147 (N_12147,N_11984,N_11993);
nor U12148 (N_12148,N_11827,N_11939);
nor U12149 (N_12149,N_11819,N_11955);
xnor U12150 (N_12150,N_11903,N_11916);
and U12151 (N_12151,N_11995,N_11847);
xor U12152 (N_12152,N_11893,N_11938);
nand U12153 (N_12153,N_11927,N_11906);
or U12154 (N_12154,N_11827,N_11951);
nor U12155 (N_12155,N_11890,N_11827);
or U12156 (N_12156,N_11821,N_11886);
nand U12157 (N_12157,N_11869,N_11864);
nand U12158 (N_12158,N_11939,N_11997);
or U12159 (N_12159,N_11971,N_11845);
xor U12160 (N_12160,N_11987,N_11854);
nand U12161 (N_12161,N_11991,N_11985);
nor U12162 (N_12162,N_11976,N_11953);
xnor U12163 (N_12163,N_11911,N_11866);
and U12164 (N_12164,N_11965,N_11843);
nor U12165 (N_12165,N_11948,N_11980);
or U12166 (N_12166,N_11945,N_11969);
xnor U12167 (N_12167,N_11830,N_11841);
or U12168 (N_12168,N_11800,N_11822);
or U12169 (N_12169,N_11926,N_11872);
nor U12170 (N_12170,N_11923,N_11911);
or U12171 (N_12171,N_11805,N_11810);
nor U12172 (N_12172,N_11961,N_11830);
nor U12173 (N_12173,N_11841,N_11981);
xnor U12174 (N_12174,N_11912,N_11974);
and U12175 (N_12175,N_11950,N_11952);
nor U12176 (N_12176,N_11990,N_11849);
or U12177 (N_12177,N_11843,N_11854);
xor U12178 (N_12178,N_11852,N_11817);
and U12179 (N_12179,N_11832,N_11868);
and U12180 (N_12180,N_11894,N_11976);
xnor U12181 (N_12181,N_11906,N_11941);
or U12182 (N_12182,N_11810,N_11944);
or U12183 (N_12183,N_11883,N_11913);
nand U12184 (N_12184,N_11823,N_11970);
or U12185 (N_12185,N_11989,N_11948);
xor U12186 (N_12186,N_11828,N_11853);
and U12187 (N_12187,N_11970,N_11853);
nand U12188 (N_12188,N_11948,N_11915);
nor U12189 (N_12189,N_11974,N_11915);
or U12190 (N_12190,N_11860,N_11955);
nor U12191 (N_12191,N_11896,N_11912);
nor U12192 (N_12192,N_11856,N_11805);
nand U12193 (N_12193,N_11837,N_11977);
or U12194 (N_12194,N_11813,N_11866);
nor U12195 (N_12195,N_11873,N_11846);
xnor U12196 (N_12196,N_11807,N_11814);
and U12197 (N_12197,N_11892,N_11890);
and U12198 (N_12198,N_11809,N_11816);
nor U12199 (N_12199,N_11989,N_11926);
nand U12200 (N_12200,N_12009,N_12033);
or U12201 (N_12201,N_12035,N_12155);
xor U12202 (N_12202,N_12113,N_12191);
or U12203 (N_12203,N_12089,N_12070);
and U12204 (N_12204,N_12180,N_12083);
xnor U12205 (N_12205,N_12114,N_12004);
nand U12206 (N_12206,N_12065,N_12162);
xor U12207 (N_12207,N_12008,N_12122);
and U12208 (N_12208,N_12138,N_12169);
nor U12209 (N_12209,N_12174,N_12166);
or U12210 (N_12210,N_12059,N_12184);
or U12211 (N_12211,N_12145,N_12023);
or U12212 (N_12212,N_12075,N_12194);
and U12213 (N_12213,N_12102,N_12044);
nor U12214 (N_12214,N_12096,N_12110);
xnor U12215 (N_12215,N_12189,N_12172);
nand U12216 (N_12216,N_12024,N_12199);
or U12217 (N_12217,N_12084,N_12177);
nand U12218 (N_12218,N_12056,N_12091);
or U12219 (N_12219,N_12055,N_12001);
and U12220 (N_12220,N_12073,N_12193);
nor U12221 (N_12221,N_12133,N_12064);
or U12222 (N_12222,N_12045,N_12063);
and U12223 (N_12223,N_12042,N_12149);
nor U12224 (N_12224,N_12049,N_12054);
and U12225 (N_12225,N_12144,N_12153);
or U12226 (N_12226,N_12074,N_12136);
xor U12227 (N_12227,N_12015,N_12118);
nand U12228 (N_12228,N_12156,N_12117);
xnor U12229 (N_12229,N_12173,N_12011);
xnor U12230 (N_12230,N_12178,N_12170);
nand U12231 (N_12231,N_12016,N_12010);
or U12232 (N_12232,N_12000,N_12098);
nor U12233 (N_12233,N_12041,N_12123);
nor U12234 (N_12234,N_12061,N_12147);
nor U12235 (N_12235,N_12040,N_12106);
or U12236 (N_12236,N_12088,N_12020);
or U12237 (N_12237,N_12012,N_12071);
xnor U12238 (N_12238,N_12120,N_12090);
nand U12239 (N_12239,N_12007,N_12132);
and U12240 (N_12240,N_12121,N_12068);
xor U12241 (N_12241,N_12058,N_12171);
and U12242 (N_12242,N_12101,N_12160);
and U12243 (N_12243,N_12053,N_12082);
and U12244 (N_12244,N_12176,N_12163);
xnor U12245 (N_12245,N_12148,N_12116);
nor U12246 (N_12246,N_12112,N_12181);
xnor U12247 (N_12247,N_12146,N_12027);
nand U12248 (N_12248,N_12046,N_12078);
or U12249 (N_12249,N_12105,N_12072);
xnor U12250 (N_12250,N_12018,N_12198);
or U12251 (N_12251,N_12167,N_12154);
or U12252 (N_12252,N_12095,N_12127);
nand U12253 (N_12253,N_12183,N_12037);
nand U12254 (N_12254,N_12187,N_12081);
and U12255 (N_12255,N_12043,N_12157);
or U12256 (N_12256,N_12125,N_12152);
or U12257 (N_12257,N_12124,N_12097);
nor U12258 (N_12258,N_12119,N_12188);
or U12259 (N_12259,N_12103,N_12062);
and U12260 (N_12260,N_12060,N_12057);
and U12261 (N_12261,N_12021,N_12052);
nor U12262 (N_12262,N_12047,N_12076);
or U12263 (N_12263,N_12161,N_12108);
or U12264 (N_12264,N_12079,N_12025);
and U12265 (N_12265,N_12107,N_12130);
nor U12266 (N_12266,N_12131,N_12067);
nand U12267 (N_12267,N_12002,N_12126);
or U12268 (N_12268,N_12017,N_12150);
and U12269 (N_12269,N_12069,N_12195);
or U12270 (N_12270,N_12026,N_12092);
nor U12271 (N_12271,N_12185,N_12077);
nor U12272 (N_12272,N_12129,N_12085);
and U12273 (N_12273,N_12151,N_12038);
nor U12274 (N_12274,N_12005,N_12109);
or U12275 (N_12275,N_12031,N_12164);
nand U12276 (N_12276,N_12036,N_12032);
and U12277 (N_12277,N_12168,N_12142);
nand U12278 (N_12278,N_12013,N_12066);
nand U12279 (N_12279,N_12019,N_12104);
xor U12280 (N_12280,N_12028,N_12190);
xnor U12281 (N_12281,N_12137,N_12141);
nor U12282 (N_12282,N_12022,N_12006);
and U12283 (N_12283,N_12143,N_12134);
nand U12284 (N_12284,N_12159,N_12030);
nor U12285 (N_12285,N_12135,N_12100);
nor U12286 (N_12286,N_12128,N_12093);
and U12287 (N_12287,N_12197,N_12029);
nand U12288 (N_12288,N_12192,N_12139);
nor U12289 (N_12289,N_12050,N_12099);
or U12290 (N_12290,N_12175,N_12014);
nand U12291 (N_12291,N_12003,N_12140);
and U12292 (N_12292,N_12111,N_12179);
nand U12293 (N_12293,N_12034,N_12115);
nor U12294 (N_12294,N_12086,N_12182);
nand U12295 (N_12295,N_12094,N_12165);
nor U12296 (N_12296,N_12158,N_12048);
or U12297 (N_12297,N_12087,N_12051);
and U12298 (N_12298,N_12196,N_12186);
xor U12299 (N_12299,N_12039,N_12080);
nor U12300 (N_12300,N_12131,N_12035);
or U12301 (N_12301,N_12037,N_12161);
nand U12302 (N_12302,N_12162,N_12037);
nand U12303 (N_12303,N_12105,N_12085);
and U12304 (N_12304,N_12191,N_12051);
nand U12305 (N_12305,N_12031,N_12063);
nand U12306 (N_12306,N_12187,N_12086);
xnor U12307 (N_12307,N_12191,N_12050);
or U12308 (N_12308,N_12015,N_12044);
or U12309 (N_12309,N_12109,N_12123);
and U12310 (N_12310,N_12108,N_12115);
xor U12311 (N_12311,N_12031,N_12123);
or U12312 (N_12312,N_12096,N_12046);
or U12313 (N_12313,N_12069,N_12038);
nor U12314 (N_12314,N_12073,N_12096);
and U12315 (N_12315,N_12040,N_12109);
nand U12316 (N_12316,N_12046,N_12076);
nand U12317 (N_12317,N_12164,N_12120);
or U12318 (N_12318,N_12103,N_12091);
and U12319 (N_12319,N_12063,N_12124);
xnor U12320 (N_12320,N_12118,N_12196);
nand U12321 (N_12321,N_12050,N_12093);
or U12322 (N_12322,N_12029,N_12097);
nand U12323 (N_12323,N_12169,N_12145);
or U12324 (N_12324,N_12190,N_12119);
or U12325 (N_12325,N_12014,N_12023);
and U12326 (N_12326,N_12181,N_12186);
or U12327 (N_12327,N_12102,N_12144);
or U12328 (N_12328,N_12182,N_12127);
and U12329 (N_12329,N_12114,N_12096);
and U12330 (N_12330,N_12000,N_12196);
nor U12331 (N_12331,N_12066,N_12140);
or U12332 (N_12332,N_12021,N_12073);
nand U12333 (N_12333,N_12046,N_12119);
or U12334 (N_12334,N_12173,N_12187);
nor U12335 (N_12335,N_12134,N_12030);
nor U12336 (N_12336,N_12111,N_12159);
nor U12337 (N_12337,N_12098,N_12163);
and U12338 (N_12338,N_12125,N_12036);
nor U12339 (N_12339,N_12129,N_12049);
and U12340 (N_12340,N_12026,N_12195);
or U12341 (N_12341,N_12120,N_12093);
nand U12342 (N_12342,N_12122,N_12097);
nor U12343 (N_12343,N_12106,N_12077);
nand U12344 (N_12344,N_12151,N_12184);
xnor U12345 (N_12345,N_12119,N_12026);
xor U12346 (N_12346,N_12003,N_12090);
xnor U12347 (N_12347,N_12038,N_12054);
or U12348 (N_12348,N_12175,N_12064);
nand U12349 (N_12349,N_12050,N_12147);
nor U12350 (N_12350,N_12142,N_12111);
and U12351 (N_12351,N_12098,N_12197);
and U12352 (N_12352,N_12062,N_12054);
nand U12353 (N_12353,N_12094,N_12088);
nor U12354 (N_12354,N_12097,N_12076);
or U12355 (N_12355,N_12096,N_12199);
nor U12356 (N_12356,N_12028,N_12083);
nor U12357 (N_12357,N_12003,N_12104);
nand U12358 (N_12358,N_12027,N_12184);
xnor U12359 (N_12359,N_12180,N_12109);
or U12360 (N_12360,N_12076,N_12128);
xor U12361 (N_12361,N_12110,N_12054);
nor U12362 (N_12362,N_12005,N_12063);
nor U12363 (N_12363,N_12013,N_12128);
and U12364 (N_12364,N_12144,N_12135);
nand U12365 (N_12365,N_12018,N_12124);
and U12366 (N_12366,N_12014,N_12029);
xnor U12367 (N_12367,N_12037,N_12061);
nand U12368 (N_12368,N_12013,N_12117);
or U12369 (N_12369,N_12018,N_12195);
and U12370 (N_12370,N_12097,N_12144);
nor U12371 (N_12371,N_12012,N_12101);
nor U12372 (N_12372,N_12163,N_12043);
nand U12373 (N_12373,N_12070,N_12059);
nor U12374 (N_12374,N_12105,N_12195);
or U12375 (N_12375,N_12119,N_12159);
nand U12376 (N_12376,N_12136,N_12020);
nor U12377 (N_12377,N_12123,N_12101);
or U12378 (N_12378,N_12135,N_12134);
or U12379 (N_12379,N_12006,N_12101);
nand U12380 (N_12380,N_12118,N_12062);
xor U12381 (N_12381,N_12047,N_12184);
nor U12382 (N_12382,N_12050,N_12043);
nand U12383 (N_12383,N_12132,N_12100);
xnor U12384 (N_12384,N_12106,N_12066);
or U12385 (N_12385,N_12155,N_12054);
xnor U12386 (N_12386,N_12146,N_12014);
xnor U12387 (N_12387,N_12180,N_12195);
nor U12388 (N_12388,N_12153,N_12005);
nor U12389 (N_12389,N_12161,N_12052);
and U12390 (N_12390,N_12149,N_12054);
or U12391 (N_12391,N_12162,N_12027);
xor U12392 (N_12392,N_12007,N_12120);
and U12393 (N_12393,N_12142,N_12098);
nor U12394 (N_12394,N_12004,N_12023);
or U12395 (N_12395,N_12157,N_12117);
nor U12396 (N_12396,N_12122,N_12117);
xnor U12397 (N_12397,N_12140,N_12013);
xor U12398 (N_12398,N_12093,N_12114);
nand U12399 (N_12399,N_12136,N_12149);
or U12400 (N_12400,N_12240,N_12252);
xnor U12401 (N_12401,N_12228,N_12303);
or U12402 (N_12402,N_12395,N_12205);
and U12403 (N_12403,N_12298,N_12321);
nand U12404 (N_12404,N_12317,N_12238);
nor U12405 (N_12405,N_12275,N_12312);
xnor U12406 (N_12406,N_12387,N_12365);
and U12407 (N_12407,N_12210,N_12237);
nor U12408 (N_12408,N_12230,N_12284);
xnor U12409 (N_12409,N_12366,N_12300);
nand U12410 (N_12410,N_12227,N_12364);
nor U12411 (N_12411,N_12213,N_12305);
nor U12412 (N_12412,N_12229,N_12201);
and U12413 (N_12413,N_12242,N_12335);
nor U12414 (N_12414,N_12200,N_12330);
and U12415 (N_12415,N_12338,N_12336);
or U12416 (N_12416,N_12307,N_12322);
nor U12417 (N_12417,N_12225,N_12398);
xnor U12418 (N_12418,N_12260,N_12209);
xnor U12419 (N_12419,N_12306,N_12292);
or U12420 (N_12420,N_12232,N_12358);
and U12421 (N_12421,N_12318,N_12320);
and U12422 (N_12422,N_12382,N_12219);
xnor U12423 (N_12423,N_12344,N_12396);
nor U12424 (N_12424,N_12270,N_12278);
or U12425 (N_12425,N_12286,N_12223);
and U12426 (N_12426,N_12363,N_12394);
nand U12427 (N_12427,N_12215,N_12206);
or U12428 (N_12428,N_12296,N_12380);
nand U12429 (N_12429,N_12362,N_12202);
xor U12430 (N_12430,N_12257,N_12354);
xor U12431 (N_12431,N_12341,N_12258);
nand U12432 (N_12432,N_12309,N_12231);
nand U12433 (N_12433,N_12248,N_12283);
nand U12434 (N_12434,N_12261,N_12323);
nand U12435 (N_12435,N_12385,N_12218);
and U12436 (N_12436,N_12333,N_12379);
and U12437 (N_12437,N_12288,N_12376);
nand U12438 (N_12438,N_12374,N_12253);
and U12439 (N_12439,N_12384,N_12381);
or U12440 (N_12440,N_12246,N_12235);
nand U12441 (N_12441,N_12327,N_12311);
and U12442 (N_12442,N_12370,N_12247);
xor U12443 (N_12443,N_12272,N_12373);
and U12444 (N_12444,N_12388,N_12291);
nand U12445 (N_12445,N_12371,N_12222);
and U12446 (N_12446,N_12269,N_12273);
nor U12447 (N_12447,N_12244,N_12359);
xnor U12448 (N_12448,N_12256,N_12264);
nand U12449 (N_12449,N_12226,N_12343);
xor U12450 (N_12450,N_12266,N_12353);
nor U12451 (N_12451,N_12314,N_12351);
or U12452 (N_12452,N_12375,N_12313);
and U12453 (N_12453,N_12308,N_12294);
xnor U12454 (N_12454,N_12319,N_12290);
or U12455 (N_12455,N_12243,N_12368);
or U12456 (N_12456,N_12204,N_12271);
nand U12457 (N_12457,N_12331,N_12262);
and U12458 (N_12458,N_12295,N_12268);
nor U12459 (N_12459,N_12399,N_12282);
xor U12460 (N_12460,N_12301,N_12357);
nor U12461 (N_12461,N_12337,N_12236);
nand U12462 (N_12462,N_12233,N_12241);
and U12463 (N_12463,N_12392,N_12287);
nand U12464 (N_12464,N_12208,N_12285);
xor U12465 (N_12465,N_12281,N_12342);
nor U12466 (N_12466,N_12310,N_12378);
xor U12467 (N_12467,N_12332,N_12390);
and U12468 (N_12468,N_12265,N_12249);
nand U12469 (N_12469,N_12346,N_12355);
nor U12470 (N_12470,N_12280,N_12367);
or U12471 (N_12471,N_12239,N_12315);
and U12472 (N_12472,N_12369,N_12224);
and U12473 (N_12473,N_12277,N_12212);
or U12474 (N_12474,N_12214,N_12276);
nand U12475 (N_12475,N_12383,N_12245);
or U12476 (N_12476,N_12326,N_12203);
xnor U12477 (N_12477,N_12274,N_12293);
and U12478 (N_12478,N_12234,N_12334);
nand U12479 (N_12479,N_12267,N_12220);
xor U12480 (N_12480,N_12348,N_12347);
nand U12481 (N_12481,N_12360,N_12329);
xor U12482 (N_12482,N_12393,N_12349);
nor U12483 (N_12483,N_12350,N_12339);
nor U12484 (N_12484,N_12372,N_12361);
nor U12485 (N_12485,N_12299,N_12389);
or U12486 (N_12486,N_12259,N_12302);
nor U12487 (N_12487,N_12352,N_12356);
or U12488 (N_12488,N_12325,N_12255);
or U12489 (N_12489,N_12216,N_12386);
xor U12490 (N_12490,N_12289,N_12211);
nor U12491 (N_12491,N_12345,N_12377);
xnor U12492 (N_12492,N_12324,N_12207);
and U12493 (N_12493,N_12217,N_12391);
and U12494 (N_12494,N_12263,N_12251);
or U12495 (N_12495,N_12397,N_12304);
or U12496 (N_12496,N_12316,N_12297);
nor U12497 (N_12497,N_12328,N_12254);
xnor U12498 (N_12498,N_12340,N_12250);
and U12499 (N_12499,N_12221,N_12279);
and U12500 (N_12500,N_12387,N_12376);
xor U12501 (N_12501,N_12347,N_12321);
xor U12502 (N_12502,N_12342,N_12246);
or U12503 (N_12503,N_12363,N_12331);
and U12504 (N_12504,N_12332,N_12212);
nor U12505 (N_12505,N_12210,N_12233);
and U12506 (N_12506,N_12375,N_12390);
and U12507 (N_12507,N_12397,N_12283);
nand U12508 (N_12508,N_12295,N_12248);
nand U12509 (N_12509,N_12287,N_12267);
and U12510 (N_12510,N_12363,N_12235);
nor U12511 (N_12511,N_12299,N_12247);
or U12512 (N_12512,N_12357,N_12376);
or U12513 (N_12513,N_12235,N_12361);
xnor U12514 (N_12514,N_12272,N_12328);
and U12515 (N_12515,N_12396,N_12225);
nand U12516 (N_12516,N_12367,N_12271);
xnor U12517 (N_12517,N_12299,N_12287);
or U12518 (N_12518,N_12300,N_12215);
or U12519 (N_12519,N_12226,N_12271);
nor U12520 (N_12520,N_12317,N_12269);
nor U12521 (N_12521,N_12314,N_12382);
nand U12522 (N_12522,N_12281,N_12287);
and U12523 (N_12523,N_12232,N_12398);
and U12524 (N_12524,N_12227,N_12374);
and U12525 (N_12525,N_12249,N_12323);
nor U12526 (N_12526,N_12338,N_12213);
or U12527 (N_12527,N_12240,N_12349);
and U12528 (N_12528,N_12202,N_12338);
and U12529 (N_12529,N_12284,N_12345);
and U12530 (N_12530,N_12275,N_12344);
or U12531 (N_12531,N_12345,N_12210);
nor U12532 (N_12532,N_12293,N_12270);
nor U12533 (N_12533,N_12373,N_12242);
or U12534 (N_12534,N_12281,N_12296);
nand U12535 (N_12535,N_12342,N_12247);
or U12536 (N_12536,N_12275,N_12314);
nor U12537 (N_12537,N_12381,N_12392);
xnor U12538 (N_12538,N_12348,N_12393);
nor U12539 (N_12539,N_12266,N_12243);
or U12540 (N_12540,N_12344,N_12366);
and U12541 (N_12541,N_12352,N_12341);
nand U12542 (N_12542,N_12274,N_12253);
and U12543 (N_12543,N_12320,N_12342);
nand U12544 (N_12544,N_12293,N_12345);
nor U12545 (N_12545,N_12320,N_12324);
or U12546 (N_12546,N_12292,N_12204);
nand U12547 (N_12547,N_12320,N_12360);
nor U12548 (N_12548,N_12307,N_12238);
and U12549 (N_12549,N_12233,N_12275);
and U12550 (N_12550,N_12398,N_12376);
xnor U12551 (N_12551,N_12384,N_12229);
and U12552 (N_12552,N_12363,N_12242);
and U12553 (N_12553,N_12385,N_12396);
or U12554 (N_12554,N_12375,N_12374);
nand U12555 (N_12555,N_12251,N_12265);
nor U12556 (N_12556,N_12202,N_12344);
xor U12557 (N_12557,N_12221,N_12360);
and U12558 (N_12558,N_12354,N_12315);
and U12559 (N_12559,N_12375,N_12392);
or U12560 (N_12560,N_12348,N_12327);
and U12561 (N_12561,N_12241,N_12240);
nand U12562 (N_12562,N_12279,N_12290);
nand U12563 (N_12563,N_12251,N_12340);
nand U12564 (N_12564,N_12358,N_12307);
and U12565 (N_12565,N_12379,N_12242);
and U12566 (N_12566,N_12200,N_12253);
nor U12567 (N_12567,N_12312,N_12357);
nor U12568 (N_12568,N_12258,N_12371);
and U12569 (N_12569,N_12268,N_12371);
and U12570 (N_12570,N_12213,N_12325);
nand U12571 (N_12571,N_12292,N_12305);
or U12572 (N_12572,N_12340,N_12233);
nand U12573 (N_12573,N_12220,N_12315);
or U12574 (N_12574,N_12345,N_12226);
nor U12575 (N_12575,N_12289,N_12290);
xnor U12576 (N_12576,N_12209,N_12287);
nand U12577 (N_12577,N_12314,N_12311);
nor U12578 (N_12578,N_12261,N_12331);
xnor U12579 (N_12579,N_12272,N_12233);
nor U12580 (N_12580,N_12217,N_12358);
or U12581 (N_12581,N_12230,N_12343);
nor U12582 (N_12582,N_12232,N_12250);
nor U12583 (N_12583,N_12319,N_12214);
xor U12584 (N_12584,N_12244,N_12283);
and U12585 (N_12585,N_12326,N_12280);
nand U12586 (N_12586,N_12362,N_12208);
nor U12587 (N_12587,N_12249,N_12266);
nand U12588 (N_12588,N_12357,N_12371);
nand U12589 (N_12589,N_12379,N_12360);
xor U12590 (N_12590,N_12238,N_12290);
or U12591 (N_12591,N_12312,N_12380);
or U12592 (N_12592,N_12381,N_12259);
xor U12593 (N_12593,N_12337,N_12346);
nand U12594 (N_12594,N_12347,N_12322);
xnor U12595 (N_12595,N_12201,N_12289);
or U12596 (N_12596,N_12217,N_12203);
xor U12597 (N_12597,N_12241,N_12206);
nor U12598 (N_12598,N_12278,N_12345);
nor U12599 (N_12599,N_12302,N_12398);
and U12600 (N_12600,N_12524,N_12499);
nor U12601 (N_12601,N_12598,N_12563);
nor U12602 (N_12602,N_12576,N_12578);
nor U12603 (N_12603,N_12527,N_12487);
nor U12604 (N_12604,N_12519,N_12450);
xnor U12605 (N_12605,N_12407,N_12402);
and U12606 (N_12606,N_12416,N_12496);
nor U12607 (N_12607,N_12458,N_12534);
or U12608 (N_12608,N_12425,N_12506);
nor U12609 (N_12609,N_12514,N_12501);
xnor U12610 (N_12610,N_12565,N_12522);
or U12611 (N_12611,N_12401,N_12415);
nor U12612 (N_12612,N_12595,N_12538);
or U12613 (N_12613,N_12568,N_12446);
nor U12614 (N_12614,N_12422,N_12488);
xnor U12615 (N_12615,N_12433,N_12594);
or U12616 (N_12616,N_12587,N_12532);
nor U12617 (N_12617,N_12596,N_12404);
nand U12618 (N_12618,N_12477,N_12569);
nor U12619 (N_12619,N_12517,N_12471);
nor U12620 (N_12620,N_12434,N_12489);
xnor U12621 (N_12621,N_12573,N_12561);
nor U12622 (N_12622,N_12559,N_12406);
xnor U12623 (N_12623,N_12462,N_12591);
xnor U12624 (N_12624,N_12507,N_12555);
or U12625 (N_12625,N_12544,N_12479);
and U12626 (N_12626,N_12592,N_12583);
nor U12627 (N_12627,N_12585,N_12593);
xnor U12628 (N_12628,N_12432,N_12579);
nor U12629 (N_12629,N_12581,N_12494);
nor U12630 (N_12630,N_12562,N_12413);
xor U12631 (N_12631,N_12481,N_12580);
nand U12632 (N_12632,N_12497,N_12537);
and U12633 (N_12633,N_12550,N_12521);
or U12634 (N_12634,N_12525,N_12539);
and U12635 (N_12635,N_12536,N_12574);
xor U12636 (N_12636,N_12528,N_12518);
xor U12637 (N_12637,N_12451,N_12505);
nand U12638 (N_12638,N_12546,N_12428);
and U12639 (N_12639,N_12504,N_12473);
xor U12640 (N_12640,N_12548,N_12468);
and U12641 (N_12641,N_12449,N_12436);
nor U12642 (N_12642,N_12426,N_12557);
nand U12643 (N_12643,N_12582,N_12408);
xnor U12644 (N_12644,N_12540,N_12466);
xor U12645 (N_12645,N_12414,N_12438);
xor U12646 (N_12646,N_12552,N_12455);
nor U12647 (N_12647,N_12543,N_12502);
or U12648 (N_12648,N_12599,N_12470);
and U12649 (N_12649,N_12560,N_12431);
nor U12650 (N_12650,N_12558,N_12590);
nor U12651 (N_12651,N_12570,N_12495);
and U12652 (N_12652,N_12472,N_12589);
nand U12653 (N_12653,N_12551,N_12509);
and U12654 (N_12654,N_12443,N_12515);
nor U12655 (N_12655,N_12584,N_12498);
nand U12656 (N_12656,N_12491,N_12435);
or U12657 (N_12657,N_12424,N_12447);
or U12658 (N_12658,N_12508,N_12500);
or U12659 (N_12659,N_12427,N_12530);
nand U12660 (N_12660,N_12531,N_12547);
and U12661 (N_12661,N_12465,N_12549);
xnor U12662 (N_12662,N_12533,N_12445);
or U12663 (N_12663,N_12474,N_12448);
nor U12664 (N_12664,N_12577,N_12480);
and U12665 (N_12665,N_12571,N_12418);
or U12666 (N_12666,N_12456,N_12457);
nor U12667 (N_12667,N_12483,N_12588);
or U12668 (N_12668,N_12510,N_12529);
or U12669 (N_12669,N_12556,N_12511);
nor U12670 (N_12670,N_12463,N_12545);
xor U12671 (N_12671,N_12400,N_12441);
and U12672 (N_12672,N_12410,N_12503);
xnor U12673 (N_12673,N_12490,N_12542);
xnor U12674 (N_12674,N_12437,N_12464);
nand U12675 (N_12675,N_12484,N_12412);
nand U12676 (N_12676,N_12460,N_12564);
xor U12677 (N_12677,N_12423,N_12467);
nor U12678 (N_12678,N_12421,N_12442);
nand U12679 (N_12679,N_12478,N_12513);
nor U12680 (N_12680,N_12520,N_12419);
nor U12681 (N_12681,N_12567,N_12411);
nor U12682 (N_12682,N_12409,N_12586);
nor U12683 (N_12683,N_12512,N_12523);
nand U12684 (N_12684,N_12461,N_12485);
xnor U12685 (N_12685,N_12475,N_12430);
nor U12686 (N_12686,N_12403,N_12566);
nand U12687 (N_12687,N_12452,N_12493);
nand U12688 (N_12688,N_12439,N_12454);
nor U12689 (N_12689,N_12516,N_12440);
or U12690 (N_12690,N_12444,N_12476);
or U12691 (N_12691,N_12554,N_12492);
or U12692 (N_12692,N_12469,N_12597);
nor U12693 (N_12693,N_12420,N_12459);
and U12694 (N_12694,N_12405,N_12417);
nor U12695 (N_12695,N_12429,N_12453);
nand U12696 (N_12696,N_12575,N_12541);
nor U12697 (N_12697,N_12553,N_12482);
xnor U12698 (N_12698,N_12535,N_12526);
nand U12699 (N_12699,N_12572,N_12486);
or U12700 (N_12700,N_12500,N_12496);
xnor U12701 (N_12701,N_12533,N_12472);
nand U12702 (N_12702,N_12503,N_12457);
nand U12703 (N_12703,N_12557,N_12470);
xnor U12704 (N_12704,N_12599,N_12441);
or U12705 (N_12705,N_12412,N_12435);
nand U12706 (N_12706,N_12591,N_12504);
xnor U12707 (N_12707,N_12471,N_12414);
xor U12708 (N_12708,N_12541,N_12450);
nand U12709 (N_12709,N_12576,N_12456);
nand U12710 (N_12710,N_12496,N_12531);
nor U12711 (N_12711,N_12577,N_12531);
and U12712 (N_12712,N_12401,N_12575);
nor U12713 (N_12713,N_12424,N_12425);
nor U12714 (N_12714,N_12520,N_12489);
and U12715 (N_12715,N_12415,N_12438);
nand U12716 (N_12716,N_12472,N_12496);
nand U12717 (N_12717,N_12573,N_12534);
and U12718 (N_12718,N_12582,N_12564);
xor U12719 (N_12719,N_12480,N_12417);
or U12720 (N_12720,N_12539,N_12519);
nor U12721 (N_12721,N_12434,N_12533);
or U12722 (N_12722,N_12529,N_12511);
or U12723 (N_12723,N_12408,N_12404);
nor U12724 (N_12724,N_12542,N_12588);
xor U12725 (N_12725,N_12526,N_12419);
nor U12726 (N_12726,N_12467,N_12521);
nand U12727 (N_12727,N_12540,N_12492);
or U12728 (N_12728,N_12512,N_12489);
and U12729 (N_12729,N_12408,N_12424);
nand U12730 (N_12730,N_12548,N_12588);
or U12731 (N_12731,N_12418,N_12550);
and U12732 (N_12732,N_12543,N_12548);
xnor U12733 (N_12733,N_12500,N_12411);
nor U12734 (N_12734,N_12468,N_12490);
nor U12735 (N_12735,N_12550,N_12556);
nor U12736 (N_12736,N_12567,N_12400);
or U12737 (N_12737,N_12419,N_12417);
or U12738 (N_12738,N_12413,N_12450);
nor U12739 (N_12739,N_12422,N_12597);
or U12740 (N_12740,N_12509,N_12492);
nand U12741 (N_12741,N_12520,N_12445);
xor U12742 (N_12742,N_12500,N_12469);
xor U12743 (N_12743,N_12571,N_12543);
and U12744 (N_12744,N_12478,N_12417);
nand U12745 (N_12745,N_12584,N_12431);
and U12746 (N_12746,N_12538,N_12541);
nand U12747 (N_12747,N_12484,N_12419);
or U12748 (N_12748,N_12424,N_12472);
nor U12749 (N_12749,N_12488,N_12406);
nor U12750 (N_12750,N_12566,N_12441);
xnor U12751 (N_12751,N_12431,N_12495);
xor U12752 (N_12752,N_12469,N_12552);
or U12753 (N_12753,N_12440,N_12518);
xor U12754 (N_12754,N_12560,N_12497);
xor U12755 (N_12755,N_12476,N_12568);
nand U12756 (N_12756,N_12469,N_12470);
nor U12757 (N_12757,N_12457,N_12512);
nor U12758 (N_12758,N_12466,N_12492);
nor U12759 (N_12759,N_12561,N_12418);
nor U12760 (N_12760,N_12569,N_12433);
or U12761 (N_12761,N_12495,N_12598);
xnor U12762 (N_12762,N_12447,N_12513);
and U12763 (N_12763,N_12413,N_12537);
nand U12764 (N_12764,N_12437,N_12472);
or U12765 (N_12765,N_12539,N_12425);
nor U12766 (N_12766,N_12577,N_12538);
xor U12767 (N_12767,N_12443,N_12584);
nor U12768 (N_12768,N_12555,N_12407);
nand U12769 (N_12769,N_12552,N_12439);
nand U12770 (N_12770,N_12517,N_12526);
nand U12771 (N_12771,N_12530,N_12498);
or U12772 (N_12772,N_12557,N_12447);
or U12773 (N_12773,N_12576,N_12516);
xnor U12774 (N_12774,N_12515,N_12591);
nand U12775 (N_12775,N_12442,N_12436);
nand U12776 (N_12776,N_12513,N_12556);
nand U12777 (N_12777,N_12561,N_12508);
xnor U12778 (N_12778,N_12542,N_12414);
nand U12779 (N_12779,N_12428,N_12474);
xnor U12780 (N_12780,N_12520,N_12533);
and U12781 (N_12781,N_12458,N_12417);
nor U12782 (N_12782,N_12477,N_12555);
nand U12783 (N_12783,N_12467,N_12535);
xnor U12784 (N_12784,N_12505,N_12565);
or U12785 (N_12785,N_12517,N_12514);
xor U12786 (N_12786,N_12524,N_12550);
and U12787 (N_12787,N_12561,N_12407);
and U12788 (N_12788,N_12586,N_12464);
nor U12789 (N_12789,N_12422,N_12511);
xor U12790 (N_12790,N_12466,N_12588);
and U12791 (N_12791,N_12472,N_12440);
xor U12792 (N_12792,N_12549,N_12542);
xnor U12793 (N_12793,N_12451,N_12561);
or U12794 (N_12794,N_12541,N_12471);
xor U12795 (N_12795,N_12473,N_12595);
xnor U12796 (N_12796,N_12540,N_12541);
nand U12797 (N_12797,N_12440,N_12405);
xor U12798 (N_12798,N_12590,N_12513);
nand U12799 (N_12799,N_12437,N_12524);
or U12800 (N_12800,N_12769,N_12706);
nand U12801 (N_12801,N_12675,N_12610);
xor U12802 (N_12802,N_12739,N_12701);
nor U12803 (N_12803,N_12760,N_12779);
nand U12804 (N_12804,N_12679,N_12792);
or U12805 (N_12805,N_12607,N_12793);
nand U12806 (N_12806,N_12733,N_12713);
nor U12807 (N_12807,N_12752,N_12676);
and U12808 (N_12808,N_12641,N_12776);
or U12809 (N_12809,N_12666,N_12753);
nor U12810 (N_12810,N_12750,N_12609);
xor U12811 (N_12811,N_12672,N_12797);
nor U12812 (N_12812,N_12747,N_12684);
nor U12813 (N_12813,N_12765,N_12766);
or U12814 (N_12814,N_12748,N_12657);
nor U12815 (N_12815,N_12741,N_12649);
nand U12816 (N_12816,N_12788,N_12756);
or U12817 (N_12817,N_12658,N_12730);
nor U12818 (N_12818,N_12611,N_12694);
xor U12819 (N_12819,N_12763,N_12700);
and U12820 (N_12820,N_12715,N_12754);
xnor U12821 (N_12821,N_12600,N_12755);
and U12822 (N_12822,N_12671,N_12630);
and U12823 (N_12823,N_12697,N_12791);
xor U12824 (N_12824,N_12691,N_12648);
and U12825 (N_12825,N_12708,N_12709);
nor U12826 (N_12826,N_12742,N_12795);
xnor U12827 (N_12827,N_12743,N_12744);
nand U12828 (N_12828,N_12794,N_12703);
nor U12829 (N_12829,N_12652,N_12686);
nor U12830 (N_12830,N_12645,N_12674);
nand U12831 (N_12831,N_12624,N_12665);
nand U12832 (N_12832,N_12746,N_12762);
xnor U12833 (N_12833,N_12711,N_12618);
nor U12834 (N_12834,N_12654,N_12650);
nand U12835 (N_12835,N_12728,N_12617);
or U12836 (N_12836,N_12693,N_12628);
or U12837 (N_12837,N_12781,N_12629);
and U12838 (N_12838,N_12775,N_12616);
or U12839 (N_12839,N_12623,N_12651);
and U12840 (N_12840,N_12782,N_12667);
or U12841 (N_12841,N_12710,N_12780);
nor U12842 (N_12842,N_12695,N_12723);
nand U12843 (N_12843,N_12720,N_12613);
xnor U12844 (N_12844,N_12758,N_12699);
and U12845 (N_12845,N_12642,N_12719);
or U12846 (N_12846,N_12614,N_12688);
or U12847 (N_12847,N_12656,N_12660);
or U12848 (N_12848,N_12778,N_12721);
xnor U12849 (N_12849,N_12736,N_12659);
nand U12850 (N_12850,N_12751,N_12771);
xnor U12851 (N_12851,N_12673,N_12646);
nor U12852 (N_12852,N_12683,N_12682);
nor U12853 (N_12853,N_12789,N_12612);
nand U12854 (N_12854,N_12638,N_12664);
or U12855 (N_12855,N_12786,N_12772);
or U12856 (N_12856,N_12790,N_12640);
xnor U12857 (N_12857,N_12653,N_12687);
and U12858 (N_12858,N_12783,N_12681);
xor U12859 (N_12859,N_12689,N_12707);
xor U12860 (N_12860,N_12716,N_12661);
and U12861 (N_12861,N_12690,N_12669);
nand U12862 (N_12862,N_12725,N_12768);
nand U12863 (N_12863,N_12636,N_12685);
nand U12864 (N_12864,N_12738,N_12740);
xnor U12865 (N_12865,N_12620,N_12670);
xnor U12866 (N_12866,N_12632,N_12634);
xnor U12867 (N_12867,N_12732,N_12605);
nor U12868 (N_12868,N_12677,N_12601);
nand U12869 (N_12869,N_12608,N_12680);
nand U12870 (N_12870,N_12718,N_12626);
and U12871 (N_12871,N_12622,N_12714);
nor U12872 (N_12872,N_12767,N_12784);
and U12873 (N_12873,N_12717,N_12655);
nand U12874 (N_12874,N_12724,N_12734);
xnor U12875 (N_12875,N_12643,N_12668);
nor U12876 (N_12876,N_12727,N_12785);
xor U12877 (N_12877,N_12726,N_12663);
xor U12878 (N_12878,N_12604,N_12606);
nand U12879 (N_12879,N_12749,N_12639);
and U12880 (N_12880,N_12712,N_12745);
or U12881 (N_12881,N_12737,N_12770);
or U12882 (N_12882,N_12704,N_12602);
nor U12883 (N_12883,N_12722,N_12774);
nand U12884 (N_12884,N_12799,N_12627);
xnor U12885 (N_12885,N_12696,N_12798);
and U12886 (N_12886,N_12662,N_12678);
or U12887 (N_12887,N_12757,N_12764);
or U12888 (N_12888,N_12759,N_12621);
xnor U12889 (N_12889,N_12692,N_12647);
xnor U12890 (N_12890,N_12787,N_12705);
and U12891 (N_12891,N_12637,N_12625);
nand U12892 (N_12892,N_12698,N_12644);
xnor U12893 (N_12893,N_12761,N_12796);
and U12894 (N_12894,N_12603,N_12735);
xnor U12895 (N_12895,N_12777,N_12633);
nor U12896 (N_12896,N_12702,N_12729);
or U12897 (N_12897,N_12773,N_12731);
nor U12898 (N_12898,N_12631,N_12619);
nor U12899 (N_12899,N_12635,N_12615);
nand U12900 (N_12900,N_12739,N_12689);
nand U12901 (N_12901,N_12685,N_12621);
and U12902 (N_12902,N_12732,N_12748);
or U12903 (N_12903,N_12610,N_12776);
xnor U12904 (N_12904,N_12619,N_12613);
and U12905 (N_12905,N_12736,N_12721);
or U12906 (N_12906,N_12665,N_12630);
or U12907 (N_12907,N_12781,N_12630);
nor U12908 (N_12908,N_12683,N_12764);
and U12909 (N_12909,N_12644,N_12755);
nor U12910 (N_12910,N_12768,N_12671);
or U12911 (N_12911,N_12700,N_12650);
xor U12912 (N_12912,N_12771,N_12628);
or U12913 (N_12913,N_12702,N_12629);
or U12914 (N_12914,N_12795,N_12696);
nor U12915 (N_12915,N_12706,N_12655);
and U12916 (N_12916,N_12793,N_12758);
nand U12917 (N_12917,N_12660,N_12798);
nand U12918 (N_12918,N_12649,N_12776);
xor U12919 (N_12919,N_12610,N_12787);
nor U12920 (N_12920,N_12776,N_12775);
and U12921 (N_12921,N_12635,N_12690);
and U12922 (N_12922,N_12618,N_12797);
nand U12923 (N_12923,N_12672,N_12683);
nor U12924 (N_12924,N_12746,N_12750);
nand U12925 (N_12925,N_12701,N_12710);
nand U12926 (N_12926,N_12667,N_12719);
nand U12927 (N_12927,N_12634,N_12759);
or U12928 (N_12928,N_12674,N_12746);
nor U12929 (N_12929,N_12641,N_12675);
nand U12930 (N_12930,N_12699,N_12719);
nand U12931 (N_12931,N_12753,N_12619);
nand U12932 (N_12932,N_12603,N_12783);
or U12933 (N_12933,N_12642,N_12617);
and U12934 (N_12934,N_12628,N_12656);
nand U12935 (N_12935,N_12762,N_12725);
and U12936 (N_12936,N_12784,N_12715);
and U12937 (N_12937,N_12672,N_12773);
xnor U12938 (N_12938,N_12622,N_12732);
or U12939 (N_12939,N_12773,N_12681);
and U12940 (N_12940,N_12699,N_12743);
nor U12941 (N_12941,N_12643,N_12703);
and U12942 (N_12942,N_12669,N_12703);
nand U12943 (N_12943,N_12683,N_12668);
nor U12944 (N_12944,N_12602,N_12707);
nand U12945 (N_12945,N_12648,N_12711);
nor U12946 (N_12946,N_12633,N_12672);
and U12947 (N_12947,N_12757,N_12605);
or U12948 (N_12948,N_12752,N_12695);
nand U12949 (N_12949,N_12615,N_12747);
or U12950 (N_12950,N_12631,N_12686);
nor U12951 (N_12951,N_12713,N_12691);
nand U12952 (N_12952,N_12642,N_12648);
nor U12953 (N_12953,N_12619,N_12601);
and U12954 (N_12954,N_12690,N_12665);
nor U12955 (N_12955,N_12681,N_12785);
and U12956 (N_12956,N_12675,N_12662);
or U12957 (N_12957,N_12774,N_12627);
xor U12958 (N_12958,N_12606,N_12701);
or U12959 (N_12959,N_12673,N_12695);
and U12960 (N_12960,N_12762,N_12603);
or U12961 (N_12961,N_12798,N_12761);
or U12962 (N_12962,N_12766,N_12705);
xnor U12963 (N_12963,N_12771,N_12698);
or U12964 (N_12964,N_12627,N_12721);
and U12965 (N_12965,N_12613,N_12631);
or U12966 (N_12966,N_12616,N_12633);
or U12967 (N_12967,N_12767,N_12697);
nor U12968 (N_12968,N_12697,N_12664);
nand U12969 (N_12969,N_12628,N_12797);
nand U12970 (N_12970,N_12761,N_12733);
or U12971 (N_12971,N_12765,N_12652);
or U12972 (N_12972,N_12614,N_12717);
and U12973 (N_12973,N_12605,N_12628);
nand U12974 (N_12974,N_12748,N_12691);
xnor U12975 (N_12975,N_12642,N_12747);
xnor U12976 (N_12976,N_12631,N_12627);
nand U12977 (N_12977,N_12715,N_12792);
nand U12978 (N_12978,N_12677,N_12699);
nand U12979 (N_12979,N_12601,N_12771);
or U12980 (N_12980,N_12686,N_12731);
nand U12981 (N_12981,N_12757,N_12760);
and U12982 (N_12982,N_12762,N_12787);
and U12983 (N_12983,N_12756,N_12772);
and U12984 (N_12984,N_12634,N_12700);
or U12985 (N_12985,N_12779,N_12671);
nor U12986 (N_12986,N_12738,N_12705);
and U12987 (N_12987,N_12762,N_12706);
xnor U12988 (N_12988,N_12696,N_12629);
nand U12989 (N_12989,N_12764,N_12779);
nand U12990 (N_12990,N_12734,N_12662);
nor U12991 (N_12991,N_12713,N_12743);
nand U12992 (N_12992,N_12697,N_12646);
xnor U12993 (N_12993,N_12711,N_12691);
nand U12994 (N_12994,N_12681,N_12601);
or U12995 (N_12995,N_12794,N_12750);
xor U12996 (N_12996,N_12691,N_12708);
and U12997 (N_12997,N_12730,N_12696);
and U12998 (N_12998,N_12652,N_12631);
xnor U12999 (N_12999,N_12634,N_12791);
and U13000 (N_13000,N_12969,N_12882);
or U13001 (N_13001,N_12830,N_12886);
or U13002 (N_13002,N_12850,N_12845);
and U13003 (N_13003,N_12883,N_12881);
xnor U13004 (N_13004,N_12874,N_12937);
or U13005 (N_13005,N_12916,N_12909);
nand U13006 (N_13006,N_12933,N_12961);
and U13007 (N_13007,N_12953,N_12977);
and U13008 (N_13008,N_12905,N_12938);
and U13009 (N_13009,N_12818,N_12889);
nor U13010 (N_13010,N_12992,N_12834);
nor U13011 (N_13011,N_12800,N_12808);
nand U13012 (N_13012,N_12993,N_12939);
nor U13013 (N_13013,N_12803,N_12946);
nand U13014 (N_13014,N_12998,N_12848);
nand U13015 (N_13015,N_12892,N_12866);
nand U13016 (N_13016,N_12825,N_12989);
nand U13017 (N_13017,N_12828,N_12870);
or U13018 (N_13018,N_12832,N_12964);
or U13019 (N_13019,N_12943,N_12861);
and U13020 (N_13020,N_12922,N_12862);
nor U13021 (N_13021,N_12934,N_12910);
nor U13022 (N_13022,N_12954,N_12813);
nand U13023 (N_13023,N_12844,N_12987);
or U13024 (N_13024,N_12947,N_12841);
and U13025 (N_13025,N_12885,N_12871);
nand U13026 (N_13026,N_12991,N_12996);
nor U13027 (N_13027,N_12948,N_12847);
nand U13028 (N_13028,N_12801,N_12944);
and U13029 (N_13029,N_12923,N_12928);
nand U13030 (N_13030,N_12936,N_12864);
nand U13031 (N_13031,N_12994,N_12884);
nand U13032 (N_13032,N_12903,N_12853);
or U13033 (N_13033,N_12831,N_12887);
or U13034 (N_13034,N_12986,N_12907);
xor U13035 (N_13035,N_12880,N_12817);
xor U13036 (N_13036,N_12972,N_12959);
and U13037 (N_13037,N_12918,N_12904);
nor U13038 (N_13038,N_12901,N_12863);
or U13039 (N_13039,N_12966,N_12902);
nand U13040 (N_13040,N_12915,N_12980);
xor U13041 (N_13041,N_12958,N_12812);
nand U13042 (N_13042,N_12890,N_12900);
or U13043 (N_13043,N_12979,N_12925);
or U13044 (N_13044,N_12995,N_12842);
nand U13045 (N_13045,N_12868,N_12877);
nor U13046 (N_13046,N_12806,N_12962);
xnor U13047 (N_13047,N_12897,N_12858);
nand U13048 (N_13048,N_12895,N_12974);
and U13049 (N_13049,N_12839,N_12835);
and U13050 (N_13050,N_12810,N_12988);
and U13051 (N_13051,N_12978,N_12804);
or U13052 (N_13052,N_12956,N_12965);
nand U13053 (N_13053,N_12836,N_12814);
and U13054 (N_13054,N_12950,N_12869);
and U13055 (N_13055,N_12932,N_12908);
nor U13056 (N_13056,N_12906,N_12935);
nand U13057 (N_13057,N_12878,N_12855);
xor U13058 (N_13058,N_12949,N_12893);
xnor U13059 (N_13059,N_12963,N_12967);
or U13060 (N_13060,N_12894,N_12815);
xor U13061 (N_13061,N_12985,N_12941);
or U13062 (N_13062,N_12924,N_12945);
nor U13063 (N_13063,N_12824,N_12930);
xor U13064 (N_13064,N_12919,N_12872);
or U13065 (N_13065,N_12816,N_12957);
and U13066 (N_13066,N_12827,N_12968);
and U13067 (N_13067,N_12809,N_12876);
nand U13068 (N_13068,N_12807,N_12976);
or U13069 (N_13069,N_12990,N_12920);
xnor U13070 (N_13070,N_12837,N_12819);
xor U13071 (N_13071,N_12849,N_12971);
and U13072 (N_13072,N_12840,N_12982);
nand U13073 (N_13073,N_12888,N_12865);
nor U13074 (N_13074,N_12826,N_12873);
and U13075 (N_13075,N_12926,N_12896);
and U13076 (N_13076,N_12838,N_12940);
or U13077 (N_13077,N_12917,N_12952);
or U13078 (N_13078,N_12913,N_12856);
and U13079 (N_13079,N_12811,N_12822);
nor U13080 (N_13080,N_12914,N_12833);
nor U13081 (N_13081,N_12805,N_12875);
or U13082 (N_13082,N_12879,N_12820);
nor U13083 (N_13083,N_12891,N_12843);
and U13084 (N_13084,N_12942,N_12927);
nand U13085 (N_13085,N_12846,N_12852);
nand U13086 (N_13086,N_12975,N_12860);
xnor U13087 (N_13087,N_12899,N_12981);
and U13088 (N_13088,N_12983,N_12951);
nor U13089 (N_13089,N_12859,N_12851);
nor U13090 (N_13090,N_12854,N_12973);
or U13091 (N_13091,N_12898,N_12921);
nand U13092 (N_13092,N_12997,N_12823);
and U13093 (N_13093,N_12802,N_12929);
and U13094 (N_13094,N_12911,N_12867);
or U13095 (N_13095,N_12912,N_12931);
nor U13096 (N_13096,N_12960,N_12857);
and U13097 (N_13097,N_12984,N_12821);
xnor U13098 (N_13098,N_12970,N_12955);
and U13099 (N_13099,N_12829,N_12999);
or U13100 (N_13100,N_12990,N_12915);
xor U13101 (N_13101,N_12944,N_12818);
and U13102 (N_13102,N_12870,N_12917);
and U13103 (N_13103,N_12963,N_12848);
nor U13104 (N_13104,N_12805,N_12929);
xnor U13105 (N_13105,N_12836,N_12933);
nor U13106 (N_13106,N_12945,N_12875);
nand U13107 (N_13107,N_12866,N_12989);
nor U13108 (N_13108,N_12993,N_12811);
xor U13109 (N_13109,N_12919,N_12875);
and U13110 (N_13110,N_12873,N_12825);
nand U13111 (N_13111,N_12837,N_12914);
nand U13112 (N_13112,N_12802,N_12900);
xor U13113 (N_13113,N_12844,N_12825);
nand U13114 (N_13114,N_12923,N_12887);
nand U13115 (N_13115,N_12971,N_12824);
and U13116 (N_13116,N_12946,N_12957);
or U13117 (N_13117,N_12821,N_12806);
nor U13118 (N_13118,N_12970,N_12865);
and U13119 (N_13119,N_12856,N_12842);
nand U13120 (N_13120,N_12857,N_12892);
nand U13121 (N_13121,N_12899,N_12822);
nor U13122 (N_13122,N_12983,N_12887);
or U13123 (N_13123,N_12848,N_12906);
or U13124 (N_13124,N_12942,N_12908);
nand U13125 (N_13125,N_12832,N_12996);
or U13126 (N_13126,N_12841,N_12871);
or U13127 (N_13127,N_12847,N_12874);
xor U13128 (N_13128,N_12840,N_12925);
nand U13129 (N_13129,N_12960,N_12902);
and U13130 (N_13130,N_12859,N_12959);
xor U13131 (N_13131,N_12941,N_12831);
nor U13132 (N_13132,N_12848,N_12956);
or U13133 (N_13133,N_12954,N_12853);
and U13134 (N_13134,N_12861,N_12810);
or U13135 (N_13135,N_12854,N_12988);
nand U13136 (N_13136,N_12956,N_12882);
and U13137 (N_13137,N_12947,N_12994);
nor U13138 (N_13138,N_12813,N_12827);
nand U13139 (N_13139,N_12887,N_12970);
xor U13140 (N_13140,N_12973,N_12804);
or U13141 (N_13141,N_12891,N_12854);
xnor U13142 (N_13142,N_12836,N_12831);
nand U13143 (N_13143,N_12967,N_12903);
nor U13144 (N_13144,N_12985,N_12952);
nand U13145 (N_13145,N_12850,N_12808);
xor U13146 (N_13146,N_12844,N_12890);
nand U13147 (N_13147,N_12965,N_12806);
or U13148 (N_13148,N_12872,N_12831);
nand U13149 (N_13149,N_12940,N_12914);
nor U13150 (N_13150,N_12810,N_12806);
xnor U13151 (N_13151,N_12808,N_12976);
nand U13152 (N_13152,N_12964,N_12900);
and U13153 (N_13153,N_12997,N_12824);
and U13154 (N_13154,N_12970,N_12848);
xnor U13155 (N_13155,N_12966,N_12820);
and U13156 (N_13156,N_12855,N_12995);
xnor U13157 (N_13157,N_12896,N_12931);
or U13158 (N_13158,N_12907,N_12883);
nand U13159 (N_13159,N_12998,N_12906);
or U13160 (N_13160,N_12889,N_12829);
nor U13161 (N_13161,N_12968,N_12946);
nand U13162 (N_13162,N_12995,N_12802);
or U13163 (N_13163,N_12905,N_12804);
or U13164 (N_13164,N_12967,N_12970);
or U13165 (N_13165,N_12951,N_12899);
nand U13166 (N_13166,N_12818,N_12865);
or U13167 (N_13167,N_12835,N_12853);
nand U13168 (N_13168,N_12885,N_12892);
or U13169 (N_13169,N_12834,N_12880);
xnor U13170 (N_13170,N_12843,N_12970);
nand U13171 (N_13171,N_12989,N_12877);
nand U13172 (N_13172,N_12805,N_12816);
or U13173 (N_13173,N_12901,N_12896);
or U13174 (N_13174,N_12819,N_12869);
nor U13175 (N_13175,N_12932,N_12967);
or U13176 (N_13176,N_12884,N_12999);
nand U13177 (N_13177,N_12964,N_12898);
or U13178 (N_13178,N_12998,N_12855);
xor U13179 (N_13179,N_12898,N_12910);
and U13180 (N_13180,N_12979,N_12936);
and U13181 (N_13181,N_12913,N_12886);
nand U13182 (N_13182,N_12947,N_12906);
nand U13183 (N_13183,N_12826,N_12904);
nand U13184 (N_13184,N_12853,N_12907);
or U13185 (N_13185,N_12959,N_12855);
xor U13186 (N_13186,N_12851,N_12953);
and U13187 (N_13187,N_12827,N_12834);
nand U13188 (N_13188,N_12973,N_12989);
xnor U13189 (N_13189,N_12811,N_12878);
xnor U13190 (N_13190,N_12966,N_12908);
and U13191 (N_13191,N_12899,N_12931);
or U13192 (N_13192,N_12852,N_12906);
nor U13193 (N_13193,N_12843,N_12883);
nor U13194 (N_13194,N_12986,N_12853);
nor U13195 (N_13195,N_12865,N_12915);
nor U13196 (N_13196,N_12824,N_12826);
nand U13197 (N_13197,N_12923,N_12869);
xor U13198 (N_13198,N_12890,N_12911);
nor U13199 (N_13199,N_12934,N_12931);
and U13200 (N_13200,N_13017,N_13172);
nor U13201 (N_13201,N_13118,N_13151);
nand U13202 (N_13202,N_13163,N_13139);
xnor U13203 (N_13203,N_13137,N_13158);
and U13204 (N_13204,N_13079,N_13060);
nand U13205 (N_13205,N_13164,N_13083);
xor U13206 (N_13206,N_13180,N_13178);
and U13207 (N_13207,N_13111,N_13001);
and U13208 (N_13208,N_13073,N_13153);
nand U13209 (N_13209,N_13145,N_13182);
nand U13210 (N_13210,N_13088,N_13189);
and U13211 (N_13211,N_13062,N_13167);
or U13212 (N_13212,N_13121,N_13161);
nand U13213 (N_13213,N_13074,N_13106);
nand U13214 (N_13214,N_13039,N_13041);
or U13215 (N_13215,N_13067,N_13115);
and U13216 (N_13216,N_13091,N_13169);
nor U13217 (N_13217,N_13126,N_13096);
nor U13218 (N_13218,N_13036,N_13147);
nor U13219 (N_13219,N_13144,N_13000);
or U13220 (N_13220,N_13197,N_13141);
or U13221 (N_13221,N_13042,N_13176);
or U13222 (N_13222,N_13047,N_13069);
nor U13223 (N_13223,N_13045,N_13087);
and U13224 (N_13224,N_13011,N_13085);
or U13225 (N_13225,N_13092,N_13159);
and U13226 (N_13226,N_13123,N_13082);
and U13227 (N_13227,N_13077,N_13051);
xnor U13228 (N_13228,N_13008,N_13029);
xor U13229 (N_13229,N_13193,N_13136);
nand U13230 (N_13230,N_13099,N_13084);
and U13231 (N_13231,N_13095,N_13194);
nand U13232 (N_13232,N_13049,N_13196);
and U13233 (N_13233,N_13076,N_13005);
xor U13234 (N_13234,N_13179,N_13109);
or U13235 (N_13235,N_13059,N_13097);
xor U13236 (N_13236,N_13043,N_13192);
and U13237 (N_13237,N_13154,N_13038);
nor U13238 (N_13238,N_13015,N_13174);
xnor U13239 (N_13239,N_13021,N_13132);
nand U13240 (N_13240,N_13127,N_13177);
or U13241 (N_13241,N_13046,N_13168);
or U13242 (N_13242,N_13101,N_13064);
nand U13243 (N_13243,N_13171,N_13102);
or U13244 (N_13244,N_13034,N_13068);
nand U13245 (N_13245,N_13090,N_13048);
nand U13246 (N_13246,N_13198,N_13003);
nand U13247 (N_13247,N_13129,N_13185);
xor U13248 (N_13248,N_13070,N_13033);
and U13249 (N_13249,N_13071,N_13030);
or U13250 (N_13250,N_13012,N_13050);
nor U13251 (N_13251,N_13114,N_13055);
xnor U13252 (N_13252,N_13026,N_13009);
xor U13253 (N_13253,N_13103,N_13120);
nand U13254 (N_13254,N_13190,N_13010);
and U13255 (N_13255,N_13181,N_13130);
and U13256 (N_13256,N_13063,N_13066);
xnor U13257 (N_13257,N_13104,N_13122);
nor U13258 (N_13258,N_13173,N_13037);
nor U13259 (N_13259,N_13175,N_13072);
xnor U13260 (N_13260,N_13191,N_13150);
nand U13261 (N_13261,N_13162,N_13116);
or U13262 (N_13262,N_13032,N_13052);
or U13263 (N_13263,N_13149,N_13044);
xnor U13264 (N_13264,N_13094,N_13016);
xnor U13265 (N_13265,N_13157,N_13004);
xnor U13266 (N_13266,N_13143,N_13019);
and U13267 (N_13267,N_13022,N_13020);
or U13268 (N_13268,N_13142,N_13183);
nor U13269 (N_13269,N_13018,N_13089);
and U13270 (N_13270,N_13075,N_13093);
nand U13271 (N_13271,N_13006,N_13057);
nor U13272 (N_13272,N_13140,N_13187);
xnor U13273 (N_13273,N_13078,N_13113);
and U13274 (N_13274,N_13024,N_13119);
or U13275 (N_13275,N_13128,N_13013);
xnor U13276 (N_13276,N_13054,N_13014);
nor U13277 (N_13277,N_13061,N_13035);
nor U13278 (N_13278,N_13166,N_13135);
or U13279 (N_13279,N_13156,N_13138);
nor U13280 (N_13280,N_13028,N_13131);
nand U13281 (N_13281,N_13152,N_13065);
or U13282 (N_13282,N_13184,N_13040);
nand U13283 (N_13283,N_13160,N_13108);
and U13284 (N_13284,N_13025,N_13110);
or U13285 (N_13285,N_13100,N_13170);
xnor U13286 (N_13286,N_13002,N_13081);
nor U13287 (N_13287,N_13133,N_13165);
nor U13288 (N_13288,N_13098,N_13124);
xor U13289 (N_13289,N_13155,N_13105);
nor U13290 (N_13290,N_13186,N_13195);
or U13291 (N_13291,N_13027,N_13056);
nand U13292 (N_13292,N_13112,N_13117);
or U13293 (N_13293,N_13125,N_13146);
nor U13294 (N_13294,N_13053,N_13058);
nor U13295 (N_13295,N_13080,N_13007);
nand U13296 (N_13296,N_13107,N_13199);
or U13297 (N_13297,N_13188,N_13148);
or U13298 (N_13298,N_13134,N_13023);
nand U13299 (N_13299,N_13086,N_13031);
xnor U13300 (N_13300,N_13115,N_13182);
xnor U13301 (N_13301,N_13022,N_13115);
and U13302 (N_13302,N_13166,N_13026);
nor U13303 (N_13303,N_13161,N_13040);
or U13304 (N_13304,N_13085,N_13133);
nand U13305 (N_13305,N_13056,N_13033);
or U13306 (N_13306,N_13189,N_13041);
nand U13307 (N_13307,N_13196,N_13163);
nand U13308 (N_13308,N_13155,N_13122);
or U13309 (N_13309,N_13188,N_13035);
and U13310 (N_13310,N_13116,N_13156);
and U13311 (N_13311,N_13002,N_13192);
and U13312 (N_13312,N_13030,N_13121);
and U13313 (N_13313,N_13159,N_13024);
or U13314 (N_13314,N_13133,N_13160);
and U13315 (N_13315,N_13004,N_13179);
or U13316 (N_13316,N_13055,N_13006);
or U13317 (N_13317,N_13067,N_13151);
or U13318 (N_13318,N_13060,N_13006);
nor U13319 (N_13319,N_13038,N_13060);
xor U13320 (N_13320,N_13195,N_13103);
xnor U13321 (N_13321,N_13109,N_13115);
nor U13322 (N_13322,N_13194,N_13139);
nand U13323 (N_13323,N_13010,N_13073);
or U13324 (N_13324,N_13133,N_13009);
nor U13325 (N_13325,N_13072,N_13165);
or U13326 (N_13326,N_13064,N_13030);
nand U13327 (N_13327,N_13081,N_13155);
nor U13328 (N_13328,N_13149,N_13139);
xor U13329 (N_13329,N_13186,N_13087);
nor U13330 (N_13330,N_13071,N_13148);
and U13331 (N_13331,N_13185,N_13094);
nor U13332 (N_13332,N_13000,N_13026);
nor U13333 (N_13333,N_13167,N_13038);
nor U13334 (N_13334,N_13023,N_13033);
and U13335 (N_13335,N_13108,N_13145);
or U13336 (N_13336,N_13165,N_13027);
xor U13337 (N_13337,N_13118,N_13179);
and U13338 (N_13338,N_13176,N_13105);
or U13339 (N_13339,N_13039,N_13095);
nor U13340 (N_13340,N_13079,N_13075);
xnor U13341 (N_13341,N_13135,N_13150);
nor U13342 (N_13342,N_13047,N_13171);
and U13343 (N_13343,N_13197,N_13152);
nor U13344 (N_13344,N_13053,N_13039);
or U13345 (N_13345,N_13157,N_13174);
or U13346 (N_13346,N_13126,N_13162);
nor U13347 (N_13347,N_13113,N_13045);
or U13348 (N_13348,N_13058,N_13131);
nand U13349 (N_13349,N_13182,N_13124);
xor U13350 (N_13350,N_13038,N_13055);
xor U13351 (N_13351,N_13076,N_13187);
and U13352 (N_13352,N_13186,N_13102);
xnor U13353 (N_13353,N_13105,N_13016);
xor U13354 (N_13354,N_13178,N_13035);
nand U13355 (N_13355,N_13073,N_13004);
nand U13356 (N_13356,N_13065,N_13122);
or U13357 (N_13357,N_13199,N_13141);
nor U13358 (N_13358,N_13185,N_13186);
nand U13359 (N_13359,N_13094,N_13073);
and U13360 (N_13360,N_13147,N_13022);
and U13361 (N_13361,N_13096,N_13147);
xnor U13362 (N_13362,N_13141,N_13123);
or U13363 (N_13363,N_13167,N_13105);
xnor U13364 (N_13364,N_13000,N_13086);
or U13365 (N_13365,N_13154,N_13162);
and U13366 (N_13366,N_13080,N_13061);
nor U13367 (N_13367,N_13168,N_13076);
and U13368 (N_13368,N_13184,N_13056);
xnor U13369 (N_13369,N_13184,N_13014);
and U13370 (N_13370,N_13141,N_13149);
and U13371 (N_13371,N_13036,N_13027);
nor U13372 (N_13372,N_13186,N_13114);
or U13373 (N_13373,N_13172,N_13005);
and U13374 (N_13374,N_13098,N_13025);
nor U13375 (N_13375,N_13126,N_13103);
and U13376 (N_13376,N_13126,N_13052);
xor U13377 (N_13377,N_13108,N_13171);
and U13378 (N_13378,N_13073,N_13054);
nor U13379 (N_13379,N_13101,N_13181);
nand U13380 (N_13380,N_13005,N_13065);
and U13381 (N_13381,N_13141,N_13092);
xnor U13382 (N_13382,N_13138,N_13063);
and U13383 (N_13383,N_13092,N_13130);
xnor U13384 (N_13384,N_13020,N_13046);
nor U13385 (N_13385,N_13094,N_13191);
nor U13386 (N_13386,N_13130,N_13185);
nor U13387 (N_13387,N_13112,N_13120);
xor U13388 (N_13388,N_13032,N_13008);
nor U13389 (N_13389,N_13190,N_13093);
xor U13390 (N_13390,N_13122,N_13068);
nand U13391 (N_13391,N_13174,N_13145);
nand U13392 (N_13392,N_13071,N_13124);
or U13393 (N_13393,N_13010,N_13006);
and U13394 (N_13394,N_13065,N_13171);
nor U13395 (N_13395,N_13034,N_13137);
nand U13396 (N_13396,N_13048,N_13097);
xnor U13397 (N_13397,N_13127,N_13113);
or U13398 (N_13398,N_13060,N_13117);
xnor U13399 (N_13399,N_13113,N_13071);
nor U13400 (N_13400,N_13241,N_13237);
nand U13401 (N_13401,N_13243,N_13232);
nand U13402 (N_13402,N_13223,N_13257);
and U13403 (N_13403,N_13274,N_13212);
nand U13404 (N_13404,N_13305,N_13316);
and U13405 (N_13405,N_13272,N_13297);
or U13406 (N_13406,N_13326,N_13294);
xor U13407 (N_13407,N_13224,N_13354);
or U13408 (N_13408,N_13395,N_13310);
nand U13409 (N_13409,N_13377,N_13250);
nor U13410 (N_13410,N_13365,N_13235);
xor U13411 (N_13411,N_13315,N_13280);
and U13412 (N_13412,N_13393,N_13293);
or U13413 (N_13413,N_13277,N_13309);
xor U13414 (N_13414,N_13317,N_13286);
nand U13415 (N_13415,N_13343,N_13350);
nand U13416 (N_13416,N_13370,N_13281);
nand U13417 (N_13417,N_13225,N_13355);
and U13418 (N_13418,N_13245,N_13296);
xor U13419 (N_13419,N_13204,N_13353);
nor U13420 (N_13420,N_13288,N_13252);
xnor U13421 (N_13421,N_13383,N_13229);
xnor U13422 (N_13422,N_13319,N_13337);
xnor U13423 (N_13423,N_13398,N_13330);
nor U13424 (N_13424,N_13282,N_13234);
xor U13425 (N_13425,N_13262,N_13357);
xnor U13426 (N_13426,N_13363,N_13263);
xnor U13427 (N_13427,N_13338,N_13375);
nand U13428 (N_13428,N_13331,N_13248);
nor U13429 (N_13429,N_13356,N_13368);
and U13430 (N_13430,N_13372,N_13379);
xnor U13431 (N_13431,N_13351,N_13251);
and U13432 (N_13432,N_13240,N_13301);
nor U13433 (N_13433,N_13226,N_13246);
xor U13434 (N_13434,N_13266,N_13289);
nand U13435 (N_13435,N_13295,N_13244);
nor U13436 (N_13436,N_13347,N_13270);
and U13437 (N_13437,N_13340,N_13360);
and U13438 (N_13438,N_13218,N_13265);
and U13439 (N_13439,N_13376,N_13279);
xor U13440 (N_13440,N_13336,N_13221);
or U13441 (N_13441,N_13322,N_13371);
nor U13442 (N_13442,N_13346,N_13313);
nor U13443 (N_13443,N_13276,N_13390);
nand U13444 (N_13444,N_13230,N_13219);
xor U13445 (N_13445,N_13332,N_13238);
and U13446 (N_13446,N_13287,N_13222);
xor U13447 (N_13447,N_13200,N_13299);
xnor U13448 (N_13448,N_13284,N_13373);
nor U13449 (N_13449,N_13256,N_13311);
xnor U13450 (N_13450,N_13369,N_13359);
xor U13451 (N_13451,N_13324,N_13334);
xnor U13452 (N_13452,N_13308,N_13304);
or U13453 (N_13453,N_13307,N_13385);
or U13454 (N_13454,N_13278,N_13302);
nand U13455 (N_13455,N_13291,N_13389);
and U13456 (N_13456,N_13348,N_13202);
xnor U13457 (N_13457,N_13314,N_13341);
xor U13458 (N_13458,N_13211,N_13387);
nor U13459 (N_13459,N_13335,N_13358);
nand U13460 (N_13460,N_13327,N_13220);
or U13461 (N_13461,N_13328,N_13203);
nand U13462 (N_13462,N_13258,N_13349);
and U13463 (N_13463,N_13303,N_13259);
xor U13464 (N_13464,N_13207,N_13275);
nor U13465 (N_13465,N_13344,N_13397);
nand U13466 (N_13466,N_13228,N_13396);
xnor U13467 (N_13467,N_13333,N_13381);
nor U13468 (N_13468,N_13391,N_13271);
nand U13469 (N_13469,N_13283,N_13323);
nand U13470 (N_13470,N_13267,N_13364);
nand U13471 (N_13471,N_13210,N_13362);
xnor U13472 (N_13472,N_13386,N_13361);
or U13473 (N_13473,N_13269,N_13366);
nor U13474 (N_13474,N_13345,N_13233);
xor U13475 (N_13475,N_13249,N_13382);
nand U13476 (N_13476,N_13285,N_13206);
and U13477 (N_13477,N_13213,N_13378);
and U13478 (N_13478,N_13318,N_13321);
or U13479 (N_13479,N_13352,N_13253);
nand U13480 (N_13480,N_13261,N_13300);
nor U13481 (N_13481,N_13388,N_13216);
nor U13482 (N_13482,N_13306,N_13273);
nand U13483 (N_13483,N_13247,N_13205);
nor U13484 (N_13484,N_13342,N_13214);
and U13485 (N_13485,N_13380,N_13236);
or U13486 (N_13486,N_13399,N_13339);
nand U13487 (N_13487,N_13292,N_13392);
or U13488 (N_13488,N_13374,N_13254);
nand U13489 (N_13489,N_13264,N_13227);
nand U13490 (N_13490,N_13239,N_13312);
nor U13491 (N_13491,N_13384,N_13298);
or U13492 (N_13492,N_13268,N_13320);
nor U13493 (N_13493,N_13329,N_13394);
or U13494 (N_13494,N_13255,N_13217);
or U13495 (N_13495,N_13231,N_13325);
nor U13496 (N_13496,N_13215,N_13209);
and U13497 (N_13497,N_13201,N_13367);
nand U13498 (N_13498,N_13208,N_13260);
xor U13499 (N_13499,N_13290,N_13242);
nand U13500 (N_13500,N_13213,N_13290);
or U13501 (N_13501,N_13229,N_13243);
nand U13502 (N_13502,N_13392,N_13210);
or U13503 (N_13503,N_13202,N_13378);
xor U13504 (N_13504,N_13267,N_13202);
nor U13505 (N_13505,N_13207,N_13369);
nor U13506 (N_13506,N_13304,N_13247);
and U13507 (N_13507,N_13207,N_13367);
or U13508 (N_13508,N_13317,N_13222);
nor U13509 (N_13509,N_13335,N_13270);
or U13510 (N_13510,N_13353,N_13206);
nor U13511 (N_13511,N_13243,N_13203);
nand U13512 (N_13512,N_13393,N_13302);
nand U13513 (N_13513,N_13377,N_13283);
or U13514 (N_13514,N_13259,N_13299);
or U13515 (N_13515,N_13262,N_13375);
and U13516 (N_13516,N_13252,N_13316);
nand U13517 (N_13517,N_13292,N_13336);
nand U13518 (N_13518,N_13345,N_13273);
or U13519 (N_13519,N_13363,N_13355);
and U13520 (N_13520,N_13302,N_13341);
xor U13521 (N_13521,N_13240,N_13232);
and U13522 (N_13522,N_13336,N_13372);
or U13523 (N_13523,N_13396,N_13334);
or U13524 (N_13524,N_13319,N_13305);
xor U13525 (N_13525,N_13247,N_13200);
or U13526 (N_13526,N_13370,N_13277);
nor U13527 (N_13527,N_13371,N_13328);
nand U13528 (N_13528,N_13217,N_13399);
nand U13529 (N_13529,N_13249,N_13384);
or U13530 (N_13530,N_13346,N_13284);
or U13531 (N_13531,N_13367,N_13384);
or U13532 (N_13532,N_13317,N_13259);
and U13533 (N_13533,N_13380,N_13205);
or U13534 (N_13534,N_13374,N_13251);
or U13535 (N_13535,N_13322,N_13260);
xor U13536 (N_13536,N_13350,N_13331);
nor U13537 (N_13537,N_13256,N_13325);
nand U13538 (N_13538,N_13290,N_13214);
and U13539 (N_13539,N_13325,N_13239);
and U13540 (N_13540,N_13327,N_13308);
nor U13541 (N_13541,N_13300,N_13296);
or U13542 (N_13542,N_13271,N_13327);
nor U13543 (N_13543,N_13275,N_13287);
xnor U13544 (N_13544,N_13262,N_13330);
nand U13545 (N_13545,N_13237,N_13331);
xor U13546 (N_13546,N_13355,N_13258);
nor U13547 (N_13547,N_13220,N_13302);
xnor U13548 (N_13548,N_13288,N_13212);
xor U13549 (N_13549,N_13335,N_13219);
nand U13550 (N_13550,N_13235,N_13280);
nor U13551 (N_13551,N_13317,N_13299);
or U13552 (N_13552,N_13326,N_13271);
xor U13553 (N_13553,N_13384,N_13210);
nor U13554 (N_13554,N_13281,N_13287);
nand U13555 (N_13555,N_13219,N_13291);
or U13556 (N_13556,N_13270,N_13285);
nor U13557 (N_13557,N_13393,N_13214);
xnor U13558 (N_13558,N_13366,N_13289);
nor U13559 (N_13559,N_13256,N_13296);
nand U13560 (N_13560,N_13298,N_13278);
nand U13561 (N_13561,N_13363,N_13303);
xnor U13562 (N_13562,N_13359,N_13394);
or U13563 (N_13563,N_13227,N_13381);
or U13564 (N_13564,N_13246,N_13275);
and U13565 (N_13565,N_13292,N_13393);
or U13566 (N_13566,N_13321,N_13207);
nand U13567 (N_13567,N_13385,N_13354);
nor U13568 (N_13568,N_13220,N_13365);
nor U13569 (N_13569,N_13382,N_13324);
nand U13570 (N_13570,N_13200,N_13310);
nand U13571 (N_13571,N_13394,N_13323);
or U13572 (N_13572,N_13351,N_13277);
or U13573 (N_13573,N_13246,N_13234);
xor U13574 (N_13574,N_13368,N_13285);
nor U13575 (N_13575,N_13260,N_13333);
and U13576 (N_13576,N_13395,N_13313);
nand U13577 (N_13577,N_13280,N_13320);
and U13578 (N_13578,N_13204,N_13307);
and U13579 (N_13579,N_13330,N_13375);
nand U13580 (N_13580,N_13297,N_13204);
and U13581 (N_13581,N_13287,N_13252);
nor U13582 (N_13582,N_13374,N_13360);
xnor U13583 (N_13583,N_13278,N_13256);
xnor U13584 (N_13584,N_13343,N_13393);
xor U13585 (N_13585,N_13324,N_13289);
nor U13586 (N_13586,N_13242,N_13216);
nor U13587 (N_13587,N_13395,N_13382);
nor U13588 (N_13588,N_13207,N_13327);
xnor U13589 (N_13589,N_13394,N_13315);
and U13590 (N_13590,N_13209,N_13230);
and U13591 (N_13591,N_13351,N_13334);
and U13592 (N_13592,N_13225,N_13258);
xnor U13593 (N_13593,N_13243,N_13274);
nand U13594 (N_13594,N_13351,N_13212);
and U13595 (N_13595,N_13394,N_13321);
and U13596 (N_13596,N_13368,N_13217);
and U13597 (N_13597,N_13215,N_13284);
nor U13598 (N_13598,N_13382,N_13338);
nand U13599 (N_13599,N_13314,N_13242);
nor U13600 (N_13600,N_13422,N_13488);
and U13601 (N_13601,N_13432,N_13483);
xor U13602 (N_13602,N_13508,N_13489);
nand U13603 (N_13603,N_13474,N_13435);
and U13604 (N_13604,N_13498,N_13541);
nor U13605 (N_13605,N_13579,N_13490);
and U13606 (N_13606,N_13412,N_13537);
nand U13607 (N_13607,N_13589,N_13401);
xor U13608 (N_13608,N_13507,N_13462);
and U13609 (N_13609,N_13561,N_13469);
or U13610 (N_13610,N_13506,N_13487);
and U13611 (N_13611,N_13406,N_13492);
xor U13612 (N_13612,N_13529,N_13505);
xor U13613 (N_13613,N_13570,N_13598);
xor U13614 (N_13614,N_13468,N_13404);
or U13615 (N_13615,N_13517,N_13534);
or U13616 (N_13616,N_13554,N_13439);
nor U13617 (N_13617,N_13527,N_13512);
or U13618 (N_13618,N_13459,N_13580);
nor U13619 (N_13619,N_13495,N_13430);
or U13620 (N_13620,N_13592,N_13409);
nand U13621 (N_13621,N_13516,N_13450);
or U13622 (N_13622,N_13520,N_13472);
xor U13623 (N_13623,N_13445,N_13466);
xor U13624 (N_13624,N_13535,N_13560);
nand U13625 (N_13625,N_13440,N_13567);
nor U13626 (N_13626,N_13452,N_13577);
nand U13627 (N_13627,N_13426,N_13416);
and U13628 (N_13628,N_13475,N_13515);
nor U13629 (N_13629,N_13513,N_13509);
and U13630 (N_13630,N_13407,N_13429);
nand U13631 (N_13631,N_13478,N_13565);
xor U13632 (N_13632,N_13599,N_13420);
nor U13633 (N_13633,N_13413,N_13476);
nor U13634 (N_13634,N_13502,N_13411);
xnor U13635 (N_13635,N_13514,N_13403);
and U13636 (N_13636,N_13425,N_13482);
or U13637 (N_13637,N_13437,N_13595);
nand U13638 (N_13638,N_13551,N_13470);
xor U13639 (N_13639,N_13464,N_13456);
or U13640 (N_13640,N_13491,N_13446);
nand U13641 (N_13641,N_13451,N_13581);
nor U13642 (N_13642,N_13503,N_13461);
nand U13643 (N_13643,N_13547,N_13524);
or U13644 (N_13644,N_13557,N_13518);
nor U13645 (N_13645,N_13553,N_13572);
and U13646 (N_13646,N_13463,N_13571);
nand U13647 (N_13647,N_13415,N_13423);
and U13648 (N_13648,N_13428,N_13582);
or U13649 (N_13649,N_13528,N_13438);
and U13650 (N_13650,N_13418,N_13526);
nor U13651 (N_13651,N_13484,N_13583);
and U13652 (N_13652,N_13477,N_13596);
xnor U13653 (N_13653,N_13563,N_13540);
xor U13654 (N_13654,N_13419,N_13574);
nor U13655 (N_13655,N_13500,N_13555);
xor U13656 (N_13656,N_13447,N_13511);
xor U13657 (N_13657,N_13400,N_13575);
and U13658 (N_13658,N_13434,N_13442);
or U13659 (N_13659,N_13414,N_13441);
nor U13660 (N_13660,N_13473,N_13543);
nand U13661 (N_13661,N_13550,N_13467);
nand U13662 (N_13662,N_13471,N_13559);
nand U13663 (N_13663,N_13569,N_13402);
and U13664 (N_13664,N_13525,N_13530);
or U13665 (N_13665,N_13594,N_13427);
nor U13666 (N_13666,N_13539,N_13504);
nand U13667 (N_13667,N_13584,N_13501);
or U13668 (N_13668,N_13533,N_13458);
xnor U13669 (N_13669,N_13552,N_13497);
or U13670 (N_13670,N_13433,N_13522);
nand U13671 (N_13671,N_13573,N_13424);
nor U13672 (N_13672,N_13480,N_13556);
nand U13673 (N_13673,N_13597,N_13481);
nor U13674 (N_13674,N_13590,N_13443);
or U13675 (N_13675,N_13405,N_13593);
and U13676 (N_13676,N_13586,N_13521);
and U13677 (N_13677,N_13564,N_13531);
xor U13678 (N_13678,N_13465,N_13496);
or U13679 (N_13679,N_13460,N_13454);
and U13680 (N_13680,N_13548,N_13578);
or U13681 (N_13681,N_13431,N_13421);
nand U13682 (N_13682,N_13436,N_13449);
and U13683 (N_13683,N_13562,N_13455);
xor U13684 (N_13684,N_13493,N_13566);
and U13685 (N_13685,N_13417,N_13549);
or U13686 (N_13686,N_13494,N_13510);
nand U13687 (N_13687,N_13546,N_13536);
nor U13688 (N_13688,N_13519,N_13558);
nor U13689 (N_13689,N_13457,N_13486);
nor U13690 (N_13690,N_13542,N_13485);
or U13691 (N_13691,N_13453,N_13448);
or U13692 (N_13692,N_13479,N_13568);
nand U13693 (N_13693,N_13576,N_13444);
and U13694 (N_13694,N_13410,N_13591);
and U13695 (N_13695,N_13585,N_13538);
nor U13696 (N_13696,N_13408,N_13545);
nor U13697 (N_13697,N_13587,N_13499);
and U13698 (N_13698,N_13532,N_13523);
or U13699 (N_13699,N_13544,N_13588);
or U13700 (N_13700,N_13487,N_13415);
nand U13701 (N_13701,N_13516,N_13429);
nand U13702 (N_13702,N_13589,N_13499);
or U13703 (N_13703,N_13424,N_13545);
and U13704 (N_13704,N_13417,N_13441);
and U13705 (N_13705,N_13583,N_13496);
or U13706 (N_13706,N_13456,N_13427);
and U13707 (N_13707,N_13561,N_13424);
nand U13708 (N_13708,N_13416,N_13482);
or U13709 (N_13709,N_13592,N_13501);
xnor U13710 (N_13710,N_13569,N_13416);
xor U13711 (N_13711,N_13411,N_13424);
or U13712 (N_13712,N_13574,N_13579);
or U13713 (N_13713,N_13487,N_13485);
xor U13714 (N_13714,N_13596,N_13591);
and U13715 (N_13715,N_13502,N_13480);
nand U13716 (N_13716,N_13553,N_13417);
and U13717 (N_13717,N_13454,N_13421);
or U13718 (N_13718,N_13432,N_13438);
and U13719 (N_13719,N_13490,N_13563);
nor U13720 (N_13720,N_13545,N_13434);
or U13721 (N_13721,N_13527,N_13400);
or U13722 (N_13722,N_13406,N_13504);
or U13723 (N_13723,N_13550,N_13452);
nor U13724 (N_13724,N_13590,N_13497);
and U13725 (N_13725,N_13532,N_13480);
and U13726 (N_13726,N_13426,N_13462);
or U13727 (N_13727,N_13559,N_13486);
and U13728 (N_13728,N_13475,N_13471);
and U13729 (N_13729,N_13561,N_13451);
nor U13730 (N_13730,N_13418,N_13596);
xnor U13731 (N_13731,N_13469,N_13427);
xor U13732 (N_13732,N_13547,N_13477);
and U13733 (N_13733,N_13421,N_13580);
and U13734 (N_13734,N_13536,N_13521);
nor U13735 (N_13735,N_13593,N_13534);
xnor U13736 (N_13736,N_13402,N_13416);
xor U13737 (N_13737,N_13405,N_13453);
and U13738 (N_13738,N_13428,N_13538);
nand U13739 (N_13739,N_13524,N_13417);
or U13740 (N_13740,N_13497,N_13442);
nor U13741 (N_13741,N_13536,N_13401);
and U13742 (N_13742,N_13556,N_13566);
xor U13743 (N_13743,N_13411,N_13485);
nor U13744 (N_13744,N_13503,N_13530);
and U13745 (N_13745,N_13457,N_13511);
nor U13746 (N_13746,N_13451,N_13541);
nand U13747 (N_13747,N_13469,N_13522);
or U13748 (N_13748,N_13505,N_13484);
xor U13749 (N_13749,N_13499,N_13572);
and U13750 (N_13750,N_13451,N_13402);
xor U13751 (N_13751,N_13580,N_13511);
nor U13752 (N_13752,N_13553,N_13594);
nor U13753 (N_13753,N_13429,N_13538);
nand U13754 (N_13754,N_13419,N_13513);
nand U13755 (N_13755,N_13511,N_13520);
or U13756 (N_13756,N_13504,N_13536);
and U13757 (N_13757,N_13517,N_13427);
and U13758 (N_13758,N_13490,N_13516);
and U13759 (N_13759,N_13407,N_13493);
xor U13760 (N_13760,N_13475,N_13550);
xor U13761 (N_13761,N_13507,N_13588);
xnor U13762 (N_13762,N_13552,N_13504);
nand U13763 (N_13763,N_13486,N_13494);
and U13764 (N_13764,N_13439,N_13454);
and U13765 (N_13765,N_13538,N_13500);
or U13766 (N_13766,N_13455,N_13449);
or U13767 (N_13767,N_13506,N_13541);
nor U13768 (N_13768,N_13447,N_13403);
and U13769 (N_13769,N_13420,N_13435);
and U13770 (N_13770,N_13572,N_13458);
xor U13771 (N_13771,N_13502,N_13570);
and U13772 (N_13772,N_13593,N_13501);
xnor U13773 (N_13773,N_13430,N_13523);
and U13774 (N_13774,N_13509,N_13479);
and U13775 (N_13775,N_13526,N_13538);
xor U13776 (N_13776,N_13584,N_13407);
nor U13777 (N_13777,N_13546,N_13408);
and U13778 (N_13778,N_13455,N_13441);
and U13779 (N_13779,N_13453,N_13551);
nor U13780 (N_13780,N_13561,N_13458);
and U13781 (N_13781,N_13505,N_13434);
nand U13782 (N_13782,N_13415,N_13570);
nor U13783 (N_13783,N_13530,N_13468);
and U13784 (N_13784,N_13516,N_13428);
or U13785 (N_13785,N_13495,N_13406);
xor U13786 (N_13786,N_13479,N_13455);
or U13787 (N_13787,N_13462,N_13491);
nor U13788 (N_13788,N_13482,N_13503);
xnor U13789 (N_13789,N_13500,N_13415);
nor U13790 (N_13790,N_13484,N_13478);
nand U13791 (N_13791,N_13585,N_13418);
nor U13792 (N_13792,N_13499,N_13500);
nor U13793 (N_13793,N_13517,N_13557);
nor U13794 (N_13794,N_13431,N_13500);
or U13795 (N_13795,N_13490,N_13476);
or U13796 (N_13796,N_13466,N_13517);
nor U13797 (N_13797,N_13438,N_13454);
xnor U13798 (N_13798,N_13559,N_13495);
nand U13799 (N_13799,N_13578,N_13573);
nand U13800 (N_13800,N_13790,N_13786);
or U13801 (N_13801,N_13606,N_13727);
xnor U13802 (N_13802,N_13646,N_13741);
or U13803 (N_13803,N_13629,N_13749);
nand U13804 (N_13804,N_13753,N_13695);
nor U13805 (N_13805,N_13623,N_13783);
xor U13806 (N_13806,N_13723,N_13674);
and U13807 (N_13807,N_13728,N_13720);
nor U13808 (N_13808,N_13784,N_13652);
or U13809 (N_13809,N_13611,N_13719);
or U13810 (N_13810,N_13656,N_13733);
xor U13811 (N_13811,N_13613,N_13602);
and U13812 (N_13812,N_13707,N_13673);
nand U13813 (N_13813,N_13600,N_13792);
nor U13814 (N_13814,N_13654,N_13717);
nor U13815 (N_13815,N_13650,N_13740);
or U13816 (N_13816,N_13761,N_13665);
xnor U13817 (N_13817,N_13730,N_13678);
and U13818 (N_13818,N_13704,N_13752);
nand U13819 (N_13819,N_13735,N_13605);
or U13820 (N_13820,N_13635,N_13785);
nor U13821 (N_13821,N_13725,N_13647);
xor U13822 (N_13822,N_13660,N_13697);
xor U13823 (N_13823,N_13690,N_13636);
nor U13824 (N_13824,N_13743,N_13758);
and U13825 (N_13825,N_13683,N_13769);
nor U13826 (N_13826,N_13661,N_13764);
or U13827 (N_13827,N_13700,N_13778);
nor U13828 (N_13828,N_13767,N_13676);
and U13829 (N_13829,N_13742,N_13655);
xor U13830 (N_13830,N_13691,N_13619);
and U13831 (N_13831,N_13601,N_13737);
nand U13832 (N_13832,N_13639,N_13696);
and U13833 (N_13833,N_13625,N_13620);
and U13834 (N_13834,N_13750,N_13645);
or U13835 (N_13835,N_13771,N_13603);
nor U13836 (N_13836,N_13713,N_13644);
xor U13837 (N_13837,N_13712,N_13662);
or U13838 (N_13838,N_13618,N_13773);
xnor U13839 (N_13839,N_13687,N_13608);
xor U13840 (N_13840,N_13798,N_13693);
nor U13841 (N_13841,N_13616,N_13666);
or U13842 (N_13842,N_13780,N_13711);
and U13843 (N_13843,N_13765,N_13757);
nand U13844 (N_13844,N_13682,N_13722);
xor U13845 (N_13845,N_13747,N_13714);
nor U13846 (N_13846,N_13793,N_13795);
or U13847 (N_13847,N_13788,N_13648);
and U13848 (N_13848,N_13659,N_13726);
or U13849 (N_13849,N_13679,N_13718);
nor U13850 (N_13850,N_13776,N_13705);
and U13851 (N_13851,N_13781,N_13689);
nand U13852 (N_13852,N_13617,N_13703);
or U13853 (N_13853,N_13710,N_13754);
nand U13854 (N_13854,N_13732,N_13751);
nor U13855 (N_13855,N_13643,N_13614);
nand U13856 (N_13856,N_13663,N_13729);
or U13857 (N_13857,N_13615,N_13685);
or U13858 (N_13858,N_13692,N_13760);
and U13859 (N_13859,N_13734,N_13649);
nor U13860 (N_13860,N_13799,N_13738);
or U13861 (N_13861,N_13634,N_13797);
or U13862 (N_13862,N_13671,N_13770);
or U13863 (N_13863,N_13657,N_13624);
or U13864 (N_13864,N_13622,N_13702);
xor U13865 (N_13865,N_13664,N_13604);
xnor U13866 (N_13866,N_13610,N_13774);
nand U13867 (N_13867,N_13746,N_13745);
and U13868 (N_13868,N_13791,N_13653);
nand U13869 (N_13869,N_13759,N_13609);
xnor U13870 (N_13870,N_13768,N_13724);
nand U13871 (N_13871,N_13675,N_13755);
or U13872 (N_13872,N_13607,N_13736);
nor U13873 (N_13873,N_13677,N_13744);
nor U13874 (N_13874,N_13694,N_13688);
and U13875 (N_13875,N_13638,N_13762);
and U13876 (N_13876,N_13640,N_13698);
or U13877 (N_13877,N_13651,N_13716);
or U13878 (N_13878,N_13642,N_13630);
or U13879 (N_13879,N_13739,N_13701);
or U13880 (N_13880,N_13756,N_13748);
nand U13881 (N_13881,N_13721,N_13779);
or U13882 (N_13882,N_13627,N_13680);
and U13883 (N_13883,N_13628,N_13668);
nor U13884 (N_13884,N_13626,N_13777);
or U13885 (N_13885,N_13612,N_13709);
nand U13886 (N_13886,N_13672,N_13708);
nand U13887 (N_13887,N_13686,N_13731);
nor U13888 (N_13888,N_13796,N_13681);
nand U13889 (N_13889,N_13782,N_13772);
and U13890 (N_13890,N_13766,N_13669);
or U13891 (N_13891,N_13775,N_13763);
xor U13892 (N_13892,N_13715,N_13637);
xnor U13893 (N_13893,N_13684,N_13794);
xnor U13894 (N_13894,N_13670,N_13632);
and U13895 (N_13895,N_13667,N_13706);
and U13896 (N_13896,N_13699,N_13621);
nand U13897 (N_13897,N_13631,N_13787);
nand U13898 (N_13898,N_13658,N_13789);
or U13899 (N_13899,N_13633,N_13641);
and U13900 (N_13900,N_13606,N_13682);
nand U13901 (N_13901,N_13667,N_13775);
and U13902 (N_13902,N_13652,N_13726);
nand U13903 (N_13903,N_13791,N_13681);
or U13904 (N_13904,N_13650,N_13731);
nand U13905 (N_13905,N_13746,N_13680);
and U13906 (N_13906,N_13662,N_13606);
and U13907 (N_13907,N_13774,N_13673);
or U13908 (N_13908,N_13676,N_13776);
and U13909 (N_13909,N_13719,N_13742);
nand U13910 (N_13910,N_13622,N_13600);
xor U13911 (N_13911,N_13614,N_13759);
nand U13912 (N_13912,N_13728,N_13608);
or U13913 (N_13913,N_13747,N_13791);
nand U13914 (N_13914,N_13618,N_13602);
nor U13915 (N_13915,N_13657,N_13604);
or U13916 (N_13916,N_13710,N_13773);
or U13917 (N_13917,N_13715,N_13692);
and U13918 (N_13918,N_13756,N_13715);
and U13919 (N_13919,N_13761,N_13740);
nor U13920 (N_13920,N_13697,N_13741);
xor U13921 (N_13921,N_13712,N_13673);
xnor U13922 (N_13922,N_13773,N_13707);
nor U13923 (N_13923,N_13620,N_13788);
nand U13924 (N_13924,N_13675,N_13728);
nor U13925 (N_13925,N_13764,N_13666);
nand U13926 (N_13926,N_13623,N_13645);
xnor U13927 (N_13927,N_13735,N_13760);
and U13928 (N_13928,N_13721,N_13651);
or U13929 (N_13929,N_13685,N_13655);
or U13930 (N_13930,N_13606,N_13702);
nor U13931 (N_13931,N_13741,N_13691);
nand U13932 (N_13932,N_13612,N_13613);
or U13933 (N_13933,N_13659,N_13685);
nor U13934 (N_13934,N_13733,N_13696);
or U13935 (N_13935,N_13775,N_13627);
and U13936 (N_13936,N_13785,N_13651);
and U13937 (N_13937,N_13694,N_13608);
nor U13938 (N_13938,N_13754,N_13650);
nor U13939 (N_13939,N_13615,N_13664);
nor U13940 (N_13940,N_13694,N_13652);
and U13941 (N_13941,N_13665,N_13745);
nor U13942 (N_13942,N_13690,N_13633);
xor U13943 (N_13943,N_13696,N_13603);
and U13944 (N_13944,N_13753,N_13732);
nor U13945 (N_13945,N_13661,N_13623);
and U13946 (N_13946,N_13783,N_13664);
or U13947 (N_13947,N_13623,N_13641);
and U13948 (N_13948,N_13643,N_13628);
and U13949 (N_13949,N_13725,N_13716);
nor U13950 (N_13950,N_13740,N_13757);
nand U13951 (N_13951,N_13741,N_13730);
and U13952 (N_13952,N_13615,N_13768);
or U13953 (N_13953,N_13621,N_13623);
or U13954 (N_13954,N_13646,N_13784);
and U13955 (N_13955,N_13686,N_13685);
and U13956 (N_13956,N_13793,N_13799);
xor U13957 (N_13957,N_13777,N_13650);
or U13958 (N_13958,N_13648,N_13790);
nand U13959 (N_13959,N_13794,N_13775);
xor U13960 (N_13960,N_13657,N_13630);
or U13961 (N_13961,N_13703,N_13719);
nand U13962 (N_13962,N_13720,N_13719);
xnor U13963 (N_13963,N_13688,N_13658);
nor U13964 (N_13964,N_13746,N_13760);
nor U13965 (N_13965,N_13718,N_13723);
xnor U13966 (N_13966,N_13795,N_13654);
or U13967 (N_13967,N_13743,N_13682);
nor U13968 (N_13968,N_13698,N_13772);
nand U13969 (N_13969,N_13636,N_13677);
xor U13970 (N_13970,N_13697,N_13785);
nand U13971 (N_13971,N_13736,N_13648);
xor U13972 (N_13972,N_13679,N_13796);
xnor U13973 (N_13973,N_13651,N_13622);
xnor U13974 (N_13974,N_13746,N_13718);
and U13975 (N_13975,N_13670,N_13797);
nor U13976 (N_13976,N_13717,N_13758);
nand U13977 (N_13977,N_13624,N_13654);
or U13978 (N_13978,N_13644,N_13664);
or U13979 (N_13979,N_13644,N_13603);
xnor U13980 (N_13980,N_13663,N_13758);
or U13981 (N_13981,N_13736,N_13692);
nand U13982 (N_13982,N_13654,N_13636);
nor U13983 (N_13983,N_13735,N_13732);
and U13984 (N_13984,N_13613,N_13733);
or U13985 (N_13985,N_13635,N_13768);
xor U13986 (N_13986,N_13603,N_13683);
nor U13987 (N_13987,N_13727,N_13710);
nor U13988 (N_13988,N_13677,N_13795);
xor U13989 (N_13989,N_13664,N_13762);
nor U13990 (N_13990,N_13748,N_13602);
nand U13991 (N_13991,N_13775,N_13603);
xor U13992 (N_13992,N_13618,N_13669);
nand U13993 (N_13993,N_13779,N_13675);
or U13994 (N_13994,N_13652,N_13772);
xnor U13995 (N_13995,N_13755,N_13746);
xor U13996 (N_13996,N_13775,N_13772);
nor U13997 (N_13997,N_13712,N_13627);
xnor U13998 (N_13998,N_13632,N_13601);
or U13999 (N_13999,N_13748,N_13688);
or U14000 (N_14000,N_13866,N_13835);
nand U14001 (N_14001,N_13906,N_13935);
nor U14002 (N_14002,N_13887,N_13910);
and U14003 (N_14003,N_13991,N_13878);
nor U14004 (N_14004,N_13972,N_13955);
nand U14005 (N_14005,N_13858,N_13947);
or U14006 (N_14006,N_13949,N_13933);
or U14007 (N_14007,N_13822,N_13813);
xor U14008 (N_14008,N_13953,N_13876);
and U14009 (N_14009,N_13980,N_13862);
and U14010 (N_14010,N_13979,N_13860);
or U14011 (N_14011,N_13803,N_13809);
or U14012 (N_14012,N_13936,N_13856);
or U14013 (N_14013,N_13994,N_13962);
nand U14014 (N_14014,N_13900,N_13837);
and U14015 (N_14015,N_13896,N_13913);
or U14016 (N_14016,N_13880,N_13873);
nand U14017 (N_14017,N_13865,N_13969);
nand U14018 (N_14018,N_13902,N_13937);
nor U14019 (N_14019,N_13911,N_13893);
nand U14020 (N_14020,N_13990,N_13855);
nor U14021 (N_14021,N_13874,N_13807);
or U14022 (N_14022,N_13829,N_13879);
nor U14023 (N_14023,N_13869,N_13812);
and U14024 (N_14024,N_13882,N_13989);
xor U14025 (N_14025,N_13877,N_13982);
or U14026 (N_14026,N_13944,N_13908);
xnor U14027 (N_14027,N_13864,N_13888);
or U14028 (N_14028,N_13828,N_13915);
or U14029 (N_14029,N_13988,N_13857);
nand U14030 (N_14030,N_13974,N_13904);
and U14031 (N_14031,N_13886,N_13965);
xor U14032 (N_14032,N_13917,N_13931);
xor U14033 (N_14033,N_13916,N_13832);
xor U14034 (N_14034,N_13814,N_13872);
xnor U14035 (N_14035,N_13836,N_13957);
or U14036 (N_14036,N_13901,N_13859);
and U14037 (N_14037,N_13995,N_13960);
and U14038 (N_14038,N_13800,N_13889);
nor U14039 (N_14039,N_13824,N_13970);
xor U14040 (N_14040,N_13940,N_13923);
or U14041 (N_14041,N_13964,N_13843);
nand U14042 (N_14042,N_13976,N_13847);
nor U14043 (N_14043,N_13881,N_13833);
or U14044 (N_14044,N_13986,N_13998);
nor U14045 (N_14045,N_13918,N_13909);
nor U14046 (N_14046,N_13884,N_13852);
nor U14047 (N_14047,N_13867,N_13892);
or U14048 (N_14048,N_13977,N_13929);
or U14049 (N_14049,N_13871,N_13930);
or U14050 (N_14050,N_13959,N_13820);
nand U14051 (N_14051,N_13932,N_13823);
xnor U14052 (N_14052,N_13868,N_13985);
and U14053 (N_14053,N_13842,N_13973);
xnor U14054 (N_14054,N_13815,N_13920);
nor U14055 (N_14055,N_13841,N_13897);
or U14056 (N_14056,N_13907,N_13961);
xnor U14057 (N_14057,N_13895,N_13848);
and U14058 (N_14058,N_13952,N_13921);
xor U14059 (N_14059,N_13950,N_13826);
nor U14060 (N_14060,N_13846,N_13967);
nor U14061 (N_14061,N_13924,N_13899);
nand U14062 (N_14062,N_13999,N_13870);
or U14063 (N_14063,N_13840,N_13975);
xnor U14064 (N_14064,N_13958,N_13861);
xnor U14065 (N_14065,N_13928,N_13968);
and U14066 (N_14066,N_13898,N_13997);
nand U14067 (N_14067,N_13853,N_13905);
or U14068 (N_14068,N_13926,N_13922);
or U14069 (N_14069,N_13983,N_13802);
nor U14070 (N_14070,N_13943,N_13831);
nand U14071 (N_14071,N_13939,N_13816);
and U14072 (N_14072,N_13817,N_13844);
and U14073 (N_14073,N_13992,N_13914);
or U14074 (N_14074,N_13850,N_13963);
nor U14075 (N_14075,N_13805,N_13891);
nor U14076 (N_14076,N_13938,N_13821);
nor U14077 (N_14077,N_13927,N_13954);
or U14078 (N_14078,N_13801,N_13942);
nor U14079 (N_14079,N_13854,N_13948);
or U14080 (N_14080,N_13984,N_13811);
nor U14081 (N_14081,N_13981,N_13806);
nand U14082 (N_14082,N_13941,N_13808);
or U14083 (N_14083,N_13925,N_13919);
or U14084 (N_14084,N_13978,N_13912);
nor U14085 (N_14085,N_13956,N_13903);
and U14086 (N_14086,N_13934,N_13883);
nor U14087 (N_14087,N_13834,N_13830);
or U14088 (N_14088,N_13825,N_13827);
nand U14089 (N_14089,N_13951,N_13971);
xnor U14090 (N_14090,N_13804,N_13863);
xnor U14091 (N_14091,N_13851,N_13819);
or U14092 (N_14092,N_13890,N_13987);
or U14093 (N_14093,N_13945,N_13946);
and U14094 (N_14094,N_13818,N_13839);
nand U14095 (N_14095,N_13810,N_13996);
xnor U14096 (N_14096,N_13838,N_13993);
nand U14097 (N_14097,N_13966,N_13845);
nand U14098 (N_14098,N_13885,N_13849);
and U14099 (N_14099,N_13894,N_13875);
xnor U14100 (N_14100,N_13978,N_13888);
and U14101 (N_14101,N_13843,N_13968);
or U14102 (N_14102,N_13879,N_13972);
and U14103 (N_14103,N_13898,N_13811);
xnor U14104 (N_14104,N_13820,N_13925);
and U14105 (N_14105,N_13951,N_13839);
and U14106 (N_14106,N_13819,N_13977);
or U14107 (N_14107,N_13805,N_13968);
xor U14108 (N_14108,N_13917,N_13958);
nor U14109 (N_14109,N_13832,N_13824);
or U14110 (N_14110,N_13901,N_13825);
nor U14111 (N_14111,N_13923,N_13948);
nor U14112 (N_14112,N_13876,N_13862);
nand U14113 (N_14113,N_13960,N_13863);
or U14114 (N_14114,N_13837,N_13929);
nand U14115 (N_14115,N_13905,N_13833);
xnor U14116 (N_14116,N_13925,N_13842);
nand U14117 (N_14117,N_13928,N_13923);
nand U14118 (N_14118,N_13913,N_13997);
nor U14119 (N_14119,N_13842,N_13876);
xor U14120 (N_14120,N_13985,N_13827);
and U14121 (N_14121,N_13925,N_13931);
or U14122 (N_14122,N_13969,N_13872);
nor U14123 (N_14123,N_13814,N_13893);
or U14124 (N_14124,N_13966,N_13943);
xnor U14125 (N_14125,N_13803,N_13841);
and U14126 (N_14126,N_13887,N_13923);
nor U14127 (N_14127,N_13940,N_13885);
or U14128 (N_14128,N_13924,N_13988);
xor U14129 (N_14129,N_13940,N_13891);
xor U14130 (N_14130,N_13814,N_13958);
nor U14131 (N_14131,N_13820,N_13821);
nand U14132 (N_14132,N_13890,N_13896);
xnor U14133 (N_14133,N_13892,N_13861);
and U14134 (N_14134,N_13985,N_13844);
xor U14135 (N_14135,N_13979,N_13852);
nand U14136 (N_14136,N_13825,N_13932);
nand U14137 (N_14137,N_13802,N_13990);
xor U14138 (N_14138,N_13958,N_13835);
and U14139 (N_14139,N_13806,N_13863);
nand U14140 (N_14140,N_13865,N_13838);
xnor U14141 (N_14141,N_13812,N_13906);
or U14142 (N_14142,N_13989,N_13828);
and U14143 (N_14143,N_13921,N_13879);
nand U14144 (N_14144,N_13929,N_13815);
or U14145 (N_14145,N_13897,N_13800);
and U14146 (N_14146,N_13964,N_13846);
xnor U14147 (N_14147,N_13930,N_13893);
xnor U14148 (N_14148,N_13994,N_13922);
xnor U14149 (N_14149,N_13822,N_13820);
xnor U14150 (N_14150,N_13868,N_13943);
xor U14151 (N_14151,N_13846,N_13848);
xor U14152 (N_14152,N_13984,N_13829);
nor U14153 (N_14153,N_13995,N_13861);
nand U14154 (N_14154,N_13933,N_13953);
and U14155 (N_14155,N_13904,N_13953);
nor U14156 (N_14156,N_13957,N_13969);
and U14157 (N_14157,N_13852,N_13837);
nand U14158 (N_14158,N_13916,N_13977);
xor U14159 (N_14159,N_13828,N_13809);
and U14160 (N_14160,N_13827,N_13861);
nor U14161 (N_14161,N_13816,N_13837);
or U14162 (N_14162,N_13977,N_13902);
nand U14163 (N_14163,N_13907,N_13923);
nand U14164 (N_14164,N_13925,N_13800);
nor U14165 (N_14165,N_13909,N_13910);
xnor U14166 (N_14166,N_13995,N_13880);
nor U14167 (N_14167,N_13901,N_13873);
or U14168 (N_14168,N_13864,N_13877);
xor U14169 (N_14169,N_13995,N_13818);
and U14170 (N_14170,N_13959,N_13937);
nor U14171 (N_14171,N_13822,N_13927);
nor U14172 (N_14172,N_13814,N_13875);
xor U14173 (N_14173,N_13999,N_13961);
nand U14174 (N_14174,N_13880,N_13897);
or U14175 (N_14175,N_13924,N_13856);
xor U14176 (N_14176,N_13850,N_13924);
xnor U14177 (N_14177,N_13846,N_13913);
nor U14178 (N_14178,N_13904,N_13834);
nor U14179 (N_14179,N_13814,N_13867);
nor U14180 (N_14180,N_13802,N_13870);
nor U14181 (N_14181,N_13852,N_13964);
nor U14182 (N_14182,N_13971,N_13849);
nand U14183 (N_14183,N_13829,N_13863);
xor U14184 (N_14184,N_13826,N_13926);
xnor U14185 (N_14185,N_13846,N_13898);
and U14186 (N_14186,N_13969,N_13976);
nor U14187 (N_14187,N_13879,N_13903);
nor U14188 (N_14188,N_13990,N_13826);
nor U14189 (N_14189,N_13899,N_13987);
or U14190 (N_14190,N_13928,N_13880);
and U14191 (N_14191,N_13984,N_13953);
nor U14192 (N_14192,N_13852,N_13871);
nor U14193 (N_14193,N_13817,N_13893);
xnor U14194 (N_14194,N_13861,N_13884);
or U14195 (N_14195,N_13939,N_13837);
and U14196 (N_14196,N_13938,N_13904);
xnor U14197 (N_14197,N_13950,N_13942);
and U14198 (N_14198,N_13818,N_13848);
nand U14199 (N_14199,N_13819,N_13995);
nor U14200 (N_14200,N_14070,N_14054);
nor U14201 (N_14201,N_14082,N_14081);
or U14202 (N_14202,N_14022,N_14020);
xnor U14203 (N_14203,N_14125,N_14103);
nor U14204 (N_14204,N_14027,N_14132);
or U14205 (N_14205,N_14000,N_14075);
or U14206 (N_14206,N_14138,N_14071);
xnor U14207 (N_14207,N_14056,N_14151);
nand U14208 (N_14208,N_14077,N_14120);
nand U14209 (N_14209,N_14042,N_14137);
or U14210 (N_14210,N_14154,N_14113);
xor U14211 (N_14211,N_14044,N_14096);
xnor U14212 (N_14212,N_14122,N_14017);
xnor U14213 (N_14213,N_14085,N_14074);
and U14214 (N_14214,N_14139,N_14136);
nor U14215 (N_14215,N_14172,N_14186);
and U14216 (N_14216,N_14062,N_14149);
xnor U14217 (N_14217,N_14018,N_14049);
xnor U14218 (N_14218,N_14182,N_14058);
nor U14219 (N_14219,N_14097,N_14107);
and U14220 (N_14220,N_14142,N_14194);
xnor U14221 (N_14221,N_14073,N_14173);
xor U14222 (N_14222,N_14144,N_14159);
and U14223 (N_14223,N_14087,N_14008);
nand U14224 (N_14224,N_14118,N_14199);
xnor U14225 (N_14225,N_14140,N_14175);
nor U14226 (N_14226,N_14197,N_14048);
or U14227 (N_14227,N_14162,N_14038);
nand U14228 (N_14228,N_14116,N_14148);
nand U14229 (N_14229,N_14080,N_14112);
xor U14230 (N_14230,N_14036,N_14191);
nor U14231 (N_14231,N_14164,N_14127);
nand U14232 (N_14232,N_14009,N_14089);
and U14233 (N_14233,N_14052,N_14179);
xor U14234 (N_14234,N_14043,N_14066);
xnor U14235 (N_14235,N_14180,N_14196);
nand U14236 (N_14236,N_14030,N_14079);
and U14237 (N_14237,N_14006,N_14057);
nand U14238 (N_14238,N_14005,N_14069);
or U14239 (N_14239,N_14126,N_14152);
nor U14240 (N_14240,N_14101,N_14031);
or U14241 (N_14241,N_14021,N_14195);
nor U14242 (N_14242,N_14192,N_14121);
nand U14243 (N_14243,N_14061,N_14090);
nor U14244 (N_14244,N_14059,N_14165);
nand U14245 (N_14245,N_14041,N_14032);
and U14246 (N_14246,N_14171,N_14166);
xnor U14247 (N_14247,N_14010,N_14190);
nor U14248 (N_14248,N_14123,N_14067);
xnor U14249 (N_14249,N_14146,N_14007);
xor U14250 (N_14250,N_14039,N_14093);
nor U14251 (N_14251,N_14115,N_14108);
nor U14252 (N_14252,N_14037,N_14011);
nor U14253 (N_14253,N_14019,N_14014);
or U14254 (N_14254,N_14117,N_14034);
or U14255 (N_14255,N_14084,N_14178);
nand U14256 (N_14256,N_14029,N_14040);
or U14257 (N_14257,N_14102,N_14114);
nor U14258 (N_14258,N_14033,N_14076);
xnor U14259 (N_14259,N_14092,N_14198);
nand U14260 (N_14260,N_14060,N_14012);
and U14261 (N_14261,N_14083,N_14193);
nand U14262 (N_14262,N_14141,N_14187);
nor U14263 (N_14263,N_14065,N_14174);
and U14264 (N_14264,N_14156,N_14153);
nand U14265 (N_14265,N_14001,N_14072);
nor U14266 (N_14266,N_14150,N_14003);
nand U14267 (N_14267,N_14086,N_14104);
or U14268 (N_14268,N_14157,N_14185);
and U14269 (N_14269,N_14002,N_14013);
and U14270 (N_14270,N_14133,N_14028);
or U14271 (N_14271,N_14068,N_14091);
and U14272 (N_14272,N_14099,N_14169);
nor U14273 (N_14273,N_14158,N_14045);
xor U14274 (N_14274,N_14064,N_14105);
or U14275 (N_14275,N_14168,N_14109);
or U14276 (N_14276,N_14119,N_14177);
nand U14277 (N_14277,N_14094,N_14035);
nor U14278 (N_14278,N_14161,N_14163);
nor U14279 (N_14279,N_14095,N_14189);
nand U14280 (N_14280,N_14015,N_14025);
nor U14281 (N_14281,N_14134,N_14026);
or U14282 (N_14282,N_14131,N_14130);
xnor U14283 (N_14283,N_14053,N_14160);
and U14284 (N_14284,N_14016,N_14181);
nor U14285 (N_14285,N_14145,N_14143);
and U14286 (N_14286,N_14147,N_14047);
and U14287 (N_14287,N_14188,N_14176);
nor U14288 (N_14288,N_14023,N_14170);
and U14289 (N_14289,N_14167,N_14088);
nand U14290 (N_14290,N_14111,N_14184);
nor U14291 (N_14291,N_14024,N_14129);
and U14292 (N_14292,N_14100,N_14110);
and U14293 (N_14293,N_14055,N_14063);
and U14294 (N_14294,N_14004,N_14183);
nor U14295 (N_14295,N_14106,N_14050);
and U14296 (N_14296,N_14135,N_14051);
or U14297 (N_14297,N_14098,N_14078);
xor U14298 (N_14298,N_14155,N_14124);
nand U14299 (N_14299,N_14128,N_14046);
nand U14300 (N_14300,N_14165,N_14105);
or U14301 (N_14301,N_14053,N_14036);
or U14302 (N_14302,N_14013,N_14157);
and U14303 (N_14303,N_14057,N_14100);
nor U14304 (N_14304,N_14057,N_14185);
and U14305 (N_14305,N_14079,N_14001);
or U14306 (N_14306,N_14151,N_14055);
or U14307 (N_14307,N_14117,N_14078);
xnor U14308 (N_14308,N_14019,N_14092);
nand U14309 (N_14309,N_14053,N_14060);
xor U14310 (N_14310,N_14131,N_14189);
nor U14311 (N_14311,N_14043,N_14158);
or U14312 (N_14312,N_14021,N_14074);
and U14313 (N_14313,N_14138,N_14101);
nor U14314 (N_14314,N_14041,N_14007);
and U14315 (N_14315,N_14027,N_14170);
xor U14316 (N_14316,N_14154,N_14105);
or U14317 (N_14317,N_14003,N_14008);
xnor U14318 (N_14318,N_14191,N_14132);
nor U14319 (N_14319,N_14020,N_14151);
or U14320 (N_14320,N_14079,N_14103);
xnor U14321 (N_14321,N_14177,N_14025);
and U14322 (N_14322,N_14073,N_14133);
and U14323 (N_14323,N_14117,N_14021);
or U14324 (N_14324,N_14039,N_14008);
nand U14325 (N_14325,N_14147,N_14005);
nand U14326 (N_14326,N_14129,N_14112);
and U14327 (N_14327,N_14017,N_14016);
or U14328 (N_14328,N_14171,N_14088);
and U14329 (N_14329,N_14076,N_14081);
nand U14330 (N_14330,N_14121,N_14171);
or U14331 (N_14331,N_14080,N_14175);
nor U14332 (N_14332,N_14116,N_14155);
or U14333 (N_14333,N_14091,N_14197);
xor U14334 (N_14334,N_14029,N_14199);
xor U14335 (N_14335,N_14152,N_14125);
nor U14336 (N_14336,N_14096,N_14199);
or U14337 (N_14337,N_14025,N_14178);
and U14338 (N_14338,N_14050,N_14195);
and U14339 (N_14339,N_14067,N_14073);
xor U14340 (N_14340,N_14070,N_14105);
and U14341 (N_14341,N_14056,N_14110);
xor U14342 (N_14342,N_14054,N_14097);
and U14343 (N_14343,N_14192,N_14177);
xnor U14344 (N_14344,N_14141,N_14072);
nor U14345 (N_14345,N_14098,N_14186);
nor U14346 (N_14346,N_14064,N_14148);
xnor U14347 (N_14347,N_14004,N_14106);
nor U14348 (N_14348,N_14105,N_14115);
xor U14349 (N_14349,N_14185,N_14082);
and U14350 (N_14350,N_14112,N_14087);
nand U14351 (N_14351,N_14179,N_14134);
nand U14352 (N_14352,N_14024,N_14102);
and U14353 (N_14353,N_14013,N_14180);
and U14354 (N_14354,N_14107,N_14167);
nand U14355 (N_14355,N_14084,N_14146);
xor U14356 (N_14356,N_14160,N_14068);
or U14357 (N_14357,N_14089,N_14063);
nor U14358 (N_14358,N_14060,N_14030);
and U14359 (N_14359,N_14143,N_14090);
nand U14360 (N_14360,N_14166,N_14131);
xnor U14361 (N_14361,N_14063,N_14163);
nor U14362 (N_14362,N_14166,N_14180);
and U14363 (N_14363,N_14066,N_14061);
or U14364 (N_14364,N_14157,N_14115);
nand U14365 (N_14365,N_14174,N_14110);
nand U14366 (N_14366,N_14163,N_14108);
nand U14367 (N_14367,N_14015,N_14075);
nand U14368 (N_14368,N_14026,N_14033);
or U14369 (N_14369,N_14186,N_14108);
nand U14370 (N_14370,N_14112,N_14125);
nor U14371 (N_14371,N_14050,N_14031);
nor U14372 (N_14372,N_14165,N_14029);
xor U14373 (N_14373,N_14116,N_14137);
or U14374 (N_14374,N_14055,N_14076);
nand U14375 (N_14375,N_14069,N_14108);
nor U14376 (N_14376,N_14114,N_14044);
xnor U14377 (N_14377,N_14140,N_14010);
and U14378 (N_14378,N_14197,N_14111);
or U14379 (N_14379,N_14049,N_14062);
nand U14380 (N_14380,N_14190,N_14054);
and U14381 (N_14381,N_14182,N_14024);
nand U14382 (N_14382,N_14002,N_14035);
nor U14383 (N_14383,N_14137,N_14046);
xnor U14384 (N_14384,N_14098,N_14007);
nor U14385 (N_14385,N_14193,N_14132);
nand U14386 (N_14386,N_14096,N_14150);
and U14387 (N_14387,N_14188,N_14053);
nor U14388 (N_14388,N_14185,N_14099);
xnor U14389 (N_14389,N_14102,N_14140);
nor U14390 (N_14390,N_14086,N_14116);
xnor U14391 (N_14391,N_14077,N_14045);
nor U14392 (N_14392,N_14099,N_14133);
nand U14393 (N_14393,N_14105,N_14044);
nand U14394 (N_14394,N_14138,N_14016);
nor U14395 (N_14395,N_14114,N_14186);
xnor U14396 (N_14396,N_14017,N_14133);
or U14397 (N_14397,N_14138,N_14034);
nor U14398 (N_14398,N_14075,N_14156);
nor U14399 (N_14399,N_14038,N_14089);
nand U14400 (N_14400,N_14208,N_14293);
nor U14401 (N_14401,N_14322,N_14229);
nor U14402 (N_14402,N_14292,N_14327);
or U14403 (N_14403,N_14269,N_14386);
or U14404 (N_14404,N_14226,N_14276);
nor U14405 (N_14405,N_14300,N_14200);
and U14406 (N_14406,N_14360,N_14353);
and U14407 (N_14407,N_14241,N_14301);
and U14408 (N_14408,N_14221,N_14315);
or U14409 (N_14409,N_14263,N_14347);
or U14410 (N_14410,N_14278,N_14264);
or U14411 (N_14411,N_14374,N_14329);
xor U14412 (N_14412,N_14385,N_14381);
nand U14413 (N_14413,N_14289,N_14238);
or U14414 (N_14414,N_14320,N_14261);
and U14415 (N_14415,N_14215,N_14230);
nand U14416 (N_14416,N_14216,N_14399);
nand U14417 (N_14417,N_14205,N_14325);
and U14418 (N_14418,N_14224,N_14368);
xor U14419 (N_14419,N_14288,N_14249);
nor U14420 (N_14420,N_14319,N_14335);
xnor U14421 (N_14421,N_14384,N_14375);
nor U14422 (N_14422,N_14212,N_14234);
and U14423 (N_14423,N_14377,N_14390);
nand U14424 (N_14424,N_14214,N_14354);
xnor U14425 (N_14425,N_14338,N_14206);
nor U14426 (N_14426,N_14350,N_14201);
nand U14427 (N_14427,N_14253,N_14240);
xnor U14428 (N_14428,N_14337,N_14294);
nand U14429 (N_14429,N_14233,N_14244);
nand U14430 (N_14430,N_14317,N_14366);
or U14431 (N_14431,N_14286,N_14334);
nand U14432 (N_14432,N_14314,N_14239);
or U14433 (N_14433,N_14252,N_14380);
xor U14434 (N_14434,N_14248,N_14348);
xor U14435 (N_14435,N_14372,N_14296);
or U14436 (N_14436,N_14344,N_14243);
and U14437 (N_14437,N_14291,N_14257);
nand U14438 (N_14438,N_14357,N_14247);
nand U14439 (N_14439,N_14265,N_14379);
and U14440 (N_14440,N_14340,N_14280);
and U14441 (N_14441,N_14295,N_14262);
nor U14442 (N_14442,N_14367,N_14306);
and U14443 (N_14443,N_14259,N_14299);
or U14444 (N_14444,N_14395,N_14342);
and U14445 (N_14445,N_14333,N_14378);
nand U14446 (N_14446,N_14250,N_14392);
nand U14447 (N_14447,N_14323,N_14330);
nand U14448 (N_14448,N_14313,N_14321);
nor U14449 (N_14449,N_14236,N_14270);
nand U14450 (N_14450,N_14345,N_14284);
nor U14451 (N_14451,N_14363,N_14213);
and U14452 (N_14452,N_14343,N_14272);
nor U14453 (N_14453,N_14237,N_14290);
or U14454 (N_14454,N_14332,N_14246);
or U14455 (N_14455,N_14268,N_14397);
nor U14456 (N_14456,N_14203,N_14308);
or U14457 (N_14457,N_14307,N_14324);
and U14458 (N_14458,N_14369,N_14376);
nand U14459 (N_14459,N_14339,N_14225);
or U14460 (N_14460,N_14383,N_14254);
nor U14461 (N_14461,N_14305,N_14382);
nor U14462 (N_14462,N_14266,N_14207);
xor U14463 (N_14463,N_14298,N_14287);
or U14464 (N_14464,N_14228,N_14318);
nand U14465 (N_14465,N_14311,N_14396);
and U14466 (N_14466,N_14365,N_14393);
nand U14467 (N_14467,N_14231,N_14312);
nand U14468 (N_14468,N_14222,N_14336);
nand U14469 (N_14469,N_14391,N_14245);
or U14470 (N_14470,N_14362,N_14364);
and U14471 (N_14471,N_14359,N_14217);
and U14472 (N_14472,N_14210,N_14341);
nand U14473 (N_14473,N_14346,N_14389);
xnor U14474 (N_14474,N_14356,N_14388);
or U14475 (N_14475,N_14303,N_14309);
or U14476 (N_14476,N_14218,N_14227);
nand U14477 (N_14477,N_14398,N_14371);
nor U14478 (N_14478,N_14275,N_14328);
nand U14479 (N_14479,N_14267,N_14279);
xnor U14480 (N_14480,N_14302,N_14209);
nand U14481 (N_14481,N_14283,N_14204);
and U14482 (N_14482,N_14361,N_14271);
nor U14483 (N_14483,N_14310,N_14387);
nor U14484 (N_14484,N_14258,N_14297);
nand U14485 (N_14485,N_14220,N_14281);
xor U14486 (N_14486,N_14331,N_14304);
and U14487 (N_14487,N_14223,N_14316);
nor U14488 (N_14488,N_14326,N_14232);
and U14489 (N_14489,N_14282,N_14260);
nand U14490 (N_14490,N_14242,N_14351);
and U14491 (N_14491,N_14352,N_14394);
nor U14492 (N_14492,N_14251,N_14256);
nand U14493 (N_14493,N_14277,N_14255);
nand U14494 (N_14494,N_14235,N_14285);
nor U14495 (N_14495,N_14274,N_14370);
xnor U14496 (N_14496,N_14211,N_14219);
nor U14497 (N_14497,N_14358,N_14355);
xor U14498 (N_14498,N_14273,N_14202);
nand U14499 (N_14499,N_14349,N_14373);
xor U14500 (N_14500,N_14299,N_14240);
nor U14501 (N_14501,N_14398,N_14349);
and U14502 (N_14502,N_14323,N_14313);
nor U14503 (N_14503,N_14376,N_14302);
and U14504 (N_14504,N_14349,N_14338);
and U14505 (N_14505,N_14205,N_14203);
nor U14506 (N_14506,N_14398,N_14389);
xnor U14507 (N_14507,N_14399,N_14281);
xnor U14508 (N_14508,N_14364,N_14353);
xor U14509 (N_14509,N_14326,N_14348);
and U14510 (N_14510,N_14318,N_14382);
and U14511 (N_14511,N_14331,N_14352);
xor U14512 (N_14512,N_14213,N_14390);
nor U14513 (N_14513,N_14218,N_14205);
nor U14514 (N_14514,N_14364,N_14320);
nor U14515 (N_14515,N_14366,N_14320);
or U14516 (N_14516,N_14327,N_14283);
nand U14517 (N_14517,N_14299,N_14274);
xor U14518 (N_14518,N_14379,N_14395);
xnor U14519 (N_14519,N_14356,N_14208);
or U14520 (N_14520,N_14337,N_14244);
nor U14521 (N_14521,N_14340,N_14226);
and U14522 (N_14522,N_14334,N_14310);
and U14523 (N_14523,N_14399,N_14327);
nor U14524 (N_14524,N_14229,N_14240);
or U14525 (N_14525,N_14258,N_14334);
nand U14526 (N_14526,N_14393,N_14245);
and U14527 (N_14527,N_14224,N_14383);
nor U14528 (N_14528,N_14236,N_14393);
and U14529 (N_14529,N_14390,N_14362);
and U14530 (N_14530,N_14388,N_14321);
nor U14531 (N_14531,N_14267,N_14351);
and U14532 (N_14532,N_14385,N_14215);
xor U14533 (N_14533,N_14208,N_14398);
nand U14534 (N_14534,N_14336,N_14207);
or U14535 (N_14535,N_14275,N_14320);
and U14536 (N_14536,N_14364,N_14207);
nor U14537 (N_14537,N_14265,N_14373);
nor U14538 (N_14538,N_14318,N_14395);
nand U14539 (N_14539,N_14301,N_14233);
or U14540 (N_14540,N_14337,N_14306);
or U14541 (N_14541,N_14215,N_14278);
nor U14542 (N_14542,N_14206,N_14382);
and U14543 (N_14543,N_14208,N_14322);
xor U14544 (N_14544,N_14240,N_14391);
xnor U14545 (N_14545,N_14313,N_14283);
and U14546 (N_14546,N_14272,N_14322);
xor U14547 (N_14547,N_14222,N_14340);
nor U14548 (N_14548,N_14237,N_14205);
or U14549 (N_14549,N_14244,N_14351);
nand U14550 (N_14550,N_14255,N_14393);
nor U14551 (N_14551,N_14311,N_14264);
nor U14552 (N_14552,N_14386,N_14224);
and U14553 (N_14553,N_14294,N_14399);
nor U14554 (N_14554,N_14214,N_14230);
nor U14555 (N_14555,N_14315,N_14312);
nor U14556 (N_14556,N_14361,N_14380);
nor U14557 (N_14557,N_14247,N_14236);
xor U14558 (N_14558,N_14379,N_14368);
and U14559 (N_14559,N_14314,N_14218);
nand U14560 (N_14560,N_14254,N_14282);
and U14561 (N_14561,N_14315,N_14259);
or U14562 (N_14562,N_14367,N_14209);
nand U14563 (N_14563,N_14349,N_14391);
or U14564 (N_14564,N_14309,N_14335);
nor U14565 (N_14565,N_14226,N_14210);
or U14566 (N_14566,N_14200,N_14237);
and U14567 (N_14567,N_14266,N_14390);
nand U14568 (N_14568,N_14323,N_14374);
xor U14569 (N_14569,N_14340,N_14231);
nand U14570 (N_14570,N_14264,N_14294);
nand U14571 (N_14571,N_14288,N_14325);
or U14572 (N_14572,N_14269,N_14327);
nand U14573 (N_14573,N_14209,N_14214);
or U14574 (N_14574,N_14348,N_14399);
xnor U14575 (N_14575,N_14211,N_14336);
or U14576 (N_14576,N_14272,N_14300);
nor U14577 (N_14577,N_14237,N_14338);
or U14578 (N_14578,N_14298,N_14299);
xnor U14579 (N_14579,N_14382,N_14299);
xor U14580 (N_14580,N_14369,N_14334);
or U14581 (N_14581,N_14287,N_14388);
and U14582 (N_14582,N_14217,N_14282);
nand U14583 (N_14583,N_14225,N_14293);
xor U14584 (N_14584,N_14319,N_14380);
xnor U14585 (N_14585,N_14367,N_14284);
nand U14586 (N_14586,N_14235,N_14280);
xnor U14587 (N_14587,N_14326,N_14269);
nor U14588 (N_14588,N_14282,N_14280);
nand U14589 (N_14589,N_14284,N_14264);
nand U14590 (N_14590,N_14390,N_14257);
xor U14591 (N_14591,N_14228,N_14206);
and U14592 (N_14592,N_14251,N_14264);
and U14593 (N_14593,N_14344,N_14277);
or U14594 (N_14594,N_14268,N_14291);
or U14595 (N_14595,N_14397,N_14280);
or U14596 (N_14596,N_14266,N_14308);
and U14597 (N_14597,N_14377,N_14373);
nand U14598 (N_14598,N_14361,N_14258);
or U14599 (N_14599,N_14399,N_14347);
nor U14600 (N_14600,N_14419,N_14514);
nand U14601 (N_14601,N_14483,N_14448);
or U14602 (N_14602,N_14443,N_14585);
xor U14603 (N_14603,N_14450,N_14428);
nand U14604 (N_14604,N_14439,N_14577);
xor U14605 (N_14605,N_14520,N_14491);
nand U14606 (N_14606,N_14526,N_14493);
nor U14607 (N_14607,N_14413,N_14554);
nor U14608 (N_14608,N_14567,N_14513);
or U14609 (N_14609,N_14405,N_14432);
nor U14610 (N_14610,N_14541,N_14598);
nand U14611 (N_14611,N_14403,N_14519);
nand U14612 (N_14612,N_14478,N_14505);
xnor U14613 (N_14613,N_14453,N_14445);
and U14614 (N_14614,N_14442,N_14480);
and U14615 (N_14615,N_14431,N_14500);
nor U14616 (N_14616,N_14412,N_14589);
or U14617 (N_14617,N_14596,N_14415);
xnor U14618 (N_14618,N_14578,N_14551);
nor U14619 (N_14619,N_14416,N_14459);
nor U14620 (N_14620,N_14456,N_14475);
nor U14621 (N_14621,N_14438,N_14401);
xnor U14622 (N_14622,N_14467,N_14407);
xor U14623 (N_14623,N_14454,N_14540);
or U14624 (N_14624,N_14477,N_14455);
or U14625 (N_14625,N_14574,N_14510);
nand U14626 (N_14626,N_14521,N_14498);
or U14627 (N_14627,N_14511,N_14528);
or U14628 (N_14628,N_14408,N_14565);
and U14629 (N_14629,N_14468,N_14588);
nor U14630 (N_14630,N_14563,N_14400);
nor U14631 (N_14631,N_14460,N_14522);
and U14632 (N_14632,N_14470,N_14487);
xnor U14633 (N_14633,N_14469,N_14446);
xor U14634 (N_14634,N_14580,N_14536);
nor U14635 (N_14635,N_14489,N_14492);
or U14636 (N_14636,N_14523,N_14471);
or U14637 (N_14637,N_14462,N_14584);
nand U14638 (N_14638,N_14527,N_14576);
or U14639 (N_14639,N_14444,N_14441);
nand U14640 (N_14640,N_14575,N_14484);
nand U14641 (N_14641,N_14423,N_14414);
nand U14642 (N_14642,N_14564,N_14476);
nor U14643 (N_14643,N_14549,N_14566);
and U14644 (N_14644,N_14424,N_14546);
nor U14645 (N_14645,N_14482,N_14552);
nand U14646 (N_14646,N_14425,N_14494);
or U14647 (N_14647,N_14518,N_14508);
nand U14648 (N_14648,N_14561,N_14461);
or U14649 (N_14649,N_14464,N_14599);
and U14650 (N_14650,N_14555,N_14499);
and U14651 (N_14651,N_14557,N_14593);
xnor U14652 (N_14652,N_14586,N_14537);
and U14653 (N_14653,N_14422,N_14558);
xnor U14654 (N_14654,N_14581,N_14507);
and U14655 (N_14655,N_14426,N_14474);
nor U14656 (N_14656,N_14421,N_14569);
or U14657 (N_14657,N_14559,N_14449);
or U14658 (N_14658,N_14486,N_14597);
or U14659 (N_14659,N_14573,N_14587);
or U14660 (N_14660,N_14595,N_14544);
xor U14661 (N_14661,N_14506,N_14437);
and U14662 (N_14662,N_14447,N_14504);
nand U14663 (N_14663,N_14495,N_14545);
and U14664 (N_14664,N_14420,N_14556);
or U14665 (N_14665,N_14531,N_14579);
nor U14666 (N_14666,N_14570,N_14524);
xor U14667 (N_14667,N_14479,N_14560);
xnor U14668 (N_14668,N_14472,N_14533);
xnor U14669 (N_14669,N_14451,N_14502);
nor U14670 (N_14670,N_14402,N_14535);
or U14671 (N_14671,N_14434,N_14547);
or U14672 (N_14672,N_14488,N_14463);
or U14673 (N_14673,N_14503,N_14538);
nor U14674 (N_14674,N_14530,N_14457);
and U14675 (N_14675,N_14568,N_14571);
or U14676 (N_14676,N_14430,N_14406);
and U14677 (N_14677,N_14516,N_14572);
and U14678 (N_14678,N_14473,N_14512);
or U14679 (N_14679,N_14417,N_14592);
xor U14680 (N_14680,N_14436,N_14404);
nand U14681 (N_14681,N_14590,N_14515);
or U14682 (N_14682,N_14583,N_14427);
nor U14683 (N_14683,N_14532,N_14525);
and U14684 (N_14684,N_14517,N_14465);
nand U14685 (N_14685,N_14429,N_14529);
and U14686 (N_14686,N_14553,N_14485);
xnor U14687 (N_14687,N_14418,N_14550);
or U14688 (N_14688,N_14433,N_14466);
nor U14689 (N_14689,N_14452,N_14534);
xnor U14690 (N_14690,N_14542,N_14497);
or U14691 (N_14691,N_14411,N_14548);
or U14692 (N_14692,N_14458,N_14582);
or U14693 (N_14693,N_14562,N_14591);
nand U14694 (N_14694,N_14509,N_14410);
nor U14695 (N_14695,N_14496,N_14435);
or U14696 (N_14696,N_14594,N_14409);
or U14697 (N_14697,N_14490,N_14543);
and U14698 (N_14698,N_14440,N_14539);
nand U14699 (N_14699,N_14481,N_14501);
xnor U14700 (N_14700,N_14514,N_14537);
and U14701 (N_14701,N_14595,N_14594);
xor U14702 (N_14702,N_14431,N_14482);
and U14703 (N_14703,N_14598,N_14590);
xnor U14704 (N_14704,N_14540,N_14537);
and U14705 (N_14705,N_14495,N_14500);
or U14706 (N_14706,N_14488,N_14595);
or U14707 (N_14707,N_14497,N_14584);
nor U14708 (N_14708,N_14535,N_14455);
xnor U14709 (N_14709,N_14482,N_14422);
and U14710 (N_14710,N_14454,N_14551);
nand U14711 (N_14711,N_14456,N_14517);
nand U14712 (N_14712,N_14579,N_14506);
nor U14713 (N_14713,N_14444,N_14528);
and U14714 (N_14714,N_14423,N_14597);
or U14715 (N_14715,N_14537,N_14579);
nand U14716 (N_14716,N_14401,N_14497);
nor U14717 (N_14717,N_14585,N_14491);
nor U14718 (N_14718,N_14480,N_14406);
nor U14719 (N_14719,N_14448,N_14488);
xor U14720 (N_14720,N_14479,N_14451);
or U14721 (N_14721,N_14476,N_14483);
nor U14722 (N_14722,N_14573,N_14566);
and U14723 (N_14723,N_14469,N_14475);
and U14724 (N_14724,N_14568,N_14504);
nor U14725 (N_14725,N_14546,N_14542);
and U14726 (N_14726,N_14458,N_14525);
or U14727 (N_14727,N_14573,N_14568);
nor U14728 (N_14728,N_14594,N_14425);
or U14729 (N_14729,N_14502,N_14514);
and U14730 (N_14730,N_14515,N_14551);
nor U14731 (N_14731,N_14499,N_14532);
or U14732 (N_14732,N_14463,N_14562);
or U14733 (N_14733,N_14536,N_14490);
xnor U14734 (N_14734,N_14515,N_14465);
xnor U14735 (N_14735,N_14480,N_14579);
or U14736 (N_14736,N_14484,N_14420);
or U14737 (N_14737,N_14465,N_14486);
nor U14738 (N_14738,N_14481,N_14445);
nor U14739 (N_14739,N_14500,N_14567);
xor U14740 (N_14740,N_14460,N_14452);
and U14741 (N_14741,N_14526,N_14558);
nand U14742 (N_14742,N_14557,N_14454);
and U14743 (N_14743,N_14587,N_14546);
xnor U14744 (N_14744,N_14462,N_14443);
nor U14745 (N_14745,N_14570,N_14503);
nor U14746 (N_14746,N_14483,N_14409);
or U14747 (N_14747,N_14587,N_14450);
nand U14748 (N_14748,N_14586,N_14580);
nand U14749 (N_14749,N_14565,N_14585);
nand U14750 (N_14750,N_14436,N_14449);
nor U14751 (N_14751,N_14423,N_14552);
or U14752 (N_14752,N_14419,N_14550);
nand U14753 (N_14753,N_14445,N_14561);
nor U14754 (N_14754,N_14419,N_14463);
and U14755 (N_14755,N_14471,N_14437);
and U14756 (N_14756,N_14517,N_14547);
xnor U14757 (N_14757,N_14405,N_14475);
xor U14758 (N_14758,N_14424,N_14588);
or U14759 (N_14759,N_14487,N_14417);
nor U14760 (N_14760,N_14434,N_14514);
or U14761 (N_14761,N_14429,N_14473);
or U14762 (N_14762,N_14419,N_14495);
xor U14763 (N_14763,N_14598,N_14535);
or U14764 (N_14764,N_14409,N_14412);
or U14765 (N_14765,N_14587,N_14404);
nor U14766 (N_14766,N_14493,N_14535);
nor U14767 (N_14767,N_14465,N_14585);
nand U14768 (N_14768,N_14526,N_14490);
xnor U14769 (N_14769,N_14584,N_14402);
xor U14770 (N_14770,N_14485,N_14459);
xor U14771 (N_14771,N_14538,N_14492);
nor U14772 (N_14772,N_14440,N_14555);
or U14773 (N_14773,N_14510,N_14436);
nand U14774 (N_14774,N_14408,N_14411);
and U14775 (N_14775,N_14447,N_14479);
or U14776 (N_14776,N_14588,N_14419);
nand U14777 (N_14777,N_14503,N_14545);
nor U14778 (N_14778,N_14570,N_14554);
and U14779 (N_14779,N_14545,N_14442);
nand U14780 (N_14780,N_14538,N_14585);
xnor U14781 (N_14781,N_14537,N_14428);
nor U14782 (N_14782,N_14574,N_14454);
nand U14783 (N_14783,N_14585,N_14486);
xor U14784 (N_14784,N_14416,N_14586);
and U14785 (N_14785,N_14559,N_14597);
nand U14786 (N_14786,N_14500,N_14483);
and U14787 (N_14787,N_14522,N_14489);
nand U14788 (N_14788,N_14517,N_14427);
and U14789 (N_14789,N_14454,N_14527);
and U14790 (N_14790,N_14537,N_14455);
nor U14791 (N_14791,N_14424,N_14405);
xnor U14792 (N_14792,N_14480,N_14466);
nor U14793 (N_14793,N_14504,N_14499);
xor U14794 (N_14794,N_14522,N_14470);
nor U14795 (N_14795,N_14578,N_14547);
or U14796 (N_14796,N_14476,N_14427);
nand U14797 (N_14797,N_14444,N_14578);
nor U14798 (N_14798,N_14567,N_14452);
xnor U14799 (N_14799,N_14475,N_14417);
nor U14800 (N_14800,N_14714,N_14649);
xnor U14801 (N_14801,N_14762,N_14735);
and U14802 (N_14802,N_14718,N_14668);
nor U14803 (N_14803,N_14766,N_14682);
xnor U14804 (N_14804,N_14721,N_14773);
xor U14805 (N_14805,N_14733,N_14713);
nand U14806 (N_14806,N_14729,N_14663);
nand U14807 (N_14807,N_14661,N_14738);
xor U14808 (N_14808,N_14676,N_14761);
and U14809 (N_14809,N_14754,N_14653);
or U14810 (N_14810,N_14765,N_14785);
or U14811 (N_14811,N_14700,N_14793);
and U14812 (N_14812,N_14730,N_14657);
or U14813 (N_14813,N_14671,N_14731);
or U14814 (N_14814,N_14605,N_14734);
xnor U14815 (N_14815,N_14618,N_14737);
and U14816 (N_14816,N_14712,N_14614);
xor U14817 (N_14817,N_14710,N_14757);
nor U14818 (N_14818,N_14615,N_14781);
nand U14819 (N_14819,N_14770,N_14672);
and U14820 (N_14820,N_14795,N_14637);
nand U14821 (N_14821,N_14675,N_14646);
xnor U14822 (N_14822,N_14604,N_14651);
nor U14823 (N_14823,N_14679,N_14621);
xor U14824 (N_14824,N_14704,N_14607);
or U14825 (N_14825,N_14736,N_14626);
xor U14826 (N_14826,N_14799,N_14789);
or U14827 (N_14827,N_14719,N_14644);
nor U14828 (N_14828,N_14708,N_14778);
and U14829 (N_14829,N_14658,N_14774);
and U14830 (N_14830,N_14791,N_14788);
nand U14831 (N_14831,N_14709,N_14655);
or U14832 (N_14832,N_14716,N_14643);
nand U14833 (N_14833,N_14724,N_14727);
xnor U14834 (N_14834,N_14715,N_14640);
nand U14835 (N_14835,N_14698,N_14687);
and U14836 (N_14836,N_14650,N_14688);
and U14837 (N_14837,N_14798,N_14767);
or U14838 (N_14838,N_14622,N_14697);
nand U14839 (N_14839,N_14691,N_14630);
nor U14840 (N_14840,N_14602,N_14629);
nor U14841 (N_14841,N_14683,N_14685);
nor U14842 (N_14842,N_14780,N_14612);
nor U14843 (N_14843,N_14690,N_14786);
nand U14844 (N_14844,N_14775,N_14636);
xor U14845 (N_14845,N_14673,N_14641);
or U14846 (N_14846,N_14705,N_14656);
nand U14847 (N_14847,N_14723,N_14634);
and U14848 (N_14848,N_14739,N_14701);
nor U14849 (N_14849,N_14628,N_14776);
nand U14850 (N_14850,N_14702,N_14662);
and U14851 (N_14851,N_14642,N_14681);
or U14852 (N_14852,N_14611,N_14794);
and U14853 (N_14853,N_14792,N_14744);
nand U14854 (N_14854,N_14728,N_14711);
nand U14855 (N_14855,N_14667,N_14763);
and U14856 (N_14856,N_14722,N_14783);
or U14857 (N_14857,N_14624,N_14747);
nor U14858 (N_14858,N_14769,N_14619);
nor U14859 (N_14859,N_14695,N_14703);
xor U14860 (N_14860,N_14601,N_14760);
nor U14861 (N_14861,N_14678,N_14694);
nand U14862 (N_14862,N_14750,N_14693);
nor U14863 (N_14863,N_14732,N_14666);
xnor U14864 (N_14864,N_14742,N_14755);
and U14865 (N_14865,N_14680,N_14647);
nor U14866 (N_14866,N_14743,N_14686);
xor U14867 (N_14867,N_14740,N_14768);
or U14868 (N_14868,N_14677,N_14771);
nor U14869 (N_14869,N_14660,N_14608);
nand U14870 (N_14870,N_14670,N_14790);
or U14871 (N_14871,N_14669,N_14772);
or U14872 (N_14872,N_14684,N_14610);
nor U14873 (N_14873,N_14631,N_14758);
xnor U14874 (N_14874,N_14692,N_14613);
or U14875 (N_14875,N_14689,N_14664);
nand U14876 (N_14876,N_14674,N_14759);
nor U14877 (N_14877,N_14777,N_14706);
and U14878 (N_14878,N_14764,N_14751);
and U14879 (N_14879,N_14741,N_14717);
nand U14880 (N_14880,N_14797,N_14659);
or U14881 (N_14881,N_14696,N_14633);
nor U14882 (N_14882,N_14652,N_14746);
or U14883 (N_14883,N_14707,N_14725);
or U14884 (N_14884,N_14616,N_14620);
and U14885 (N_14885,N_14645,N_14627);
or U14886 (N_14886,N_14782,N_14639);
or U14887 (N_14887,N_14603,N_14752);
or U14888 (N_14888,N_14632,N_14665);
or U14889 (N_14889,N_14796,N_14606);
or U14890 (N_14890,N_14756,N_14638);
nand U14891 (N_14891,N_14787,N_14648);
nor U14892 (N_14892,N_14623,N_14753);
nor U14893 (N_14893,N_14609,N_14720);
or U14894 (N_14894,N_14617,N_14749);
and U14895 (N_14895,N_14779,N_14699);
and U14896 (N_14896,N_14600,N_14748);
or U14897 (N_14897,N_14745,N_14784);
nor U14898 (N_14898,N_14625,N_14635);
nand U14899 (N_14899,N_14654,N_14726);
xnor U14900 (N_14900,N_14625,N_14670);
or U14901 (N_14901,N_14640,N_14772);
and U14902 (N_14902,N_14693,N_14734);
and U14903 (N_14903,N_14733,N_14652);
and U14904 (N_14904,N_14699,N_14666);
xor U14905 (N_14905,N_14790,N_14787);
xnor U14906 (N_14906,N_14771,N_14605);
nor U14907 (N_14907,N_14778,N_14756);
and U14908 (N_14908,N_14746,N_14695);
or U14909 (N_14909,N_14672,N_14755);
or U14910 (N_14910,N_14665,N_14753);
and U14911 (N_14911,N_14628,N_14662);
nand U14912 (N_14912,N_14662,N_14667);
xor U14913 (N_14913,N_14795,N_14777);
nand U14914 (N_14914,N_14771,N_14723);
nand U14915 (N_14915,N_14752,N_14694);
or U14916 (N_14916,N_14799,N_14635);
and U14917 (N_14917,N_14642,N_14711);
nor U14918 (N_14918,N_14753,N_14786);
xor U14919 (N_14919,N_14610,N_14782);
and U14920 (N_14920,N_14679,N_14782);
and U14921 (N_14921,N_14625,N_14639);
xnor U14922 (N_14922,N_14783,N_14702);
nand U14923 (N_14923,N_14700,N_14641);
and U14924 (N_14924,N_14783,N_14602);
and U14925 (N_14925,N_14786,N_14765);
or U14926 (N_14926,N_14764,N_14722);
nand U14927 (N_14927,N_14704,N_14752);
or U14928 (N_14928,N_14604,N_14623);
xor U14929 (N_14929,N_14696,N_14668);
and U14930 (N_14930,N_14679,N_14628);
nor U14931 (N_14931,N_14666,N_14690);
nor U14932 (N_14932,N_14665,N_14741);
xor U14933 (N_14933,N_14739,N_14691);
nor U14934 (N_14934,N_14799,N_14605);
xor U14935 (N_14935,N_14640,N_14674);
nand U14936 (N_14936,N_14736,N_14679);
nor U14937 (N_14937,N_14652,N_14685);
and U14938 (N_14938,N_14722,N_14701);
or U14939 (N_14939,N_14778,N_14695);
nor U14940 (N_14940,N_14730,N_14767);
nor U14941 (N_14941,N_14684,N_14699);
nor U14942 (N_14942,N_14697,N_14719);
and U14943 (N_14943,N_14621,N_14710);
nor U14944 (N_14944,N_14743,N_14690);
and U14945 (N_14945,N_14639,N_14720);
nor U14946 (N_14946,N_14601,N_14729);
nor U14947 (N_14947,N_14638,N_14731);
and U14948 (N_14948,N_14620,N_14729);
nand U14949 (N_14949,N_14748,N_14783);
nor U14950 (N_14950,N_14725,N_14794);
nor U14951 (N_14951,N_14660,N_14798);
nor U14952 (N_14952,N_14670,N_14607);
nand U14953 (N_14953,N_14601,N_14742);
or U14954 (N_14954,N_14614,N_14616);
and U14955 (N_14955,N_14734,N_14625);
and U14956 (N_14956,N_14605,N_14773);
or U14957 (N_14957,N_14620,N_14629);
nor U14958 (N_14958,N_14778,N_14656);
or U14959 (N_14959,N_14771,N_14624);
and U14960 (N_14960,N_14767,N_14631);
and U14961 (N_14961,N_14716,N_14672);
or U14962 (N_14962,N_14762,N_14618);
nand U14963 (N_14963,N_14639,N_14771);
and U14964 (N_14964,N_14640,N_14624);
xor U14965 (N_14965,N_14732,N_14662);
xor U14966 (N_14966,N_14794,N_14645);
or U14967 (N_14967,N_14622,N_14776);
xor U14968 (N_14968,N_14768,N_14673);
nor U14969 (N_14969,N_14706,N_14705);
and U14970 (N_14970,N_14738,N_14703);
or U14971 (N_14971,N_14684,N_14774);
xor U14972 (N_14972,N_14763,N_14768);
or U14973 (N_14973,N_14688,N_14631);
and U14974 (N_14974,N_14609,N_14789);
xor U14975 (N_14975,N_14619,N_14652);
and U14976 (N_14976,N_14734,N_14703);
nor U14977 (N_14977,N_14766,N_14608);
nand U14978 (N_14978,N_14645,N_14702);
and U14979 (N_14979,N_14674,N_14703);
nand U14980 (N_14980,N_14679,N_14727);
xnor U14981 (N_14981,N_14767,N_14722);
or U14982 (N_14982,N_14630,N_14775);
nand U14983 (N_14983,N_14704,N_14605);
and U14984 (N_14984,N_14758,N_14739);
and U14985 (N_14985,N_14605,N_14779);
and U14986 (N_14986,N_14760,N_14704);
nor U14987 (N_14987,N_14709,N_14622);
nand U14988 (N_14988,N_14686,N_14762);
and U14989 (N_14989,N_14688,N_14726);
or U14990 (N_14990,N_14664,N_14611);
nor U14991 (N_14991,N_14743,N_14758);
xor U14992 (N_14992,N_14712,N_14693);
and U14993 (N_14993,N_14613,N_14684);
xnor U14994 (N_14994,N_14737,N_14660);
nor U14995 (N_14995,N_14613,N_14602);
xor U14996 (N_14996,N_14603,N_14693);
nor U14997 (N_14997,N_14693,N_14641);
or U14998 (N_14998,N_14680,N_14602);
and U14999 (N_14999,N_14710,N_14620);
xor U15000 (N_15000,N_14963,N_14988);
and U15001 (N_15001,N_14850,N_14964);
nor U15002 (N_15002,N_14950,N_14918);
nand U15003 (N_15003,N_14965,N_14823);
nor U15004 (N_15004,N_14805,N_14994);
xnor U15005 (N_15005,N_14920,N_14906);
xor U15006 (N_15006,N_14949,N_14861);
nand U15007 (N_15007,N_14890,N_14970);
nand U15008 (N_15008,N_14904,N_14808);
xnor U15009 (N_15009,N_14814,N_14903);
and U15010 (N_15010,N_14824,N_14930);
nand U15011 (N_15011,N_14907,N_14831);
and U15012 (N_15012,N_14835,N_14853);
nand U15013 (N_15013,N_14945,N_14860);
nand U15014 (N_15014,N_14877,N_14826);
nor U15015 (N_15015,N_14924,N_14966);
xnor U15016 (N_15016,N_14923,N_14961);
xnor U15017 (N_15017,N_14957,N_14883);
xor U15018 (N_15018,N_14955,N_14810);
nor U15019 (N_15019,N_14940,N_14978);
nand U15020 (N_15020,N_14857,N_14977);
nand U15021 (N_15021,N_14820,N_14913);
or U15022 (N_15022,N_14954,N_14878);
nor U15023 (N_15023,N_14933,N_14973);
nor U15024 (N_15024,N_14919,N_14827);
xor U15025 (N_15025,N_14927,N_14894);
nor U15026 (N_15026,N_14901,N_14999);
nor U15027 (N_15027,N_14881,N_14889);
or U15028 (N_15028,N_14873,N_14862);
or U15029 (N_15029,N_14819,N_14884);
or U15030 (N_15030,N_14993,N_14944);
xnor U15031 (N_15031,N_14854,N_14971);
nor U15032 (N_15032,N_14836,N_14837);
xor U15033 (N_15033,N_14981,N_14912);
xor U15034 (N_15034,N_14991,N_14951);
or U15035 (N_15035,N_14905,N_14852);
nand U15036 (N_15036,N_14958,N_14975);
or U15037 (N_15037,N_14804,N_14932);
and U15038 (N_15038,N_14897,N_14813);
xor U15039 (N_15039,N_14845,N_14847);
or U15040 (N_15040,N_14856,N_14926);
nor U15041 (N_15041,N_14983,N_14886);
nor U15042 (N_15042,N_14997,N_14867);
and U15043 (N_15043,N_14969,N_14888);
nor U15044 (N_15044,N_14896,N_14815);
or U15045 (N_15045,N_14870,N_14938);
or U15046 (N_15046,N_14990,N_14960);
and U15047 (N_15047,N_14830,N_14911);
xor U15048 (N_15048,N_14967,N_14895);
nand U15049 (N_15049,N_14974,N_14979);
nand U15050 (N_15050,N_14803,N_14909);
or U15051 (N_15051,N_14807,N_14855);
or U15052 (N_15052,N_14832,N_14834);
nor U15053 (N_15053,N_14874,N_14929);
or U15054 (N_15054,N_14843,N_14908);
xnor U15055 (N_15055,N_14900,N_14863);
nand U15056 (N_15056,N_14892,N_14921);
nor U15057 (N_15057,N_14898,N_14809);
and U15058 (N_15058,N_14828,N_14917);
and U15059 (N_15059,N_14865,N_14996);
nor U15060 (N_15060,N_14992,N_14995);
or U15061 (N_15061,N_14839,N_14869);
nor U15062 (N_15062,N_14866,N_14915);
nand U15063 (N_15063,N_14887,N_14982);
xnor U15064 (N_15064,N_14942,N_14914);
nor U15065 (N_15065,N_14800,N_14976);
nor U15066 (N_15066,N_14816,N_14821);
xnor U15067 (N_15067,N_14956,N_14818);
nor U15068 (N_15068,N_14806,N_14851);
nor U15069 (N_15069,N_14941,N_14962);
nor U15070 (N_15070,N_14943,N_14980);
or U15071 (N_15071,N_14959,N_14880);
and U15072 (N_15072,N_14931,N_14953);
xnor U15073 (N_15073,N_14802,N_14848);
or U15074 (N_15074,N_14939,N_14833);
and U15075 (N_15075,N_14849,N_14858);
nand U15076 (N_15076,N_14893,N_14868);
xnor U15077 (N_15077,N_14902,N_14948);
and U15078 (N_15078,N_14998,N_14871);
or U15079 (N_15079,N_14891,N_14935);
nor U15080 (N_15080,N_14952,N_14859);
nand U15081 (N_15081,N_14986,N_14882);
nand U15082 (N_15082,N_14936,N_14846);
xor U15083 (N_15083,N_14876,N_14937);
nand U15084 (N_15084,N_14910,N_14879);
nand U15085 (N_15085,N_14825,N_14812);
nand U15086 (N_15086,N_14842,N_14985);
nor U15087 (N_15087,N_14801,N_14968);
and U15088 (N_15088,N_14872,N_14989);
or U15089 (N_15089,N_14811,N_14841);
nand U15090 (N_15090,N_14916,N_14925);
or U15091 (N_15091,N_14864,N_14822);
xor U15092 (N_15092,N_14885,N_14844);
or U15093 (N_15093,N_14934,N_14838);
nand U15094 (N_15094,N_14984,N_14987);
or U15095 (N_15095,N_14840,N_14922);
or U15096 (N_15096,N_14829,N_14817);
nand U15097 (N_15097,N_14972,N_14875);
nand U15098 (N_15098,N_14946,N_14947);
xor U15099 (N_15099,N_14899,N_14928);
and U15100 (N_15100,N_14882,N_14961);
nor U15101 (N_15101,N_14988,N_14940);
xnor U15102 (N_15102,N_14917,N_14874);
or U15103 (N_15103,N_14806,N_14817);
xnor U15104 (N_15104,N_14942,N_14835);
or U15105 (N_15105,N_14978,N_14847);
xnor U15106 (N_15106,N_14883,N_14953);
and U15107 (N_15107,N_14825,N_14803);
or U15108 (N_15108,N_14841,N_14859);
and U15109 (N_15109,N_14999,N_14857);
nor U15110 (N_15110,N_14966,N_14813);
and U15111 (N_15111,N_14992,N_14889);
nor U15112 (N_15112,N_14831,N_14974);
nand U15113 (N_15113,N_14900,N_14832);
and U15114 (N_15114,N_14853,N_14932);
and U15115 (N_15115,N_14836,N_14847);
nand U15116 (N_15116,N_14927,N_14966);
nor U15117 (N_15117,N_14898,N_14878);
and U15118 (N_15118,N_14910,N_14947);
nand U15119 (N_15119,N_14855,N_14969);
xnor U15120 (N_15120,N_14916,N_14883);
and U15121 (N_15121,N_14984,N_14941);
xor U15122 (N_15122,N_14891,N_14956);
and U15123 (N_15123,N_14840,N_14841);
nor U15124 (N_15124,N_14827,N_14901);
or U15125 (N_15125,N_14918,N_14955);
and U15126 (N_15126,N_14804,N_14975);
nand U15127 (N_15127,N_14892,N_14996);
and U15128 (N_15128,N_14913,N_14862);
nor U15129 (N_15129,N_14868,N_14856);
or U15130 (N_15130,N_14975,N_14935);
or U15131 (N_15131,N_14827,N_14957);
or U15132 (N_15132,N_14995,N_14865);
xnor U15133 (N_15133,N_14955,N_14822);
nor U15134 (N_15134,N_14826,N_14847);
or U15135 (N_15135,N_14810,N_14903);
nand U15136 (N_15136,N_14994,N_14888);
and U15137 (N_15137,N_14890,N_14834);
nor U15138 (N_15138,N_14943,N_14989);
nor U15139 (N_15139,N_14856,N_14855);
nand U15140 (N_15140,N_14943,N_14946);
or U15141 (N_15141,N_14967,N_14989);
or U15142 (N_15142,N_14906,N_14859);
nand U15143 (N_15143,N_14888,N_14899);
or U15144 (N_15144,N_14839,N_14966);
nand U15145 (N_15145,N_14867,N_14892);
nor U15146 (N_15146,N_14807,N_14856);
or U15147 (N_15147,N_14971,N_14828);
nor U15148 (N_15148,N_14976,N_14823);
or U15149 (N_15149,N_14928,N_14869);
nand U15150 (N_15150,N_14802,N_14871);
nand U15151 (N_15151,N_14912,N_14868);
or U15152 (N_15152,N_14936,N_14905);
xnor U15153 (N_15153,N_14937,N_14935);
nand U15154 (N_15154,N_14835,N_14995);
and U15155 (N_15155,N_14961,N_14916);
nand U15156 (N_15156,N_14993,N_14815);
nand U15157 (N_15157,N_14900,N_14968);
or U15158 (N_15158,N_14833,N_14979);
nand U15159 (N_15159,N_14837,N_14818);
and U15160 (N_15160,N_14976,N_14864);
nor U15161 (N_15161,N_14838,N_14957);
nand U15162 (N_15162,N_14990,N_14833);
or U15163 (N_15163,N_14977,N_14826);
and U15164 (N_15164,N_14868,N_14979);
or U15165 (N_15165,N_14878,N_14953);
or U15166 (N_15166,N_14995,N_14953);
nand U15167 (N_15167,N_14863,N_14812);
nand U15168 (N_15168,N_14910,N_14821);
and U15169 (N_15169,N_14983,N_14934);
or U15170 (N_15170,N_14993,N_14976);
nor U15171 (N_15171,N_14921,N_14977);
or U15172 (N_15172,N_14809,N_14993);
or U15173 (N_15173,N_14893,N_14940);
or U15174 (N_15174,N_14811,N_14865);
xnor U15175 (N_15175,N_14893,N_14801);
or U15176 (N_15176,N_14926,N_14885);
nand U15177 (N_15177,N_14891,N_14984);
xnor U15178 (N_15178,N_14901,N_14883);
or U15179 (N_15179,N_14917,N_14869);
or U15180 (N_15180,N_14829,N_14803);
xnor U15181 (N_15181,N_14862,N_14941);
nand U15182 (N_15182,N_14963,N_14880);
xor U15183 (N_15183,N_14973,N_14903);
nand U15184 (N_15184,N_14835,N_14890);
nor U15185 (N_15185,N_14938,N_14955);
xnor U15186 (N_15186,N_14916,N_14865);
nor U15187 (N_15187,N_14846,N_14818);
or U15188 (N_15188,N_14871,N_14880);
and U15189 (N_15189,N_14850,N_14884);
nor U15190 (N_15190,N_14887,N_14976);
and U15191 (N_15191,N_14933,N_14941);
and U15192 (N_15192,N_14808,N_14964);
and U15193 (N_15193,N_14968,N_14829);
nand U15194 (N_15194,N_14960,N_14858);
xnor U15195 (N_15195,N_14840,N_14821);
nor U15196 (N_15196,N_14975,N_14988);
nand U15197 (N_15197,N_14869,N_14811);
nand U15198 (N_15198,N_14827,N_14967);
and U15199 (N_15199,N_14876,N_14806);
nand U15200 (N_15200,N_15098,N_15025);
nor U15201 (N_15201,N_15177,N_15002);
nand U15202 (N_15202,N_15023,N_15007);
nand U15203 (N_15203,N_15166,N_15170);
or U15204 (N_15204,N_15157,N_15184);
xor U15205 (N_15205,N_15021,N_15001);
nor U15206 (N_15206,N_15044,N_15128);
nand U15207 (N_15207,N_15140,N_15014);
nor U15208 (N_15208,N_15058,N_15005);
nand U15209 (N_15209,N_15103,N_15163);
nor U15210 (N_15210,N_15075,N_15082);
nand U15211 (N_15211,N_15095,N_15053);
xnor U15212 (N_15212,N_15091,N_15046);
or U15213 (N_15213,N_15059,N_15174);
or U15214 (N_15214,N_15189,N_15169);
and U15215 (N_15215,N_15136,N_15097);
xnor U15216 (N_15216,N_15137,N_15070);
and U15217 (N_15217,N_15067,N_15181);
xor U15218 (N_15218,N_15020,N_15084);
nor U15219 (N_15219,N_15042,N_15194);
nand U15220 (N_15220,N_15175,N_15145);
nor U15221 (N_15221,N_15028,N_15065);
xnor U15222 (N_15222,N_15093,N_15073);
nand U15223 (N_15223,N_15167,N_15118);
or U15224 (N_15224,N_15120,N_15016);
nor U15225 (N_15225,N_15133,N_15012);
xor U15226 (N_15226,N_15198,N_15032);
nand U15227 (N_15227,N_15050,N_15147);
nand U15228 (N_15228,N_15154,N_15105);
or U15229 (N_15229,N_15109,N_15164);
or U15230 (N_15230,N_15022,N_15078);
nand U15231 (N_15231,N_15188,N_15008);
or U15232 (N_15232,N_15106,N_15009);
nand U15233 (N_15233,N_15116,N_15179);
or U15234 (N_15234,N_15015,N_15013);
nor U15235 (N_15235,N_15038,N_15102);
xor U15236 (N_15236,N_15076,N_15165);
nand U15237 (N_15237,N_15158,N_15191);
or U15238 (N_15238,N_15132,N_15026);
or U15239 (N_15239,N_15135,N_15148);
or U15240 (N_15240,N_15161,N_15143);
nor U15241 (N_15241,N_15192,N_15096);
nand U15242 (N_15242,N_15049,N_15153);
or U15243 (N_15243,N_15069,N_15024);
nor U15244 (N_15244,N_15045,N_15077);
xnor U15245 (N_15245,N_15017,N_15115);
or U15246 (N_15246,N_15149,N_15139);
xor U15247 (N_15247,N_15003,N_15151);
nor U15248 (N_15248,N_15036,N_15122);
or U15249 (N_15249,N_15010,N_15054);
nand U15250 (N_15250,N_15186,N_15071);
or U15251 (N_15251,N_15112,N_15123);
xor U15252 (N_15252,N_15138,N_15094);
or U15253 (N_15253,N_15029,N_15035);
xor U15254 (N_15254,N_15144,N_15155);
or U15255 (N_15255,N_15006,N_15197);
nor U15256 (N_15256,N_15004,N_15039);
nand U15257 (N_15257,N_15159,N_15027);
xor U15258 (N_15258,N_15108,N_15030);
nand U15259 (N_15259,N_15099,N_15168);
nor U15260 (N_15260,N_15126,N_15083);
nor U15261 (N_15261,N_15111,N_15055);
nand U15262 (N_15262,N_15092,N_15033);
xnor U15263 (N_15263,N_15068,N_15113);
or U15264 (N_15264,N_15130,N_15187);
nor U15265 (N_15265,N_15152,N_15171);
xnor U15266 (N_15266,N_15195,N_15019);
nand U15267 (N_15267,N_15119,N_15041);
or U15268 (N_15268,N_15162,N_15101);
nand U15269 (N_15269,N_15088,N_15063);
nor U15270 (N_15270,N_15156,N_15086);
nand U15271 (N_15271,N_15125,N_15121);
or U15272 (N_15272,N_15127,N_15142);
nor U15273 (N_15273,N_15089,N_15114);
nand U15274 (N_15274,N_15062,N_15000);
nor U15275 (N_15275,N_15104,N_15011);
or U15276 (N_15276,N_15185,N_15129);
and U15277 (N_15277,N_15090,N_15066);
and U15278 (N_15278,N_15196,N_15056);
or U15279 (N_15279,N_15080,N_15048);
nor U15280 (N_15280,N_15110,N_15172);
or U15281 (N_15281,N_15131,N_15031);
nand U15282 (N_15282,N_15085,N_15183);
xor U15283 (N_15283,N_15146,N_15087);
nor U15284 (N_15284,N_15117,N_15072);
or U15285 (N_15285,N_15141,N_15100);
nor U15286 (N_15286,N_15193,N_15018);
or U15287 (N_15287,N_15124,N_15081);
nand U15288 (N_15288,N_15180,N_15064);
or U15289 (N_15289,N_15057,N_15107);
nor U15290 (N_15290,N_15182,N_15061);
nand U15291 (N_15291,N_15052,N_15199);
xnor U15292 (N_15292,N_15040,N_15037);
xnor U15293 (N_15293,N_15060,N_15173);
nand U15294 (N_15294,N_15190,N_15178);
xor U15295 (N_15295,N_15079,N_15051);
nand U15296 (N_15296,N_15150,N_15043);
xnor U15297 (N_15297,N_15074,N_15034);
or U15298 (N_15298,N_15047,N_15134);
xor U15299 (N_15299,N_15176,N_15160);
nand U15300 (N_15300,N_15115,N_15122);
nor U15301 (N_15301,N_15046,N_15010);
nor U15302 (N_15302,N_15115,N_15162);
and U15303 (N_15303,N_15121,N_15147);
xor U15304 (N_15304,N_15041,N_15051);
and U15305 (N_15305,N_15071,N_15058);
xor U15306 (N_15306,N_15098,N_15138);
nor U15307 (N_15307,N_15114,N_15190);
xor U15308 (N_15308,N_15158,N_15111);
and U15309 (N_15309,N_15134,N_15044);
and U15310 (N_15310,N_15034,N_15188);
nand U15311 (N_15311,N_15181,N_15080);
nor U15312 (N_15312,N_15125,N_15147);
and U15313 (N_15313,N_15118,N_15094);
xnor U15314 (N_15314,N_15068,N_15084);
and U15315 (N_15315,N_15063,N_15020);
xor U15316 (N_15316,N_15101,N_15056);
xor U15317 (N_15317,N_15193,N_15078);
and U15318 (N_15318,N_15092,N_15108);
nor U15319 (N_15319,N_15048,N_15026);
and U15320 (N_15320,N_15139,N_15115);
nor U15321 (N_15321,N_15115,N_15051);
xor U15322 (N_15322,N_15156,N_15148);
nor U15323 (N_15323,N_15042,N_15157);
and U15324 (N_15324,N_15082,N_15152);
nand U15325 (N_15325,N_15069,N_15170);
or U15326 (N_15326,N_15156,N_15122);
nand U15327 (N_15327,N_15186,N_15041);
nand U15328 (N_15328,N_15013,N_15084);
nand U15329 (N_15329,N_15053,N_15052);
nor U15330 (N_15330,N_15163,N_15004);
nand U15331 (N_15331,N_15009,N_15102);
xor U15332 (N_15332,N_15178,N_15007);
nand U15333 (N_15333,N_15168,N_15003);
or U15334 (N_15334,N_15007,N_15171);
nand U15335 (N_15335,N_15003,N_15006);
nand U15336 (N_15336,N_15008,N_15141);
xnor U15337 (N_15337,N_15042,N_15113);
xnor U15338 (N_15338,N_15146,N_15041);
xnor U15339 (N_15339,N_15105,N_15043);
xor U15340 (N_15340,N_15005,N_15023);
nand U15341 (N_15341,N_15058,N_15129);
or U15342 (N_15342,N_15173,N_15130);
or U15343 (N_15343,N_15174,N_15060);
or U15344 (N_15344,N_15020,N_15164);
or U15345 (N_15345,N_15096,N_15099);
or U15346 (N_15346,N_15142,N_15135);
and U15347 (N_15347,N_15083,N_15081);
nor U15348 (N_15348,N_15108,N_15122);
xnor U15349 (N_15349,N_15117,N_15083);
xnor U15350 (N_15350,N_15075,N_15016);
and U15351 (N_15351,N_15056,N_15082);
or U15352 (N_15352,N_15064,N_15133);
nor U15353 (N_15353,N_15134,N_15079);
and U15354 (N_15354,N_15130,N_15149);
nand U15355 (N_15355,N_15074,N_15067);
nor U15356 (N_15356,N_15109,N_15182);
and U15357 (N_15357,N_15012,N_15079);
and U15358 (N_15358,N_15059,N_15040);
nor U15359 (N_15359,N_15098,N_15187);
nor U15360 (N_15360,N_15117,N_15081);
and U15361 (N_15361,N_15188,N_15050);
nand U15362 (N_15362,N_15037,N_15030);
nand U15363 (N_15363,N_15039,N_15060);
nand U15364 (N_15364,N_15068,N_15157);
nor U15365 (N_15365,N_15117,N_15180);
or U15366 (N_15366,N_15162,N_15058);
or U15367 (N_15367,N_15149,N_15010);
xor U15368 (N_15368,N_15131,N_15135);
nor U15369 (N_15369,N_15018,N_15020);
nor U15370 (N_15370,N_15188,N_15194);
or U15371 (N_15371,N_15033,N_15145);
or U15372 (N_15372,N_15095,N_15089);
and U15373 (N_15373,N_15165,N_15153);
or U15374 (N_15374,N_15086,N_15141);
nand U15375 (N_15375,N_15105,N_15183);
or U15376 (N_15376,N_15167,N_15011);
and U15377 (N_15377,N_15111,N_15145);
or U15378 (N_15378,N_15101,N_15194);
or U15379 (N_15379,N_15155,N_15167);
and U15380 (N_15380,N_15032,N_15143);
or U15381 (N_15381,N_15026,N_15027);
nand U15382 (N_15382,N_15173,N_15152);
or U15383 (N_15383,N_15064,N_15061);
nand U15384 (N_15384,N_15072,N_15042);
or U15385 (N_15385,N_15012,N_15162);
nand U15386 (N_15386,N_15143,N_15080);
nand U15387 (N_15387,N_15064,N_15161);
nor U15388 (N_15388,N_15041,N_15181);
or U15389 (N_15389,N_15138,N_15069);
nor U15390 (N_15390,N_15070,N_15034);
or U15391 (N_15391,N_15185,N_15078);
and U15392 (N_15392,N_15061,N_15033);
xnor U15393 (N_15393,N_15057,N_15197);
and U15394 (N_15394,N_15133,N_15177);
xor U15395 (N_15395,N_15181,N_15059);
or U15396 (N_15396,N_15092,N_15046);
and U15397 (N_15397,N_15109,N_15035);
nor U15398 (N_15398,N_15126,N_15176);
nor U15399 (N_15399,N_15027,N_15035);
xor U15400 (N_15400,N_15226,N_15205);
nand U15401 (N_15401,N_15313,N_15295);
or U15402 (N_15402,N_15257,N_15362);
or U15403 (N_15403,N_15261,N_15213);
nand U15404 (N_15404,N_15386,N_15218);
xnor U15405 (N_15405,N_15384,N_15368);
nand U15406 (N_15406,N_15350,N_15298);
nand U15407 (N_15407,N_15397,N_15279);
or U15408 (N_15408,N_15234,N_15381);
or U15409 (N_15409,N_15260,N_15270);
nand U15410 (N_15410,N_15389,N_15275);
xnor U15411 (N_15411,N_15282,N_15366);
or U15412 (N_15412,N_15277,N_15332);
and U15413 (N_15413,N_15237,N_15251);
or U15414 (N_15414,N_15307,N_15399);
nor U15415 (N_15415,N_15278,N_15239);
nor U15416 (N_15416,N_15266,N_15243);
xor U15417 (N_15417,N_15301,N_15342);
or U15418 (N_15418,N_15391,N_15352);
xnor U15419 (N_15419,N_15367,N_15273);
nor U15420 (N_15420,N_15259,N_15244);
nand U15421 (N_15421,N_15292,N_15358);
nor U15422 (N_15422,N_15258,N_15222);
xnor U15423 (N_15423,N_15291,N_15221);
xnor U15424 (N_15424,N_15371,N_15289);
nand U15425 (N_15425,N_15286,N_15379);
xnor U15426 (N_15426,N_15363,N_15232);
nor U15427 (N_15427,N_15223,N_15348);
nand U15428 (N_15428,N_15281,N_15250);
or U15429 (N_15429,N_15327,N_15320);
or U15430 (N_15430,N_15268,N_15328);
and U15431 (N_15431,N_15267,N_15207);
nand U15432 (N_15432,N_15249,N_15308);
nor U15433 (N_15433,N_15231,N_15297);
nand U15434 (N_15434,N_15290,N_15293);
nor U15435 (N_15435,N_15382,N_15321);
or U15436 (N_15436,N_15316,N_15233);
or U15437 (N_15437,N_15387,N_15309);
nand U15438 (N_15438,N_15303,N_15253);
nor U15439 (N_15439,N_15378,N_15353);
xor U15440 (N_15440,N_15317,N_15256);
and U15441 (N_15441,N_15325,N_15288);
or U15442 (N_15442,N_15326,N_15377);
nand U15443 (N_15443,N_15246,N_15370);
nand U15444 (N_15444,N_15361,N_15340);
and U15445 (N_15445,N_15294,N_15283);
nor U15446 (N_15446,N_15375,N_15214);
nor U15447 (N_15447,N_15343,N_15346);
or U15448 (N_15448,N_15240,N_15312);
nor U15449 (N_15449,N_15311,N_15322);
nor U15450 (N_15450,N_15235,N_15210);
and U15451 (N_15451,N_15225,N_15330);
or U15452 (N_15452,N_15242,N_15365);
and U15453 (N_15453,N_15344,N_15349);
nand U15454 (N_15454,N_15241,N_15238);
and U15455 (N_15455,N_15236,N_15300);
xnor U15456 (N_15456,N_15206,N_15254);
xor U15457 (N_15457,N_15395,N_15310);
and U15458 (N_15458,N_15360,N_15219);
or U15459 (N_15459,N_15398,N_15285);
nand U15460 (N_15460,N_15336,N_15247);
nand U15461 (N_15461,N_15319,N_15357);
and U15462 (N_15462,N_15262,N_15209);
xnor U15463 (N_15463,N_15369,N_15202);
and U15464 (N_15464,N_15211,N_15263);
and U15465 (N_15465,N_15302,N_15335);
nor U15466 (N_15466,N_15208,N_15315);
or U15467 (N_15467,N_15341,N_15380);
nand U15468 (N_15468,N_15334,N_15396);
nand U15469 (N_15469,N_15345,N_15200);
nor U15470 (N_15470,N_15333,N_15212);
or U15471 (N_15471,N_15299,N_15351);
nand U15472 (N_15472,N_15383,N_15255);
nor U15473 (N_15473,N_15393,N_15372);
or U15474 (N_15474,N_15274,N_15216);
nor U15475 (N_15475,N_15359,N_15376);
nor U15476 (N_15476,N_15364,N_15356);
nor U15477 (N_15477,N_15339,N_15269);
or U15478 (N_15478,N_15373,N_15272);
nor U15479 (N_15479,N_15228,N_15276);
or U15480 (N_15480,N_15201,N_15329);
or U15481 (N_15481,N_15347,N_15331);
xor U15482 (N_15482,N_15252,N_15217);
and U15483 (N_15483,N_15394,N_15248);
xnor U15484 (N_15484,N_15203,N_15224);
xnor U15485 (N_15485,N_15385,N_15306);
xnor U15486 (N_15486,N_15388,N_15390);
or U15487 (N_15487,N_15337,N_15374);
xor U15488 (N_15488,N_15296,N_15305);
nand U15489 (N_15489,N_15287,N_15265);
nor U15490 (N_15490,N_15284,N_15355);
nand U15491 (N_15491,N_15304,N_15227);
nor U15492 (N_15492,N_15338,N_15314);
xor U15493 (N_15493,N_15204,N_15392);
or U15494 (N_15494,N_15271,N_15220);
and U15495 (N_15495,N_15245,N_15324);
nand U15496 (N_15496,N_15318,N_15229);
xor U15497 (N_15497,N_15264,N_15280);
nand U15498 (N_15498,N_15323,N_15354);
or U15499 (N_15499,N_15230,N_15215);
or U15500 (N_15500,N_15319,N_15226);
nand U15501 (N_15501,N_15239,N_15301);
nand U15502 (N_15502,N_15225,N_15321);
or U15503 (N_15503,N_15399,N_15370);
xor U15504 (N_15504,N_15304,N_15341);
nand U15505 (N_15505,N_15373,N_15334);
or U15506 (N_15506,N_15226,N_15287);
nor U15507 (N_15507,N_15362,N_15377);
nor U15508 (N_15508,N_15361,N_15329);
or U15509 (N_15509,N_15398,N_15300);
xnor U15510 (N_15510,N_15233,N_15227);
nand U15511 (N_15511,N_15304,N_15210);
nand U15512 (N_15512,N_15227,N_15200);
xor U15513 (N_15513,N_15237,N_15337);
nand U15514 (N_15514,N_15262,N_15321);
or U15515 (N_15515,N_15394,N_15310);
nand U15516 (N_15516,N_15375,N_15232);
or U15517 (N_15517,N_15347,N_15295);
or U15518 (N_15518,N_15215,N_15243);
nand U15519 (N_15519,N_15394,N_15281);
nand U15520 (N_15520,N_15273,N_15378);
and U15521 (N_15521,N_15211,N_15239);
nor U15522 (N_15522,N_15395,N_15239);
nor U15523 (N_15523,N_15222,N_15380);
and U15524 (N_15524,N_15253,N_15348);
and U15525 (N_15525,N_15269,N_15256);
xnor U15526 (N_15526,N_15254,N_15223);
xor U15527 (N_15527,N_15351,N_15229);
xor U15528 (N_15528,N_15315,N_15347);
nand U15529 (N_15529,N_15399,N_15328);
and U15530 (N_15530,N_15297,N_15295);
and U15531 (N_15531,N_15332,N_15382);
nand U15532 (N_15532,N_15301,N_15378);
nand U15533 (N_15533,N_15239,N_15342);
and U15534 (N_15534,N_15207,N_15354);
or U15535 (N_15535,N_15328,N_15386);
nor U15536 (N_15536,N_15283,N_15246);
nor U15537 (N_15537,N_15332,N_15280);
or U15538 (N_15538,N_15229,N_15328);
xnor U15539 (N_15539,N_15232,N_15246);
nor U15540 (N_15540,N_15359,N_15342);
nor U15541 (N_15541,N_15371,N_15258);
or U15542 (N_15542,N_15274,N_15379);
nor U15543 (N_15543,N_15363,N_15391);
xor U15544 (N_15544,N_15343,N_15275);
xnor U15545 (N_15545,N_15390,N_15242);
nand U15546 (N_15546,N_15273,N_15320);
or U15547 (N_15547,N_15369,N_15370);
nand U15548 (N_15548,N_15235,N_15345);
nand U15549 (N_15549,N_15358,N_15209);
or U15550 (N_15550,N_15257,N_15314);
and U15551 (N_15551,N_15264,N_15386);
nor U15552 (N_15552,N_15351,N_15288);
and U15553 (N_15553,N_15222,N_15344);
or U15554 (N_15554,N_15296,N_15231);
xnor U15555 (N_15555,N_15213,N_15394);
xnor U15556 (N_15556,N_15252,N_15384);
nand U15557 (N_15557,N_15214,N_15367);
nand U15558 (N_15558,N_15364,N_15334);
nand U15559 (N_15559,N_15274,N_15227);
xnor U15560 (N_15560,N_15211,N_15381);
nand U15561 (N_15561,N_15238,N_15261);
nand U15562 (N_15562,N_15362,N_15311);
or U15563 (N_15563,N_15246,N_15226);
nor U15564 (N_15564,N_15375,N_15264);
nand U15565 (N_15565,N_15394,N_15349);
and U15566 (N_15566,N_15236,N_15347);
xor U15567 (N_15567,N_15320,N_15313);
nand U15568 (N_15568,N_15310,N_15393);
and U15569 (N_15569,N_15214,N_15330);
and U15570 (N_15570,N_15346,N_15296);
and U15571 (N_15571,N_15357,N_15230);
xnor U15572 (N_15572,N_15314,N_15221);
or U15573 (N_15573,N_15275,N_15357);
or U15574 (N_15574,N_15314,N_15347);
xor U15575 (N_15575,N_15206,N_15284);
and U15576 (N_15576,N_15373,N_15337);
or U15577 (N_15577,N_15274,N_15333);
xor U15578 (N_15578,N_15215,N_15270);
nor U15579 (N_15579,N_15258,N_15202);
xnor U15580 (N_15580,N_15347,N_15330);
or U15581 (N_15581,N_15225,N_15259);
nor U15582 (N_15582,N_15236,N_15331);
or U15583 (N_15583,N_15288,N_15289);
nor U15584 (N_15584,N_15247,N_15200);
and U15585 (N_15585,N_15338,N_15254);
xnor U15586 (N_15586,N_15396,N_15237);
nor U15587 (N_15587,N_15366,N_15215);
or U15588 (N_15588,N_15242,N_15389);
nand U15589 (N_15589,N_15285,N_15259);
nand U15590 (N_15590,N_15315,N_15316);
or U15591 (N_15591,N_15299,N_15396);
nand U15592 (N_15592,N_15306,N_15295);
or U15593 (N_15593,N_15291,N_15387);
nand U15594 (N_15594,N_15281,N_15397);
and U15595 (N_15595,N_15353,N_15286);
xor U15596 (N_15596,N_15209,N_15363);
xor U15597 (N_15597,N_15279,N_15323);
xnor U15598 (N_15598,N_15300,N_15269);
and U15599 (N_15599,N_15365,N_15291);
or U15600 (N_15600,N_15481,N_15521);
or U15601 (N_15601,N_15570,N_15493);
and U15602 (N_15602,N_15402,N_15465);
nand U15603 (N_15603,N_15562,N_15523);
or U15604 (N_15604,N_15573,N_15431);
nand U15605 (N_15605,N_15418,N_15507);
or U15606 (N_15606,N_15584,N_15526);
nor U15607 (N_15607,N_15408,N_15564);
nand U15608 (N_15608,N_15458,N_15425);
nand U15609 (N_15609,N_15490,N_15576);
xnor U15610 (N_15610,N_15597,N_15435);
nand U15611 (N_15611,N_15582,N_15437);
and U15612 (N_15612,N_15417,N_15532);
and U15613 (N_15613,N_15555,N_15447);
nand U15614 (N_15614,N_15580,N_15459);
or U15615 (N_15615,N_15598,N_15444);
xnor U15616 (N_15616,N_15515,N_15462);
or U15617 (N_15617,N_15478,N_15593);
nor U15618 (N_15618,N_15529,N_15571);
nor U15619 (N_15619,N_15439,N_15453);
and U15620 (N_15620,N_15494,N_15446);
nand U15621 (N_15621,N_15590,N_15499);
or U15622 (N_15622,N_15419,N_15471);
nor U15623 (N_15623,N_15544,N_15440);
nor U15624 (N_15624,N_15583,N_15401);
nand U15625 (N_15625,N_15487,N_15513);
nand U15626 (N_15626,N_15498,N_15484);
and U15627 (N_15627,N_15533,N_15579);
or U15628 (N_15628,N_15540,N_15561);
or U15629 (N_15629,N_15551,N_15543);
or U15630 (N_15630,N_15516,N_15511);
nor U15631 (N_15631,N_15438,N_15518);
xor U15632 (N_15632,N_15424,N_15483);
nor U15633 (N_15633,N_15406,N_15514);
xnor U15634 (N_15634,N_15452,N_15577);
or U15635 (N_15635,N_15448,N_15509);
nor U15636 (N_15636,N_15432,N_15434);
xor U15637 (N_15637,N_15468,N_15574);
and U15638 (N_15638,N_15457,N_15489);
or U15639 (N_15639,N_15430,N_15560);
or U15640 (N_15640,N_15488,N_15474);
xnor U15641 (N_15641,N_15569,N_15536);
nor U15642 (N_15642,N_15445,N_15528);
and U15643 (N_15643,N_15556,N_15545);
xor U15644 (N_15644,N_15589,N_15442);
nand U15645 (N_15645,N_15594,N_15491);
nor U15646 (N_15646,N_15596,N_15591);
xor U15647 (N_15647,N_15541,N_15415);
or U15648 (N_15648,N_15421,N_15512);
nand U15649 (N_15649,N_15428,N_15524);
xnor U15650 (N_15650,N_15429,N_15595);
nand U15651 (N_15651,N_15568,N_15403);
and U15652 (N_15652,N_15449,N_15531);
or U15653 (N_15653,N_15492,N_15517);
nand U15654 (N_15654,N_15522,N_15539);
nor U15655 (N_15655,N_15548,N_15405);
and U15656 (N_15656,N_15495,N_15400);
nand U15657 (N_15657,N_15411,N_15506);
nand U15658 (N_15658,N_15476,N_15479);
or U15659 (N_15659,N_15451,N_15500);
or U15660 (N_15660,N_15472,N_15423);
xnor U15661 (N_15661,N_15463,N_15588);
xor U15662 (N_15662,N_15546,N_15565);
nand U15663 (N_15663,N_15480,N_15537);
or U15664 (N_15664,N_15592,N_15534);
xnor U15665 (N_15665,N_15455,N_15443);
and U15666 (N_15666,N_15497,N_15466);
xor U15667 (N_15667,N_15510,N_15550);
xor U15668 (N_15668,N_15409,N_15585);
xor U15669 (N_15669,N_15502,N_15486);
nor U15670 (N_15670,N_15504,N_15578);
or U15671 (N_15671,N_15575,N_15549);
xnor U15672 (N_15672,N_15441,N_15460);
xnor U15673 (N_15673,N_15520,N_15436);
xor U15674 (N_15674,N_15547,N_15473);
nor U15675 (N_15675,N_15559,N_15535);
and U15676 (N_15676,N_15530,N_15505);
xnor U15677 (N_15677,N_15450,N_15566);
or U15678 (N_15678,N_15426,N_15538);
nor U15679 (N_15679,N_15477,N_15412);
nor U15680 (N_15680,N_15542,N_15422);
nand U15681 (N_15681,N_15599,N_15420);
xor U15682 (N_15682,N_15503,N_15554);
nand U15683 (N_15683,N_15414,N_15416);
nor U15684 (N_15684,N_15501,N_15558);
nand U15685 (N_15685,N_15482,N_15467);
or U15686 (N_15686,N_15525,N_15410);
nor U15687 (N_15687,N_15404,N_15519);
nand U15688 (N_15688,N_15427,N_15527);
and U15689 (N_15689,N_15433,N_15407);
nor U15690 (N_15690,N_15552,N_15563);
or U15691 (N_15691,N_15461,N_15456);
nand U15692 (N_15692,N_15587,N_15557);
and U15693 (N_15693,N_15508,N_15485);
xor U15694 (N_15694,N_15572,N_15567);
nor U15695 (N_15695,N_15475,N_15464);
nor U15696 (N_15696,N_15581,N_15454);
xor U15697 (N_15697,N_15413,N_15496);
or U15698 (N_15698,N_15553,N_15469);
nand U15699 (N_15699,N_15470,N_15586);
nor U15700 (N_15700,N_15426,N_15549);
or U15701 (N_15701,N_15420,N_15476);
nor U15702 (N_15702,N_15446,N_15503);
nor U15703 (N_15703,N_15485,N_15549);
xnor U15704 (N_15704,N_15448,N_15406);
xor U15705 (N_15705,N_15403,N_15511);
nor U15706 (N_15706,N_15573,N_15578);
and U15707 (N_15707,N_15597,N_15526);
nor U15708 (N_15708,N_15498,N_15529);
or U15709 (N_15709,N_15572,N_15437);
xor U15710 (N_15710,N_15478,N_15586);
nand U15711 (N_15711,N_15513,N_15529);
nand U15712 (N_15712,N_15477,N_15569);
and U15713 (N_15713,N_15564,N_15556);
nand U15714 (N_15714,N_15440,N_15470);
nand U15715 (N_15715,N_15458,N_15577);
or U15716 (N_15716,N_15553,N_15506);
xor U15717 (N_15717,N_15557,N_15589);
nor U15718 (N_15718,N_15543,N_15461);
xnor U15719 (N_15719,N_15552,N_15550);
and U15720 (N_15720,N_15416,N_15535);
and U15721 (N_15721,N_15512,N_15408);
or U15722 (N_15722,N_15535,N_15526);
or U15723 (N_15723,N_15432,N_15522);
xnor U15724 (N_15724,N_15451,N_15581);
nand U15725 (N_15725,N_15532,N_15517);
and U15726 (N_15726,N_15480,N_15533);
and U15727 (N_15727,N_15481,N_15422);
xor U15728 (N_15728,N_15490,N_15593);
nor U15729 (N_15729,N_15572,N_15541);
xnor U15730 (N_15730,N_15495,N_15599);
xor U15731 (N_15731,N_15564,N_15451);
or U15732 (N_15732,N_15411,N_15516);
and U15733 (N_15733,N_15523,N_15472);
nand U15734 (N_15734,N_15552,N_15501);
nand U15735 (N_15735,N_15553,N_15450);
or U15736 (N_15736,N_15567,N_15408);
nand U15737 (N_15737,N_15485,N_15444);
and U15738 (N_15738,N_15505,N_15430);
nand U15739 (N_15739,N_15590,N_15543);
and U15740 (N_15740,N_15400,N_15529);
and U15741 (N_15741,N_15412,N_15550);
or U15742 (N_15742,N_15509,N_15544);
and U15743 (N_15743,N_15593,N_15485);
nor U15744 (N_15744,N_15408,N_15413);
nor U15745 (N_15745,N_15464,N_15595);
nand U15746 (N_15746,N_15591,N_15593);
or U15747 (N_15747,N_15547,N_15526);
xnor U15748 (N_15748,N_15524,N_15527);
xor U15749 (N_15749,N_15567,N_15496);
nand U15750 (N_15750,N_15438,N_15548);
or U15751 (N_15751,N_15487,N_15423);
nand U15752 (N_15752,N_15527,N_15435);
nand U15753 (N_15753,N_15559,N_15460);
nand U15754 (N_15754,N_15517,N_15458);
or U15755 (N_15755,N_15403,N_15411);
nand U15756 (N_15756,N_15445,N_15402);
xnor U15757 (N_15757,N_15527,N_15536);
and U15758 (N_15758,N_15410,N_15575);
or U15759 (N_15759,N_15596,N_15415);
nor U15760 (N_15760,N_15592,N_15505);
and U15761 (N_15761,N_15444,N_15552);
nor U15762 (N_15762,N_15440,N_15545);
and U15763 (N_15763,N_15487,N_15575);
xor U15764 (N_15764,N_15440,N_15438);
nand U15765 (N_15765,N_15588,N_15533);
and U15766 (N_15766,N_15540,N_15459);
xor U15767 (N_15767,N_15417,N_15542);
nor U15768 (N_15768,N_15495,N_15471);
or U15769 (N_15769,N_15426,N_15512);
or U15770 (N_15770,N_15512,N_15486);
nand U15771 (N_15771,N_15546,N_15476);
and U15772 (N_15772,N_15517,N_15521);
nand U15773 (N_15773,N_15532,N_15496);
nand U15774 (N_15774,N_15574,N_15595);
nand U15775 (N_15775,N_15415,N_15458);
nor U15776 (N_15776,N_15556,N_15429);
or U15777 (N_15777,N_15436,N_15509);
and U15778 (N_15778,N_15472,N_15512);
or U15779 (N_15779,N_15429,N_15570);
xnor U15780 (N_15780,N_15474,N_15410);
xnor U15781 (N_15781,N_15415,N_15506);
xor U15782 (N_15782,N_15598,N_15443);
and U15783 (N_15783,N_15577,N_15540);
xnor U15784 (N_15784,N_15454,N_15536);
xor U15785 (N_15785,N_15520,N_15552);
nand U15786 (N_15786,N_15446,N_15473);
nand U15787 (N_15787,N_15537,N_15527);
nand U15788 (N_15788,N_15426,N_15499);
xnor U15789 (N_15789,N_15471,N_15553);
nand U15790 (N_15790,N_15445,N_15437);
nor U15791 (N_15791,N_15471,N_15590);
nor U15792 (N_15792,N_15446,N_15496);
and U15793 (N_15793,N_15556,N_15483);
xnor U15794 (N_15794,N_15508,N_15443);
or U15795 (N_15795,N_15571,N_15533);
nand U15796 (N_15796,N_15401,N_15480);
nor U15797 (N_15797,N_15528,N_15546);
or U15798 (N_15798,N_15516,N_15478);
nor U15799 (N_15799,N_15579,N_15518);
xnor U15800 (N_15800,N_15632,N_15621);
xnor U15801 (N_15801,N_15760,N_15716);
or U15802 (N_15802,N_15757,N_15660);
xnor U15803 (N_15803,N_15623,N_15655);
or U15804 (N_15804,N_15736,N_15616);
nand U15805 (N_15805,N_15618,N_15619);
or U15806 (N_15806,N_15725,N_15675);
or U15807 (N_15807,N_15723,N_15607);
nand U15808 (N_15808,N_15764,N_15708);
or U15809 (N_15809,N_15696,N_15690);
xnor U15810 (N_15810,N_15699,N_15653);
xnor U15811 (N_15811,N_15729,N_15719);
or U15812 (N_15812,N_15768,N_15672);
or U15813 (N_15813,N_15774,N_15783);
and U15814 (N_15814,N_15628,N_15746);
and U15815 (N_15815,N_15649,N_15750);
xor U15816 (N_15816,N_15674,N_15798);
nor U15817 (N_15817,N_15691,N_15638);
or U15818 (N_15818,N_15755,N_15778);
xor U15819 (N_15819,N_15753,N_15614);
and U15820 (N_15820,N_15600,N_15782);
nand U15821 (N_15821,N_15777,N_15739);
nand U15822 (N_15822,N_15605,N_15694);
nor U15823 (N_15823,N_15609,N_15771);
nand U15824 (N_15824,N_15667,N_15790);
or U15825 (N_15825,N_15787,N_15712);
and U15826 (N_15826,N_15747,N_15652);
or U15827 (N_15827,N_15610,N_15637);
nor U15828 (N_15828,N_15612,N_15641);
or U15829 (N_15829,N_15608,N_15743);
nand U15830 (N_15830,N_15733,N_15727);
and U15831 (N_15831,N_15715,N_15786);
nor U15832 (N_15832,N_15713,N_15745);
or U15833 (N_15833,N_15781,N_15681);
or U15834 (N_15834,N_15766,N_15748);
and U15835 (N_15835,N_15758,N_15737);
nand U15836 (N_15836,N_15684,N_15731);
or U15837 (N_15837,N_15689,N_15756);
nor U15838 (N_15838,N_15680,N_15685);
and U15839 (N_15839,N_15738,N_15613);
nand U15840 (N_15840,N_15763,N_15668);
or U15841 (N_15841,N_15686,N_15657);
or U15842 (N_15842,N_15794,N_15734);
nand U15843 (N_15843,N_15617,N_15629);
nor U15844 (N_15844,N_15742,N_15700);
nor U15845 (N_15845,N_15762,N_15604);
xor U15846 (N_15846,N_15722,N_15635);
nand U15847 (N_15847,N_15773,N_15759);
and U15848 (N_15848,N_15706,N_15669);
and U15849 (N_15849,N_15606,N_15772);
xnor U15850 (N_15850,N_15761,N_15789);
and U15851 (N_15851,N_15648,N_15702);
xor U15852 (N_15852,N_15697,N_15640);
or U15853 (N_15853,N_15647,N_15797);
nand U15854 (N_15854,N_15658,N_15650);
nand U15855 (N_15855,N_15665,N_15707);
and U15856 (N_15856,N_15646,N_15688);
xnor U15857 (N_15857,N_15779,N_15683);
nor U15858 (N_15858,N_15661,N_15677);
and U15859 (N_15859,N_15726,N_15780);
xnor U15860 (N_15860,N_15717,N_15670);
nand U15861 (N_15861,N_15754,N_15718);
and U15862 (N_15862,N_15631,N_15732);
xor U15863 (N_15863,N_15744,N_15749);
or U15864 (N_15864,N_15626,N_15704);
nand U15865 (N_15865,N_15662,N_15633);
or U15866 (N_15866,N_15791,N_15703);
and U15867 (N_15867,N_15721,N_15687);
xnor U15868 (N_15868,N_15678,N_15642);
nor U15869 (N_15869,N_15735,N_15651);
xnor U15870 (N_15870,N_15785,N_15793);
and U15871 (N_15871,N_15714,N_15784);
xor U15872 (N_15872,N_15692,N_15656);
nand U15873 (N_15873,N_15644,N_15636);
or U15874 (N_15874,N_15671,N_15679);
or U15875 (N_15875,N_15602,N_15625);
nor U15876 (N_15876,N_15615,N_15711);
and U15877 (N_15877,N_15601,N_15799);
xor U15878 (N_15878,N_15659,N_15724);
or U15879 (N_15879,N_15695,N_15620);
or U15880 (N_15880,N_15682,N_15630);
xnor U15881 (N_15881,N_15709,N_15765);
or U15882 (N_15882,N_15795,N_15639);
and U15883 (N_15883,N_15751,N_15622);
and U15884 (N_15884,N_15740,N_15664);
xor U15885 (N_15885,N_15770,N_15730);
nand U15886 (N_15886,N_15728,N_15701);
nand U15887 (N_15887,N_15663,N_15627);
xnor U15888 (N_15888,N_15676,N_15720);
xor U15889 (N_15889,N_15752,N_15767);
or U15890 (N_15890,N_15788,N_15769);
nand U15891 (N_15891,N_15710,N_15693);
xor U15892 (N_15892,N_15775,N_15673);
or U15893 (N_15893,N_15666,N_15603);
nand U15894 (N_15894,N_15705,N_15741);
and U15895 (N_15895,N_15792,N_15645);
nand U15896 (N_15896,N_15776,N_15698);
and U15897 (N_15897,N_15634,N_15643);
nand U15898 (N_15898,N_15624,N_15796);
xor U15899 (N_15899,N_15654,N_15611);
nand U15900 (N_15900,N_15649,N_15640);
xnor U15901 (N_15901,N_15742,N_15693);
and U15902 (N_15902,N_15720,N_15635);
or U15903 (N_15903,N_15662,N_15657);
nand U15904 (N_15904,N_15776,N_15630);
xor U15905 (N_15905,N_15781,N_15705);
or U15906 (N_15906,N_15712,N_15660);
or U15907 (N_15907,N_15646,N_15768);
nand U15908 (N_15908,N_15777,N_15672);
nor U15909 (N_15909,N_15711,N_15650);
and U15910 (N_15910,N_15780,N_15652);
nand U15911 (N_15911,N_15618,N_15749);
or U15912 (N_15912,N_15696,N_15701);
xnor U15913 (N_15913,N_15682,N_15635);
xor U15914 (N_15914,N_15739,N_15732);
or U15915 (N_15915,N_15777,N_15776);
nor U15916 (N_15916,N_15709,N_15716);
xor U15917 (N_15917,N_15786,N_15681);
nor U15918 (N_15918,N_15743,N_15658);
nand U15919 (N_15919,N_15610,N_15703);
and U15920 (N_15920,N_15600,N_15751);
nor U15921 (N_15921,N_15618,N_15602);
nor U15922 (N_15922,N_15767,N_15634);
and U15923 (N_15923,N_15610,N_15658);
or U15924 (N_15924,N_15655,N_15783);
nor U15925 (N_15925,N_15798,N_15666);
xnor U15926 (N_15926,N_15605,N_15756);
and U15927 (N_15927,N_15639,N_15676);
or U15928 (N_15928,N_15735,N_15729);
or U15929 (N_15929,N_15705,N_15611);
and U15930 (N_15930,N_15747,N_15793);
nor U15931 (N_15931,N_15783,N_15745);
nand U15932 (N_15932,N_15606,N_15671);
and U15933 (N_15933,N_15755,N_15795);
xor U15934 (N_15934,N_15792,N_15692);
xnor U15935 (N_15935,N_15714,N_15660);
nor U15936 (N_15936,N_15747,N_15791);
and U15937 (N_15937,N_15749,N_15724);
nand U15938 (N_15938,N_15738,N_15614);
and U15939 (N_15939,N_15637,N_15605);
and U15940 (N_15940,N_15778,N_15703);
nor U15941 (N_15941,N_15795,N_15614);
or U15942 (N_15942,N_15740,N_15610);
and U15943 (N_15943,N_15762,N_15610);
xnor U15944 (N_15944,N_15690,N_15692);
nand U15945 (N_15945,N_15706,N_15623);
and U15946 (N_15946,N_15615,N_15797);
nor U15947 (N_15947,N_15790,N_15600);
or U15948 (N_15948,N_15773,N_15639);
and U15949 (N_15949,N_15701,N_15748);
nand U15950 (N_15950,N_15639,N_15718);
nand U15951 (N_15951,N_15606,N_15651);
nand U15952 (N_15952,N_15788,N_15796);
nand U15953 (N_15953,N_15612,N_15772);
nand U15954 (N_15954,N_15783,N_15703);
nor U15955 (N_15955,N_15655,N_15798);
or U15956 (N_15956,N_15658,N_15611);
nor U15957 (N_15957,N_15632,N_15606);
and U15958 (N_15958,N_15759,N_15730);
xnor U15959 (N_15959,N_15770,N_15712);
and U15960 (N_15960,N_15683,N_15691);
nor U15961 (N_15961,N_15785,N_15721);
nand U15962 (N_15962,N_15714,N_15617);
or U15963 (N_15963,N_15630,N_15716);
nand U15964 (N_15964,N_15607,N_15743);
nand U15965 (N_15965,N_15608,N_15790);
and U15966 (N_15966,N_15714,N_15719);
xnor U15967 (N_15967,N_15702,N_15750);
and U15968 (N_15968,N_15659,N_15662);
or U15969 (N_15969,N_15667,N_15698);
xor U15970 (N_15970,N_15731,N_15740);
or U15971 (N_15971,N_15632,N_15657);
nand U15972 (N_15972,N_15649,N_15671);
nor U15973 (N_15973,N_15684,N_15738);
nor U15974 (N_15974,N_15682,N_15698);
nand U15975 (N_15975,N_15786,N_15644);
nand U15976 (N_15976,N_15789,N_15794);
or U15977 (N_15977,N_15755,N_15791);
nand U15978 (N_15978,N_15647,N_15681);
nor U15979 (N_15979,N_15786,N_15712);
and U15980 (N_15980,N_15682,N_15763);
or U15981 (N_15981,N_15665,N_15762);
or U15982 (N_15982,N_15692,N_15731);
or U15983 (N_15983,N_15695,N_15704);
xor U15984 (N_15984,N_15642,N_15672);
nor U15985 (N_15985,N_15657,N_15693);
nand U15986 (N_15986,N_15750,N_15758);
and U15987 (N_15987,N_15764,N_15611);
xnor U15988 (N_15988,N_15690,N_15658);
nand U15989 (N_15989,N_15688,N_15773);
nor U15990 (N_15990,N_15661,N_15617);
and U15991 (N_15991,N_15768,N_15690);
or U15992 (N_15992,N_15655,N_15741);
nor U15993 (N_15993,N_15733,N_15661);
and U15994 (N_15994,N_15608,N_15621);
and U15995 (N_15995,N_15664,N_15657);
or U15996 (N_15996,N_15676,N_15747);
nor U15997 (N_15997,N_15763,N_15708);
or U15998 (N_15998,N_15694,N_15797);
nor U15999 (N_15999,N_15601,N_15641);
or U16000 (N_16000,N_15856,N_15848);
nor U16001 (N_16001,N_15801,N_15835);
xnor U16002 (N_16002,N_15991,N_15807);
xnor U16003 (N_16003,N_15983,N_15923);
xnor U16004 (N_16004,N_15827,N_15960);
nand U16005 (N_16005,N_15888,N_15806);
or U16006 (N_16006,N_15855,N_15828);
or U16007 (N_16007,N_15915,N_15861);
nor U16008 (N_16008,N_15805,N_15898);
nor U16009 (N_16009,N_15867,N_15893);
nor U16010 (N_16010,N_15813,N_15838);
nand U16011 (N_16011,N_15850,N_15945);
and U16012 (N_16012,N_15944,N_15843);
nor U16013 (N_16013,N_15953,N_15849);
nand U16014 (N_16014,N_15975,N_15882);
or U16015 (N_16015,N_15967,N_15938);
or U16016 (N_16016,N_15876,N_15917);
or U16017 (N_16017,N_15931,N_15844);
and U16018 (N_16018,N_15878,N_15842);
and U16019 (N_16019,N_15839,N_15971);
nor U16020 (N_16020,N_15961,N_15852);
and U16021 (N_16021,N_15851,N_15918);
xor U16022 (N_16022,N_15956,N_15997);
or U16023 (N_16023,N_15959,N_15815);
xor U16024 (N_16024,N_15955,N_15820);
nor U16025 (N_16025,N_15906,N_15934);
nand U16026 (N_16026,N_15845,N_15870);
and U16027 (N_16027,N_15987,N_15834);
and U16028 (N_16028,N_15930,N_15885);
nand U16029 (N_16029,N_15872,N_15899);
nor U16030 (N_16030,N_15869,N_15884);
nand U16031 (N_16031,N_15935,N_15940);
or U16032 (N_16032,N_15816,N_15988);
xnor U16033 (N_16033,N_15963,N_15980);
nand U16034 (N_16034,N_15951,N_15920);
or U16035 (N_16035,N_15912,N_15803);
or U16036 (N_16036,N_15978,N_15836);
or U16037 (N_16037,N_15986,N_15868);
or U16038 (N_16038,N_15990,N_15942);
xor U16039 (N_16039,N_15947,N_15928);
nand U16040 (N_16040,N_15857,N_15901);
nor U16041 (N_16041,N_15823,N_15907);
or U16042 (N_16042,N_15933,N_15913);
or U16043 (N_16043,N_15896,N_15902);
and U16044 (N_16044,N_15969,N_15995);
nand U16045 (N_16045,N_15859,N_15883);
and U16046 (N_16046,N_15965,N_15922);
xnor U16047 (N_16047,N_15874,N_15911);
xnor U16048 (N_16048,N_15804,N_15858);
nor U16049 (N_16049,N_15962,N_15829);
or U16050 (N_16050,N_15847,N_15921);
xnor U16051 (N_16051,N_15914,N_15808);
nand U16052 (N_16052,N_15841,N_15900);
xor U16053 (N_16053,N_15864,N_15817);
or U16054 (N_16054,N_15974,N_15826);
xor U16055 (N_16055,N_15875,N_15863);
or U16056 (N_16056,N_15948,N_15865);
nor U16057 (N_16057,N_15905,N_15927);
or U16058 (N_16058,N_15814,N_15985);
or U16059 (N_16059,N_15891,N_15998);
xor U16060 (N_16060,N_15964,N_15831);
xor U16061 (N_16061,N_15825,N_15818);
or U16062 (N_16062,N_15809,N_15968);
nor U16063 (N_16063,N_15994,N_15887);
nand U16064 (N_16064,N_15800,N_15866);
nand U16065 (N_16065,N_15984,N_15954);
or U16066 (N_16066,N_15993,N_15970);
and U16067 (N_16067,N_15949,N_15976);
nor U16068 (N_16068,N_15925,N_15924);
xor U16069 (N_16069,N_15910,N_15939);
nor U16070 (N_16070,N_15904,N_15981);
nor U16071 (N_16071,N_15821,N_15941);
xnor U16072 (N_16072,N_15919,N_15819);
nand U16073 (N_16073,N_15890,N_15946);
or U16074 (N_16074,N_15812,N_15926);
or U16075 (N_16075,N_15811,N_15889);
nor U16076 (N_16076,N_15862,N_15873);
nand U16077 (N_16077,N_15886,N_15802);
and U16078 (N_16078,N_15895,N_15982);
xnor U16079 (N_16079,N_15871,N_15881);
nor U16080 (N_16080,N_15822,N_15854);
or U16081 (N_16081,N_15860,N_15832);
nand U16082 (N_16082,N_15973,N_15996);
nor U16083 (N_16083,N_15992,N_15833);
xnor U16084 (N_16084,N_15846,N_15972);
and U16085 (N_16085,N_15999,N_15903);
nor U16086 (N_16086,N_15830,N_15880);
or U16087 (N_16087,N_15916,N_15957);
nor U16088 (N_16088,N_15909,N_15937);
nand U16089 (N_16089,N_15877,N_15879);
and U16090 (N_16090,N_15966,N_15977);
xnor U16091 (N_16091,N_15894,N_15908);
nor U16092 (N_16092,N_15979,N_15932);
xor U16093 (N_16093,N_15824,N_15952);
nand U16094 (N_16094,N_15840,N_15950);
nor U16095 (N_16095,N_15853,N_15958);
nand U16096 (N_16096,N_15936,N_15929);
and U16097 (N_16097,N_15989,N_15943);
xnor U16098 (N_16098,N_15897,N_15892);
nor U16099 (N_16099,N_15810,N_15837);
or U16100 (N_16100,N_15965,N_15839);
and U16101 (N_16101,N_15939,N_15865);
xor U16102 (N_16102,N_15825,N_15949);
xnor U16103 (N_16103,N_15924,N_15993);
and U16104 (N_16104,N_15880,N_15896);
nand U16105 (N_16105,N_15885,N_15991);
and U16106 (N_16106,N_15868,N_15804);
and U16107 (N_16107,N_15938,N_15895);
nor U16108 (N_16108,N_15990,N_15811);
or U16109 (N_16109,N_15969,N_15871);
or U16110 (N_16110,N_15853,N_15943);
or U16111 (N_16111,N_15891,N_15865);
xor U16112 (N_16112,N_15850,N_15842);
nand U16113 (N_16113,N_15938,N_15864);
or U16114 (N_16114,N_15964,N_15962);
nor U16115 (N_16115,N_15950,N_15970);
xor U16116 (N_16116,N_15871,N_15928);
nor U16117 (N_16117,N_15941,N_15970);
xor U16118 (N_16118,N_15800,N_15824);
xnor U16119 (N_16119,N_15892,N_15821);
or U16120 (N_16120,N_15932,N_15910);
or U16121 (N_16121,N_15927,N_15978);
or U16122 (N_16122,N_15953,N_15918);
nor U16123 (N_16123,N_15940,N_15817);
nand U16124 (N_16124,N_15854,N_15852);
nor U16125 (N_16125,N_15921,N_15843);
nor U16126 (N_16126,N_15932,N_15937);
and U16127 (N_16127,N_15878,N_15872);
and U16128 (N_16128,N_15997,N_15865);
xnor U16129 (N_16129,N_15998,N_15953);
xor U16130 (N_16130,N_15861,N_15957);
and U16131 (N_16131,N_15966,N_15816);
or U16132 (N_16132,N_15895,N_15846);
and U16133 (N_16133,N_15801,N_15993);
and U16134 (N_16134,N_15842,N_15855);
nor U16135 (N_16135,N_15811,N_15817);
or U16136 (N_16136,N_15951,N_15973);
nand U16137 (N_16137,N_15882,N_15895);
xor U16138 (N_16138,N_15816,N_15970);
and U16139 (N_16139,N_15946,N_15926);
and U16140 (N_16140,N_15965,N_15854);
xor U16141 (N_16141,N_15992,N_15975);
nor U16142 (N_16142,N_15932,N_15881);
or U16143 (N_16143,N_15867,N_15859);
and U16144 (N_16144,N_15942,N_15979);
and U16145 (N_16145,N_15915,N_15851);
and U16146 (N_16146,N_15921,N_15881);
nand U16147 (N_16147,N_15955,N_15841);
or U16148 (N_16148,N_15875,N_15849);
xnor U16149 (N_16149,N_15956,N_15803);
nand U16150 (N_16150,N_15999,N_15996);
xnor U16151 (N_16151,N_15898,N_15870);
and U16152 (N_16152,N_15826,N_15872);
nand U16153 (N_16153,N_15878,N_15953);
nor U16154 (N_16154,N_15924,N_15948);
nand U16155 (N_16155,N_15875,N_15873);
and U16156 (N_16156,N_15897,N_15858);
and U16157 (N_16157,N_15802,N_15959);
and U16158 (N_16158,N_15961,N_15979);
xor U16159 (N_16159,N_15864,N_15950);
xor U16160 (N_16160,N_15995,N_15866);
nand U16161 (N_16161,N_15905,N_15917);
and U16162 (N_16162,N_15984,N_15854);
xor U16163 (N_16163,N_15887,N_15988);
and U16164 (N_16164,N_15975,N_15861);
nor U16165 (N_16165,N_15950,N_15832);
or U16166 (N_16166,N_15948,N_15815);
nor U16167 (N_16167,N_15941,N_15816);
and U16168 (N_16168,N_15883,N_15916);
nor U16169 (N_16169,N_15912,N_15850);
and U16170 (N_16170,N_15841,N_15818);
or U16171 (N_16171,N_15901,N_15858);
nand U16172 (N_16172,N_15952,N_15941);
nor U16173 (N_16173,N_15983,N_15879);
and U16174 (N_16174,N_15945,N_15944);
and U16175 (N_16175,N_15804,N_15890);
xor U16176 (N_16176,N_15924,N_15801);
xor U16177 (N_16177,N_15872,N_15956);
and U16178 (N_16178,N_15876,N_15892);
nor U16179 (N_16179,N_15830,N_15970);
nand U16180 (N_16180,N_15971,N_15882);
nor U16181 (N_16181,N_15853,N_15830);
and U16182 (N_16182,N_15992,N_15885);
nand U16183 (N_16183,N_15832,N_15993);
nor U16184 (N_16184,N_15817,N_15903);
nor U16185 (N_16185,N_15995,N_15929);
nand U16186 (N_16186,N_15948,N_15986);
nand U16187 (N_16187,N_15949,N_15851);
nor U16188 (N_16188,N_15930,N_15836);
nand U16189 (N_16189,N_15910,N_15953);
nand U16190 (N_16190,N_15971,N_15895);
or U16191 (N_16191,N_15880,N_15877);
xor U16192 (N_16192,N_15886,N_15823);
xor U16193 (N_16193,N_15948,N_15826);
nor U16194 (N_16194,N_15999,N_15918);
xnor U16195 (N_16195,N_15933,N_15976);
xor U16196 (N_16196,N_15885,N_15824);
nand U16197 (N_16197,N_15931,N_15963);
xor U16198 (N_16198,N_15890,N_15990);
xor U16199 (N_16199,N_15891,N_15911);
nand U16200 (N_16200,N_16116,N_16152);
or U16201 (N_16201,N_16100,N_16015);
xor U16202 (N_16202,N_16041,N_16154);
nor U16203 (N_16203,N_16123,N_16143);
xnor U16204 (N_16204,N_16137,N_16027);
nand U16205 (N_16205,N_16058,N_16082);
nand U16206 (N_16206,N_16102,N_16035);
nor U16207 (N_16207,N_16159,N_16182);
and U16208 (N_16208,N_16156,N_16008);
and U16209 (N_16209,N_16083,N_16073);
nor U16210 (N_16210,N_16016,N_16090);
nand U16211 (N_16211,N_16032,N_16080);
or U16212 (N_16212,N_16050,N_16163);
xnor U16213 (N_16213,N_16081,N_16071);
nand U16214 (N_16214,N_16107,N_16186);
and U16215 (N_16215,N_16004,N_16070);
nand U16216 (N_16216,N_16195,N_16164);
xnor U16217 (N_16217,N_16197,N_16108);
nor U16218 (N_16218,N_16188,N_16088);
and U16219 (N_16219,N_16181,N_16189);
xor U16220 (N_16220,N_16112,N_16003);
nor U16221 (N_16221,N_16104,N_16007);
or U16222 (N_16222,N_16132,N_16084);
xnor U16223 (N_16223,N_16130,N_16095);
xor U16224 (N_16224,N_16006,N_16078);
or U16225 (N_16225,N_16134,N_16075);
nor U16226 (N_16226,N_16117,N_16145);
or U16227 (N_16227,N_16039,N_16149);
or U16228 (N_16228,N_16002,N_16093);
and U16229 (N_16229,N_16063,N_16165);
xnor U16230 (N_16230,N_16173,N_16171);
nand U16231 (N_16231,N_16185,N_16176);
nand U16232 (N_16232,N_16076,N_16061);
xnor U16233 (N_16233,N_16120,N_16036);
nor U16234 (N_16234,N_16121,N_16133);
nand U16235 (N_16235,N_16119,N_16077);
or U16236 (N_16236,N_16045,N_16018);
nand U16237 (N_16237,N_16196,N_16001);
nor U16238 (N_16238,N_16177,N_16193);
xnor U16239 (N_16239,N_16109,N_16026);
xor U16240 (N_16240,N_16122,N_16151);
or U16241 (N_16241,N_16030,N_16037);
or U16242 (N_16242,N_16013,N_16067);
nor U16243 (N_16243,N_16113,N_16064);
nand U16244 (N_16244,N_16147,N_16072);
nor U16245 (N_16245,N_16153,N_16166);
nand U16246 (N_16246,N_16025,N_16011);
and U16247 (N_16247,N_16172,N_16146);
or U16248 (N_16248,N_16128,N_16096);
nand U16249 (N_16249,N_16161,N_16180);
or U16250 (N_16250,N_16136,N_16126);
nand U16251 (N_16251,N_16135,N_16158);
xor U16252 (N_16252,N_16056,N_16183);
nand U16253 (N_16253,N_16057,N_16010);
or U16254 (N_16254,N_16139,N_16065);
xor U16255 (N_16255,N_16097,N_16044);
or U16256 (N_16256,N_16019,N_16020);
xor U16257 (N_16257,N_16021,N_16086);
or U16258 (N_16258,N_16052,N_16051);
nor U16259 (N_16259,N_16029,N_16110);
nor U16260 (N_16260,N_16014,N_16190);
or U16261 (N_16261,N_16114,N_16033);
or U16262 (N_16262,N_16024,N_16111);
and U16263 (N_16263,N_16142,N_16048);
or U16264 (N_16264,N_16184,N_16055);
and U16265 (N_16265,N_16160,N_16125);
and U16266 (N_16266,N_16047,N_16099);
xor U16267 (N_16267,N_16169,N_16103);
nand U16268 (N_16268,N_16144,N_16157);
and U16269 (N_16269,N_16167,N_16101);
and U16270 (N_16270,N_16060,N_16092);
nor U16271 (N_16271,N_16162,N_16066);
or U16272 (N_16272,N_16148,N_16040);
xor U16273 (N_16273,N_16046,N_16068);
xor U16274 (N_16274,N_16106,N_16105);
nor U16275 (N_16275,N_16138,N_16028);
and U16276 (N_16276,N_16062,N_16054);
and U16277 (N_16277,N_16031,N_16053);
and U16278 (N_16278,N_16098,N_16175);
and U16279 (N_16279,N_16191,N_16198);
and U16280 (N_16280,N_16091,N_16174);
or U16281 (N_16281,N_16049,N_16192);
or U16282 (N_16282,N_16155,N_16127);
nand U16283 (N_16283,N_16087,N_16179);
or U16284 (N_16284,N_16009,N_16194);
xnor U16285 (N_16285,N_16043,N_16094);
nand U16286 (N_16286,N_16089,N_16059);
and U16287 (N_16287,N_16131,N_16038);
or U16288 (N_16288,N_16042,N_16022);
and U16289 (N_16289,N_16085,N_16118);
nand U16290 (N_16290,N_16168,N_16199);
or U16291 (N_16291,N_16034,N_16012);
or U16292 (N_16292,N_16129,N_16079);
and U16293 (N_16293,N_16115,N_16124);
or U16294 (N_16294,N_16074,N_16140);
nand U16295 (N_16295,N_16187,N_16150);
xor U16296 (N_16296,N_16141,N_16069);
and U16297 (N_16297,N_16178,N_16023);
or U16298 (N_16298,N_16005,N_16000);
nand U16299 (N_16299,N_16017,N_16170);
xnor U16300 (N_16300,N_16149,N_16083);
nor U16301 (N_16301,N_16077,N_16055);
or U16302 (N_16302,N_16003,N_16044);
and U16303 (N_16303,N_16137,N_16195);
or U16304 (N_16304,N_16082,N_16106);
xor U16305 (N_16305,N_16046,N_16001);
and U16306 (N_16306,N_16152,N_16151);
xor U16307 (N_16307,N_16148,N_16017);
or U16308 (N_16308,N_16159,N_16152);
and U16309 (N_16309,N_16194,N_16123);
and U16310 (N_16310,N_16128,N_16032);
or U16311 (N_16311,N_16017,N_16048);
or U16312 (N_16312,N_16127,N_16007);
nand U16313 (N_16313,N_16062,N_16086);
nand U16314 (N_16314,N_16074,N_16110);
xnor U16315 (N_16315,N_16053,N_16177);
xnor U16316 (N_16316,N_16056,N_16079);
and U16317 (N_16317,N_16077,N_16171);
xnor U16318 (N_16318,N_16005,N_16081);
or U16319 (N_16319,N_16154,N_16089);
xnor U16320 (N_16320,N_16160,N_16116);
nor U16321 (N_16321,N_16079,N_16077);
nand U16322 (N_16322,N_16187,N_16174);
and U16323 (N_16323,N_16069,N_16075);
nor U16324 (N_16324,N_16169,N_16071);
nor U16325 (N_16325,N_16066,N_16126);
and U16326 (N_16326,N_16064,N_16187);
nor U16327 (N_16327,N_16070,N_16015);
nand U16328 (N_16328,N_16019,N_16095);
nor U16329 (N_16329,N_16018,N_16011);
nand U16330 (N_16330,N_16126,N_16045);
xnor U16331 (N_16331,N_16104,N_16146);
nand U16332 (N_16332,N_16145,N_16153);
xor U16333 (N_16333,N_16176,N_16043);
and U16334 (N_16334,N_16129,N_16084);
and U16335 (N_16335,N_16161,N_16171);
and U16336 (N_16336,N_16018,N_16124);
nor U16337 (N_16337,N_16124,N_16157);
nand U16338 (N_16338,N_16049,N_16148);
and U16339 (N_16339,N_16143,N_16094);
xor U16340 (N_16340,N_16124,N_16068);
or U16341 (N_16341,N_16145,N_16069);
and U16342 (N_16342,N_16127,N_16133);
and U16343 (N_16343,N_16187,N_16134);
nor U16344 (N_16344,N_16159,N_16102);
xnor U16345 (N_16345,N_16105,N_16158);
nor U16346 (N_16346,N_16189,N_16136);
or U16347 (N_16347,N_16082,N_16010);
xnor U16348 (N_16348,N_16117,N_16005);
nand U16349 (N_16349,N_16024,N_16016);
nand U16350 (N_16350,N_16117,N_16044);
nand U16351 (N_16351,N_16055,N_16094);
nand U16352 (N_16352,N_16170,N_16184);
nand U16353 (N_16353,N_16166,N_16040);
nand U16354 (N_16354,N_16163,N_16032);
nor U16355 (N_16355,N_16040,N_16016);
xor U16356 (N_16356,N_16126,N_16065);
and U16357 (N_16357,N_16063,N_16142);
and U16358 (N_16358,N_16091,N_16118);
or U16359 (N_16359,N_16179,N_16078);
nor U16360 (N_16360,N_16071,N_16183);
nand U16361 (N_16361,N_16147,N_16094);
or U16362 (N_16362,N_16023,N_16161);
nand U16363 (N_16363,N_16044,N_16009);
nand U16364 (N_16364,N_16090,N_16123);
xor U16365 (N_16365,N_16057,N_16088);
nand U16366 (N_16366,N_16191,N_16013);
and U16367 (N_16367,N_16069,N_16157);
nand U16368 (N_16368,N_16189,N_16137);
or U16369 (N_16369,N_16030,N_16059);
xnor U16370 (N_16370,N_16159,N_16082);
nand U16371 (N_16371,N_16005,N_16192);
or U16372 (N_16372,N_16033,N_16152);
xnor U16373 (N_16373,N_16055,N_16023);
nor U16374 (N_16374,N_16020,N_16158);
and U16375 (N_16375,N_16198,N_16091);
nand U16376 (N_16376,N_16124,N_16081);
xnor U16377 (N_16377,N_16174,N_16059);
xor U16378 (N_16378,N_16102,N_16146);
xor U16379 (N_16379,N_16071,N_16113);
xnor U16380 (N_16380,N_16150,N_16194);
nand U16381 (N_16381,N_16185,N_16116);
or U16382 (N_16382,N_16101,N_16003);
xor U16383 (N_16383,N_16148,N_16122);
and U16384 (N_16384,N_16024,N_16070);
xnor U16385 (N_16385,N_16089,N_16118);
nor U16386 (N_16386,N_16139,N_16072);
nand U16387 (N_16387,N_16168,N_16188);
or U16388 (N_16388,N_16143,N_16074);
and U16389 (N_16389,N_16037,N_16047);
xor U16390 (N_16390,N_16102,N_16135);
nand U16391 (N_16391,N_16142,N_16130);
nor U16392 (N_16392,N_16028,N_16186);
xor U16393 (N_16393,N_16142,N_16151);
nand U16394 (N_16394,N_16082,N_16181);
nor U16395 (N_16395,N_16168,N_16174);
nand U16396 (N_16396,N_16047,N_16147);
and U16397 (N_16397,N_16099,N_16153);
or U16398 (N_16398,N_16038,N_16094);
or U16399 (N_16399,N_16159,N_16195);
xor U16400 (N_16400,N_16386,N_16327);
xor U16401 (N_16401,N_16261,N_16213);
xor U16402 (N_16402,N_16267,N_16361);
nand U16403 (N_16403,N_16339,N_16312);
or U16404 (N_16404,N_16342,N_16380);
nor U16405 (N_16405,N_16337,N_16377);
and U16406 (N_16406,N_16356,N_16202);
or U16407 (N_16407,N_16371,N_16279);
nor U16408 (N_16408,N_16247,N_16310);
xnor U16409 (N_16409,N_16203,N_16357);
and U16410 (N_16410,N_16262,N_16218);
xor U16411 (N_16411,N_16311,N_16334);
xnor U16412 (N_16412,N_16251,N_16200);
or U16413 (N_16413,N_16393,N_16343);
xor U16414 (N_16414,N_16244,N_16346);
or U16415 (N_16415,N_16300,N_16397);
and U16416 (N_16416,N_16323,N_16225);
nor U16417 (N_16417,N_16298,N_16389);
or U16418 (N_16418,N_16315,N_16217);
xnor U16419 (N_16419,N_16235,N_16201);
nor U16420 (N_16420,N_16350,N_16347);
xor U16421 (N_16421,N_16237,N_16272);
and U16422 (N_16422,N_16212,N_16306);
and U16423 (N_16423,N_16216,N_16324);
and U16424 (N_16424,N_16253,N_16211);
or U16425 (N_16425,N_16325,N_16336);
xor U16426 (N_16426,N_16234,N_16372);
nand U16427 (N_16427,N_16296,N_16359);
and U16428 (N_16428,N_16264,N_16290);
and U16429 (N_16429,N_16326,N_16246);
nand U16430 (N_16430,N_16270,N_16275);
nand U16431 (N_16431,N_16266,N_16369);
or U16432 (N_16432,N_16368,N_16238);
or U16433 (N_16433,N_16245,N_16373);
nand U16434 (N_16434,N_16243,N_16291);
nor U16435 (N_16435,N_16385,N_16379);
nand U16436 (N_16436,N_16332,N_16257);
and U16437 (N_16437,N_16233,N_16320);
or U16438 (N_16438,N_16208,N_16232);
xnor U16439 (N_16439,N_16329,N_16220);
nor U16440 (N_16440,N_16294,N_16219);
nor U16441 (N_16441,N_16252,N_16207);
nand U16442 (N_16442,N_16328,N_16285);
and U16443 (N_16443,N_16307,N_16249);
nor U16444 (N_16444,N_16367,N_16283);
or U16445 (N_16445,N_16317,N_16231);
or U16446 (N_16446,N_16210,N_16351);
nand U16447 (N_16447,N_16333,N_16378);
nor U16448 (N_16448,N_16281,N_16365);
nor U16449 (N_16449,N_16360,N_16230);
nor U16450 (N_16450,N_16286,N_16354);
xor U16451 (N_16451,N_16364,N_16239);
and U16452 (N_16452,N_16394,N_16215);
nor U16453 (N_16453,N_16335,N_16288);
nor U16454 (N_16454,N_16277,N_16299);
nand U16455 (N_16455,N_16370,N_16301);
and U16456 (N_16456,N_16255,N_16304);
nand U16457 (N_16457,N_16388,N_16226);
or U16458 (N_16458,N_16248,N_16375);
or U16459 (N_16459,N_16223,N_16269);
xor U16460 (N_16460,N_16314,N_16331);
and U16461 (N_16461,N_16263,N_16322);
xor U16462 (N_16462,N_16353,N_16383);
xor U16463 (N_16463,N_16268,N_16293);
nor U16464 (N_16464,N_16287,N_16305);
or U16465 (N_16465,N_16362,N_16258);
nor U16466 (N_16466,N_16391,N_16295);
nor U16467 (N_16467,N_16227,N_16292);
nand U16468 (N_16468,N_16302,N_16387);
nand U16469 (N_16469,N_16338,N_16297);
xnor U16470 (N_16470,N_16363,N_16276);
and U16471 (N_16471,N_16384,N_16348);
nor U16472 (N_16472,N_16345,N_16396);
or U16473 (N_16473,N_16399,N_16381);
nand U16474 (N_16474,N_16341,N_16374);
and U16475 (N_16475,N_16256,N_16308);
and U16476 (N_16476,N_16390,N_16289);
and U16477 (N_16477,N_16214,N_16282);
and U16478 (N_16478,N_16340,N_16358);
nand U16479 (N_16479,N_16240,N_16355);
and U16480 (N_16480,N_16259,N_16204);
nor U16481 (N_16481,N_16274,N_16209);
or U16482 (N_16482,N_16330,N_16309);
xnor U16483 (N_16483,N_16224,N_16278);
and U16484 (N_16484,N_16398,N_16392);
and U16485 (N_16485,N_16229,N_16313);
xnor U16486 (N_16486,N_16280,N_16366);
nand U16487 (N_16487,N_16273,N_16228);
and U16488 (N_16488,N_16376,N_16265);
nand U16489 (N_16489,N_16260,N_16316);
and U16490 (N_16490,N_16271,N_16382);
or U16491 (N_16491,N_16206,N_16221);
and U16492 (N_16492,N_16318,N_16321);
and U16493 (N_16493,N_16250,N_16236);
nor U16494 (N_16494,N_16349,N_16303);
and U16495 (N_16495,N_16242,N_16222);
or U16496 (N_16496,N_16395,N_16344);
or U16497 (N_16497,N_16254,N_16352);
xnor U16498 (N_16498,N_16205,N_16319);
or U16499 (N_16499,N_16241,N_16284);
or U16500 (N_16500,N_16355,N_16353);
and U16501 (N_16501,N_16347,N_16321);
nor U16502 (N_16502,N_16310,N_16327);
or U16503 (N_16503,N_16329,N_16352);
and U16504 (N_16504,N_16201,N_16380);
xor U16505 (N_16505,N_16382,N_16230);
nor U16506 (N_16506,N_16264,N_16361);
and U16507 (N_16507,N_16352,N_16279);
nor U16508 (N_16508,N_16231,N_16393);
nand U16509 (N_16509,N_16356,N_16364);
and U16510 (N_16510,N_16293,N_16309);
xor U16511 (N_16511,N_16258,N_16388);
nor U16512 (N_16512,N_16291,N_16278);
nand U16513 (N_16513,N_16375,N_16251);
and U16514 (N_16514,N_16224,N_16225);
nor U16515 (N_16515,N_16237,N_16244);
nand U16516 (N_16516,N_16372,N_16251);
xnor U16517 (N_16517,N_16327,N_16302);
xor U16518 (N_16518,N_16381,N_16337);
and U16519 (N_16519,N_16276,N_16370);
nand U16520 (N_16520,N_16320,N_16396);
xor U16521 (N_16521,N_16349,N_16213);
nand U16522 (N_16522,N_16382,N_16217);
or U16523 (N_16523,N_16329,N_16213);
nor U16524 (N_16524,N_16252,N_16383);
or U16525 (N_16525,N_16276,N_16395);
nor U16526 (N_16526,N_16260,N_16393);
nand U16527 (N_16527,N_16358,N_16276);
and U16528 (N_16528,N_16307,N_16288);
xor U16529 (N_16529,N_16303,N_16299);
xnor U16530 (N_16530,N_16380,N_16207);
or U16531 (N_16531,N_16374,N_16222);
nand U16532 (N_16532,N_16346,N_16355);
or U16533 (N_16533,N_16382,N_16250);
xor U16534 (N_16534,N_16239,N_16319);
or U16535 (N_16535,N_16286,N_16310);
nand U16536 (N_16536,N_16217,N_16328);
and U16537 (N_16537,N_16316,N_16317);
or U16538 (N_16538,N_16376,N_16200);
nor U16539 (N_16539,N_16313,N_16365);
and U16540 (N_16540,N_16356,N_16320);
nor U16541 (N_16541,N_16225,N_16232);
nand U16542 (N_16542,N_16325,N_16295);
or U16543 (N_16543,N_16341,N_16267);
nand U16544 (N_16544,N_16205,N_16286);
nand U16545 (N_16545,N_16343,N_16210);
xnor U16546 (N_16546,N_16252,N_16319);
and U16547 (N_16547,N_16239,N_16353);
or U16548 (N_16548,N_16234,N_16314);
xor U16549 (N_16549,N_16363,N_16251);
or U16550 (N_16550,N_16214,N_16213);
xnor U16551 (N_16551,N_16366,N_16278);
nor U16552 (N_16552,N_16373,N_16353);
and U16553 (N_16553,N_16228,N_16374);
or U16554 (N_16554,N_16338,N_16267);
nor U16555 (N_16555,N_16259,N_16364);
nor U16556 (N_16556,N_16207,N_16381);
xnor U16557 (N_16557,N_16241,N_16301);
xor U16558 (N_16558,N_16337,N_16346);
xor U16559 (N_16559,N_16222,N_16323);
nand U16560 (N_16560,N_16331,N_16267);
xnor U16561 (N_16561,N_16381,N_16349);
and U16562 (N_16562,N_16210,N_16392);
and U16563 (N_16563,N_16353,N_16305);
and U16564 (N_16564,N_16272,N_16238);
nor U16565 (N_16565,N_16381,N_16354);
and U16566 (N_16566,N_16222,N_16232);
or U16567 (N_16567,N_16285,N_16312);
nor U16568 (N_16568,N_16377,N_16212);
and U16569 (N_16569,N_16375,N_16274);
and U16570 (N_16570,N_16354,N_16378);
xor U16571 (N_16571,N_16277,N_16222);
and U16572 (N_16572,N_16363,N_16285);
nor U16573 (N_16573,N_16365,N_16390);
nand U16574 (N_16574,N_16365,N_16389);
nor U16575 (N_16575,N_16394,N_16273);
and U16576 (N_16576,N_16271,N_16323);
xor U16577 (N_16577,N_16201,N_16311);
nor U16578 (N_16578,N_16355,N_16361);
xnor U16579 (N_16579,N_16272,N_16337);
xor U16580 (N_16580,N_16207,N_16337);
or U16581 (N_16581,N_16263,N_16259);
or U16582 (N_16582,N_16313,N_16265);
nor U16583 (N_16583,N_16215,N_16276);
nor U16584 (N_16584,N_16318,N_16242);
xor U16585 (N_16585,N_16332,N_16221);
nand U16586 (N_16586,N_16303,N_16363);
and U16587 (N_16587,N_16215,N_16356);
or U16588 (N_16588,N_16246,N_16202);
or U16589 (N_16589,N_16292,N_16247);
or U16590 (N_16590,N_16274,N_16300);
nor U16591 (N_16591,N_16241,N_16242);
or U16592 (N_16592,N_16398,N_16295);
nor U16593 (N_16593,N_16270,N_16348);
nor U16594 (N_16594,N_16290,N_16296);
nor U16595 (N_16595,N_16336,N_16368);
or U16596 (N_16596,N_16243,N_16260);
xor U16597 (N_16597,N_16349,N_16335);
and U16598 (N_16598,N_16344,N_16367);
and U16599 (N_16599,N_16367,N_16322);
nand U16600 (N_16600,N_16472,N_16417);
or U16601 (N_16601,N_16520,N_16431);
nor U16602 (N_16602,N_16465,N_16597);
xnor U16603 (N_16603,N_16411,N_16462);
xnor U16604 (N_16604,N_16437,N_16412);
nand U16605 (N_16605,N_16568,N_16413);
nor U16606 (N_16606,N_16428,N_16476);
xor U16607 (N_16607,N_16557,N_16502);
and U16608 (N_16608,N_16584,N_16471);
xor U16609 (N_16609,N_16489,N_16575);
or U16610 (N_16610,N_16421,N_16510);
and U16611 (N_16611,N_16400,N_16565);
xor U16612 (N_16612,N_16403,N_16481);
or U16613 (N_16613,N_16509,N_16461);
or U16614 (N_16614,N_16493,N_16596);
nand U16615 (N_16615,N_16422,N_16537);
nor U16616 (N_16616,N_16562,N_16579);
nor U16617 (N_16617,N_16441,N_16416);
nand U16618 (N_16618,N_16521,N_16410);
nor U16619 (N_16619,N_16547,N_16420);
and U16620 (N_16620,N_16540,N_16552);
and U16621 (N_16621,N_16452,N_16598);
xor U16622 (N_16622,N_16508,N_16494);
nor U16623 (N_16623,N_16429,N_16451);
xnor U16624 (N_16624,N_16513,N_16427);
and U16625 (N_16625,N_16514,N_16570);
and U16626 (N_16626,N_16546,N_16402);
or U16627 (N_16627,N_16517,N_16566);
or U16628 (N_16628,N_16443,N_16561);
nand U16629 (N_16629,N_16445,N_16444);
xnor U16630 (N_16630,N_16544,N_16446);
and U16631 (N_16631,N_16539,N_16555);
or U16632 (N_16632,N_16496,N_16483);
nand U16633 (N_16633,N_16586,N_16577);
nand U16634 (N_16634,N_16573,N_16543);
or U16635 (N_16635,N_16458,N_16529);
or U16636 (N_16636,N_16487,N_16564);
xnor U16637 (N_16637,N_16470,N_16409);
nand U16638 (N_16638,N_16426,N_16559);
nor U16639 (N_16639,N_16455,N_16459);
xnor U16640 (N_16640,N_16556,N_16599);
or U16641 (N_16641,N_16475,N_16524);
or U16642 (N_16642,N_16518,N_16504);
nor U16643 (N_16643,N_16419,N_16450);
or U16644 (N_16644,N_16490,N_16534);
and U16645 (N_16645,N_16477,N_16523);
nand U16646 (N_16646,N_16589,N_16506);
xor U16647 (N_16647,N_16585,N_16560);
xor U16648 (N_16648,N_16482,N_16460);
nor U16649 (N_16649,N_16525,N_16554);
or U16650 (N_16650,N_16594,N_16473);
and U16651 (N_16651,N_16418,N_16480);
nand U16652 (N_16652,N_16574,N_16478);
xnor U16653 (N_16653,N_16583,N_16425);
and U16654 (N_16654,N_16528,N_16563);
nor U16655 (N_16655,N_16515,N_16414);
xnor U16656 (N_16656,N_16438,N_16501);
nand U16657 (N_16657,N_16590,N_16538);
xnor U16658 (N_16658,N_16466,N_16591);
xnor U16659 (N_16659,N_16434,N_16580);
nand U16660 (N_16660,N_16595,N_16469);
nand U16661 (N_16661,N_16497,N_16440);
nor U16662 (N_16662,N_16516,N_16484);
and U16663 (N_16663,N_16454,N_16522);
xnor U16664 (N_16664,N_16535,N_16433);
xor U16665 (N_16665,N_16581,N_16542);
and U16666 (N_16666,N_16404,N_16532);
nand U16667 (N_16667,N_16408,N_16582);
and U16668 (N_16668,N_16526,N_16572);
nand U16669 (N_16669,N_16519,N_16512);
and U16670 (N_16670,N_16491,N_16549);
nor U16671 (N_16671,N_16474,N_16553);
nand U16672 (N_16672,N_16578,N_16463);
nand U16673 (N_16673,N_16531,N_16533);
xnor U16674 (N_16674,N_16423,N_16449);
xnor U16675 (N_16675,N_16569,N_16503);
or U16676 (N_16676,N_16406,N_16576);
nand U16677 (N_16677,N_16498,N_16405);
xnor U16678 (N_16678,N_16550,N_16424);
or U16679 (N_16679,N_16486,N_16432);
nor U16680 (N_16680,N_16430,N_16464);
or U16681 (N_16681,N_16505,N_16468);
nand U16682 (N_16682,N_16567,N_16407);
xnor U16683 (N_16683,N_16587,N_16447);
nor U16684 (N_16684,N_16401,N_16495);
nand U16685 (N_16685,N_16541,N_16593);
nand U16686 (N_16686,N_16571,N_16492);
nor U16687 (N_16687,N_16551,N_16527);
xnor U16688 (N_16688,N_16415,N_16435);
and U16689 (N_16689,N_16488,N_16439);
nor U16690 (N_16690,N_16545,N_16485);
nand U16691 (N_16691,N_16588,N_16530);
and U16692 (N_16692,N_16456,N_16467);
nand U16693 (N_16693,N_16511,N_16499);
or U16694 (N_16694,N_16558,N_16500);
xnor U16695 (N_16695,N_16436,N_16507);
xnor U16696 (N_16696,N_16448,N_16592);
nand U16697 (N_16697,N_16536,N_16457);
nor U16698 (N_16698,N_16453,N_16548);
or U16699 (N_16699,N_16479,N_16442);
xor U16700 (N_16700,N_16596,N_16417);
nor U16701 (N_16701,N_16551,N_16538);
or U16702 (N_16702,N_16438,N_16433);
nand U16703 (N_16703,N_16447,N_16586);
nand U16704 (N_16704,N_16425,N_16453);
xor U16705 (N_16705,N_16406,N_16423);
and U16706 (N_16706,N_16542,N_16543);
nand U16707 (N_16707,N_16493,N_16542);
or U16708 (N_16708,N_16428,N_16400);
and U16709 (N_16709,N_16523,N_16557);
and U16710 (N_16710,N_16529,N_16558);
nor U16711 (N_16711,N_16541,N_16474);
nand U16712 (N_16712,N_16402,N_16528);
nor U16713 (N_16713,N_16534,N_16510);
or U16714 (N_16714,N_16530,N_16454);
xnor U16715 (N_16715,N_16459,N_16500);
xor U16716 (N_16716,N_16484,N_16417);
xnor U16717 (N_16717,N_16565,N_16425);
and U16718 (N_16718,N_16490,N_16599);
and U16719 (N_16719,N_16469,N_16541);
or U16720 (N_16720,N_16432,N_16417);
nor U16721 (N_16721,N_16489,N_16465);
and U16722 (N_16722,N_16558,N_16453);
nor U16723 (N_16723,N_16417,N_16446);
nor U16724 (N_16724,N_16452,N_16546);
and U16725 (N_16725,N_16531,N_16470);
and U16726 (N_16726,N_16411,N_16484);
or U16727 (N_16727,N_16599,N_16568);
or U16728 (N_16728,N_16540,N_16557);
xor U16729 (N_16729,N_16488,N_16473);
xor U16730 (N_16730,N_16424,N_16590);
nand U16731 (N_16731,N_16437,N_16462);
xnor U16732 (N_16732,N_16513,N_16525);
or U16733 (N_16733,N_16587,N_16520);
nor U16734 (N_16734,N_16482,N_16551);
and U16735 (N_16735,N_16575,N_16561);
nand U16736 (N_16736,N_16524,N_16421);
nor U16737 (N_16737,N_16517,N_16568);
nand U16738 (N_16738,N_16419,N_16455);
xor U16739 (N_16739,N_16435,N_16597);
and U16740 (N_16740,N_16567,N_16432);
nor U16741 (N_16741,N_16451,N_16427);
xnor U16742 (N_16742,N_16411,N_16425);
xor U16743 (N_16743,N_16473,N_16585);
or U16744 (N_16744,N_16460,N_16595);
nand U16745 (N_16745,N_16522,N_16505);
and U16746 (N_16746,N_16522,N_16418);
nand U16747 (N_16747,N_16407,N_16459);
or U16748 (N_16748,N_16462,N_16503);
and U16749 (N_16749,N_16581,N_16551);
and U16750 (N_16750,N_16485,N_16471);
nand U16751 (N_16751,N_16446,N_16452);
xnor U16752 (N_16752,N_16463,N_16441);
or U16753 (N_16753,N_16423,N_16442);
nand U16754 (N_16754,N_16475,N_16503);
nor U16755 (N_16755,N_16485,N_16443);
or U16756 (N_16756,N_16550,N_16454);
and U16757 (N_16757,N_16406,N_16415);
nand U16758 (N_16758,N_16454,N_16457);
nand U16759 (N_16759,N_16478,N_16584);
nor U16760 (N_16760,N_16552,N_16476);
and U16761 (N_16761,N_16474,N_16492);
and U16762 (N_16762,N_16532,N_16520);
nor U16763 (N_16763,N_16467,N_16495);
nor U16764 (N_16764,N_16525,N_16465);
nor U16765 (N_16765,N_16539,N_16547);
or U16766 (N_16766,N_16452,N_16442);
nor U16767 (N_16767,N_16533,N_16554);
nor U16768 (N_16768,N_16586,N_16544);
xnor U16769 (N_16769,N_16566,N_16573);
or U16770 (N_16770,N_16460,N_16409);
nor U16771 (N_16771,N_16569,N_16530);
nand U16772 (N_16772,N_16581,N_16582);
nand U16773 (N_16773,N_16449,N_16493);
nand U16774 (N_16774,N_16418,N_16417);
xnor U16775 (N_16775,N_16565,N_16442);
xnor U16776 (N_16776,N_16597,N_16575);
or U16777 (N_16777,N_16402,N_16460);
and U16778 (N_16778,N_16536,N_16515);
xor U16779 (N_16779,N_16537,N_16458);
or U16780 (N_16780,N_16590,N_16443);
or U16781 (N_16781,N_16499,N_16402);
and U16782 (N_16782,N_16433,N_16475);
or U16783 (N_16783,N_16582,N_16552);
nor U16784 (N_16784,N_16585,N_16574);
nand U16785 (N_16785,N_16409,N_16407);
nor U16786 (N_16786,N_16592,N_16450);
xnor U16787 (N_16787,N_16599,N_16507);
xnor U16788 (N_16788,N_16580,N_16507);
or U16789 (N_16789,N_16437,N_16529);
and U16790 (N_16790,N_16420,N_16474);
and U16791 (N_16791,N_16473,N_16411);
nand U16792 (N_16792,N_16454,N_16567);
or U16793 (N_16793,N_16515,N_16430);
or U16794 (N_16794,N_16450,N_16577);
and U16795 (N_16795,N_16488,N_16544);
and U16796 (N_16796,N_16543,N_16521);
nand U16797 (N_16797,N_16562,N_16590);
or U16798 (N_16798,N_16522,N_16514);
xnor U16799 (N_16799,N_16441,N_16569);
xnor U16800 (N_16800,N_16766,N_16743);
nand U16801 (N_16801,N_16651,N_16746);
and U16802 (N_16802,N_16715,N_16693);
or U16803 (N_16803,N_16750,N_16729);
and U16804 (N_16804,N_16642,N_16763);
nand U16805 (N_16805,N_16633,N_16726);
xor U16806 (N_16806,N_16640,N_16770);
and U16807 (N_16807,N_16728,N_16778);
or U16808 (N_16808,N_16739,N_16676);
xor U16809 (N_16809,N_16732,N_16742);
nand U16810 (N_16810,N_16677,N_16667);
xnor U16811 (N_16811,N_16737,N_16777);
and U16812 (N_16812,N_16784,N_16669);
nand U16813 (N_16813,N_16782,N_16736);
and U16814 (N_16814,N_16789,N_16656);
or U16815 (N_16815,N_16691,N_16794);
and U16816 (N_16816,N_16688,N_16659);
nand U16817 (N_16817,N_16622,N_16675);
or U16818 (N_16818,N_16653,N_16685);
nand U16819 (N_16819,N_16634,N_16648);
or U16820 (N_16820,N_16627,N_16623);
nand U16821 (N_16821,N_16722,N_16745);
nor U16822 (N_16822,N_16717,N_16628);
or U16823 (N_16823,N_16658,N_16703);
nand U16824 (N_16824,N_16684,N_16681);
xor U16825 (N_16825,N_16682,N_16613);
nand U16826 (N_16826,N_16604,N_16711);
or U16827 (N_16827,N_16609,N_16748);
nand U16828 (N_16828,N_16665,N_16654);
xor U16829 (N_16829,N_16649,N_16647);
nor U16830 (N_16830,N_16643,N_16673);
nand U16831 (N_16831,N_16702,N_16731);
or U16832 (N_16832,N_16662,N_16701);
nor U16833 (N_16833,N_16707,N_16605);
and U16834 (N_16834,N_16683,N_16758);
nand U16835 (N_16835,N_16601,N_16674);
nand U16836 (N_16836,N_16757,N_16626);
or U16837 (N_16837,N_16760,N_16754);
or U16838 (N_16838,N_16720,N_16775);
xnor U16839 (N_16839,N_16617,N_16695);
nor U16840 (N_16840,N_16637,N_16621);
or U16841 (N_16841,N_16773,N_16641);
and U16842 (N_16842,N_16759,N_16706);
or U16843 (N_16843,N_16797,N_16644);
nor U16844 (N_16844,N_16713,N_16664);
nor U16845 (N_16845,N_16655,N_16719);
and U16846 (N_16846,N_16636,N_16671);
nand U16847 (N_16847,N_16632,N_16646);
xor U16848 (N_16848,N_16793,N_16630);
xor U16849 (N_16849,N_16710,N_16749);
nor U16850 (N_16850,N_16735,N_16716);
nor U16851 (N_16851,N_16768,N_16699);
and U16852 (N_16852,N_16698,N_16666);
or U16853 (N_16853,N_16756,N_16786);
xor U16854 (N_16854,N_16704,N_16725);
and U16855 (N_16855,N_16602,N_16718);
or U16856 (N_16856,N_16614,N_16697);
xor U16857 (N_16857,N_16796,N_16600);
xnor U16858 (N_16858,N_16690,N_16752);
or U16859 (N_16859,N_16753,N_16687);
xor U16860 (N_16860,N_16791,N_16638);
and U16861 (N_16861,N_16694,N_16783);
nand U16862 (N_16862,N_16755,N_16708);
nand U16863 (N_16863,N_16700,N_16714);
nand U16864 (N_16864,N_16639,N_16615);
xnor U16865 (N_16865,N_16727,N_16792);
nand U16866 (N_16866,N_16663,N_16764);
nand U16867 (N_16867,N_16787,N_16771);
and U16868 (N_16868,N_16661,N_16776);
or U16869 (N_16869,N_16680,N_16744);
and U16870 (N_16870,N_16747,N_16774);
xor U16871 (N_16871,N_16686,N_16650);
nor U16872 (N_16872,N_16618,N_16689);
and U16873 (N_16873,N_16781,N_16733);
xnor U16874 (N_16874,N_16741,N_16761);
nand U16875 (N_16875,N_16705,N_16620);
xnor U16876 (N_16876,N_16606,N_16611);
nand U16877 (N_16877,N_16678,N_16734);
xor U16878 (N_16878,N_16635,N_16712);
nand U16879 (N_16879,N_16723,N_16660);
and U16880 (N_16880,N_16779,N_16692);
nand U16881 (N_16881,N_16619,N_16645);
and U16882 (N_16882,N_16785,N_16629);
xor U16883 (N_16883,N_16709,N_16788);
and U16884 (N_16884,N_16612,N_16624);
xnor U16885 (N_16885,N_16625,N_16610);
xnor U16886 (N_16886,N_16751,N_16631);
xor U16887 (N_16887,N_16721,N_16608);
and U16888 (N_16888,N_16652,N_16762);
and U16889 (N_16889,N_16730,N_16780);
and U16890 (N_16890,N_16679,N_16724);
or U16891 (N_16891,N_16769,N_16798);
and U16892 (N_16892,N_16790,N_16607);
xor U16893 (N_16893,N_16696,N_16670);
nor U16894 (N_16894,N_16672,N_16668);
or U16895 (N_16895,N_16616,N_16657);
nand U16896 (N_16896,N_16738,N_16772);
nand U16897 (N_16897,N_16767,N_16765);
nor U16898 (N_16898,N_16740,N_16799);
xor U16899 (N_16899,N_16603,N_16795);
and U16900 (N_16900,N_16753,N_16745);
or U16901 (N_16901,N_16627,N_16608);
and U16902 (N_16902,N_16657,N_16650);
nand U16903 (N_16903,N_16728,N_16612);
xor U16904 (N_16904,N_16603,N_16729);
xnor U16905 (N_16905,N_16727,N_16746);
or U16906 (N_16906,N_16789,N_16749);
or U16907 (N_16907,N_16705,N_16711);
nor U16908 (N_16908,N_16712,N_16769);
or U16909 (N_16909,N_16761,N_16726);
xnor U16910 (N_16910,N_16662,N_16668);
nand U16911 (N_16911,N_16707,N_16781);
nand U16912 (N_16912,N_16791,N_16751);
xnor U16913 (N_16913,N_16729,N_16679);
or U16914 (N_16914,N_16645,N_16606);
nor U16915 (N_16915,N_16759,N_16765);
and U16916 (N_16916,N_16794,N_16640);
nand U16917 (N_16917,N_16731,N_16633);
nor U16918 (N_16918,N_16684,N_16793);
xor U16919 (N_16919,N_16603,N_16736);
nor U16920 (N_16920,N_16686,N_16776);
nor U16921 (N_16921,N_16780,N_16604);
and U16922 (N_16922,N_16677,N_16653);
nand U16923 (N_16923,N_16795,N_16641);
nand U16924 (N_16924,N_16783,N_16665);
and U16925 (N_16925,N_16761,N_16615);
xor U16926 (N_16926,N_16735,N_16701);
xor U16927 (N_16927,N_16762,N_16761);
or U16928 (N_16928,N_16787,N_16608);
xor U16929 (N_16929,N_16677,N_16621);
nor U16930 (N_16930,N_16620,N_16707);
nand U16931 (N_16931,N_16724,N_16699);
xor U16932 (N_16932,N_16705,N_16645);
and U16933 (N_16933,N_16658,N_16648);
or U16934 (N_16934,N_16652,N_16749);
or U16935 (N_16935,N_16681,N_16635);
nand U16936 (N_16936,N_16606,N_16790);
xor U16937 (N_16937,N_16759,N_16699);
nand U16938 (N_16938,N_16745,N_16613);
or U16939 (N_16939,N_16665,N_16608);
and U16940 (N_16940,N_16719,N_16796);
or U16941 (N_16941,N_16699,N_16695);
nor U16942 (N_16942,N_16610,N_16632);
nand U16943 (N_16943,N_16616,N_16600);
or U16944 (N_16944,N_16636,N_16601);
or U16945 (N_16945,N_16787,N_16798);
and U16946 (N_16946,N_16694,N_16607);
nand U16947 (N_16947,N_16633,N_16681);
or U16948 (N_16948,N_16764,N_16610);
and U16949 (N_16949,N_16702,N_16698);
or U16950 (N_16950,N_16732,N_16674);
nor U16951 (N_16951,N_16777,N_16611);
xor U16952 (N_16952,N_16683,N_16752);
or U16953 (N_16953,N_16728,N_16624);
xor U16954 (N_16954,N_16737,N_16740);
or U16955 (N_16955,N_16736,N_16670);
nand U16956 (N_16956,N_16676,N_16664);
or U16957 (N_16957,N_16796,N_16697);
nand U16958 (N_16958,N_16760,N_16756);
xor U16959 (N_16959,N_16707,N_16629);
nor U16960 (N_16960,N_16680,N_16630);
nand U16961 (N_16961,N_16752,N_16614);
or U16962 (N_16962,N_16798,N_16718);
xor U16963 (N_16963,N_16772,N_16627);
nor U16964 (N_16964,N_16612,N_16793);
or U16965 (N_16965,N_16610,N_16645);
or U16966 (N_16966,N_16625,N_16710);
and U16967 (N_16967,N_16620,N_16656);
xnor U16968 (N_16968,N_16649,N_16756);
nor U16969 (N_16969,N_16622,N_16705);
xor U16970 (N_16970,N_16745,N_16751);
nand U16971 (N_16971,N_16659,N_16719);
and U16972 (N_16972,N_16761,N_16788);
or U16973 (N_16973,N_16737,N_16682);
and U16974 (N_16974,N_16764,N_16798);
and U16975 (N_16975,N_16772,N_16636);
nand U16976 (N_16976,N_16765,N_16738);
xnor U16977 (N_16977,N_16667,N_16641);
and U16978 (N_16978,N_16732,N_16632);
nor U16979 (N_16979,N_16784,N_16791);
and U16980 (N_16980,N_16611,N_16614);
nor U16981 (N_16981,N_16795,N_16772);
or U16982 (N_16982,N_16623,N_16700);
nand U16983 (N_16983,N_16716,N_16607);
or U16984 (N_16984,N_16678,N_16640);
or U16985 (N_16985,N_16694,N_16635);
nand U16986 (N_16986,N_16793,N_16663);
xor U16987 (N_16987,N_16676,N_16682);
nor U16988 (N_16988,N_16677,N_16616);
nor U16989 (N_16989,N_16602,N_16758);
nand U16990 (N_16990,N_16742,N_16711);
xnor U16991 (N_16991,N_16736,N_16731);
nand U16992 (N_16992,N_16649,N_16682);
nor U16993 (N_16993,N_16783,N_16688);
and U16994 (N_16994,N_16684,N_16633);
or U16995 (N_16995,N_16609,N_16649);
nand U16996 (N_16996,N_16693,N_16616);
xnor U16997 (N_16997,N_16700,N_16672);
nand U16998 (N_16998,N_16640,N_16611);
or U16999 (N_16999,N_16642,N_16760);
or U17000 (N_17000,N_16857,N_16866);
xnor U17001 (N_17001,N_16948,N_16932);
nand U17002 (N_17002,N_16911,N_16899);
and U17003 (N_17003,N_16918,N_16954);
nand U17004 (N_17004,N_16843,N_16930);
xor U17005 (N_17005,N_16811,N_16879);
xor U17006 (N_17006,N_16847,N_16939);
and U17007 (N_17007,N_16810,N_16975);
xnor U17008 (N_17008,N_16838,N_16873);
xnor U17009 (N_17009,N_16963,N_16987);
nand U17010 (N_17010,N_16988,N_16924);
xnor U17011 (N_17011,N_16931,N_16890);
nor U17012 (N_17012,N_16898,N_16950);
nand U17013 (N_17013,N_16983,N_16974);
xor U17014 (N_17014,N_16962,N_16804);
nor U17015 (N_17015,N_16929,N_16822);
or U17016 (N_17016,N_16845,N_16894);
and U17017 (N_17017,N_16969,N_16826);
nor U17018 (N_17018,N_16961,N_16882);
xor U17019 (N_17019,N_16947,N_16900);
xnor U17020 (N_17020,N_16957,N_16968);
nor U17021 (N_17021,N_16992,N_16925);
and U17022 (N_17022,N_16986,N_16909);
nor U17023 (N_17023,N_16885,N_16807);
nand U17024 (N_17024,N_16858,N_16896);
or U17025 (N_17025,N_16995,N_16808);
and U17026 (N_17026,N_16914,N_16904);
and U17027 (N_17027,N_16891,N_16846);
nor U17028 (N_17028,N_16883,N_16952);
and U17029 (N_17029,N_16941,N_16852);
nand U17030 (N_17030,N_16981,N_16820);
xor U17031 (N_17031,N_16874,N_16990);
nand U17032 (N_17032,N_16831,N_16823);
nor U17033 (N_17033,N_16921,N_16869);
and U17034 (N_17034,N_16870,N_16850);
and U17035 (N_17035,N_16901,N_16915);
nand U17036 (N_17036,N_16926,N_16958);
and U17037 (N_17037,N_16828,N_16818);
xor U17038 (N_17038,N_16844,N_16906);
and U17039 (N_17039,N_16993,N_16825);
and U17040 (N_17040,N_16877,N_16977);
xor U17041 (N_17041,N_16938,N_16856);
xor U17042 (N_17042,N_16907,N_16934);
and U17043 (N_17043,N_16878,N_16966);
nand U17044 (N_17044,N_16884,N_16935);
nand U17045 (N_17045,N_16861,N_16839);
nor U17046 (N_17046,N_16859,N_16860);
nor U17047 (N_17047,N_16864,N_16815);
and U17048 (N_17048,N_16871,N_16985);
and U17049 (N_17049,N_16835,N_16976);
nor U17050 (N_17050,N_16994,N_16979);
nor U17051 (N_17051,N_16999,N_16972);
nand U17052 (N_17052,N_16951,N_16821);
xnor U17053 (N_17053,N_16991,N_16830);
nand U17054 (N_17054,N_16980,N_16943);
nand U17055 (N_17055,N_16881,N_16893);
or U17056 (N_17056,N_16997,N_16889);
nand U17057 (N_17057,N_16888,N_16827);
nor U17058 (N_17058,N_16989,N_16910);
xnor U17059 (N_17059,N_16875,N_16868);
nand U17060 (N_17060,N_16848,N_16892);
nor U17061 (N_17061,N_16801,N_16937);
or U17062 (N_17062,N_16876,N_16933);
and U17063 (N_17063,N_16834,N_16944);
and U17064 (N_17064,N_16945,N_16862);
or U17065 (N_17065,N_16905,N_16813);
or U17066 (N_17066,N_16978,N_16984);
and U17067 (N_17067,N_16959,N_16922);
or U17068 (N_17068,N_16956,N_16895);
or U17069 (N_17069,N_16982,N_16946);
and U17070 (N_17070,N_16927,N_16902);
xor U17071 (N_17071,N_16824,N_16840);
or U17072 (N_17072,N_16996,N_16837);
xnor U17073 (N_17073,N_16940,N_16903);
or U17074 (N_17074,N_16923,N_16819);
nand U17075 (N_17075,N_16809,N_16872);
xor U17076 (N_17076,N_16998,N_16897);
nor U17077 (N_17077,N_16865,N_16964);
or U17078 (N_17078,N_16863,N_16971);
nand U17079 (N_17079,N_16805,N_16967);
and U17080 (N_17080,N_16836,N_16854);
nand U17081 (N_17081,N_16829,N_16851);
xnor U17082 (N_17082,N_16880,N_16806);
nand U17083 (N_17083,N_16965,N_16853);
and U17084 (N_17084,N_16800,N_16936);
xnor U17085 (N_17085,N_16833,N_16919);
xnor U17086 (N_17086,N_16842,N_16841);
xnor U17087 (N_17087,N_16812,N_16814);
nand U17088 (N_17088,N_16802,N_16886);
xnor U17089 (N_17089,N_16849,N_16920);
nor U17090 (N_17090,N_16928,N_16960);
xnor U17091 (N_17091,N_16942,N_16803);
nand U17092 (N_17092,N_16949,N_16867);
nand U17093 (N_17093,N_16816,N_16887);
nand U17094 (N_17094,N_16953,N_16955);
nor U17095 (N_17095,N_16973,N_16855);
and U17096 (N_17096,N_16970,N_16817);
nor U17097 (N_17097,N_16912,N_16832);
and U17098 (N_17098,N_16913,N_16908);
xor U17099 (N_17099,N_16916,N_16917);
or U17100 (N_17100,N_16913,N_16927);
nor U17101 (N_17101,N_16831,N_16934);
nand U17102 (N_17102,N_16991,N_16821);
nand U17103 (N_17103,N_16913,N_16930);
xnor U17104 (N_17104,N_16866,N_16842);
nand U17105 (N_17105,N_16948,N_16858);
nor U17106 (N_17106,N_16933,N_16884);
nor U17107 (N_17107,N_16863,N_16817);
and U17108 (N_17108,N_16908,N_16975);
nand U17109 (N_17109,N_16976,N_16993);
xor U17110 (N_17110,N_16858,N_16876);
or U17111 (N_17111,N_16994,N_16847);
nor U17112 (N_17112,N_16883,N_16866);
and U17113 (N_17113,N_16892,N_16971);
nor U17114 (N_17114,N_16832,N_16834);
xor U17115 (N_17115,N_16986,N_16859);
xnor U17116 (N_17116,N_16917,N_16918);
nor U17117 (N_17117,N_16958,N_16817);
nand U17118 (N_17118,N_16870,N_16959);
and U17119 (N_17119,N_16985,N_16843);
xnor U17120 (N_17120,N_16896,N_16922);
nand U17121 (N_17121,N_16944,N_16818);
nand U17122 (N_17122,N_16842,N_16979);
nand U17123 (N_17123,N_16983,N_16946);
nor U17124 (N_17124,N_16991,N_16870);
or U17125 (N_17125,N_16997,N_16843);
nor U17126 (N_17126,N_16946,N_16810);
xor U17127 (N_17127,N_16871,N_16841);
xnor U17128 (N_17128,N_16854,N_16930);
or U17129 (N_17129,N_16837,N_16882);
xor U17130 (N_17130,N_16886,N_16870);
and U17131 (N_17131,N_16872,N_16804);
and U17132 (N_17132,N_16856,N_16949);
nand U17133 (N_17133,N_16938,N_16993);
and U17134 (N_17134,N_16894,N_16810);
nor U17135 (N_17135,N_16973,N_16847);
nor U17136 (N_17136,N_16960,N_16892);
and U17137 (N_17137,N_16826,N_16802);
nand U17138 (N_17138,N_16936,N_16972);
and U17139 (N_17139,N_16906,N_16992);
nor U17140 (N_17140,N_16966,N_16899);
or U17141 (N_17141,N_16900,N_16985);
nor U17142 (N_17142,N_16926,N_16831);
nor U17143 (N_17143,N_16906,N_16828);
and U17144 (N_17144,N_16839,N_16940);
nand U17145 (N_17145,N_16803,N_16946);
or U17146 (N_17146,N_16984,N_16883);
nand U17147 (N_17147,N_16853,N_16841);
nand U17148 (N_17148,N_16819,N_16910);
or U17149 (N_17149,N_16848,N_16913);
and U17150 (N_17150,N_16900,N_16941);
or U17151 (N_17151,N_16947,N_16963);
and U17152 (N_17152,N_16899,N_16905);
or U17153 (N_17153,N_16860,N_16903);
or U17154 (N_17154,N_16887,N_16938);
nor U17155 (N_17155,N_16886,N_16928);
nor U17156 (N_17156,N_16913,N_16892);
nand U17157 (N_17157,N_16959,N_16899);
nand U17158 (N_17158,N_16851,N_16847);
and U17159 (N_17159,N_16800,N_16910);
nand U17160 (N_17160,N_16854,N_16880);
nor U17161 (N_17161,N_16950,N_16855);
nor U17162 (N_17162,N_16939,N_16835);
and U17163 (N_17163,N_16873,N_16974);
and U17164 (N_17164,N_16905,N_16913);
xnor U17165 (N_17165,N_16976,N_16931);
nor U17166 (N_17166,N_16968,N_16918);
nand U17167 (N_17167,N_16954,N_16912);
xor U17168 (N_17168,N_16896,N_16868);
or U17169 (N_17169,N_16829,N_16824);
nor U17170 (N_17170,N_16970,N_16997);
xnor U17171 (N_17171,N_16818,N_16847);
xor U17172 (N_17172,N_16890,N_16884);
nand U17173 (N_17173,N_16967,N_16828);
nor U17174 (N_17174,N_16916,N_16825);
xnor U17175 (N_17175,N_16921,N_16974);
or U17176 (N_17176,N_16980,N_16937);
nor U17177 (N_17177,N_16991,N_16825);
nor U17178 (N_17178,N_16865,N_16983);
or U17179 (N_17179,N_16819,N_16998);
and U17180 (N_17180,N_16949,N_16850);
nand U17181 (N_17181,N_16904,N_16909);
nor U17182 (N_17182,N_16813,N_16914);
or U17183 (N_17183,N_16870,N_16916);
nor U17184 (N_17184,N_16999,N_16905);
xor U17185 (N_17185,N_16825,N_16814);
and U17186 (N_17186,N_16893,N_16835);
or U17187 (N_17187,N_16866,N_16888);
or U17188 (N_17188,N_16859,N_16983);
and U17189 (N_17189,N_16930,N_16887);
nand U17190 (N_17190,N_16957,N_16807);
xor U17191 (N_17191,N_16980,N_16910);
nand U17192 (N_17192,N_16914,N_16934);
and U17193 (N_17193,N_16883,N_16802);
and U17194 (N_17194,N_16941,N_16998);
nand U17195 (N_17195,N_16965,N_16997);
nor U17196 (N_17196,N_16863,N_16993);
or U17197 (N_17197,N_16942,N_16801);
and U17198 (N_17198,N_16899,N_16808);
or U17199 (N_17199,N_16813,N_16919);
xor U17200 (N_17200,N_17031,N_17166);
or U17201 (N_17201,N_17142,N_17116);
and U17202 (N_17202,N_17147,N_17187);
nor U17203 (N_17203,N_17173,N_17161);
xor U17204 (N_17204,N_17030,N_17089);
nor U17205 (N_17205,N_17131,N_17169);
nor U17206 (N_17206,N_17056,N_17097);
nor U17207 (N_17207,N_17047,N_17082);
nand U17208 (N_17208,N_17025,N_17157);
nand U17209 (N_17209,N_17191,N_17062);
and U17210 (N_17210,N_17046,N_17003);
xor U17211 (N_17211,N_17016,N_17118);
and U17212 (N_17212,N_17154,N_17023);
or U17213 (N_17213,N_17127,N_17069);
xor U17214 (N_17214,N_17102,N_17149);
nand U17215 (N_17215,N_17073,N_17092);
or U17216 (N_17216,N_17034,N_17172);
nor U17217 (N_17217,N_17179,N_17115);
and U17218 (N_17218,N_17086,N_17010);
xnor U17219 (N_17219,N_17117,N_17024);
or U17220 (N_17220,N_17129,N_17111);
and U17221 (N_17221,N_17193,N_17153);
nor U17222 (N_17222,N_17052,N_17167);
xor U17223 (N_17223,N_17171,N_17194);
nor U17224 (N_17224,N_17064,N_17095);
nand U17225 (N_17225,N_17038,N_17192);
xnor U17226 (N_17226,N_17158,N_17007);
nor U17227 (N_17227,N_17144,N_17159);
nor U17228 (N_17228,N_17145,N_17168);
xor U17229 (N_17229,N_17164,N_17195);
or U17230 (N_17230,N_17124,N_17143);
nand U17231 (N_17231,N_17136,N_17040);
and U17232 (N_17232,N_17151,N_17140);
xor U17233 (N_17233,N_17088,N_17074);
and U17234 (N_17234,N_17122,N_17036);
and U17235 (N_17235,N_17049,N_17042);
nor U17236 (N_17236,N_17113,N_17180);
nand U17237 (N_17237,N_17099,N_17170);
and U17238 (N_17238,N_17156,N_17197);
nor U17239 (N_17239,N_17126,N_17104);
nand U17240 (N_17240,N_17001,N_17015);
or U17241 (N_17241,N_17044,N_17027);
xor U17242 (N_17242,N_17132,N_17119);
nor U17243 (N_17243,N_17160,N_17028);
nor U17244 (N_17244,N_17041,N_17125);
xnor U17245 (N_17245,N_17083,N_17189);
nor U17246 (N_17246,N_17130,N_17176);
nand U17247 (N_17247,N_17012,N_17021);
nor U17248 (N_17248,N_17079,N_17045);
nand U17249 (N_17249,N_17076,N_17061);
xnor U17250 (N_17250,N_17181,N_17190);
and U17251 (N_17251,N_17055,N_17066);
nand U17252 (N_17252,N_17043,N_17105);
or U17253 (N_17253,N_17093,N_17121);
nor U17254 (N_17254,N_17196,N_17020);
nand U17255 (N_17255,N_17063,N_17002);
nand U17256 (N_17256,N_17098,N_17058);
nand U17257 (N_17257,N_17078,N_17094);
and U17258 (N_17258,N_17008,N_17146);
nand U17259 (N_17259,N_17152,N_17100);
nor U17260 (N_17260,N_17006,N_17013);
nand U17261 (N_17261,N_17048,N_17184);
or U17262 (N_17262,N_17178,N_17128);
or U17263 (N_17263,N_17199,N_17103);
or U17264 (N_17264,N_17060,N_17134);
and U17265 (N_17265,N_17004,N_17057);
nand U17266 (N_17266,N_17150,N_17174);
xnor U17267 (N_17267,N_17072,N_17009);
nand U17268 (N_17268,N_17050,N_17039);
and U17269 (N_17269,N_17123,N_17087);
or U17270 (N_17270,N_17011,N_17175);
nand U17271 (N_17271,N_17026,N_17109);
nor U17272 (N_17272,N_17120,N_17022);
nand U17273 (N_17273,N_17139,N_17133);
nor U17274 (N_17274,N_17188,N_17018);
nor U17275 (N_17275,N_17141,N_17075);
or U17276 (N_17276,N_17107,N_17077);
or U17277 (N_17277,N_17080,N_17096);
xnor U17278 (N_17278,N_17035,N_17110);
and U17279 (N_17279,N_17198,N_17148);
nand U17280 (N_17280,N_17091,N_17033);
nand U17281 (N_17281,N_17177,N_17070);
and U17282 (N_17282,N_17014,N_17163);
nand U17283 (N_17283,N_17051,N_17183);
xor U17284 (N_17284,N_17138,N_17101);
nand U17285 (N_17285,N_17068,N_17182);
xnor U17286 (N_17286,N_17137,N_17005);
nor U17287 (N_17287,N_17155,N_17032);
or U17288 (N_17288,N_17090,N_17114);
nor U17289 (N_17289,N_17162,N_17017);
nor U17290 (N_17290,N_17165,N_17185);
and U17291 (N_17291,N_17108,N_17054);
and U17292 (N_17292,N_17037,N_17065);
and U17293 (N_17293,N_17106,N_17081);
nor U17294 (N_17294,N_17135,N_17186);
and U17295 (N_17295,N_17085,N_17053);
or U17296 (N_17296,N_17019,N_17112);
or U17297 (N_17297,N_17084,N_17059);
nor U17298 (N_17298,N_17000,N_17029);
and U17299 (N_17299,N_17067,N_17071);
nand U17300 (N_17300,N_17095,N_17130);
nor U17301 (N_17301,N_17089,N_17197);
or U17302 (N_17302,N_17132,N_17172);
or U17303 (N_17303,N_17153,N_17158);
nor U17304 (N_17304,N_17146,N_17131);
nor U17305 (N_17305,N_17120,N_17138);
xnor U17306 (N_17306,N_17044,N_17040);
and U17307 (N_17307,N_17182,N_17188);
xor U17308 (N_17308,N_17181,N_17083);
and U17309 (N_17309,N_17118,N_17116);
nor U17310 (N_17310,N_17089,N_17166);
xnor U17311 (N_17311,N_17139,N_17091);
and U17312 (N_17312,N_17059,N_17064);
nor U17313 (N_17313,N_17013,N_17130);
xor U17314 (N_17314,N_17140,N_17044);
xor U17315 (N_17315,N_17168,N_17118);
or U17316 (N_17316,N_17060,N_17066);
nor U17317 (N_17317,N_17159,N_17181);
nor U17318 (N_17318,N_17046,N_17042);
and U17319 (N_17319,N_17003,N_17001);
or U17320 (N_17320,N_17012,N_17051);
nand U17321 (N_17321,N_17073,N_17126);
or U17322 (N_17322,N_17142,N_17190);
or U17323 (N_17323,N_17029,N_17064);
nor U17324 (N_17324,N_17162,N_17181);
nor U17325 (N_17325,N_17054,N_17080);
nor U17326 (N_17326,N_17194,N_17109);
xnor U17327 (N_17327,N_17073,N_17158);
or U17328 (N_17328,N_17045,N_17023);
or U17329 (N_17329,N_17160,N_17084);
or U17330 (N_17330,N_17163,N_17087);
or U17331 (N_17331,N_17033,N_17076);
nand U17332 (N_17332,N_17063,N_17041);
and U17333 (N_17333,N_17184,N_17031);
xor U17334 (N_17334,N_17126,N_17086);
or U17335 (N_17335,N_17195,N_17166);
and U17336 (N_17336,N_17051,N_17186);
or U17337 (N_17337,N_17005,N_17140);
xor U17338 (N_17338,N_17106,N_17186);
nand U17339 (N_17339,N_17116,N_17150);
nor U17340 (N_17340,N_17195,N_17137);
nor U17341 (N_17341,N_17196,N_17068);
and U17342 (N_17342,N_17057,N_17066);
xor U17343 (N_17343,N_17153,N_17060);
or U17344 (N_17344,N_17193,N_17087);
nand U17345 (N_17345,N_17100,N_17002);
xor U17346 (N_17346,N_17000,N_17177);
or U17347 (N_17347,N_17068,N_17192);
xnor U17348 (N_17348,N_17144,N_17055);
or U17349 (N_17349,N_17145,N_17114);
xor U17350 (N_17350,N_17079,N_17151);
nor U17351 (N_17351,N_17078,N_17110);
or U17352 (N_17352,N_17150,N_17006);
xnor U17353 (N_17353,N_17046,N_17073);
xnor U17354 (N_17354,N_17000,N_17050);
or U17355 (N_17355,N_17038,N_17187);
or U17356 (N_17356,N_17042,N_17141);
or U17357 (N_17357,N_17068,N_17140);
xor U17358 (N_17358,N_17184,N_17035);
nand U17359 (N_17359,N_17003,N_17038);
and U17360 (N_17360,N_17048,N_17025);
or U17361 (N_17361,N_17145,N_17060);
or U17362 (N_17362,N_17059,N_17085);
or U17363 (N_17363,N_17061,N_17085);
or U17364 (N_17364,N_17148,N_17088);
or U17365 (N_17365,N_17022,N_17188);
nand U17366 (N_17366,N_17140,N_17064);
and U17367 (N_17367,N_17011,N_17012);
or U17368 (N_17368,N_17134,N_17022);
nand U17369 (N_17369,N_17171,N_17107);
xnor U17370 (N_17370,N_17093,N_17073);
xor U17371 (N_17371,N_17131,N_17075);
or U17372 (N_17372,N_17109,N_17095);
xor U17373 (N_17373,N_17135,N_17170);
nand U17374 (N_17374,N_17049,N_17029);
or U17375 (N_17375,N_17178,N_17016);
xnor U17376 (N_17376,N_17075,N_17042);
or U17377 (N_17377,N_17013,N_17153);
or U17378 (N_17378,N_17198,N_17108);
nor U17379 (N_17379,N_17022,N_17014);
and U17380 (N_17380,N_17000,N_17165);
nor U17381 (N_17381,N_17135,N_17157);
nand U17382 (N_17382,N_17005,N_17195);
nand U17383 (N_17383,N_17171,N_17031);
or U17384 (N_17384,N_17152,N_17184);
nand U17385 (N_17385,N_17046,N_17092);
or U17386 (N_17386,N_17179,N_17127);
or U17387 (N_17387,N_17062,N_17131);
xnor U17388 (N_17388,N_17163,N_17108);
nand U17389 (N_17389,N_17072,N_17166);
or U17390 (N_17390,N_17078,N_17082);
nand U17391 (N_17391,N_17055,N_17153);
and U17392 (N_17392,N_17040,N_17122);
xnor U17393 (N_17393,N_17123,N_17118);
and U17394 (N_17394,N_17012,N_17149);
or U17395 (N_17395,N_17063,N_17005);
xnor U17396 (N_17396,N_17057,N_17141);
xor U17397 (N_17397,N_17126,N_17039);
nor U17398 (N_17398,N_17141,N_17103);
nor U17399 (N_17399,N_17036,N_17029);
nand U17400 (N_17400,N_17285,N_17306);
nand U17401 (N_17401,N_17391,N_17376);
xnor U17402 (N_17402,N_17219,N_17368);
or U17403 (N_17403,N_17202,N_17214);
nand U17404 (N_17404,N_17209,N_17207);
nor U17405 (N_17405,N_17257,N_17266);
and U17406 (N_17406,N_17387,N_17394);
and U17407 (N_17407,N_17329,N_17226);
xnor U17408 (N_17408,N_17340,N_17256);
nand U17409 (N_17409,N_17277,N_17327);
nand U17410 (N_17410,N_17361,N_17284);
and U17411 (N_17411,N_17262,N_17255);
nor U17412 (N_17412,N_17320,N_17396);
and U17413 (N_17413,N_17310,N_17279);
xnor U17414 (N_17414,N_17352,N_17382);
and U17415 (N_17415,N_17349,N_17213);
nor U17416 (N_17416,N_17205,N_17260);
or U17417 (N_17417,N_17232,N_17305);
nor U17418 (N_17418,N_17316,N_17222);
or U17419 (N_17419,N_17235,N_17204);
and U17420 (N_17420,N_17392,N_17223);
and U17421 (N_17421,N_17244,N_17292);
xor U17422 (N_17422,N_17275,N_17220);
xnor U17423 (N_17423,N_17290,N_17215);
xor U17424 (N_17424,N_17318,N_17337);
nor U17425 (N_17425,N_17228,N_17383);
xor U17426 (N_17426,N_17286,N_17379);
nand U17427 (N_17427,N_17242,N_17324);
nor U17428 (N_17428,N_17388,N_17304);
xnor U17429 (N_17429,N_17236,N_17201);
nor U17430 (N_17430,N_17385,N_17200);
nor U17431 (N_17431,N_17356,N_17339);
and U17432 (N_17432,N_17321,N_17303);
or U17433 (N_17433,N_17347,N_17332);
nand U17434 (N_17434,N_17393,N_17312);
nor U17435 (N_17435,N_17246,N_17291);
nand U17436 (N_17436,N_17359,N_17237);
xor U17437 (N_17437,N_17380,N_17250);
nor U17438 (N_17438,N_17240,N_17363);
xor U17439 (N_17439,N_17398,N_17243);
xor U17440 (N_17440,N_17323,N_17357);
or U17441 (N_17441,N_17289,N_17252);
or U17442 (N_17442,N_17268,N_17390);
nand U17443 (N_17443,N_17206,N_17267);
or U17444 (N_17444,N_17314,N_17384);
nor U17445 (N_17445,N_17366,N_17328);
or U17446 (N_17446,N_17374,N_17338);
nor U17447 (N_17447,N_17360,N_17227);
and U17448 (N_17448,N_17353,N_17258);
xor U17449 (N_17449,N_17253,N_17254);
or U17450 (N_17450,N_17265,N_17355);
nor U17451 (N_17451,N_17269,N_17221);
and U17452 (N_17452,N_17224,N_17386);
nand U17453 (N_17453,N_17333,N_17283);
nand U17454 (N_17454,N_17342,N_17208);
nand U17455 (N_17455,N_17271,N_17238);
and U17456 (N_17456,N_17302,N_17296);
nor U17457 (N_17457,N_17395,N_17365);
nand U17458 (N_17458,N_17293,N_17375);
and U17459 (N_17459,N_17231,N_17278);
xnor U17460 (N_17460,N_17239,N_17325);
or U17461 (N_17461,N_17288,N_17245);
nand U17462 (N_17462,N_17343,N_17354);
nand U17463 (N_17463,N_17210,N_17270);
xnor U17464 (N_17464,N_17287,N_17319);
nor U17465 (N_17465,N_17261,N_17203);
nand U17466 (N_17466,N_17317,N_17341);
nor U17467 (N_17467,N_17218,N_17370);
and U17468 (N_17468,N_17330,N_17350);
or U17469 (N_17469,N_17399,N_17276);
and U17470 (N_17470,N_17348,N_17248);
nor U17471 (N_17471,N_17282,N_17241);
nor U17472 (N_17472,N_17378,N_17273);
xnor U17473 (N_17473,N_17322,N_17281);
and U17474 (N_17474,N_17367,N_17313);
and U17475 (N_17475,N_17225,N_17345);
nor U17476 (N_17476,N_17344,N_17216);
and U17477 (N_17477,N_17247,N_17315);
or U17478 (N_17478,N_17294,N_17295);
or U17479 (N_17479,N_17373,N_17211);
xnor U17480 (N_17480,N_17233,N_17307);
or U17481 (N_17481,N_17336,N_17251);
and U17482 (N_17482,N_17259,N_17263);
or U17483 (N_17483,N_17331,N_17346);
and U17484 (N_17484,N_17229,N_17297);
and U17485 (N_17485,N_17364,N_17274);
nor U17486 (N_17486,N_17377,N_17230);
nor U17487 (N_17487,N_17369,N_17381);
and U17488 (N_17488,N_17389,N_17362);
nor U17489 (N_17489,N_17351,N_17334);
nor U17490 (N_17490,N_17234,N_17272);
or U17491 (N_17491,N_17299,N_17212);
xor U17492 (N_17492,N_17372,N_17397);
xnor U17493 (N_17493,N_17311,N_17308);
or U17494 (N_17494,N_17309,N_17326);
xnor U17495 (N_17495,N_17358,N_17280);
or U17496 (N_17496,N_17249,N_17298);
xor U17497 (N_17497,N_17300,N_17217);
and U17498 (N_17498,N_17301,N_17371);
and U17499 (N_17499,N_17335,N_17264);
or U17500 (N_17500,N_17285,N_17277);
and U17501 (N_17501,N_17284,N_17241);
nand U17502 (N_17502,N_17288,N_17256);
nor U17503 (N_17503,N_17298,N_17358);
and U17504 (N_17504,N_17254,N_17399);
or U17505 (N_17505,N_17212,N_17359);
nor U17506 (N_17506,N_17344,N_17359);
nand U17507 (N_17507,N_17341,N_17326);
nor U17508 (N_17508,N_17283,N_17309);
xor U17509 (N_17509,N_17295,N_17332);
nand U17510 (N_17510,N_17289,N_17269);
nor U17511 (N_17511,N_17204,N_17346);
nand U17512 (N_17512,N_17378,N_17283);
and U17513 (N_17513,N_17225,N_17322);
and U17514 (N_17514,N_17292,N_17219);
and U17515 (N_17515,N_17284,N_17216);
or U17516 (N_17516,N_17277,N_17293);
and U17517 (N_17517,N_17299,N_17209);
nor U17518 (N_17518,N_17254,N_17355);
or U17519 (N_17519,N_17308,N_17316);
or U17520 (N_17520,N_17337,N_17352);
nor U17521 (N_17521,N_17297,N_17290);
nand U17522 (N_17522,N_17367,N_17309);
nor U17523 (N_17523,N_17332,N_17334);
nand U17524 (N_17524,N_17270,N_17347);
and U17525 (N_17525,N_17201,N_17345);
or U17526 (N_17526,N_17204,N_17333);
nand U17527 (N_17527,N_17261,N_17228);
xor U17528 (N_17528,N_17249,N_17390);
xnor U17529 (N_17529,N_17271,N_17324);
or U17530 (N_17530,N_17338,N_17322);
and U17531 (N_17531,N_17325,N_17361);
and U17532 (N_17532,N_17215,N_17301);
xnor U17533 (N_17533,N_17379,N_17308);
nor U17534 (N_17534,N_17306,N_17214);
nor U17535 (N_17535,N_17252,N_17376);
nand U17536 (N_17536,N_17345,N_17209);
and U17537 (N_17537,N_17315,N_17383);
or U17538 (N_17538,N_17373,N_17245);
xnor U17539 (N_17539,N_17284,N_17242);
and U17540 (N_17540,N_17349,N_17245);
xor U17541 (N_17541,N_17398,N_17224);
and U17542 (N_17542,N_17313,N_17217);
nand U17543 (N_17543,N_17225,N_17238);
nor U17544 (N_17544,N_17305,N_17365);
nand U17545 (N_17545,N_17388,N_17244);
xor U17546 (N_17546,N_17323,N_17384);
nor U17547 (N_17547,N_17246,N_17281);
or U17548 (N_17548,N_17349,N_17385);
nand U17549 (N_17549,N_17260,N_17241);
nor U17550 (N_17550,N_17253,N_17394);
and U17551 (N_17551,N_17359,N_17228);
nand U17552 (N_17552,N_17260,N_17333);
nand U17553 (N_17553,N_17353,N_17360);
nor U17554 (N_17554,N_17210,N_17321);
xor U17555 (N_17555,N_17229,N_17305);
or U17556 (N_17556,N_17281,N_17221);
nor U17557 (N_17557,N_17284,N_17308);
xor U17558 (N_17558,N_17211,N_17200);
and U17559 (N_17559,N_17363,N_17322);
nor U17560 (N_17560,N_17257,N_17370);
nor U17561 (N_17561,N_17395,N_17383);
nand U17562 (N_17562,N_17320,N_17302);
and U17563 (N_17563,N_17390,N_17215);
and U17564 (N_17564,N_17350,N_17292);
nand U17565 (N_17565,N_17320,N_17364);
or U17566 (N_17566,N_17382,N_17291);
or U17567 (N_17567,N_17394,N_17271);
and U17568 (N_17568,N_17312,N_17315);
and U17569 (N_17569,N_17299,N_17389);
xor U17570 (N_17570,N_17366,N_17295);
or U17571 (N_17571,N_17291,N_17227);
nand U17572 (N_17572,N_17305,N_17341);
and U17573 (N_17573,N_17254,N_17361);
or U17574 (N_17574,N_17253,N_17282);
or U17575 (N_17575,N_17219,N_17263);
xor U17576 (N_17576,N_17305,N_17368);
xor U17577 (N_17577,N_17367,N_17338);
nor U17578 (N_17578,N_17382,N_17362);
and U17579 (N_17579,N_17351,N_17265);
or U17580 (N_17580,N_17389,N_17211);
and U17581 (N_17581,N_17361,N_17335);
and U17582 (N_17582,N_17213,N_17350);
and U17583 (N_17583,N_17236,N_17378);
or U17584 (N_17584,N_17245,N_17336);
xnor U17585 (N_17585,N_17255,N_17210);
nand U17586 (N_17586,N_17228,N_17349);
xnor U17587 (N_17587,N_17265,N_17234);
nand U17588 (N_17588,N_17314,N_17295);
nor U17589 (N_17589,N_17232,N_17367);
or U17590 (N_17590,N_17299,N_17242);
xnor U17591 (N_17591,N_17297,N_17226);
xor U17592 (N_17592,N_17329,N_17249);
xnor U17593 (N_17593,N_17215,N_17233);
nor U17594 (N_17594,N_17248,N_17377);
nor U17595 (N_17595,N_17200,N_17363);
and U17596 (N_17596,N_17267,N_17258);
nand U17597 (N_17597,N_17314,N_17229);
nor U17598 (N_17598,N_17215,N_17265);
and U17599 (N_17599,N_17201,N_17351);
nand U17600 (N_17600,N_17576,N_17475);
or U17601 (N_17601,N_17577,N_17422);
nor U17602 (N_17602,N_17508,N_17500);
nor U17603 (N_17603,N_17499,N_17466);
xor U17604 (N_17604,N_17518,N_17497);
nand U17605 (N_17605,N_17540,N_17558);
xnor U17606 (N_17606,N_17566,N_17505);
nor U17607 (N_17607,N_17568,N_17457);
and U17608 (N_17608,N_17517,N_17541);
nor U17609 (N_17609,N_17592,N_17491);
xor U17610 (N_17610,N_17573,N_17461);
and U17611 (N_17611,N_17570,N_17595);
and U17612 (N_17612,N_17522,N_17582);
nand U17613 (N_17613,N_17429,N_17597);
or U17614 (N_17614,N_17528,N_17591);
nor U17615 (N_17615,N_17534,N_17453);
nand U17616 (N_17616,N_17504,N_17551);
nor U17617 (N_17617,N_17478,N_17542);
nand U17618 (N_17618,N_17445,N_17472);
and U17619 (N_17619,N_17520,N_17511);
and U17620 (N_17620,N_17503,N_17436);
nand U17621 (N_17621,N_17572,N_17507);
nand U17622 (N_17622,N_17408,N_17424);
or U17623 (N_17623,N_17409,N_17562);
and U17624 (N_17624,N_17585,N_17479);
nor U17625 (N_17625,N_17513,N_17404);
or U17626 (N_17626,N_17543,N_17403);
or U17627 (N_17627,N_17406,N_17578);
and U17628 (N_17628,N_17455,N_17527);
and U17629 (N_17629,N_17529,N_17432);
nand U17630 (N_17630,N_17579,N_17548);
nand U17631 (N_17631,N_17456,N_17593);
or U17632 (N_17632,N_17599,N_17598);
nand U17633 (N_17633,N_17571,N_17483);
or U17634 (N_17634,N_17416,N_17468);
nand U17635 (N_17635,N_17430,N_17405);
nand U17636 (N_17636,N_17485,N_17559);
xor U17637 (N_17637,N_17428,N_17512);
and U17638 (N_17638,N_17427,N_17470);
and U17639 (N_17639,N_17484,N_17425);
nor U17640 (N_17640,N_17426,N_17423);
xnor U17641 (N_17641,N_17531,N_17496);
xnor U17642 (N_17642,N_17567,N_17526);
xor U17643 (N_17643,N_17437,N_17557);
and U17644 (N_17644,N_17596,N_17501);
xnor U17645 (N_17645,N_17494,N_17469);
xnor U17646 (N_17646,N_17441,N_17417);
nor U17647 (N_17647,N_17574,N_17550);
and U17648 (N_17648,N_17546,N_17462);
xnor U17649 (N_17649,N_17509,N_17400);
nor U17650 (N_17650,N_17487,N_17476);
nand U17651 (N_17651,N_17510,N_17556);
xor U17652 (N_17652,N_17449,N_17467);
xnor U17653 (N_17653,N_17459,N_17502);
nand U17654 (N_17654,N_17435,N_17533);
xnor U17655 (N_17655,N_17565,N_17547);
xor U17656 (N_17656,N_17473,N_17521);
xor U17657 (N_17657,N_17458,N_17495);
or U17658 (N_17658,N_17587,N_17535);
and U17659 (N_17659,N_17401,N_17460);
nand U17660 (N_17660,N_17444,N_17482);
and U17661 (N_17661,N_17536,N_17433);
or U17662 (N_17662,N_17538,N_17464);
nor U17663 (N_17663,N_17465,N_17580);
nor U17664 (N_17664,N_17523,N_17537);
and U17665 (N_17665,N_17442,N_17515);
xor U17666 (N_17666,N_17563,N_17418);
or U17667 (N_17667,N_17569,N_17506);
nand U17668 (N_17668,N_17519,N_17560);
nand U17669 (N_17669,N_17584,N_17588);
nor U17670 (N_17670,N_17490,N_17481);
nand U17671 (N_17671,N_17413,N_17514);
nor U17672 (N_17672,N_17415,N_17471);
and U17673 (N_17673,N_17452,N_17564);
or U17674 (N_17674,N_17492,N_17554);
xor U17675 (N_17675,N_17488,N_17553);
nand U17676 (N_17676,N_17421,N_17447);
or U17677 (N_17677,N_17463,N_17486);
nand U17678 (N_17678,N_17443,N_17489);
or U17679 (N_17679,N_17414,N_17454);
nand U17680 (N_17680,N_17589,N_17561);
and U17681 (N_17681,N_17450,N_17419);
or U17682 (N_17682,N_17594,N_17439);
xnor U17683 (N_17683,N_17477,N_17431);
nor U17684 (N_17684,N_17539,N_17480);
nand U17685 (N_17685,N_17549,N_17410);
or U17686 (N_17686,N_17532,N_17446);
or U17687 (N_17687,N_17555,N_17525);
or U17688 (N_17688,N_17434,N_17474);
xor U17689 (N_17689,N_17516,N_17583);
nand U17690 (N_17690,N_17544,N_17412);
nor U17691 (N_17691,N_17438,N_17407);
nor U17692 (N_17692,N_17545,N_17448);
xnor U17693 (N_17693,N_17524,N_17440);
and U17694 (N_17694,N_17402,N_17590);
or U17695 (N_17695,N_17530,N_17552);
nand U17696 (N_17696,N_17420,N_17493);
nand U17697 (N_17697,N_17451,N_17581);
xnor U17698 (N_17698,N_17498,N_17586);
xor U17699 (N_17699,N_17575,N_17411);
or U17700 (N_17700,N_17530,N_17476);
or U17701 (N_17701,N_17576,N_17580);
xnor U17702 (N_17702,N_17464,N_17522);
xnor U17703 (N_17703,N_17589,N_17553);
nand U17704 (N_17704,N_17451,N_17544);
nor U17705 (N_17705,N_17428,N_17589);
or U17706 (N_17706,N_17517,N_17540);
or U17707 (N_17707,N_17416,N_17590);
nand U17708 (N_17708,N_17502,N_17470);
nor U17709 (N_17709,N_17588,N_17438);
nor U17710 (N_17710,N_17515,N_17505);
and U17711 (N_17711,N_17419,N_17468);
nand U17712 (N_17712,N_17477,N_17418);
xor U17713 (N_17713,N_17584,N_17575);
nand U17714 (N_17714,N_17404,N_17435);
and U17715 (N_17715,N_17446,N_17536);
nand U17716 (N_17716,N_17438,N_17509);
xnor U17717 (N_17717,N_17517,N_17436);
or U17718 (N_17718,N_17583,N_17552);
xnor U17719 (N_17719,N_17567,N_17555);
nand U17720 (N_17720,N_17452,N_17432);
nor U17721 (N_17721,N_17522,N_17520);
or U17722 (N_17722,N_17563,N_17526);
nand U17723 (N_17723,N_17405,N_17414);
xor U17724 (N_17724,N_17463,N_17501);
nand U17725 (N_17725,N_17554,N_17568);
and U17726 (N_17726,N_17529,N_17590);
and U17727 (N_17727,N_17461,N_17465);
or U17728 (N_17728,N_17534,N_17458);
and U17729 (N_17729,N_17473,N_17544);
or U17730 (N_17730,N_17582,N_17587);
nand U17731 (N_17731,N_17579,N_17539);
or U17732 (N_17732,N_17504,N_17429);
xnor U17733 (N_17733,N_17470,N_17567);
or U17734 (N_17734,N_17467,N_17547);
or U17735 (N_17735,N_17533,N_17598);
and U17736 (N_17736,N_17599,N_17400);
xor U17737 (N_17737,N_17545,N_17599);
xnor U17738 (N_17738,N_17595,N_17437);
nand U17739 (N_17739,N_17470,N_17576);
nand U17740 (N_17740,N_17511,N_17467);
and U17741 (N_17741,N_17535,N_17568);
nor U17742 (N_17742,N_17459,N_17505);
nor U17743 (N_17743,N_17499,N_17599);
and U17744 (N_17744,N_17498,N_17509);
nor U17745 (N_17745,N_17579,N_17453);
nor U17746 (N_17746,N_17517,N_17547);
nor U17747 (N_17747,N_17553,N_17433);
and U17748 (N_17748,N_17401,N_17473);
xor U17749 (N_17749,N_17530,N_17504);
and U17750 (N_17750,N_17457,N_17471);
or U17751 (N_17751,N_17445,N_17459);
xnor U17752 (N_17752,N_17509,N_17547);
nor U17753 (N_17753,N_17470,N_17591);
nand U17754 (N_17754,N_17464,N_17490);
nand U17755 (N_17755,N_17505,N_17418);
xnor U17756 (N_17756,N_17424,N_17543);
xnor U17757 (N_17757,N_17486,N_17556);
nand U17758 (N_17758,N_17598,N_17517);
or U17759 (N_17759,N_17448,N_17529);
nor U17760 (N_17760,N_17438,N_17472);
xnor U17761 (N_17761,N_17597,N_17567);
nor U17762 (N_17762,N_17509,N_17576);
or U17763 (N_17763,N_17419,N_17555);
xor U17764 (N_17764,N_17536,N_17434);
nand U17765 (N_17765,N_17533,N_17586);
nand U17766 (N_17766,N_17448,N_17474);
xnor U17767 (N_17767,N_17555,N_17459);
or U17768 (N_17768,N_17471,N_17414);
and U17769 (N_17769,N_17440,N_17471);
or U17770 (N_17770,N_17585,N_17424);
xor U17771 (N_17771,N_17440,N_17486);
or U17772 (N_17772,N_17490,N_17436);
xnor U17773 (N_17773,N_17508,N_17538);
xor U17774 (N_17774,N_17520,N_17418);
xnor U17775 (N_17775,N_17440,N_17542);
and U17776 (N_17776,N_17505,N_17467);
xnor U17777 (N_17777,N_17584,N_17491);
and U17778 (N_17778,N_17568,N_17513);
xor U17779 (N_17779,N_17486,N_17482);
nand U17780 (N_17780,N_17415,N_17506);
xnor U17781 (N_17781,N_17568,N_17532);
and U17782 (N_17782,N_17576,N_17467);
nand U17783 (N_17783,N_17581,N_17413);
and U17784 (N_17784,N_17559,N_17576);
nand U17785 (N_17785,N_17546,N_17580);
xnor U17786 (N_17786,N_17590,N_17578);
xor U17787 (N_17787,N_17463,N_17517);
nor U17788 (N_17788,N_17593,N_17489);
and U17789 (N_17789,N_17537,N_17497);
nand U17790 (N_17790,N_17406,N_17421);
or U17791 (N_17791,N_17592,N_17514);
and U17792 (N_17792,N_17538,N_17510);
nor U17793 (N_17793,N_17455,N_17425);
xor U17794 (N_17794,N_17402,N_17465);
xnor U17795 (N_17795,N_17512,N_17470);
nand U17796 (N_17796,N_17547,N_17532);
and U17797 (N_17797,N_17544,N_17496);
nor U17798 (N_17798,N_17544,N_17599);
and U17799 (N_17799,N_17597,N_17578);
xor U17800 (N_17800,N_17684,N_17669);
nand U17801 (N_17801,N_17775,N_17627);
or U17802 (N_17802,N_17625,N_17740);
or U17803 (N_17803,N_17710,N_17634);
and U17804 (N_17804,N_17778,N_17753);
xnor U17805 (N_17805,N_17748,N_17781);
nand U17806 (N_17806,N_17703,N_17730);
nand U17807 (N_17807,N_17648,N_17605);
xor U17808 (N_17808,N_17642,N_17606);
xor U17809 (N_17809,N_17737,N_17711);
nor U17810 (N_17810,N_17796,N_17609);
or U17811 (N_17811,N_17664,N_17666);
or U17812 (N_17812,N_17745,N_17799);
or U17813 (N_17813,N_17688,N_17665);
nand U17814 (N_17814,N_17706,N_17747);
and U17815 (N_17815,N_17749,N_17783);
nand U17816 (N_17816,N_17617,N_17601);
xnor U17817 (N_17817,N_17659,N_17776);
nand U17818 (N_17818,N_17717,N_17785);
or U17819 (N_17819,N_17699,N_17779);
xor U17820 (N_17820,N_17720,N_17768);
nand U17821 (N_17821,N_17772,N_17741);
and U17822 (N_17822,N_17789,N_17687);
or U17823 (N_17823,N_17724,N_17707);
nor U17824 (N_17824,N_17610,N_17673);
nand U17825 (N_17825,N_17769,N_17639);
nand U17826 (N_17826,N_17655,N_17645);
and U17827 (N_17827,N_17794,N_17679);
nand U17828 (N_17828,N_17692,N_17672);
nor U17829 (N_17829,N_17670,N_17722);
xor U17830 (N_17830,N_17628,N_17758);
and U17831 (N_17831,N_17675,N_17721);
nand U17832 (N_17832,N_17759,N_17698);
nor U17833 (N_17833,N_17764,N_17602);
nand U17834 (N_17834,N_17654,N_17715);
nor U17835 (N_17835,N_17790,N_17668);
nor U17836 (N_17836,N_17784,N_17621);
and U17837 (N_17837,N_17690,N_17786);
xnor U17838 (N_17838,N_17643,N_17638);
xor U17839 (N_17839,N_17713,N_17716);
or U17840 (N_17840,N_17732,N_17693);
nand U17841 (N_17841,N_17614,N_17653);
or U17842 (N_17842,N_17705,N_17736);
nor U17843 (N_17843,N_17657,N_17742);
nor U17844 (N_17844,N_17682,N_17782);
nor U17845 (N_17845,N_17700,N_17636);
and U17846 (N_17846,N_17680,N_17656);
nand U17847 (N_17847,N_17754,N_17704);
xor U17848 (N_17848,N_17734,N_17774);
or U17849 (N_17849,N_17795,N_17708);
nor U17850 (N_17850,N_17702,N_17647);
nand U17851 (N_17851,N_17600,N_17773);
nor U17852 (N_17852,N_17616,N_17723);
nor U17853 (N_17853,N_17622,N_17735);
and U17854 (N_17854,N_17607,N_17685);
or U17855 (N_17855,N_17650,N_17671);
or U17856 (N_17856,N_17660,N_17752);
nand U17857 (N_17857,N_17603,N_17651);
and U17858 (N_17858,N_17683,N_17677);
and U17859 (N_17859,N_17726,N_17714);
xor U17860 (N_17860,N_17739,N_17760);
nand U17861 (N_17861,N_17765,N_17644);
or U17862 (N_17862,N_17797,N_17751);
xnor U17863 (N_17863,N_17676,N_17631);
and U17864 (N_17864,N_17767,N_17623);
and U17865 (N_17865,N_17697,N_17728);
nand U17866 (N_17866,N_17691,N_17712);
nor U17867 (N_17867,N_17719,N_17780);
xnor U17868 (N_17868,N_17618,N_17725);
and U17869 (N_17869,N_17608,N_17750);
or U17870 (N_17870,N_17770,N_17663);
xnor U17871 (N_17871,N_17718,N_17755);
nor U17872 (N_17872,N_17701,N_17633);
nor U17873 (N_17873,N_17761,N_17766);
nand U17874 (N_17874,N_17630,N_17694);
and U17875 (N_17875,N_17788,N_17635);
or U17876 (N_17876,N_17624,N_17738);
nand U17877 (N_17877,N_17729,N_17787);
nor U17878 (N_17878,N_17727,N_17613);
nor U17879 (N_17879,N_17695,N_17632);
xnor U17880 (N_17880,N_17646,N_17667);
xor U17881 (N_17881,N_17756,N_17743);
nand U17882 (N_17882,N_17777,N_17757);
nand U17883 (N_17883,N_17612,N_17744);
nand U17884 (N_17884,N_17637,N_17674);
and U17885 (N_17885,N_17686,N_17661);
and U17886 (N_17886,N_17798,N_17731);
nand U17887 (N_17887,N_17793,N_17763);
or U17888 (N_17888,N_17619,N_17762);
and U17889 (N_17889,N_17746,N_17662);
or U17890 (N_17890,N_17641,N_17791);
and U17891 (N_17891,N_17658,N_17640);
and U17892 (N_17892,N_17620,N_17792);
xnor U17893 (N_17893,N_17709,N_17611);
and U17894 (N_17894,N_17733,N_17689);
or U17895 (N_17895,N_17696,N_17681);
or U17896 (N_17896,N_17626,N_17629);
nor U17897 (N_17897,N_17771,N_17649);
or U17898 (N_17898,N_17604,N_17678);
nor U17899 (N_17899,N_17615,N_17652);
nand U17900 (N_17900,N_17749,N_17738);
nor U17901 (N_17901,N_17726,N_17785);
xor U17902 (N_17902,N_17785,N_17706);
xnor U17903 (N_17903,N_17677,N_17631);
and U17904 (N_17904,N_17784,N_17679);
nand U17905 (N_17905,N_17603,N_17702);
nor U17906 (N_17906,N_17640,N_17785);
nor U17907 (N_17907,N_17624,N_17669);
xnor U17908 (N_17908,N_17640,N_17681);
or U17909 (N_17909,N_17703,N_17775);
nor U17910 (N_17910,N_17601,N_17685);
nor U17911 (N_17911,N_17798,N_17609);
xor U17912 (N_17912,N_17739,N_17748);
xnor U17913 (N_17913,N_17621,N_17637);
xnor U17914 (N_17914,N_17623,N_17720);
and U17915 (N_17915,N_17702,N_17733);
or U17916 (N_17916,N_17750,N_17712);
and U17917 (N_17917,N_17674,N_17751);
and U17918 (N_17918,N_17783,N_17692);
or U17919 (N_17919,N_17740,N_17700);
xnor U17920 (N_17920,N_17736,N_17762);
and U17921 (N_17921,N_17694,N_17712);
xor U17922 (N_17922,N_17719,N_17698);
xnor U17923 (N_17923,N_17794,N_17734);
and U17924 (N_17924,N_17652,N_17728);
xnor U17925 (N_17925,N_17606,N_17776);
nand U17926 (N_17926,N_17709,N_17715);
nand U17927 (N_17927,N_17794,N_17753);
or U17928 (N_17928,N_17791,N_17644);
nor U17929 (N_17929,N_17603,N_17796);
and U17930 (N_17930,N_17654,N_17672);
or U17931 (N_17931,N_17680,N_17677);
or U17932 (N_17932,N_17762,N_17695);
nand U17933 (N_17933,N_17726,N_17754);
nand U17934 (N_17934,N_17746,N_17689);
xor U17935 (N_17935,N_17701,N_17626);
xor U17936 (N_17936,N_17609,N_17739);
nor U17937 (N_17937,N_17637,N_17752);
or U17938 (N_17938,N_17704,N_17735);
nor U17939 (N_17939,N_17763,N_17670);
nand U17940 (N_17940,N_17613,N_17668);
or U17941 (N_17941,N_17632,N_17674);
nand U17942 (N_17942,N_17706,N_17621);
or U17943 (N_17943,N_17730,N_17633);
or U17944 (N_17944,N_17657,N_17632);
nor U17945 (N_17945,N_17633,N_17657);
nor U17946 (N_17946,N_17617,N_17644);
nand U17947 (N_17947,N_17643,N_17733);
or U17948 (N_17948,N_17793,N_17622);
xor U17949 (N_17949,N_17633,N_17629);
and U17950 (N_17950,N_17735,N_17729);
nand U17951 (N_17951,N_17797,N_17680);
nand U17952 (N_17952,N_17781,N_17618);
and U17953 (N_17953,N_17712,N_17686);
nand U17954 (N_17954,N_17603,N_17637);
xnor U17955 (N_17955,N_17743,N_17753);
or U17956 (N_17956,N_17787,N_17730);
nor U17957 (N_17957,N_17737,N_17601);
nor U17958 (N_17958,N_17793,N_17673);
nor U17959 (N_17959,N_17632,N_17683);
and U17960 (N_17960,N_17794,N_17683);
nor U17961 (N_17961,N_17608,N_17665);
xnor U17962 (N_17962,N_17731,N_17670);
xnor U17963 (N_17963,N_17695,N_17767);
or U17964 (N_17964,N_17761,N_17740);
xnor U17965 (N_17965,N_17708,N_17667);
or U17966 (N_17966,N_17757,N_17707);
nor U17967 (N_17967,N_17600,N_17656);
nand U17968 (N_17968,N_17700,N_17753);
and U17969 (N_17969,N_17712,N_17690);
nor U17970 (N_17970,N_17637,N_17648);
xnor U17971 (N_17971,N_17784,N_17743);
and U17972 (N_17972,N_17614,N_17645);
and U17973 (N_17973,N_17683,N_17687);
nor U17974 (N_17974,N_17608,N_17606);
nand U17975 (N_17975,N_17729,N_17667);
and U17976 (N_17976,N_17671,N_17690);
and U17977 (N_17977,N_17787,N_17661);
nor U17978 (N_17978,N_17777,N_17609);
nor U17979 (N_17979,N_17792,N_17621);
or U17980 (N_17980,N_17673,N_17716);
nor U17981 (N_17981,N_17644,N_17653);
nor U17982 (N_17982,N_17780,N_17624);
xnor U17983 (N_17983,N_17790,N_17737);
xor U17984 (N_17984,N_17705,N_17694);
xor U17985 (N_17985,N_17732,N_17641);
xnor U17986 (N_17986,N_17645,N_17745);
or U17987 (N_17987,N_17620,N_17725);
nor U17988 (N_17988,N_17786,N_17770);
xnor U17989 (N_17989,N_17652,N_17689);
and U17990 (N_17990,N_17793,N_17731);
nand U17991 (N_17991,N_17796,N_17643);
nor U17992 (N_17992,N_17773,N_17611);
or U17993 (N_17993,N_17610,N_17676);
or U17994 (N_17994,N_17678,N_17790);
nor U17995 (N_17995,N_17668,N_17707);
nand U17996 (N_17996,N_17652,N_17608);
xor U17997 (N_17997,N_17769,N_17785);
xnor U17998 (N_17998,N_17748,N_17709);
nor U17999 (N_17999,N_17619,N_17626);
xnor U18000 (N_18000,N_17852,N_17880);
nor U18001 (N_18001,N_17883,N_17895);
xnor U18002 (N_18002,N_17942,N_17952);
or U18003 (N_18003,N_17807,N_17937);
or U18004 (N_18004,N_17948,N_17832);
or U18005 (N_18005,N_17874,N_17847);
and U18006 (N_18006,N_17823,N_17935);
nand U18007 (N_18007,N_17958,N_17955);
or U18008 (N_18008,N_17882,N_17875);
nor U18009 (N_18009,N_17985,N_17914);
xor U18010 (N_18010,N_17850,N_17876);
xor U18011 (N_18011,N_17970,N_17949);
nor U18012 (N_18012,N_17996,N_17956);
nor U18013 (N_18013,N_17826,N_17978);
or U18014 (N_18014,N_17809,N_17897);
or U18015 (N_18015,N_17909,N_17974);
nor U18016 (N_18016,N_17884,N_17979);
or U18017 (N_18017,N_17907,N_17997);
and U18018 (N_18018,N_17924,N_17941);
and U18019 (N_18019,N_17857,N_17841);
xor U18020 (N_18020,N_17873,N_17911);
nand U18021 (N_18021,N_17969,N_17959);
and U18022 (N_18022,N_17851,N_17886);
nor U18023 (N_18023,N_17889,N_17861);
nand U18024 (N_18024,N_17939,N_17840);
and U18025 (N_18025,N_17928,N_17819);
or U18026 (N_18026,N_17825,N_17957);
or U18027 (N_18027,N_17870,N_17910);
nor U18028 (N_18028,N_17922,N_17971);
xor U18029 (N_18029,N_17860,N_17842);
and U18030 (N_18030,N_17920,N_17871);
nand U18031 (N_18031,N_17991,N_17918);
xnor U18032 (N_18032,N_17810,N_17872);
and U18033 (N_18033,N_17856,N_17834);
and U18034 (N_18034,N_17829,N_17862);
nor U18035 (N_18035,N_17866,N_17990);
or U18036 (N_18036,N_17953,N_17986);
and U18037 (N_18037,N_17845,N_17858);
xnor U18038 (N_18038,N_17988,N_17863);
or U18039 (N_18039,N_17802,N_17905);
nand U18040 (N_18040,N_17814,N_17805);
xnor U18041 (N_18041,N_17963,N_17867);
nand U18042 (N_18042,N_17902,N_17891);
or U18043 (N_18043,N_17936,N_17833);
nand U18044 (N_18044,N_17919,N_17906);
and U18045 (N_18045,N_17831,N_17967);
nor U18046 (N_18046,N_17878,N_17830);
nor U18047 (N_18047,N_17813,N_17839);
or U18048 (N_18048,N_17938,N_17943);
and U18049 (N_18049,N_17898,N_17903);
and U18050 (N_18050,N_17994,N_17993);
or U18051 (N_18051,N_17844,N_17975);
xnor U18052 (N_18052,N_17923,N_17801);
nor U18053 (N_18053,N_17999,N_17917);
and U18054 (N_18054,N_17981,N_17859);
and U18055 (N_18055,N_17811,N_17894);
nand U18056 (N_18056,N_17890,N_17879);
or U18057 (N_18057,N_17968,N_17806);
nor U18058 (N_18058,N_17820,N_17838);
xor U18059 (N_18059,N_17822,N_17881);
or U18060 (N_18060,N_17925,N_17989);
nand U18061 (N_18061,N_17940,N_17932);
nand U18062 (N_18062,N_17992,N_17836);
or U18063 (N_18063,N_17916,N_17817);
nand U18064 (N_18064,N_17926,N_17960);
and U18065 (N_18065,N_17855,N_17885);
and U18066 (N_18066,N_17853,N_17913);
and U18067 (N_18067,N_17908,N_17892);
or U18068 (N_18068,N_17901,N_17854);
or U18069 (N_18069,N_17984,N_17899);
or U18070 (N_18070,N_17973,N_17998);
and U18071 (N_18071,N_17944,N_17828);
nor U18072 (N_18072,N_17951,N_17869);
nor U18073 (N_18073,N_17846,N_17900);
and U18074 (N_18074,N_17837,N_17921);
or U18075 (N_18075,N_17945,N_17868);
nor U18076 (N_18076,N_17934,N_17930);
xnor U18077 (N_18077,N_17965,N_17933);
xor U18078 (N_18078,N_17976,N_17864);
nor U18079 (N_18079,N_17824,N_17912);
xnor U18080 (N_18080,N_17929,N_17954);
xnor U18081 (N_18081,N_17849,N_17865);
or U18082 (N_18082,N_17808,N_17947);
or U18083 (N_18083,N_17982,N_17893);
xnor U18084 (N_18084,N_17816,N_17804);
and U18085 (N_18085,N_17983,N_17888);
nor U18086 (N_18086,N_17961,N_17972);
nand U18087 (N_18087,N_17950,N_17995);
nand U18088 (N_18088,N_17843,N_17896);
xnor U18089 (N_18089,N_17821,N_17931);
and U18090 (N_18090,N_17977,N_17915);
xnor U18091 (N_18091,N_17877,N_17964);
xnor U18092 (N_18092,N_17987,N_17966);
or U18093 (N_18093,N_17835,N_17818);
xor U18094 (N_18094,N_17815,N_17887);
nand U18095 (N_18095,N_17803,N_17848);
nand U18096 (N_18096,N_17946,N_17980);
xor U18097 (N_18097,N_17927,N_17904);
nand U18098 (N_18098,N_17962,N_17827);
and U18099 (N_18099,N_17812,N_17800);
nor U18100 (N_18100,N_17954,N_17903);
xor U18101 (N_18101,N_17805,N_17853);
and U18102 (N_18102,N_17825,N_17878);
and U18103 (N_18103,N_17866,N_17911);
and U18104 (N_18104,N_17806,N_17986);
xor U18105 (N_18105,N_17948,N_17842);
nor U18106 (N_18106,N_17968,N_17841);
or U18107 (N_18107,N_17803,N_17981);
or U18108 (N_18108,N_17928,N_17991);
or U18109 (N_18109,N_17975,N_17813);
nand U18110 (N_18110,N_17969,N_17871);
or U18111 (N_18111,N_17832,N_17985);
nand U18112 (N_18112,N_17923,N_17932);
nor U18113 (N_18113,N_17896,N_17834);
xor U18114 (N_18114,N_17867,N_17857);
nand U18115 (N_18115,N_17929,N_17985);
nand U18116 (N_18116,N_17837,N_17802);
nand U18117 (N_18117,N_17999,N_17880);
and U18118 (N_18118,N_17947,N_17954);
nand U18119 (N_18119,N_17959,N_17939);
nand U18120 (N_18120,N_17997,N_17878);
xor U18121 (N_18121,N_17819,N_17827);
nand U18122 (N_18122,N_17859,N_17845);
or U18123 (N_18123,N_17813,N_17916);
and U18124 (N_18124,N_17875,N_17991);
and U18125 (N_18125,N_17988,N_17895);
and U18126 (N_18126,N_17913,N_17931);
nor U18127 (N_18127,N_17824,N_17817);
xor U18128 (N_18128,N_17981,N_17995);
nand U18129 (N_18129,N_17817,N_17809);
xnor U18130 (N_18130,N_17985,N_17872);
and U18131 (N_18131,N_17804,N_17883);
nand U18132 (N_18132,N_17990,N_17896);
and U18133 (N_18133,N_17935,N_17868);
xor U18134 (N_18134,N_17838,N_17897);
nor U18135 (N_18135,N_17870,N_17866);
and U18136 (N_18136,N_17811,N_17962);
nor U18137 (N_18137,N_17833,N_17905);
or U18138 (N_18138,N_17952,N_17841);
nor U18139 (N_18139,N_17958,N_17978);
xor U18140 (N_18140,N_17833,N_17923);
nand U18141 (N_18141,N_17904,N_17875);
nor U18142 (N_18142,N_17998,N_17815);
xnor U18143 (N_18143,N_17878,N_17964);
xnor U18144 (N_18144,N_17838,N_17893);
nand U18145 (N_18145,N_17970,N_17994);
nor U18146 (N_18146,N_17814,N_17992);
nor U18147 (N_18147,N_17821,N_17958);
xnor U18148 (N_18148,N_17858,N_17976);
xor U18149 (N_18149,N_17987,N_17889);
and U18150 (N_18150,N_17979,N_17812);
nor U18151 (N_18151,N_17919,N_17920);
nor U18152 (N_18152,N_17938,N_17840);
xnor U18153 (N_18153,N_17914,N_17945);
or U18154 (N_18154,N_17951,N_17801);
nor U18155 (N_18155,N_17901,N_17951);
xnor U18156 (N_18156,N_17965,N_17952);
and U18157 (N_18157,N_17850,N_17860);
and U18158 (N_18158,N_17966,N_17945);
nor U18159 (N_18159,N_17885,N_17961);
xor U18160 (N_18160,N_17883,N_17928);
nor U18161 (N_18161,N_17928,N_17888);
or U18162 (N_18162,N_17863,N_17914);
and U18163 (N_18163,N_17967,N_17906);
and U18164 (N_18164,N_17835,N_17963);
nand U18165 (N_18165,N_17861,N_17865);
or U18166 (N_18166,N_17816,N_17928);
xor U18167 (N_18167,N_17835,N_17860);
or U18168 (N_18168,N_17962,N_17890);
and U18169 (N_18169,N_17812,N_17975);
and U18170 (N_18170,N_17881,N_17850);
and U18171 (N_18171,N_17861,N_17941);
xnor U18172 (N_18172,N_17894,N_17979);
xor U18173 (N_18173,N_17984,N_17838);
nand U18174 (N_18174,N_17823,N_17920);
xor U18175 (N_18175,N_17970,N_17901);
or U18176 (N_18176,N_17955,N_17896);
nand U18177 (N_18177,N_17916,N_17911);
xor U18178 (N_18178,N_17930,N_17883);
xor U18179 (N_18179,N_17963,N_17918);
nor U18180 (N_18180,N_17896,N_17818);
nand U18181 (N_18181,N_17924,N_17897);
or U18182 (N_18182,N_17931,N_17996);
nor U18183 (N_18183,N_17827,N_17813);
xnor U18184 (N_18184,N_17992,N_17894);
and U18185 (N_18185,N_17874,N_17877);
xor U18186 (N_18186,N_17820,N_17819);
nand U18187 (N_18187,N_17956,N_17987);
or U18188 (N_18188,N_17996,N_17948);
or U18189 (N_18189,N_17977,N_17965);
nor U18190 (N_18190,N_17964,N_17972);
xnor U18191 (N_18191,N_17894,N_17854);
or U18192 (N_18192,N_17956,N_17891);
and U18193 (N_18193,N_17931,N_17987);
nand U18194 (N_18194,N_17947,N_17935);
and U18195 (N_18195,N_17900,N_17977);
xor U18196 (N_18196,N_17875,N_17816);
or U18197 (N_18197,N_17892,N_17819);
or U18198 (N_18198,N_17941,N_17998);
and U18199 (N_18199,N_17919,N_17959);
and U18200 (N_18200,N_18102,N_18053);
and U18201 (N_18201,N_18022,N_18087);
xnor U18202 (N_18202,N_18111,N_18026);
or U18203 (N_18203,N_18161,N_18007);
nand U18204 (N_18204,N_18166,N_18067);
or U18205 (N_18205,N_18002,N_18016);
nor U18206 (N_18206,N_18080,N_18034);
nor U18207 (N_18207,N_18155,N_18120);
xnor U18208 (N_18208,N_18189,N_18044);
or U18209 (N_18209,N_18116,N_18049);
nor U18210 (N_18210,N_18184,N_18057);
or U18211 (N_18211,N_18181,N_18153);
xnor U18212 (N_18212,N_18165,N_18112);
and U18213 (N_18213,N_18142,N_18186);
nor U18214 (N_18214,N_18188,N_18000);
and U18215 (N_18215,N_18079,N_18129);
xor U18216 (N_18216,N_18084,N_18163);
or U18217 (N_18217,N_18004,N_18150);
nand U18218 (N_18218,N_18020,N_18170);
nor U18219 (N_18219,N_18193,N_18177);
xor U18220 (N_18220,N_18009,N_18179);
and U18221 (N_18221,N_18117,N_18063);
xor U18222 (N_18222,N_18023,N_18038);
or U18223 (N_18223,N_18115,N_18088);
nor U18224 (N_18224,N_18171,N_18172);
nor U18225 (N_18225,N_18035,N_18024);
nand U18226 (N_18226,N_18013,N_18059);
or U18227 (N_18227,N_18138,N_18083);
xnor U18228 (N_18228,N_18137,N_18182);
and U18229 (N_18229,N_18113,N_18109);
or U18230 (N_18230,N_18176,N_18040);
nor U18231 (N_18231,N_18028,N_18073);
nand U18232 (N_18232,N_18062,N_18173);
nand U18233 (N_18233,N_18042,N_18151);
nor U18234 (N_18234,N_18148,N_18114);
nor U18235 (N_18235,N_18123,N_18124);
or U18236 (N_18236,N_18082,N_18036);
xor U18237 (N_18237,N_18106,N_18043);
xnor U18238 (N_18238,N_18191,N_18012);
xor U18239 (N_18239,N_18046,N_18101);
nor U18240 (N_18240,N_18064,N_18144);
nand U18241 (N_18241,N_18019,N_18003);
and U18242 (N_18242,N_18135,N_18066);
nor U18243 (N_18243,N_18133,N_18199);
or U18244 (N_18244,N_18090,N_18131);
or U18245 (N_18245,N_18055,N_18006);
nor U18246 (N_18246,N_18010,N_18018);
xnor U18247 (N_18247,N_18168,N_18098);
nor U18248 (N_18248,N_18056,N_18195);
nor U18249 (N_18249,N_18132,N_18011);
nor U18250 (N_18250,N_18078,N_18190);
nor U18251 (N_18251,N_18118,N_18174);
xnor U18252 (N_18252,N_18180,N_18110);
or U18253 (N_18253,N_18141,N_18074);
and U18254 (N_18254,N_18052,N_18050);
nand U18255 (N_18255,N_18198,N_18158);
nand U18256 (N_18256,N_18029,N_18122);
nor U18257 (N_18257,N_18121,N_18167);
or U18258 (N_18258,N_18068,N_18089);
xnor U18259 (N_18259,N_18025,N_18145);
or U18260 (N_18260,N_18054,N_18081);
nand U18261 (N_18261,N_18146,N_18143);
nand U18262 (N_18262,N_18149,N_18070);
nand U18263 (N_18263,N_18126,N_18128);
xor U18264 (N_18264,N_18162,N_18060);
xnor U18265 (N_18265,N_18157,N_18021);
nand U18266 (N_18266,N_18094,N_18017);
or U18267 (N_18267,N_18105,N_18093);
or U18268 (N_18268,N_18095,N_18069);
or U18269 (N_18269,N_18072,N_18075);
nand U18270 (N_18270,N_18048,N_18139);
and U18271 (N_18271,N_18183,N_18096);
nor U18272 (N_18272,N_18085,N_18061);
xnor U18273 (N_18273,N_18071,N_18001);
nor U18274 (N_18274,N_18108,N_18107);
or U18275 (N_18275,N_18027,N_18152);
xnor U18276 (N_18276,N_18104,N_18051);
nor U18277 (N_18277,N_18041,N_18154);
or U18278 (N_18278,N_18032,N_18130);
nand U18279 (N_18279,N_18008,N_18086);
and U18280 (N_18280,N_18197,N_18015);
xor U18281 (N_18281,N_18125,N_18091);
or U18282 (N_18282,N_18103,N_18187);
or U18283 (N_18283,N_18119,N_18194);
and U18284 (N_18284,N_18005,N_18039);
or U18285 (N_18285,N_18076,N_18185);
nor U18286 (N_18286,N_18045,N_18037);
or U18287 (N_18287,N_18058,N_18014);
nand U18288 (N_18288,N_18160,N_18030);
nor U18289 (N_18289,N_18178,N_18192);
and U18290 (N_18290,N_18136,N_18047);
or U18291 (N_18291,N_18147,N_18175);
and U18292 (N_18292,N_18169,N_18031);
or U18293 (N_18293,N_18196,N_18127);
or U18294 (N_18294,N_18100,N_18092);
or U18295 (N_18295,N_18164,N_18140);
and U18296 (N_18296,N_18033,N_18159);
nand U18297 (N_18297,N_18065,N_18097);
nor U18298 (N_18298,N_18134,N_18077);
xor U18299 (N_18299,N_18156,N_18099);
and U18300 (N_18300,N_18080,N_18074);
or U18301 (N_18301,N_18183,N_18093);
and U18302 (N_18302,N_18037,N_18185);
nor U18303 (N_18303,N_18132,N_18157);
xnor U18304 (N_18304,N_18083,N_18123);
nor U18305 (N_18305,N_18079,N_18111);
and U18306 (N_18306,N_18024,N_18080);
nand U18307 (N_18307,N_18010,N_18109);
or U18308 (N_18308,N_18035,N_18152);
nor U18309 (N_18309,N_18190,N_18106);
nor U18310 (N_18310,N_18096,N_18187);
or U18311 (N_18311,N_18065,N_18193);
or U18312 (N_18312,N_18128,N_18193);
and U18313 (N_18313,N_18164,N_18147);
nand U18314 (N_18314,N_18177,N_18089);
and U18315 (N_18315,N_18127,N_18186);
xor U18316 (N_18316,N_18009,N_18157);
nor U18317 (N_18317,N_18084,N_18108);
or U18318 (N_18318,N_18159,N_18138);
or U18319 (N_18319,N_18182,N_18049);
xnor U18320 (N_18320,N_18098,N_18136);
xnor U18321 (N_18321,N_18036,N_18191);
nand U18322 (N_18322,N_18129,N_18046);
xor U18323 (N_18323,N_18017,N_18134);
xor U18324 (N_18324,N_18017,N_18172);
nand U18325 (N_18325,N_18023,N_18082);
nor U18326 (N_18326,N_18173,N_18052);
and U18327 (N_18327,N_18011,N_18060);
and U18328 (N_18328,N_18142,N_18013);
and U18329 (N_18329,N_18014,N_18077);
nand U18330 (N_18330,N_18013,N_18038);
nor U18331 (N_18331,N_18166,N_18008);
nand U18332 (N_18332,N_18111,N_18048);
and U18333 (N_18333,N_18125,N_18004);
or U18334 (N_18334,N_18086,N_18184);
nor U18335 (N_18335,N_18165,N_18121);
and U18336 (N_18336,N_18105,N_18188);
and U18337 (N_18337,N_18001,N_18179);
or U18338 (N_18338,N_18150,N_18110);
and U18339 (N_18339,N_18194,N_18131);
nor U18340 (N_18340,N_18056,N_18060);
nand U18341 (N_18341,N_18189,N_18109);
nand U18342 (N_18342,N_18146,N_18182);
or U18343 (N_18343,N_18094,N_18180);
nor U18344 (N_18344,N_18046,N_18130);
or U18345 (N_18345,N_18119,N_18023);
nand U18346 (N_18346,N_18012,N_18059);
or U18347 (N_18347,N_18007,N_18177);
or U18348 (N_18348,N_18014,N_18174);
nor U18349 (N_18349,N_18010,N_18048);
nand U18350 (N_18350,N_18034,N_18093);
or U18351 (N_18351,N_18108,N_18162);
xnor U18352 (N_18352,N_18101,N_18164);
nand U18353 (N_18353,N_18109,N_18014);
or U18354 (N_18354,N_18059,N_18123);
nand U18355 (N_18355,N_18002,N_18054);
nor U18356 (N_18356,N_18134,N_18199);
xor U18357 (N_18357,N_18061,N_18040);
and U18358 (N_18358,N_18037,N_18034);
nor U18359 (N_18359,N_18028,N_18091);
nand U18360 (N_18360,N_18189,N_18080);
nand U18361 (N_18361,N_18130,N_18104);
and U18362 (N_18362,N_18117,N_18119);
xnor U18363 (N_18363,N_18032,N_18118);
and U18364 (N_18364,N_18154,N_18046);
xor U18365 (N_18365,N_18160,N_18175);
or U18366 (N_18366,N_18008,N_18033);
nor U18367 (N_18367,N_18063,N_18026);
and U18368 (N_18368,N_18191,N_18094);
xor U18369 (N_18369,N_18045,N_18089);
and U18370 (N_18370,N_18135,N_18021);
nand U18371 (N_18371,N_18123,N_18007);
and U18372 (N_18372,N_18142,N_18191);
xor U18373 (N_18373,N_18112,N_18088);
and U18374 (N_18374,N_18024,N_18132);
and U18375 (N_18375,N_18156,N_18050);
nand U18376 (N_18376,N_18020,N_18061);
and U18377 (N_18377,N_18022,N_18069);
and U18378 (N_18378,N_18005,N_18138);
and U18379 (N_18379,N_18159,N_18090);
nor U18380 (N_18380,N_18103,N_18017);
nand U18381 (N_18381,N_18074,N_18031);
and U18382 (N_18382,N_18033,N_18181);
and U18383 (N_18383,N_18085,N_18158);
nor U18384 (N_18384,N_18195,N_18025);
and U18385 (N_18385,N_18145,N_18141);
nor U18386 (N_18386,N_18082,N_18005);
xnor U18387 (N_18387,N_18024,N_18147);
nor U18388 (N_18388,N_18157,N_18113);
and U18389 (N_18389,N_18186,N_18143);
nor U18390 (N_18390,N_18196,N_18161);
xor U18391 (N_18391,N_18156,N_18063);
nand U18392 (N_18392,N_18086,N_18127);
or U18393 (N_18393,N_18019,N_18157);
nor U18394 (N_18394,N_18018,N_18124);
or U18395 (N_18395,N_18005,N_18192);
nand U18396 (N_18396,N_18136,N_18088);
or U18397 (N_18397,N_18128,N_18179);
nand U18398 (N_18398,N_18025,N_18088);
and U18399 (N_18399,N_18096,N_18041);
xnor U18400 (N_18400,N_18393,N_18211);
xor U18401 (N_18401,N_18209,N_18361);
and U18402 (N_18402,N_18318,N_18220);
xor U18403 (N_18403,N_18308,N_18249);
and U18404 (N_18404,N_18208,N_18265);
nand U18405 (N_18405,N_18229,N_18330);
nor U18406 (N_18406,N_18346,N_18356);
nor U18407 (N_18407,N_18203,N_18268);
nand U18408 (N_18408,N_18289,N_18215);
nor U18409 (N_18409,N_18399,N_18284);
and U18410 (N_18410,N_18364,N_18368);
nor U18411 (N_18411,N_18230,N_18285);
and U18412 (N_18412,N_18254,N_18282);
xor U18413 (N_18413,N_18232,N_18326);
and U18414 (N_18414,N_18267,N_18328);
and U18415 (N_18415,N_18351,N_18359);
xor U18416 (N_18416,N_18336,N_18358);
nor U18417 (N_18417,N_18286,N_18387);
and U18418 (N_18418,N_18288,N_18389);
nand U18419 (N_18419,N_18367,N_18247);
nor U18420 (N_18420,N_18227,N_18245);
xnor U18421 (N_18421,N_18325,N_18292);
and U18422 (N_18422,N_18372,N_18222);
xor U18423 (N_18423,N_18278,N_18272);
and U18424 (N_18424,N_18269,N_18250);
and U18425 (N_18425,N_18300,N_18397);
nand U18426 (N_18426,N_18264,N_18243);
nor U18427 (N_18427,N_18304,N_18213);
nand U18428 (N_18428,N_18378,N_18369);
nand U18429 (N_18429,N_18201,N_18307);
and U18430 (N_18430,N_18241,N_18331);
and U18431 (N_18431,N_18316,N_18355);
nor U18432 (N_18432,N_18248,N_18332);
nand U18433 (N_18433,N_18348,N_18321);
xnor U18434 (N_18434,N_18386,N_18382);
or U18435 (N_18435,N_18204,N_18370);
xor U18436 (N_18436,N_18212,N_18380);
or U18437 (N_18437,N_18329,N_18337);
or U18438 (N_18438,N_18236,N_18324);
xnor U18439 (N_18439,N_18216,N_18275);
nand U18440 (N_18440,N_18218,N_18357);
nor U18441 (N_18441,N_18327,N_18224);
or U18442 (N_18442,N_18223,N_18258);
xnor U18443 (N_18443,N_18373,N_18237);
nor U18444 (N_18444,N_18235,N_18277);
nand U18445 (N_18445,N_18392,N_18352);
and U18446 (N_18446,N_18394,N_18252);
xor U18447 (N_18447,N_18262,N_18260);
and U18448 (N_18448,N_18345,N_18225);
or U18449 (N_18449,N_18334,N_18293);
and U18450 (N_18450,N_18256,N_18266);
xnor U18451 (N_18451,N_18360,N_18362);
or U18452 (N_18452,N_18319,N_18383);
nor U18453 (N_18453,N_18276,N_18313);
and U18454 (N_18454,N_18390,N_18379);
or U18455 (N_18455,N_18296,N_18338);
nand U18456 (N_18456,N_18271,N_18315);
nor U18457 (N_18457,N_18287,N_18365);
nor U18458 (N_18458,N_18202,N_18283);
nor U18459 (N_18459,N_18312,N_18333);
nor U18460 (N_18460,N_18206,N_18349);
and U18461 (N_18461,N_18376,N_18305);
nand U18462 (N_18462,N_18261,N_18263);
and U18463 (N_18463,N_18375,N_18238);
xnor U18464 (N_18464,N_18253,N_18342);
nor U18465 (N_18465,N_18309,N_18233);
nor U18466 (N_18466,N_18294,N_18384);
nor U18467 (N_18467,N_18366,N_18371);
and U18468 (N_18468,N_18335,N_18255);
or U18469 (N_18469,N_18205,N_18207);
and U18470 (N_18470,N_18314,N_18317);
xor U18471 (N_18471,N_18299,N_18302);
nor U18472 (N_18472,N_18242,N_18303);
and U18473 (N_18473,N_18234,N_18320);
nor U18474 (N_18474,N_18214,N_18339);
and U18475 (N_18475,N_18310,N_18217);
nand U18476 (N_18476,N_18279,N_18340);
nand U18477 (N_18477,N_18374,N_18219);
xor U18478 (N_18478,N_18274,N_18398);
or U18479 (N_18479,N_18377,N_18251);
nand U18480 (N_18480,N_18270,N_18280);
or U18481 (N_18481,N_18343,N_18341);
nor U18482 (N_18482,N_18347,N_18388);
and U18483 (N_18483,N_18200,N_18259);
xor U18484 (N_18484,N_18396,N_18391);
nand U18485 (N_18485,N_18221,N_18228);
nor U18486 (N_18486,N_18385,N_18244);
nor U18487 (N_18487,N_18381,N_18344);
or U18488 (N_18488,N_18322,N_18350);
and U18489 (N_18489,N_18306,N_18354);
and U18490 (N_18490,N_18297,N_18301);
nand U18491 (N_18491,N_18298,N_18210);
nand U18492 (N_18492,N_18353,N_18311);
nand U18493 (N_18493,N_18246,N_18363);
xor U18494 (N_18494,N_18295,N_18281);
xor U18495 (N_18495,N_18290,N_18231);
and U18496 (N_18496,N_18257,N_18395);
nand U18497 (N_18497,N_18291,N_18226);
and U18498 (N_18498,N_18323,N_18240);
xor U18499 (N_18499,N_18273,N_18239);
nand U18500 (N_18500,N_18353,N_18346);
nand U18501 (N_18501,N_18336,N_18266);
and U18502 (N_18502,N_18340,N_18213);
and U18503 (N_18503,N_18336,N_18395);
xnor U18504 (N_18504,N_18230,N_18380);
or U18505 (N_18505,N_18241,N_18306);
nor U18506 (N_18506,N_18272,N_18252);
nand U18507 (N_18507,N_18347,N_18377);
nor U18508 (N_18508,N_18327,N_18386);
nand U18509 (N_18509,N_18258,N_18302);
or U18510 (N_18510,N_18345,N_18311);
xor U18511 (N_18511,N_18333,N_18316);
nand U18512 (N_18512,N_18288,N_18301);
or U18513 (N_18513,N_18298,N_18328);
nor U18514 (N_18514,N_18259,N_18331);
and U18515 (N_18515,N_18233,N_18273);
and U18516 (N_18516,N_18320,N_18342);
nor U18517 (N_18517,N_18398,N_18390);
or U18518 (N_18518,N_18212,N_18372);
nor U18519 (N_18519,N_18392,N_18327);
nor U18520 (N_18520,N_18294,N_18286);
or U18521 (N_18521,N_18336,N_18279);
nor U18522 (N_18522,N_18350,N_18319);
xnor U18523 (N_18523,N_18242,N_18306);
nor U18524 (N_18524,N_18333,N_18276);
or U18525 (N_18525,N_18210,N_18360);
nor U18526 (N_18526,N_18222,N_18360);
or U18527 (N_18527,N_18225,N_18236);
nor U18528 (N_18528,N_18280,N_18306);
nor U18529 (N_18529,N_18365,N_18379);
or U18530 (N_18530,N_18265,N_18212);
nor U18531 (N_18531,N_18329,N_18243);
nand U18532 (N_18532,N_18339,N_18231);
nor U18533 (N_18533,N_18365,N_18274);
nor U18534 (N_18534,N_18303,N_18323);
xnor U18535 (N_18535,N_18258,N_18209);
and U18536 (N_18536,N_18279,N_18231);
nand U18537 (N_18537,N_18280,N_18246);
or U18538 (N_18538,N_18264,N_18263);
xor U18539 (N_18539,N_18248,N_18362);
nor U18540 (N_18540,N_18313,N_18359);
nand U18541 (N_18541,N_18218,N_18362);
and U18542 (N_18542,N_18274,N_18313);
xor U18543 (N_18543,N_18269,N_18311);
xor U18544 (N_18544,N_18261,N_18266);
and U18545 (N_18545,N_18288,N_18385);
and U18546 (N_18546,N_18293,N_18259);
xor U18547 (N_18547,N_18211,N_18382);
xor U18548 (N_18548,N_18256,N_18281);
and U18549 (N_18549,N_18321,N_18200);
nor U18550 (N_18550,N_18311,N_18340);
xor U18551 (N_18551,N_18253,N_18371);
and U18552 (N_18552,N_18226,N_18311);
or U18553 (N_18553,N_18277,N_18273);
nor U18554 (N_18554,N_18284,N_18236);
nand U18555 (N_18555,N_18232,N_18222);
nor U18556 (N_18556,N_18260,N_18336);
or U18557 (N_18557,N_18276,N_18246);
xnor U18558 (N_18558,N_18351,N_18386);
or U18559 (N_18559,N_18319,N_18263);
nand U18560 (N_18560,N_18370,N_18284);
or U18561 (N_18561,N_18304,N_18238);
or U18562 (N_18562,N_18286,N_18232);
nand U18563 (N_18563,N_18314,N_18355);
xor U18564 (N_18564,N_18391,N_18264);
and U18565 (N_18565,N_18358,N_18225);
and U18566 (N_18566,N_18340,N_18328);
xnor U18567 (N_18567,N_18242,N_18228);
and U18568 (N_18568,N_18388,N_18247);
or U18569 (N_18569,N_18283,N_18226);
xnor U18570 (N_18570,N_18322,N_18333);
nand U18571 (N_18571,N_18287,N_18331);
nor U18572 (N_18572,N_18300,N_18381);
xor U18573 (N_18573,N_18220,N_18345);
or U18574 (N_18574,N_18349,N_18363);
nand U18575 (N_18575,N_18392,N_18318);
xnor U18576 (N_18576,N_18280,N_18315);
xnor U18577 (N_18577,N_18383,N_18354);
nor U18578 (N_18578,N_18337,N_18211);
xnor U18579 (N_18579,N_18353,N_18240);
or U18580 (N_18580,N_18356,N_18225);
xor U18581 (N_18581,N_18337,N_18261);
xnor U18582 (N_18582,N_18355,N_18397);
and U18583 (N_18583,N_18390,N_18297);
xor U18584 (N_18584,N_18305,N_18236);
xnor U18585 (N_18585,N_18208,N_18365);
nor U18586 (N_18586,N_18390,N_18334);
and U18587 (N_18587,N_18271,N_18200);
nor U18588 (N_18588,N_18370,N_18352);
and U18589 (N_18589,N_18207,N_18300);
nand U18590 (N_18590,N_18259,N_18332);
xor U18591 (N_18591,N_18294,N_18390);
xnor U18592 (N_18592,N_18342,N_18302);
and U18593 (N_18593,N_18245,N_18220);
nand U18594 (N_18594,N_18304,N_18326);
nor U18595 (N_18595,N_18245,N_18388);
and U18596 (N_18596,N_18355,N_18231);
xor U18597 (N_18597,N_18274,N_18322);
nor U18598 (N_18598,N_18399,N_18342);
nand U18599 (N_18599,N_18257,N_18204);
and U18600 (N_18600,N_18563,N_18496);
and U18601 (N_18601,N_18436,N_18495);
and U18602 (N_18602,N_18596,N_18407);
nand U18603 (N_18603,N_18548,N_18587);
nand U18604 (N_18604,N_18443,N_18557);
xor U18605 (N_18605,N_18498,N_18491);
and U18606 (N_18606,N_18466,N_18578);
xnor U18607 (N_18607,N_18489,N_18520);
and U18608 (N_18608,N_18431,N_18534);
xnor U18609 (N_18609,N_18475,N_18595);
nand U18610 (N_18610,N_18451,N_18525);
xnor U18611 (N_18611,N_18493,N_18552);
and U18612 (N_18612,N_18476,N_18486);
and U18613 (N_18613,N_18425,N_18459);
xnor U18614 (N_18614,N_18565,N_18598);
nor U18615 (N_18615,N_18411,N_18438);
nand U18616 (N_18616,N_18434,N_18429);
xnor U18617 (N_18617,N_18492,N_18577);
and U18618 (N_18618,N_18482,N_18424);
xnor U18619 (N_18619,N_18551,N_18437);
and U18620 (N_18620,N_18469,N_18535);
nand U18621 (N_18621,N_18541,N_18410);
or U18622 (N_18622,N_18441,N_18597);
nand U18623 (N_18623,N_18536,N_18470);
or U18624 (N_18624,N_18453,N_18522);
nor U18625 (N_18625,N_18422,N_18403);
nor U18626 (N_18626,N_18582,N_18572);
nor U18627 (N_18627,N_18526,N_18583);
and U18628 (N_18628,N_18550,N_18440);
and U18629 (N_18629,N_18544,N_18448);
nor U18630 (N_18630,N_18539,N_18442);
or U18631 (N_18631,N_18439,N_18400);
xor U18632 (N_18632,N_18527,N_18462);
xnor U18633 (N_18633,N_18432,N_18511);
or U18634 (N_18634,N_18545,N_18450);
nor U18635 (N_18635,N_18487,N_18404);
nand U18636 (N_18636,N_18455,N_18497);
nand U18637 (N_18637,N_18447,N_18558);
or U18638 (N_18638,N_18415,N_18433);
nand U18639 (N_18639,N_18519,N_18500);
nand U18640 (N_18640,N_18494,N_18481);
nor U18641 (N_18641,N_18428,N_18546);
nand U18642 (N_18642,N_18401,N_18584);
xor U18643 (N_18643,N_18559,N_18423);
nand U18644 (N_18644,N_18588,N_18514);
nor U18645 (N_18645,N_18521,N_18513);
xnor U18646 (N_18646,N_18484,N_18524);
xor U18647 (N_18647,N_18419,N_18561);
or U18648 (N_18648,N_18483,N_18599);
and U18649 (N_18649,N_18471,N_18567);
nand U18650 (N_18650,N_18594,N_18512);
xnor U18651 (N_18651,N_18532,N_18490);
nand U18652 (N_18652,N_18509,N_18414);
nor U18653 (N_18653,N_18538,N_18580);
nand U18654 (N_18654,N_18408,N_18454);
nand U18655 (N_18655,N_18473,N_18406);
nor U18656 (N_18656,N_18508,N_18555);
and U18657 (N_18657,N_18590,N_18474);
and U18658 (N_18658,N_18435,N_18554);
xnor U18659 (N_18659,N_18560,N_18488);
or U18660 (N_18660,N_18542,N_18571);
nand U18661 (N_18661,N_18477,N_18591);
or U18662 (N_18662,N_18518,N_18402);
nand U18663 (N_18663,N_18456,N_18515);
and U18664 (N_18664,N_18413,N_18416);
or U18665 (N_18665,N_18468,N_18576);
and U18666 (N_18666,N_18480,N_18505);
xor U18667 (N_18667,N_18446,N_18449);
and U18668 (N_18668,N_18517,N_18507);
or U18669 (N_18669,N_18549,N_18569);
nor U18670 (N_18670,N_18503,N_18537);
and U18671 (N_18671,N_18444,N_18501);
nor U18672 (N_18672,N_18523,N_18478);
nor U18673 (N_18673,N_18463,N_18516);
and U18674 (N_18674,N_18593,N_18543);
and U18675 (N_18675,N_18467,N_18530);
or U18676 (N_18676,N_18430,N_18573);
nand U18677 (N_18677,N_18540,N_18412);
xor U18678 (N_18678,N_18421,N_18409);
xnor U18679 (N_18679,N_18510,N_18592);
nor U18680 (N_18680,N_18585,N_18589);
xnor U18681 (N_18681,N_18445,N_18418);
and U18682 (N_18682,N_18458,N_18420);
nand U18683 (N_18683,N_18553,N_18547);
and U18684 (N_18684,N_18586,N_18427);
or U18685 (N_18685,N_18528,N_18457);
nand U18686 (N_18686,N_18504,N_18574);
or U18687 (N_18687,N_18566,N_18405);
nor U18688 (N_18688,N_18579,N_18499);
nor U18689 (N_18689,N_18564,N_18479);
or U18690 (N_18690,N_18570,N_18575);
or U18691 (N_18691,N_18417,N_18460);
nand U18692 (N_18692,N_18426,N_18506);
or U18693 (N_18693,N_18581,N_18531);
or U18694 (N_18694,N_18452,N_18502);
and U18695 (N_18695,N_18461,N_18464);
or U18696 (N_18696,N_18485,N_18562);
or U18697 (N_18697,N_18533,N_18465);
or U18698 (N_18698,N_18529,N_18556);
and U18699 (N_18699,N_18568,N_18472);
or U18700 (N_18700,N_18407,N_18524);
xnor U18701 (N_18701,N_18432,N_18507);
and U18702 (N_18702,N_18528,N_18446);
nand U18703 (N_18703,N_18573,N_18418);
nor U18704 (N_18704,N_18505,N_18431);
or U18705 (N_18705,N_18416,N_18578);
and U18706 (N_18706,N_18434,N_18471);
and U18707 (N_18707,N_18583,N_18589);
nor U18708 (N_18708,N_18400,N_18562);
or U18709 (N_18709,N_18587,N_18514);
nand U18710 (N_18710,N_18413,N_18504);
or U18711 (N_18711,N_18419,N_18421);
and U18712 (N_18712,N_18456,N_18442);
or U18713 (N_18713,N_18492,N_18581);
xnor U18714 (N_18714,N_18416,N_18550);
nand U18715 (N_18715,N_18490,N_18570);
and U18716 (N_18716,N_18527,N_18552);
or U18717 (N_18717,N_18443,N_18529);
xnor U18718 (N_18718,N_18550,N_18408);
nand U18719 (N_18719,N_18421,N_18466);
or U18720 (N_18720,N_18598,N_18593);
nand U18721 (N_18721,N_18429,N_18590);
nor U18722 (N_18722,N_18592,N_18449);
or U18723 (N_18723,N_18414,N_18523);
and U18724 (N_18724,N_18451,N_18435);
nor U18725 (N_18725,N_18406,N_18444);
xor U18726 (N_18726,N_18404,N_18564);
nand U18727 (N_18727,N_18563,N_18529);
xor U18728 (N_18728,N_18530,N_18536);
nor U18729 (N_18729,N_18497,N_18506);
or U18730 (N_18730,N_18444,N_18487);
and U18731 (N_18731,N_18505,N_18550);
and U18732 (N_18732,N_18552,N_18451);
or U18733 (N_18733,N_18484,N_18408);
nor U18734 (N_18734,N_18484,N_18435);
nand U18735 (N_18735,N_18465,N_18573);
xnor U18736 (N_18736,N_18493,N_18542);
nor U18737 (N_18737,N_18465,N_18586);
and U18738 (N_18738,N_18420,N_18558);
nor U18739 (N_18739,N_18425,N_18498);
or U18740 (N_18740,N_18518,N_18593);
xnor U18741 (N_18741,N_18410,N_18580);
and U18742 (N_18742,N_18534,N_18441);
nand U18743 (N_18743,N_18583,N_18500);
or U18744 (N_18744,N_18527,N_18477);
and U18745 (N_18745,N_18406,N_18407);
nand U18746 (N_18746,N_18451,N_18439);
and U18747 (N_18747,N_18504,N_18479);
nor U18748 (N_18748,N_18494,N_18528);
or U18749 (N_18749,N_18418,N_18521);
nand U18750 (N_18750,N_18456,N_18431);
or U18751 (N_18751,N_18522,N_18558);
xnor U18752 (N_18752,N_18425,N_18520);
nor U18753 (N_18753,N_18465,N_18482);
or U18754 (N_18754,N_18527,N_18555);
and U18755 (N_18755,N_18456,N_18418);
nand U18756 (N_18756,N_18495,N_18408);
nor U18757 (N_18757,N_18554,N_18585);
and U18758 (N_18758,N_18566,N_18520);
or U18759 (N_18759,N_18570,N_18523);
nand U18760 (N_18760,N_18511,N_18562);
nand U18761 (N_18761,N_18561,N_18500);
and U18762 (N_18762,N_18576,N_18432);
xnor U18763 (N_18763,N_18490,N_18544);
nand U18764 (N_18764,N_18496,N_18482);
or U18765 (N_18765,N_18559,N_18556);
nor U18766 (N_18766,N_18599,N_18448);
xnor U18767 (N_18767,N_18474,N_18557);
nand U18768 (N_18768,N_18537,N_18449);
nand U18769 (N_18769,N_18416,N_18465);
and U18770 (N_18770,N_18571,N_18457);
nor U18771 (N_18771,N_18573,N_18579);
nand U18772 (N_18772,N_18552,N_18440);
xor U18773 (N_18773,N_18418,N_18498);
and U18774 (N_18774,N_18400,N_18444);
nand U18775 (N_18775,N_18467,N_18501);
xnor U18776 (N_18776,N_18584,N_18572);
nor U18777 (N_18777,N_18436,N_18529);
xnor U18778 (N_18778,N_18529,N_18521);
or U18779 (N_18779,N_18448,N_18507);
nand U18780 (N_18780,N_18469,N_18501);
nand U18781 (N_18781,N_18405,N_18438);
nor U18782 (N_18782,N_18561,N_18567);
or U18783 (N_18783,N_18541,N_18459);
and U18784 (N_18784,N_18599,N_18574);
nor U18785 (N_18785,N_18468,N_18446);
or U18786 (N_18786,N_18592,N_18406);
and U18787 (N_18787,N_18520,N_18567);
or U18788 (N_18788,N_18529,N_18507);
xnor U18789 (N_18789,N_18416,N_18545);
xor U18790 (N_18790,N_18459,N_18536);
nor U18791 (N_18791,N_18417,N_18475);
xnor U18792 (N_18792,N_18454,N_18581);
nand U18793 (N_18793,N_18481,N_18433);
nor U18794 (N_18794,N_18407,N_18490);
xor U18795 (N_18795,N_18528,N_18487);
and U18796 (N_18796,N_18518,N_18458);
nand U18797 (N_18797,N_18424,N_18409);
nand U18798 (N_18798,N_18460,N_18554);
or U18799 (N_18799,N_18468,N_18598);
and U18800 (N_18800,N_18692,N_18746);
xor U18801 (N_18801,N_18650,N_18779);
xor U18802 (N_18802,N_18681,N_18720);
or U18803 (N_18803,N_18765,N_18639);
nand U18804 (N_18804,N_18687,N_18603);
and U18805 (N_18805,N_18641,N_18677);
nor U18806 (N_18806,N_18704,N_18792);
or U18807 (N_18807,N_18689,N_18742);
xor U18808 (N_18808,N_18736,N_18698);
nand U18809 (N_18809,N_18789,N_18732);
nor U18810 (N_18810,N_18691,N_18718);
and U18811 (N_18811,N_18622,N_18714);
xnor U18812 (N_18812,N_18662,N_18686);
or U18813 (N_18813,N_18702,N_18608);
xor U18814 (N_18814,N_18793,N_18672);
nor U18815 (N_18815,N_18657,N_18602);
xnor U18816 (N_18816,N_18629,N_18785);
xnor U18817 (N_18817,N_18607,N_18617);
xnor U18818 (N_18818,N_18798,N_18624);
and U18819 (N_18819,N_18740,N_18761);
or U18820 (N_18820,N_18620,N_18794);
nor U18821 (N_18821,N_18665,N_18751);
xnor U18822 (N_18822,N_18713,N_18621);
xnor U18823 (N_18823,N_18735,N_18690);
and U18824 (N_18824,N_18762,N_18684);
or U18825 (N_18825,N_18717,N_18786);
nand U18826 (N_18826,N_18769,N_18683);
and U18827 (N_18827,N_18707,N_18680);
and U18828 (N_18828,N_18634,N_18752);
or U18829 (N_18829,N_18640,N_18763);
or U18830 (N_18830,N_18754,N_18637);
nand U18831 (N_18831,N_18638,N_18749);
nor U18832 (N_18832,N_18695,N_18726);
nor U18833 (N_18833,N_18737,N_18618);
nor U18834 (N_18834,N_18758,N_18630);
and U18835 (N_18835,N_18612,N_18674);
or U18836 (N_18836,N_18780,N_18697);
xor U18837 (N_18837,N_18604,N_18666);
and U18838 (N_18838,N_18781,N_18659);
xor U18839 (N_18839,N_18649,N_18653);
xor U18840 (N_18840,N_18741,N_18635);
nor U18841 (N_18841,N_18727,N_18766);
and U18842 (N_18842,N_18772,N_18699);
and U18843 (N_18843,N_18631,N_18719);
nand U18844 (N_18844,N_18633,N_18611);
nand U18845 (N_18845,N_18623,N_18656);
and U18846 (N_18846,N_18605,N_18614);
nand U18847 (N_18847,N_18744,N_18663);
or U18848 (N_18848,N_18627,N_18642);
xor U18849 (N_18849,N_18722,N_18668);
and U18850 (N_18850,N_18700,N_18658);
and U18851 (N_18851,N_18628,N_18787);
nand U18852 (N_18852,N_18711,N_18784);
nand U18853 (N_18853,N_18788,N_18685);
xor U18854 (N_18854,N_18750,N_18679);
nor U18855 (N_18855,N_18748,N_18613);
and U18856 (N_18856,N_18701,N_18770);
nand U18857 (N_18857,N_18673,N_18790);
nor U18858 (N_18858,N_18670,N_18773);
and U18859 (N_18859,N_18644,N_18647);
xor U18860 (N_18860,N_18723,N_18799);
nand U18861 (N_18861,N_18768,N_18775);
and U18862 (N_18862,N_18706,N_18678);
and U18863 (N_18863,N_18708,N_18664);
and U18864 (N_18864,N_18716,N_18648);
or U18865 (N_18865,N_18676,N_18710);
xnor U18866 (N_18866,N_18636,N_18694);
or U18867 (N_18867,N_18777,N_18729);
or U18868 (N_18868,N_18767,N_18712);
nor U18869 (N_18869,N_18652,N_18625);
nor U18870 (N_18870,N_18733,N_18738);
or U18871 (N_18871,N_18693,N_18705);
xnor U18872 (N_18872,N_18646,N_18675);
or U18873 (N_18873,N_18771,N_18724);
nand U18874 (N_18874,N_18601,N_18776);
nand U18875 (N_18875,N_18669,N_18600);
nor U18876 (N_18876,N_18660,N_18759);
or U18877 (N_18877,N_18728,N_18651);
nand U18878 (N_18878,N_18721,N_18655);
or U18879 (N_18879,N_18696,N_18615);
nor U18880 (N_18880,N_18610,N_18626);
and U18881 (N_18881,N_18682,N_18760);
xnor U18882 (N_18882,N_18778,N_18730);
nand U18883 (N_18883,N_18725,N_18703);
or U18884 (N_18884,N_18606,N_18645);
nand U18885 (N_18885,N_18632,N_18796);
nor U18886 (N_18886,N_18709,N_18643);
or U18887 (N_18887,N_18619,N_18743);
nor U18888 (N_18888,N_18661,N_18671);
nor U18889 (N_18889,N_18774,N_18745);
xnor U18890 (N_18890,N_18791,N_18715);
xor U18891 (N_18891,N_18753,N_18757);
nor U18892 (N_18892,N_18667,N_18739);
nor U18893 (N_18893,N_18755,N_18783);
nor U18894 (N_18894,N_18688,N_18609);
or U18895 (N_18895,N_18756,N_18654);
nor U18896 (N_18896,N_18734,N_18795);
or U18897 (N_18897,N_18764,N_18616);
or U18898 (N_18898,N_18782,N_18731);
nand U18899 (N_18899,N_18797,N_18747);
nand U18900 (N_18900,N_18650,N_18749);
and U18901 (N_18901,N_18661,N_18726);
xnor U18902 (N_18902,N_18701,N_18729);
and U18903 (N_18903,N_18647,N_18779);
xnor U18904 (N_18904,N_18768,N_18788);
or U18905 (N_18905,N_18731,N_18684);
nor U18906 (N_18906,N_18658,N_18670);
nand U18907 (N_18907,N_18708,N_18600);
and U18908 (N_18908,N_18757,N_18747);
nand U18909 (N_18909,N_18624,N_18615);
or U18910 (N_18910,N_18716,N_18614);
or U18911 (N_18911,N_18782,N_18617);
nor U18912 (N_18912,N_18679,N_18608);
or U18913 (N_18913,N_18666,N_18681);
and U18914 (N_18914,N_18792,N_18630);
and U18915 (N_18915,N_18659,N_18650);
nor U18916 (N_18916,N_18688,N_18608);
and U18917 (N_18917,N_18798,N_18716);
nor U18918 (N_18918,N_18641,N_18794);
nor U18919 (N_18919,N_18780,N_18615);
nor U18920 (N_18920,N_18722,N_18784);
nand U18921 (N_18921,N_18714,N_18603);
nand U18922 (N_18922,N_18764,N_18797);
xnor U18923 (N_18923,N_18648,N_18605);
nor U18924 (N_18924,N_18743,N_18644);
or U18925 (N_18925,N_18709,N_18698);
and U18926 (N_18926,N_18718,N_18698);
and U18927 (N_18927,N_18740,N_18643);
nor U18928 (N_18928,N_18734,N_18694);
nor U18929 (N_18929,N_18646,N_18660);
nand U18930 (N_18930,N_18650,N_18637);
nor U18931 (N_18931,N_18791,N_18614);
nor U18932 (N_18932,N_18779,N_18626);
or U18933 (N_18933,N_18776,N_18635);
nand U18934 (N_18934,N_18612,N_18608);
nor U18935 (N_18935,N_18752,N_18646);
or U18936 (N_18936,N_18686,N_18741);
nor U18937 (N_18937,N_18707,N_18630);
or U18938 (N_18938,N_18663,N_18610);
and U18939 (N_18939,N_18611,N_18649);
and U18940 (N_18940,N_18790,N_18725);
and U18941 (N_18941,N_18768,N_18716);
or U18942 (N_18942,N_18789,N_18641);
xor U18943 (N_18943,N_18797,N_18761);
nor U18944 (N_18944,N_18760,N_18770);
xnor U18945 (N_18945,N_18734,N_18781);
or U18946 (N_18946,N_18769,N_18671);
or U18947 (N_18947,N_18655,N_18683);
or U18948 (N_18948,N_18621,N_18652);
xnor U18949 (N_18949,N_18752,N_18694);
nor U18950 (N_18950,N_18652,N_18764);
or U18951 (N_18951,N_18722,N_18734);
or U18952 (N_18952,N_18641,N_18705);
nand U18953 (N_18953,N_18767,N_18666);
nor U18954 (N_18954,N_18637,N_18649);
nor U18955 (N_18955,N_18724,N_18748);
nand U18956 (N_18956,N_18637,N_18628);
and U18957 (N_18957,N_18643,N_18678);
or U18958 (N_18958,N_18782,N_18712);
nor U18959 (N_18959,N_18736,N_18755);
and U18960 (N_18960,N_18787,N_18701);
nand U18961 (N_18961,N_18721,N_18600);
or U18962 (N_18962,N_18675,N_18691);
nor U18963 (N_18963,N_18742,N_18651);
and U18964 (N_18964,N_18759,N_18748);
nor U18965 (N_18965,N_18665,N_18606);
nand U18966 (N_18966,N_18651,N_18645);
or U18967 (N_18967,N_18685,N_18701);
nand U18968 (N_18968,N_18618,N_18747);
and U18969 (N_18969,N_18698,N_18795);
nor U18970 (N_18970,N_18725,N_18710);
nand U18971 (N_18971,N_18622,N_18607);
and U18972 (N_18972,N_18671,N_18746);
nand U18973 (N_18973,N_18649,N_18742);
and U18974 (N_18974,N_18682,N_18604);
xor U18975 (N_18975,N_18671,N_18721);
nor U18976 (N_18976,N_18794,N_18757);
xor U18977 (N_18977,N_18684,N_18788);
nor U18978 (N_18978,N_18721,N_18699);
xor U18979 (N_18979,N_18600,N_18740);
xnor U18980 (N_18980,N_18690,N_18760);
nor U18981 (N_18981,N_18798,N_18631);
xor U18982 (N_18982,N_18616,N_18657);
and U18983 (N_18983,N_18677,N_18614);
nand U18984 (N_18984,N_18761,N_18644);
and U18985 (N_18985,N_18649,N_18677);
or U18986 (N_18986,N_18601,N_18747);
nand U18987 (N_18987,N_18791,N_18736);
and U18988 (N_18988,N_18766,N_18759);
xor U18989 (N_18989,N_18650,N_18777);
and U18990 (N_18990,N_18754,N_18682);
nor U18991 (N_18991,N_18700,N_18686);
nor U18992 (N_18992,N_18630,N_18607);
or U18993 (N_18993,N_18614,N_18665);
or U18994 (N_18994,N_18611,N_18681);
xor U18995 (N_18995,N_18791,N_18690);
nand U18996 (N_18996,N_18723,N_18777);
xnor U18997 (N_18997,N_18727,N_18714);
nand U18998 (N_18998,N_18757,N_18779);
xnor U18999 (N_18999,N_18688,N_18763);
xnor U19000 (N_19000,N_18888,N_18806);
and U19001 (N_19001,N_18892,N_18854);
nand U19002 (N_19002,N_18984,N_18915);
nor U19003 (N_19003,N_18966,N_18909);
nor U19004 (N_19004,N_18846,N_18977);
nor U19005 (N_19005,N_18911,N_18994);
nand U19006 (N_19006,N_18919,N_18851);
and U19007 (N_19007,N_18906,N_18896);
or U19008 (N_19008,N_18813,N_18980);
xor U19009 (N_19009,N_18926,N_18927);
xor U19010 (N_19010,N_18916,N_18820);
nand U19011 (N_19011,N_18940,N_18997);
xor U19012 (N_19012,N_18925,N_18952);
or U19013 (N_19013,N_18941,N_18974);
xor U19014 (N_19014,N_18862,N_18898);
nor U19015 (N_19015,N_18955,N_18903);
nand U19016 (N_19016,N_18805,N_18876);
or U19017 (N_19017,N_18943,N_18938);
or U19018 (N_19018,N_18970,N_18928);
xnor U19019 (N_19019,N_18939,N_18870);
xor U19020 (N_19020,N_18991,N_18864);
xor U19021 (N_19021,N_18821,N_18914);
xor U19022 (N_19022,N_18924,N_18845);
and U19023 (N_19023,N_18954,N_18891);
nand U19024 (N_19024,N_18814,N_18887);
and U19025 (N_19025,N_18883,N_18899);
and U19026 (N_19026,N_18942,N_18834);
and U19027 (N_19027,N_18848,N_18957);
xnor U19028 (N_19028,N_18830,N_18872);
nor U19029 (N_19029,N_18843,N_18996);
nand U19030 (N_19030,N_18975,N_18958);
nand U19031 (N_19031,N_18929,N_18852);
xnor U19032 (N_19032,N_18871,N_18857);
nand U19033 (N_19033,N_18837,N_18890);
and U19034 (N_19034,N_18815,N_18930);
and U19035 (N_19035,N_18819,N_18983);
nor U19036 (N_19036,N_18986,N_18901);
nand U19037 (N_19037,N_18987,N_18858);
or U19038 (N_19038,N_18885,N_18880);
xnor U19039 (N_19039,N_18882,N_18913);
xnor U19040 (N_19040,N_18812,N_18921);
and U19041 (N_19041,N_18817,N_18900);
and U19042 (N_19042,N_18968,N_18842);
nand U19043 (N_19043,N_18973,N_18948);
xor U19044 (N_19044,N_18964,N_18895);
or U19045 (N_19045,N_18935,N_18945);
nor U19046 (N_19046,N_18985,N_18893);
or U19047 (N_19047,N_18875,N_18831);
and U19048 (N_19048,N_18801,N_18894);
and U19049 (N_19049,N_18979,N_18879);
or U19050 (N_19050,N_18931,N_18838);
xor U19051 (N_19051,N_18947,N_18804);
nor U19052 (N_19052,N_18972,N_18951);
nand U19053 (N_19053,N_18990,N_18839);
or U19054 (N_19054,N_18803,N_18978);
and U19055 (N_19055,N_18910,N_18937);
nor U19056 (N_19056,N_18855,N_18802);
nor U19057 (N_19057,N_18853,N_18999);
nand U19058 (N_19058,N_18841,N_18933);
nand U19059 (N_19059,N_18993,N_18998);
nor U19060 (N_19060,N_18823,N_18902);
xnor U19061 (N_19061,N_18917,N_18861);
or U19062 (N_19062,N_18967,N_18962);
nand U19063 (N_19063,N_18976,N_18950);
nor U19064 (N_19064,N_18856,N_18859);
and U19065 (N_19065,N_18992,N_18995);
or U19066 (N_19066,N_18877,N_18835);
or U19067 (N_19067,N_18811,N_18961);
nand U19068 (N_19068,N_18989,N_18869);
xnor U19069 (N_19069,N_18816,N_18953);
and U19070 (N_19070,N_18907,N_18822);
and U19071 (N_19071,N_18868,N_18826);
nand U19072 (N_19072,N_18918,N_18920);
nor U19073 (N_19073,N_18828,N_18897);
nor U19074 (N_19074,N_18827,N_18946);
nand U19075 (N_19075,N_18981,N_18922);
nand U19076 (N_19076,N_18889,N_18849);
xor U19077 (N_19077,N_18800,N_18836);
and U19078 (N_19078,N_18908,N_18960);
nor U19079 (N_19079,N_18884,N_18818);
and U19080 (N_19080,N_18833,N_18959);
and U19081 (N_19081,N_18944,N_18956);
and U19082 (N_19082,N_18904,N_18824);
and U19083 (N_19083,N_18982,N_18963);
or U19084 (N_19084,N_18832,N_18936);
nand U19085 (N_19085,N_18912,N_18844);
nor U19086 (N_19086,N_18807,N_18949);
nor U19087 (N_19087,N_18923,N_18825);
nor U19088 (N_19088,N_18810,N_18971);
and U19089 (N_19089,N_18969,N_18878);
or U19090 (N_19090,N_18829,N_18905);
or U19091 (N_19091,N_18934,N_18886);
nand U19092 (N_19092,N_18860,N_18873);
nor U19093 (N_19093,N_18867,N_18847);
or U19094 (N_19094,N_18988,N_18840);
nor U19095 (N_19095,N_18850,N_18881);
nor U19096 (N_19096,N_18863,N_18865);
or U19097 (N_19097,N_18809,N_18965);
nor U19098 (N_19098,N_18866,N_18874);
or U19099 (N_19099,N_18808,N_18932);
nand U19100 (N_19100,N_18955,N_18922);
xnor U19101 (N_19101,N_18971,N_18894);
nand U19102 (N_19102,N_18954,N_18877);
xor U19103 (N_19103,N_18880,N_18937);
nand U19104 (N_19104,N_18846,N_18854);
xnor U19105 (N_19105,N_18963,N_18841);
or U19106 (N_19106,N_18850,N_18973);
xor U19107 (N_19107,N_18835,N_18813);
and U19108 (N_19108,N_18934,N_18993);
and U19109 (N_19109,N_18923,N_18810);
xnor U19110 (N_19110,N_18963,N_18932);
and U19111 (N_19111,N_18818,N_18817);
nor U19112 (N_19112,N_18811,N_18850);
xor U19113 (N_19113,N_18905,N_18959);
xor U19114 (N_19114,N_18928,N_18964);
nor U19115 (N_19115,N_18921,N_18925);
nand U19116 (N_19116,N_18820,N_18926);
xnor U19117 (N_19117,N_18813,N_18987);
xor U19118 (N_19118,N_18971,N_18803);
nor U19119 (N_19119,N_18849,N_18832);
nand U19120 (N_19120,N_18852,N_18841);
xor U19121 (N_19121,N_18881,N_18948);
nand U19122 (N_19122,N_18826,N_18928);
or U19123 (N_19123,N_18836,N_18802);
and U19124 (N_19124,N_18816,N_18930);
and U19125 (N_19125,N_18996,N_18978);
and U19126 (N_19126,N_18940,N_18822);
and U19127 (N_19127,N_18919,N_18975);
nor U19128 (N_19128,N_18998,N_18989);
and U19129 (N_19129,N_18984,N_18861);
xnor U19130 (N_19130,N_18823,N_18930);
nand U19131 (N_19131,N_18936,N_18813);
and U19132 (N_19132,N_18967,N_18861);
xor U19133 (N_19133,N_18883,N_18848);
nor U19134 (N_19134,N_18867,N_18944);
xor U19135 (N_19135,N_18848,N_18939);
or U19136 (N_19136,N_18928,N_18914);
xnor U19137 (N_19137,N_18993,N_18897);
or U19138 (N_19138,N_18878,N_18894);
xor U19139 (N_19139,N_18978,N_18869);
nand U19140 (N_19140,N_18973,N_18879);
nor U19141 (N_19141,N_18978,N_18825);
nor U19142 (N_19142,N_18880,N_18928);
nor U19143 (N_19143,N_18976,N_18909);
nand U19144 (N_19144,N_18805,N_18917);
nand U19145 (N_19145,N_18887,N_18849);
and U19146 (N_19146,N_18826,N_18865);
and U19147 (N_19147,N_18896,N_18855);
nor U19148 (N_19148,N_18910,N_18988);
nor U19149 (N_19149,N_18866,N_18962);
or U19150 (N_19150,N_18976,N_18917);
nand U19151 (N_19151,N_18846,N_18802);
xor U19152 (N_19152,N_18986,N_18938);
or U19153 (N_19153,N_18884,N_18970);
and U19154 (N_19154,N_18885,N_18871);
xor U19155 (N_19155,N_18861,N_18882);
and U19156 (N_19156,N_18940,N_18907);
nor U19157 (N_19157,N_18835,N_18816);
xor U19158 (N_19158,N_18927,N_18969);
xor U19159 (N_19159,N_18879,N_18971);
and U19160 (N_19160,N_18824,N_18926);
and U19161 (N_19161,N_18855,N_18992);
nor U19162 (N_19162,N_18838,N_18993);
xor U19163 (N_19163,N_18852,N_18804);
or U19164 (N_19164,N_18888,N_18895);
xnor U19165 (N_19165,N_18875,N_18851);
xnor U19166 (N_19166,N_18926,N_18921);
nor U19167 (N_19167,N_18896,N_18904);
xnor U19168 (N_19168,N_18878,N_18873);
xnor U19169 (N_19169,N_18875,N_18973);
and U19170 (N_19170,N_18997,N_18972);
and U19171 (N_19171,N_18890,N_18908);
or U19172 (N_19172,N_18937,N_18986);
and U19173 (N_19173,N_18813,N_18848);
or U19174 (N_19174,N_18899,N_18978);
nand U19175 (N_19175,N_18885,N_18813);
xor U19176 (N_19176,N_18826,N_18946);
xor U19177 (N_19177,N_18919,N_18970);
xor U19178 (N_19178,N_18848,N_18997);
nand U19179 (N_19179,N_18813,N_18800);
or U19180 (N_19180,N_18895,N_18926);
xnor U19181 (N_19181,N_18857,N_18855);
nor U19182 (N_19182,N_18931,N_18924);
and U19183 (N_19183,N_18871,N_18856);
nor U19184 (N_19184,N_18915,N_18886);
or U19185 (N_19185,N_18891,N_18899);
nor U19186 (N_19186,N_18901,N_18908);
and U19187 (N_19187,N_18953,N_18841);
xor U19188 (N_19188,N_18854,N_18988);
and U19189 (N_19189,N_18982,N_18955);
and U19190 (N_19190,N_18870,N_18948);
xor U19191 (N_19191,N_18877,N_18846);
and U19192 (N_19192,N_18887,N_18913);
nand U19193 (N_19193,N_18840,N_18815);
and U19194 (N_19194,N_18984,N_18996);
or U19195 (N_19195,N_18984,N_18928);
xor U19196 (N_19196,N_18930,N_18900);
or U19197 (N_19197,N_18941,N_18885);
nand U19198 (N_19198,N_18901,N_18873);
and U19199 (N_19199,N_18994,N_18851);
or U19200 (N_19200,N_19047,N_19195);
or U19201 (N_19201,N_19171,N_19057);
nand U19202 (N_19202,N_19070,N_19050);
xnor U19203 (N_19203,N_19083,N_19187);
xnor U19204 (N_19204,N_19006,N_19080);
nor U19205 (N_19205,N_19129,N_19052);
and U19206 (N_19206,N_19003,N_19102);
nand U19207 (N_19207,N_19156,N_19071);
and U19208 (N_19208,N_19024,N_19114);
or U19209 (N_19209,N_19142,N_19173);
xnor U19210 (N_19210,N_19038,N_19026);
xnor U19211 (N_19211,N_19113,N_19034);
and U19212 (N_19212,N_19064,N_19176);
or U19213 (N_19213,N_19163,N_19108);
xnor U19214 (N_19214,N_19067,N_19196);
or U19215 (N_19215,N_19058,N_19051);
nor U19216 (N_19216,N_19030,N_19045);
or U19217 (N_19217,N_19007,N_19144);
xor U19218 (N_19218,N_19110,N_19090);
nand U19219 (N_19219,N_19043,N_19012);
nor U19220 (N_19220,N_19033,N_19086);
and U19221 (N_19221,N_19094,N_19005);
and U19222 (N_19222,N_19008,N_19096);
nand U19223 (N_19223,N_19170,N_19032);
xnor U19224 (N_19224,N_19097,N_19158);
and U19225 (N_19225,N_19085,N_19036);
or U19226 (N_19226,N_19035,N_19157);
nor U19227 (N_19227,N_19040,N_19133);
xnor U19228 (N_19228,N_19134,N_19117);
and U19229 (N_19229,N_19078,N_19151);
or U19230 (N_19230,N_19153,N_19087);
nand U19231 (N_19231,N_19135,N_19081);
and U19232 (N_19232,N_19009,N_19194);
nand U19233 (N_19233,N_19186,N_19073);
and U19234 (N_19234,N_19139,N_19075);
or U19235 (N_19235,N_19140,N_19178);
xor U19236 (N_19236,N_19168,N_19189);
xor U19237 (N_19237,N_19041,N_19183);
or U19238 (N_19238,N_19104,N_19002);
xnor U19239 (N_19239,N_19084,N_19031);
or U19240 (N_19240,N_19105,N_19018);
xnor U19241 (N_19241,N_19164,N_19021);
xor U19242 (N_19242,N_19175,N_19120);
xnor U19243 (N_19243,N_19112,N_19049);
nor U19244 (N_19244,N_19020,N_19025);
nor U19245 (N_19245,N_19115,N_19082);
nor U19246 (N_19246,N_19028,N_19180);
xor U19247 (N_19247,N_19065,N_19132);
xnor U19248 (N_19248,N_19055,N_19068);
or U19249 (N_19249,N_19143,N_19023);
and U19250 (N_19250,N_19056,N_19042);
xnor U19251 (N_19251,N_19010,N_19019);
or U19252 (N_19252,N_19066,N_19193);
or U19253 (N_19253,N_19107,N_19063);
nor U19254 (N_19254,N_19177,N_19017);
nand U19255 (N_19255,N_19122,N_19123);
or U19256 (N_19256,N_19093,N_19188);
nor U19257 (N_19257,N_19076,N_19014);
xor U19258 (N_19258,N_19152,N_19013);
and U19259 (N_19259,N_19167,N_19111);
xnor U19260 (N_19260,N_19191,N_19100);
xnor U19261 (N_19261,N_19146,N_19150);
xor U19262 (N_19262,N_19099,N_19062);
nand U19263 (N_19263,N_19181,N_19190);
and U19264 (N_19264,N_19128,N_19118);
nand U19265 (N_19265,N_19103,N_19127);
or U19266 (N_19266,N_19079,N_19141);
xor U19267 (N_19267,N_19027,N_19131);
xor U19268 (N_19268,N_19145,N_19199);
or U19269 (N_19269,N_19088,N_19121);
xor U19270 (N_19270,N_19054,N_19148);
xnor U19271 (N_19271,N_19048,N_19172);
nor U19272 (N_19272,N_19072,N_19037);
or U19273 (N_19273,N_19197,N_19106);
nand U19274 (N_19274,N_19069,N_19059);
nand U19275 (N_19275,N_19162,N_19001);
nor U19276 (N_19276,N_19169,N_19077);
nor U19277 (N_19277,N_19179,N_19182);
nand U19278 (N_19278,N_19126,N_19044);
nand U19279 (N_19279,N_19125,N_19109);
and U19280 (N_19280,N_19060,N_19000);
and U19281 (N_19281,N_19119,N_19095);
nand U19282 (N_19282,N_19136,N_19101);
nor U19283 (N_19283,N_19161,N_19130);
and U19284 (N_19284,N_19098,N_19004);
xnor U19285 (N_19285,N_19022,N_19185);
and U19286 (N_19286,N_19053,N_19016);
or U19287 (N_19287,N_19149,N_19147);
nor U19288 (N_19288,N_19046,N_19159);
or U19289 (N_19289,N_19091,N_19174);
xor U19290 (N_19290,N_19137,N_19011);
nand U19291 (N_19291,N_19154,N_19092);
nor U19292 (N_19292,N_19039,N_19089);
xor U19293 (N_19293,N_19160,N_19192);
nand U19294 (N_19294,N_19124,N_19184);
and U19295 (N_19295,N_19138,N_19061);
xor U19296 (N_19296,N_19029,N_19155);
and U19297 (N_19297,N_19015,N_19116);
xor U19298 (N_19298,N_19074,N_19166);
nor U19299 (N_19299,N_19165,N_19198);
nand U19300 (N_19300,N_19149,N_19067);
and U19301 (N_19301,N_19055,N_19062);
or U19302 (N_19302,N_19003,N_19015);
nand U19303 (N_19303,N_19071,N_19038);
nor U19304 (N_19304,N_19039,N_19085);
xor U19305 (N_19305,N_19066,N_19005);
and U19306 (N_19306,N_19055,N_19142);
nor U19307 (N_19307,N_19081,N_19075);
xor U19308 (N_19308,N_19086,N_19028);
nand U19309 (N_19309,N_19033,N_19197);
xor U19310 (N_19310,N_19047,N_19050);
or U19311 (N_19311,N_19073,N_19065);
xor U19312 (N_19312,N_19079,N_19051);
nand U19313 (N_19313,N_19077,N_19000);
xor U19314 (N_19314,N_19176,N_19061);
nand U19315 (N_19315,N_19060,N_19016);
xor U19316 (N_19316,N_19187,N_19144);
or U19317 (N_19317,N_19145,N_19068);
xnor U19318 (N_19318,N_19110,N_19199);
nor U19319 (N_19319,N_19007,N_19185);
or U19320 (N_19320,N_19045,N_19144);
or U19321 (N_19321,N_19013,N_19023);
nand U19322 (N_19322,N_19192,N_19010);
nor U19323 (N_19323,N_19019,N_19139);
or U19324 (N_19324,N_19040,N_19026);
or U19325 (N_19325,N_19095,N_19003);
xnor U19326 (N_19326,N_19099,N_19006);
and U19327 (N_19327,N_19098,N_19173);
nor U19328 (N_19328,N_19156,N_19023);
nand U19329 (N_19329,N_19059,N_19171);
nand U19330 (N_19330,N_19049,N_19177);
nor U19331 (N_19331,N_19144,N_19073);
nand U19332 (N_19332,N_19156,N_19151);
nand U19333 (N_19333,N_19073,N_19012);
nor U19334 (N_19334,N_19151,N_19003);
and U19335 (N_19335,N_19080,N_19007);
and U19336 (N_19336,N_19156,N_19078);
nor U19337 (N_19337,N_19108,N_19082);
xor U19338 (N_19338,N_19044,N_19114);
nand U19339 (N_19339,N_19000,N_19120);
or U19340 (N_19340,N_19113,N_19092);
and U19341 (N_19341,N_19030,N_19155);
and U19342 (N_19342,N_19113,N_19150);
and U19343 (N_19343,N_19096,N_19140);
nor U19344 (N_19344,N_19003,N_19160);
xor U19345 (N_19345,N_19086,N_19017);
nand U19346 (N_19346,N_19122,N_19128);
nor U19347 (N_19347,N_19128,N_19059);
and U19348 (N_19348,N_19183,N_19126);
nand U19349 (N_19349,N_19181,N_19012);
or U19350 (N_19350,N_19000,N_19063);
nand U19351 (N_19351,N_19127,N_19117);
nor U19352 (N_19352,N_19100,N_19023);
nor U19353 (N_19353,N_19064,N_19155);
nand U19354 (N_19354,N_19107,N_19194);
and U19355 (N_19355,N_19018,N_19162);
nand U19356 (N_19356,N_19164,N_19062);
nand U19357 (N_19357,N_19186,N_19113);
xnor U19358 (N_19358,N_19060,N_19046);
nand U19359 (N_19359,N_19055,N_19164);
and U19360 (N_19360,N_19011,N_19199);
xor U19361 (N_19361,N_19095,N_19025);
and U19362 (N_19362,N_19030,N_19031);
xor U19363 (N_19363,N_19082,N_19093);
xnor U19364 (N_19364,N_19129,N_19060);
nor U19365 (N_19365,N_19179,N_19170);
xor U19366 (N_19366,N_19180,N_19086);
nand U19367 (N_19367,N_19004,N_19034);
xor U19368 (N_19368,N_19096,N_19110);
xnor U19369 (N_19369,N_19041,N_19042);
xnor U19370 (N_19370,N_19149,N_19001);
xnor U19371 (N_19371,N_19062,N_19103);
nand U19372 (N_19372,N_19160,N_19095);
nand U19373 (N_19373,N_19133,N_19191);
nor U19374 (N_19374,N_19173,N_19189);
xor U19375 (N_19375,N_19001,N_19007);
and U19376 (N_19376,N_19010,N_19117);
xor U19377 (N_19377,N_19054,N_19087);
nand U19378 (N_19378,N_19057,N_19059);
xor U19379 (N_19379,N_19072,N_19193);
nor U19380 (N_19380,N_19173,N_19038);
or U19381 (N_19381,N_19049,N_19024);
nor U19382 (N_19382,N_19156,N_19065);
nand U19383 (N_19383,N_19134,N_19080);
nand U19384 (N_19384,N_19142,N_19004);
and U19385 (N_19385,N_19078,N_19081);
nand U19386 (N_19386,N_19051,N_19140);
or U19387 (N_19387,N_19175,N_19010);
nand U19388 (N_19388,N_19006,N_19141);
nand U19389 (N_19389,N_19043,N_19109);
xor U19390 (N_19390,N_19158,N_19095);
and U19391 (N_19391,N_19182,N_19133);
nor U19392 (N_19392,N_19045,N_19021);
or U19393 (N_19393,N_19169,N_19018);
or U19394 (N_19394,N_19056,N_19139);
nand U19395 (N_19395,N_19160,N_19117);
xnor U19396 (N_19396,N_19129,N_19018);
and U19397 (N_19397,N_19116,N_19131);
or U19398 (N_19398,N_19036,N_19003);
xor U19399 (N_19399,N_19117,N_19189);
nand U19400 (N_19400,N_19350,N_19229);
xor U19401 (N_19401,N_19363,N_19394);
nor U19402 (N_19402,N_19273,N_19348);
nand U19403 (N_19403,N_19380,N_19296);
xor U19404 (N_19404,N_19376,N_19366);
and U19405 (N_19405,N_19212,N_19244);
nor U19406 (N_19406,N_19237,N_19333);
nor U19407 (N_19407,N_19369,N_19241);
nand U19408 (N_19408,N_19365,N_19374);
or U19409 (N_19409,N_19291,N_19217);
nor U19410 (N_19410,N_19269,N_19274);
xor U19411 (N_19411,N_19377,N_19253);
xnor U19412 (N_19412,N_19246,N_19283);
or U19413 (N_19413,N_19250,N_19387);
nand U19414 (N_19414,N_19265,N_19251);
or U19415 (N_19415,N_19203,N_19230);
and U19416 (N_19416,N_19359,N_19316);
or U19417 (N_19417,N_19208,N_19224);
or U19418 (N_19418,N_19351,N_19354);
nand U19419 (N_19419,N_19367,N_19298);
or U19420 (N_19420,N_19293,N_19297);
nor U19421 (N_19421,N_19397,N_19344);
nand U19422 (N_19422,N_19356,N_19288);
nand U19423 (N_19423,N_19308,N_19232);
or U19424 (N_19424,N_19370,N_19318);
xnor U19425 (N_19425,N_19225,N_19384);
xor U19426 (N_19426,N_19242,N_19341);
nand U19427 (N_19427,N_19227,N_19235);
nor U19428 (N_19428,N_19202,N_19236);
xnor U19429 (N_19429,N_19313,N_19393);
xor U19430 (N_19430,N_19254,N_19275);
xnor U19431 (N_19431,N_19259,N_19331);
nand U19432 (N_19432,N_19292,N_19210);
and U19433 (N_19433,N_19271,N_19299);
or U19434 (N_19434,N_19379,N_19270);
nor U19435 (N_19435,N_19392,N_19205);
or U19436 (N_19436,N_19383,N_19303);
nand U19437 (N_19437,N_19305,N_19262);
nor U19438 (N_19438,N_19226,N_19304);
nand U19439 (N_19439,N_19260,N_19228);
nor U19440 (N_19440,N_19249,N_19219);
nor U19441 (N_19441,N_19314,N_19239);
or U19442 (N_19442,N_19209,N_19216);
nor U19443 (N_19443,N_19223,N_19207);
and U19444 (N_19444,N_19362,N_19222);
or U19445 (N_19445,N_19231,N_19214);
and U19446 (N_19446,N_19256,N_19211);
xor U19447 (N_19447,N_19263,N_19347);
nor U19448 (N_19448,N_19302,N_19276);
nor U19449 (N_19449,N_19220,N_19311);
and U19450 (N_19450,N_19278,N_19391);
nand U19451 (N_19451,N_19364,N_19357);
and U19452 (N_19452,N_19353,N_19307);
xnor U19453 (N_19453,N_19372,N_19201);
and U19454 (N_19454,N_19346,N_19215);
or U19455 (N_19455,N_19355,N_19280);
and U19456 (N_19456,N_19324,N_19310);
and U19457 (N_19457,N_19396,N_19248);
xnor U19458 (N_19458,N_19309,N_19300);
and U19459 (N_19459,N_19252,N_19336);
nand U19460 (N_19460,N_19319,N_19247);
or U19461 (N_19461,N_19358,N_19334);
and U19462 (N_19462,N_19321,N_19345);
nand U19463 (N_19463,N_19294,N_19378);
or U19464 (N_19464,N_19389,N_19323);
or U19465 (N_19465,N_19390,N_19386);
nand U19466 (N_19466,N_19206,N_19281);
nand U19467 (N_19467,N_19385,N_19330);
xnor U19468 (N_19468,N_19267,N_19261);
nor U19469 (N_19469,N_19282,N_19315);
nor U19470 (N_19470,N_19360,N_19257);
or U19471 (N_19471,N_19221,N_19327);
nor U19472 (N_19472,N_19238,N_19340);
or U19473 (N_19473,N_19375,N_19290);
nand U19474 (N_19474,N_19200,N_19258);
nor U19475 (N_19475,N_19343,N_19325);
xor U19476 (N_19476,N_19233,N_19285);
or U19477 (N_19477,N_19255,N_19213);
or U19478 (N_19478,N_19399,N_19240);
nand U19479 (N_19479,N_19301,N_19349);
and U19480 (N_19480,N_19245,N_19320);
or U19481 (N_19481,N_19371,N_19289);
and U19482 (N_19482,N_19398,N_19266);
nor U19483 (N_19483,N_19368,N_19326);
xnor U19484 (N_19484,N_19279,N_19317);
or U19485 (N_19485,N_19395,N_19352);
and U19486 (N_19486,N_19204,N_19268);
xnor U19487 (N_19487,N_19342,N_19337);
or U19488 (N_19488,N_19361,N_19306);
and U19489 (N_19489,N_19329,N_19287);
or U19490 (N_19490,N_19338,N_19322);
or U19491 (N_19491,N_19388,N_19286);
nor U19492 (N_19492,N_19234,N_19264);
xnor U19493 (N_19493,N_19328,N_19243);
nor U19494 (N_19494,N_19295,N_19335);
or U19495 (N_19495,N_19272,N_19277);
xor U19496 (N_19496,N_19381,N_19218);
nand U19497 (N_19497,N_19332,N_19284);
nor U19498 (N_19498,N_19339,N_19312);
xor U19499 (N_19499,N_19373,N_19382);
xnor U19500 (N_19500,N_19314,N_19299);
nor U19501 (N_19501,N_19395,N_19285);
or U19502 (N_19502,N_19233,N_19320);
nand U19503 (N_19503,N_19385,N_19203);
nand U19504 (N_19504,N_19349,N_19316);
and U19505 (N_19505,N_19393,N_19263);
or U19506 (N_19506,N_19217,N_19227);
and U19507 (N_19507,N_19353,N_19329);
xor U19508 (N_19508,N_19366,N_19201);
nor U19509 (N_19509,N_19377,N_19240);
nand U19510 (N_19510,N_19332,N_19369);
xor U19511 (N_19511,N_19298,N_19335);
and U19512 (N_19512,N_19341,N_19380);
nand U19513 (N_19513,N_19203,N_19206);
and U19514 (N_19514,N_19362,N_19293);
nor U19515 (N_19515,N_19281,N_19392);
xnor U19516 (N_19516,N_19345,N_19398);
nand U19517 (N_19517,N_19366,N_19299);
or U19518 (N_19518,N_19245,N_19282);
nor U19519 (N_19519,N_19328,N_19209);
nor U19520 (N_19520,N_19304,N_19225);
xor U19521 (N_19521,N_19234,N_19299);
nor U19522 (N_19522,N_19314,N_19238);
nor U19523 (N_19523,N_19315,N_19252);
or U19524 (N_19524,N_19318,N_19344);
or U19525 (N_19525,N_19375,N_19232);
and U19526 (N_19526,N_19244,N_19329);
nand U19527 (N_19527,N_19372,N_19287);
xnor U19528 (N_19528,N_19341,N_19226);
or U19529 (N_19529,N_19267,N_19214);
or U19530 (N_19530,N_19214,N_19301);
and U19531 (N_19531,N_19373,N_19372);
nor U19532 (N_19532,N_19248,N_19233);
nand U19533 (N_19533,N_19215,N_19246);
nor U19534 (N_19534,N_19237,N_19319);
and U19535 (N_19535,N_19320,N_19259);
nand U19536 (N_19536,N_19344,N_19231);
or U19537 (N_19537,N_19307,N_19343);
xnor U19538 (N_19538,N_19280,N_19266);
xor U19539 (N_19539,N_19307,N_19351);
xor U19540 (N_19540,N_19329,N_19342);
and U19541 (N_19541,N_19332,N_19365);
nand U19542 (N_19542,N_19370,N_19367);
xor U19543 (N_19543,N_19395,N_19253);
or U19544 (N_19544,N_19267,N_19266);
and U19545 (N_19545,N_19263,N_19326);
xnor U19546 (N_19546,N_19366,N_19214);
xnor U19547 (N_19547,N_19253,N_19273);
or U19548 (N_19548,N_19336,N_19235);
and U19549 (N_19549,N_19371,N_19297);
or U19550 (N_19550,N_19376,N_19302);
nand U19551 (N_19551,N_19308,N_19310);
and U19552 (N_19552,N_19335,N_19222);
or U19553 (N_19553,N_19330,N_19200);
xor U19554 (N_19554,N_19268,N_19350);
or U19555 (N_19555,N_19217,N_19290);
nand U19556 (N_19556,N_19301,N_19286);
or U19557 (N_19557,N_19370,N_19271);
nand U19558 (N_19558,N_19365,N_19317);
xnor U19559 (N_19559,N_19215,N_19287);
xnor U19560 (N_19560,N_19278,N_19242);
nand U19561 (N_19561,N_19392,N_19239);
and U19562 (N_19562,N_19203,N_19340);
xnor U19563 (N_19563,N_19338,N_19298);
nand U19564 (N_19564,N_19288,N_19234);
nor U19565 (N_19565,N_19302,N_19213);
and U19566 (N_19566,N_19272,N_19206);
nand U19567 (N_19567,N_19257,N_19326);
or U19568 (N_19568,N_19258,N_19396);
nand U19569 (N_19569,N_19205,N_19271);
xnor U19570 (N_19570,N_19240,N_19266);
nand U19571 (N_19571,N_19302,N_19255);
xnor U19572 (N_19572,N_19349,N_19302);
and U19573 (N_19573,N_19231,N_19392);
or U19574 (N_19574,N_19269,N_19344);
or U19575 (N_19575,N_19380,N_19265);
and U19576 (N_19576,N_19372,N_19204);
nand U19577 (N_19577,N_19291,N_19243);
and U19578 (N_19578,N_19211,N_19263);
or U19579 (N_19579,N_19366,N_19320);
xor U19580 (N_19580,N_19389,N_19305);
or U19581 (N_19581,N_19251,N_19354);
xnor U19582 (N_19582,N_19234,N_19208);
or U19583 (N_19583,N_19283,N_19388);
and U19584 (N_19584,N_19261,N_19383);
and U19585 (N_19585,N_19342,N_19206);
xnor U19586 (N_19586,N_19321,N_19262);
and U19587 (N_19587,N_19364,N_19283);
or U19588 (N_19588,N_19255,N_19393);
and U19589 (N_19589,N_19283,N_19267);
and U19590 (N_19590,N_19316,N_19340);
or U19591 (N_19591,N_19287,N_19259);
nor U19592 (N_19592,N_19316,N_19233);
nor U19593 (N_19593,N_19296,N_19348);
and U19594 (N_19594,N_19273,N_19395);
xnor U19595 (N_19595,N_19223,N_19348);
or U19596 (N_19596,N_19357,N_19250);
nand U19597 (N_19597,N_19321,N_19236);
or U19598 (N_19598,N_19292,N_19352);
nor U19599 (N_19599,N_19342,N_19373);
and U19600 (N_19600,N_19502,N_19493);
nor U19601 (N_19601,N_19437,N_19562);
xor U19602 (N_19602,N_19411,N_19584);
and U19603 (N_19603,N_19540,N_19499);
nor U19604 (N_19604,N_19462,N_19429);
nor U19605 (N_19605,N_19569,N_19466);
xor U19606 (N_19606,N_19432,N_19537);
nand U19607 (N_19607,N_19505,N_19443);
nor U19608 (N_19608,N_19550,N_19450);
nor U19609 (N_19609,N_19551,N_19401);
and U19610 (N_19610,N_19589,N_19406);
and U19611 (N_19611,N_19568,N_19439);
nand U19612 (N_19612,N_19488,N_19442);
or U19613 (N_19613,N_19496,N_19507);
nor U19614 (N_19614,N_19572,N_19487);
nor U19615 (N_19615,N_19449,N_19420);
xor U19616 (N_19616,N_19517,N_19549);
and U19617 (N_19617,N_19417,N_19409);
or U19618 (N_19618,N_19457,N_19486);
and U19619 (N_19619,N_19510,N_19580);
xor U19620 (N_19620,N_19599,N_19467);
nor U19621 (N_19621,N_19552,N_19460);
and U19622 (N_19622,N_19593,N_19404);
xor U19623 (N_19623,N_19577,N_19465);
nand U19624 (N_19624,N_19490,N_19590);
xnor U19625 (N_19625,N_19500,N_19533);
nor U19626 (N_19626,N_19515,N_19554);
xor U19627 (N_19627,N_19452,N_19513);
nor U19628 (N_19628,N_19415,N_19514);
or U19629 (N_19629,N_19586,N_19545);
and U19630 (N_19630,N_19553,N_19476);
nor U19631 (N_19631,N_19530,N_19436);
nor U19632 (N_19632,N_19451,N_19543);
or U19633 (N_19633,N_19475,N_19403);
nor U19634 (N_19634,N_19596,N_19573);
xnor U19635 (N_19635,N_19509,N_19520);
xor U19636 (N_19636,N_19532,N_19419);
xor U19637 (N_19637,N_19592,N_19548);
xor U19638 (N_19638,N_19542,N_19574);
or U19639 (N_19639,N_19434,N_19501);
nand U19640 (N_19640,N_19561,N_19423);
nor U19641 (N_19641,N_19564,N_19508);
nand U19642 (N_19642,N_19494,N_19511);
or U19643 (N_19643,N_19512,N_19595);
or U19644 (N_19644,N_19425,N_19481);
nand U19645 (N_19645,N_19570,N_19519);
nor U19646 (N_19646,N_19521,N_19414);
and U19647 (N_19647,N_19472,N_19497);
xnor U19648 (N_19648,N_19474,N_19407);
xnor U19649 (N_19649,N_19527,N_19485);
nor U19650 (N_19650,N_19518,N_19525);
or U19651 (N_19651,N_19453,N_19558);
and U19652 (N_19652,N_19422,N_19428);
xnor U19653 (N_19653,N_19463,N_19426);
xor U19654 (N_19654,N_19412,N_19479);
nor U19655 (N_19655,N_19544,N_19546);
or U19656 (N_19656,N_19456,N_19566);
and U19657 (N_19657,N_19563,N_19455);
xnor U19658 (N_19658,N_19498,N_19582);
nor U19659 (N_19659,N_19579,N_19459);
nor U19660 (N_19660,N_19531,N_19441);
or U19661 (N_19661,N_19516,N_19492);
xor U19662 (N_19662,N_19597,N_19478);
xnor U19663 (N_19663,N_19424,N_19405);
and U19664 (N_19664,N_19576,N_19468);
xor U19665 (N_19665,N_19433,N_19524);
nand U19666 (N_19666,N_19484,N_19440);
and U19667 (N_19667,N_19565,N_19473);
or U19668 (N_19668,N_19464,N_19445);
or U19669 (N_19669,N_19523,N_19557);
nand U19670 (N_19670,N_19400,N_19482);
nor U19671 (N_19671,N_19461,N_19491);
and U19672 (N_19672,N_19402,N_19416);
nor U19673 (N_19673,N_19526,N_19454);
or U19674 (N_19674,N_19534,N_19421);
or U19675 (N_19675,N_19470,N_19547);
nand U19676 (N_19676,N_19581,N_19435);
or U19677 (N_19677,N_19431,N_19591);
and U19678 (N_19678,N_19418,N_19560);
xnor U19679 (N_19679,N_19413,N_19598);
nand U19680 (N_19680,N_19458,N_19444);
xor U19681 (N_19681,N_19448,N_19559);
xor U19682 (N_19682,N_19471,N_19556);
nand U19683 (N_19683,N_19588,N_19541);
xnor U19684 (N_19684,N_19483,N_19585);
xor U19685 (N_19685,N_19587,N_19410);
nand U19686 (N_19686,N_19430,N_19535);
and U19687 (N_19687,N_19495,N_19446);
nor U19688 (N_19688,N_19555,N_19536);
nand U19689 (N_19689,N_19427,N_19438);
nand U19690 (N_19690,N_19539,N_19529);
nand U19691 (N_19691,N_19594,N_19503);
or U19692 (N_19692,N_19583,N_19528);
or U19693 (N_19693,N_19567,N_19408);
and U19694 (N_19694,N_19480,N_19575);
xnor U19695 (N_19695,N_19447,N_19504);
nor U19696 (N_19696,N_19469,N_19571);
or U19697 (N_19697,N_19538,N_19477);
or U19698 (N_19698,N_19578,N_19506);
nor U19699 (N_19699,N_19522,N_19489);
xnor U19700 (N_19700,N_19536,N_19578);
and U19701 (N_19701,N_19511,N_19447);
nor U19702 (N_19702,N_19522,N_19408);
or U19703 (N_19703,N_19458,N_19519);
xnor U19704 (N_19704,N_19430,N_19457);
and U19705 (N_19705,N_19554,N_19564);
nand U19706 (N_19706,N_19444,N_19536);
nor U19707 (N_19707,N_19582,N_19423);
xor U19708 (N_19708,N_19416,N_19572);
xnor U19709 (N_19709,N_19582,N_19513);
xor U19710 (N_19710,N_19457,N_19418);
or U19711 (N_19711,N_19521,N_19577);
nor U19712 (N_19712,N_19453,N_19429);
nor U19713 (N_19713,N_19479,N_19577);
or U19714 (N_19714,N_19450,N_19514);
nor U19715 (N_19715,N_19424,N_19437);
xor U19716 (N_19716,N_19545,N_19528);
xor U19717 (N_19717,N_19499,N_19577);
nand U19718 (N_19718,N_19540,N_19569);
nor U19719 (N_19719,N_19591,N_19433);
and U19720 (N_19720,N_19558,N_19463);
and U19721 (N_19721,N_19424,N_19488);
nand U19722 (N_19722,N_19449,N_19489);
nand U19723 (N_19723,N_19459,N_19521);
and U19724 (N_19724,N_19417,N_19451);
nor U19725 (N_19725,N_19417,N_19511);
nand U19726 (N_19726,N_19435,N_19483);
nand U19727 (N_19727,N_19481,N_19551);
xnor U19728 (N_19728,N_19439,N_19443);
or U19729 (N_19729,N_19481,N_19452);
xor U19730 (N_19730,N_19493,N_19468);
xnor U19731 (N_19731,N_19451,N_19547);
xor U19732 (N_19732,N_19501,N_19515);
or U19733 (N_19733,N_19558,N_19485);
and U19734 (N_19734,N_19523,N_19537);
and U19735 (N_19735,N_19593,N_19545);
or U19736 (N_19736,N_19560,N_19407);
nor U19737 (N_19737,N_19528,N_19496);
nand U19738 (N_19738,N_19471,N_19432);
xor U19739 (N_19739,N_19408,N_19517);
nand U19740 (N_19740,N_19464,N_19457);
or U19741 (N_19741,N_19549,N_19504);
xnor U19742 (N_19742,N_19408,N_19566);
xor U19743 (N_19743,N_19546,N_19422);
and U19744 (N_19744,N_19594,N_19508);
and U19745 (N_19745,N_19555,N_19558);
xor U19746 (N_19746,N_19552,N_19597);
nand U19747 (N_19747,N_19485,N_19501);
nand U19748 (N_19748,N_19451,N_19560);
and U19749 (N_19749,N_19574,N_19425);
nor U19750 (N_19750,N_19415,N_19482);
xor U19751 (N_19751,N_19409,N_19473);
nor U19752 (N_19752,N_19549,N_19433);
nor U19753 (N_19753,N_19425,N_19553);
nand U19754 (N_19754,N_19439,N_19425);
and U19755 (N_19755,N_19591,N_19494);
xor U19756 (N_19756,N_19534,N_19587);
nor U19757 (N_19757,N_19567,N_19517);
or U19758 (N_19758,N_19561,N_19576);
nor U19759 (N_19759,N_19461,N_19471);
and U19760 (N_19760,N_19436,N_19521);
nand U19761 (N_19761,N_19573,N_19514);
xnor U19762 (N_19762,N_19471,N_19416);
and U19763 (N_19763,N_19514,N_19473);
or U19764 (N_19764,N_19410,N_19407);
or U19765 (N_19765,N_19422,N_19429);
xor U19766 (N_19766,N_19531,N_19440);
nor U19767 (N_19767,N_19522,N_19411);
nor U19768 (N_19768,N_19590,N_19472);
nand U19769 (N_19769,N_19598,N_19550);
nand U19770 (N_19770,N_19417,N_19445);
xnor U19771 (N_19771,N_19545,N_19580);
and U19772 (N_19772,N_19569,N_19520);
and U19773 (N_19773,N_19552,N_19596);
nand U19774 (N_19774,N_19587,N_19589);
and U19775 (N_19775,N_19488,N_19514);
nor U19776 (N_19776,N_19529,N_19528);
and U19777 (N_19777,N_19421,N_19484);
nand U19778 (N_19778,N_19456,N_19556);
xnor U19779 (N_19779,N_19419,N_19459);
nor U19780 (N_19780,N_19425,N_19562);
and U19781 (N_19781,N_19435,N_19437);
or U19782 (N_19782,N_19548,N_19507);
nand U19783 (N_19783,N_19426,N_19401);
and U19784 (N_19784,N_19400,N_19464);
xor U19785 (N_19785,N_19515,N_19558);
nand U19786 (N_19786,N_19567,N_19472);
or U19787 (N_19787,N_19423,N_19410);
and U19788 (N_19788,N_19468,N_19403);
nor U19789 (N_19789,N_19449,N_19425);
and U19790 (N_19790,N_19585,N_19527);
and U19791 (N_19791,N_19595,N_19444);
and U19792 (N_19792,N_19463,N_19541);
nor U19793 (N_19793,N_19442,N_19498);
nor U19794 (N_19794,N_19449,N_19542);
xor U19795 (N_19795,N_19476,N_19441);
nor U19796 (N_19796,N_19500,N_19528);
and U19797 (N_19797,N_19502,N_19471);
nand U19798 (N_19798,N_19561,N_19427);
xnor U19799 (N_19799,N_19428,N_19467);
nand U19800 (N_19800,N_19732,N_19775);
xor U19801 (N_19801,N_19702,N_19785);
nor U19802 (N_19802,N_19784,N_19722);
xnor U19803 (N_19803,N_19710,N_19641);
nand U19804 (N_19804,N_19758,N_19723);
xnor U19805 (N_19805,N_19781,N_19706);
or U19806 (N_19806,N_19741,N_19639);
xor U19807 (N_19807,N_19675,N_19672);
or U19808 (N_19808,N_19795,N_19765);
and U19809 (N_19809,N_19657,N_19633);
xnor U19810 (N_19810,N_19792,N_19767);
or U19811 (N_19811,N_19618,N_19786);
nor U19812 (N_19812,N_19678,N_19681);
nand U19813 (N_19813,N_19776,N_19659);
nor U19814 (N_19814,N_19747,N_19616);
or U19815 (N_19815,N_19717,N_19773);
and U19816 (N_19816,N_19654,N_19794);
nor U19817 (N_19817,N_19661,N_19606);
nor U19818 (N_19818,N_19688,N_19696);
nand U19819 (N_19819,N_19620,N_19768);
and U19820 (N_19820,N_19662,N_19656);
or U19821 (N_19821,N_19651,N_19714);
and U19822 (N_19822,N_19730,N_19629);
and U19823 (N_19823,N_19752,N_19671);
or U19824 (N_19824,N_19729,N_19685);
or U19825 (N_19825,N_19783,N_19631);
nand U19826 (N_19826,N_19771,N_19621);
xnor U19827 (N_19827,N_19611,N_19780);
nand U19828 (N_19828,N_19782,N_19777);
nand U19829 (N_19829,N_19721,N_19740);
nand U19830 (N_19830,N_19649,N_19716);
nand U19831 (N_19831,N_19738,N_19610);
xnor U19832 (N_19832,N_19701,N_19724);
and U19833 (N_19833,N_19684,N_19600);
and U19834 (N_19834,N_19719,N_19769);
nand U19835 (N_19835,N_19602,N_19687);
nor U19836 (N_19836,N_19759,N_19609);
and U19837 (N_19837,N_19756,N_19680);
nor U19838 (N_19838,N_19770,N_19615);
nand U19839 (N_19839,N_19778,N_19601);
nand U19840 (N_19840,N_19617,N_19718);
xnor U19841 (N_19841,N_19734,N_19625);
nor U19842 (N_19842,N_19699,N_19622);
and U19843 (N_19843,N_19733,N_19604);
or U19844 (N_19844,N_19636,N_19664);
or U19845 (N_19845,N_19712,N_19720);
xnor U19846 (N_19846,N_19709,N_19796);
nor U19847 (N_19847,N_19731,N_19772);
nor U19848 (N_19848,N_19605,N_19644);
nor U19849 (N_19849,N_19739,N_19787);
nor U19850 (N_19850,N_19623,N_19630);
nand U19851 (N_19851,N_19726,N_19670);
xor U19852 (N_19852,N_19725,N_19643);
xnor U19853 (N_19853,N_19647,N_19637);
xnor U19854 (N_19854,N_19648,N_19750);
and U19855 (N_19855,N_19763,N_19612);
nand U19856 (N_19856,N_19757,N_19632);
nor U19857 (N_19857,N_19789,N_19735);
xnor U19858 (N_19858,N_19744,N_19603);
nand U19859 (N_19859,N_19798,N_19779);
and U19860 (N_19860,N_19627,N_19715);
and U19861 (N_19861,N_19634,N_19624);
and U19862 (N_19862,N_19658,N_19799);
and U19863 (N_19863,N_19665,N_19628);
or U19864 (N_19864,N_19761,N_19727);
xor U19865 (N_19865,N_19743,N_19746);
xnor U19866 (N_19866,N_19690,N_19790);
xor U19867 (N_19867,N_19797,N_19660);
nor U19868 (N_19868,N_19693,N_19686);
xnor U19869 (N_19869,N_19754,N_19673);
xor U19870 (N_19870,N_19676,N_19691);
nand U19871 (N_19871,N_19703,N_19793);
xnor U19872 (N_19872,N_19642,N_19652);
nor U19873 (N_19873,N_19791,N_19774);
xnor U19874 (N_19874,N_19764,N_19704);
or U19875 (N_19875,N_19638,N_19708);
nand U19876 (N_19876,N_19650,N_19745);
xor U19877 (N_19877,N_19753,N_19698);
and U19878 (N_19878,N_19626,N_19697);
or U19879 (N_19879,N_19683,N_19653);
or U19880 (N_19880,N_19667,N_19668);
or U19881 (N_19881,N_19762,N_19695);
nor U19882 (N_19882,N_19635,N_19760);
or U19883 (N_19883,N_19694,N_19679);
or U19884 (N_19884,N_19728,N_19608);
nor U19885 (N_19885,N_19619,N_19640);
nor U19886 (N_19886,N_19713,N_19669);
or U19887 (N_19887,N_19646,N_19755);
nand U19888 (N_19888,N_19645,N_19748);
and U19889 (N_19889,N_19614,N_19707);
nand U19890 (N_19890,N_19742,N_19689);
or U19891 (N_19891,N_19700,N_19682);
xor U19892 (N_19892,N_19751,N_19788);
or U19893 (N_19893,N_19655,N_19737);
nor U19894 (N_19894,N_19674,N_19666);
xnor U19895 (N_19895,N_19705,N_19736);
xnor U19896 (N_19896,N_19692,N_19663);
and U19897 (N_19897,N_19749,N_19613);
nand U19898 (N_19898,N_19607,N_19766);
or U19899 (N_19899,N_19677,N_19711);
xnor U19900 (N_19900,N_19724,N_19702);
xor U19901 (N_19901,N_19679,N_19616);
nand U19902 (N_19902,N_19732,N_19785);
or U19903 (N_19903,N_19750,N_19733);
nor U19904 (N_19904,N_19606,N_19636);
nor U19905 (N_19905,N_19618,N_19678);
and U19906 (N_19906,N_19791,N_19651);
or U19907 (N_19907,N_19607,N_19675);
nand U19908 (N_19908,N_19693,N_19796);
xor U19909 (N_19909,N_19624,N_19696);
or U19910 (N_19910,N_19723,N_19752);
xnor U19911 (N_19911,N_19730,N_19789);
xnor U19912 (N_19912,N_19679,N_19696);
or U19913 (N_19913,N_19636,N_19672);
and U19914 (N_19914,N_19680,N_19654);
nand U19915 (N_19915,N_19728,N_19629);
or U19916 (N_19916,N_19771,N_19647);
and U19917 (N_19917,N_19678,N_19791);
nand U19918 (N_19918,N_19748,N_19659);
xnor U19919 (N_19919,N_19607,N_19753);
and U19920 (N_19920,N_19738,N_19743);
or U19921 (N_19921,N_19687,N_19623);
xnor U19922 (N_19922,N_19637,N_19618);
or U19923 (N_19923,N_19640,N_19781);
and U19924 (N_19924,N_19639,N_19627);
or U19925 (N_19925,N_19603,N_19736);
or U19926 (N_19926,N_19680,N_19732);
and U19927 (N_19927,N_19770,N_19709);
nand U19928 (N_19928,N_19632,N_19736);
or U19929 (N_19929,N_19799,N_19644);
and U19930 (N_19930,N_19685,N_19621);
xor U19931 (N_19931,N_19756,N_19744);
nor U19932 (N_19932,N_19755,N_19688);
or U19933 (N_19933,N_19756,N_19761);
nand U19934 (N_19934,N_19635,N_19768);
nor U19935 (N_19935,N_19788,N_19601);
or U19936 (N_19936,N_19651,N_19758);
nand U19937 (N_19937,N_19681,N_19742);
and U19938 (N_19938,N_19643,N_19601);
xnor U19939 (N_19939,N_19691,N_19643);
and U19940 (N_19940,N_19666,N_19617);
nand U19941 (N_19941,N_19770,N_19643);
nand U19942 (N_19942,N_19759,N_19651);
nand U19943 (N_19943,N_19714,N_19725);
nand U19944 (N_19944,N_19635,N_19604);
and U19945 (N_19945,N_19778,N_19794);
nand U19946 (N_19946,N_19767,N_19726);
nor U19947 (N_19947,N_19656,N_19681);
nor U19948 (N_19948,N_19653,N_19663);
nor U19949 (N_19949,N_19793,N_19754);
nor U19950 (N_19950,N_19683,N_19609);
and U19951 (N_19951,N_19769,N_19697);
nand U19952 (N_19952,N_19717,N_19766);
nor U19953 (N_19953,N_19602,N_19675);
or U19954 (N_19954,N_19618,N_19792);
xor U19955 (N_19955,N_19699,N_19744);
and U19956 (N_19956,N_19633,N_19767);
nor U19957 (N_19957,N_19648,N_19771);
nand U19958 (N_19958,N_19767,N_19685);
xnor U19959 (N_19959,N_19715,N_19676);
or U19960 (N_19960,N_19779,N_19677);
xnor U19961 (N_19961,N_19759,N_19770);
and U19962 (N_19962,N_19680,N_19784);
and U19963 (N_19963,N_19782,N_19720);
or U19964 (N_19964,N_19681,N_19693);
nor U19965 (N_19965,N_19728,N_19699);
xor U19966 (N_19966,N_19776,N_19685);
nand U19967 (N_19967,N_19677,N_19705);
nand U19968 (N_19968,N_19666,N_19775);
or U19969 (N_19969,N_19673,N_19799);
nand U19970 (N_19970,N_19704,N_19673);
nor U19971 (N_19971,N_19638,N_19729);
xor U19972 (N_19972,N_19776,N_19779);
and U19973 (N_19973,N_19696,N_19703);
or U19974 (N_19974,N_19662,N_19612);
xnor U19975 (N_19975,N_19662,N_19631);
nand U19976 (N_19976,N_19702,N_19656);
and U19977 (N_19977,N_19639,N_19718);
nand U19978 (N_19978,N_19738,N_19754);
or U19979 (N_19979,N_19620,N_19784);
nand U19980 (N_19980,N_19773,N_19623);
nand U19981 (N_19981,N_19706,N_19738);
nor U19982 (N_19982,N_19787,N_19616);
nand U19983 (N_19983,N_19688,N_19770);
nor U19984 (N_19984,N_19628,N_19744);
nand U19985 (N_19985,N_19774,N_19628);
nand U19986 (N_19986,N_19719,N_19644);
and U19987 (N_19987,N_19687,N_19725);
xnor U19988 (N_19988,N_19665,N_19732);
xnor U19989 (N_19989,N_19648,N_19664);
xor U19990 (N_19990,N_19788,N_19737);
nand U19991 (N_19991,N_19725,N_19717);
nor U19992 (N_19992,N_19642,N_19701);
xor U19993 (N_19993,N_19738,N_19744);
xor U19994 (N_19994,N_19620,N_19624);
or U19995 (N_19995,N_19626,N_19672);
nand U19996 (N_19996,N_19680,N_19640);
nand U19997 (N_19997,N_19602,N_19708);
nor U19998 (N_19998,N_19633,N_19717);
and U19999 (N_19999,N_19720,N_19631);
or U20000 (N_20000,N_19994,N_19833);
nor U20001 (N_20001,N_19878,N_19811);
xnor U20002 (N_20002,N_19835,N_19890);
and U20003 (N_20003,N_19989,N_19889);
and U20004 (N_20004,N_19856,N_19942);
xnor U20005 (N_20005,N_19933,N_19941);
nand U20006 (N_20006,N_19844,N_19903);
xor U20007 (N_20007,N_19803,N_19988);
nand U20008 (N_20008,N_19888,N_19852);
nand U20009 (N_20009,N_19805,N_19965);
nor U20010 (N_20010,N_19993,N_19914);
nand U20011 (N_20011,N_19821,N_19998);
nor U20012 (N_20012,N_19885,N_19945);
or U20013 (N_20013,N_19930,N_19800);
or U20014 (N_20014,N_19936,N_19912);
and U20015 (N_20015,N_19983,N_19915);
or U20016 (N_20016,N_19971,N_19947);
or U20017 (N_20017,N_19809,N_19935);
nand U20018 (N_20018,N_19975,N_19827);
nand U20019 (N_20019,N_19812,N_19831);
or U20020 (N_20020,N_19834,N_19946);
nand U20021 (N_20021,N_19931,N_19876);
or U20022 (N_20022,N_19963,N_19979);
and U20023 (N_20023,N_19860,N_19828);
nand U20024 (N_20024,N_19956,N_19958);
nor U20025 (N_20025,N_19985,N_19817);
and U20026 (N_20026,N_19891,N_19948);
nor U20027 (N_20027,N_19986,N_19850);
or U20028 (N_20028,N_19925,N_19918);
and U20029 (N_20029,N_19801,N_19858);
and U20030 (N_20030,N_19937,N_19870);
xor U20031 (N_20031,N_19882,N_19953);
nand U20032 (N_20032,N_19845,N_19934);
or U20033 (N_20033,N_19922,N_19893);
xor U20034 (N_20034,N_19892,N_19902);
and U20035 (N_20035,N_19978,N_19807);
nor U20036 (N_20036,N_19961,N_19977);
xor U20037 (N_20037,N_19967,N_19932);
and U20038 (N_20038,N_19949,N_19887);
nor U20039 (N_20039,N_19830,N_19943);
and U20040 (N_20040,N_19940,N_19897);
xor U20041 (N_20041,N_19984,N_19841);
or U20042 (N_20042,N_19901,N_19847);
xor U20043 (N_20043,N_19871,N_19881);
nor U20044 (N_20044,N_19944,N_19906);
and U20045 (N_20045,N_19866,N_19968);
nor U20046 (N_20046,N_19981,N_19895);
xor U20047 (N_20047,N_19883,N_19825);
or U20048 (N_20048,N_19861,N_19962);
and U20049 (N_20049,N_19859,N_19910);
and U20050 (N_20050,N_19960,N_19957);
nand U20051 (N_20051,N_19884,N_19992);
nor U20052 (N_20052,N_19873,N_19829);
nand U20053 (N_20053,N_19969,N_19813);
nand U20054 (N_20054,N_19973,N_19818);
nor U20055 (N_20055,N_19880,N_19904);
nand U20056 (N_20056,N_19974,N_19819);
xnor U20057 (N_20057,N_19877,N_19972);
and U20058 (N_20058,N_19980,N_19919);
nand U20059 (N_20059,N_19837,N_19836);
nand U20060 (N_20060,N_19802,N_19874);
nor U20061 (N_20061,N_19926,N_19854);
or U20062 (N_20062,N_19900,N_19929);
xnor U20063 (N_20063,N_19938,N_19954);
and U20064 (N_20064,N_19851,N_19997);
and U20065 (N_20065,N_19822,N_19909);
or U20066 (N_20066,N_19959,N_19843);
and U20067 (N_20067,N_19868,N_19886);
and U20068 (N_20068,N_19982,N_19864);
nor U20069 (N_20069,N_19966,N_19816);
and U20070 (N_20070,N_19894,N_19928);
and U20071 (N_20071,N_19939,N_19995);
xnor U20072 (N_20072,N_19848,N_19826);
nor U20073 (N_20073,N_19863,N_19867);
or U20074 (N_20074,N_19950,N_19808);
nand U20075 (N_20075,N_19879,N_19899);
or U20076 (N_20076,N_19842,N_19921);
or U20077 (N_20077,N_19832,N_19896);
xnor U20078 (N_20078,N_19853,N_19804);
or U20079 (N_20079,N_19857,N_19849);
and U20080 (N_20080,N_19996,N_19970);
xnor U20081 (N_20081,N_19955,N_19991);
nand U20082 (N_20082,N_19964,N_19840);
and U20083 (N_20083,N_19913,N_19990);
xnor U20084 (N_20084,N_19924,N_19907);
xor U20085 (N_20085,N_19824,N_19862);
and U20086 (N_20086,N_19927,N_19814);
xor U20087 (N_20087,N_19905,N_19806);
or U20088 (N_20088,N_19999,N_19815);
or U20089 (N_20089,N_19917,N_19838);
and U20090 (N_20090,N_19920,N_19869);
xnor U20091 (N_20091,N_19976,N_19951);
nand U20092 (N_20092,N_19839,N_19952);
nor U20093 (N_20093,N_19908,N_19875);
nor U20094 (N_20094,N_19855,N_19923);
xor U20095 (N_20095,N_19810,N_19898);
nand U20096 (N_20096,N_19865,N_19846);
xnor U20097 (N_20097,N_19916,N_19872);
nand U20098 (N_20098,N_19911,N_19987);
and U20099 (N_20099,N_19823,N_19820);
and U20100 (N_20100,N_19923,N_19866);
nand U20101 (N_20101,N_19975,N_19876);
nand U20102 (N_20102,N_19995,N_19979);
or U20103 (N_20103,N_19813,N_19948);
or U20104 (N_20104,N_19910,N_19857);
xnor U20105 (N_20105,N_19958,N_19942);
xnor U20106 (N_20106,N_19826,N_19829);
nor U20107 (N_20107,N_19940,N_19854);
or U20108 (N_20108,N_19891,N_19867);
nand U20109 (N_20109,N_19919,N_19984);
and U20110 (N_20110,N_19928,N_19808);
nor U20111 (N_20111,N_19972,N_19920);
and U20112 (N_20112,N_19917,N_19926);
xnor U20113 (N_20113,N_19890,N_19924);
or U20114 (N_20114,N_19807,N_19971);
nand U20115 (N_20115,N_19960,N_19873);
and U20116 (N_20116,N_19877,N_19875);
or U20117 (N_20117,N_19933,N_19931);
nand U20118 (N_20118,N_19962,N_19865);
xor U20119 (N_20119,N_19809,N_19993);
nor U20120 (N_20120,N_19980,N_19882);
and U20121 (N_20121,N_19966,N_19866);
nand U20122 (N_20122,N_19866,N_19940);
or U20123 (N_20123,N_19985,N_19869);
xor U20124 (N_20124,N_19879,N_19997);
and U20125 (N_20125,N_19923,N_19936);
xnor U20126 (N_20126,N_19921,N_19907);
or U20127 (N_20127,N_19889,N_19867);
and U20128 (N_20128,N_19913,N_19896);
nor U20129 (N_20129,N_19926,N_19994);
nand U20130 (N_20130,N_19960,N_19946);
or U20131 (N_20131,N_19861,N_19916);
nor U20132 (N_20132,N_19880,N_19923);
or U20133 (N_20133,N_19882,N_19833);
and U20134 (N_20134,N_19951,N_19989);
or U20135 (N_20135,N_19884,N_19829);
xnor U20136 (N_20136,N_19886,N_19835);
nor U20137 (N_20137,N_19830,N_19864);
xnor U20138 (N_20138,N_19968,N_19936);
and U20139 (N_20139,N_19900,N_19906);
nand U20140 (N_20140,N_19872,N_19918);
nor U20141 (N_20141,N_19842,N_19831);
and U20142 (N_20142,N_19883,N_19833);
or U20143 (N_20143,N_19974,N_19939);
and U20144 (N_20144,N_19986,N_19969);
nor U20145 (N_20145,N_19958,N_19997);
nand U20146 (N_20146,N_19835,N_19872);
and U20147 (N_20147,N_19859,N_19857);
xor U20148 (N_20148,N_19879,N_19948);
nor U20149 (N_20149,N_19914,N_19933);
nand U20150 (N_20150,N_19906,N_19863);
or U20151 (N_20151,N_19856,N_19825);
nand U20152 (N_20152,N_19874,N_19875);
and U20153 (N_20153,N_19873,N_19941);
nor U20154 (N_20154,N_19975,N_19965);
or U20155 (N_20155,N_19879,N_19823);
xnor U20156 (N_20156,N_19907,N_19923);
and U20157 (N_20157,N_19849,N_19860);
nor U20158 (N_20158,N_19973,N_19996);
nor U20159 (N_20159,N_19874,N_19918);
xnor U20160 (N_20160,N_19987,N_19932);
or U20161 (N_20161,N_19994,N_19911);
or U20162 (N_20162,N_19994,N_19856);
and U20163 (N_20163,N_19984,N_19910);
xnor U20164 (N_20164,N_19853,N_19908);
and U20165 (N_20165,N_19906,N_19854);
or U20166 (N_20166,N_19963,N_19832);
and U20167 (N_20167,N_19836,N_19958);
nor U20168 (N_20168,N_19973,N_19902);
xnor U20169 (N_20169,N_19873,N_19824);
xnor U20170 (N_20170,N_19859,N_19809);
nor U20171 (N_20171,N_19934,N_19909);
nand U20172 (N_20172,N_19961,N_19967);
and U20173 (N_20173,N_19941,N_19959);
xor U20174 (N_20174,N_19958,N_19953);
nor U20175 (N_20175,N_19923,N_19894);
xnor U20176 (N_20176,N_19880,N_19991);
nand U20177 (N_20177,N_19846,N_19985);
or U20178 (N_20178,N_19830,N_19848);
and U20179 (N_20179,N_19892,N_19837);
xnor U20180 (N_20180,N_19848,N_19853);
nor U20181 (N_20181,N_19900,N_19865);
xor U20182 (N_20182,N_19933,N_19910);
nand U20183 (N_20183,N_19803,N_19901);
or U20184 (N_20184,N_19958,N_19825);
or U20185 (N_20185,N_19961,N_19950);
nor U20186 (N_20186,N_19891,N_19997);
and U20187 (N_20187,N_19848,N_19859);
nand U20188 (N_20188,N_19806,N_19956);
nor U20189 (N_20189,N_19956,N_19916);
nand U20190 (N_20190,N_19984,N_19939);
or U20191 (N_20191,N_19967,N_19874);
nor U20192 (N_20192,N_19815,N_19824);
xnor U20193 (N_20193,N_19951,N_19845);
nor U20194 (N_20194,N_19830,N_19904);
xnor U20195 (N_20195,N_19881,N_19838);
and U20196 (N_20196,N_19867,N_19900);
xor U20197 (N_20197,N_19888,N_19857);
nor U20198 (N_20198,N_19810,N_19903);
nand U20199 (N_20199,N_19813,N_19954);
nand U20200 (N_20200,N_20170,N_20147);
and U20201 (N_20201,N_20165,N_20120);
xor U20202 (N_20202,N_20175,N_20127);
xor U20203 (N_20203,N_20145,N_20029);
nand U20204 (N_20204,N_20198,N_20140);
or U20205 (N_20205,N_20099,N_20049);
nand U20206 (N_20206,N_20061,N_20011);
and U20207 (N_20207,N_20015,N_20042);
and U20208 (N_20208,N_20133,N_20155);
or U20209 (N_20209,N_20173,N_20027);
nand U20210 (N_20210,N_20081,N_20050);
xor U20211 (N_20211,N_20076,N_20067);
or U20212 (N_20212,N_20113,N_20051);
nand U20213 (N_20213,N_20153,N_20197);
nor U20214 (N_20214,N_20199,N_20169);
and U20215 (N_20215,N_20040,N_20053);
nand U20216 (N_20216,N_20037,N_20137);
and U20217 (N_20217,N_20186,N_20152);
nand U20218 (N_20218,N_20012,N_20097);
and U20219 (N_20219,N_20154,N_20024);
or U20220 (N_20220,N_20148,N_20026);
nor U20221 (N_20221,N_20104,N_20036);
or U20222 (N_20222,N_20072,N_20074);
nand U20223 (N_20223,N_20022,N_20008);
and U20224 (N_20224,N_20183,N_20045);
and U20225 (N_20225,N_20160,N_20002);
and U20226 (N_20226,N_20192,N_20082);
nor U20227 (N_20227,N_20054,N_20089);
or U20228 (N_20228,N_20064,N_20098);
nor U20229 (N_20229,N_20052,N_20003);
or U20230 (N_20230,N_20041,N_20117);
xor U20231 (N_20231,N_20185,N_20060);
nand U20232 (N_20232,N_20068,N_20124);
xor U20233 (N_20233,N_20078,N_20126);
and U20234 (N_20234,N_20058,N_20069);
nand U20235 (N_20235,N_20146,N_20095);
and U20236 (N_20236,N_20073,N_20034);
xor U20237 (N_20237,N_20167,N_20163);
xor U20238 (N_20238,N_20014,N_20010);
nor U20239 (N_20239,N_20108,N_20056);
or U20240 (N_20240,N_20071,N_20013);
or U20241 (N_20241,N_20000,N_20087);
nor U20242 (N_20242,N_20066,N_20080);
nor U20243 (N_20243,N_20059,N_20122);
xor U20244 (N_20244,N_20180,N_20116);
xnor U20245 (N_20245,N_20166,N_20189);
xor U20246 (N_20246,N_20107,N_20128);
or U20247 (N_20247,N_20179,N_20031);
nor U20248 (N_20248,N_20090,N_20168);
and U20249 (N_20249,N_20130,N_20001);
nor U20250 (N_20250,N_20009,N_20038);
and U20251 (N_20251,N_20193,N_20057);
nand U20252 (N_20252,N_20079,N_20190);
nor U20253 (N_20253,N_20141,N_20084);
or U20254 (N_20254,N_20184,N_20156);
nor U20255 (N_20255,N_20083,N_20018);
nand U20256 (N_20256,N_20149,N_20023);
and U20257 (N_20257,N_20096,N_20101);
or U20258 (N_20258,N_20062,N_20070);
or U20259 (N_20259,N_20043,N_20159);
nor U20260 (N_20260,N_20187,N_20158);
or U20261 (N_20261,N_20016,N_20085);
and U20262 (N_20262,N_20030,N_20119);
nor U20263 (N_20263,N_20188,N_20177);
nor U20264 (N_20264,N_20077,N_20161);
xnor U20265 (N_20265,N_20150,N_20109);
or U20266 (N_20266,N_20005,N_20102);
nand U20267 (N_20267,N_20004,N_20176);
xnor U20268 (N_20268,N_20093,N_20194);
nand U20269 (N_20269,N_20020,N_20118);
or U20270 (N_20270,N_20181,N_20094);
xnor U20271 (N_20271,N_20103,N_20063);
or U20272 (N_20272,N_20172,N_20017);
and U20273 (N_20273,N_20196,N_20138);
xor U20274 (N_20274,N_20065,N_20135);
xnor U20275 (N_20275,N_20021,N_20139);
and U20276 (N_20276,N_20088,N_20171);
nor U20277 (N_20277,N_20164,N_20131);
nand U20278 (N_20278,N_20157,N_20143);
nand U20279 (N_20279,N_20006,N_20055);
nor U20280 (N_20280,N_20182,N_20007);
or U20281 (N_20281,N_20110,N_20132);
nor U20282 (N_20282,N_20129,N_20039);
and U20283 (N_20283,N_20178,N_20033);
xnor U20284 (N_20284,N_20162,N_20123);
nor U20285 (N_20285,N_20174,N_20121);
nand U20286 (N_20286,N_20114,N_20195);
or U20287 (N_20287,N_20019,N_20047);
nor U20288 (N_20288,N_20032,N_20100);
nor U20289 (N_20289,N_20044,N_20125);
xor U20290 (N_20290,N_20035,N_20086);
nor U20291 (N_20291,N_20134,N_20106);
xnor U20292 (N_20292,N_20028,N_20191);
or U20293 (N_20293,N_20112,N_20115);
or U20294 (N_20294,N_20092,N_20136);
or U20295 (N_20295,N_20048,N_20075);
nand U20296 (N_20296,N_20142,N_20151);
or U20297 (N_20297,N_20091,N_20025);
nor U20298 (N_20298,N_20046,N_20144);
nor U20299 (N_20299,N_20105,N_20111);
or U20300 (N_20300,N_20180,N_20098);
and U20301 (N_20301,N_20154,N_20147);
and U20302 (N_20302,N_20016,N_20024);
nor U20303 (N_20303,N_20105,N_20171);
nand U20304 (N_20304,N_20061,N_20090);
nor U20305 (N_20305,N_20104,N_20105);
or U20306 (N_20306,N_20131,N_20183);
and U20307 (N_20307,N_20128,N_20015);
or U20308 (N_20308,N_20106,N_20025);
nor U20309 (N_20309,N_20012,N_20039);
nor U20310 (N_20310,N_20028,N_20193);
and U20311 (N_20311,N_20055,N_20155);
nor U20312 (N_20312,N_20142,N_20110);
xor U20313 (N_20313,N_20185,N_20036);
xor U20314 (N_20314,N_20199,N_20063);
nor U20315 (N_20315,N_20056,N_20048);
and U20316 (N_20316,N_20061,N_20047);
and U20317 (N_20317,N_20117,N_20084);
or U20318 (N_20318,N_20039,N_20150);
or U20319 (N_20319,N_20092,N_20050);
xnor U20320 (N_20320,N_20073,N_20153);
and U20321 (N_20321,N_20138,N_20124);
and U20322 (N_20322,N_20036,N_20121);
and U20323 (N_20323,N_20112,N_20073);
nand U20324 (N_20324,N_20068,N_20015);
nor U20325 (N_20325,N_20025,N_20129);
or U20326 (N_20326,N_20145,N_20007);
or U20327 (N_20327,N_20012,N_20117);
nand U20328 (N_20328,N_20065,N_20057);
xor U20329 (N_20329,N_20067,N_20143);
nand U20330 (N_20330,N_20058,N_20198);
and U20331 (N_20331,N_20082,N_20137);
and U20332 (N_20332,N_20116,N_20156);
xnor U20333 (N_20333,N_20195,N_20048);
nor U20334 (N_20334,N_20073,N_20165);
and U20335 (N_20335,N_20179,N_20081);
or U20336 (N_20336,N_20034,N_20185);
nand U20337 (N_20337,N_20078,N_20090);
nand U20338 (N_20338,N_20166,N_20144);
or U20339 (N_20339,N_20064,N_20094);
nand U20340 (N_20340,N_20090,N_20065);
or U20341 (N_20341,N_20160,N_20015);
nor U20342 (N_20342,N_20124,N_20024);
nand U20343 (N_20343,N_20073,N_20130);
and U20344 (N_20344,N_20109,N_20107);
or U20345 (N_20345,N_20092,N_20022);
nor U20346 (N_20346,N_20176,N_20172);
and U20347 (N_20347,N_20022,N_20042);
or U20348 (N_20348,N_20151,N_20147);
nand U20349 (N_20349,N_20080,N_20082);
and U20350 (N_20350,N_20110,N_20026);
nand U20351 (N_20351,N_20015,N_20036);
and U20352 (N_20352,N_20051,N_20085);
or U20353 (N_20353,N_20138,N_20191);
nand U20354 (N_20354,N_20168,N_20018);
and U20355 (N_20355,N_20045,N_20069);
xor U20356 (N_20356,N_20142,N_20086);
and U20357 (N_20357,N_20133,N_20149);
nand U20358 (N_20358,N_20143,N_20050);
or U20359 (N_20359,N_20132,N_20024);
xor U20360 (N_20360,N_20058,N_20006);
nor U20361 (N_20361,N_20171,N_20073);
nand U20362 (N_20362,N_20152,N_20172);
nor U20363 (N_20363,N_20143,N_20069);
nand U20364 (N_20364,N_20072,N_20100);
and U20365 (N_20365,N_20080,N_20158);
nand U20366 (N_20366,N_20033,N_20143);
and U20367 (N_20367,N_20009,N_20095);
nor U20368 (N_20368,N_20049,N_20037);
or U20369 (N_20369,N_20152,N_20197);
or U20370 (N_20370,N_20186,N_20148);
xor U20371 (N_20371,N_20006,N_20109);
or U20372 (N_20372,N_20001,N_20005);
and U20373 (N_20373,N_20086,N_20029);
nand U20374 (N_20374,N_20163,N_20099);
or U20375 (N_20375,N_20173,N_20151);
nand U20376 (N_20376,N_20185,N_20147);
and U20377 (N_20377,N_20097,N_20178);
nor U20378 (N_20378,N_20118,N_20166);
nor U20379 (N_20379,N_20151,N_20180);
nor U20380 (N_20380,N_20112,N_20199);
or U20381 (N_20381,N_20095,N_20018);
or U20382 (N_20382,N_20189,N_20024);
or U20383 (N_20383,N_20114,N_20170);
nor U20384 (N_20384,N_20130,N_20019);
nand U20385 (N_20385,N_20061,N_20163);
or U20386 (N_20386,N_20003,N_20018);
or U20387 (N_20387,N_20126,N_20119);
nor U20388 (N_20388,N_20121,N_20126);
or U20389 (N_20389,N_20067,N_20164);
nand U20390 (N_20390,N_20137,N_20056);
nor U20391 (N_20391,N_20194,N_20188);
or U20392 (N_20392,N_20027,N_20112);
xor U20393 (N_20393,N_20189,N_20052);
or U20394 (N_20394,N_20171,N_20086);
xnor U20395 (N_20395,N_20076,N_20154);
nand U20396 (N_20396,N_20166,N_20049);
nand U20397 (N_20397,N_20010,N_20034);
and U20398 (N_20398,N_20085,N_20198);
xnor U20399 (N_20399,N_20144,N_20160);
or U20400 (N_20400,N_20268,N_20214);
xnor U20401 (N_20401,N_20232,N_20242);
and U20402 (N_20402,N_20200,N_20269);
nand U20403 (N_20403,N_20288,N_20384);
or U20404 (N_20404,N_20292,N_20320);
nor U20405 (N_20405,N_20371,N_20306);
and U20406 (N_20406,N_20248,N_20243);
nand U20407 (N_20407,N_20287,N_20224);
nand U20408 (N_20408,N_20213,N_20303);
nor U20409 (N_20409,N_20328,N_20314);
nand U20410 (N_20410,N_20207,N_20256);
or U20411 (N_20411,N_20250,N_20298);
xnor U20412 (N_20412,N_20376,N_20259);
xnor U20413 (N_20413,N_20286,N_20291);
and U20414 (N_20414,N_20323,N_20229);
or U20415 (N_20415,N_20319,N_20349);
or U20416 (N_20416,N_20249,N_20329);
nor U20417 (N_20417,N_20341,N_20392);
or U20418 (N_20418,N_20223,N_20344);
and U20419 (N_20419,N_20300,N_20258);
xnor U20420 (N_20420,N_20369,N_20296);
and U20421 (N_20421,N_20273,N_20277);
and U20422 (N_20422,N_20297,N_20343);
or U20423 (N_20423,N_20363,N_20218);
xor U20424 (N_20424,N_20347,N_20210);
nor U20425 (N_20425,N_20271,N_20342);
nor U20426 (N_20426,N_20237,N_20310);
xor U20427 (N_20427,N_20348,N_20365);
and U20428 (N_20428,N_20331,N_20275);
nor U20429 (N_20429,N_20370,N_20366);
nand U20430 (N_20430,N_20318,N_20230);
and U20431 (N_20431,N_20236,N_20357);
nand U20432 (N_20432,N_20265,N_20350);
xor U20433 (N_20433,N_20219,N_20260);
nor U20434 (N_20434,N_20202,N_20355);
nand U20435 (N_20435,N_20381,N_20389);
nor U20436 (N_20436,N_20374,N_20262);
nor U20437 (N_20437,N_20239,N_20336);
and U20438 (N_20438,N_20380,N_20330);
and U20439 (N_20439,N_20217,N_20373);
and U20440 (N_20440,N_20386,N_20352);
xnor U20441 (N_20441,N_20215,N_20245);
xnor U20442 (N_20442,N_20295,N_20235);
nand U20443 (N_20443,N_20255,N_20308);
or U20444 (N_20444,N_20383,N_20240);
and U20445 (N_20445,N_20302,N_20231);
and U20446 (N_20446,N_20375,N_20382);
and U20447 (N_20447,N_20356,N_20247);
nor U20448 (N_20448,N_20315,N_20278);
and U20449 (N_20449,N_20252,N_20238);
or U20450 (N_20450,N_20335,N_20226);
or U20451 (N_20451,N_20206,N_20251);
nand U20452 (N_20452,N_20393,N_20264);
or U20453 (N_20453,N_20304,N_20267);
nor U20454 (N_20454,N_20339,N_20385);
nor U20455 (N_20455,N_20326,N_20305);
or U20456 (N_20456,N_20313,N_20301);
xor U20457 (N_20457,N_20281,N_20390);
and U20458 (N_20458,N_20216,N_20276);
nor U20459 (N_20459,N_20307,N_20391);
xnor U20460 (N_20460,N_20358,N_20332);
xor U20461 (N_20461,N_20254,N_20324);
xnor U20462 (N_20462,N_20204,N_20354);
nor U20463 (N_20463,N_20345,N_20211);
nor U20464 (N_20464,N_20377,N_20233);
or U20465 (N_20465,N_20234,N_20333);
xor U20466 (N_20466,N_20261,N_20398);
and U20467 (N_20467,N_20325,N_20244);
nand U20468 (N_20468,N_20212,N_20316);
nand U20469 (N_20469,N_20241,N_20272);
nand U20470 (N_20470,N_20317,N_20222);
nand U20471 (N_20471,N_20399,N_20337);
nand U20472 (N_20472,N_20209,N_20327);
or U20473 (N_20473,N_20227,N_20208);
nor U20474 (N_20474,N_20334,N_20294);
nand U20475 (N_20475,N_20279,N_20274);
nor U20476 (N_20476,N_20283,N_20362);
xnor U20477 (N_20477,N_20397,N_20282);
and U20478 (N_20478,N_20290,N_20280);
xor U20479 (N_20479,N_20387,N_20312);
or U20480 (N_20480,N_20321,N_20379);
nand U20481 (N_20481,N_20395,N_20284);
nand U20482 (N_20482,N_20201,N_20253);
nand U20483 (N_20483,N_20289,N_20394);
nand U20484 (N_20484,N_20228,N_20353);
nand U20485 (N_20485,N_20270,N_20299);
xor U20486 (N_20486,N_20257,N_20322);
or U20487 (N_20487,N_20388,N_20346);
nand U20488 (N_20488,N_20263,N_20293);
nor U20489 (N_20489,N_20372,N_20367);
or U20490 (N_20490,N_20396,N_20360);
and U20491 (N_20491,N_20359,N_20309);
or U20492 (N_20492,N_20246,N_20266);
and U20493 (N_20493,N_20351,N_20364);
and U20494 (N_20494,N_20378,N_20361);
nand U20495 (N_20495,N_20340,N_20221);
or U20496 (N_20496,N_20225,N_20338);
and U20497 (N_20497,N_20205,N_20311);
and U20498 (N_20498,N_20220,N_20285);
xor U20499 (N_20499,N_20203,N_20368);
xnor U20500 (N_20500,N_20228,N_20209);
xor U20501 (N_20501,N_20219,N_20354);
xor U20502 (N_20502,N_20389,N_20203);
nor U20503 (N_20503,N_20308,N_20390);
nor U20504 (N_20504,N_20313,N_20249);
nor U20505 (N_20505,N_20275,N_20234);
and U20506 (N_20506,N_20328,N_20256);
and U20507 (N_20507,N_20241,N_20291);
nor U20508 (N_20508,N_20280,N_20353);
nand U20509 (N_20509,N_20232,N_20326);
or U20510 (N_20510,N_20322,N_20371);
or U20511 (N_20511,N_20224,N_20303);
nor U20512 (N_20512,N_20315,N_20280);
xor U20513 (N_20513,N_20310,N_20333);
nor U20514 (N_20514,N_20357,N_20350);
nand U20515 (N_20515,N_20263,N_20285);
nand U20516 (N_20516,N_20380,N_20332);
nand U20517 (N_20517,N_20265,N_20399);
nor U20518 (N_20518,N_20255,N_20298);
nand U20519 (N_20519,N_20269,N_20382);
and U20520 (N_20520,N_20316,N_20311);
and U20521 (N_20521,N_20362,N_20301);
xnor U20522 (N_20522,N_20319,N_20385);
xnor U20523 (N_20523,N_20293,N_20246);
and U20524 (N_20524,N_20356,N_20282);
nor U20525 (N_20525,N_20351,N_20310);
xor U20526 (N_20526,N_20272,N_20334);
xnor U20527 (N_20527,N_20248,N_20373);
xor U20528 (N_20528,N_20302,N_20219);
or U20529 (N_20529,N_20368,N_20313);
xor U20530 (N_20530,N_20380,N_20321);
nand U20531 (N_20531,N_20395,N_20387);
xor U20532 (N_20532,N_20358,N_20250);
nand U20533 (N_20533,N_20201,N_20298);
nor U20534 (N_20534,N_20345,N_20214);
and U20535 (N_20535,N_20323,N_20304);
xnor U20536 (N_20536,N_20221,N_20355);
xnor U20537 (N_20537,N_20293,N_20265);
nand U20538 (N_20538,N_20210,N_20218);
and U20539 (N_20539,N_20316,N_20250);
xnor U20540 (N_20540,N_20275,N_20291);
xor U20541 (N_20541,N_20361,N_20347);
nand U20542 (N_20542,N_20267,N_20337);
or U20543 (N_20543,N_20215,N_20344);
nor U20544 (N_20544,N_20200,N_20208);
or U20545 (N_20545,N_20314,N_20392);
nand U20546 (N_20546,N_20267,N_20212);
nand U20547 (N_20547,N_20360,N_20210);
or U20548 (N_20548,N_20323,N_20288);
nand U20549 (N_20549,N_20336,N_20241);
nand U20550 (N_20550,N_20351,N_20253);
nor U20551 (N_20551,N_20296,N_20310);
and U20552 (N_20552,N_20292,N_20204);
or U20553 (N_20553,N_20348,N_20270);
xor U20554 (N_20554,N_20394,N_20307);
nand U20555 (N_20555,N_20288,N_20242);
nor U20556 (N_20556,N_20260,N_20302);
xnor U20557 (N_20557,N_20211,N_20337);
nor U20558 (N_20558,N_20350,N_20393);
xnor U20559 (N_20559,N_20339,N_20211);
nand U20560 (N_20560,N_20358,N_20270);
nand U20561 (N_20561,N_20221,N_20210);
nand U20562 (N_20562,N_20211,N_20274);
xor U20563 (N_20563,N_20266,N_20233);
nand U20564 (N_20564,N_20206,N_20305);
nor U20565 (N_20565,N_20351,N_20372);
xor U20566 (N_20566,N_20286,N_20393);
nand U20567 (N_20567,N_20388,N_20245);
nand U20568 (N_20568,N_20368,N_20380);
or U20569 (N_20569,N_20204,N_20283);
and U20570 (N_20570,N_20349,N_20351);
xor U20571 (N_20571,N_20277,N_20354);
xor U20572 (N_20572,N_20221,N_20273);
xnor U20573 (N_20573,N_20311,N_20238);
or U20574 (N_20574,N_20285,N_20317);
or U20575 (N_20575,N_20357,N_20239);
or U20576 (N_20576,N_20284,N_20349);
nand U20577 (N_20577,N_20355,N_20241);
nor U20578 (N_20578,N_20284,N_20326);
and U20579 (N_20579,N_20372,N_20278);
nand U20580 (N_20580,N_20258,N_20295);
xor U20581 (N_20581,N_20323,N_20306);
and U20582 (N_20582,N_20398,N_20307);
nand U20583 (N_20583,N_20338,N_20213);
or U20584 (N_20584,N_20247,N_20398);
xor U20585 (N_20585,N_20345,N_20394);
and U20586 (N_20586,N_20296,N_20211);
and U20587 (N_20587,N_20337,N_20253);
xor U20588 (N_20588,N_20336,N_20206);
and U20589 (N_20589,N_20214,N_20213);
or U20590 (N_20590,N_20284,N_20225);
nand U20591 (N_20591,N_20234,N_20200);
or U20592 (N_20592,N_20274,N_20223);
nand U20593 (N_20593,N_20278,N_20251);
and U20594 (N_20594,N_20373,N_20347);
and U20595 (N_20595,N_20341,N_20313);
or U20596 (N_20596,N_20255,N_20381);
or U20597 (N_20597,N_20245,N_20201);
and U20598 (N_20598,N_20279,N_20379);
or U20599 (N_20599,N_20333,N_20396);
or U20600 (N_20600,N_20430,N_20511);
or U20601 (N_20601,N_20539,N_20563);
or U20602 (N_20602,N_20596,N_20433);
xnor U20603 (N_20603,N_20410,N_20400);
or U20604 (N_20604,N_20469,N_20422);
and U20605 (N_20605,N_20488,N_20543);
and U20606 (N_20606,N_20567,N_20444);
xnor U20607 (N_20607,N_20598,N_20440);
and U20608 (N_20608,N_20575,N_20536);
nor U20609 (N_20609,N_20558,N_20416);
or U20610 (N_20610,N_20492,N_20589);
nand U20611 (N_20611,N_20427,N_20428);
nor U20612 (N_20612,N_20419,N_20459);
xor U20613 (N_20613,N_20496,N_20415);
and U20614 (N_20614,N_20445,N_20561);
and U20615 (N_20615,N_20437,N_20557);
or U20616 (N_20616,N_20538,N_20578);
and U20617 (N_20617,N_20541,N_20592);
and U20618 (N_20618,N_20441,N_20546);
xor U20619 (N_20619,N_20485,N_20523);
xor U20620 (N_20620,N_20521,N_20581);
or U20621 (N_20621,N_20443,N_20417);
or U20622 (N_20622,N_20528,N_20436);
or U20623 (N_20623,N_20452,N_20507);
xor U20624 (N_20624,N_20549,N_20510);
nor U20625 (N_20625,N_20401,N_20553);
nand U20626 (N_20626,N_20587,N_20402);
or U20627 (N_20627,N_20503,N_20451);
xor U20628 (N_20628,N_20475,N_20421);
nand U20629 (N_20629,N_20454,N_20411);
or U20630 (N_20630,N_20471,N_20467);
or U20631 (N_20631,N_20499,N_20453);
or U20632 (N_20632,N_20590,N_20569);
or U20633 (N_20633,N_20423,N_20534);
or U20634 (N_20634,N_20464,N_20491);
or U20635 (N_20635,N_20424,N_20431);
nand U20636 (N_20636,N_20479,N_20593);
nor U20637 (N_20637,N_20588,N_20500);
nand U20638 (N_20638,N_20525,N_20474);
or U20639 (N_20639,N_20448,N_20489);
or U20640 (N_20640,N_20458,N_20572);
nand U20641 (N_20641,N_20484,N_20420);
nor U20642 (N_20642,N_20591,N_20520);
xor U20643 (N_20643,N_20403,N_20586);
and U20644 (N_20644,N_20568,N_20442);
nand U20645 (N_20645,N_20514,N_20426);
xnor U20646 (N_20646,N_20527,N_20405);
nand U20647 (N_20647,N_20535,N_20599);
xnor U20648 (N_20648,N_20434,N_20493);
and U20649 (N_20649,N_20466,N_20579);
or U20650 (N_20650,N_20460,N_20574);
or U20651 (N_20651,N_20583,N_20494);
and U20652 (N_20652,N_20495,N_20542);
or U20653 (N_20653,N_20446,N_20513);
nor U20654 (N_20654,N_20515,N_20532);
nor U20655 (N_20655,N_20470,N_20463);
nand U20656 (N_20656,N_20526,N_20449);
xor U20657 (N_20657,N_20425,N_20486);
nor U20658 (N_20658,N_20461,N_20450);
nand U20659 (N_20659,N_20516,N_20435);
nand U20660 (N_20660,N_20522,N_20518);
nor U20661 (N_20661,N_20533,N_20529);
xnor U20662 (N_20662,N_20455,N_20508);
and U20663 (N_20663,N_20597,N_20438);
nand U20664 (N_20664,N_20481,N_20512);
nor U20665 (N_20665,N_20478,N_20555);
nor U20666 (N_20666,N_20480,N_20509);
nand U20667 (N_20667,N_20498,N_20545);
nor U20668 (N_20668,N_20407,N_20559);
nand U20669 (N_20669,N_20432,N_20580);
or U20670 (N_20670,N_20462,N_20406);
or U20671 (N_20671,N_20456,N_20413);
and U20672 (N_20672,N_20560,N_20577);
nor U20673 (N_20673,N_20550,N_20408);
or U20674 (N_20674,N_20473,N_20564);
nor U20675 (N_20675,N_20412,N_20487);
or U20676 (N_20676,N_20504,N_20562);
nor U20677 (N_20677,N_20594,N_20404);
or U20678 (N_20678,N_20570,N_20585);
nor U20679 (N_20679,N_20418,N_20468);
nor U20680 (N_20680,N_20573,N_20531);
nor U20681 (N_20681,N_20490,N_20519);
nor U20682 (N_20682,N_20565,N_20571);
and U20683 (N_20683,N_20439,N_20505);
nand U20684 (N_20684,N_20556,N_20457);
nor U20685 (N_20685,N_20497,N_20566);
and U20686 (N_20686,N_20544,N_20552);
nor U20687 (N_20687,N_20429,N_20548);
and U20688 (N_20688,N_20409,N_20483);
or U20689 (N_20689,N_20501,N_20584);
and U20690 (N_20690,N_20482,N_20517);
or U20691 (N_20691,N_20414,N_20447);
and U20692 (N_20692,N_20530,N_20582);
and U20693 (N_20693,N_20502,N_20595);
or U20694 (N_20694,N_20551,N_20537);
and U20695 (N_20695,N_20540,N_20476);
or U20696 (N_20696,N_20477,N_20472);
or U20697 (N_20697,N_20576,N_20465);
and U20698 (N_20698,N_20524,N_20506);
or U20699 (N_20699,N_20554,N_20547);
nand U20700 (N_20700,N_20591,N_20558);
nor U20701 (N_20701,N_20544,N_20458);
and U20702 (N_20702,N_20567,N_20540);
or U20703 (N_20703,N_20595,N_20427);
nand U20704 (N_20704,N_20405,N_20408);
or U20705 (N_20705,N_20402,N_20433);
xnor U20706 (N_20706,N_20467,N_20451);
nand U20707 (N_20707,N_20564,N_20482);
or U20708 (N_20708,N_20533,N_20420);
xor U20709 (N_20709,N_20463,N_20410);
xnor U20710 (N_20710,N_20521,N_20441);
nand U20711 (N_20711,N_20559,N_20594);
nand U20712 (N_20712,N_20433,N_20540);
or U20713 (N_20713,N_20519,N_20585);
nand U20714 (N_20714,N_20540,N_20411);
nor U20715 (N_20715,N_20425,N_20599);
or U20716 (N_20716,N_20584,N_20556);
nand U20717 (N_20717,N_20532,N_20594);
nor U20718 (N_20718,N_20572,N_20476);
nor U20719 (N_20719,N_20470,N_20500);
nand U20720 (N_20720,N_20536,N_20449);
nand U20721 (N_20721,N_20587,N_20463);
nor U20722 (N_20722,N_20472,N_20496);
or U20723 (N_20723,N_20462,N_20409);
and U20724 (N_20724,N_20500,N_20461);
or U20725 (N_20725,N_20438,N_20432);
nand U20726 (N_20726,N_20569,N_20483);
nor U20727 (N_20727,N_20527,N_20579);
nor U20728 (N_20728,N_20426,N_20468);
nor U20729 (N_20729,N_20550,N_20570);
xor U20730 (N_20730,N_20403,N_20489);
or U20731 (N_20731,N_20423,N_20405);
nor U20732 (N_20732,N_20497,N_20570);
nand U20733 (N_20733,N_20584,N_20555);
nor U20734 (N_20734,N_20496,N_20505);
and U20735 (N_20735,N_20435,N_20482);
or U20736 (N_20736,N_20436,N_20580);
nor U20737 (N_20737,N_20539,N_20577);
nor U20738 (N_20738,N_20596,N_20570);
or U20739 (N_20739,N_20564,N_20419);
nor U20740 (N_20740,N_20421,N_20595);
xnor U20741 (N_20741,N_20403,N_20426);
xnor U20742 (N_20742,N_20444,N_20538);
nor U20743 (N_20743,N_20448,N_20461);
xor U20744 (N_20744,N_20529,N_20566);
nor U20745 (N_20745,N_20408,N_20409);
xor U20746 (N_20746,N_20592,N_20433);
or U20747 (N_20747,N_20528,N_20426);
or U20748 (N_20748,N_20598,N_20411);
xnor U20749 (N_20749,N_20529,N_20477);
nor U20750 (N_20750,N_20514,N_20490);
or U20751 (N_20751,N_20545,N_20513);
nand U20752 (N_20752,N_20418,N_20543);
or U20753 (N_20753,N_20499,N_20594);
and U20754 (N_20754,N_20499,N_20558);
and U20755 (N_20755,N_20576,N_20480);
or U20756 (N_20756,N_20500,N_20498);
nor U20757 (N_20757,N_20536,N_20547);
xnor U20758 (N_20758,N_20422,N_20411);
and U20759 (N_20759,N_20504,N_20454);
nor U20760 (N_20760,N_20591,N_20424);
or U20761 (N_20761,N_20437,N_20408);
and U20762 (N_20762,N_20466,N_20545);
xnor U20763 (N_20763,N_20473,N_20533);
xor U20764 (N_20764,N_20504,N_20475);
xnor U20765 (N_20765,N_20501,N_20544);
and U20766 (N_20766,N_20417,N_20434);
nor U20767 (N_20767,N_20546,N_20577);
and U20768 (N_20768,N_20593,N_20527);
xor U20769 (N_20769,N_20452,N_20569);
and U20770 (N_20770,N_20556,N_20478);
and U20771 (N_20771,N_20463,N_20464);
xnor U20772 (N_20772,N_20454,N_20457);
nor U20773 (N_20773,N_20417,N_20568);
xor U20774 (N_20774,N_20432,N_20566);
and U20775 (N_20775,N_20524,N_20599);
nor U20776 (N_20776,N_20583,N_20511);
xor U20777 (N_20777,N_20456,N_20560);
or U20778 (N_20778,N_20452,N_20582);
and U20779 (N_20779,N_20421,N_20558);
xor U20780 (N_20780,N_20558,N_20593);
and U20781 (N_20781,N_20573,N_20554);
xor U20782 (N_20782,N_20514,N_20575);
xor U20783 (N_20783,N_20546,N_20581);
nand U20784 (N_20784,N_20593,N_20560);
nor U20785 (N_20785,N_20414,N_20583);
nand U20786 (N_20786,N_20449,N_20400);
and U20787 (N_20787,N_20453,N_20448);
nand U20788 (N_20788,N_20557,N_20532);
and U20789 (N_20789,N_20539,N_20417);
and U20790 (N_20790,N_20587,N_20514);
and U20791 (N_20791,N_20498,N_20417);
xor U20792 (N_20792,N_20574,N_20468);
xor U20793 (N_20793,N_20541,N_20479);
nor U20794 (N_20794,N_20464,N_20525);
or U20795 (N_20795,N_20457,N_20478);
and U20796 (N_20796,N_20587,N_20517);
xor U20797 (N_20797,N_20497,N_20513);
and U20798 (N_20798,N_20533,N_20527);
and U20799 (N_20799,N_20445,N_20531);
xnor U20800 (N_20800,N_20623,N_20663);
nand U20801 (N_20801,N_20631,N_20657);
nor U20802 (N_20802,N_20789,N_20673);
nand U20803 (N_20803,N_20772,N_20783);
xor U20804 (N_20804,N_20616,N_20645);
xnor U20805 (N_20805,N_20785,N_20640);
or U20806 (N_20806,N_20709,N_20672);
nor U20807 (N_20807,N_20792,N_20749);
and U20808 (N_20808,N_20779,N_20681);
xnor U20809 (N_20809,N_20702,N_20771);
or U20810 (N_20810,N_20786,N_20793);
xnor U20811 (N_20811,N_20668,N_20740);
and U20812 (N_20812,N_20676,N_20731);
xnor U20813 (N_20813,N_20797,N_20699);
nor U20814 (N_20814,N_20670,N_20647);
nor U20815 (N_20815,N_20698,N_20764);
xnor U20816 (N_20816,N_20794,N_20608);
and U20817 (N_20817,N_20648,N_20653);
nor U20818 (N_20818,N_20644,N_20639);
and U20819 (N_20819,N_20715,N_20742);
nor U20820 (N_20820,N_20726,N_20627);
xnor U20821 (N_20821,N_20674,N_20641);
nand U20822 (N_20822,N_20790,N_20739);
or U20823 (N_20823,N_20635,N_20752);
xor U20824 (N_20824,N_20620,N_20705);
and U20825 (N_20825,N_20777,N_20706);
xnor U20826 (N_20826,N_20602,N_20795);
or U20827 (N_20827,N_20666,N_20667);
nor U20828 (N_20828,N_20614,N_20721);
and U20829 (N_20829,N_20680,N_20655);
xnor U20830 (N_20830,N_20691,N_20751);
or U20831 (N_20831,N_20671,N_20708);
or U20832 (N_20832,N_20775,N_20625);
xnor U20833 (N_20833,N_20665,N_20651);
and U20834 (N_20834,N_20615,N_20610);
xnor U20835 (N_20835,N_20688,N_20707);
nor U20836 (N_20836,N_20601,N_20609);
and U20837 (N_20837,N_20778,N_20743);
and U20838 (N_20838,N_20662,N_20661);
nor U20839 (N_20839,N_20768,N_20745);
nor U20840 (N_20840,N_20711,N_20788);
nand U20841 (N_20841,N_20619,N_20798);
and U20842 (N_20842,N_20762,N_20652);
or U20843 (N_20843,N_20622,N_20738);
nor U20844 (N_20844,N_20679,N_20678);
xor U20845 (N_20845,N_20704,N_20780);
nor U20846 (N_20846,N_20677,N_20659);
and U20847 (N_20847,N_20696,N_20643);
xnor U20848 (N_20848,N_20621,N_20741);
xor U20849 (N_20849,N_20729,N_20730);
and U20850 (N_20850,N_20685,N_20710);
nand U20851 (N_20851,N_20719,N_20763);
or U20852 (N_20852,N_20753,N_20720);
or U20853 (N_20853,N_20723,N_20716);
xnor U20854 (N_20854,N_20755,N_20646);
or U20855 (N_20855,N_20660,N_20791);
or U20856 (N_20856,N_20747,N_20724);
or U20857 (N_20857,N_20617,N_20628);
nor U20858 (N_20858,N_20611,N_20634);
nor U20859 (N_20859,N_20769,N_20746);
nor U20860 (N_20860,N_20612,N_20733);
xnor U20861 (N_20861,N_20656,N_20664);
and U20862 (N_20862,N_20757,N_20748);
or U20863 (N_20863,N_20694,N_20682);
nand U20864 (N_20864,N_20781,N_20613);
or U20865 (N_20865,N_20796,N_20692);
and U20866 (N_20866,N_20630,N_20776);
xnor U20867 (N_20867,N_20684,N_20606);
and U20868 (N_20868,N_20759,N_20600);
nand U20869 (N_20869,N_20675,N_20799);
nand U20870 (N_20870,N_20722,N_20744);
xnor U20871 (N_20871,N_20618,N_20642);
and U20872 (N_20872,N_20767,N_20638);
nor U20873 (N_20873,N_20603,N_20633);
and U20874 (N_20874,N_20787,N_20725);
nand U20875 (N_20875,N_20649,N_20784);
or U20876 (N_20876,N_20736,N_20607);
xnor U20877 (N_20877,N_20605,N_20756);
and U20878 (N_20878,N_20773,N_20650);
and U20879 (N_20879,N_20687,N_20782);
xor U20880 (N_20880,N_20750,N_20712);
nand U20881 (N_20881,N_20701,N_20713);
and U20882 (N_20882,N_20765,N_20629);
and U20883 (N_20883,N_20626,N_20636);
nand U20884 (N_20884,N_20718,N_20669);
nor U20885 (N_20885,N_20654,N_20758);
nor U20886 (N_20886,N_20737,N_20658);
or U20887 (N_20887,N_20766,N_20632);
nand U20888 (N_20888,N_20760,N_20761);
nor U20889 (N_20889,N_20604,N_20732);
and U20890 (N_20890,N_20689,N_20686);
nand U20891 (N_20891,N_20770,N_20703);
nor U20892 (N_20892,N_20624,N_20695);
or U20893 (N_20893,N_20734,N_20683);
nor U20894 (N_20894,N_20754,N_20637);
nor U20895 (N_20895,N_20714,N_20700);
nor U20896 (N_20896,N_20717,N_20697);
xnor U20897 (N_20897,N_20735,N_20727);
and U20898 (N_20898,N_20693,N_20774);
xor U20899 (N_20899,N_20690,N_20728);
nor U20900 (N_20900,N_20733,N_20753);
nor U20901 (N_20901,N_20602,N_20679);
or U20902 (N_20902,N_20659,N_20607);
nand U20903 (N_20903,N_20737,N_20636);
nor U20904 (N_20904,N_20620,N_20644);
nor U20905 (N_20905,N_20736,N_20725);
and U20906 (N_20906,N_20738,N_20733);
or U20907 (N_20907,N_20759,N_20793);
xnor U20908 (N_20908,N_20747,N_20709);
or U20909 (N_20909,N_20642,N_20739);
and U20910 (N_20910,N_20720,N_20733);
nor U20911 (N_20911,N_20647,N_20720);
or U20912 (N_20912,N_20653,N_20705);
nand U20913 (N_20913,N_20699,N_20723);
nand U20914 (N_20914,N_20621,N_20757);
nor U20915 (N_20915,N_20629,N_20780);
or U20916 (N_20916,N_20734,N_20702);
nand U20917 (N_20917,N_20742,N_20768);
nor U20918 (N_20918,N_20730,N_20653);
xnor U20919 (N_20919,N_20733,N_20747);
xnor U20920 (N_20920,N_20767,N_20739);
nand U20921 (N_20921,N_20651,N_20629);
nor U20922 (N_20922,N_20649,N_20644);
nand U20923 (N_20923,N_20625,N_20764);
xnor U20924 (N_20924,N_20772,N_20660);
nand U20925 (N_20925,N_20715,N_20676);
xor U20926 (N_20926,N_20664,N_20602);
and U20927 (N_20927,N_20747,N_20632);
nor U20928 (N_20928,N_20751,N_20622);
nor U20929 (N_20929,N_20651,N_20603);
or U20930 (N_20930,N_20707,N_20695);
xnor U20931 (N_20931,N_20766,N_20684);
nand U20932 (N_20932,N_20767,N_20628);
nor U20933 (N_20933,N_20664,N_20642);
nor U20934 (N_20934,N_20778,N_20618);
nor U20935 (N_20935,N_20628,N_20763);
xor U20936 (N_20936,N_20775,N_20724);
and U20937 (N_20937,N_20761,N_20686);
nor U20938 (N_20938,N_20669,N_20640);
xor U20939 (N_20939,N_20735,N_20610);
or U20940 (N_20940,N_20720,N_20649);
xnor U20941 (N_20941,N_20628,N_20758);
nor U20942 (N_20942,N_20754,N_20641);
nand U20943 (N_20943,N_20723,N_20776);
nor U20944 (N_20944,N_20684,N_20713);
nand U20945 (N_20945,N_20797,N_20771);
or U20946 (N_20946,N_20633,N_20728);
and U20947 (N_20947,N_20720,N_20786);
nand U20948 (N_20948,N_20686,N_20667);
or U20949 (N_20949,N_20712,N_20788);
nand U20950 (N_20950,N_20798,N_20673);
nand U20951 (N_20951,N_20627,N_20610);
xor U20952 (N_20952,N_20731,N_20613);
or U20953 (N_20953,N_20610,N_20717);
xnor U20954 (N_20954,N_20613,N_20643);
or U20955 (N_20955,N_20616,N_20737);
nor U20956 (N_20956,N_20748,N_20621);
xnor U20957 (N_20957,N_20716,N_20706);
nor U20958 (N_20958,N_20610,N_20787);
nor U20959 (N_20959,N_20672,N_20707);
or U20960 (N_20960,N_20758,N_20601);
nand U20961 (N_20961,N_20691,N_20684);
and U20962 (N_20962,N_20728,N_20622);
xor U20963 (N_20963,N_20771,N_20793);
nor U20964 (N_20964,N_20663,N_20602);
and U20965 (N_20965,N_20666,N_20659);
or U20966 (N_20966,N_20719,N_20640);
or U20967 (N_20967,N_20634,N_20749);
or U20968 (N_20968,N_20773,N_20754);
nand U20969 (N_20969,N_20649,N_20663);
or U20970 (N_20970,N_20698,N_20741);
nor U20971 (N_20971,N_20781,N_20784);
or U20972 (N_20972,N_20625,N_20770);
nand U20973 (N_20973,N_20753,N_20758);
nor U20974 (N_20974,N_20660,N_20707);
nand U20975 (N_20975,N_20646,N_20750);
xor U20976 (N_20976,N_20666,N_20782);
nand U20977 (N_20977,N_20759,N_20616);
or U20978 (N_20978,N_20605,N_20723);
nand U20979 (N_20979,N_20735,N_20649);
and U20980 (N_20980,N_20719,N_20710);
nor U20981 (N_20981,N_20762,N_20653);
nor U20982 (N_20982,N_20710,N_20627);
and U20983 (N_20983,N_20684,N_20611);
nor U20984 (N_20984,N_20702,N_20615);
and U20985 (N_20985,N_20662,N_20606);
nor U20986 (N_20986,N_20651,N_20735);
and U20987 (N_20987,N_20732,N_20602);
and U20988 (N_20988,N_20696,N_20738);
and U20989 (N_20989,N_20796,N_20642);
and U20990 (N_20990,N_20735,N_20631);
xnor U20991 (N_20991,N_20742,N_20624);
or U20992 (N_20992,N_20729,N_20621);
or U20993 (N_20993,N_20633,N_20699);
xor U20994 (N_20994,N_20673,N_20732);
xor U20995 (N_20995,N_20742,N_20776);
nand U20996 (N_20996,N_20793,N_20615);
and U20997 (N_20997,N_20795,N_20735);
and U20998 (N_20998,N_20778,N_20648);
or U20999 (N_20999,N_20728,N_20737);
nor U21000 (N_21000,N_20882,N_20963);
and U21001 (N_21001,N_20931,N_20807);
nor U21002 (N_21002,N_20809,N_20964);
xnor U21003 (N_21003,N_20880,N_20858);
nor U21004 (N_21004,N_20961,N_20924);
or U21005 (N_21005,N_20861,N_20838);
or U21006 (N_21006,N_20958,N_20933);
and U21007 (N_21007,N_20881,N_20935);
xor U21008 (N_21008,N_20986,N_20821);
nor U21009 (N_21009,N_20818,N_20955);
or U21010 (N_21010,N_20890,N_20868);
nand U21011 (N_21011,N_20857,N_20817);
nor U21012 (N_21012,N_20897,N_20895);
nor U21013 (N_21013,N_20984,N_20810);
xnor U21014 (N_21014,N_20846,N_20912);
nand U21015 (N_21015,N_20865,N_20878);
nand U21016 (N_21016,N_20820,N_20854);
or U21017 (N_21017,N_20979,N_20823);
xnor U21018 (N_21018,N_20939,N_20938);
or U21019 (N_21019,N_20894,N_20937);
and U21020 (N_21020,N_20951,N_20953);
and U21021 (N_21021,N_20903,N_20833);
nor U21022 (N_21022,N_20896,N_20832);
and U21023 (N_21023,N_20994,N_20981);
nand U21024 (N_21024,N_20972,N_20826);
nand U21025 (N_21025,N_20926,N_20987);
and U21026 (N_21026,N_20840,N_20869);
nor U21027 (N_21027,N_20872,N_20891);
nor U21028 (N_21028,N_20803,N_20808);
nand U21029 (N_21029,N_20847,N_20804);
and U21030 (N_21030,N_20813,N_20916);
xor U21031 (N_21031,N_20980,N_20806);
nor U21032 (N_21032,N_20900,N_20998);
nor U21033 (N_21033,N_20862,N_20859);
or U21034 (N_21034,N_20919,N_20936);
nand U21035 (N_21035,N_20814,N_20829);
and U21036 (N_21036,N_20822,N_20956);
xnor U21037 (N_21037,N_20883,N_20876);
and U21038 (N_21038,N_20929,N_20834);
or U21039 (N_21039,N_20989,N_20904);
or U21040 (N_21040,N_20921,N_20949);
nand U21041 (N_21041,N_20856,N_20850);
xnor U21042 (N_21042,N_20928,N_20874);
nor U21043 (N_21043,N_20837,N_20830);
or U21044 (N_21044,N_20948,N_20892);
nand U21045 (N_21045,N_20879,N_20932);
xnor U21046 (N_21046,N_20993,N_20884);
nand U21047 (N_21047,N_20934,N_20811);
nand U21048 (N_21048,N_20995,N_20920);
xor U21049 (N_21049,N_20898,N_20970);
nand U21050 (N_21050,N_20950,N_20971);
xor U21051 (N_21051,N_20819,N_20905);
and U21052 (N_21052,N_20852,N_20901);
or U21053 (N_21053,N_20923,N_20836);
xor U21054 (N_21054,N_20845,N_20990);
nor U21055 (N_21055,N_20983,N_20805);
xnor U21056 (N_21056,N_20875,N_20962);
nand U21057 (N_21057,N_20812,N_20801);
or U21058 (N_21058,N_20855,N_20841);
and U21059 (N_21059,N_20988,N_20902);
nand U21060 (N_21060,N_20945,N_20952);
and U21061 (N_21061,N_20835,N_20968);
xnor U21062 (N_21062,N_20886,N_20888);
nor U21063 (N_21063,N_20844,N_20839);
nor U21064 (N_21064,N_20992,N_20893);
and U21065 (N_21065,N_20967,N_20915);
and U21066 (N_21066,N_20885,N_20960);
and U21067 (N_21067,N_20969,N_20918);
nand U21068 (N_21068,N_20991,N_20975);
nand U21069 (N_21069,N_20870,N_20940);
and U21070 (N_21070,N_20899,N_20867);
or U21071 (N_21071,N_20873,N_20907);
or U21072 (N_21072,N_20906,N_20978);
nand U21073 (N_21073,N_20941,N_20911);
nand U21074 (N_21074,N_20831,N_20871);
nor U21075 (N_21075,N_20843,N_20877);
and U21076 (N_21076,N_20889,N_20944);
or U21077 (N_21077,N_20913,N_20974);
nor U21078 (N_21078,N_20909,N_20947);
or U21079 (N_21079,N_20942,N_20977);
and U21080 (N_21080,N_20828,N_20914);
or U21081 (N_21081,N_20946,N_20849);
xor U21082 (N_21082,N_20997,N_20800);
or U21083 (N_21083,N_20853,N_20908);
or U21084 (N_21084,N_20917,N_20866);
and U21085 (N_21085,N_20860,N_20910);
xnor U21086 (N_21086,N_20976,N_20851);
and U21087 (N_21087,N_20965,N_20887);
and U21088 (N_21088,N_20954,N_20943);
nand U21089 (N_21089,N_20816,N_20827);
nor U21090 (N_21090,N_20815,N_20802);
nor U21091 (N_21091,N_20864,N_20922);
nor U21092 (N_21092,N_20927,N_20842);
and U21093 (N_21093,N_20930,N_20959);
nor U21094 (N_21094,N_20999,N_20966);
xnor U21095 (N_21095,N_20824,N_20848);
or U21096 (N_21096,N_20825,N_20925);
xor U21097 (N_21097,N_20982,N_20957);
or U21098 (N_21098,N_20985,N_20863);
or U21099 (N_21099,N_20973,N_20996);
and U21100 (N_21100,N_20937,N_20833);
nand U21101 (N_21101,N_20821,N_20906);
xnor U21102 (N_21102,N_20960,N_20929);
and U21103 (N_21103,N_20835,N_20975);
or U21104 (N_21104,N_20821,N_20996);
or U21105 (N_21105,N_20979,N_20834);
nor U21106 (N_21106,N_20820,N_20800);
nand U21107 (N_21107,N_20898,N_20964);
xnor U21108 (N_21108,N_20882,N_20872);
or U21109 (N_21109,N_20994,N_20849);
xnor U21110 (N_21110,N_20823,N_20836);
or U21111 (N_21111,N_20841,N_20952);
nand U21112 (N_21112,N_20888,N_20907);
nor U21113 (N_21113,N_20925,N_20814);
nor U21114 (N_21114,N_20987,N_20905);
nor U21115 (N_21115,N_20971,N_20977);
xnor U21116 (N_21116,N_20887,N_20834);
xnor U21117 (N_21117,N_20973,N_20910);
nor U21118 (N_21118,N_20911,N_20880);
or U21119 (N_21119,N_20907,N_20849);
nor U21120 (N_21120,N_20806,N_20897);
and U21121 (N_21121,N_20948,N_20814);
nand U21122 (N_21122,N_20836,N_20905);
nand U21123 (N_21123,N_20878,N_20892);
nor U21124 (N_21124,N_20998,N_20820);
and U21125 (N_21125,N_20878,N_20914);
xor U21126 (N_21126,N_20967,N_20976);
xnor U21127 (N_21127,N_20843,N_20827);
nand U21128 (N_21128,N_20822,N_20889);
nor U21129 (N_21129,N_20936,N_20818);
nor U21130 (N_21130,N_20932,N_20998);
and U21131 (N_21131,N_20801,N_20861);
or U21132 (N_21132,N_20852,N_20837);
xor U21133 (N_21133,N_20909,N_20977);
nor U21134 (N_21134,N_20942,N_20897);
nand U21135 (N_21135,N_20821,N_20938);
xnor U21136 (N_21136,N_20978,N_20981);
nor U21137 (N_21137,N_20852,N_20926);
and U21138 (N_21138,N_20981,N_20925);
xnor U21139 (N_21139,N_20812,N_20846);
or U21140 (N_21140,N_20846,N_20897);
or U21141 (N_21141,N_20866,N_20888);
nor U21142 (N_21142,N_20821,N_20990);
nand U21143 (N_21143,N_20970,N_20850);
nor U21144 (N_21144,N_20972,N_20843);
or U21145 (N_21145,N_20994,N_20801);
and U21146 (N_21146,N_20802,N_20848);
xor U21147 (N_21147,N_20934,N_20851);
xnor U21148 (N_21148,N_20961,N_20829);
nor U21149 (N_21149,N_20827,N_20857);
and U21150 (N_21150,N_20844,N_20906);
nor U21151 (N_21151,N_20982,N_20973);
nor U21152 (N_21152,N_20879,N_20842);
xnor U21153 (N_21153,N_20937,N_20848);
nor U21154 (N_21154,N_20989,N_20915);
nand U21155 (N_21155,N_20974,N_20844);
nand U21156 (N_21156,N_20948,N_20928);
nor U21157 (N_21157,N_20969,N_20947);
or U21158 (N_21158,N_20905,N_20931);
and U21159 (N_21159,N_20870,N_20975);
or U21160 (N_21160,N_20891,N_20958);
and U21161 (N_21161,N_20807,N_20971);
or U21162 (N_21162,N_20862,N_20882);
xor U21163 (N_21163,N_20843,N_20977);
nand U21164 (N_21164,N_20998,N_20893);
nor U21165 (N_21165,N_20873,N_20910);
nor U21166 (N_21166,N_20886,N_20953);
nand U21167 (N_21167,N_20811,N_20985);
nand U21168 (N_21168,N_20814,N_20939);
nand U21169 (N_21169,N_20828,N_20912);
nor U21170 (N_21170,N_20912,N_20833);
or U21171 (N_21171,N_20836,N_20961);
nand U21172 (N_21172,N_20872,N_20972);
nand U21173 (N_21173,N_20885,N_20906);
nor U21174 (N_21174,N_20999,N_20822);
nand U21175 (N_21175,N_20865,N_20954);
xor U21176 (N_21176,N_20911,N_20853);
nand U21177 (N_21177,N_20926,N_20920);
xor U21178 (N_21178,N_20947,N_20900);
nor U21179 (N_21179,N_20860,N_20838);
or U21180 (N_21180,N_20931,N_20993);
and U21181 (N_21181,N_20803,N_20958);
or U21182 (N_21182,N_20929,N_20987);
or U21183 (N_21183,N_20876,N_20892);
and U21184 (N_21184,N_20916,N_20957);
xnor U21185 (N_21185,N_20837,N_20868);
xnor U21186 (N_21186,N_20988,N_20961);
xor U21187 (N_21187,N_20880,N_20997);
and U21188 (N_21188,N_20816,N_20924);
nand U21189 (N_21189,N_20841,N_20866);
and U21190 (N_21190,N_20828,N_20959);
nor U21191 (N_21191,N_20852,N_20851);
nor U21192 (N_21192,N_20906,N_20904);
and U21193 (N_21193,N_20827,N_20866);
and U21194 (N_21194,N_20956,N_20877);
nand U21195 (N_21195,N_20880,N_20923);
nor U21196 (N_21196,N_20993,N_20871);
nand U21197 (N_21197,N_20944,N_20858);
nor U21198 (N_21198,N_20899,N_20858);
and U21199 (N_21199,N_20809,N_20931);
xor U21200 (N_21200,N_21107,N_21034);
nand U21201 (N_21201,N_21036,N_21105);
xor U21202 (N_21202,N_21148,N_21160);
or U21203 (N_21203,N_21101,N_21018);
or U21204 (N_21204,N_21130,N_21135);
xnor U21205 (N_21205,N_21067,N_21031);
xor U21206 (N_21206,N_21080,N_21171);
or U21207 (N_21207,N_21129,N_21089);
nand U21208 (N_21208,N_21045,N_21185);
xor U21209 (N_21209,N_21112,N_21024);
nor U21210 (N_21210,N_21058,N_21143);
nand U21211 (N_21211,N_21104,N_21139);
or U21212 (N_21212,N_21108,N_21082);
xor U21213 (N_21213,N_21153,N_21176);
and U21214 (N_21214,N_21035,N_21057);
or U21215 (N_21215,N_21099,N_21137);
and U21216 (N_21216,N_21109,N_21020);
nor U21217 (N_21217,N_21144,N_21097);
or U21218 (N_21218,N_21198,N_21116);
xnor U21219 (N_21219,N_21155,N_21103);
xnor U21220 (N_21220,N_21170,N_21190);
nor U21221 (N_21221,N_21021,N_21147);
or U21222 (N_21222,N_21124,N_21004);
or U21223 (N_21223,N_21092,N_21076);
xnor U21224 (N_21224,N_21118,N_21110);
xor U21225 (N_21225,N_21027,N_21093);
nor U21226 (N_21226,N_21111,N_21022);
or U21227 (N_21227,N_21085,N_21043);
xor U21228 (N_21228,N_21166,N_21090);
or U21229 (N_21229,N_21011,N_21182);
nand U21230 (N_21230,N_21046,N_21158);
nand U21231 (N_21231,N_21087,N_21121);
or U21232 (N_21232,N_21049,N_21125);
nand U21233 (N_21233,N_21019,N_21029);
and U21234 (N_21234,N_21005,N_21002);
nor U21235 (N_21235,N_21042,N_21047);
nand U21236 (N_21236,N_21123,N_21165);
xor U21237 (N_21237,N_21113,N_21075);
xnor U21238 (N_21238,N_21114,N_21007);
or U21239 (N_21239,N_21079,N_21181);
and U21240 (N_21240,N_21056,N_21050);
and U21241 (N_21241,N_21066,N_21194);
nand U21242 (N_21242,N_21064,N_21174);
or U21243 (N_21243,N_21126,N_21167);
or U21244 (N_21244,N_21017,N_21122);
xor U21245 (N_21245,N_21133,N_21052);
and U21246 (N_21246,N_21177,N_21175);
and U21247 (N_21247,N_21070,N_21154);
nor U21248 (N_21248,N_21168,N_21051);
nor U21249 (N_21249,N_21159,N_21040);
nor U21250 (N_21250,N_21078,N_21131);
nand U21251 (N_21251,N_21119,N_21013);
nand U21252 (N_21252,N_21033,N_21138);
or U21253 (N_21253,N_21014,N_21161);
nor U21254 (N_21254,N_21003,N_21074);
and U21255 (N_21255,N_21163,N_21100);
nand U21256 (N_21256,N_21009,N_21142);
nor U21257 (N_21257,N_21102,N_21127);
and U21258 (N_21258,N_21053,N_21150);
xor U21259 (N_21259,N_21012,N_21063);
and U21260 (N_21260,N_21071,N_21032);
or U21261 (N_21261,N_21026,N_21146);
nand U21262 (N_21262,N_21086,N_21088);
xor U21263 (N_21263,N_21059,N_21193);
or U21264 (N_21264,N_21008,N_21072);
or U21265 (N_21265,N_21096,N_21023);
or U21266 (N_21266,N_21081,N_21179);
or U21267 (N_21267,N_21128,N_21197);
or U21268 (N_21268,N_21169,N_21192);
or U21269 (N_21269,N_21001,N_21028);
nor U21270 (N_21270,N_21149,N_21120);
xnor U21271 (N_21271,N_21025,N_21037);
and U21272 (N_21272,N_21164,N_21136);
xnor U21273 (N_21273,N_21196,N_21069);
nor U21274 (N_21274,N_21187,N_21195);
xnor U21275 (N_21275,N_21162,N_21178);
nand U21276 (N_21276,N_21173,N_21186);
nor U21277 (N_21277,N_21073,N_21041);
xor U21278 (N_21278,N_21180,N_21189);
and U21279 (N_21279,N_21134,N_21140);
nand U21280 (N_21280,N_21084,N_21077);
nor U21281 (N_21281,N_21106,N_21055);
nand U21282 (N_21282,N_21183,N_21191);
nor U21283 (N_21283,N_21000,N_21157);
nor U21284 (N_21284,N_21095,N_21068);
or U21285 (N_21285,N_21152,N_21094);
or U21286 (N_21286,N_21117,N_21141);
nor U21287 (N_21287,N_21151,N_21091);
nor U21288 (N_21288,N_21010,N_21145);
and U21289 (N_21289,N_21015,N_21062);
xnor U21290 (N_21290,N_21038,N_21048);
and U21291 (N_21291,N_21065,N_21060);
or U21292 (N_21292,N_21132,N_21115);
xnor U21293 (N_21293,N_21054,N_21172);
nand U21294 (N_21294,N_21188,N_21006);
nor U21295 (N_21295,N_21039,N_21083);
nor U21296 (N_21296,N_21156,N_21061);
nand U21297 (N_21297,N_21199,N_21016);
xor U21298 (N_21298,N_21030,N_21184);
or U21299 (N_21299,N_21098,N_21044);
xor U21300 (N_21300,N_21179,N_21001);
nand U21301 (N_21301,N_21182,N_21198);
xnor U21302 (N_21302,N_21042,N_21112);
or U21303 (N_21303,N_21043,N_21026);
nor U21304 (N_21304,N_21150,N_21197);
nand U21305 (N_21305,N_21172,N_21036);
and U21306 (N_21306,N_21130,N_21196);
nand U21307 (N_21307,N_21185,N_21155);
nand U21308 (N_21308,N_21166,N_21047);
or U21309 (N_21309,N_21143,N_21015);
nand U21310 (N_21310,N_21115,N_21122);
nor U21311 (N_21311,N_21154,N_21165);
nor U21312 (N_21312,N_21198,N_21157);
xor U21313 (N_21313,N_21154,N_21185);
nand U21314 (N_21314,N_21176,N_21184);
nand U21315 (N_21315,N_21028,N_21075);
xor U21316 (N_21316,N_21111,N_21152);
and U21317 (N_21317,N_21147,N_21043);
or U21318 (N_21318,N_21147,N_21115);
nand U21319 (N_21319,N_21170,N_21178);
nand U21320 (N_21320,N_21146,N_21013);
xor U21321 (N_21321,N_21054,N_21175);
and U21322 (N_21322,N_21107,N_21071);
xnor U21323 (N_21323,N_21198,N_21083);
or U21324 (N_21324,N_21038,N_21138);
nor U21325 (N_21325,N_21029,N_21047);
and U21326 (N_21326,N_21106,N_21142);
xnor U21327 (N_21327,N_21092,N_21023);
and U21328 (N_21328,N_21176,N_21084);
and U21329 (N_21329,N_21185,N_21098);
or U21330 (N_21330,N_21016,N_21068);
nor U21331 (N_21331,N_21101,N_21185);
nand U21332 (N_21332,N_21059,N_21097);
nor U21333 (N_21333,N_21140,N_21036);
or U21334 (N_21334,N_21010,N_21088);
nand U21335 (N_21335,N_21199,N_21116);
or U21336 (N_21336,N_21093,N_21062);
or U21337 (N_21337,N_21182,N_21061);
xnor U21338 (N_21338,N_21132,N_21071);
nand U21339 (N_21339,N_21076,N_21064);
and U21340 (N_21340,N_21052,N_21115);
nor U21341 (N_21341,N_21165,N_21037);
and U21342 (N_21342,N_21003,N_21052);
nor U21343 (N_21343,N_21028,N_21187);
xnor U21344 (N_21344,N_21192,N_21098);
nor U21345 (N_21345,N_21030,N_21157);
nor U21346 (N_21346,N_21148,N_21161);
nand U21347 (N_21347,N_21165,N_21068);
and U21348 (N_21348,N_21166,N_21119);
nand U21349 (N_21349,N_21122,N_21195);
and U21350 (N_21350,N_21134,N_21047);
nor U21351 (N_21351,N_21167,N_21035);
and U21352 (N_21352,N_21189,N_21170);
nand U21353 (N_21353,N_21099,N_21157);
xor U21354 (N_21354,N_21130,N_21182);
or U21355 (N_21355,N_21061,N_21110);
nand U21356 (N_21356,N_21072,N_21127);
and U21357 (N_21357,N_21177,N_21017);
and U21358 (N_21358,N_21126,N_21002);
or U21359 (N_21359,N_21094,N_21056);
nor U21360 (N_21360,N_21137,N_21060);
or U21361 (N_21361,N_21014,N_21095);
and U21362 (N_21362,N_21143,N_21170);
xnor U21363 (N_21363,N_21163,N_21020);
and U21364 (N_21364,N_21111,N_21033);
nand U21365 (N_21365,N_21122,N_21194);
and U21366 (N_21366,N_21036,N_21135);
or U21367 (N_21367,N_21142,N_21125);
nor U21368 (N_21368,N_21078,N_21112);
xor U21369 (N_21369,N_21079,N_21020);
or U21370 (N_21370,N_21188,N_21161);
nor U21371 (N_21371,N_21078,N_21156);
or U21372 (N_21372,N_21046,N_21078);
nand U21373 (N_21373,N_21054,N_21098);
or U21374 (N_21374,N_21195,N_21027);
nor U21375 (N_21375,N_21168,N_21042);
xnor U21376 (N_21376,N_21119,N_21185);
nand U21377 (N_21377,N_21198,N_21020);
nand U21378 (N_21378,N_21150,N_21087);
xor U21379 (N_21379,N_21021,N_21034);
nand U21380 (N_21380,N_21084,N_21119);
xnor U21381 (N_21381,N_21035,N_21045);
or U21382 (N_21382,N_21009,N_21030);
and U21383 (N_21383,N_21056,N_21137);
xor U21384 (N_21384,N_21028,N_21076);
xor U21385 (N_21385,N_21070,N_21129);
xnor U21386 (N_21386,N_21009,N_21183);
nor U21387 (N_21387,N_21063,N_21103);
xnor U21388 (N_21388,N_21161,N_21166);
or U21389 (N_21389,N_21137,N_21087);
nor U21390 (N_21390,N_21177,N_21107);
nor U21391 (N_21391,N_21045,N_21098);
or U21392 (N_21392,N_21038,N_21010);
nor U21393 (N_21393,N_21195,N_21001);
nand U21394 (N_21394,N_21144,N_21003);
nand U21395 (N_21395,N_21058,N_21139);
nor U21396 (N_21396,N_21003,N_21059);
nor U21397 (N_21397,N_21137,N_21037);
nor U21398 (N_21398,N_21029,N_21168);
nor U21399 (N_21399,N_21076,N_21131);
and U21400 (N_21400,N_21371,N_21310);
or U21401 (N_21401,N_21282,N_21389);
and U21402 (N_21402,N_21369,N_21252);
xor U21403 (N_21403,N_21388,N_21319);
or U21404 (N_21404,N_21262,N_21358);
xor U21405 (N_21405,N_21368,N_21226);
nand U21406 (N_21406,N_21311,N_21210);
xor U21407 (N_21407,N_21292,N_21268);
nor U21408 (N_21408,N_21378,N_21295);
nand U21409 (N_21409,N_21259,N_21370);
or U21410 (N_21410,N_21318,N_21242);
and U21411 (N_21411,N_21314,N_21263);
and U21412 (N_21412,N_21356,N_21208);
xor U21413 (N_21413,N_21360,N_21216);
and U21414 (N_21414,N_21205,N_21246);
or U21415 (N_21415,N_21331,N_21346);
nand U21416 (N_21416,N_21261,N_21281);
nor U21417 (N_21417,N_21296,N_21219);
nand U21418 (N_21418,N_21313,N_21302);
nand U21419 (N_21419,N_21234,N_21275);
nor U21420 (N_21420,N_21278,N_21238);
nor U21421 (N_21421,N_21345,N_21276);
or U21422 (N_21422,N_21377,N_21309);
or U21423 (N_21423,N_21376,N_21243);
nor U21424 (N_21424,N_21301,N_21227);
or U21425 (N_21425,N_21362,N_21340);
or U21426 (N_21426,N_21273,N_21218);
and U21427 (N_21427,N_21298,N_21339);
nor U21428 (N_21428,N_21260,N_21272);
nor U21429 (N_21429,N_21223,N_21351);
xor U21430 (N_21430,N_21287,N_21332);
nand U21431 (N_21431,N_21220,N_21211);
and U21432 (N_21432,N_21231,N_21250);
nor U21433 (N_21433,N_21303,N_21365);
nor U21434 (N_21434,N_21217,N_21255);
nor U21435 (N_21435,N_21229,N_21321);
or U21436 (N_21436,N_21395,N_21241);
nand U21437 (N_21437,N_21209,N_21341);
and U21438 (N_21438,N_21324,N_21256);
and U21439 (N_21439,N_21290,N_21251);
or U21440 (N_21440,N_21326,N_21240);
xnor U21441 (N_21441,N_21359,N_21233);
nor U21442 (N_21442,N_21304,N_21366);
or U21443 (N_21443,N_21399,N_21285);
and U21444 (N_21444,N_21288,N_21380);
or U21445 (N_21445,N_21397,N_21320);
or U21446 (N_21446,N_21232,N_21271);
xor U21447 (N_21447,N_21327,N_21312);
nor U21448 (N_21448,N_21322,N_21347);
xnor U21449 (N_21449,N_21213,N_21280);
or U21450 (N_21450,N_21387,N_21247);
xnor U21451 (N_21451,N_21283,N_21249);
nor U21452 (N_21452,N_21315,N_21375);
xnor U21453 (N_21453,N_21230,N_21239);
nand U21454 (N_21454,N_21221,N_21350);
xor U21455 (N_21455,N_21386,N_21373);
nand U21456 (N_21456,N_21338,N_21269);
xnor U21457 (N_21457,N_21352,N_21367);
and U21458 (N_21458,N_21294,N_21267);
xor U21459 (N_21459,N_21323,N_21214);
nor U21460 (N_21460,N_21335,N_21307);
and U21461 (N_21461,N_21200,N_21390);
nor U21462 (N_21462,N_21265,N_21382);
or U21463 (N_21463,N_21383,N_21245);
or U21464 (N_21464,N_21353,N_21306);
or U21465 (N_21465,N_21325,N_21206);
and U21466 (N_21466,N_21224,N_21349);
xor U21467 (N_21467,N_21329,N_21244);
or U21468 (N_21468,N_21277,N_21379);
and U21469 (N_21469,N_21279,N_21364);
nor U21470 (N_21470,N_21328,N_21308);
and U21471 (N_21471,N_21330,N_21201);
nand U21472 (N_21472,N_21222,N_21337);
nand U21473 (N_21473,N_21264,N_21385);
xnor U21474 (N_21474,N_21357,N_21336);
or U21475 (N_21475,N_21228,N_21354);
nor U21476 (N_21476,N_21372,N_21284);
nor U21477 (N_21477,N_21253,N_21289);
nand U21478 (N_21478,N_21394,N_21333);
nand U21479 (N_21479,N_21225,N_21235);
nor U21480 (N_21480,N_21305,N_21299);
or U21481 (N_21481,N_21363,N_21202);
nor U21482 (N_21482,N_21266,N_21342);
nor U21483 (N_21483,N_21334,N_21348);
or U21484 (N_21484,N_21291,N_21392);
and U21485 (N_21485,N_21398,N_21286);
or U21486 (N_21486,N_21270,N_21317);
nand U21487 (N_21487,N_21361,N_21215);
xnor U21488 (N_21488,N_21204,N_21343);
nor U21489 (N_21489,N_21254,N_21355);
xor U21490 (N_21490,N_21374,N_21293);
and U21491 (N_21491,N_21248,N_21344);
or U21492 (N_21492,N_21207,N_21258);
nand U21493 (N_21493,N_21237,N_21381);
or U21494 (N_21494,N_21396,N_21300);
nor U21495 (N_21495,N_21384,N_21212);
and U21496 (N_21496,N_21274,N_21391);
xnor U21497 (N_21497,N_21257,N_21316);
nand U21498 (N_21498,N_21203,N_21236);
nand U21499 (N_21499,N_21393,N_21297);
and U21500 (N_21500,N_21391,N_21397);
nand U21501 (N_21501,N_21242,N_21320);
nor U21502 (N_21502,N_21248,N_21220);
nand U21503 (N_21503,N_21379,N_21242);
xor U21504 (N_21504,N_21367,N_21299);
xnor U21505 (N_21505,N_21305,N_21313);
xnor U21506 (N_21506,N_21357,N_21350);
and U21507 (N_21507,N_21395,N_21323);
nand U21508 (N_21508,N_21300,N_21308);
nand U21509 (N_21509,N_21263,N_21319);
or U21510 (N_21510,N_21262,N_21254);
xor U21511 (N_21511,N_21324,N_21372);
xor U21512 (N_21512,N_21206,N_21320);
nor U21513 (N_21513,N_21231,N_21371);
and U21514 (N_21514,N_21305,N_21214);
or U21515 (N_21515,N_21359,N_21398);
nand U21516 (N_21516,N_21314,N_21226);
and U21517 (N_21517,N_21348,N_21200);
nand U21518 (N_21518,N_21214,N_21392);
xnor U21519 (N_21519,N_21250,N_21314);
nor U21520 (N_21520,N_21257,N_21205);
nand U21521 (N_21521,N_21312,N_21381);
and U21522 (N_21522,N_21276,N_21283);
nor U21523 (N_21523,N_21234,N_21240);
nand U21524 (N_21524,N_21248,N_21331);
and U21525 (N_21525,N_21366,N_21247);
nor U21526 (N_21526,N_21274,N_21276);
nor U21527 (N_21527,N_21228,N_21314);
xor U21528 (N_21528,N_21263,N_21244);
and U21529 (N_21529,N_21323,N_21373);
nor U21530 (N_21530,N_21277,N_21327);
nand U21531 (N_21531,N_21237,N_21390);
nand U21532 (N_21532,N_21336,N_21366);
xor U21533 (N_21533,N_21234,N_21394);
or U21534 (N_21534,N_21218,N_21243);
and U21535 (N_21535,N_21395,N_21285);
or U21536 (N_21536,N_21376,N_21285);
xnor U21537 (N_21537,N_21364,N_21204);
and U21538 (N_21538,N_21284,N_21388);
or U21539 (N_21539,N_21293,N_21384);
nor U21540 (N_21540,N_21352,N_21236);
nand U21541 (N_21541,N_21246,N_21207);
nand U21542 (N_21542,N_21341,N_21364);
nand U21543 (N_21543,N_21351,N_21284);
and U21544 (N_21544,N_21273,N_21381);
or U21545 (N_21545,N_21265,N_21261);
nand U21546 (N_21546,N_21334,N_21352);
and U21547 (N_21547,N_21263,N_21385);
and U21548 (N_21548,N_21342,N_21233);
nor U21549 (N_21549,N_21375,N_21347);
and U21550 (N_21550,N_21232,N_21398);
or U21551 (N_21551,N_21241,N_21343);
and U21552 (N_21552,N_21350,N_21325);
nand U21553 (N_21553,N_21396,N_21363);
and U21554 (N_21554,N_21367,N_21235);
nand U21555 (N_21555,N_21248,N_21334);
or U21556 (N_21556,N_21381,N_21244);
nor U21557 (N_21557,N_21258,N_21315);
nand U21558 (N_21558,N_21223,N_21322);
nor U21559 (N_21559,N_21245,N_21399);
nor U21560 (N_21560,N_21313,N_21342);
xnor U21561 (N_21561,N_21329,N_21315);
nand U21562 (N_21562,N_21256,N_21287);
nand U21563 (N_21563,N_21360,N_21341);
or U21564 (N_21564,N_21341,N_21393);
nand U21565 (N_21565,N_21341,N_21374);
or U21566 (N_21566,N_21317,N_21292);
xnor U21567 (N_21567,N_21333,N_21281);
and U21568 (N_21568,N_21354,N_21353);
nand U21569 (N_21569,N_21386,N_21247);
xor U21570 (N_21570,N_21345,N_21390);
and U21571 (N_21571,N_21314,N_21362);
xor U21572 (N_21572,N_21230,N_21371);
nor U21573 (N_21573,N_21216,N_21278);
nand U21574 (N_21574,N_21382,N_21235);
nand U21575 (N_21575,N_21259,N_21373);
nor U21576 (N_21576,N_21211,N_21347);
nor U21577 (N_21577,N_21281,N_21309);
nor U21578 (N_21578,N_21341,N_21310);
nor U21579 (N_21579,N_21322,N_21346);
nor U21580 (N_21580,N_21319,N_21385);
xnor U21581 (N_21581,N_21351,N_21336);
nand U21582 (N_21582,N_21311,N_21376);
or U21583 (N_21583,N_21253,N_21237);
nor U21584 (N_21584,N_21395,N_21281);
nand U21585 (N_21585,N_21329,N_21374);
and U21586 (N_21586,N_21211,N_21331);
xnor U21587 (N_21587,N_21319,N_21240);
or U21588 (N_21588,N_21207,N_21353);
or U21589 (N_21589,N_21264,N_21269);
and U21590 (N_21590,N_21204,N_21385);
and U21591 (N_21591,N_21357,N_21352);
xor U21592 (N_21592,N_21319,N_21223);
nor U21593 (N_21593,N_21388,N_21215);
and U21594 (N_21594,N_21392,N_21318);
and U21595 (N_21595,N_21200,N_21346);
or U21596 (N_21596,N_21306,N_21253);
nand U21597 (N_21597,N_21353,N_21237);
or U21598 (N_21598,N_21351,N_21269);
xnor U21599 (N_21599,N_21289,N_21366);
xor U21600 (N_21600,N_21407,N_21596);
nand U21601 (N_21601,N_21501,N_21569);
nor U21602 (N_21602,N_21576,N_21554);
nor U21603 (N_21603,N_21500,N_21475);
or U21604 (N_21604,N_21541,N_21577);
xnor U21605 (N_21605,N_21545,N_21564);
or U21606 (N_21606,N_21493,N_21486);
xnor U21607 (N_21607,N_21425,N_21424);
nor U21608 (N_21608,N_21597,N_21474);
and U21609 (N_21609,N_21411,N_21444);
and U21610 (N_21610,N_21415,N_21400);
or U21611 (N_21611,N_21506,N_21497);
xor U21612 (N_21612,N_21520,N_21478);
nand U21613 (N_21613,N_21439,N_21409);
xor U21614 (N_21614,N_21448,N_21463);
nand U21615 (N_21615,N_21533,N_21591);
or U21616 (N_21616,N_21530,N_21406);
xnor U21617 (N_21617,N_21588,N_21437);
nor U21618 (N_21618,N_21538,N_21492);
and U21619 (N_21619,N_21494,N_21401);
nand U21620 (N_21620,N_21562,N_21477);
nor U21621 (N_21621,N_21580,N_21540);
and U21622 (N_21622,N_21466,N_21495);
xor U21623 (N_21623,N_21468,N_21485);
nand U21624 (N_21624,N_21547,N_21481);
nor U21625 (N_21625,N_21514,N_21458);
nand U21626 (N_21626,N_21404,N_21574);
xor U21627 (N_21627,N_21402,N_21509);
or U21628 (N_21628,N_21535,N_21452);
xnor U21629 (N_21629,N_21465,N_21594);
xnor U21630 (N_21630,N_21449,N_21410);
xor U21631 (N_21631,N_21542,N_21546);
xnor U21632 (N_21632,N_21421,N_21453);
xor U21633 (N_21633,N_21549,N_21435);
and U21634 (N_21634,N_21440,N_21483);
nand U21635 (N_21635,N_21570,N_21592);
or U21636 (N_21636,N_21460,N_21482);
xor U21637 (N_21637,N_21510,N_21568);
nand U21638 (N_21638,N_21419,N_21584);
nor U21639 (N_21639,N_21445,N_21462);
nor U21640 (N_21640,N_21499,N_21472);
or U21641 (N_21641,N_21505,N_21470);
or U21642 (N_21642,N_21442,N_21422);
or U21643 (N_21643,N_21512,N_21555);
nand U21644 (N_21644,N_21480,N_21525);
nand U21645 (N_21645,N_21586,N_21469);
nand U21646 (N_21646,N_21417,N_21504);
or U21647 (N_21647,N_21456,N_21523);
xor U21648 (N_21648,N_21587,N_21521);
and U21649 (N_21649,N_21551,N_21450);
xor U21650 (N_21650,N_21560,N_21519);
nand U21651 (N_21651,N_21490,N_21461);
nor U21652 (N_21652,N_21516,N_21429);
nor U21653 (N_21653,N_21479,N_21464);
xnor U21654 (N_21654,N_21511,N_21573);
nand U21655 (N_21655,N_21488,N_21590);
and U21656 (N_21656,N_21471,N_21473);
xor U21657 (N_21657,N_21585,N_21572);
nand U21658 (N_21658,N_21503,N_21524);
or U21659 (N_21659,N_21565,N_21476);
or U21660 (N_21660,N_21566,N_21534);
and U21661 (N_21661,N_21518,N_21467);
nand U21662 (N_21662,N_21502,N_21548);
nand U21663 (N_21663,N_21430,N_21438);
or U21664 (N_21664,N_21522,N_21418);
nand U21665 (N_21665,N_21583,N_21526);
or U21666 (N_21666,N_21539,N_21454);
or U21667 (N_21667,N_21552,N_21599);
or U21668 (N_21668,N_21423,N_21558);
xnor U21669 (N_21669,N_21537,N_21544);
or U21670 (N_21670,N_21543,N_21455);
nor U21671 (N_21671,N_21427,N_21527);
or U21672 (N_21672,N_21536,N_21405);
and U21673 (N_21673,N_21428,N_21420);
and U21674 (N_21674,N_21561,N_21559);
nor U21675 (N_21675,N_21431,N_21507);
nand U21676 (N_21676,N_21403,N_21443);
nand U21677 (N_21677,N_21426,N_21434);
and U21678 (N_21678,N_21532,N_21595);
nor U21679 (N_21679,N_21412,N_21557);
or U21680 (N_21680,N_21441,N_21416);
nor U21681 (N_21681,N_21556,N_21487);
xnor U21682 (N_21682,N_21589,N_21579);
nor U21683 (N_21683,N_21498,N_21451);
nand U21684 (N_21684,N_21459,N_21578);
and U21685 (N_21685,N_21489,N_21553);
and U21686 (N_21686,N_21446,N_21457);
and U21687 (N_21687,N_21550,N_21529);
xor U21688 (N_21688,N_21433,N_21528);
nor U21689 (N_21689,N_21513,N_21575);
xnor U21690 (N_21690,N_21571,N_21593);
xor U21691 (N_21691,N_21436,N_21508);
xor U21692 (N_21692,N_21447,N_21598);
or U21693 (N_21693,N_21432,N_21491);
or U21694 (N_21694,N_21413,N_21515);
or U21695 (N_21695,N_21567,N_21531);
nand U21696 (N_21696,N_21496,N_21484);
and U21697 (N_21697,N_21563,N_21582);
or U21698 (N_21698,N_21408,N_21517);
and U21699 (N_21699,N_21414,N_21581);
xnor U21700 (N_21700,N_21544,N_21484);
nand U21701 (N_21701,N_21454,N_21592);
and U21702 (N_21702,N_21436,N_21411);
nand U21703 (N_21703,N_21464,N_21596);
or U21704 (N_21704,N_21435,N_21586);
xor U21705 (N_21705,N_21532,N_21468);
and U21706 (N_21706,N_21594,N_21482);
or U21707 (N_21707,N_21496,N_21512);
nand U21708 (N_21708,N_21560,N_21439);
nand U21709 (N_21709,N_21544,N_21409);
xnor U21710 (N_21710,N_21509,N_21500);
and U21711 (N_21711,N_21534,N_21428);
nand U21712 (N_21712,N_21417,N_21495);
nand U21713 (N_21713,N_21532,N_21543);
nand U21714 (N_21714,N_21469,N_21562);
and U21715 (N_21715,N_21513,N_21415);
nor U21716 (N_21716,N_21519,N_21463);
nor U21717 (N_21717,N_21536,N_21450);
or U21718 (N_21718,N_21515,N_21517);
nand U21719 (N_21719,N_21404,N_21466);
and U21720 (N_21720,N_21401,N_21415);
and U21721 (N_21721,N_21521,N_21579);
or U21722 (N_21722,N_21494,N_21555);
xnor U21723 (N_21723,N_21502,N_21464);
nand U21724 (N_21724,N_21471,N_21579);
xor U21725 (N_21725,N_21466,N_21560);
and U21726 (N_21726,N_21438,N_21586);
xor U21727 (N_21727,N_21551,N_21554);
and U21728 (N_21728,N_21567,N_21468);
and U21729 (N_21729,N_21552,N_21545);
nand U21730 (N_21730,N_21598,N_21534);
or U21731 (N_21731,N_21407,N_21575);
nand U21732 (N_21732,N_21585,N_21428);
or U21733 (N_21733,N_21521,N_21504);
or U21734 (N_21734,N_21592,N_21409);
nand U21735 (N_21735,N_21540,N_21594);
or U21736 (N_21736,N_21513,N_21528);
nor U21737 (N_21737,N_21530,N_21439);
nor U21738 (N_21738,N_21494,N_21508);
xnor U21739 (N_21739,N_21572,N_21587);
or U21740 (N_21740,N_21450,N_21434);
and U21741 (N_21741,N_21434,N_21591);
nand U21742 (N_21742,N_21491,N_21516);
xnor U21743 (N_21743,N_21569,N_21532);
or U21744 (N_21744,N_21458,N_21498);
nand U21745 (N_21745,N_21428,N_21445);
nand U21746 (N_21746,N_21597,N_21402);
nor U21747 (N_21747,N_21471,N_21485);
nor U21748 (N_21748,N_21526,N_21543);
nand U21749 (N_21749,N_21491,N_21587);
xor U21750 (N_21750,N_21403,N_21486);
or U21751 (N_21751,N_21433,N_21417);
nor U21752 (N_21752,N_21494,N_21403);
xnor U21753 (N_21753,N_21505,N_21559);
nand U21754 (N_21754,N_21453,N_21579);
or U21755 (N_21755,N_21457,N_21525);
and U21756 (N_21756,N_21543,N_21582);
xor U21757 (N_21757,N_21550,N_21427);
nand U21758 (N_21758,N_21526,N_21498);
nand U21759 (N_21759,N_21523,N_21473);
xnor U21760 (N_21760,N_21538,N_21559);
nand U21761 (N_21761,N_21436,N_21490);
nand U21762 (N_21762,N_21581,N_21402);
xor U21763 (N_21763,N_21565,N_21457);
xnor U21764 (N_21764,N_21599,N_21517);
nor U21765 (N_21765,N_21546,N_21461);
and U21766 (N_21766,N_21560,N_21419);
nand U21767 (N_21767,N_21480,N_21488);
xnor U21768 (N_21768,N_21430,N_21428);
nand U21769 (N_21769,N_21409,N_21421);
or U21770 (N_21770,N_21407,N_21590);
and U21771 (N_21771,N_21539,N_21584);
nor U21772 (N_21772,N_21510,N_21594);
nand U21773 (N_21773,N_21585,N_21501);
and U21774 (N_21774,N_21507,N_21591);
nand U21775 (N_21775,N_21518,N_21598);
and U21776 (N_21776,N_21592,N_21469);
and U21777 (N_21777,N_21496,N_21405);
and U21778 (N_21778,N_21537,N_21480);
xor U21779 (N_21779,N_21560,N_21561);
nand U21780 (N_21780,N_21469,N_21492);
nor U21781 (N_21781,N_21595,N_21477);
nand U21782 (N_21782,N_21424,N_21509);
or U21783 (N_21783,N_21579,N_21592);
nor U21784 (N_21784,N_21489,N_21483);
and U21785 (N_21785,N_21408,N_21475);
nand U21786 (N_21786,N_21487,N_21488);
and U21787 (N_21787,N_21504,N_21455);
nand U21788 (N_21788,N_21563,N_21537);
nand U21789 (N_21789,N_21541,N_21514);
or U21790 (N_21790,N_21434,N_21473);
nor U21791 (N_21791,N_21504,N_21485);
nand U21792 (N_21792,N_21500,N_21497);
nor U21793 (N_21793,N_21491,N_21599);
xnor U21794 (N_21794,N_21489,N_21401);
nand U21795 (N_21795,N_21441,N_21482);
nor U21796 (N_21796,N_21574,N_21499);
or U21797 (N_21797,N_21544,N_21540);
or U21798 (N_21798,N_21532,N_21596);
or U21799 (N_21799,N_21461,N_21413);
xor U21800 (N_21800,N_21751,N_21630);
nand U21801 (N_21801,N_21662,N_21767);
nor U21802 (N_21802,N_21671,N_21749);
nor U21803 (N_21803,N_21753,N_21648);
nor U21804 (N_21804,N_21719,N_21601);
xnor U21805 (N_21805,N_21620,N_21645);
xor U21806 (N_21806,N_21661,N_21781);
or U21807 (N_21807,N_21738,N_21794);
or U21808 (N_21808,N_21640,N_21747);
or U21809 (N_21809,N_21611,N_21663);
or U21810 (N_21810,N_21652,N_21702);
xnor U21811 (N_21811,N_21780,N_21672);
xor U21812 (N_21812,N_21743,N_21769);
and U21813 (N_21813,N_21618,N_21735);
or U21814 (N_21814,N_21647,N_21690);
and U21815 (N_21815,N_21632,N_21609);
nor U21816 (N_21816,N_21759,N_21750);
nor U21817 (N_21817,N_21772,N_21740);
and U21818 (N_21818,N_21783,N_21797);
or U21819 (N_21819,N_21739,N_21737);
nand U21820 (N_21820,N_21674,N_21606);
nor U21821 (N_21821,N_21777,N_21697);
nor U21822 (N_21822,N_21669,N_21685);
nand U21823 (N_21823,N_21649,N_21733);
nor U21824 (N_21824,N_21614,N_21725);
or U21825 (N_21825,N_21600,N_21720);
nand U21826 (N_21826,N_21605,N_21756);
or U21827 (N_21827,N_21704,N_21604);
and U21828 (N_21828,N_21686,N_21643);
nand U21829 (N_21829,N_21608,N_21754);
and U21830 (N_21830,N_21795,N_21633);
or U21831 (N_21831,N_21658,N_21667);
nand U21832 (N_21832,N_21722,N_21710);
nor U21833 (N_21833,N_21746,N_21634);
and U21834 (N_21834,N_21682,N_21785);
xnor U21835 (N_21835,N_21791,N_21731);
or U21836 (N_21836,N_21761,N_21692);
or U21837 (N_21837,N_21615,N_21617);
nor U21838 (N_21838,N_21745,N_21677);
nor U21839 (N_21839,N_21706,N_21727);
nand U21840 (N_21840,N_21712,N_21639);
xnor U21841 (N_21841,N_21717,N_21748);
or U21842 (N_21842,N_21638,N_21776);
and U21843 (N_21843,N_21689,N_21798);
or U21844 (N_21844,N_21603,N_21721);
or U21845 (N_21845,N_21701,N_21644);
and U21846 (N_21846,N_21724,N_21773);
or U21847 (N_21847,N_21708,N_21679);
and U21848 (N_21848,N_21660,N_21665);
or U21849 (N_21849,N_21709,N_21782);
xnor U21850 (N_21850,N_21616,N_21680);
xor U21851 (N_21851,N_21683,N_21637);
nand U21852 (N_21852,N_21757,N_21651);
xor U21853 (N_21853,N_21625,N_21728);
or U21854 (N_21854,N_21636,N_21755);
nor U21855 (N_21855,N_21778,N_21768);
nand U21856 (N_21856,N_21726,N_21681);
and U21857 (N_21857,N_21742,N_21673);
nand U21858 (N_21858,N_21627,N_21707);
nand U21859 (N_21859,N_21695,N_21734);
and U21860 (N_21860,N_21610,N_21779);
nor U21861 (N_21861,N_21729,N_21602);
xnor U21862 (N_21862,N_21718,N_21657);
or U21863 (N_21863,N_21732,N_21659);
nand U21864 (N_21864,N_21656,N_21675);
xnor U21865 (N_21865,N_21763,N_21796);
nor U21866 (N_21866,N_21622,N_21666);
nand U21867 (N_21867,N_21765,N_21621);
and U21868 (N_21868,N_21786,N_21771);
xor U21869 (N_21869,N_21684,N_21678);
xor U21870 (N_21870,N_21696,N_21770);
xnor U21871 (N_21871,N_21760,N_21799);
or U21872 (N_21872,N_21758,N_21676);
or U21873 (N_21873,N_21793,N_21654);
nor U21874 (N_21874,N_21619,N_21668);
nor U21875 (N_21875,N_21752,N_21653);
nor U21876 (N_21876,N_21766,N_21700);
nor U21877 (N_21877,N_21642,N_21714);
nand U21878 (N_21878,N_21792,N_21705);
or U21879 (N_21879,N_21784,N_21641);
xnor U21880 (N_21880,N_21613,N_21715);
nand U21881 (N_21881,N_21744,N_21713);
or U21882 (N_21882,N_21730,N_21741);
and U21883 (N_21883,N_21762,N_21650);
nand U21884 (N_21884,N_21789,N_21711);
xor U21885 (N_21885,N_21764,N_21703);
xor U21886 (N_21886,N_21687,N_21635);
nand U21887 (N_21887,N_21664,N_21626);
nor U21888 (N_21888,N_21736,N_21624);
and U21889 (N_21889,N_21788,N_21607);
nand U21890 (N_21890,N_21790,N_21691);
and U21891 (N_21891,N_21698,N_21612);
and U21892 (N_21892,N_21774,N_21716);
and U21893 (N_21893,N_21628,N_21775);
or U21894 (N_21894,N_21631,N_21723);
nand U21895 (N_21895,N_21623,N_21699);
or U21896 (N_21896,N_21655,N_21646);
xor U21897 (N_21897,N_21629,N_21688);
xnor U21898 (N_21898,N_21670,N_21694);
nor U21899 (N_21899,N_21787,N_21693);
nand U21900 (N_21900,N_21606,N_21759);
nor U21901 (N_21901,N_21745,N_21696);
xor U21902 (N_21902,N_21619,N_21685);
nand U21903 (N_21903,N_21781,N_21633);
nand U21904 (N_21904,N_21699,N_21652);
nor U21905 (N_21905,N_21685,N_21742);
or U21906 (N_21906,N_21791,N_21612);
nand U21907 (N_21907,N_21783,N_21734);
and U21908 (N_21908,N_21675,N_21717);
and U21909 (N_21909,N_21733,N_21628);
nand U21910 (N_21910,N_21735,N_21660);
and U21911 (N_21911,N_21798,N_21781);
or U21912 (N_21912,N_21766,N_21664);
and U21913 (N_21913,N_21697,N_21778);
nor U21914 (N_21914,N_21657,N_21619);
nand U21915 (N_21915,N_21718,N_21698);
xnor U21916 (N_21916,N_21674,N_21643);
and U21917 (N_21917,N_21640,N_21690);
and U21918 (N_21918,N_21640,N_21746);
and U21919 (N_21919,N_21649,N_21718);
nand U21920 (N_21920,N_21772,N_21662);
and U21921 (N_21921,N_21783,N_21653);
nand U21922 (N_21922,N_21771,N_21709);
or U21923 (N_21923,N_21686,N_21768);
nor U21924 (N_21924,N_21688,N_21740);
nand U21925 (N_21925,N_21635,N_21608);
xnor U21926 (N_21926,N_21788,N_21790);
or U21927 (N_21927,N_21753,N_21745);
xnor U21928 (N_21928,N_21776,N_21613);
nand U21929 (N_21929,N_21774,N_21787);
xor U21930 (N_21930,N_21637,N_21699);
xor U21931 (N_21931,N_21728,N_21692);
or U21932 (N_21932,N_21785,N_21659);
xnor U21933 (N_21933,N_21701,N_21734);
nor U21934 (N_21934,N_21744,N_21664);
nor U21935 (N_21935,N_21600,N_21764);
nor U21936 (N_21936,N_21676,N_21708);
or U21937 (N_21937,N_21676,N_21697);
nand U21938 (N_21938,N_21664,N_21792);
xnor U21939 (N_21939,N_21769,N_21726);
and U21940 (N_21940,N_21710,N_21797);
and U21941 (N_21941,N_21640,N_21631);
and U21942 (N_21942,N_21639,N_21614);
xnor U21943 (N_21943,N_21676,N_21669);
nor U21944 (N_21944,N_21760,N_21657);
and U21945 (N_21945,N_21748,N_21792);
or U21946 (N_21946,N_21665,N_21795);
or U21947 (N_21947,N_21756,N_21705);
xnor U21948 (N_21948,N_21669,N_21635);
xor U21949 (N_21949,N_21775,N_21687);
and U21950 (N_21950,N_21741,N_21637);
or U21951 (N_21951,N_21656,N_21670);
nor U21952 (N_21952,N_21708,N_21620);
and U21953 (N_21953,N_21727,N_21749);
nor U21954 (N_21954,N_21630,N_21658);
nor U21955 (N_21955,N_21763,N_21709);
and U21956 (N_21956,N_21619,N_21616);
nor U21957 (N_21957,N_21738,N_21745);
xor U21958 (N_21958,N_21702,N_21725);
and U21959 (N_21959,N_21656,N_21798);
nor U21960 (N_21960,N_21740,N_21761);
nand U21961 (N_21961,N_21795,N_21724);
xnor U21962 (N_21962,N_21773,N_21721);
or U21963 (N_21963,N_21663,N_21795);
xnor U21964 (N_21964,N_21653,N_21614);
xor U21965 (N_21965,N_21617,N_21748);
nor U21966 (N_21966,N_21718,N_21693);
and U21967 (N_21967,N_21608,N_21788);
nand U21968 (N_21968,N_21656,N_21769);
or U21969 (N_21969,N_21669,N_21653);
nand U21970 (N_21970,N_21791,N_21778);
xnor U21971 (N_21971,N_21699,N_21630);
xor U21972 (N_21972,N_21643,N_21754);
and U21973 (N_21973,N_21786,N_21653);
xor U21974 (N_21974,N_21742,N_21747);
nand U21975 (N_21975,N_21626,N_21630);
and U21976 (N_21976,N_21676,N_21679);
xor U21977 (N_21977,N_21603,N_21763);
nand U21978 (N_21978,N_21687,N_21674);
or U21979 (N_21979,N_21652,N_21611);
xnor U21980 (N_21980,N_21793,N_21719);
nor U21981 (N_21981,N_21755,N_21672);
xnor U21982 (N_21982,N_21761,N_21714);
xnor U21983 (N_21983,N_21727,N_21656);
nor U21984 (N_21984,N_21762,N_21660);
xnor U21985 (N_21985,N_21762,N_21680);
or U21986 (N_21986,N_21657,N_21656);
nand U21987 (N_21987,N_21631,N_21653);
xor U21988 (N_21988,N_21614,N_21624);
and U21989 (N_21989,N_21672,N_21647);
or U21990 (N_21990,N_21796,N_21730);
nand U21991 (N_21991,N_21637,N_21724);
xnor U21992 (N_21992,N_21629,N_21615);
and U21993 (N_21993,N_21691,N_21775);
nand U21994 (N_21994,N_21756,N_21710);
nand U21995 (N_21995,N_21797,N_21684);
xor U21996 (N_21996,N_21615,N_21676);
or U21997 (N_21997,N_21623,N_21665);
and U21998 (N_21998,N_21661,N_21703);
nor U21999 (N_21999,N_21629,N_21744);
xnor U22000 (N_22000,N_21863,N_21934);
nand U22001 (N_22001,N_21947,N_21936);
or U22002 (N_22002,N_21959,N_21957);
and U22003 (N_22003,N_21826,N_21940);
nand U22004 (N_22004,N_21835,N_21926);
and U22005 (N_22005,N_21800,N_21931);
xnor U22006 (N_22006,N_21991,N_21939);
nor U22007 (N_22007,N_21900,N_21841);
nor U22008 (N_22008,N_21852,N_21971);
xor U22009 (N_22009,N_21869,N_21961);
or U22010 (N_22010,N_21986,N_21903);
or U22011 (N_22011,N_21945,N_21833);
xor U22012 (N_22012,N_21875,N_21840);
nor U22013 (N_22013,N_21870,N_21972);
nor U22014 (N_22014,N_21982,N_21809);
or U22015 (N_22015,N_21878,N_21912);
nand U22016 (N_22016,N_21853,N_21948);
and U22017 (N_22017,N_21861,N_21846);
or U22018 (N_22018,N_21886,N_21816);
nand U22019 (N_22019,N_21932,N_21985);
nor U22020 (N_22020,N_21915,N_21801);
nand U22021 (N_22021,N_21894,N_21808);
nor U22022 (N_22022,N_21996,N_21973);
or U22023 (N_22023,N_21879,N_21922);
or U22024 (N_22024,N_21876,N_21997);
or U22025 (N_22025,N_21845,N_21938);
nand U22026 (N_22026,N_21976,N_21956);
nor U22027 (N_22027,N_21871,N_21943);
and U22028 (N_22028,N_21824,N_21812);
nand U22029 (N_22029,N_21814,N_21930);
and U22030 (N_22030,N_21950,N_21838);
nor U22031 (N_22031,N_21919,N_21828);
or U22032 (N_22032,N_21974,N_21983);
and U22033 (N_22033,N_21963,N_21803);
nor U22034 (N_22034,N_21859,N_21905);
and U22035 (N_22035,N_21810,N_21860);
xor U22036 (N_22036,N_21916,N_21832);
or U22037 (N_22037,N_21891,N_21952);
or U22038 (N_22038,N_21975,N_21818);
nor U22039 (N_22039,N_21901,N_21981);
nor U22040 (N_22040,N_21949,N_21898);
or U22041 (N_22041,N_21904,N_21881);
and U22042 (N_22042,N_21849,N_21872);
xnor U22043 (N_22043,N_21909,N_21842);
nand U22044 (N_22044,N_21937,N_21998);
and U22045 (N_22045,N_21914,N_21817);
nand U22046 (N_22046,N_21933,N_21837);
nor U22047 (N_22047,N_21865,N_21893);
and U22048 (N_22048,N_21850,N_21887);
xnor U22049 (N_22049,N_21944,N_21807);
xor U22050 (N_22050,N_21908,N_21966);
and U22051 (N_22051,N_21854,N_21899);
nand U22052 (N_22052,N_21951,N_21862);
or U22053 (N_22053,N_21987,N_21970);
nand U22054 (N_22054,N_21896,N_21913);
xnor U22055 (N_22055,N_21942,N_21918);
nand U22056 (N_22056,N_21839,N_21968);
nor U22057 (N_22057,N_21873,N_21990);
xnor U22058 (N_22058,N_21941,N_21874);
xnor U22059 (N_22059,N_21897,N_21925);
and U22060 (N_22060,N_21980,N_21880);
xnor U22061 (N_22061,N_21829,N_21962);
nand U22062 (N_22062,N_21965,N_21844);
or U22063 (N_22063,N_21855,N_21902);
xnor U22064 (N_22064,N_21946,N_21906);
or U22065 (N_22065,N_21834,N_21917);
xor U22066 (N_22066,N_21954,N_21984);
and U22067 (N_22067,N_21993,N_21836);
nand U22068 (N_22068,N_21977,N_21989);
and U22069 (N_22069,N_21802,N_21994);
nand U22070 (N_22070,N_21907,N_21847);
and U22071 (N_22071,N_21864,N_21921);
nand U22072 (N_22072,N_21848,N_21992);
or U22073 (N_22073,N_21960,N_21929);
nand U22074 (N_22074,N_21964,N_21806);
or U22075 (N_22075,N_21811,N_21953);
xor U22076 (N_22076,N_21822,N_21856);
nand U22077 (N_22077,N_21884,N_21851);
nor U22078 (N_22078,N_21923,N_21967);
and U22079 (N_22079,N_21978,N_21920);
xor U22080 (N_22080,N_21999,N_21969);
and U22081 (N_22081,N_21831,N_21877);
or U22082 (N_22082,N_21815,N_21928);
nor U22083 (N_22083,N_21890,N_21958);
or U22084 (N_22084,N_21866,N_21882);
nor U22085 (N_22085,N_21823,N_21885);
xnor U22086 (N_22086,N_21827,N_21883);
nand U22087 (N_22087,N_21868,N_21927);
xor U22088 (N_22088,N_21867,N_21910);
xnor U22089 (N_22089,N_21830,N_21857);
xnor U22090 (N_22090,N_21820,N_21843);
nand U22091 (N_22091,N_21924,N_21955);
xnor U22092 (N_22092,N_21819,N_21813);
or U22093 (N_22093,N_21805,N_21995);
or U22094 (N_22094,N_21825,N_21858);
or U22095 (N_22095,N_21888,N_21988);
nor U22096 (N_22096,N_21935,N_21895);
nor U22097 (N_22097,N_21911,N_21892);
xor U22098 (N_22098,N_21821,N_21979);
or U22099 (N_22099,N_21804,N_21889);
xnor U22100 (N_22100,N_21989,N_21899);
and U22101 (N_22101,N_21927,N_21892);
nand U22102 (N_22102,N_21950,N_21859);
xnor U22103 (N_22103,N_21931,N_21977);
nor U22104 (N_22104,N_21930,N_21999);
nand U22105 (N_22105,N_21959,N_21820);
or U22106 (N_22106,N_21969,N_21858);
nor U22107 (N_22107,N_21992,N_21988);
and U22108 (N_22108,N_21802,N_21936);
nor U22109 (N_22109,N_21836,N_21930);
xnor U22110 (N_22110,N_21830,N_21930);
and U22111 (N_22111,N_21878,N_21948);
nand U22112 (N_22112,N_21857,N_21942);
and U22113 (N_22113,N_21891,N_21892);
nor U22114 (N_22114,N_21857,N_21863);
xnor U22115 (N_22115,N_21878,N_21970);
and U22116 (N_22116,N_21874,N_21802);
nand U22117 (N_22117,N_21837,N_21819);
or U22118 (N_22118,N_21894,N_21868);
or U22119 (N_22119,N_21923,N_21947);
or U22120 (N_22120,N_21833,N_21954);
nor U22121 (N_22121,N_21804,N_21912);
xor U22122 (N_22122,N_21832,N_21858);
or U22123 (N_22123,N_21866,N_21943);
nor U22124 (N_22124,N_21989,N_21877);
xor U22125 (N_22125,N_21946,N_21990);
nand U22126 (N_22126,N_21829,N_21822);
or U22127 (N_22127,N_21946,N_21862);
nand U22128 (N_22128,N_21968,N_21900);
or U22129 (N_22129,N_21948,N_21922);
or U22130 (N_22130,N_21838,N_21913);
and U22131 (N_22131,N_21972,N_21913);
nand U22132 (N_22132,N_21936,N_21836);
nand U22133 (N_22133,N_21878,N_21991);
and U22134 (N_22134,N_21954,N_21951);
xnor U22135 (N_22135,N_21991,N_21846);
or U22136 (N_22136,N_21910,N_21880);
nand U22137 (N_22137,N_21840,N_21893);
xor U22138 (N_22138,N_21999,N_21833);
nor U22139 (N_22139,N_21956,N_21966);
or U22140 (N_22140,N_21932,N_21908);
xor U22141 (N_22141,N_21841,N_21968);
nand U22142 (N_22142,N_21953,N_21865);
nand U22143 (N_22143,N_21876,N_21949);
or U22144 (N_22144,N_21890,N_21949);
nor U22145 (N_22145,N_21981,N_21860);
nand U22146 (N_22146,N_21959,N_21981);
nor U22147 (N_22147,N_21984,N_21885);
nor U22148 (N_22148,N_21976,N_21910);
xor U22149 (N_22149,N_21901,N_21870);
and U22150 (N_22150,N_21800,N_21805);
xor U22151 (N_22151,N_21945,N_21999);
nor U22152 (N_22152,N_21982,N_21895);
or U22153 (N_22153,N_21989,N_21934);
nor U22154 (N_22154,N_21885,N_21900);
nor U22155 (N_22155,N_21809,N_21902);
or U22156 (N_22156,N_21834,N_21810);
or U22157 (N_22157,N_21807,N_21815);
xnor U22158 (N_22158,N_21959,N_21943);
and U22159 (N_22159,N_21877,N_21984);
nor U22160 (N_22160,N_21989,N_21974);
and U22161 (N_22161,N_21949,N_21922);
nor U22162 (N_22162,N_21832,N_21962);
and U22163 (N_22163,N_21859,N_21964);
and U22164 (N_22164,N_21881,N_21887);
nor U22165 (N_22165,N_21893,N_21926);
nor U22166 (N_22166,N_21922,N_21904);
nor U22167 (N_22167,N_21898,N_21853);
or U22168 (N_22168,N_21901,N_21919);
nor U22169 (N_22169,N_21811,N_21822);
xnor U22170 (N_22170,N_21991,N_21852);
or U22171 (N_22171,N_21940,N_21837);
nor U22172 (N_22172,N_21904,N_21905);
nand U22173 (N_22173,N_21918,N_21810);
and U22174 (N_22174,N_21811,N_21907);
nand U22175 (N_22175,N_21914,N_21847);
nand U22176 (N_22176,N_21971,N_21858);
and U22177 (N_22177,N_21988,N_21976);
xor U22178 (N_22178,N_21820,N_21905);
xor U22179 (N_22179,N_21873,N_21927);
and U22180 (N_22180,N_21926,N_21889);
nand U22181 (N_22181,N_21880,N_21860);
or U22182 (N_22182,N_21996,N_21915);
xor U22183 (N_22183,N_21907,N_21943);
nand U22184 (N_22184,N_21875,N_21809);
and U22185 (N_22185,N_21883,N_21847);
or U22186 (N_22186,N_21874,N_21861);
xnor U22187 (N_22187,N_21977,N_21998);
or U22188 (N_22188,N_21955,N_21820);
xor U22189 (N_22189,N_21978,N_21869);
nor U22190 (N_22190,N_21963,N_21954);
nand U22191 (N_22191,N_21944,N_21863);
or U22192 (N_22192,N_21987,N_21976);
xor U22193 (N_22193,N_21886,N_21994);
xnor U22194 (N_22194,N_21881,N_21849);
or U22195 (N_22195,N_21990,N_21859);
or U22196 (N_22196,N_21919,N_21870);
and U22197 (N_22197,N_21969,N_21914);
xnor U22198 (N_22198,N_21995,N_21983);
nand U22199 (N_22199,N_21899,N_21910);
or U22200 (N_22200,N_22029,N_22160);
nand U22201 (N_22201,N_22133,N_22169);
and U22202 (N_22202,N_22127,N_22054);
nor U22203 (N_22203,N_22101,N_22149);
and U22204 (N_22204,N_22091,N_22147);
and U22205 (N_22205,N_22037,N_22035);
nand U22206 (N_22206,N_22064,N_22023);
nand U22207 (N_22207,N_22123,N_22115);
or U22208 (N_22208,N_22012,N_22103);
and U22209 (N_22209,N_22145,N_22051);
nor U22210 (N_22210,N_22005,N_22027);
nand U22211 (N_22211,N_22017,N_22063);
xor U22212 (N_22212,N_22087,N_22191);
nand U22213 (N_22213,N_22040,N_22121);
and U22214 (N_22214,N_22096,N_22173);
nand U22215 (N_22215,N_22004,N_22020);
or U22216 (N_22216,N_22010,N_22107);
nand U22217 (N_22217,N_22168,N_22136);
xnor U22218 (N_22218,N_22084,N_22082);
xnor U22219 (N_22219,N_22003,N_22086);
or U22220 (N_22220,N_22157,N_22179);
xor U22221 (N_22221,N_22083,N_22182);
nand U22222 (N_22222,N_22112,N_22022);
or U22223 (N_22223,N_22034,N_22011);
xor U22224 (N_22224,N_22069,N_22060);
nand U22225 (N_22225,N_22198,N_22164);
and U22226 (N_22226,N_22106,N_22065);
or U22227 (N_22227,N_22178,N_22071);
and U22228 (N_22228,N_22124,N_22076);
nand U22229 (N_22229,N_22199,N_22097);
xor U22230 (N_22230,N_22153,N_22174);
or U22231 (N_22231,N_22151,N_22187);
xnor U22232 (N_22232,N_22013,N_22036);
or U22233 (N_22233,N_22067,N_22156);
xnor U22234 (N_22234,N_22059,N_22080);
or U22235 (N_22235,N_22105,N_22166);
xor U22236 (N_22236,N_22062,N_22146);
nand U22237 (N_22237,N_22049,N_22077);
or U22238 (N_22238,N_22090,N_22102);
xor U22239 (N_22239,N_22032,N_22038);
and U22240 (N_22240,N_22066,N_22162);
or U22241 (N_22241,N_22093,N_22184);
xor U22242 (N_22242,N_22000,N_22095);
or U22243 (N_22243,N_22197,N_22129);
or U22244 (N_22244,N_22039,N_22055);
nand U22245 (N_22245,N_22117,N_22158);
and U22246 (N_22246,N_22172,N_22144);
or U22247 (N_22247,N_22094,N_22092);
nand U22248 (N_22248,N_22061,N_22050);
xor U22249 (N_22249,N_22175,N_22108);
or U22250 (N_22250,N_22152,N_22183);
xor U22251 (N_22251,N_22002,N_22193);
nor U22252 (N_22252,N_22070,N_22137);
and U22253 (N_22253,N_22044,N_22014);
nor U22254 (N_22254,N_22181,N_22155);
and U22255 (N_22255,N_22078,N_22185);
xor U22256 (N_22256,N_22116,N_22056);
nor U22257 (N_22257,N_22189,N_22159);
nand U22258 (N_22258,N_22100,N_22072);
or U22259 (N_22259,N_22041,N_22104);
xor U22260 (N_22260,N_22141,N_22001);
nor U22261 (N_22261,N_22131,N_22163);
nor U22262 (N_22262,N_22120,N_22114);
and U22263 (N_22263,N_22068,N_22109);
nor U22264 (N_22264,N_22007,N_22188);
and U22265 (N_22265,N_22006,N_22122);
nor U22266 (N_22266,N_22088,N_22053);
xnor U22267 (N_22267,N_22042,N_22110);
nand U22268 (N_22268,N_22030,N_22143);
or U22269 (N_22269,N_22138,N_22089);
and U22270 (N_22270,N_22154,N_22161);
nand U22271 (N_22271,N_22167,N_22028);
nand U22272 (N_22272,N_22186,N_22177);
or U22273 (N_22273,N_22008,N_22045);
nor U22274 (N_22274,N_22194,N_22118);
nand U22275 (N_22275,N_22074,N_22170);
and U22276 (N_22276,N_22135,N_22180);
nor U22277 (N_22277,N_22058,N_22099);
and U22278 (N_22278,N_22125,N_22130);
xor U22279 (N_22279,N_22081,N_22165);
and U22280 (N_22280,N_22190,N_22113);
nor U22281 (N_22281,N_22196,N_22192);
xnor U22282 (N_22282,N_22057,N_22009);
xor U22283 (N_22283,N_22024,N_22018);
nand U22284 (N_22284,N_22128,N_22073);
and U22285 (N_22285,N_22026,N_22098);
nand U22286 (N_22286,N_22148,N_22176);
xnor U22287 (N_22287,N_22142,N_22021);
nand U22288 (N_22288,N_22048,N_22171);
or U22289 (N_22289,N_22139,N_22079);
nand U22290 (N_22290,N_22016,N_22134);
or U22291 (N_22291,N_22195,N_22015);
or U22292 (N_22292,N_22019,N_22150);
or U22293 (N_22293,N_22033,N_22043);
xor U22294 (N_22294,N_22047,N_22119);
nand U22295 (N_22295,N_22025,N_22126);
nand U22296 (N_22296,N_22140,N_22031);
xnor U22297 (N_22297,N_22085,N_22111);
and U22298 (N_22298,N_22132,N_22052);
nor U22299 (N_22299,N_22046,N_22075);
xor U22300 (N_22300,N_22011,N_22084);
xnor U22301 (N_22301,N_22102,N_22033);
nor U22302 (N_22302,N_22158,N_22134);
nor U22303 (N_22303,N_22025,N_22124);
or U22304 (N_22304,N_22144,N_22079);
xnor U22305 (N_22305,N_22147,N_22025);
xnor U22306 (N_22306,N_22008,N_22096);
nand U22307 (N_22307,N_22134,N_22131);
xor U22308 (N_22308,N_22095,N_22187);
and U22309 (N_22309,N_22179,N_22001);
xnor U22310 (N_22310,N_22188,N_22105);
xor U22311 (N_22311,N_22053,N_22137);
nand U22312 (N_22312,N_22043,N_22038);
nand U22313 (N_22313,N_22151,N_22100);
and U22314 (N_22314,N_22086,N_22160);
or U22315 (N_22315,N_22002,N_22016);
xor U22316 (N_22316,N_22052,N_22162);
nor U22317 (N_22317,N_22175,N_22141);
nor U22318 (N_22318,N_22148,N_22116);
xnor U22319 (N_22319,N_22159,N_22130);
xnor U22320 (N_22320,N_22053,N_22112);
and U22321 (N_22321,N_22078,N_22049);
nand U22322 (N_22322,N_22107,N_22049);
or U22323 (N_22323,N_22025,N_22160);
and U22324 (N_22324,N_22025,N_22063);
nand U22325 (N_22325,N_22059,N_22149);
nor U22326 (N_22326,N_22137,N_22143);
xor U22327 (N_22327,N_22012,N_22114);
and U22328 (N_22328,N_22074,N_22131);
nor U22329 (N_22329,N_22068,N_22134);
or U22330 (N_22330,N_22067,N_22008);
nor U22331 (N_22331,N_22129,N_22101);
nand U22332 (N_22332,N_22117,N_22114);
nand U22333 (N_22333,N_22093,N_22078);
or U22334 (N_22334,N_22119,N_22131);
xor U22335 (N_22335,N_22174,N_22088);
nand U22336 (N_22336,N_22025,N_22026);
and U22337 (N_22337,N_22076,N_22025);
xnor U22338 (N_22338,N_22070,N_22039);
and U22339 (N_22339,N_22180,N_22101);
xnor U22340 (N_22340,N_22113,N_22133);
or U22341 (N_22341,N_22117,N_22054);
nand U22342 (N_22342,N_22171,N_22199);
or U22343 (N_22343,N_22033,N_22142);
and U22344 (N_22344,N_22025,N_22036);
xnor U22345 (N_22345,N_22104,N_22161);
nor U22346 (N_22346,N_22021,N_22064);
or U22347 (N_22347,N_22123,N_22032);
nor U22348 (N_22348,N_22059,N_22104);
nor U22349 (N_22349,N_22093,N_22109);
and U22350 (N_22350,N_22171,N_22023);
nand U22351 (N_22351,N_22038,N_22137);
xor U22352 (N_22352,N_22133,N_22042);
nand U22353 (N_22353,N_22086,N_22158);
nand U22354 (N_22354,N_22184,N_22119);
nor U22355 (N_22355,N_22169,N_22194);
nand U22356 (N_22356,N_22197,N_22150);
nand U22357 (N_22357,N_22044,N_22120);
and U22358 (N_22358,N_22196,N_22049);
xor U22359 (N_22359,N_22128,N_22044);
nor U22360 (N_22360,N_22199,N_22044);
nor U22361 (N_22361,N_22179,N_22035);
and U22362 (N_22362,N_22161,N_22052);
or U22363 (N_22363,N_22003,N_22069);
and U22364 (N_22364,N_22015,N_22080);
nand U22365 (N_22365,N_22148,N_22047);
and U22366 (N_22366,N_22063,N_22189);
nor U22367 (N_22367,N_22116,N_22068);
and U22368 (N_22368,N_22111,N_22039);
or U22369 (N_22369,N_22125,N_22002);
or U22370 (N_22370,N_22046,N_22165);
xnor U22371 (N_22371,N_22081,N_22105);
nor U22372 (N_22372,N_22010,N_22116);
nand U22373 (N_22373,N_22154,N_22001);
nor U22374 (N_22374,N_22131,N_22165);
and U22375 (N_22375,N_22188,N_22133);
xnor U22376 (N_22376,N_22071,N_22037);
or U22377 (N_22377,N_22181,N_22032);
xor U22378 (N_22378,N_22080,N_22171);
nor U22379 (N_22379,N_22144,N_22083);
and U22380 (N_22380,N_22188,N_22189);
xor U22381 (N_22381,N_22037,N_22001);
and U22382 (N_22382,N_22004,N_22037);
xnor U22383 (N_22383,N_22159,N_22060);
xor U22384 (N_22384,N_22122,N_22061);
nor U22385 (N_22385,N_22162,N_22160);
or U22386 (N_22386,N_22095,N_22061);
xor U22387 (N_22387,N_22038,N_22102);
nor U22388 (N_22388,N_22114,N_22118);
and U22389 (N_22389,N_22113,N_22063);
nor U22390 (N_22390,N_22008,N_22097);
and U22391 (N_22391,N_22074,N_22049);
or U22392 (N_22392,N_22012,N_22081);
or U22393 (N_22393,N_22004,N_22115);
and U22394 (N_22394,N_22044,N_22137);
nor U22395 (N_22395,N_22033,N_22126);
nor U22396 (N_22396,N_22078,N_22118);
nor U22397 (N_22397,N_22143,N_22060);
or U22398 (N_22398,N_22152,N_22016);
nor U22399 (N_22399,N_22169,N_22053);
and U22400 (N_22400,N_22229,N_22287);
and U22401 (N_22401,N_22213,N_22360);
and U22402 (N_22402,N_22324,N_22286);
nand U22403 (N_22403,N_22228,N_22334);
xor U22404 (N_22404,N_22302,N_22277);
and U22405 (N_22405,N_22327,N_22364);
xor U22406 (N_22406,N_22268,N_22217);
and U22407 (N_22407,N_22250,N_22280);
xor U22408 (N_22408,N_22244,N_22206);
or U22409 (N_22409,N_22380,N_22224);
or U22410 (N_22410,N_22245,N_22220);
nand U22411 (N_22411,N_22341,N_22314);
xnor U22412 (N_22412,N_22271,N_22330);
or U22413 (N_22413,N_22331,N_22305);
nand U22414 (N_22414,N_22316,N_22375);
and U22415 (N_22415,N_22320,N_22219);
nor U22416 (N_22416,N_22209,N_22263);
and U22417 (N_22417,N_22221,N_22311);
nand U22418 (N_22418,N_22378,N_22211);
xor U22419 (N_22419,N_22256,N_22355);
nand U22420 (N_22420,N_22387,N_22201);
xor U22421 (N_22421,N_22281,N_22299);
nor U22422 (N_22422,N_22267,N_22264);
and U22423 (N_22423,N_22390,N_22363);
or U22424 (N_22424,N_22313,N_22322);
and U22425 (N_22425,N_22352,N_22356);
or U22426 (N_22426,N_22207,N_22232);
nand U22427 (N_22427,N_22237,N_22365);
and U22428 (N_22428,N_22369,N_22321);
nand U22429 (N_22429,N_22293,N_22292);
nor U22430 (N_22430,N_22307,N_22389);
nor U22431 (N_22431,N_22298,N_22301);
nand U22432 (N_22432,N_22214,N_22241);
and U22433 (N_22433,N_22384,N_22223);
nor U22434 (N_22434,N_22349,N_22273);
and U22435 (N_22435,N_22383,N_22372);
or U22436 (N_22436,N_22336,N_22391);
and U22437 (N_22437,N_22367,N_22253);
xnor U22438 (N_22438,N_22265,N_22353);
nand U22439 (N_22439,N_22239,N_22278);
nand U22440 (N_22440,N_22381,N_22394);
and U22441 (N_22441,N_22399,N_22258);
nand U22442 (N_22442,N_22257,N_22251);
nand U22443 (N_22443,N_22344,N_22315);
nand U22444 (N_22444,N_22275,N_22386);
xor U22445 (N_22445,N_22368,N_22233);
nand U22446 (N_22446,N_22359,N_22385);
xnor U22447 (N_22447,N_22238,N_22342);
nor U22448 (N_22448,N_22395,N_22222);
or U22449 (N_22449,N_22347,N_22376);
nor U22450 (N_22450,N_22205,N_22397);
or U22451 (N_22451,N_22304,N_22242);
nand U22452 (N_22452,N_22358,N_22300);
or U22453 (N_22453,N_22335,N_22296);
or U22454 (N_22454,N_22323,N_22261);
xnor U22455 (N_22455,N_22284,N_22246);
nand U22456 (N_22456,N_22306,N_22260);
xnor U22457 (N_22457,N_22318,N_22294);
nor U22458 (N_22458,N_22252,N_22283);
nor U22459 (N_22459,N_22329,N_22231);
nor U22460 (N_22460,N_22297,N_22377);
or U22461 (N_22461,N_22343,N_22203);
nor U22462 (N_22462,N_22393,N_22398);
xor U22463 (N_22463,N_22351,N_22370);
or U22464 (N_22464,N_22202,N_22262);
and U22465 (N_22465,N_22215,N_22357);
xor U22466 (N_22466,N_22210,N_22362);
or U22467 (N_22467,N_22354,N_22333);
and U22468 (N_22468,N_22276,N_22332);
and U22469 (N_22469,N_22325,N_22279);
nor U22470 (N_22470,N_22312,N_22388);
or U22471 (N_22471,N_22240,N_22326);
nor U22472 (N_22472,N_22303,N_22212);
xor U22473 (N_22473,N_22339,N_22289);
or U22474 (N_22474,N_22282,N_22235);
and U22475 (N_22475,N_22288,N_22337);
nand U22476 (N_22476,N_22200,N_22226);
xnor U22477 (N_22477,N_22225,N_22361);
nor U22478 (N_22478,N_22348,N_22295);
nand U22479 (N_22479,N_22204,N_22227);
nand U22480 (N_22480,N_22243,N_22270);
nand U22481 (N_22481,N_22346,N_22308);
nand U22482 (N_22482,N_22319,N_22340);
nand U22483 (N_22483,N_22230,N_22234);
nor U22484 (N_22484,N_22216,N_22247);
nand U22485 (N_22485,N_22350,N_22328);
nor U22486 (N_22486,N_22373,N_22254);
xnor U22487 (N_22487,N_22249,N_22366);
nor U22488 (N_22488,N_22274,N_22396);
or U22489 (N_22489,N_22255,N_22248);
nor U22490 (N_22490,N_22266,N_22290);
nand U22491 (N_22491,N_22285,N_22310);
nand U22492 (N_22492,N_22218,N_22392);
nor U22493 (N_22493,N_22208,N_22345);
nand U22494 (N_22494,N_22236,N_22259);
nor U22495 (N_22495,N_22317,N_22379);
nor U22496 (N_22496,N_22272,N_22371);
and U22497 (N_22497,N_22382,N_22309);
xor U22498 (N_22498,N_22269,N_22291);
or U22499 (N_22499,N_22338,N_22374);
nor U22500 (N_22500,N_22354,N_22201);
and U22501 (N_22501,N_22230,N_22371);
xor U22502 (N_22502,N_22220,N_22232);
or U22503 (N_22503,N_22260,N_22221);
nor U22504 (N_22504,N_22237,N_22364);
and U22505 (N_22505,N_22233,N_22268);
nor U22506 (N_22506,N_22246,N_22286);
nor U22507 (N_22507,N_22283,N_22376);
nand U22508 (N_22508,N_22390,N_22206);
or U22509 (N_22509,N_22281,N_22370);
nor U22510 (N_22510,N_22271,N_22251);
xnor U22511 (N_22511,N_22222,N_22283);
or U22512 (N_22512,N_22265,N_22235);
xor U22513 (N_22513,N_22349,N_22399);
and U22514 (N_22514,N_22237,N_22327);
nor U22515 (N_22515,N_22379,N_22329);
nand U22516 (N_22516,N_22301,N_22312);
or U22517 (N_22517,N_22303,N_22396);
nor U22518 (N_22518,N_22322,N_22275);
or U22519 (N_22519,N_22219,N_22290);
or U22520 (N_22520,N_22330,N_22300);
and U22521 (N_22521,N_22203,N_22248);
nand U22522 (N_22522,N_22302,N_22246);
nor U22523 (N_22523,N_22335,N_22371);
nor U22524 (N_22524,N_22287,N_22285);
nor U22525 (N_22525,N_22335,N_22336);
xor U22526 (N_22526,N_22383,N_22398);
or U22527 (N_22527,N_22268,N_22257);
nand U22528 (N_22528,N_22382,N_22339);
nand U22529 (N_22529,N_22374,N_22208);
and U22530 (N_22530,N_22336,N_22353);
or U22531 (N_22531,N_22303,N_22317);
or U22532 (N_22532,N_22335,N_22212);
and U22533 (N_22533,N_22315,N_22393);
xor U22534 (N_22534,N_22222,N_22248);
xor U22535 (N_22535,N_22363,N_22297);
nor U22536 (N_22536,N_22287,N_22328);
nor U22537 (N_22537,N_22212,N_22288);
nand U22538 (N_22538,N_22248,N_22219);
xnor U22539 (N_22539,N_22326,N_22320);
nand U22540 (N_22540,N_22237,N_22350);
and U22541 (N_22541,N_22276,N_22262);
and U22542 (N_22542,N_22214,N_22354);
nand U22543 (N_22543,N_22313,N_22344);
nor U22544 (N_22544,N_22211,N_22203);
nand U22545 (N_22545,N_22298,N_22293);
or U22546 (N_22546,N_22339,N_22261);
and U22547 (N_22547,N_22272,N_22291);
or U22548 (N_22548,N_22331,N_22279);
xnor U22549 (N_22549,N_22396,N_22350);
nand U22550 (N_22550,N_22200,N_22381);
or U22551 (N_22551,N_22364,N_22354);
and U22552 (N_22552,N_22205,N_22249);
or U22553 (N_22553,N_22248,N_22258);
xnor U22554 (N_22554,N_22278,N_22365);
or U22555 (N_22555,N_22212,N_22269);
nor U22556 (N_22556,N_22366,N_22299);
nor U22557 (N_22557,N_22352,N_22216);
xnor U22558 (N_22558,N_22293,N_22250);
nor U22559 (N_22559,N_22364,N_22347);
xor U22560 (N_22560,N_22249,N_22363);
and U22561 (N_22561,N_22241,N_22233);
nor U22562 (N_22562,N_22235,N_22262);
nor U22563 (N_22563,N_22221,N_22203);
xor U22564 (N_22564,N_22377,N_22396);
and U22565 (N_22565,N_22280,N_22228);
xor U22566 (N_22566,N_22369,N_22203);
nand U22567 (N_22567,N_22328,N_22358);
nor U22568 (N_22568,N_22374,N_22260);
nor U22569 (N_22569,N_22381,N_22254);
nand U22570 (N_22570,N_22222,N_22239);
and U22571 (N_22571,N_22293,N_22393);
or U22572 (N_22572,N_22385,N_22395);
and U22573 (N_22573,N_22230,N_22297);
or U22574 (N_22574,N_22249,N_22287);
nor U22575 (N_22575,N_22273,N_22202);
xor U22576 (N_22576,N_22252,N_22361);
or U22577 (N_22577,N_22242,N_22283);
nand U22578 (N_22578,N_22222,N_22217);
xnor U22579 (N_22579,N_22242,N_22360);
nor U22580 (N_22580,N_22292,N_22391);
xor U22581 (N_22581,N_22230,N_22311);
nor U22582 (N_22582,N_22391,N_22317);
nand U22583 (N_22583,N_22237,N_22211);
and U22584 (N_22584,N_22399,N_22240);
and U22585 (N_22585,N_22206,N_22220);
nor U22586 (N_22586,N_22235,N_22331);
and U22587 (N_22587,N_22290,N_22236);
nor U22588 (N_22588,N_22243,N_22260);
or U22589 (N_22589,N_22302,N_22362);
or U22590 (N_22590,N_22328,N_22266);
and U22591 (N_22591,N_22342,N_22286);
or U22592 (N_22592,N_22261,N_22337);
nand U22593 (N_22593,N_22293,N_22353);
nor U22594 (N_22594,N_22321,N_22303);
and U22595 (N_22595,N_22273,N_22346);
and U22596 (N_22596,N_22397,N_22299);
nand U22597 (N_22597,N_22229,N_22383);
nor U22598 (N_22598,N_22249,N_22231);
nor U22599 (N_22599,N_22221,N_22303);
and U22600 (N_22600,N_22574,N_22545);
nand U22601 (N_22601,N_22493,N_22515);
xnor U22602 (N_22602,N_22536,N_22594);
and U22603 (N_22603,N_22461,N_22540);
and U22604 (N_22604,N_22592,N_22570);
nand U22605 (N_22605,N_22478,N_22460);
nor U22606 (N_22606,N_22528,N_22514);
nand U22607 (N_22607,N_22572,N_22524);
or U22608 (N_22608,N_22546,N_22464);
and U22609 (N_22609,N_22486,N_22596);
nand U22610 (N_22610,N_22549,N_22561);
and U22611 (N_22611,N_22521,N_22569);
xor U22612 (N_22612,N_22440,N_22492);
xor U22613 (N_22613,N_22522,N_22428);
and U22614 (N_22614,N_22500,N_22562);
and U22615 (N_22615,N_22523,N_22418);
xnor U22616 (N_22616,N_22404,N_22436);
and U22617 (N_22617,N_22482,N_22576);
nand U22618 (N_22618,N_22502,N_22425);
nor U22619 (N_22619,N_22438,N_22581);
nor U22620 (N_22620,N_22547,N_22580);
nand U22621 (N_22621,N_22408,N_22503);
nor U22622 (N_22622,N_22585,N_22504);
or U22623 (N_22623,N_22535,N_22566);
nor U22624 (N_22624,N_22597,N_22488);
nor U22625 (N_22625,N_22445,N_22573);
or U22626 (N_22626,N_22485,N_22589);
nand U22627 (N_22627,N_22400,N_22577);
nand U22628 (N_22628,N_22409,N_22453);
xor U22629 (N_22629,N_22419,N_22458);
nand U22630 (N_22630,N_22582,N_22477);
xnor U22631 (N_22631,N_22530,N_22431);
nand U22632 (N_22632,N_22527,N_22497);
or U22633 (N_22633,N_22519,N_22417);
nand U22634 (N_22634,N_22402,N_22447);
xnor U22635 (N_22635,N_22529,N_22587);
nor U22636 (N_22636,N_22463,N_22434);
or U22637 (N_22637,N_22469,N_22498);
nor U22638 (N_22638,N_22505,N_22411);
xnor U22639 (N_22639,N_22552,N_22538);
nor U22640 (N_22640,N_22533,N_22490);
nor U22641 (N_22641,N_22583,N_22520);
and U22642 (N_22642,N_22548,N_22508);
xor U22643 (N_22643,N_22451,N_22537);
nor U22644 (N_22644,N_22414,N_22517);
nor U22645 (N_22645,N_22420,N_22446);
xnor U22646 (N_22646,N_22443,N_22454);
nand U22647 (N_22647,N_22432,N_22467);
and U22648 (N_22648,N_22450,N_22471);
nand U22649 (N_22649,N_22466,N_22511);
and U22650 (N_22650,N_22456,N_22416);
nand U22651 (N_22651,N_22513,N_22544);
xor U22652 (N_22652,N_22413,N_22484);
or U22653 (N_22653,N_22584,N_22421);
and U22654 (N_22654,N_22586,N_22422);
nand U22655 (N_22655,N_22483,N_22579);
and U22656 (N_22656,N_22439,N_22495);
xor U22657 (N_22657,N_22541,N_22433);
xnor U22658 (N_22658,N_22560,N_22526);
nand U22659 (N_22659,N_22598,N_22465);
nor U22660 (N_22660,N_22501,N_22506);
and U22661 (N_22661,N_22557,N_22479);
nor U22662 (N_22662,N_22542,N_22468);
or U22663 (N_22663,N_22424,N_22470);
or U22664 (N_22664,N_22578,N_22455);
nor U22665 (N_22665,N_22472,N_22430);
xnor U22666 (N_22666,N_22588,N_22599);
and U22667 (N_22667,N_22567,N_22437);
or U22668 (N_22668,N_22565,N_22449);
nor U22669 (N_22669,N_22555,N_22423);
nand U22670 (N_22670,N_22539,N_22550);
nand U22671 (N_22671,N_22516,N_22457);
nand U22672 (N_22672,N_22494,N_22429);
and U22673 (N_22673,N_22435,N_22412);
and U22674 (N_22674,N_22489,N_22462);
nor U22675 (N_22675,N_22553,N_22452);
nor U22676 (N_22676,N_22407,N_22448);
xnor U22677 (N_22677,N_22481,N_22558);
and U22678 (N_22678,N_22531,N_22534);
or U22679 (N_22679,N_22487,N_22563);
nor U22680 (N_22680,N_22401,N_22590);
and U22681 (N_22681,N_22510,N_22476);
xor U22682 (N_22682,N_22499,N_22442);
or U22683 (N_22683,N_22474,N_22543);
and U22684 (N_22684,N_22525,N_22551);
or U22685 (N_22685,N_22571,N_22403);
xnor U22686 (N_22686,N_22554,N_22473);
or U22687 (N_22687,N_22559,N_22568);
or U22688 (N_22688,N_22444,N_22475);
or U22689 (N_22689,N_22496,N_22575);
xnor U22690 (N_22690,N_22593,N_22512);
and U22691 (N_22691,N_22595,N_22441);
nor U22692 (N_22692,N_22556,N_22459);
nor U22693 (N_22693,N_22509,N_22564);
nor U22694 (N_22694,N_22427,N_22480);
nor U22695 (N_22695,N_22532,N_22406);
nand U22696 (N_22696,N_22415,N_22410);
and U22697 (N_22697,N_22405,N_22491);
or U22698 (N_22698,N_22591,N_22426);
xor U22699 (N_22699,N_22518,N_22507);
xnor U22700 (N_22700,N_22446,N_22439);
xor U22701 (N_22701,N_22499,N_22485);
nand U22702 (N_22702,N_22558,N_22430);
or U22703 (N_22703,N_22524,N_22544);
and U22704 (N_22704,N_22507,N_22558);
nor U22705 (N_22705,N_22557,N_22522);
xnor U22706 (N_22706,N_22595,N_22556);
nand U22707 (N_22707,N_22448,N_22567);
and U22708 (N_22708,N_22456,N_22499);
and U22709 (N_22709,N_22594,N_22579);
nor U22710 (N_22710,N_22530,N_22556);
and U22711 (N_22711,N_22538,N_22530);
xor U22712 (N_22712,N_22450,N_22599);
xnor U22713 (N_22713,N_22451,N_22401);
or U22714 (N_22714,N_22495,N_22525);
or U22715 (N_22715,N_22430,N_22467);
or U22716 (N_22716,N_22585,N_22495);
nor U22717 (N_22717,N_22577,N_22452);
nor U22718 (N_22718,N_22482,N_22502);
xor U22719 (N_22719,N_22509,N_22526);
and U22720 (N_22720,N_22581,N_22575);
nor U22721 (N_22721,N_22502,N_22534);
nor U22722 (N_22722,N_22563,N_22408);
nor U22723 (N_22723,N_22545,N_22405);
or U22724 (N_22724,N_22494,N_22405);
nor U22725 (N_22725,N_22468,N_22573);
xor U22726 (N_22726,N_22498,N_22481);
xor U22727 (N_22727,N_22526,N_22406);
nand U22728 (N_22728,N_22420,N_22585);
or U22729 (N_22729,N_22476,N_22500);
or U22730 (N_22730,N_22462,N_22444);
nand U22731 (N_22731,N_22481,N_22414);
nand U22732 (N_22732,N_22462,N_22473);
nand U22733 (N_22733,N_22589,N_22456);
and U22734 (N_22734,N_22570,N_22512);
and U22735 (N_22735,N_22500,N_22556);
nand U22736 (N_22736,N_22452,N_22582);
and U22737 (N_22737,N_22420,N_22425);
and U22738 (N_22738,N_22499,N_22467);
and U22739 (N_22739,N_22544,N_22469);
nor U22740 (N_22740,N_22569,N_22597);
and U22741 (N_22741,N_22533,N_22459);
xnor U22742 (N_22742,N_22513,N_22552);
or U22743 (N_22743,N_22543,N_22490);
nand U22744 (N_22744,N_22547,N_22597);
and U22745 (N_22745,N_22455,N_22466);
xor U22746 (N_22746,N_22451,N_22566);
nand U22747 (N_22747,N_22490,N_22400);
nand U22748 (N_22748,N_22463,N_22521);
and U22749 (N_22749,N_22412,N_22598);
xnor U22750 (N_22750,N_22597,N_22485);
nand U22751 (N_22751,N_22410,N_22574);
nor U22752 (N_22752,N_22482,N_22462);
or U22753 (N_22753,N_22461,N_22424);
nand U22754 (N_22754,N_22568,N_22414);
and U22755 (N_22755,N_22582,N_22520);
nand U22756 (N_22756,N_22458,N_22429);
xor U22757 (N_22757,N_22420,N_22572);
nor U22758 (N_22758,N_22438,N_22588);
nor U22759 (N_22759,N_22465,N_22536);
or U22760 (N_22760,N_22436,N_22545);
xnor U22761 (N_22761,N_22453,N_22404);
and U22762 (N_22762,N_22557,N_22592);
nor U22763 (N_22763,N_22434,N_22516);
or U22764 (N_22764,N_22443,N_22493);
or U22765 (N_22765,N_22549,N_22580);
and U22766 (N_22766,N_22420,N_22552);
and U22767 (N_22767,N_22496,N_22488);
nand U22768 (N_22768,N_22596,N_22526);
and U22769 (N_22769,N_22413,N_22401);
and U22770 (N_22770,N_22591,N_22534);
nor U22771 (N_22771,N_22560,N_22470);
xor U22772 (N_22772,N_22423,N_22419);
nor U22773 (N_22773,N_22568,N_22567);
or U22774 (N_22774,N_22470,N_22480);
nand U22775 (N_22775,N_22545,N_22424);
nand U22776 (N_22776,N_22585,N_22409);
nor U22777 (N_22777,N_22417,N_22520);
nor U22778 (N_22778,N_22551,N_22410);
and U22779 (N_22779,N_22552,N_22489);
nand U22780 (N_22780,N_22501,N_22491);
xor U22781 (N_22781,N_22599,N_22540);
and U22782 (N_22782,N_22457,N_22475);
nor U22783 (N_22783,N_22440,N_22571);
xnor U22784 (N_22784,N_22530,N_22524);
nand U22785 (N_22785,N_22422,N_22539);
and U22786 (N_22786,N_22552,N_22507);
xor U22787 (N_22787,N_22443,N_22594);
and U22788 (N_22788,N_22599,N_22473);
nor U22789 (N_22789,N_22519,N_22539);
and U22790 (N_22790,N_22556,N_22541);
nor U22791 (N_22791,N_22466,N_22429);
and U22792 (N_22792,N_22411,N_22575);
nor U22793 (N_22793,N_22438,N_22488);
nand U22794 (N_22794,N_22443,N_22468);
and U22795 (N_22795,N_22454,N_22502);
xor U22796 (N_22796,N_22438,N_22460);
and U22797 (N_22797,N_22472,N_22492);
nand U22798 (N_22798,N_22439,N_22403);
or U22799 (N_22799,N_22581,N_22407);
nor U22800 (N_22800,N_22718,N_22701);
or U22801 (N_22801,N_22727,N_22615);
or U22802 (N_22802,N_22662,N_22765);
or U22803 (N_22803,N_22744,N_22725);
nand U22804 (N_22804,N_22714,N_22600);
or U22805 (N_22805,N_22677,N_22777);
nor U22806 (N_22806,N_22657,N_22645);
and U22807 (N_22807,N_22712,N_22736);
nand U22808 (N_22808,N_22604,N_22702);
nor U22809 (N_22809,N_22745,N_22617);
nor U22810 (N_22810,N_22709,N_22748);
or U22811 (N_22811,N_22774,N_22775);
nand U22812 (N_22812,N_22637,N_22618);
xor U22813 (N_22813,N_22755,N_22644);
or U22814 (N_22814,N_22738,N_22666);
nand U22815 (N_22815,N_22758,N_22678);
and U22816 (N_22816,N_22746,N_22768);
nor U22817 (N_22817,N_22631,N_22628);
nor U22818 (N_22818,N_22747,N_22793);
or U22819 (N_22819,N_22616,N_22764);
xnor U22820 (N_22820,N_22750,N_22782);
nor U22821 (N_22821,N_22681,N_22717);
or U22822 (N_22822,N_22694,N_22625);
xnor U22823 (N_22823,N_22708,N_22756);
and U22824 (N_22824,N_22691,N_22606);
or U22825 (N_22825,N_22672,N_22649);
xnor U22826 (N_22826,N_22737,N_22733);
nand U22827 (N_22827,N_22647,N_22608);
nor U22828 (N_22828,N_22661,N_22794);
nand U22829 (N_22829,N_22638,N_22707);
nor U22830 (N_22830,N_22773,N_22713);
and U22831 (N_22831,N_22669,N_22726);
xor U22832 (N_22832,N_22673,N_22633);
nand U22833 (N_22833,N_22721,N_22619);
or U22834 (N_22834,N_22620,N_22705);
nor U22835 (N_22835,N_22656,N_22760);
xnor U22836 (N_22836,N_22622,N_22728);
nand U22837 (N_22837,N_22697,N_22766);
nor U22838 (N_22838,N_22719,N_22663);
and U22839 (N_22839,N_22770,N_22761);
nor U22840 (N_22840,N_22660,N_22641);
and U22841 (N_22841,N_22687,N_22698);
nor U22842 (N_22842,N_22646,N_22602);
and U22843 (N_22843,N_22632,N_22611);
xnor U22844 (N_22844,N_22706,N_22634);
or U22845 (N_22845,N_22688,N_22715);
nand U22846 (N_22846,N_22724,N_22796);
xor U22847 (N_22847,N_22772,N_22786);
nor U22848 (N_22848,N_22704,N_22729);
nor U22849 (N_22849,N_22730,N_22659);
nand U22850 (N_22850,N_22603,N_22742);
and U22851 (N_22851,N_22609,N_22612);
or U22852 (N_22852,N_22689,N_22665);
nor U22853 (N_22853,N_22734,N_22664);
or U22854 (N_22854,N_22754,N_22642);
nor U22855 (N_22855,N_22605,N_22759);
nor U22856 (N_22856,N_22679,N_22739);
and U22857 (N_22857,N_22716,N_22703);
nor U22858 (N_22858,N_22696,N_22654);
nand U22859 (N_22859,N_22627,N_22787);
nor U22860 (N_22860,N_22683,N_22751);
or U22861 (N_22861,N_22720,N_22731);
nor U22862 (N_22862,N_22797,N_22763);
and U22863 (N_22863,N_22798,N_22629);
nor U22864 (N_22864,N_22630,N_22675);
nand U22865 (N_22865,N_22684,N_22643);
nor U22866 (N_22866,N_22732,N_22690);
and U22867 (N_22867,N_22648,N_22785);
or U22868 (N_22868,N_22762,N_22607);
nor U22869 (N_22869,N_22613,N_22740);
and U22870 (N_22870,N_22790,N_22636);
nor U22871 (N_22871,N_22621,N_22655);
xnor U22872 (N_22872,N_22614,N_22780);
nor U22873 (N_22873,N_22735,N_22753);
nor U22874 (N_22874,N_22791,N_22640);
or U22875 (N_22875,N_22653,N_22799);
nor U22876 (N_22876,N_22769,N_22695);
or U22877 (N_22877,N_22781,N_22741);
or U22878 (N_22878,N_22711,N_22778);
or U22879 (N_22879,N_22710,N_22651);
nor U22880 (N_22880,N_22685,N_22693);
and U22881 (N_22881,N_22624,N_22752);
or U22882 (N_22882,N_22635,N_22784);
and U22883 (N_22883,N_22674,N_22757);
or U22884 (N_22884,N_22771,N_22692);
nand U22885 (N_22885,N_22671,N_22667);
xor U22886 (N_22886,N_22783,N_22749);
xnor U22887 (N_22887,N_22792,N_22788);
xnor U22888 (N_22888,N_22779,N_22743);
and U22889 (N_22889,N_22658,N_22686);
or U22890 (N_22890,N_22680,N_22789);
nor U22891 (N_22891,N_22795,N_22601);
or U22892 (N_22892,N_22776,N_22670);
and U22893 (N_22893,N_22650,N_22699);
xnor U22894 (N_22894,N_22626,N_22652);
or U22895 (N_22895,N_22639,N_22700);
nor U22896 (N_22896,N_22722,N_22767);
nor U22897 (N_22897,N_22668,N_22682);
nand U22898 (N_22898,N_22676,N_22623);
nand U22899 (N_22899,N_22723,N_22610);
and U22900 (N_22900,N_22623,N_22718);
xnor U22901 (N_22901,N_22785,N_22767);
xor U22902 (N_22902,N_22689,N_22706);
nor U22903 (N_22903,N_22776,N_22777);
and U22904 (N_22904,N_22604,N_22786);
or U22905 (N_22905,N_22775,N_22677);
xnor U22906 (N_22906,N_22647,N_22734);
and U22907 (N_22907,N_22759,N_22652);
or U22908 (N_22908,N_22793,N_22629);
nand U22909 (N_22909,N_22694,N_22754);
and U22910 (N_22910,N_22793,N_22678);
xor U22911 (N_22911,N_22633,N_22649);
nand U22912 (N_22912,N_22781,N_22662);
xnor U22913 (N_22913,N_22799,N_22645);
nor U22914 (N_22914,N_22625,N_22707);
and U22915 (N_22915,N_22688,N_22696);
xnor U22916 (N_22916,N_22732,N_22791);
xor U22917 (N_22917,N_22793,N_22614);
and U22918 (N_22918,N_22736,N_22699);
or U22919 (N_22919,N_22658,N_22769);
or U22920 (N_22920,N_22606,N_22679);
nand U22921 (N_22921,N_22645,N_22636);
nor U22922 (N_22922,N_22628,N_22798);
nor U22923 (N_22923,N_22731,N_22771);
nand U22924 (N_22924,N_22690,N_22739);
or U22925 (N_22925,N_22698,N_22695);
xor U22926 (N_22926,N_22653,N_22797);
nand U22927 (N_22927,N_22671,N_22676);
nand U22928 (N_22928,N_22618,N_22626);
nor U22929 (N_22929,N_22720,N_22788);
nor U22930 (N_22930,N_22647,N_22685);
xnor U22931 (N_22931,N_22724,N_22730);
nor U22932 (N_22932,N_22708,N_22799);
xnor U22933 (N_22933,N_22723,N_22612);
and U22934 (N_22934,N_22677,N_22621);
or U22935 (N_22935,N_22743,N_22748);
and U22936 (N_22936,N_22744,N_22687);
nand U22937 (N_22937,N_22703,N_22640);
nand U22938 (N_22938,N_22769,N_22627);
nand U22939 (N_22939,N_22770,N_22718);
nand U22940 (N_22940,N_22685,N_22723);
and U22941 (N_22941,N_22619,N_22600);
nor U22942 (N_22942,N_22674,N_22642);
nor U22943 (N_22943,N_22677,N_22620);
nand U22944 (N_22944,N_22779,N_22714);
or U22945 (N_22945,N_22651,N_22750);
and U22946 (N_22946,N_22780,N_22741);
or U22947 (N_22947,N_22753,N_22766);
and U22948 (N_22948,N_22767,N_22720);
and U22949 (N_22949,N_22795,N_22729);
xnor U22950 (N_22950,N_22758,N_22617);
nand U22951 (N_22951,N_22692,N_22774);
nand U22952 (N_22952,N_22737,N_22625);
xor U22953 (N_22953,N_22712,N_22633);
and U22954 (N_22954,N_22691,N_22627);
xnor U22955 (N_22955,N_22642,N_22600);
nor U22956 (N_22956,N_22630,N_22606);
or U22957 (N_22957,N_22639,N_22624);
nor U22958 (N_22958,N_22728,N_22693);
nand U22959 (N_22959,N_22756,N_22706);
xor U22960 (N_22960,N_22698,N_22646);
and U22961 (N_22961,N_22624,N_22763);
nand U22962 (N_22962,N_22646,N_22664);
and U22963 (N_22963,N_22775,N_22699);
and U22964 (N_22964,N_22624,N_22724);
and U22965 (N_22965,N_22756,N_22734);
or U22966 (N_22966,N_22689,N_22692);
and U22967 (N_22967,N_22682,N_22704);
nand U22968 (N_22968,N_22680,N_22763);
nand U22969 (N_22969,N_22608,N_22632);
or U22970 (N_22970,N_22761,N_22678);
xnor U22971 (N_22971,N_22712,N_22726);
or U22972 (N_22972,N_22791,N_22731);
or U22973 (N_22973,N_22630,N_22615);
nand U22974 (N_22974,N_22768,N_22682);
xor U22975 (N_22975,N_22783,N_22757);
xnor U22976 (N_22976,N_22705,N_22654);
nor U22977 (N_22977,N_22623,N_22784);
or U22978 (N_22978,N_22692,N_22651);
and U22979 (N_22979,N_22697,N_22717);
or U22980 (N_22980,N_22716,N_22654);
or U22981 (N_22981,N_22610,N_22791);
and U22982 (N_22982,N_22634,N_22657);
xnor U22983 (N_22983,N_22622,N_22709);
nand U22984 (N_22984,N_22722,N_22625);
nor U22985 (N_22985,N_22701,N_22623);
xnor U22986 (N_22986,N_22624,N_22615);
nand U22987 (N_22987,N_22717,N_22696);
and U22988 (N_22988,N_22683,N_22601);
and U22989 (N_22989,N_22658,N_22696);
xor U22990 (N_22990,N_22716,N_22633);
xor U22991 (N_22991,N_22764,N_22690);
and U22992 (N_22992,N_22640,N_22619);
nor U22993 (N_22993,N_22702,N_22762);
xor U22994 (N_22994,N_22625,N_22770);
and U22995 (N_22995,N_22670,N_22770);
xnor U22996 (N_22996,N_22693,N_22740);
nand U22997 (N_22997,N_22702,N_22680);
and U22998 (N_22998,N_22782,N_22611);
or U22999 (N_22999,N_22796,N_22789);
xor U23000 (N_23000,N_22874,N_22903);
or U23001 (N_23001,N_22930,N_22894);
and U23002 (N_23002,N_22837,N_22970);
xor U23003 (N_23003,N_22909,N_22927);
or U23004 (N_23004,N_22811,N_22917);
nand U23005 (N_23005,N_22934,N_22882);
or U23006 (N_23006,N_22900,N_22980);
and U23007 (N_23007,N_22905,N_22999);
or U23008 (N_23008,N_22820,N_22801);
and U23009 (N_23009,N_22857,N_22908);
or U23010 (N_23010,N_22924,N_22845);
xor U23011 (N_23011,N_22975,N_22869);
or U23012 (N_23012,N_22814,N_22942);
nand U23013 (N_23013,N_22881,N_22846);
or U23014 (N_23014,N_22863,N_22895);
and U23015 (N_23015,N_22870,N_22810);
and U23016 (N_23016,N_22952,N_22890);
nand U23017 (N_23017,N_22955,N_22947);
nor U23018 (N_23018,N_22834,N_22819);
or U23019 (N_23019,N_22974,N_22809);
nand U23020 (N_23020,N_22830,N_22827);
or U23021 (N_23021,N_22919,N_22828);
nor U23022 (N_23022,N_22914,N_22841);
or U23023 (N_23023,N_22944,N_22943);
and U23024 (N_23024,N_22893,N_22899);
and U23025 (N_23025,N_22864,N_22994);
and U23026 (N_23026,N_22860,N_22879);
xnor U23027 (N_23027,N_22997,N_22978);
nor U23028 (N_23028,N_22992,N_22995);
nor U23029 (N_23029,N_22902,N_22824);
nand U23030 (N_23030,N_22948,N_22812);
nor U23031 (N_23031,N_22865,N_22853);
nor U23032 (N_23032,N_22805,N_22977);
and U23033 (N_23033,N_22911,N_22958);
xnor U23034 (N_23034,N_22949,N_22898);
and U23035 (N_23035,N_22959,N_22872);
and U23036 (N_23036,N_22907,N_22804);
or U23037 (N_23037,N_22839,N_22962);
nand U23038 (N_23038,N_22968,N_22877);
nor U23039 (N_23039,N_22876,N_22953);
nand U23040 (N_23040,N_22913,N_22951);
or U23041 (N_23041,N_22939,N_22825);
and U23042 (N_23042,N_22843,N_22896);
nand U23043 (N_23043,N_22831,N_22973);
nor U23044 (N_23044,N_22840,N_22883);
and U23045 (N_23045,N_22996,N_22813);
nand U23046 (N_23046,N_22929,N_22802);
nor U23047 (N_23047,N_22868,N_22931);
nor U23048 (N_23048,N_22842,N_22822);
or U23049 (N_23049,N_22885,N_22983);
or U23050 (N_23050,N_22928,N_22850);
nor U23051 (N_23051,N_22847,N_22904);
xnor U23052 (N_23052,N_22818,N_22817);
nand U23053 (N_23053,N_22856,N_22960);
xnor U23054 (N_23054,N_22887,N_22932);
nor U23055 (N_23055,N_22862,N_22815);
nand U23056 (N_23056,N_22915,N_22852);
or U23057 (N_23057,N_22910,N_22961);
or U23058 (N_23058,N_22901,N_22984);
and U23059 (N_23059,N_22867,N_22963);
nand U23060 (N_23060,N_22821,N_22967);
nand U23061 (N_23061,N_22981,N_22964);
nand U23062 (N_23062,N_22807,N_22855);
nor U23063 (N_23063,N_22888,N_22803);
and U23064 (N_23064,N_22991,N_22806);
xnor U23065 (N_23065,N_22808,N_22940);
nand U23066 (N_23066,N_22848,N_22859);
xnor U23067 (N_23067,N_22954,N_22880);
xor U23068 (N_23068,N_22826,N_22987);
xor U23069 (N_23069,N_22912,N_22971);
nand U23070 (N_23070,N_22993,N_22936);
or U23071 (N_23071,N_22937,N_22886);
nor U23072 (N_23072,N_22851,N_22823);
nand U23073 (N_23073,N_22941,N_22921);
and U23074 (N_23074,N_22878,N_22982);
or U23075 (N_23075,N_22926,N_22989);
or U23076 (N_23076,N_22935,N_22950);
and U23077 (N_23077,N_22829,N_22891);
and U23078 (N_23078,N_22844,N_22972);
xor U23079 (N_23079,N_22998,N_22836);
and U23080 (N_23080,N_22849,N_22922);
and U23081 (N_23081,N_22892,N_22835);
xor U23082 (N_23082,N_22906,N_22925);
nor U23083 (N_23083,N_22838,N_22985);
nor U23084 (N_23084,N_22988,N_22889);
xnor U23085 (N_23085,N_22875,N_22832);
or U23086 (N_23086,N_22873,N_22866);
and U23087 (N_23087,N_22816,N_22854);
or U23088 (N_23088,N_22923,N_22871);
nor U23089 (N_23089,N_22986,N_22916);
xor U23090 (N_23090,N_22858,N_22800);
and U23091 (N_23091,N_22920,N_22966);
or U23092 (N_23092,N_22945,N_22918);
nor U23093 (N_23093,N_22861,N_22946);
nor U23094 (N_23094,N_22965,N_22933);
and U23095 (N_23095,N_22938,N_22884);
and U23096 (N_23096,N_22956,N_22897);
xor U23097 (N_23097,N_22969,N_22976);
nor U23098 (N_23098,N_22990,N_22833);
xnor U23099 (N_23099,N_22957,N_22979);
nand U23100 (N_23100,N_22819,N_22966);
and U23101 (N_23101,N_22875,N_22846);
and U23102 (N_23102,N_22808,N_22905);
xor U23103 (N_23103,N_22862,N_22914);
nor U23104 (N_23104,N_22849,N_22857);
nor U23105 (N_23105,N_22893,N_22878);
nor U23106 (N_23106,N_22824,N_22961);
xor U23107 (N_23107,N_22905,N_22860);
nor U23108 (N_23108,N_22891,N_22939);
nor U23109 (N_23109,N_22979,N_22864);
and U23110 (N_23110,N_22934,N_22802);
nor U23111 (N_23111,N_22844,N_22994);
nor U23112 (N_23112,N_22883,N_22929);
nor U23113 (N_23113,N_22856,N_22803);
nand U23114 (N_23114,N_22978,N_22829);
or U23115 (N_23115,N_22851,N_22998);
xor U23116 (N_23116,N_22921,N_22960);
xor U23117 (N_23117,N_22841,N_22984);
nand U23118 (N_23118,N_22993,N_22977);
nand U23119 (N_23119,N_22947,N_22802);
nor U23120 (N_23120,N_22949,N_22844);
or U23121 (N_23121,N_22896,N_22807);
xnor U23122 (N_23122,N_22899,N_22977);
or U23123 (N_23123,N_22875,N_22959);
or U23124 (N_23124,N_22855,N_22835);
nand U23125 (N_23125,N_22812,N_22878);
or U23126 (N_23126,N_22851,N_22873);
nor U23127 (N_23127,N_22841,N_22898);
nand U23128 (N_23128,N_22954,N_22903);
nor U23129 (N_23129,N_22891,N_22819);
or U23130 (N_23130,N_22836,N_22858);
or U23131 (N_23131,N_22963,N_22859);
nand U23132 (N_23132,N_22936,N_22867);
and U23133 (N_23133,N_22876,N_22822);
nor U23134 (N_23134,N_22943,N_22989);
nor U23135 (N_23135,N_22975,N_22840);
nor U23136 (N_23136,N_22981,N_22929);
xor U23137 (N_23137,N_22897,N_22826);
and U23138 (N_23138,N_22925,N_22816);
or U23139 (N_23139,N_22946,N_22875);
and U23140 (N_23140,N_22869,N_22880);
xor U23141 (N_23141,N_22808,N_22914);
nand U23142 (N_23142,N_22875,N_22867);
and U23143 (N_23143,N_22891,N_22856);
nand U23144 (N_23144,N_22996,N_22875);
xnor U23145 (N_23145,N_22910,N_22851);
or U23146 (N_23146,N_22926,N_22928);
and U23147 (N_23147,N_22958,N_22816);
nand U23148 (N_23148,N_22883,N_22932);
xnor U23149 (N_23149,N_22850,N_22803);
xnor U23150 (N_23150,N_22870,N_22957);
or U23151 (N_23151,N_22983,N_22912);
xnor U23152 (N_23152,N_22851,N_22820);
or U23153 (N_23153,N_22848,N_22985);
nand U23154 (N_23154,N_22812,N_22976);
nand U23155 (N_23155,N_22966,N_22924);
or U23156 (N_23156,N_22942,N_22880);
xor U23157 (N_23157,N_22950,N_22802);
xor U23158 (N_23158,N_22961,N_22825);
nor U23159 (N_23159,N_22903,N_22850);
nor U23160 (N_23160,N_22803,N_22810);
nor U23161 (N_23161,N_22911,N_22851);
or U23162 (N_23162,N_22805,N_22953);
xor U23163 (N_23163,N_22901,N_22945);
xor U23164 (N_23164,N_22850,N_22971);
nand U23165 (N_23165,N_22805,N_22886);
xnor U23166 (N_23166,N_22863,N_22860);
and U23167 (N_23167,N_22942,N_22812);
xnor U23168 (N_23168,N_22821,N_22908);
nor U23169 (N_23169,N_22952,N_22921);
nand U23170 (N_23170,N_22864,N_22802);
and U23171 (N_23171,N_22859,N_22890);
or U23172 (N_23172,N_22975,N_22838);
nand U23173 (N_23173,N_22816,N_22857);
and U23174 (N_23174,N_22838,N_22992);
xnor U23175 (N_23175,N_22813,N_22853);
and U23176 (N_23176,N_22872,N_22880);
or U23177 (N_23177,N_22826,N_22845);
or U23178 (N_23178,N_22854,N_22892);
or U23179 (N_23179,N_22838,N_22935);
or U23180 (N_23180,N_22879,N_22912);
or U23181 (N_23181,N_22942,N_22990);
nand U23182 (N_23182,N_22812,N_22907);
nand U23183 (N_23183,N_22917,N_22882);
nor U23184 (N_23184,N_22949,N_22890);
nor U23185 (N_23185,N_22876,N_22815);
nand U23186 (N_23186,N_22929,N_22906);
nand U23187 (N_23187,N_22829,N_22981);
nor U23188 (N_23188,N_22826,N_22853);
nand U23189 (N_23189,N_22871,N_22809);
or U23190 (N_23190,N_22877,N_22826);
xnor U23191 (N_23191,N_22975,N_22906);
nand U23192 (N_23192,N_22910,N_22879);
and U23193 (N_23193,N_22889,N_22891);
nand U23194 (N_23194,N_22898,N_22943);
or U23195 (N_23195,N_22867,N_22856);
nor U23196 (N_23196,N_22986,N_22908);
xnor U23197 (N_23197,N_22953,N_22874);
or U23198 (N_23198,N_22833,N_22883);
xnor U23199 (N_23199,N_22938,N_22924);
nand U23200 (N_23200,N_23171,N_23056);
nand U23201 (N_23201,N_23191,N_23125);
xor U23202 (N_23202,N_23166,N_23022);
xnor U23203 (N_23203,N_23088,N_23048);
xnor U23204 (N_23204,N_23103,N_23114);
nor U23205 (N_23205,N_23004,N_23001);
nand U23206 (N_23206,N_23117,N_23130);
nor U23207 (N_23207,N_23160,N_23055);
nor U23208 (N_23208,N_23159,N_23014);
xor U23209 (N_23209,N_23184,N_23134);
nor U23210 (N_23210,N_23100,N_23116);
or U23211 (N_23211,N_23192,N_23082);
and U23212 (N_23212,N_23172,N_23008);
nor U23213 (N_23213,N_23158,N_23106);
nand U23214 (N_23214,N_23046,N_23009);
xnor U23215 (N_23215,N_23075,N_23040);
nand U23216 (N_23216,N_23176,N_23094);
and U23217 (N_23217,N_23012,N_23156);
xnor U23218 (N_23218,N_23149,N_23121);
nand U23219 (N_23219,N_23150,N_23029);
nand U23220 (N_23220,N_23146,N_23143);
nand U23221 (N_23221,N_23070,N_23078);
or U23222 (N_23222,N_23093,N_23021);
and U23223 (N_23223,N_23127,N_23036);
and U23224 (N_23224,N_23039,N_23085);
nand U23225 (N_23225,N_23144,N_23193);
xnor U23226 (N_23226,N_23024,N_23069);
nor U23227 (N_23227,N_23089,N_23054);
or U23228 (N_23228,N_23157,N_23161);
nand U23229 (N_23229,N_23140,N_23076);
nor U23230 (N_23230,N_23187,N_23181);
nor U23231 (N_23231,N_23002,N_23135);
or U23232 (N_23232,N_23113,N_23091);
nor U23233 (N_23233,N_23141,N_23136);
or U23234 (N_23234,N_23190,N_23047);
and U23235 (N_23235,N_23197,N_23132);
or U23236 (N_23236,N_23018,N_23077);
or U23237 (N_23237,N_23068,N_23053);
and U23238 (N_23238,N_23196,N_23174);
and U23239 (N_23239,N_23183,N_23169);
or U23240 (N_23240,N_23118,N_23063);
xor U23241 (N_23241,N_23058,N_23071);
xnor U23242 (N_23242,N_23126,N_23119);
xor U23243 (N_23243,N_23179,N_23010);
or U23244 (N_23244,N_23067,N_23005);
or U23245 (N_23245,N_23188,N_23017);
and U23246 (N_23246,N_23041,N_23026);
and U23247 (N_23247,N_23170,N_23168);
and U23248 (N_23248,N_23045,N_23123);
or U23249 (N_23249,N_23097,N_23111);
nand U23250 (N_23250,N_23139,N_23198);
nor U23251 (N_23251,N_23037,N_23073);
or U23252 (N_23252,N_23112,N_23066);
xnor U23253 (N_23253,N_23115,N_23105);
nand U23254 (N_23254,N_23007,N_23072);
nand U23255 (N_23255,N_23081,N_23133);
xor U23256 (N_23256,N_23084,N_23167);
or U23257 (N_23257,N_23052,N_23060);
nor U23258 (N_23258,N_23110,N_23199);
or U23259 (N_23259,N_23064,N_23178);
or U23260 (N_23260,N_23180,N_23092);
nand U23261 (N_23261,N_23107,N_23099);
xor U23262 (N_23262,N_23104,N_23173);
or U23263 (N_23263,N_23131,N_23023);
xnor U23264 (N_23264,N_23163,N_23087);
and U23265 (N_23265,N_23154,N_23050);
xnor U23266 (N_23266,N_23033,N_23011);
or U23267 (N_23267,N_23030,N_23015);
nand U23268 (N_23268,N_23080,N_23034);
or U23269 (N_23269,N_23098,N_23020);
or U23270 (N_23270,N_23152,N_23162);
nand U23271 (N_23271,N_23186,N_23177);
or U23272 (N_23272,N_23000,N_23101);
nand U23273 (N_23273,N_23095,N_23025);
and U23274 (N_23274,N_23155,N_23148);
nand U23275 (N_23275,N_23016,N_23194);
nor U23276 (N_23276,N_23128,N_23027);
nand U23277 (N_23277,N_23043,N_23090);
nor U23278 (N_23278,N_23138,N_23153);
nor U23279 (N_23279,N_23142,N_23044);
xnor U23280 (N_23280,N_23108,N_23096);
nand U23281 (N_23281,N_23074,N_23065);
nand U23282 (N_23282,N_23129,N_23061);
nor U23283 (N_23283,N_23185,N_23147);
and U23284 (N_23284,N_23120,N_23189);
or U23285 (N_23285,N_23062,N_23019);
nor U23286 (N_23286,N_23109,N_23079);
or U23287 (N_23287,N_23195,N_23013);
xor U23288 (N_23288,N_23032,N_23049);
nand U23289 (N_23289,N_23124,N_23122);
and U23290 (N_23290,N_23137,N_23028);
nor U23291 (N_23291,N_23086,N_23059);
xor U23292 (N_23292,N_23175,N_23035);
nor U23293 (N_23293,N_23051,N_23145);
nand U23294 (N_23294,N_23042,N_23165);
nand U23295 (N_23295,N_23164,N_23182);
nand U23296 (N_23296,N_23031,N_23083);
and U23297 (N_23297,N_23151,N_23003);
nand U23298 (N_23298,N_23102,N_23038);
xor U23299 (N_23299,N_23006,N_23057);
xor U23300 (N_23300,N_23085,N_23175);
and U23301 (N_23301,N_23024,N_23185);
nor U23302 (N_23302,N_23077,N_23175);
xor U23303 (N_23303,N_23041,N_23112);
xnor U23304 (N_23304,N_23148,N_23199);
and U23305 (N_23305,N_23155,N_23072);
and U23306 (N_23306,N_23155,N_23181);
and U23307 (N_23307,N_23176,N_23156);
and U23308 (N_23308,N_23094,N_23199);
nand U23309 (N_23309,N_23180,N_23010);
nand U23310 (N_23310,N_23131,N_23153);
nor U23311 (N_23311,N_23149,N_23155);
and U23312 (N_23312,N_23040,N_23094);
nand U23313 (N_23313,N_23134,N_23137);
xnor U23314 (N_23314,N_23115,N_23165);
nand U23315 (N_23315,N_23179,N_23118);
nand U23316 (N_23316,N_23012,N_23155);
and U23317 (N_23317,N_23066,N_23143);
nand U23318 (N_23318,N_23115,N_23059);
or U23319 (N_23319,N_23051,N_23080);
nand U23320 (N_23320,N_23085,N_23151);
nor U23321 (N_23321,N_23009,N_23005);
xor U23322 (N_23322,N_23029,N_23023);
nor U23323 (N_23323,N_23139,N_23157);
and U23324 (N_23324,N_23179,N_23133);
or U23325 (N_23325,N_23019,N_23023);
xnor U23326 (N_23326,N_23143,N_23078);
xor U23327 (N_23327,N_23109,N_23158);
xnor U23328 (N_23328,N_23097,N_23140);
and U23329 (N_23329,N_23166,N_23044);
and U23330 (N_23330,N_23093,N_23144);
xnor U23331 (N_23331,N_23060,N_23021);
and U23332 (N_23332,N_23049,N_23071);
and U23333 (N_23333,N_23102,N_23166);
nor U23334 (N_23334,N_23154,N_23037);
xnor U23335 (N_23335,N_23134,N_23027);
nand U23336 (N_23336,N_23134,N_23136);
nand U23337 (N_23337,N_23107,N_23149);
nor U23338 (N_23338,N_23056,N_23055);
and U23339 (N_23339,N_23068,N_23037);
nand U23340 (N_23340,N_23080,N_23196);
or U23341 (N_23341,N_23105,N_23166);
nor U23342 (N_23342,N_23025,N_23087);
nand U23343 (N_23343,N_23043,N_23072);
nor U23344 (N_23344,N_23176,N_23129);
or U23345 (N_23345,N_23042,N_23001);
or U23346 (N_23346,N_23044,N_23199);
nor U23347 (N_23347,N_23010,N_23063);
or U23348 (N_23348,N_23108,N_23106);
xnor U23349 (N_23349,N_23199,N_23020);
xnor U23350 (N_23350,N_23094,N_23074);
and U23351 (N_23351,N_23152,N_23169);
and U23352 (N_23352,N_23119,N_23144);
nor U23353 (N_23353,N_23025,N_23069);
and U23354 (N_23354,N_23100,N_23073);
and U23355 (N_23355,N_23110,N_23125);
nand U23356 (N_23356,N_23131,N_23172);
xnor U23357 (N_23357,N_23028,N_23027);
nand U23358 (N_23358,N_23162,N_23155);
and U23359 (N_23359,N_23180,N_23138);
or U23360 (N_23360,N_23029,N_23140);
nor U23361 (N_23361,N_23122,N_23089);
and U23362 (N_23362,N_23150,N_23071);
nand U23363 (N_23363,N_23079,N_23005);
or U23364 (N_23364,N_23107,N_23012);
and U23365 (N_23365,N_23118,N_23099);
nand U23366 (N_23366,N_23177,N_23087);
nand U23367 (N_23367,N_23062,N_23114);
xor U23368 (N_23368,N_23067,N_23115);
nor U23369 (N_23369,N_23025,N_23163);
or U23370 (N_23370,N_23063,N_23188);
nor U23371 (N_23371,N_23114,N_23006);
nor U23372 (N_23372,N_23117,N_23177);
and U23373 (N_23373,N_23060,N_23024);
and U23374 (N_23374,N_23182,N_23124);
xnor U23375 (N_23375,N_23062,N_23098);
nand U23376 (N_23376,N_23022,N_23094);
xor U23377 (N_23377,N_23113,N_23176);
nor U23378 (N_23378,N_23076,N_23007);
or U23379 (N_23379,N_23035,N_23010);
and U23380 (N_23380,N_23025,N_23046);
or U23381 (N_23381,N_23052,N_23018);
nor U23382 (N_23382,N_23143,N_23133);
xor U23383 (N_23383,N_23112,N_23073);
nand U23384 (N_23384,N_23019,N_23037);
nor U23385 (N_23385,N_23194,N_23139);
nand U23386 (N_23386,N_23152,N_23187);
nand U23387 (N_23387,N_23071,N_23075);
or U23388 (N_23388,N_23109,N_23095);
xnor U23389 (N_23389,N_23164,N_23144);
nand U23390 (N_23390,N_23148,N_23174);
nand U23391 (N_23391,N_23001,N_23113);
and U23392 (N_23392,N_23129,N_23053);
nand U23393 (N_23393,N_23061,N_23079);
or U23394 (N_23394,N_23152,N_23046);
and U23395 (N_23395,N_23170,N_23010);
xor U23396 (N_23396,N_23098,N_23174);
and U23397 (N_23397,N_23181,N_23140);
xor U23398 (N_23398,N_23184,N_23060);
and U23399 (N_23399,N_23138,N_23128);
xor U23400 (N_23400,N_23275,N_23376);
or U23401 (N_23401,N_23348,N_23353);
xnor U23402 (N_23402,N_23207,N_23318);
nor U23403 (N_23403,N_23385,N_23242);
or U23404 (N_23404,N_23313,N_23341);
nor U23405 (N_23405,N_23265,N_23260);
and U23406 (N_23406,N_23241,N_23303);
or U23407 (N_23407,N_23309,N_23230);
and U23408 (N_23408,N_23226,N_23238);
and U23409 (N_23409,N_23356,N_23363);
or U23410 (N_23410,N_23384,N_23377);
or U23411 (N_23411,N_23335,N_23306);
and U23412 (N_23412,N_23219,N_23244);
and U23413 (N_23413,N_23327,N_23394);
or U23414 (N_23414,N_23217,N_23317);
xor U23415 (N_23415,N_23311,N_23331);
nand U23416 (N_23416,N_23337,N_23220);
xnor U23417 (N_23417,N_23386,N_23261);
nand U23418 (N_23418,N_23395,N_23300);
xor U23419 (N_23419,N_23332,N_23235);
nor U23420 (N_23420,N_23323,N_23285);
nand U23421 (N_23421,N_23329,N_23398);
or U23422 (N_23422,N_23279,N_23228);
nand U23423 (N_23423,N_23328,N_23322);
nor U23424 (N_23424,N_23283,N_23375);
xnor U23425 (N_23425,N_23397,N_23245);
or U23426 (N_23426,N_23202,N_23209);
nor U23427 (N_23427,N_23307,N_23326);
or U23428 (N_23428,N_23299,N_23374);
nand U23429 (N_23429,N_23264,N_23369);
and U23430 (N_23430,N_23297,N_23308);
nor U23431 (N_23431,N_23276,N_23214);
nand U23432 (N_23432,N_23254,N_23380);
and U23433 (N_23433,N_23273,N_23298);
and U23434 (N_23434,N_23312,N_23268);
xnor U23435 (N_23435,N_23231,N_23240);
nand U23436 (N_23436,N_23381,N_23382);
nand U23437 (N_23437,N_23224,N_23349);
or U23438 (N_23438,N_23347,N_23295);
nand U23439 (N_23439,N_23345,N_23250);
and U23440 (N_23440,N_23371,N_23296);
nor U23441 (N_23441,N_23350,N_23291);
xnor U23442 (N_23442,N_23200,N_23215);
and U23443 (N_23443,N_23257,N_23229);
nand U23444 (N_23444,N_23271,N_23222);
nor U23445 (N_23445,N_23304,N_23262);
xor U23446 (N_23446,N_23243,N_23278);
and U23447 (N_23447,N_23216,N_23320);
or U23448 (N_23448,N_23390,N_23340);
or U23449 (N_23449,N_23388,N_23379);
and U23450 (N_23450,N_23365,N_23396);
nand U23451 (N_23451,N_23355,N_23359);
nor U23452 (N_23452,N_23334,N_23248);
and U23453 (N_23453,N_23346,N_23204);
and U23454 (N_23454,N_23301,N_23258);
and U23455 (N_23455,N_23330,N_23269);
nor U23456 (N_23456,N_23344,N_23360);
nand U23457 (N_23457,N_23256,N_23373);
nand U23458 (N_23458,N_23358,N_23206);
nor U23459 (N_23459,N_23266,N_23284);
xnor U23460 (N_23460,N_23366,N_23251);
or U23461 (N_23461,N_23253,N_23393);
nand U23462 (N_23462,N_23259,N_23293);
and U23463 (N_23463,N_23392,N_23274);
or U23464 (N_23464,N_23290,N_23399);
nor U23465 (N_23465,N_23247,N_23236);
nand U23466 (N_23466,N_23315,N_23368);
nor U23467 (N_23467,N_23249,N_23294);
nor U23468 (N_23468,N_23316,N_23367);
nand U23469 (N_23469,N_23281,N_23333);
xnor U23470 (N_23470,N_23343,N_23339);
xor U23471 (N_23471,N_23282,N_23305);
xnor U23472 (N_23472,N_23223,N_23225);
nand U23473 (N_23473,N_23352,N_23314);
and U23474 (N_23474,N_23232,N_23210);
nand U23475 (N_23475,N_23213,N_23211);
nand U23476 (N_23476,N_23391,N_23288);
nand U23477 (N_23477,N_23234,N_23389);
nor U23478 (N_23478,N_23205,N_23372);
nand U23479 (N_23479,N_23324,N_23272);
nor U23480 (N_23480,N_23218,N_23287);
xnor U23481 (N_23481,N_23201,N_23321);
or U23482 (N_23482,N_23233,N_23227);
nand U23483 (N_23483,N_23255,N_23357);
nor U23484 (N_23484,N_23208,N_23263);
nand U23485 (N_23485,N_23203,N_23338);
nor U23486 (N_23486,N_23280,N_23212);
xor U23487 (N_23487,N_23286,N_23361);
nand U23488 (N_23488,N_23292,N_23246);
nor U23489 (N_23489,N_23351,N_23354);
or U23490 (N_23490,N_23362,N_23336);
nor U23491 (N_23491,N_23342,N_23364);
and U23492 (N_23492,N_23387,N_23383);
and U23493 (N_23493,N_23370,N_23221);
or U23494 (N_23494,N_23310,N_23237);
or U23495 (N_23495,N_23289,N_23277);
and U23496 (N_23496,N_23252,N_23325);
nand U23497 (N_23497,N_23378,N_23270);
nand U23498 (N_23498,N_23239,N_23302);
or U23499 (N_23499,N_23319,N_23267);
nor U23500 (N_23500,N_23319,N_23398);
or U23501 (N_23501,N_23207,N_23370);
or U23502 (N_23502,N_23205,N_23391);
nand U23503 (N_23503,N_23356,N_23200);
nand U23504 (N_23504,N_23306,N_23333);
nand U23505 (N_23505,N_23381,N_23205);
and U23506 (N_23506,N_23322,N_23321);
or U23507 (N_23507,N_23351,N_23293);
nor U23508 (N_23508,N_23260,N_23331);
xnor U23509 (N_23509,N_23220,N_23316);
nand U23510 (N_23510,N_23307,N_23303);
and U23511 (N_23511,N_23335,N_23283);
nor U23512 (N_23512,N_23326,N_23273);
nand U23513 (N_23513,N_23372,N_23223);
nand U23514 (N_23514,N_23229,N_23263);
nand U23515 (N_23515,N_23297,N_23367);
nand U23516 (N_23516,N_23336,N_23343);
nand U23517 (N_23517,N_23302,N_23370);
nor U23518 (N_23518,N_23209,N_23273);
and U23519 (N_23519,N_23238,N_23202);
nand U23520 (N_23520,N_23206,N_23283);
and U23521 (N_23521,N_23298,N_23294);
xor U23522 (N_23522,N_23225,N_23231);
nor U23523 (N_23523,N_23288,N_23310);
nand U23524 (N_23524,N_23363,N_23393);
or U23525 (N_23525,N_23252,N_23319);
and U23526 (N_23526,N_23314,N_23268);
nor U23527 (N_23527,N_23309,N_23335);
xor U23528 (N_23528,N_23356,N_23215);
or U23529 (N_23529,N_23233,N_23210);
nand U23530 (N_23530,N_23384,N_23309);
and U23531 (N_23531,N_23233,N_23243);
xnor U23532 (N_23532,N_23223,N_23224);
xor U23533 (N_23533,N_23242,N_23235);
and U23534 (N_23534,N_23360,N_23307);
or U23535 (N_23535,N_23208,N_23257);
or U23536 (N_23536,N_23259,N_23330);
nor U23537 (N_23537,N_23252,N_23372);
or U23538 (N_23538,N_23240,N_23397);
nor U23539 (N_23539,N_23374,N_23373);
nand U23540 (N_23540,N_23387,N_23302);
or U23541 (N_23541,N_23288,N_23201);
or U23542 (N_23542,N_23301,N_23272);
xor U23543 (N_23543,N_23361,N_23337);
and U23544 (N_23544,N_23280,N_23299);
and U23545 (N_23545,N_23366,N_23215);
and U23546 (N_23546,N_23243,N_23323);
nor U23547 (N_23547,N_23393,N_23230);
nor U23548 (N_23548,N_23272,N_23338);
nor U23549 (N_23549,N_23231,N_23396);
nand U23550 (N_23550,N_23257,N_23399);
nor U23551 (N_23551,N_23350,N_23395);
or U23552 (N_23552,N_23240,N_23385);
and U23553 (N_23553,N_23331,N_23388);
xnor U23554 (N_23554,N_23278,N_23349);
or U23555 (N_23555,N_23213,N_23291);
or U23556 (N_23556,N_23322,N_23256);
nand U23557 (N_23557,N_23319,N_23363);
xnor U23558 (N_23558,N_23204,N_23307);
nand U23559 (N_23559,N_23299,N_23259);
or U23560 (N_23560,N_23275,N_23223);
xor U23561 (N_23561,N_23329,N_23337);
nand U23562 (N_23562,N_23212,N_23237);
or U23563 (N_23563,N_23216,N_23265);
nand U23564 (N_23564,N_23256,N_23389);
or U23565 (N_23565,N_23387,N_23210);
and U23566 (N_23566,N_23286,N_23340);
nand U23567 (N_23567,N_23383,N_23281);
nor U23568 (N_23568,N_23329,N_23394);
nand U23569 (N_23569,N_23372,N_23203);
and U23570 (N_23570,N_23376,N_23281);
and U23571 (N_23571,N_23330,N_23395);
nand U23572 (N_23572,N_23364,N_23210);
xnor U23573 (N_23573,N_23223,N_23244);
nand U23574 (N_23574,N_23323,N_23341);
or U23575 (N_23575,N_23293,N_23283);
and U23576 (N_23576,N_23307,N_23304);
and U23577 (N_23577,N_23273,N_23328);
nor U23578 (N_23578,N_23341,N_23216);
nor U23579 (N_23579,N_23371,N_23372);
xor U23580 (N_23580,N_23294,N_23301);
nor U23581 (N_23581,N_23288,N_23232);
xor U23582 (N_23582,N_23269,N_23275);
or U23583 (N_23583,N_23318,N_23209);
xor U23584 (N_23584,N_23325,N_23322);
and U23585 (N_23585,N_23337,N_23286);
nand U23586 (N_23586,N_23246,N_23261);
nor U23587 (N_23587,N_23248,N_23290);
xor U23588 (N_23588,N_23384,N_23307);
xor U23589 (N_23589,N_23254,N_23313);
nand U23590 (N_23590,N_23288,N_23210);
xor U23591 (N_23591,N_23310,N_23264);
xnor U23592 (N_23592,N_23312,N_23260);
nor U23593 (N_23593,N_23323,N_23344);
nand U23594 (N_23594,N_23329,N_23304);
nand U23595 (N_23595,N_23200,N_23222);
xor U23596 (N_23596,N_23217,N_23221);
nor U23597 (N_23597,N_23331,N_23309);
nor U23598 (N_23598,N_23282,N_23274);
nor U23599 (N_23599,N_23239,N_23354);
xnor U23600 (N_23600,N_23562,N_23529);
or U23601 (N_23601,N_23559,N_23571);
nand U23602 (N_23602,N_23538,N_23414);
nand U23603 (N_23603,N_23478,N_23541);
nor U23604 (N_23604,N_23570,N_23532);
nor U23605 (N_23605,N_23425,N_23530);
xnor U23606 (N_23606,N_23464,N_23577);
nor U23607 (N_23607,N_23508,N_23552);
xor U23608 (N_23608,N_23515,N_23543);
nand U23609 (N_23609,N_23462,N_23485);
nand U23610 (N_23610,N_23423,N_23506);
or U23611 (N_23611,N_23525,N_23493);
xnor U23612 (N_23612,N_23488,N_23522);
xor U23613 (N_23613,N_23431,N_23470);
nor U23614 (N_23614,N_23547,N_23411);
nor U23615 (N_23615,N_23434,N_23560);
and U23616 (N_23616,N_23561,N_23444);
xor U23617 (N_23617,N_23535,N_23401);
and U23618 (N_23618,N_23494,N_23520);
nand U23619 (N_23619,N_23569,N_23474);
xor U23620 (N_23620,N_23573,N_23564);
xor U23621 (N_23621,N_23578,N_23443);
xor U23622 (N_23622,N_23481,N_23580);
nor U23623 (N_23623,N_23459,N_23471);
and U23624 (N_23624,N_23551,N_23461);
xnor U23625 (N_23625,N_23429,N_23499);
and U23626 (N_23626,N_23534,N_23544);
nor U23627 (N_23627,N_23589,N_23445);
and U23628 (N_23628,N_23507,N_23588);
xnor U23629 (N_23629,N_23486,N_23505);
or U23630 (N_23630,N_23512,N_23468);
or U23631 (N_23631,N_23587,N_23574);
nand U23632 (N_23632,N_23540,N_23526);
and U23633 (N_23633,N_23482,N_23550);
nand U23634 (N_23634,N_23473,N_23579);
xor U23635 (N_23635,N_23422,N_23413);
or U23636 (N_23636,N_23483,N_23477);
xnor U23637 (N_23637,N_23583,N_23558);
and U23638 (N_23638,N_23491,N_23517);
nand U23639 (N_23639,N_23406,N_23492);
nor U23640 (N_23640,N_23537,N_23426);
and U23641 (N_23641,N_23595,N_23451);
nand U23642 (N_23642,N_23518,N_23545);
or U23643 (N_23643,N_23584,N_23453);
nand U23644 (N_23644,N_23496,N_23549);
nand U23645 (N_23645,N_23500,N_23501);
xor U23646 (N_23646,N_23527,N_23412);
nor U23647 (N_23647,N_23441,N_23598);
nor U23648 (N_23648,N_23565,N_23465);
or U23649 (N_23649,N_23591,N_23430);
nand U23650 (N_23650,N_23460,N_23456);
xor U23651 (N_23651,N_23438,N_23531);
and U23652 (N_23652,N_23514,N_23480);
nor U23653 (N_23653,N_23467,N_23419);
nand U23654 (N_23654,N_23436,N_23400);
and U23655 (N_23655,N_23524,N_23585);
or U23656 (N_23656,N_23509,N_23404);
and U23657 (N_23657,N_23502,N_23557);
nand U23658 (N_23658,N_23446,N_23592);
nand U23659 (N_23659,N_23567,N_23432);
nor U23660 (N_23660,N_23513,N_23407);
nand U23661 (N_23661,N_23463,N_23542);
xnor U23662 (N_23662,N_23476,N_23568);
nor U23663 (N_23663,N_23455,N_23572);
nor U23664 (N_23664,N_23408,N_23487);
or U23665 (N_23665,N_23575,N_23566);
nor U23666 (N_23666,N_23586,N_23458);
and U23667 (N_23667,N_23452,N_23553);
nand U23668 (N_23668,N_23511,N_23490);
or U23669 (N_23669,N_23440,N_23439);
xor U23670 (N_23670,N_23475,N_23448);
and U23671 (N_23671,N_23597,N_23405);
nand U23672 (N_23672,N_23497,N_23555);
or U23673 (N_23673,N_23489,N_23554);
and U23674 (N_23674,N_23528,N_23437);
and U23675 (N_23675,N_23403,N_23433);
or U23676 (N_23676,N_23417,N_23420);
nand U23677 (N_23677,N_23447,N_23576);
nor U23678 (N_23678,N_23449,N_23536);
and U23679 (N_23679,N_23428,N_23410);
nand U23680 (N_23680,N_23498,N_23548);
xor U23681 (N_23681,N_23556,N_23450);
nand U23682 (N_23682,N_23454,N_23539);
and U23683 (N_23683,N_23479,N_23442);
and U23684 (N_23684,N_23590,N_23519);
nor U23685 (N_23685,N_23495,N_23472);
or U23686 (N_23686,N_23457,N_23503);
nor U23687 (N_23687,N_23415,N_23599);
nand U23688 (N_23688,N_23546,N_23469);
or U23689 (N_23689,N_23593,N_23504);
nor U23690 (N_23690,N_23581,N_23402);
xnor U23691 (N_23691,N_23582,N_23421);
nor U23692 (N_23692,N_23596,N_23466);
nor U23693 (N_23693,N_23523,N_23563);
or U23694 (N_23694,N_23416,N_23418);
nand U23695 (N_23695,N_23484,N_23424);
or U23696 (N_23696,N_23594,N_23409);
nand U23697 (N_23697,N_23533,N_23435);
nor U23698 (N_23698,N_23516,N_23427);
nor U23699 (N_23699,N_23521,N_23510);
or U23700 (N_23700,N_23480,N_23543);
or U23701 (N_23701,N_23586,N_23412);
xor U23702 (N_23702,N_23459,N_23488);
or U23703 (N_23703,N_23503,N_23480);
nor U23704 (N_23704,N_23458,N_23590);
xor U23705 (N_23705,N_23460,N_23565);
nand U23706 (N_23706,N_23585,N_23511);
and U23707 (N_23707,N_23561,N_23481);
nand U23708 (N_23708,N_23415,N_23584);
nand U23709 (N_23709,N_23526,N_23575);
nand U23710 (N_23710,N_23403,N_23435);
nor U23711 (N_23711,N_23564,N_23462);
nand U23712 (N_23712,N_23470,N_23500);
nor U23713 (N_23713,N_23454,N_23536);
nand U23714 (N_23714,N_23417,N_23533);
xnor U23715 (N_23715,N_23540,N_23405);
and U23716 (N_23716,N_23504,N_23403);
xor U23717 (N_23717,N_23585,N_23442);
nor U23718 (N_23718,N_23536,N_23594);
nand U23719 (N_23719,N_23449,N_23542);
nand U23720 (N_23720,N_23542,N_23528);
nand U23721 (N_23721,N_23572,N_23458);
nor U23722 (N_23722,N_23420,N_23480);
nor U23723 (N_23723,N_23418,N_23446);
nor U23724 (N_23724,N_23460,N_23442);
nand U23725 (N_23725,N_23540,N_23477);
and U23726 (N_23726,N_23509,N_23553);
nand U23727 (N_23727,N_23521,N_23536);
and U23728 (N_23728,N_23572,N_23510);
or U23729 (N_23729,N_23412,N_23517);
nand U23730 (N_23730,N_23531,N_23592);
and U23731 (N_23731,N_23511,N_23596);
and U23732 (N_23732,N_23497,N_23436);
nand U23733 (N_23733,N_23400,N_23549);
nand U23734 (N_23734,N_23401,N_23483);
and U23735 (N_23735,N_23461,N_23434);
nand U23736 (N_23736,N_23501,N_23447);
or U23737 (N_23737,N_23492,N_23565);
nor U23738 (N_23738,N_23434,N_23458);
nand U23739 (N_23739,N_23557,N_23485);
nand U23740 (N_23740,N_23447,N_23480);
or U23741 (N_23741,N_23592,N_23438);
nor U23742 (N_23742,N_23568,N_23442);
and U23743 (N_23743,N_23595,N_23468);
or U23744 (N_23744,N_23511,N_23457);
or U23745 (N_23745,N_23555,N_23500);
nor U23746 (N_23746,N_23430,N_23497);
or U23747 (N_23747,N_23527,N_23585);
nor U23748 (N_23748,N_23569,N_23466);
nor U23749 (N_23749,N_23504,N_23570);
nor U23750 (N_23750,N_23546,N_23495);
xor U23751 (N_23751,N_23497,N_23478);
or U23752 (N_23752,N_23527,N_23517);
nor U23753 (N_23753,N_23446,N_23429);
and U23754 (N_23754,N_23561,N_23493);
or U23755 (N_23755,N_23596,N_23525);
or U23756 (N_23756,N_23549,N_23436);
and U23757 (N_23757,N_23525,N_23452);
or U23758 (N_23758,N_23495,N_23432);
or U23759 (N_23759,N_23501,N_23438);
xor U23760 (N_23760,N_23516,N_23462);
xnor U23761 (N_23761,N_23436,N_23523);
and U23762 (N_23762,N_23519,N_23489);
nor U23763 (N_23763,N_23571,N_23411);
and U23764 (N_23764,N_23557,N_23424);
nor U23765 (N_23765,N_23470,N_23506);
xor U23766 (N_23766,N_23460,N_23415);
nand U23767 (N_23767,N_23546,N_23407);
xnor U23768 (N_23768,N_23412,N_23509);
nor U23769 (N_23769,N_23574,N_23433);
and U23770 (N_23770,N_23581,N_23573);
or U23771 (N_23771,N_23442,N_23412);
and U23772 (N_23772,N_23405,N_23422);
nor U23773 (N_23773,N_23455,N_23446);
or U23774 (N_23774,N_23540,N_23484);
or U23775 (N_23775,N_23516,N_23556);
and U23776 (N_23776,N_23483,N_23525);
and U23777 (N_23777,N_23424,N_23442);
xnor U23778 (N_23778,N_23520,N_23462);
nand U23779 (N_23779,N_23483,N_23436);
xor U23780 (N_23780,N_23542,N_23531);
and U23781 (N_23781,N_23448,N_23435);
nand U23782 (N_23782,N_23476,N_23505);
nand U23783 (N_23783,N_23412,N_23439);
or U23784 (N_23784,N_23546,N_23470);
nand U23785 (N_23785,N_23586,N_23415);
xor U23786 (N_23786,N_23401,N_23410);
xor U23787 (N_23787,N_23423,N_23473);
or U23788 (N_23788,N_23592,N_23581);
or U23789 (N_23789,N_23429,N_23510);
nor U23790 (N_23790,N_23593,N_23538);
or U23791 (N_23791,N_23473,N_23515);
nand U23792 (N_23792,N_23464,N_23578);
and U23793 (N_23793,N_23575,N_23515);
and U23794 (N_23794,N_23438,N_23528);
nor U23795 (N_23795,N_23560,N_23421);
or U23796 (N_23796,N_23530,N_23435);
xor U23797 (N_23797,N_23484,N_23470);
and U23798 (N_23798,N_23577,N_23449);
or U23799 (N_23799,N_23474,N_23549);
and U23800 (N_23800,N_23776,N_23649);
nand U23801 (N_23801,N_23770,N_23623);
or U23802 (N_23802,N_23733,N_23793);
or U23803 (N_23803,N_23774,N_23771);
and U23804 (N_23804,N_23641,N_23792);
or U23805 (N_23805,N_23690,N_23681);
nor U23806 (N_23806,N_23678,N_23672);
and U23807 (N_23807,N_23606,N_23757);
and U23808 (N_23808,N_23720,N_23766);
and U23809 (N_23809,N_23790,N_23759);
or U23810 (N_23810,N_23615,N_23740);
nor U23811 (N_23811,N_23682,N_23713);
or U23812 (N_23812,N_23786,N_23657);
nor U23813 (N_23813,N_23632,N_23687);
or U23814 (N_23814,N_23617,N_23791);
nand U23815 (N_23815,N_23778,N_23727);
nor U23816 (N_23816,N_23658,N_23679);
nand U23817 (N_23817,N_23630,N_23666);
nor U23818 (N_23818,N_23698,N_23646);
nor U23819 (N_23819,N_23633,N_23635);
nor U23820 (N_23820,N_23762,N_23744);
xor U23821 (N_23821,N_23779,N_23622);
xnor U23822 (N_23822,N_23789,N_23609);
xor U23823 (N_23823,N_23607,N_23650);
and U23824 (N_23824,N_23670,N_23704);
nand U23825 (N_23825,N_23674,N_23627);
or U23826 (N_23826,N_23725,N_23710);
xnor U23827 (N_23827,N_23602,N_23706);
nand U23828 (N_23828,N_23680,N_23783);
nor U23829 (N_23829,N_23692,N_23624);
and U23830 (N_23830,N_23717,N_23645);
nor U23831 (N_23831,N_23689,N_23749);
xor U23832 (N_23832,N_23742,N_23655);
xnor U23833 (N_23833,N_23712,N_23750);
nor U23834 (N_23834,N_23636,N_23688);
and U23835 (N_23835,N_23696,N_23787);
nor U23836 (N_23836,N_23685,N_23644);
nand U23837 (N_23837,N_23619,N_23651);
or U23838 (N_23838,N_23716,N_23686);
and U23839 (N_23839,N_23643,N_23795);
xnor U23840 (N_23840,N_23732,N_23735);
and U23841 (N_23841,N_23694,N_23768);
or U23842 (N_23842,N_23748,N_23601);
xnor U23843 (N_23843,N_23752,N_23751);
or U23844 (N_23844,N_23711,N_23603);
nand U23845 (N_23845,N_23660,N_23610);
nand U23846 (N_23846,N_23736,N_23763);
and U23847 (N_23847,N_23604,N_23767);
or U23848 (N_23848,N_23618,N_23724);
nor U23849 (N_23849,N_23760,N_23707);
and U23850 (N_23850,N_23664,N_23671);
xnor U23851 (N_23851,N_23621,N_23605);
and U23852 (N_23852,N_23616,N_23675);
or U23853 (N_23853,N_23753,N_23709);
and U23854 (N_23854,N_23654,N_23715);
or U23855 (N_23855,N_23699,N_23611);
or U23856 (N_23856,N_23745,N_23705);
nor U23857 (N_23857,N_23628,N_23673);
and U23858 (N_23858,N_23656,N_23661);
nand U23859 (N_23859,N_23648,N_23684);
xnor U23860 (N_23860,N_23798,N_23775);
or U23861 (N_23861,N_23691,N_23640);
and U23862 (N_23862,N_23755,N_23631);
and U23863 (N_23863,N_23703,N_23620);
nand U23864 (N_23864,N_23788,N_23773);
and U23865 (N_23865,N_23659,N_23634);
nor U23866 (N_23866,N_23739,N_23746);
nand U23867 (N_23867,N_23697,N_23719);
nor U23868 (N_23868,N_23723,N_23730);
nor U23869 (N_23869,N_23747,N_23608);
nor U23870 (N_23870,N_23731,N_23663);
xnor U23871 (N_23871,N_23662,N_23754);
nand U23872 (N_23872,N_23613,N_23782);
xnor U23873 (N_23873,N_23769,N_23764);
and U23874 (N_23874,N_23718,N_23668);
nor U23875 (N_23875,N_23781,N_23642);
nand U23876 (N_23876,N_23738,N_23677);
nor U23877 (N_23877,N_23784,N_23772);
nand U23878 (N_23878,N_23612,N_23729);
nand U23879 (N_23879,N_23737,N_23734);
nor U23880 (N_23880,N_23637,N_23695);
nor U23881 (N_23881,N_23614,N_23667);
nor U23882 (N_23882,N_23625,N_23653);
nand U23883 (N_23883,N_23701,N_23665);
nor U23884 (N_23884,N_23765,N_23777);
and U23885 (N_23885,N_23722,N_23756);
xor U23886 (N_23886,N_23708,N_23600);
nor U23887 (N_23887,N_23626,N_23714);
and U23888 (N_23888,N_23639,N_23702);
xor U23889 (N_23889,N_23700,N_23758);
and U23890 (N_23890,N_23652,N_23728);
xnor U23891 (N_23891,N_23721,N_23638);
and U23892 (N_23892,N_23799,N_23683);
and U23893 (N_23893,N_23785,N_23796);
xnor U23894 (N_23894,N_23629,N_23726);
and U23895 (N_23895,N_23647,N_23797);
nand U23896 (N_23896,N_23743,N_23761);
and U23897 (N_23897,N_23676,N_23780);
xnor U23898 (N_23898,N_23693,N_23741);
and U23899 (N_23899,N_23794,N_23669);
and U23900 (N_23900,N_23754,N_23705);
xnor U23901 (N_23901,N_23677,N_23627);
nand U23902 (N_23902,N_23777,N_23742);
nor U23903 (N_23903,N_23795,N_23740);
or U23904 (N_23904,N_23747,N_23633);
and U23905 (N_23905,N_23661,N_23642);
xor U23906 (N_23906,N_23704,N_23685);
and U23907 (N_23907,N_23657,N_23785);
nor U23908 (N_23908,N_23717,N_23785);
and U23909 (N_23909,N_23648,N_23770);
nand U23910 (N_23910,N_23648,N_23643);
and U23911 (N_23911,N_23695,N_23791);
nor U23912 (N_23912,N_23721,N_23689);
nor U23913 (N_23913,N_23691,N_23628);
xnor U23914 (N_23914,N_23751,N_23622);
or U23915 (N_23915,N_23761,N_23712);
or U23916 (N_23916,N_23645,N_23736);
or U23917 (N_23917,N_23620,N_23727);
nand U23918 (N_23918,N_23799,N_23626);
xor U23919 (N_23919,N_23747,N_23666);
and U23920 (N_23920,N_23716,N_23712);
and U23921 (N_23921,N_23765,N_23731);
nor U23922 (N_23922,N_23675,N_23613);
or U23923 (N_23923,N_23762,N_23702);
nor U23924 (N_23924,N_23624,N_23757);
or U23925 (N_23925,N_23791,N_23769);
and U23926 (N_23926,N_23685,N_23792);
xor U23927 (N_23927,N_23642,N_23613);
nor U23928 (N_23928,N_23651,N_23615);
xnor U23929 (N_23929,N_23714,N_23696);
nor U23930 (N_23930,N_23733,N_23650);
nand U23931 (N_23931,N_23719,N_23644);
xor U23932 (N_23932,N_23677,N_23761);
nand U23933 (N_23933,N_23690,N_23710);
nor U23934 (N_23934,N_23661,N_23776);
and U23935 (N_23935,N_23794,N_23607);
nand U23936 (N_23936,N_23753,N_23685);
nor U23937 (N_23937,N_23688,N_23798);
nand U23938 (N_23938,N_23718,N_23769);
or U23939 (N_23939,N_23675,N_23628);
nor U23940 (N_23940,N_23784,N_23779);
or U23941 (N_23941,N_23742,N_23729);
or U23942 (N_23942,N_23733,N_23736);
or U23943 (N_23943,N_23641,N_23715);
nand U23944 (N_23944,N_23780,N_23693);
or U23945 (N_23945,N_23672,N_23752);
xor U23946 (N_23946,N_23753,N_23667);
nor U23947 (N_23947,N_23627,N_23602);
or U23948 (N_23948,N_23729,N_23763);
or U23949 (N_23949,N_23685,N_23658);
xor U23950 (N_23950,N_23690,N_23615);
nand U23951 (N_23951,N_23608,N_23630);
or U23952 (N_23952,N_23788,N_23706);
nand U23953 (N_23953,N_23617,N_23604);
or U23954 (N_23954,N_23654,N_23686);
xnor U23955 (N_23955,N_23613,N_23617);
and U23956 (N_23956,N_23674,N_23763);
xor U23957 (N_23957,N_23777,N_23685);
and U23958 (N_23958,N_23641,N_23791);
and U23959 (N_23959,N_23641,N_23666);
and U23960 (N_23960,N_23794,N_23614);
nor U23961 (N_23961,N_23698,N_23629);
nor U23962 (N_23962,N_23778,N_23783);
xor U23963 (N_23963,N_23611,N_23798);
or U23964 (N_23964,N_23738,N_23680);
nand U23965 (N_23965,N_23655,N_23620);
nand U23966 (N_23966,N_23690,N_23652);
xnor U23967 (N_23967,N_23621,N_23793);
or U23968 (N_23968,N_23622,N_23770);
nand U23969 (N_23969,N_23702,N_23657);
xor U23970 (N_23970,N_23758,N_23792);
nand U23971 (N_23971,N_23619,N_23738);
and U23972 (N_23972,N_23701,N_23789);
nand U23973 (N_23973,N_23607,N_23768);
or U23974 (N_23974,N_23737,N_23713);
and U23975 (N_23975,N_23646,N_23623);
and U23976 (N_23976,N_23608,N_23685);
xnor U23977 (N_23977,N_23668,N_23679);
or U23978 (N_23978,N_23767,N_23605);
or U23979 (N_23979,N_23724,N_23732);
nand U23980 (N_23980,N_23793,N_23633);
or U23981 (N_23981,N_23711,N_23763);
or U23982 (N_23982,N_23785,N_23679);
or U23983 (N_23983,N_23751,N_23760);
nor U23984 (N_23984,N_23687,N_23681);
and U23985 (N_23985,N_23780,N_23644);
and U23986 (N_23986,N_23731,N_23653);
and U23987 (N_23987,N_23690,N_23772);
or U23988 (N_23988,N_23744,N_23799);
xnor U23989 (N_23989,N_23630,N_23753);
nor U23990 (N_23990,N_23766,N_23749);
xnor U23991 (N_23991,N_23742,N_23735);
or U23992 (N_23992,N_23652,N_23780);
nor U23993 (N_23993,N_23630,N_23794);
or U23994 (N_23994,N_23625,N_23628);
nand U23995 (N_23995,N_23712,N_23770);
or U23996 (N_23996,N_23683,N_23706);
nor U23997 (N_23997,N_23684,N_23675);
or U23998 (N_23998,N_23795,N_23779);
nand U23999 (N_23999,N_23738,N_23766);
nor U24000 (N_24000,N_23919,N_23960);
and U24001 (N_24001,N_23954,N_23903);
nand U24002 (N_24002,N_23859,N_23988);
or U24003 (N_24003,N_23856,N_23887);
and U24004 (N_24004,N_23907,N_23935);
or U24005 (N_24005,N_23983,N_23932);
xnor U24006 (N_24006,N_23839,N_23912);
or U24007 (N_24007,N_23888,N_23953);
or U24008 (N_24008,N_23924,N_23882);
nand U24009 (N_24009,N_23963,N_23858);
nand U24010 (N_24010,N_23985,N_23969);
or U24011 (N_24011,N_23914,N_23834);
or U24012 (N_24012,N_23951,N_23822);
or U24013 (N_24013,N_23892,N_23964);
or U24014 (N_24014,N_23898,N_23832);
and U24015 (N_24015,N_23923,N_23974);
nor U24016 (N_24016,N_23994,N_23833);
nor U24017 (N_24017,N_23827,N_23818);
xnor U24018 (N_24018,N_23941,N_23978);
and U24019 (N_24019,N_23893,N_23883);
xnor U24020 (N_24020,N_23920,N_23873);
nand U24021 (N_24021,N_23991,N_23910);
nand U24022 (N_24022,N_23906,N_23940);
nand U24023 (N_24023,N_23956,N_23909);
xnor U24024 (N_24024,N_23992,N_23885);
and U24025 (N_24025,N_23804,N_23810);
xnor U24026 (N_24026,N_23879,N_23880);
and U24027 (N_24027,N_23824,N_23821);
and U24028 (N_24028,N_23871,N_23847);
xnor U24029 (N_24029,N_23830,N_23840);
and U24030 (N_24030,N_23896,N_23801);
xnor U24031 (N_24031,N_23814,N_23816);
nand U24032 (N_24032,N_23876,N_23846);
xor U24033 (N_24033,N_23891,N_23843);
xnor U24034 (N_24034,N_23952,N_23889);
nand U24035 (N_24035,N_23812,N_23976);
and U24036 (N_24036,N_23990,N_23865);
nor U24037 (N_24037,N_23872,N_23894);
nand U24038 (N_24038,N_23828,N_23823);
or U24039 (N_24039,N_23886,N_23845);
xor U24040 (N_24040,N_23900,N_23805);
or U24041 (N_24041,N_23970,N_23848);
or U24042 (N_24042,N_23874,N_23977);
nand U24043 (N_24043,N_23949,N_23857);
xor U24044 (N_24044,N_23967,N_23980);
xnor U24045 (N_24045,N_23947,N_23817);
xnor U24046 (N_24046,N_23875,N_23844);
nor U24047 (N_24047,N_23945,N_23837);
nor U24048 (N_24048,N_23901,N_23939);
nand U24049 (N_24049,N_23926,N_23841);
nand U24050 (N_24050,N_23809,N_23958);
or U24051 (N_24051,N_23806,N_23937);
nor U24052 (N_24052,N_23820,N_23884);
or U24053 (N_24053,N_23895,N_23938);
xnor U24054 (N_24054,N_23966,N_23917);
nand U24055 (N_24055,N_23850,N_23968);
or U24056 (N_24056,N_23902,N_23890);
nor U24057 (N_24057,N_23864,N_23852);
and U24058 (N_24058,N_23930,N_23997);
xnor U24059 (N_24059,N_23943,N_23867);
and U24060 (N_24060,N_23948,N_23959);
and U24061 (N_24061,N_23961,N_23842);
or U24062 (N_24062,N_23829,N_23979);
or U24063 (N_24063,N_23811,N_23870);
and U24064 (N_24064,N_23929,N_23904);
nand U24065 (N_24065,N_23807,N_23957);
or U24066 (N_24066,N_23933,N_23922);
xor U24067 (N_24067,N_23862,N_23971);
xnor U24068 (N_24068,N_23911,N_23854);
nand U24069 (N_24069,N_23955,N_23921);
nor U24070 (N_24070,N_23936,N_23908);
xnor U24071 (N_24071,N_23881,N_23808);
or U24072 (N_24072,N_23946,N_23981);
xnor U24073 (N_24073,N_23982,N_23836);
nor U24074 (N_24074,N_23927,N_23826);
and U24075 (N_24075,N_23851,N_23989);
xor U24076 (N_24076,N_23972,N_23877);
nor U24077 (N_24077,N_23819,N_23897);
nand U24078 (N_24078,N_23913,N_23878);
and U24079 (N_24079,N_23998,N_23993);
xor U24080 (N_24080,N_23916,N_23986);
nand U24081 (N_24081,N_23831,N_23855);
or U24082 (N_24082,N_23868,N_23995);
xnor U24083 (N_24083,N_23863,N_23866);
and U24084 (N_24084,N_23802,N_23944);
or U24085 (N_24085,N_23962,N_23861);
nor U24086 (N_24086,N_23987,N_23925);
nor U24087 (N_24087,N_23800,N_23915);
nand U24088 (N_24088,N_23905,N_23853);
xnor U24089 (N_24089,N_23996,N_23835);
xnor U24090 (N_24090,N_23803,N_23973);
nand U24091 (N_24091,N_23899,N_23950);
and U24092 (N_24092,N_23984,N_23942);
xnor U24093 (N_24093,N_23965,N_23825);
nand U24094 (N_24094,N_23815,N_23999);
nor U24095 (N_24095,N_23934,N_23838);
or U24096 (N_24096,N_23813,N_23928);
or U24097 (N_24097,N_23931,N_23860);
nor U24098 (N_24098,N_23918,N_23869);
nand U24099 (N_24099,N_23849,N_23975);
nor U24100 (N_24100,N_23863,N_23887);
nor U24101 (N_24101,N_23953,N_23885);
xnor U24102 (N_24102,N_23819,N_23983);
or U24103 (N_24103,N_23961,N_23936);
xor U24104 (N_24104,N_23857,N_23838);
nor U24105 (N_24105,N_23882,N_23940);
xor U24106 (N_24106,N_23865,N_23881);
nor U24107 (N_24107,N_23841,N_23868);
nor U24108 (N_24108,N_23969,N_23943);
nand U24109 (N_24109,N_23872,N_23951);
and U24110 (N_24110,N_23899,N_23847);
xnor U24111 (N_24111,N_23837,N_23961);
and U24112 (N_24112,N_23903,N_23843);
and U24113 (N_24113,N_23961,N_23849);
and U24114 (N_24114,N_23975,N_23811);
or U24115 (N_24115,N_23851,N_23932);
xor U24116 (N_24116,N_23949,N_23921);
nor U24117 (N_24117,N_23961,N_23861);
nor U24118 (N_24118,N_23925,N_23945);
nand U24119 (N_24119,N_23829,N_23824);
nor U24120 (N_24120,N_23937,N_23849);
or U24121 (N_24121,N_23932,N_23988);
xor U24122 (N_24122,N_23902,N_23965);
nand U24123 (N_24123,N_23806,N_23940);
nor U24124 (N_24124,N_23803,N_23971);
xnor U24125 (N_24125,N_23896,N_23871);
and U24126 (N_24126,N_23997,N_23848);
and U24127 (N_24127,N_23837,N_23871);
nand U24128 (N_24128,N_23891,N_23945);
and U24129 (N_24129,N_23838,N_23851);
xnor U24130 (N_24130,N_23970,N_23826);
or U24131 (N_24131,N_23835,N_23914);
xnor U24132 (N_24132,N_23977,N_23800);
or U24133 (N_24133,N_23967,N_23860);
nor U24134 (N_24134,N_23846,N_23959);
and U24135 (N_24135,N_23909,N_23930);
nand U24136 (N_24136,N_23824,N_23859);
xor U24137 (N_24137,N_23944,N_23966);
nand U24138 (N_24138,N_23988,N_23832);
nand U24139 (N_24139,N_23813,N_23936);
nand U24140 (N_24140,N_23928,N_23824);
nand U24141 (N_24141,N_23867,N_23864);
or U24142 (N_24142,N_23953,N_23997);
and U24143 (N_24143,N_23984,N_23938);
and U24144 (N_24144,N_23926,N_23927);
and U24145 (N_24145,N_23920,N_23901);
and U24146 (N_24146,N_23851,N_23976);
xor U24147 (N_24147,N_23802,N_23874);
or U24148 (N_24148,N_23936,N_23833);
and U24149 (N_24149,N_23875,N_23987);
xor U24150 (N_24150,N_23880,N_23897);
and U24151 (N_24151,N_23895,N_23908);
xnor U24152 (N_24152,N_23972,N_23802);
or U24153 (N_24153,N_23946,N_23945);
and U24154 (N_24154,N_23951,N_23823);
nor U24155 (N_24155,N_23803,N_23862);
nand U24156 (N_24156,N_23836,N_23881);
or U24157 (N_24157,N_23955,N_23954);
and U24158 (N_24158,N_23910,N_23891);
and U24159 (N_24159,N_23844,N_23941);
and U24160 (N_24160,N_23812,N_23949);
and U24161 (N_24161,N_23842,N_23963);
and U24162 (N_24162,N_23860,N_23841);
nor U24163 (N_24163,N_23927,N_23942);
nand U24164 (N_24164,N_23943,N_23981);
nor U24165 (N_24165,N_23973,N_23831);
nand U24166 (N_24166,N_23850,N_23865);
nand U24167 (N_24167,N_23889,N_23809);
nand U24168 (N_24168,N_23983,N_23973);
and U24169 (N_24169,N_23848,N_23892);
and U24170 (N_24170,N_23887,N_23922);
nor U24171 (N_24171,N_23816,N_23847);
and U24172 (N_24172,N_23851,N_23954);
nor U24173 (N_24173,N_23859,N_23930);
or U24174 (N_24174,N_23961,N_23938);
nor U24175 (N_24175,N_23836,N_23888);
and U24176 (N_24176,N_23891,N_23801);
or U24177 (N_24177,N_23971,N_23860);
nand U24178 (N_24178,N_23979,N_23807);
and U24179 (N_24179,N_23960,N_23949);
or U24180 (N_24180,N_23852,N_23876);
or U24181 (N_24181,N_23986,N_23930);
and U24182 (N_24182,N_23879,N_23944);
or U24183 (N_24183,N_23993,N_23820);
and U24184 (N_24184,N_23936,N_23883);
or U24185 (N_24185,N_23891,N_23823);
nor U24186 (N_24186,N_23984,N_23897);
nand U24187 (N_24187,N_23906,N_23945);
nor U24188 (N_24188,N_23855,N_23858);
xnor U24189 (N_24189,N_23822,N_23825);
xnor U24190 (N_24190,N_23837,N_23807);
xor U24191 (N_24191,N_23856,N_23985);
nand U24192 (N_24192,N_23818,N_23980);
xnor U24193 (N_24193,N_23878,N_23856);
and U24194 (N_24194,N_23851,N_23813);
nor U24195 (N_24195,N_23914,N_23877);
xnor U24196 (N_24196,N_23941,N_23801);
nor U24197 (N_24197,N_23980,N_23986);
xor U24198 (N_24198,N_23903,N_23928);
or U24199 (N_24199,N_23835,N_23821);
xnor U24200 (N_24200,N_24186,N_24100);
xnor U24201 (N_24201,N_24187,N_24001);
xor U24202 (N_24202,N_24134,N_24080);
nor U24203 (N_24203,N_24078,N_24168);
nand U24204 (N_24204,N_24184,N_24103);
or U24205 (N_24205,N_24013,N_24069);
or U24206 (N_24206,N_24153,N_24198);
and U24207 (N_24207,N_24163,N_24067);
nand U24208 (N_24208,N_24195,N_24169);
nand U24209 (N_24209,N_24162,N_24004);
nor U24210 (N_24210,N_24130,N_24082);
or U24211 (N_24211,N_24054,N_24086);
and U24212 (N_24212,N_24056,N_24097);
xnor U24213 (N_24213,N_24114,N_24115);
xor U24214 (N_24214,N_24116,N_24154);
or U24215 (N_24215,N_24000,N_24112);
or U24216 (N_24216,N_24071,N_24111);
xnor U24217 (N_24217,N_24131,N_24096);
nand U24218 (N_24218,N_24042,N_24045);
and U24219 (N_24219,N_24025,N_24102);
xnor U24220 (N_24220,N_24147,N_24174);
and U24221 (N_24221,N_24012,N_24185);
and U24222 (N_24222,N_24008,N_24015);
or U24223 (N_24223,N_24070,N_24002);
and U24224 (N_24224,N_24181,N_24117);
xnor U24225 (N_24225,N_24140,N_24019);
nand U24226 (N_24226,N_24156,N_24160);
and U24227 (N_24227,N_24196,N_24120);
or U24228 (N_24228,N_24017,N_24074);
nand U24229 (N_24229,N_24094,N_24060);
xor U24230 (N_24230,N_24139,N_24027);
and U24231 (N_24231,N_24129,N_24044);
nand U24232 (N_24232,N_24031,N_24164);
and U24233 (N_24233,N_24090,N_24172);
or U24234 (N_24234,N_24142,N_24107);
nand U24235 (N_24235,N_24053,N_24165);
nor U24236 (N_24236,N_24144,N_24030);
or U24237 (N_24237,N_24149,N_24037);
and U24238 (N_24238,N_24141,N_24136);
or U24239 (N_24239,N_24146,N_24190);
or U24240 (N_24240,N_24182,N_24143);
nand U24241 (N_24241,N_24076,N_24121);
and U24242 (N_24242,N_24068,N_24061);
or U24243 (N_24243,N_24123,N_24039);
nand U24244 (N_24244,N_24137,N_24119);
xor U24245 (N_24245,N_24124,N_24183);
nand U24246 (N_24246,N_24050,N_24064);
nor U24247 (N_24247,N_24040,N_24171);
and U24248 (N_24248,N_24036,N_24145);
or U24249 (N_24249,N_24167,N_24072);
nand U24250 (N_24250,N_24125,N_24148);
nand U24251 (N_24251,N_24091,N_24105);
or U24252 (N_24252,N_24043,N_24109);
nand U24253 (N_24253,N_24110,N_24035);
nand U24254 (N_24254,N_24084,N_24155);
nor U24255 (N_24255,N_24159,N_24092);
and U24256 (N_24256,N_24178,N_24151);
nand U24257 (N_24257,N_24118,N_24028);
xor U24258 (N_24258,N_24089,N_24099);
nor U24259 (N_24259,N_24133,N_24087);
nand U24260 (N_24260,N_24170,N_24095);
xor U24261 (N_24261,N_24192,N_24108);
or U24262 (N_24262,N_24128,N_24180);
and U24263 (N_24263,N_24075,N_24065);
and U24264 (N_24264,N_24132,N_24157);
and U24265 (N_24265,N_24009,N_24166);
nor U24266 (N_24266,N_24049,N_24066);
and U24267 (N_24267,N_24003,N_24010);
nor U24268 (N_24268,N_24122,N_24047);
or U24269 (N_24269,N_24024,N_24011);
xor U24270 (N_24270,N_24194,N_24150);
or U24271 (N_24271,N_24063,N_24197);
or U24272 (N_24272,N_24026,N_24177);
or U24273 (N_24273,N_24046,N_24051);
xor U24274 (N_24274,N_24199,N_24113);
and U24275 (N_24275,N_24158,N_24032);
or U24276 (N_24276,N_24189,N_24104);
nand U24277 (N_24277,N_24055,N_24152);
xor U24278 (N_24278,N_24022,N_24138);
nor U24279 (N_24279,N_24034,N_24057);
xnor U24280 (N_24280,N_24081,N_24088);
and U24281 (N_24281,N_24073,N_24191);
nor U24282 (N_24282,N_24052,N_24127);
nand U24283 (N_24283,N_24041,N_24077);
and U24284 (N_24284,N_24006,N_24173);
or U24285 (N_24285,N_24188,N_24014);
and U24286 (N_24286,N_24029,N_24085);
nor U24287 (N_24287,N_24038,N_24023);
or U24288 (N_24288,N_24193,N_24126);
xor U24289 (N_24289,N_24016,N_24062);
and U24290 (N_24290,N_24005,N_24020);
xnor U24291 (N_24291,N_24135,N_24021);
nand U24292 (N_24292,N_24018,N_24048);
nor U24293 (N_24293,N_24083,N_24098);
nor U24294 (N_24294,N_24101,N_24175);
and U24295 (N_24295,N_24058,N_24161);
nor U24296 (N_24296,N_24033,N_24007);
nand U24297 (N_24297,N_24176,N_24106);
or U24298 (N_24298,N_24079,N_24179);
nor U24299 (N_24299,N_24059,N_24093);
xnor U24300 (N_24300,N_24033,N_24074);
xnor U24301 (N_24301,N_24006,N_24151);
nor U24302 (N_24302,N_24142,N_24007);
nor U24303 (N_24303,N_24027,N_24009);
nand U24304 (N_24304,N_24192,N_24194);
or U24305 (N_24305,N_24003,N_24034);
or U24306 (N_24306,N_24053,N_24164);
nor U24307 (N_24307,N_24116,N_24012);
xor U24308 (N_24308,N_24097,N_24158);
xor U24309 (N_24309,N_24014,N_24062);
xor U24310 (N_24310,N_24179,N_24198);
and U24311 (N_24311,N_24195,N_24140);
nand U24312 (N_24312,N_24149,N_24130);
xor U24313 (N_24313,N_24020,N_24006);
nand U24314 (N_24314,N_24066,N_24086);
and U24315 (N_24315,N_24123,N_24163);
nand U24316 (N_24316,N_24181,N_24068);
nand U24317 (N_24317,N_24113,N_24170);
nand U24318 (N_24318,N_24049,N_24062);
and U24319 (N_24319,N_24108,N_24142);
or U24320 (N_24320,N_24051,N_24048);
nor U24321 (N_24321,N_24080,N_24191);
or U24322 (N_24322,N_24003,N_24113);
nand U24323 (N_24323,N_24088,N_24107);
nor U24324 (N_24324,N_24186,N_24154);
nand U24325 (N_24325,N_24105,N_24085);
xnor U24326 (N_24326,N_24007,N_24165);
nor U24327 (N_24327,N_24093,N_24138);
nand U24328 (N_24328,N_24178,N_24197);
nor U24329 (N_24329,N_24112,N_24100);
nor U24330 (N_24330,N_24016,N_24193);
nor U24331 (N_24331,N_24033,N_24047);
or U24332 (N_24332,N_24059,N_24032);
xor U24333 (N_24333,N_24001,N_24015);
nor U24334 (N_24334,N_24053,N_24134);
nand U24335 (N_24335,N_24034,N_24146);
nand U24336 (N_24336,N_24160,N_24018);
or U24337 (N_24337,N_24049,N_24073);
xor U24338 (N_24338,N_24022,N_24098);
nand U24339 (N_24339,N_24163,N_24003);
or U24340 (N_24340,N_24139,N_24047);
xor U24341 (N_24341,N_24098,N_24168);
xor U24342 (N_24342,N_24162,N_24120);
xnor U24343 (N_24343,N_24162,N_24035);
or U24344 (N_24344,N_24053,N_24152);
nand U24345 (N_24345,N_24102,N_24026);
nand U24346 (N_24346,N_24044,N_24075);
and U24347 (N_24347,N_24086,N_24159);
or U24348 (N_24348,N_24098,N_24052);
xnor U24349 (N_24349,N_24053,N_24106);
xnor U24350 (N_24350,N_24186,N_24129);
nand U24351 (N_24351,N_24189,N_24134);
or U24352 (N_24352,N_24158,N_24154);
or U24353 (N_24353,N_24028,N_24023);
xnor U24354 (N_24354,N_24009,N_24033);
nand U24355 (N_24355,N_24142,N_24133);
nand U24356 (N_24356,N_24157,N_24148);
nand U24357 (N_24357,N_24187,N_24006);
or U24358 (N_24358,N_24007,N_24015);
or U24359 (N_24359,N_24064,N_24088);
or U24360 (N_24360,N_24098,N_24199);
nand U24361 (N_24361,N_24092,N_24070);
and U24362 (N_24362,N_24177,N_24055);
nand U24363 (N_24363,N_24173,N_24078);
or U24364 (N_24364,N_24179,N_24016);
nor U24365 (N_24365,N_24109,N_24189);
nand U24366 (N_24366,N_24181,N_24133);
nor U24367 (N_24367,N_24055,N_24004);
or U24368 (N_24368,N_24076,N_24036);
xor U24369 (N_24369,N_24013,N_24154);
xor U24370 (N_24370,N_24049,N_24172);
or U24371 (N_24371,N_24040,N_24084);
or U24372 (N_24372,N_24099,N_24171);
xor U24373 (N_24373,N_24170,N_24033);
xor U24374 (N_24374,N_24177,N_24136);
or U24375 (N_24375,N_24136,N_24083);
and U24376 (N_24376,N_24154,N_24163);
xnor U24377 (N_24377,N_24031,N_24145);
or U24378 (N_24378,N_24002,N_24047);
or U24379 (N_24379,N_24175,N_24070);
nand U24380 (N_24380,N_24168,N_24089);
and U24381 (N_24381,N_24028,N_24006);
and U24382 (N_24382,N_24119,N_24028);
or U24383 (N_24383,N_24007,N_24062);
or U24384 (N_24384,N_24098,N_24047);
nand U24385 (N_24385,N_24194,N_24103);
xnor U24386 (N_24386,N_24101,N_24025);
nand U24387 (N_24387,N_24050,N_24125);
or U24388 (N_24388,N_24094,N_24004);
xor U24389 (N_24389,N_24109,N_24111);
and U24390 (N_24390,N_24024,N_24186);
or U24391 (N_24391,N_24080,N_24009);
nand U24392 (N_24392,N_24139,N_24024);
or U24393 (N_24393,N_24107,N_24105);
and U24394 (N_24394,N_24091,N_24051);
xnor U24395 (N_24395,N_24135,N_24075);
or U24396 (N_24396,N_24183,N_24193);
nor U24397 (N_24397,N_24073,N_24167);
nand U24398 (N_24398,N_24043,N_24144);
nor U24399 (N_24399,N_24067,N_24174);
xnor U24400 (N_24400,N_24306,N_24331);
nand U24401 (N_24401,N_24329,N_24305);
xor U24402 (N_24402,N_24393,N_24320);
or U24403 (N_24403,N_24253,N_24359);
nor U24404 (N_24404,N_24262,N_24390);
nand U24405 (N_24405,N_24325,N_24371);
xnor U24406 (N_24406,N_24268,N_24345);
or U24407 (N_24407,N_24279,N_24340);
or U24408 (N_24408,N_24266,N_24288);
and U24409 (N_24409,N_24332,N_24337);
or U24410 (N_24410,N_24386,N_24227);
xor U24411 (N_24411,N_24293,N_24310);
nand U24412 (N_24412,N_24213,N_24252);
nor U24413 (N_24413,N_24231,N_24214);
and U24414 (N_24414,N_24243,N_24284);
nor U24415 (N_24415,N_24235,N_24241);
xor U24416 (N_24416,N_24287,N_24240);
and U24417 (N_24417,N_24391,N_24220);
nand U24418 (N_24418,N_24274,N_24398);
nand U24419 (N_24419,N_24375,N_24315);
nand U24420 (N_24420,N_24299,N_24285);
nand U24421 (N_24421,N_24369,N_24229);
nor U24422 (N_24422,N_24210,N_24349);
nor U24423 (N_24423,N_24387,N_24316);
nor U24424 (N_24424,N_24322,N_24270);
xor U24425 (N_24425,N_24264,N_24234);
and U24426 (N_24426,N_24254,N_24341);
or U24427 (N_24427,N_24292,N_24383);
and U24428 (N_24428,N_24200,N_24309);
xor U24429 (N_24429,N_24244,N_24392);
and U24430 (N_24430,N_24267,N_24312);
or U24431 (N_24431,N_24226,N_24372);
xor U24432 (N_24432,N_24248,N_24269);
or U24433 (N_24433,N_24335,N_24291);
and U24434 (N_24434,N_24265,N_24365);
xnor U24435 (N_24435,N_24208,N_24308);
nand U24436 (N_24436,N_24354,N_24295);
xnor U24437 (N_24437,N_24206,N_24237);
xnor U24438 (N_24438,N_24223,N_24294);
and U24439 (N_24439,N_24209,N_24302);
xor U24440 (N_24440,N_24389,N_24380);
nand U24441 (N_24441,N_24289,N_24319);
xor U24442 (N_24442,N_24222,N_24326);
xnor U24443 (N_24443,N_24297,N_24218);
or U24444 (N_24444,N_24352,N_24207);
or U24445 (N_24445,N_24278,N_24307);
nor U24446 (N_24446,N_24228,N_24239);
or U24447 (N_24447,N_24296,N_24358);
or U24448 (N_24448,N_24263,N_24204);
and U24449 (N_24449,N_24339,N_24355);
or U24450 (N_24450,N_24280,N_24343);
or U24451 (N_24451,N_24353,N_24216);
or U24452 (N_24452,N_24377,N_24374);
and U24453 (N_24453,N_24330,N_24211);
xnor U24454 (N_24454,N_24300,N_24271);
nor U24455 (N_24455,N_24378,N_24225);
and U24456 (N_24456,N_24394,N_24251);
nand U24457 (N_24457,N_24356,N_24348);
xor U24458 (N_24458,N_24333,N_24388);
nand U24459 (N_24459,N_24342,N_24317);
xnor U24460 (N_24460,N_24376,N_24219);
or U24461 (N_24461,N_24250,N_24367);
nor U24462 (N_24462,N_24238,N_24364);
nor U24463 (N_24463,N_24283,N_24298);
nor U24464 (N_24464,N_24236,N_24303);
nand U24465 (N_24465,N_24203,N_24314);
xnor U24466 (N_24466,N_24205,N_24382);
nor U24467 (N_24467,N_24328,N_24260);
nand U24468 (N_24468,N_24215,N_24362);
and U24469 (N_24469,N_24301,N_24272);
and U24470 (N_24470,N_24344,N_24385);
nand U24471 (N_24471,N_24217,N_24256);
xor U24472 (N_24472,N_24311,N_24336);
nor U24473 (N_24473,N_24212,N_24247);
or U24474 (N_24474,N_24224,N_24257);
xor U24475 (N_24475,N_24396,N_24276);
and U24476 (N_24476,N_24360,N_24334);
nor U24477 (N_24477,N_24259,N_24346);
nor U24478 (N_24478,N_24321,N_24232);
nor U24479 (N_24479,N_24233,N_24313);
and U24480 (N_24480,N_24273,N_24395);
nor U24481 (N_24481,N_24281,N_24338);
xor U24482 (N_24482,N_24366,N_24258);
xor U24483 (N_24483,N_24230,N_24350);
or U24484 (N_24484,N_24201,N_24323);
xor U24485 (N_24485,N_24361,N_24290);
nor U24486 (N_24486,N_24368,N_24286);
or U24487 (N_24487,N_24255,N_24202);
nand U24488 (N_24488,N_24261,N_24304);
and U24489 (N_24489,N_24277,N_24246);
and U24490 (N_24490,N_24318,N_24245);
nand U24491 (N_24491,N_24242,N_24384);
nor U24492 (N_24492,N_24347,N_24399);
and U24493 (N_24493,N_24221,N_24363);
nand U24494 (N_24494,N_24249,N_24397);
or U24495 (N_24495,N_24324,N_24381);
or U24496 (N_24496,N_24373,N_24327);
and U24497 (N_24497,N_24357,N_24351);
nor U24498 (N_24498,N_24370,N_24275);
and U24499 (N_24499,N_24379,N_24282);
or U24500 (N_24500,N_24279,N_24310);
and U24501 (N_24501,N_24333,N_24397);
nor U24502 (N_24502,N_24272,N_24353);
or U24503 (N_24503,N_24369,N_24234);
nand U24504 (N_24504,N_24349,N_24218);
xor U24505 (N_24505,N_24375,N_24397);
nand U24506 (N_24506,N_24253,N_24347);
xnor U24507 (N_24507,N_24212,N_24360);
and U24508 (N_24508,N_24348,N_24333);
nor U24509 (N_24509,N_24370,N_24391);
and U24510 (N_24510,N_24376,N_24200);
nor U24511 (N_24511,N_24341,N_24295);
or U24512 (N_24512,N_24202,N_24301);
nor U24513 (N_24513,N_24218,N_24261);
xnor U24514 (N_24514,N_24218,N_24268);
and U24515 (N_24515,N_24288,N_24286);
and U24516 (N_24516,N_24238,N_24292);
or U24517 (N_24517,N_24365,N_24379);
or U24518 (N_24518,N_24333,N_24200);
and U24519 (N_24519,N_24354,N_24222);
nand U24520 (N_24520,N_24209,N_24328);
xnor U24521 (N_24521,N_24396,N_24239);
xor U24522 (N_24522,N_24274,N_24252);
nor U24523 (N_24523,N_24391,N_24393);
nand U24524 (N_24524,N_24329,N_24351);
xor U24525 (N_24525,N_24289,N_24354);
xor U24526 (N_24526,N_24274,N_24219);
xor U24527 (N_24527,N_24270,N_24245);
or U24528 (N_24528,N_24362,N_24343);
or U24529 (N_24529,N_24303,N_24348);
and U24530 (N_24530,N_24244,N_24307);
nand U24531 (N_24531,N_24396,N_24217);
xnor U24532 (N_24532,N_24328,N_24305);
or U24533 (N_24533,N_24209,N_24260);
nand U24534 (N_24534,N_24334,N_24291);
and U24535 (N_24535,N_24304,N_24303);
and U24536 (N_24536,N_24232,N_24346);
xor U24537 (N_24537,N_24308,N_24285);
nor U24538 (N_24538,N_24209,N_24332);
and U24539 (N_24539,N_24306,N_24249);
nor U24540 (N_24540,N_24284,N_24211);
or U24541 (N_24541,N_24343,N_24318);
xor U24542 (N_24542,N_24302,N_24399);
and U24543 (N_24543,N_24326,N_24262);
nor U24544 (N_24544,N_24278,N_24398);
nor U24545 (N_24545,N_24337,N_24269);
nor U24546 (N_24546,N_24368,N_24331);
xnor U24547 (N_24547,N_24360,N_24221);
and U24548 (N_24548,N_24279,N_24233);
nand U24549 (N_24549,N_24384,N_24262);
nand U24550 (N_24550,N_24348,N_24271);
nor U24551 (N_24551,N_24313,N_24321);
nand U24552 (N_24552,N_24219,N_24213);
nand U24553 (N_24553,N_24332,N_24231);
nor U24554 (N_24554,N_24347,N_24224);
or U24555 (N_24555,N_24300,N_24335);
nor U24556 (N_24556,N_24383,N_24322);
or U24557 (N_24557,N_24247,N_24319);
and U24558 (N_24558,N_24262,N_24308);
or U24559 (N_24559,N_24232,N_24396);
and U24560 (N_24560,N_24331,N_24258);
xor U24561 (N_24561,N_24328,N_24325);
nor U24562 (N_24562,N_24201,N_24306);
xnor U24563 (N_24563,N_24201,N_24283);
or U24564 (N_24564,N_24220,N_24376);
and U24565 (N_24565,N_24251,N_24273);
xor U24566 (N_24566,N_24313,N_24299);
xnor U24567 (N_24567,N_24393,N_24358);
nor U24568 (N_24568,N_24357,N_24276);
or U24569 (N_24569,N_24237,N_24370);
nor U24570 (N_24570,N_24380,N_24239);
and U24571 (N_24571,N_24310,N_24335);
or U24572 (N_24572,N_24355,N_24231);
nand U24573 (N_24573,N_24202,N_24263);
nand U24574 (N_24574,N_24359,N_24254);
nor U24575 (N_24575,N_24298,N_24388);
or U24576 (N_24576,N_24217,N_24368);
nor U24577 (N_24577,N_24262,N_24225);
nand U24578 (N_24578,N_24208,N_24395);
nor U24579 (N_24579,N_24362,N_24294);
xnor U24580 (N_24580,N_24208,N_24357);
and U24581 (N_24581,N_24383,N_24256);
nand U24582 (N_24582,N_24251,N_24220);
or U24583 (N_24583,N_24342,N_24301);
nor U24584 (N_24584,N_24286,N_24211);
and U24585 (N_24585,N_24309,N_24290);
and U24586 (N_24586,N_24200,N_24293);
nor U24587 (N_24587,N_24244,N_24312);
and U24588 (N_24588,N_24361,N_24330);
or U24589 (N_24589,N_24320,N_24222);
and U24590 (N_24590,N_24301,N_24278);
and U24591 (N_24591,N_24330,N_24228);
xnor U24592 (N_24592,N_24314,N_24292);
or U24593 (N_24593,N_24203,N_24325);
xor U24594 (N_24594,N_24326,N_24398);
xor U24595 (N_24595,N_24393,N_24253);
or U24596 (N_24596,N_24259,N_24325);
or U24597 (N_24597,N_24333,N_24303);
or U24598 (N_24598,N_24303,N_24357);
nand U24599 (N_24599,N_24218,N_24253);
nor U24600 (N_24600,N_24482,N_24414);
xor U24601 (N_24601,N_24504,N_24539);
xnor U24602 (N_24602,N_24585,N_24583);
or U24603 (N_24603,N_24481,N_24562);
nor U24604 (N_24604,N_24542,N_24571);
or U24605 (N_24605,N_24517,N_24590);
nand U24606 (N_24606,N_24464,N_24452);
nand U24607 (N_24607,N_24572,N_24429);
or U24608 (N_24608,N_24581,N_24554);
nand U24609 (N_24609,N_24516,N_24446);
nand U24610 (N_24610,N_24480,N_24487);
and U24611 (N_24611,N_24421,N_24410);
nand U24612 (N_24612,N_24532,N_24408);
nor U24613 (N_24613,N_24503,N_24545);
and U24614 (N_24614,N_24436,N_24460);
or U24615 (N_24615,N_24588,N_24520);
or U24616 (N_24616,N_24417,N_24467);
xnor U24617 (N_24617,N_24495,N_24580);
and U24618 (N_24618,N_24568,N_24458);
or U24619 (N_24619,N_24524,N_24594);
and U24620 (N_24620,N_24519,N_24573);
nor U24621 (N_24621,N_24457,N_24549);
xnor U24622 (N_24622,N_24440,N_24409);
nor U24623 (N_24623,N_24551,N_24559);
xor U24624 (N_24624,N_24475,N_24555);
or U24625 (N_24625,N_24454,N_24547);
and U24626 (N_24626,N_24589,N_24531);
nand U24627 (N_24627,N_24578,N_24484);
nand U24628 (N_24628,N_24445,N_24598);
or U24629 (N_24629,N_24553,N_24463);
or U24630 (N_24630,N_24587,N_24478);
or U24631 (N_24631,N_24434,N_24488);
nor U24632 (N_24632,N_24413,N_24430);
xnor U24633 (N_24633,N_24405,N_24550);
and U24634 (N_24634,N_24447,N_24570);
nor U24635 (N_24635,N_24544,N_24441);
or U24636 (N_24636,N_24599,N_24534);
nor U24637 (N_24637,N_24522,N_24528);
or U24638 (N_24638,N_24462,N_24438);
or U24639 (N_24639,N_24518,N_24401);
xor U24640 (N_24640,N_24473,N_24444);
xnor U24641 (N_24641,N_24483,N_24509);
nor U24642 (N_24642,N_24492,N_24400);
or U24643 (N_24643,N_24514,N_24508);
xnor U24644 (N_24644,N_24538,N_24455);
nor U24645 (N_24645,N_24552,N_24406);
nor U24646 (N_24646,N_24437,N_24468);
or U24647 (N_24647,N_24564,N_24422);
xnor U24648 (N_24648,N_24496,N_24432);
or U24649 (N_24649,N_24443,N_24530);
or U24650 (N_24650,N_24558,N_24505);
nand U24651 (N_24651,N_24567,N_24557);
xnor U24652 (N_24652,N_24477,N_24592);
nand U24653 (N_24653,N_24593,N_24402);
or U24654 (N_24654,N_24500,N_24561);
and U24655 (N_24655,N_24511,N_24543);
nor U24656 (N_24656,N_24565,N_24575);
or U24657 (N_24657,N_24476,N_24533);
and U24658 (N_24658,N_24425,N_24537);
xor U24659 (N_24659,N_24548,N_24506);
nand U24660 (N_24660,N_24490,N_24415);
xnor U24661 (N_24661,N_24541,N_24577);
nor U24662 (N_24662,N_24527,N_24466);
nand U24663 (N_24663,N_24403,N_24502);
nor U24664 (N_24664,N_24536,N_24470);
or U24665 (N_24665,N_24521,N_24450);
or U24666 (N_24666,N_24494,N_24510);
nand U24667 (N_24667,N_24420,N_24523);
nor U24668 (N_24668,N_24404,N_24579);
or U24669 (N_24669,N_24595,N_24563);
nor U24670 (N_24670,N_24433,N_24419);
nor U24671 (N_24671,N_24449,N_24499);
and U24672 (N_24672,N_24435,N_24472);
nor U24673 (N_24673,N_24461,N_24428);
and U24674 (N_24674,N_24423,N_24569);
xor U24675 (N_24675,N_24424,N_24546);
and U24676 (N_24676,N_24439,N_24431);
or U24677 (N_24677,N_24471,N_24584);
or U24678 (N_24678,N_24540,N_24411);
or U24679 (N_24679,N_24453,N_24448);
xor U24680 (N_24680,N_24418,N_24426);
nand U24681 (N_24681,N_24416,N_24526);
nor U24682 (N_24682,N_24582,N_24586);
or U24683 (N_24683,N_24451,N_24560);
xnor U24684 (N_24684,N_24498,N_24459);
or U24685 (N_24685,N_24576,N_24497);
nand U24686 (N_24686,N_24412,N_24525);
xnor U24687 (N_24687,N_24427,N_24491);
nor U24688 (N_24688,N_24597,N_24507);
and U24689 (N_24689,N_24493,N_24535);
nor U24690 (N_24690,N_24596,N_24574);
and U24691 (N_24691,N_24513,N_24512);
xnor U24692 (N_24692,N_24489,N_24566);
and U24693 (N_24693,N_24456,N_24529);
nand U24694 (N_24694,N_24486,N_24469);
or U24695 (N_24695,N_24407,N_24501);
and U24696 (N_24696,N_24465,N_24474);
nand U24697 (N_24697,N_24442,N_24515);
or U24698 (N_24698,N_24591,N_24485);
xnor U24699 (N_24699,N_24479,N_24556);
xor U24700 (N_24700,N_24552,N_24433);
nand U24701 (N_24701,N_24412,N_24559);
or U24702 (N_24702,N_24501,N_24424);
nor U24703 (N_24703,N_24557,N_24452);
nor U24704 (N_24704,N_24410,N_24566);
xnor U24705 (N_24705,N_24526,N_24558);
xnor U24706 (N_24706,N_24598,N_24527);
xor U24707 (N_24707,N_24598,N_24591);
xnor U24708 (N_24708,N_24551,N_24435);
and U24709 (N_24709,N_24469,N_24474);
nand U24710 (N_24710,N_24411,N_24440);
nand U24711 (N_24711,N_24464,N_24532);
or U24712 (N_24712,N_24427,N_24406);
and U24713 (N_24713,N_24459,N_24512);
nor U24714 (N_24714,N_24584,N_24578);
nand U24715 (N_24715,N_24534,N_24447);
nand U24716 (N_24716,N_24556,N_24536);
nand U24717 (N_24717,N_24525,N_24474);
xnor U24718 (N_24718,N_24538,N_24412);
xnor U24719 (N_24719,N_24475,N_24511);
nor U24720 (N_24720,N_24411,N_24454);
nor U24721 (N_24721,N_24544,N_24440);
xnor U24722 (N_24722,N_24558,N_24444);
xnor U24723 (N_24723,N_24458,N_24474);
nand U24724 (N_24724,N_24508,N_24495);
xor U24725 (N_24725,N_24496,N_24419);
and U24726 (N_24726,N_24499,N_24456);
or U24727 (N_24727,N_24513,N_24411);
nor U24728 (N_24728,N_24582,N_24430);
or U24729 (N_24729,N_24438,N_24545);
nand U24730 (N_24730,N_24449,N_24570);
and U24731 (N_24731,N_24501,N_24420);
nand U24732 (N_24732,N_24471,N_24580);
xor U24733 (N_24733,N_24420,N_24434);
or U24734 (N_24734,N_24599,N_24441);
nand U24735 (N_24735,N_24482,N_24504);
nand U24736 (N_24736,N_24419,N_24521);
xnor U24737 (N_24737,N_24420,N_24419);
nor U24738 (N_24738,N_24578,N_24449);
xor U24739 (N_24739,N_24521,N_24499);
and U24740 (N_24740,N_24473,N_24400);
nor U24741 (N_24741,N_24563,N_24475);
xor U24742 (N_24742,N_24599,N_24490);
or U24743 (N_24743,N_24597,N_24451);
nand U24744 (N_24744,N_24419,N_24555);
xnor U24745 (N_24745,N_24512,N_24501);
nand U24746 (N_24746,N_24568,N_24570);
xnor U24747 (N_24747,N_24400,N_24561);
and U24748 (N_24748,N_24491,N_24468);
xnor U24749 (N_24749,N_24527,N_24432);
and U24750 (N_24750,N_24534,N_24519);
and U24751 (N_24751,N_24459,N_24585);
nand U24752 (N_24752,N_24490,N_24561);
nor U24753 (N_24753,N_24496,N_24426);
and U24754 (N_24754,N_24450,N_24489);
and U24755 (N_24755,N_24447,N_24558);
nand U24756 (N_24756,N_24435,N_24515);
and U24757 (N_24757,N_24456,N_24558);
or U24758 (N_24758,N_24580,N_24497);
xnor U24759 (N_24759,N_24490,N_24566);
xor U24760 (N_24760,N_24513,N_24525);
and U24761 (N_24761,N_24405,N_24531);
or U24762 (N_24762,N_24542,N_24471);
nand U24763 (N_24763,N_24461,N_24530);
or U24764 (N_24764,N_24536,N_24482);
nand U24765 (N_24765,N_24533,N_24519);
xor U24766 (N_24766,N_24499,N_24498);
and U24767 (N_24767,N_24552,N_24463);
or U24768 (N_24768,N_24562,N_24533);
xor U24769 (N_24769,N_24525,N_24515);
and U24770 (N_24770,N_24436,N_24512);
xor U24771 (N_24771,N_24579,N_24437);
and U24772 (N_24772,N_24575,N_24591);
or U24773 (N_24773,N_24412,N_24595);
nor U24774 (N_24774,N_24581,N_24523);
xnor U24775 (N_24775,N_24493,N_24471);
and U24776 (N_24776,N_24482,N_24499);
and U24777 (N_24777,N_24472,N_24570);
or U24778 (N_24778,N_24440,N_24505);
or U24779 (N_24779,N_24465,N_24455);
and U24780 (N_24780,N_24560,N_24425);
nand U24781 (N_24781,N_24596,N_24590);
or U24782 (N_24782,N_24547,N_24515);
nor U24783 (N_24783,N_24460,N_24485);
nor U24784 (N_24784,N_24559,N_24570);
and U24785 (N_24785,N_24417,N_24502);
or U24786 (N_24786,N_24572,N_24590);
nor U24787 (N_24787,N_24564,N_24481);
and U24788 (N_24788,N_24444,N_24452);
nor U24789 (N_24789,N_24561,N_24519);
nor U24790 (N_24790,N_24596,N_24406);
and U24791 (N_24791,N_24444,N_24544);
nand U24792 (N_24792,N_24470,N_24414);
and U24793 (N_24793,N_24494,N_24492);
or U24794 (N_24794,N_24493,N_24445);
nand U24795 (N_24795,N_24533,N_24512);
nor U24796 (N_24796,N_24405,N_24479);
and U24797 (N_24797,N_24461,N_24529);
or U24798 (N_24798,N_24440,N_24562);
nand U24799 (N_24799,N_24472,N_24429);
and U24800 (N_24800,N_24686,N_24612);
nor U24801 (N_24801,N_24792,N_24641);
xor U24802 (N_24802,N_24746,N_24694);
or U24803 (N_24803,N_24657,N_24672);
or U24804 (N_24804,N_24780,N_24692);
nor U24805 (N_24805,N_24660,N_24718);
nor U24806 (N_24806,N_24650,N_24754);
and U24807 (N_24807,N_24713,N_24779);
xor U24808 (N_24808,N_24630,N_24653);
nand U24809 (N_24809,N_24689,N_24659);
and U24810 (N_24810,N_24733,N_24710);
nand U24811 (N_24811,N_24616,N_24678);
or U24812 (N_24812,N_24787,N_24753);
and U24813 (N_24813,N_24764,N_24605);
nand U24814 (N_24814,N_24671,N_24791);
nor U24815 (N_24815,N_24609,N_24655);
nor U24816 (N_24816,N_24624,N_24626);
nor U24817 (N_24817,N_24652,N_24720);
and U24818 (N_24818,N_24656,N_24682);
or U24819 (N_24819,N_24676,N_24606);
xor U24820 (N_24820,N_24619,N_24741);
xnor U24821 (N_24821,N_24684,N_24727);
or U24822 (N_24822,N_24679,N_24739);
nand U24823 (N_24823,N_24643,N_24778);
nand U24824 (N_24824,N_24636,N_24749);
and U24825 (N_24825,N_24799,N_24726);
xnor U24826 (N_24826,N_24697,N_24771);
or U24827 (N_24827,N_24646,N_24644);
or U24828 (N_24828,N_24761,N_24707);
or U24829 (N_24829,N_24714,N_24627);
xnor U24830 (N_24830,N_24797,N_24737);
or U24831 (N_24831,N_24700,N_24736);
xnor U24832 (N_24832,N_24751,N_24766);
nand U24833 (N_24833,N_24756,N_24603);
xnor U24834 (N_24834,N_24677,N_24629);
nor U24835 (N_24835,N_24706,N_24625);
and U24836 (N_24836,N_24776,N_24798);
and U24837 (N_24837,N_24635,N_24669);
nand U24838 (N_24838,N_24649,N_24782);
and U24839 (N_24839,N_24634,N_24775);
nand U24840 (N_24840,N_24654,N_24675);
and U24841 (N_24841,N_24685,N_24683);
nand U24842 (N_24842,N_24613,N_24765);
nand U24843 (N_24843,N_24781,N_24770);
nor U24844 (N_24844,N_24786,N_24728);
nand U24845 (N_24845,N_24610,N_24690);
or U24846 (N_24846,N_24795,N_24769);
xnor U24847 (N_24847,N_24647,N_24608);
nor U24848 (N_24848,N_24658,N_24750);
or U24849 (N_24849,N_24788,N_24696);
nand U24850 (N_24850,N_24665,N_24721);
and U24851 (N_24851,N_24607,N_24789);
nand U24852 (N_24852,N_24712,N_24763);
xnor U24853 (N_24853,N_24784,N_24663);
nor U24854 (N_24854,N_24735,N_24614);
and U24855 (N_24855,N_24703,N_24680);
nor U24856 (N_24856,N_24621,N_24725);
nor U24857 (N_24857,N_24777,N_24666);
or U24858 (N_24858,N_24785,N_24699);
nor U24859 (N_24859,N_24757,N_24734);
nand U24860 (N_24860,N_24623,N_24651);
xnor U24861 (N_24861,N_24632,N_24790);
or U24862 (N_24862,N_24773,N_24732);
nand U24863 (N_24863,N_24793,N_24615);
nand U24864 (N_24864,N_24688,N_24638);
xnor U24865 (N_24865,N_24601,N_24668);
xor U24866 (N_24866,N_24722,N_24661);
xnor U24867 (N_24867,N_24717,N_24759);
xnor U24868 (N_24868,N_24611,N_24687);
or U24869 (N_24869,N_24670,N_24724);
or U24870 (N_24870,N_24617,N_24760);
or U24871 (N_24871,N_24633,N_24637);
nor U24872 (N_24872,N_24645,N_24695);
and U24873 (N_24873,N_24631,N_24752);
nor U24874 (N_24874,N_24709,N_24744);
xnor U24875 (N_24875,N_24742,N_24796);
xor U24876 (N_24876,N_24702,N_24691);
or U24877 (N_24877,N_24794,N_24783);
xor U24878 (N_24878,N_24708,N_24715);
nor U24879 (N_24879,N_24748,N_24745);
xor U24880 (N_24880,N_24639,N_24730);
or U24881 (N_24881,N_24681,N_24620);
nor U24882 (N_24882,N_24762,N_24755);
or U24883 (N_24883,N_24674,N_24604);
nand U24884 (N_24884,N_24701,N_24693);
nor U24885 (N_24885,N_24673,N_24719);
and U24886 (N_24886,N_24618,N_24602);
xnor U24887 (N_24887,N_24711,N_24662);
nand U24888 (N_24888,N_24664,N_24731);
or U24889 (N_24889,N_24642,N_24716);
xnor U24890 (N_24890,N_24774,N_24704);
or U24891 (N_24891,N_24747,N_24628);
or U24892 (N_24892,N_24723,N_24622);
and U24893 (N_24893,N_24743,N_24648);
nor U24894 (N_24894,N_24600,N_24705);
nor U24895 (N_24895,N_24768,N_24667);
nand U24896 (N_24896,N_24758,N_24738);
nand U24897 (N_24897,N_24729,N_24767);
xnor U24898 (N_24898,N_24698,N_24772);
nor U24899 (N_24899,N_24740,N_24640);
xnor U24900 (N_24900,N_24665,N_24697);
xor U24901 (N_24901,N_24780,N_24720);
or U24902 (N_24902,N_24649,N_24717);
nor U24903 (N_24903,N_24707,N_24693);
xnor U24904 (N_24904,N_24793,N_24731);
nand U24905 (N_24905,N_24636,N_24781);
nand U24906 (N_24906,N_24603,N_24643);
or U24907 (N_24907,N_24753,N_24614);
nor U24908 (N_24908,N_24766,N_24677);
nand U24909 (N_24909,N_24785,N_24696);
nor U24910 (N_24910,N_24730,N_24663);
nor U24911 (N_24911,N_24750,N_24654);
nand U24912 (N_24912,N_24798,N_24600);
nand U24913 (N_24913,N_24708,N_24662);
nor U24914 (N_24914,N_24771,N_24603);
nor U24915 (N_24915,N_24665,N_24620);
or U24916 (N_24916,N_24607,N_24702);
xor U24917 (N_24917,N_24780,N_24702);
and U24918 (N_24918,N_24790,N_24742);
nor U24919 (N_24919,N_24619,N_24612);
xnor U24920 (N_24920,N_24730,N_24601);
or U24921 (N_24921,N_24632,N_24657);
or U24922 (N_24922,N_24642,N_24789);
or U24923 (N_24923,N_24769,N_24605);
nor U24924 (N_24924,N_24730,N_24628);
nor U24925 (N_24925,N_24710,N_24739);
or U24926 (N_24926,N_24772,N_24603);
or U24927 (N_24927,N_24795,N_24648);
xor U24928 (N_24928,N_24659,N_24757);
nor U24929 (N_24929,N_24687,N_24699);
nand U24930 (N_24930,N_24666,N_24761);
or U24931 (N_24931,N_24706,N_24606);
or U24932 (N_24932,N_24629,N_24752);
xnor U24933 (N_24933,N_24643,N_24654);
nand U24934 (N_24934,N_24713,N_24641);
and U24935 (N_24935,N_24646,N_24721);
nand U24936 (N_24936,N_24794,N_24744);
xor U24937 (N_24937,N_24793,N_24796);
nor U24938 (N_24938,N_24684,N_24778);
or U24939 (N_24939,N_24668,N_24786);
nor U24940 (N_24940,N_24619,N_24742);
or U24941 (N_24941,N_24735,N_24731);
or U24942 (N_24942,N_24634,N_24691);
nand U24943 (N_24943,N_24725,N_24680);
nand U24944 (N_24944,N_24663,N_24631);
nand U24945 (N_24945,N_24671,N_24703);
xor U24946 (N_24946,N_24665,N_24686);
or U24947 (N_24947,N_24729,N_24619);
or U24948 (N_24948,N_24761,N_24770);
xor U24949 (N_24949,N_24611,N_24750);
or U24950 (N_24950,N_24713,N_24617);
or U24951 (N_24951,N_24721,N_24784);
or U24952 (N_24952,N_24727,N_24651);
and U24953 (N_24953,N_24673,N_24618);
or U24954 (N_24954,N_24750,N_24613);
and U24955 (N_24955,N_24757,N_24622);
nand U24956 (N_24956,N_24683,N_24632);
or U24957 (N_24957,N_24755,N_24786);
nand U24958 (N_24958,N_24770,N_24762);
and U24959 (N_24959,N_24674,N_24718);
xnor U24960 (N_24960,N_24734,N_24652);
xor U24961 (N_24961,N_24663,N_24607);
xnor U24962 (N_24962,N_24659,N_24676);
or U24963 (N_24963,N_24770,N_24606);
xnor U24964 (N_24964,N_24746,N_24774);
nand U24965 (N_24965,N_24729,N_24645);
nand U24966 (N_24966,N_24717,N_24677);
nor U24967 (N_24967,N_24724,N_24634);
xnor U24968 (N_24968,N_24608,N_24793);
and U24969 (N_24969,N_24601,N_24697);
and U24970 (N_24970,N_24773,N_24768);
nor U24971 (N_24971,N_24717,N_24735);
xor U24972 (N_24972,N_24715,N_24601);
nor U24973 (N_24973,N_24711,N_24757);
and U24974 (N_24974,N_24757,N_24677);
or U24975 (N_24975,N_24726,N_24632);
nand U24976 (N_24976,N_24646,N_24643);
or U24977 (N_24977,N_24752,N_24737);
nand U24978 (N_24978,N_24750,N_24644);
and U24979 (N_24979,N_24622,N_24756);
xor U24980 (N_24980,N_24658,N_24664);
and U24981 (N_24981,N_24673,N_24635);
nand U24982 (N_24982,N_24643,N_24743);
nor U24983 (N_24983,N_24722,N_24725);
and U24984 (N_24984,N_24655,N_24764);
nor U24985 (N_24985,N_24617,N_24615);
xor U24986 (N_24986,N_24773,N_24685);
or U24987 (N_24987,N_24736,N_24634);
xor U24988 (N_24988,N_24661,N_24775);
and U24989 (N_24989,N_24618,N_24765);
nand U24990 (N_24990,N_24708,N_24782);
nor U24991 (N_24991,N_24695,N_24717);
nor U24992 (N_24992,N_24726,N_24656);
and U24993 (N_24993,N_24651,N_24765);
xor U24994 (N_24994,N_24626,N_24678);
nor U24995 (N_24995,N_24796,N_24619);
nor U24996 (N_24996,N_24669,N_24783);
nor U24997 (N_24997,N_24695,N_24720);
and U24998 (N_24998,N_24744,N_24731);
nand U24999 (N_24999,N_24656,N_24798);
and UO_0 (O_0,N_24933,N_24873);
and UO_1 (O_1,N_24832,N_24901);
nor UO_2 (O_2,N_24982,N_24917);
xor UO_3 (O_3,N_24930,N_24979);
xor UO_4 (O_4,N_24907,N_24958);
or UO_5 (O_5,N_24805,N_24964);
xnor UO_6 (O_6,N_24929,N_24921);
xnor UO_7 (O_7,N_24851,N_24992);
xnor UO_8 (O_8,N_24881,N_24820);
or UO_9 (O_9,N_24926,N_24840);
nand UO_10 (O_10,N_24827,N_24807);
nand UO_11 (O_11,N_24934,N_24825);
nand UO_12 (O_12,N_24856,N_24898);
xnor UO_13 (O_13,N_24816,N_24863);
xnor UO_14 (O_14,N_24951,N_24806);
or UO_15 (O_15,N_24997,N_24976);
or UO_16 (O_16,N_24868,N_24889);
nor UO_17 (O_17,N_24937,N_24919);
xnor UO_18 (O_18,N_24974,N_24800);
nor UO_19 (O_19,N_24986,N_24936);
and UO_20 (O_20,N_24990,N_24874);
nor UO_21 (O_21,N_24989,N_24996);
and UO_22 (O_22,N_24834,N_24880);
and UO_23 (O_23,N_24962,N_24941);
nor UO_24 (O_24,N_24862,N_24826);
nor UO_25 (O_25,N_24855,N_24885);
and UO_26 (O_26,N_24954,N_24943);
and UO_27 (O_27,N_24955,N_24945);
and UO_28 (O_28,N_24886,N_24876);
or UO_29 (O_29,N_24890,N_24944);
nor UO_30 (O_30,N_24912,N_24858);
and UO_31 (O_31,N_24975,N_24870);
or UO_32 (O_32,N_24904,N_24891);
or UO_33 (O_33,N_24994,N_24985);
xor UO_34 (O_34,N_24804,N_24852);
and UO_35 (O_35,N_24847,N_24903);
and UO_36 (O_36,N_24987,N_24939);
and UO_37 (O_37,N_24893,N_24812);
nor UO_38 (O_38,N_24935,N_24818);
nor UO_39 (O_39,N_24861,N_24981);
nand UO_40 (O_40,N_24824,N_24838);
nand UO_41 (O_41,N_24931,N_24947);
or UO_42 (O_42,N_24938,N_24984);
or UO_43 (O_43,N_24978,N_24969);
or UO_44 (O_44,N_24965,N_24846);
nand UO_45 (O_45,N_24882,N_24908);
and UO_46 (O_46,N_24942,N_24869);
nand UO_47 (O_47,N_24957,N_24872);
and UO_48 (O_48,N_24822,N_24853);
nor UO_49 (O_49,N_24971,N_24854);
and UO_50 (O_50,N_24860,N_24980);
xor UO_51 (O_51,N_24879,N_24814);
nand UO_52 (O_52,N_24963,N_24956);
nand UO_53 (O_53,N_24831,N_24923);
or UO_54 (O_54,N_24914,N_24915);
nor UO_55 (O_55,N_24850,N_24928);
and UO_56 (O_56,N_24884,N_24995);
xnor UO_57 (O_57,N_24845,N_24843);
xnor UO_58 (O_58,N_24913,N_24988);
nor UO_59 (O_59,N_24911,N_24828);
or UO_60 (O_60,N_24888,N_24829);
nor UO_61 (O_61,N_24909,N_24849);
nand UO_62 (O_62,N_24906,N_24925);
nor UO_63 (O_63,N_24808,N_24837);
nand UO_64 (O_64,N_24833,N_24916);
and UO_65 (O_65,N_24966,N_24950);
xor UO_66 (O_66,N_24864,N_24859);
nor UO_67 (O_67,N_24922,N_24877);
and UO_68 (O_68,N_24823,N_24887);
nor UO_69 (O_69,N_24835,N_24927);
xnor UO_70 (O_70,N_24839,N_24910);
nand UO_71 (O_71,N_24968,N_24948);
and UO_72 (O_72,N_24866,N_24841);
and UO_73 (O_73,N_24848,N_24883);
nor UO_74 (O_74,N_24801,N_24918);
and UO_75 (O_75,N_24811,N_24932);
and UO_76 (O_76,N_24892,N_24844);
or UO_77 (O_77,N_24821,N_24993);
nand UO_78 (O_78,N_24857,N_24842);
or UO_79 (O_79,N_24952,N_24819);
xor UO_80 (O_80,N_24977,N_24894);
nand UO_81 (O_81,N_24896,N_24961);
and UO_82 (O_82,N_24953,N_24875);
xor UO_83 (O_83,N_24803,N_24920);
nor UO_84 (O_84,N_24991,N_24946);
and UO_85 (O_85,N_24865,N_24836);
or UO_86 (O_86,N_24999,N_24967);
or UO_87 (O_87,N_24972,N_24830);
nand UO_88 (O_88,N_24815,N_24895);
nor UO_89 (O_89,N_24878,N_24960);
xor UO_90 (O_90,N_24949,N_24802);
and UO_91 (O_91,N_24810,N_24902);
or UO_92 (O_92,N_24970,N_24940);
xor UO_93 (O_93,N_24809,N_24924);
and UO_94 (O_94,N_24897,N_24900);
nor UO_95 (O_95,N_24871,N_24983);
nor UO_96 (O_96,N_24817,N_24998);
nand UO_97 (O_97,N_24867,N_24899);
or UO_98 (O_98,N_24959,N_24973);
xor UO_99 (O_99,N_24905,N_24813);
or UO_100 (O_100,N_24984,N_24807);
and UO_101 (O_101,N_24812,N_24885);
xor UO_102 (O_102,N_24916,N_24854);
nor UO_103 (O_103,N_24834,N_24876);
and UO_104 (O_104,N_24833,N_24889);
nor UO_105 (O_105,N_24864,N_24801);
xnor UO_106 (O_106,N_24868,N_24835);
or UO_107 (O_107,N_24888,N_24894);
or UO_108 (O_108,N_24912,N_24861);
or UO_109 (O_109,N_24964,N_24909);
nor UO_110 (O_110,N_24998,N_24933);
or UO_111 (O_111,N_24847,N_24997);
nand UO_112 (O_112,N_24899,N_24880);
nor UO_113 (O_113,N_24914,N_24995);
nand UO_114 (O_114,N_24980,N_24987);
xnor UO_115 (O_115,N_24979,N_24809);
nor UO_116 (O_116,N_24960,N_24965);
xnor UO_117 (O_117,N_24875,N_24924);
nor UO_118 (O_118,N_24899,N_24837);
and UO_119 (O_119,N_24841,N_24887);
and UO_120 (O_120,N_24905,N_24830);
or UO_121 (O_121,N_24959,N_24862);
and UO_122 (O_122,N_24822,N_24910);
and UO_123 (O_123,N_24889,N_24848);
nand UO_124 (O_124,N_24887,N_24814);
xnor UO_125 (O_125,N_24879,N_24820);
nor UO_126 (O_126,N_24830,N_24844);
or UO_127 (O_127,N_24856,N_24806);
and UO_128 (O_128,N_24938,N_24885);
and UO_129 (O_129,N_24963,N_24858);
nand UO_130 (O_130,N_24865,N_24969);
or UO_131 (O_131,N_24984,N_24931);
and UO_132 (O_132,N_24805,N_24944);
nand UO_133 (O_133,N_24891,N_24821);
nor UO_134 (O_134,N_24895,N_24945);
nor UO_135 (O_135,N_24957,N_24853);
or UO_136 (O_136,N_24842,N_24954);
and UO_137 (O_137,N_24925,N_24944);
nor UO_138 (O_138,N_24951,N_24974);
nand UO_139 (O_139,N_24863,N_24879);
nor UO_140 (O_140,N_24860,N_24909);
xnor UO_141 (O_141,N_24920,N_24815);
and UO_142 (O_142,N_24816,N_24975);
xnor UO_143 (O_143,N_24965,N_24806);
nand UO_144 (O_144,N_24822,N_24887);
and UO_145 (O_145,N_24894,N_24893);
nand UO_146 (O_146,N_24809,N_24862);
xor UO_147 (O_147,N_24968,N_24974);
and UO_148 (O_148,N_24923,N_24909);
nor UO_149 (O_149,N_24920,N_24900);
and UO_150 (O_150,N_24988,N_24897);
nand UO_151 (O_151,N_24908,N_24935);
xnor UO_152 (O_152,N_24973,N_24825);
nand UO_153 (O_153,N_24906,N_24979);
or UO_154 (O_154,N_24836,N_24921);
or UO_155 (O_155,N_24851,N_24980);
or UO_156 (O_156,N_24955,N_24895);
nand UO_157 (O_157,N_24828,N_24896);
nand UO_158 (O_158,N_24850,N_24874);
nand UO_159 (O_159,N_24854,N_24880);
xnor UO_160 (O_160,N_24878,N_24966);
and UO_161 (O_161,N_24915,N_24960);
nor UO_162 (O_162,N_24978,N_24809);
nand UO_163 (O_163,N_24838,N_24976);
nand UO_164 (O_164,N_24927,N_24909);
xor UO_165 (O_165,N_24832,N_24916);
nor UO_166 (O_166,N_24935,N_24953);
nor UO_167 (O_167,N_24997,N_24844);
nand UO_168 (O_168,N_24924,N_24886);
xnor UO_169 (O_169,N_24923,N_24807);
nand UO_170 (O_170,N_24837,N_24937);
xor UO_171 (O_171,N_24871,N_24940);
nand UO_172 (O_172,N_24879,N_24909);
or UO_173 (O_173,N_24953,N_24833);
nor UO_174 (O_174,N_24864,N_24929);
or UO_175 (O_175,N_24944,N_24824);
and UO_176 (O_176,N_24973,N_24870);
or UO_177 (O_177,N_24976,N_24980);
or UO_178 (O_178,N_24936,N_24861);
nand UO_179 (O_179,N_24969,N_24955);
nand UO_180 (O_180,N_24893,N_24869);
nor UO_181 (O_181,N_24816,N_24872);
nand UO_182 (O_182,N_24964,N_24930);
xnor UO_183 (O_183,N_24934,N_24861);
xor UO_184 (O_184,N_24898,N_24875);
nor UO_185 (O_185,N_24924,N_24980);
nand UO_186 (O_186,N_24854,N_24856);
nor UO_187 (O_187,N_24946,N_24976);
xor UO_188 (O_188,N_24839,N_24918);
or UO_189 (O_189,N_24842,N_24804);
nor UO_190 (O_190,N_24950,N_24929);
nor UO_191 (O_191,N_24969,N_24925);
xor UO_192 (O_192,N_24814,N_24831);
xor UO_193 (O_193,N_24820,N_24842);
and UO_194 (O_194,N_24948,N_24964);
nor UO_195 (O_195,N_24867,N_24986);
or UO_196 (O_196,N_24833,N_24880);
or UO_197 (O_197,N_24964,N_24810);
nand UO_198 (O_198,N_24882,N_24928);
nand UO_199 (O_199,N_24979,N_24848);
nor UO_200 (O_200,N_24992,N_24972);
nand UO_201 (O_201,N_24831,N_24905);
nor UO_202 (O_202,N_24917,N_24977);
nand UO_203 (O_203,N_24800,N_24803);
nand UO_204 (O_204,N_24965,N_24898);
nor UO_205 (O_205,N_24994,N_24986);
xor UO_206 (O_206,N_24832,N_24898);
nor UO_207 (O_207,N_24836,N_24812);
and UO_208 (O_208,N_24969,N_24856);
xnor UO_209 (O_209,N_24880,N_24860);
xnor UO_210 (O_210,N_24800,N_24937);
xnor UO_211 (O_211,N_24942,N_24823);
nand UO_212 (O_212,N_24917,N_24827);
nor UO_213 (O_213,N_24810,N_24919);
and UO_214 (O_214,N_24838,N_24896);
and UO_215 (O_215,N_24853,N_24951);
and UO_216 (O_216,N_24848,N_24902);
nor UO_217 (O_217,N_24871,N_24810);
nand UO_218 (O_218,N_24998,N_24976);
nor UO_219 (O_219,N_24848,N_24846);
nor UO_220 (O_220,N_24920,N_24868);
nand UO_221 (O_221,N_24983,N_24988);
nand UO_222 (O_222,N_24998,N_24895);
nor UO_223 (O_223,N_24967,N_24922);
and UO_224 (O_224,N_24916,N_24892);
and UO_225 (O_225,N_24948,N_24966);
xor UO_226 (O_226,N_24844,N_24946);
or UO_227 (O_227,N_24875,N_24950);
nor UO_228 (O_228,N_24996,N_24907);
or UO_229 (O_229,N_24871,N_24870);
or UO_230 (O_230,N_24992,N_24964);
xor UO_231 (O_231,N_24937,N_24810);
nand UO_232 (O_232,N_24880,N_24870);
xor UO_233 (O_233,N_24813,N_24898);
or UO_234 (O_234,N_24938,N_24933);
nor UO_235 (O_235,N_24911,N_24926);
or UO_236 (O_236,N_24903,N_24819);
and UO_237 (O_237,N_24830,N_24989);
nor UO_238 (O_238,N_24833,N_24837);
or UO_239 (O_239,N_24867,N_24998);
xnor UO_240 (O_240,N_24935,N_24861);
and UO_241 (O_241,N_24915,N_24892);
or UO_242 (O_242,N_24994,N_24938);
and UO_243 (O_243,N_24976,N_24956);
nand UO_244 (O_244,N_24965,N_24880);
xor UO_245 (O_245,N_24965,N_24847);
xor UO_246 (O_246,N_24992,N_24959);
xnor UO_247 (O_247,N_24992,N_24893);
nor UO_248 (O_248,N_24894,N_24801);
nor UO_249 (O_249,N_24988,N_24880);
xnor UO_250 (O_250,N_24956,N_24906);
and UO_251 (O_251,N_24870,N_24898);
nand UO_252 (O_252,N_24881,N_24933);
xor UO_253 (O_253,N_24975,N_24903);
nand UO_254 (O_254,N_24854,N_24805);
nor UO_255 (O_255,N_24913,N_24930);
xor UO_256 (O_256,N_24873,N_24951);
nand UO_257 (O_257,N_24886,N_24999);
nand UO_258 (O_258,N_24818,N_24863);
and UO_259 (O_259,N_24903,N_24933);
or UO_260 (O_260,N_24940,N_24895);
xnor UO_261 (O_261,N_24924,N_24907);
or UO_262 (O_262,N_24916,N_24910);
xor UO_263 (O_263,N_24984,N_24936);
or UO_264 (O_264,N_24900,N_24936);
nand UO_265 (O_265,N_24937,N_24877);
nor UO_266 (O_266,N_24954,N_24869);
nand UO_267 (O_267,N_24817,N_24884);
or UO_268 (O_268,N_24853,N_24949);
nor UO_269 (O_269,N_24874,N_24868);
xor UO_270 (O_270,N_24988,N_24834);
nand UO_271 (O_271,N_24900,N_24986);
nand UO_272 (O_272,N_24931,N_24835);
or UO_273 (O_273,N_24962,N_24843);
nand UO_274 (O_274,N_24924,N_24965);
xnor UO_275 (O_275,N_24847,N_24835);
and UO_276 (O_276,N_24887,N_24935);
and UO_277 (O_277,N_24998,N_24942);
nor UO_278 (O_278,N_24966,N_24884);
nor UO_279 (O_279,N_24895,N_24967);
or UO_280 (O_280,N_24812,N_24816);
nor UO_281 (O_281,N_24826,N_24987);
nand UO_282 (O_282,N_24803,N_24968);
nand UO_283 (O_283,N_24886,N_24842);
or UO_284 (O_284,N_24863,N_24916);
and UO_285 (O_285,N_24832,N_24864);
and UO_286 (O_286,N_24898,N_24896);
nor UO_287 (O_287,N_24824,N_24891);
nor UO_288 (O_288,N_24884,N_24840);
nand UO_289 (O_289,N_24812,N_24928);
xnor UO_290 (O_290,N_24832,N_24809);
nor UO_291 (O_291,N_24822,N_24978);
and UO_292 (O_292,N_24811,N_24817);
xor UO_293 (O_293,N_24834,N_24960);
or UO_294 (O_294,N_24964,N_24870);
and UO_295 (O_295,N_24850,N_24945);
xnor UO_296 (O_296,N_24894,N_24835);
nand UO_297 (O_297,N_24875,N_24907);
or UO_298 (O_298,N_24978,N_24861);
nand UO_299 (O_299,N_24963,N_24803);
and UO_300 (O_300,N_24966,N_24868);
and UO_301 (O_301,N_24874,N_24996);
nand UO_302 (O_302,N_24896,N_24977);
nor UO_303 (O_303,N_24893,N_24877);
or UO_304 (O_304,N_24908,N_24947);
and UO_305 (O_305,N_24871,N_24986);
xor UO_306 (O_306,N_24920,N_24980);
nand UO_307 (O_307,N_24886,N_24910);
xor UO_308 (O_308,N_24926,N_24906);
or UO_309 (O_309,N_24894,N_24934);
xor UO_310 (O_310,N_24809,N_24860);
nand UO_311 (O_311,N_24964,N_24961);
or UO_312 (O_312,N_24810,N_24898);
and UO_313 (O_313,N_24801,N_24938);
nand UO_314 (O_314,N_24923,N_24927);
xor UO_315 (O_315,N_24861,N_24801);
or UO_316 (O_316,N_24964,N_24950);
xor UO_317 (O_317,N_24818,N_24817);
or UO_318 (O_318,N_24940,N_24904);
xor UO_319 (O_319,N_24929,N_24830);
or UO_320 (O_320,N_24926,N_24969);
xnor UO_321 (O_321,N_24823,N_24913);
xnor UO_322 (O_322,N_24897,N_24895);
xnor UO_323 (O_323,N_24905,N_24895);
or UO_324 (O_324,N_24821,N_24976);
and UO_325 (O_325,N_24950,N_24987);
nand UO_326 (O_326,N_24804,N_24887);
or UO_327 (O_327,N_24967,N_24827);
or UO_328 (O_328,N_24838,N_24832);
or UO_329 (O_329,N_24989,N_24865);
xor UO_330 (O_330,N_24954,N_24895);
and UO_331 (O_331,N_24973,N_24920);
xnor UO_332 (O_332,N_24815,N_24913);
xor UO_333 (O_333,N_24998,N_24982);
and UO_334 (O_334,N_24863,N_24827);
nand UO_335 (O_335,N_24969,N_24882);
xnor UO_336 (O_336,N_24838,N_24844);
nor UO_337 (O_337,N_24928,N_24858);
and UO_338 (O_338,N_24939,N_24871);
nor UO_339 (O_339,N_24939,N_24984);
xor UO_340 (O_340,N_24845,N_24864);
and UO_341 (O_341,N_24920,N_24826);
nand UO_342 (O_342,N_24844,N_24920);
xor UO_343 (O_343,N_24841,N_24832);
nand UO_344 (O_344,N_24928,N_24918);
nand UO_345 (O_345,N_24992,N_24981);
nor UO_346 (O_346,N_24968,N_24984);
or UO_347 (O_347,N_24933,N_24959);
or UO_348 (O_348,N_24951,N_24978);
nor UO_349 (O_349,N_24984,N_24817);
nand UO_350 (O_350,N_24846,N_24877);
and UO_351 (O_351,N_24978,N_24929);
nor UO_352 (O_352,N_24951,N_24975);
and UO_353 (O_353,N_24935,N_24814);
nand UO_354 (O_354,N_24943,N_24892);
nand UO_355 (O_355,N_24993,N_24809);
and UO_356 (O_356,N_24907,N_24934);
and UO_357 (O_357,N_24810,N_24801);
nand UO_358 (O_358,N_24987,N_24933);
and UO_359 (O_359,N_24989,N_24912);
and UO_360 (O_360,N_24974,N_24909);
nand UO_361 (O_361,N_24829,N_24916);
xor UO_362 (O_362,N_24855,N_24852);
xnor UO_363 (O_363,N_24954,N_24818);
xnor UO_364 (O_364,N_24997,N_24961);
or UO_365 (O_365,N_24898,N_24900);
and UO_366 (O_366,N_24892,N_24997);
and UO_367 (O_367,N_24822,N_24927);
nor UO_368 (O_368,N_24963,N_24941);
and UO_369 (O_369,N_24983,N_24982);
xnor UO_370 (O_370,N_24924,N_24837);
or UO_371 (O_371,N_24909,N_24945);
nor UO_372 (O_372,N_24993,N_24963);
nand UO_373 (O_373,N_24849,N_24845);
nand UO_374 (O_374,N_24918,N_24916);
or UO_375 (O_375,N_24918,N_24891);
nand UO_376 (O_376,N_24948,N_24940);
or UO_377 (O_377,N_24947,N_24905);
or UO_378 (O_378,N_24889,N_24907);
and UO_379 (O_379,N_24958,N_24845);
xnor UO_380 (O_380,N_24976,N_24841);
xor UO_381 (O_381,N_24813,N_24839);
or UO_382 (O_382,N_24980,N_24931);
or UO_383 (O_383,N_24814,N_24856);
nand UO_384 (O_384,N_24932,N_24875);
and UO_385 (O_385,N_24969,N_24922);
xnor UO_386 (O_386,N_24971,N_24917);
xnor UO_387 (O_387,N_24886,N_24885);
xor UO_388 (O_388,N_24940,N_24985);
xnor UO_389 (O_389,N_24823,N_24844);
or UO_390 (O_390,N_24918,N_24895);
and UO_391 (O_391,N_24927,N_24944);
xor UO_392 (O_392,N_24857,N_24805);
xor UO_393 (O_393,N_24999,N_24998);
nand UO_394 (O_394,N_24994,N_24932);
or UO_395 (O_395,N_24963,N_24891);
xnor UO_396 (O_396,N_24886,N_24996);
and UO_397 (O_397,N_24812,N_24846);
or UO_398 (O_398,N_24805,N_24821);
or UO_399 (O_399,N_24948,N_24849);
nand UO_400 (O_400,N_24882,N_24934);
nor UO_401 (O_401,N_24912,N_24917);
nor UO_402 (O_402,N_24906,N_24998);
or UO_403 (O_403,N_24923,N_24939);
nor UO_404 (O_404,N_24884,N_24829);
or UO_405 (O_405,N_24992,N_24895);
xor UO_406 (O_406,N_24822,N_24889);
or UO_407 (O_407,N_24900,N_24863);
xor UO_408 (O_408,N_24921,N_24811);
xor UO_409 (O_409,N_24940,N_24979);
and UO_410 (O_410,N_24893,N_24800);
xor UO_411 (O_411,N_24862,N_24825);
and UO_412 (O_412,N_24811,N_24867);
nor UO_413 (O_413,N_24896,N_24945);
nand UO_414 (O_414,N_24843,N_24965);
and UO_415 (O_415,N_24879,N_24836);
and UO_416 (O_416,N_24947,N_24956);
nor UO_417 (O_417,N_24969,N_24898);
and UO_418 (O_418,N_24945,N_24838);
nor UO_419 (O_419,N_24985,N_24900);
and UO_420 (O_420,N_24991,N_24904);
nor UO_421 (O_421,N_24836,N_24954);
and UO_422 (O_422,N_24958,N_24822);
and UO_423 (O_423,N_24937,N_24889);
or UO_424 (O_424,N_24994,N_24900);
nand UO_425 (O_425,N_24959,N_24876);
xnor UO_426 (O_426,N_24870,N_24962);
or UO_427 (O_427,N_24952,N_24986);
or UO_428 (O_428,N_24882,N_24832);
xor UO_429 (O_429,N_24990,N_24806);
xor UO_430 (O_430,N_24822,N_24961);
nand UO_431 (O_431,N_24877,N_24873);
and UO_432 (O_432,N_24842,N_24818);
nor UO_433 (O_433,N_24935,N_24888);
nand UO_434 (O_434,N_24976,N_24837);
or UO_435 (O_435,N_24811,N_24880);
nor UO_436 (O_436,N_24974,N_24877);
nand UO_437 (O_437,N_24935,N_24957);
xnor UO_438 (O_438,N_24861,N_24868);
or UO_439 (O_439,N_24856,N_24878);
and UO_440 (O_440,N_24889,N_24859);
xnor UO_441 (O_441,N_24922,N_24940);
nor UO_442 (O_442,N_24931,N_24956);
nand UO_443 (O_443,N_24820,N_24965);
and UO_444 (O_444,N_24808,N_24998);
nand UO_445 (O_445,N_24930,N_24981);
xor UO_446 (O_446,N_24907,N_24811);
nand UO_447 (O_447,N_24860,N_24828);
nand UO_448 (O_448,N_24833,N_24927);
and UO_449 (O_449,N_24859,N_24957);
nor UO_450 (O_450,N_24966,N_24805);
nor UO_451 (O_451,N_24849,N_24893);
nand UO_452 (O_452,N_24995,N_24862);
and UO_453 (O_453,N_24860,N_24879);
nor UO_454 (O_454,N_24863,N_24941);
nor UO_455 (O_455,N_24805,N_24843);
xnor UO_456 (O_456,N_24847,N_24933);
nor UO_457 (O_457,N_24873,N_24917);
nor UO_458 (O_458,N_24810,N_24867);
nand UO_459 (O_459,N_24956,N_24893);
and UO_460 (O_460,N_24923,N_24950);
nor UO_461 (O_461,N_24871,N_24888);
or UO_462 (O_462,N_24906,N_24908);
xor UO_463 (O_463,N_24890,N_24892);
xnor UO_464 (O_464,N_24878,N_24913);
nor UO_465 (O_465,N_24931,N_24823);
and UO_466 (O_466,N_24813,N_24971);
nand UO_467 (O_467,N_24994,N_24957);
xnor UO_468 (O_468,N_24818,N_24925);
nand UO_469 (O_469,N_24840,N_24873);
nand UO_470 (O_470,N_24884,N_24836);
xnor UO_471 (O_471,N_24829,N_24903);
or UO_472 (O_472,N_24881,N_24900);
or UO_473 (O_473,N_24904,N_24838);
xor UO_474 (O_474,N_24895,N_24821);
and UO_475 (O_475,N_24827,N_24914);
or UO_476 (O_476,N_24824,N_24921);
nor UO_477 (O_477,N_24969,N_24994);
nand UO_478 (O_478,N_24880,N_24937);
nor UO_479 (O_479,N_24983,N_24958);
xor UO_480 (O_480,N_24910,N_24870);
or UO_481 (O_481,N_24948,N_24836);
and UO_482 (O_482,N_24972,N_24928);
or UO_483 (O_483,N_24960,N_24806);
and UO_484 (O_484,N_24900,N_24848);
or UO_485 (O_485,N_24878,N_24956);
nand UO_486 (O_486,N_24849,N_24925);
nor UO_487 (O_487,N_24895,N_24853);
nand UO_488 (O_488,N_24887,N_24845);
xnor UO_489 (O_489,N_24911,N_24930);
or UO_490 (O_490,N_24885,N_24908);
or UO_491 (O_491,N_24807,N_24928);
or UO_492 (O_492,N_24855,N_24898);
nor UO_493 (O_493,N_24908,N_24957);
xnor UO_494 (O_494,N_24863,N_24917);
and UO_495 (O_495,N_24813,N_24872);
and UO_496 (O_496,N_24996,N_24922);
nand UO_497 (O_497,N_24895,N_24868);
xnor UO_498 (O_498,N_24881,N_24848);
and UO_499 (O_499,N_24935,N_24996);
and UO_500 (O_500,N_24887,N_24928);
xor UO_501 (O_501,N_24990,N_24921);
or UO_502 (O_502,N_24898,N_24977);
or UO_503 (O_503,N_24871,N_24876);
xor UO_504 (O_504,N_24872,N_24822);
nand UO_505 (O_505,N_24822,N_24918);
or UO_506 (O_506,N_24963,N_24817);
and UO_507 (O_507,N_24834,N_24955);
xnor UO_508 (O_508,N_24829,N_24864);
or UO_509 (O_509,N_24932,N_24966);
xor UO_510 (O_510,N_24882,N_24957);
and UO_511 (O_511,N_24951,N_24948);
and UO_512 (O_512,N_24896,N_24835);
nand UO_513 (O_513,N_24821,N_24806);
or UO_514 (O_514,N_24917,N_24807);
and UO_515 (O_515,N_24862,N_24956);
and UO_516 (O_516,N_24985,N_24884);
nand UO_517 (O_517,N_24890,N_24868);
xnor UO_518 (O_518,N_24921,N_24803);
and UO_519 (O_519,N_24915,N_24966);
nor UO_520 (O_520,N_24852,N_24885);
or UO_521 (O_521,N_24807,N_24952);
xnor UO_522 (O_522,N_24905,N_24815);
and UO_523 (O_523,N_24820,N_24917);
nand UO_524 (O_524,N_24940,N_24967);
nand UO_525 (O_525,N_24942,N_24847);
xnor UO_526 (O_526,N_24987,N_24964);
nand UO_527 (O_527,N_24831,N_24901);
and UO_528 (O_528,N_24927,N_24906);
and UO_529 (O_529,N_24995,N_24953);
xor UO_530 (O_530,N_24949,N_24933);
nand UO_531 (O_531,N_24876,N_24934);
nand UO_532 (O_532,N_24876,N_24801);
or UO_533 (O_533,N_24991,N_24892);
nand UO_534 (O_534,N_24889,N_24828);
xor UO_535 (O_535,N_24953,N_24879);
nor UO_536 (O_536,N_24803,N_24870);
nand UO_537 (O_537,N_24823,N_24814);
nand UO_538 (O_538,N_24915,N_24808);
and UO_539 (O_539,N_24860,N_24959);
nand UO_540 (O_540,N_24844,N_24954);
nor UO_541 (O_541,N_24929,N_24940);
nand UO_542 (O_542,N_24832,N_24899);
or UO_543 (O_543,N_24852,N_24833);
xor UO_544 (O_544,N_24951,N_24810);
or UO_545 (O_545,N_24907,N_24942);
nor UO_546 (O_546,N_24992,N_24866);
xnor UO_547 (O_547,N_24903,N_24924);
xnor UO_548 (O_548,N_24966,N_24936);
and UO_549 (O_549,N_24913,N_24839);
nand UO_550 (O_550,N_24935,N_24985);
nor UO_551 (O_551,N_24855,N_24817);
or UO_552 (O_552,N_24940,N_24824);
xor UO_553 (O_553,N_24966,N_24903);
nor UO_554 (O_554,N_24977,N_24949);
nand UO_555 (O_555,N_24897,N_24925);
or UO_556 (O_556,N_24846,N_24906);
nand UO_557 (O_557,N_24929,N_24986);
nand UO_558 (O_558,N_24896,N_24819);
nand UO_559 (O_559,N_24837,N_24878);
xor UO_560 (O_560,N_24818,N_24845);
and UO_561 (O_561,N_24972,N_24932);
nand UO_562 (O_562,N_24834,N_24852);
and UO_563 (O_563,N_24915,N_24867);
xor UO_564 (O_564,N_24861,N_24812);
and UO_565 (O_565,N_24879,N_24918);
xor UO_566 (O_566,N_24942,N_24911);
and UO_567 (O_567,N_24948,N_24979);
or UO_568 (O_568,N_24976,N_24979);
nand UO_569 (O_569,N_24828,N_24960);
nor UO_570 (O_570,N_24949,N_24842);
or UO_571 (O_571,N_24913,N_24904);
nand UO_572 (O_572,N_24849,N_24837);
nor UO_573 (O_573,N_24802,N_24953);
xnor UO_574 (O_574,N_24846,N_24904);
and UO_575 (O_575,N_24841,N_24942);
xnor UO_576 (O_576,N_24958,N_24865);
xor UO_577 (O_577,N_24971,N_24990);
nand UO_578 (O_578,N_24987,N_24923);
nor UO_579 (O_579,N_24803,N_24822);
xnor UO_580 (O_580,N_24984,N_24917);
nand UO_581 (O_581,N_24910,N_24858);
nand UO_582 (O_582,N_24857,N_24881);
xor UO_583 (O_583,N_24864,N_24858);
and UO_584 (O_584,N_24885,N_24959);
nand UO_585 (O_585,N_24940,N_24943);
xnor UO_586 (O_586,N_24855,N_24985);
and UO_587 (O_587,N_24822,N_24903);
nand UO_588 (O_588,N_24887,N_24875);
and UO_589 (O_589,N_24813,N_24817);
nor UO_590 (O_590,N_24971,N_24982);
and UO_591 (O_591,N_24975,N_24937);
xor UO_592 (O_592,N_24994,N_24822);
and UO_593 (O_593,N_24948,N_24839);
and UO_594 (O_594,N_24992,N_24811);
and UO_595 (O_595,N_24969,N_24831);
nand UO_596 (O_596,N_24945,N_24881);
nor UO_597 (O_597,N_24819,N_24986);
or UO_598 (O_598,N_24933,N_24922);
and UO_599 (O_599,N_24979,N_24980);
or UO_600 (O_600,N_24891,N_24819);
nand UO_601 (O_601,N_24951,N_24886);
nand UO_602 (O_602,N_24814,N_24963);
or UO_603 (O_603,N_24880,N_24876);
nor UO_604 (O_604,N_24912,N_24847);
nand UO_605 (O_605,N_24975,N_24963);
nand UO_606 (O_606,N_24984,N_24959);
nand UO_607 (O_607,N_24832,N_24913);
nand UO_608 (O_608,N_24840,N_24920);
nand UO_609 (O_609,N_24894,N_24969);
nor UO_610 (O_610,N_24877,N_24978);
nand UO_611 (O_611,N_24921,N_24885);
and UO_612 (O_612,N_24947,N_24850);
xnor UO_613 (O_613,N_24894,N_24862);
xnor UO_614 (O_614,N_24932,N_24859);
nand UO_615 (O_615,N_24899,N_24894);
or UO_616 (O_616,N_24804,N_24963);
or UO_617 (O_617,N_24811,N_24945);
nand UO_618 (O_618,N_24916,N_24995);
and UO_619 (O_619,N_24981,N_24849);
or UO_620 (O_620,N_24879,N_24910);
nand UO_621 (O_621,N_24801,N_24919);
nand UO_622 (O_622,N_24957,N_24968);
and UO_623 (O_623,N_24971,N_24953);
nand UO_624 (O_624,N_24884,N_24898);
nor UO_625 (O_625,N_24823,N_24962);
xor UO_626 (O_626,N_24904,N_24926);
nand UO_627 (O_627,N_24802,N_24820);
or UO_628 (O_628,N_24972,N_24868);
and UO_629 (O_629,N_24836,N_24875);
nand UO_630 (O_630,N_24921,N_24871);
nor UO_631 (O_631,N_24930,N_24885);
nor UO_632 (O_632,N_24861,N_24820);
nand UO_633 (O_633,N_24901,N_24870);
nand UO_634 (O_634,N_24835,N_24917);
nor UO_635 (O_635,N_24847,N_24841);
or UO_636 (O_636,N_24814,N_24885);
nor UO_637 (O_637,N_24939,N_24947);
and UO_638 (O_638,N_24950,N_24962);
or UO_639 (O_639,N_24805,N_24847);
or UO_640 (O_640,N_24829,N_24935);
xnor UO_641 (O_641,N_24818,N_24911);
nand UO_642 (O_642,N_24955,N_24947);
xnor UO_643 (O_643,N_24853,N_24856);
or UO_644 (O_644,N_24978,N_24825);
nand UO_645 (O_645,N_24818,N_24906);
and UO_646 (O_646,N_24855,N_24999);
nor UO_647 (O_647,N_24986,N_24955);
xor UO_648 (O_648,N_24947,N_24862);
xor UO_649 (O_649,N_24993,N_24830);
or UO_650 (O_650,N_24866,N_24870);
nor UO_651 (O_651,N_24855,N_24962);
nand UO_652 (O_652,N_24875,N_24864);
xnor UO_653 (O_653,N_24984,N_24882);
or UO_654 (O_654,N_24868,N_24816);
and UO_655 (O_655,N_24861,N_24884);
or UO_656 (O_656,N_24964,N_24959);
xnor UO_657 (O_657,N_24910,N_24832);
nor UO_658 (O_658,N_24981,N_24921);
nor UO_659 (O_659,N_24833,N_24810);
or UO_660 (O_660,N_24902,N_24996);
nor UO_661 (O_661,N_24937,N_24994);
or UO_662 (O_662,N_24910,N_24853);
and UO_663 (O_663,N_24977,N_24841);
and UO_664 (O_664,N_24811,N_24920);
xnor UO_665 (O_665,N_24938,N_24993);
and UO_666 (O_666,N_24917,N_24923);
or UO_667 (O_667,N_24967,N_24853);
xor UO_668 (O_668,N_24889,N_24998);
nor UO_669 (O_669,N_24951,N_24991);
and UO_670 (O_670,N_24833,N_24895);
and UO_671 (O_671,N_24944,N_24913);
and UO_672 (O_672,N_24967,N_24818);
nor UO_673 (O_673,N_24844,N_24955);
nand UO_674 (O_674,N_24984,N_24980);
xor UO_675 (O_675,N_24928,N_24934);
xnor UO_676 (O_676,N_24813,N_24856);
or UO_677 (O_677,N_24904,N_24804);
or UO_678 (O_678,N_24834,N_24992);
xnor UO_679 (O_679,N_24802,N_24801);
nor UO_680 (O_680,N_24895,N_24912);
and UO_681 (O_681,N_24923,N_24952);
or UO_682 (O_682,N_24970,N_24900);
nand UO_683 (O_683,N_24942,N_24969);
or UO_684 (O_684,N_24865,N_24952);
xnor UO_685 (O_685,N_24846,N_24990);
nor UO_686 (O_686,N_24890,N_24864);
nor UO_687 (O_687,N_24813,N_24849);
or UO_688 (O_688,N_24900,N_24830);
nor UO_689 (O_689,N_24936,N_24811);
xor UO_690 (O_690,N_24818,N_24853);
nor UO_691 (O_691,N_24923,N_24986);
and UO_692 (O_692,N_24809,N_24811);
nor UO_693 (O_693,N_24927,N_24871);
and UO_694 (O_694,N_24963,N_24980);
and UO_695 (O_695,N_24890,N_24872);
nand UO_696 (O_696,N_24908,N_24892);
xor UO_697 (O_697,N_24827,N_24891);
or UO_698 (O_698,N_24879,N_24869);
nor UO_699 (O_699,N_24911,N_24965);
xor UO_700 (O_700,N_24933,N_24930);
xnor UO_701 (O_701,N_24947,N_24872);
xor UO_702 (O_702,N_24934,N_24880);
nor UO_703 (O_703,N_24949,N_24925);
and UO_704 (O_704,N_24880,N_24823);
xnor UO_705 (O_705,N_24947,N_24856);
or UO_706 (O_706,N_24801,N_24935);
or UO_707 (O_707,N_24981,N_24957);
or UO_708 (O_708,N_24869,N_24867);
nand UO_709 (O_709,N_24851,N_24975);
nor UO_710 (O_710,N_24840,N_24820);
and UO_711 (O_711,N_24859,N_24959);
and UO_712 (O_712,N_24906,N_24922);
nor UO_713 (O_713,N_24832,N_24849);
and UO_714 (O_714,N_24883,N_24838);
or UO_715 (O_715,N_24879,N_24903);
and UO_716 (O_716,N_24973,N_24968);
or UO_717 (O_717,N_24870,N_24902);
xnor UO_718 (O_718,N_24978,N_24984);
or UO_719 (O_719,N_24876,N_24889);
or UO_720 (O_720,N_24975,N_24979);
or UO_721 (O_721,N_24975,N_24879);
nor UO_722 (O_722,N_24817,N_24894);
or UO_723 (O_723,N_24971,N_24833);
nand UO_724 (O_724,N_24803,N_24851);
and UO_725 (O_725,N_24981,N_24942);
and UO_726 (O_726,N_24965,N_24842);
nor UO_727 (O_727,N_24931,N_24988);
xor UO_728 (O_728,N_24940,N_24997);
and UO_729 (O_729,N_24980,N_24892);
nor UO_730 (O_730,N_24865,N_24825);
nand UO_731 (O_731,N_24912,N_24810);
nor UO_732 (O_732,N_24993,N_24910);
and UO_733 (O_733,N_24837,N_24972);
xor UO_734 (O_734,N_24977,N_24836);
xor UO_735 (O_735,N_24938,N_24840);
xnor UO_736 (O_736,N_24832,N_24968);
nor UO_737 (O_737,N_24862,N_24892);
and UO_738 (O_738,N_24991,N_24826);
or UO_739 (O_739,N_24945,N_24872);
nor UO_740 (O_740,N_24947,N_24940);
xor UO_741 (O_741,N_24858,N_24868);
xor UO_742 (O_742,N_24988,N_24942);
and UO_743 (O_743,N_24909,N_24939);
and UO_744 (O_744,N_24969,N_24913);
nand UO_745 (O_745,N_24861,N_24925);
nand UO_746 (O_746,N_24989,N_24812);
nand UO_747 (O_747,N_24821,N_24843);
nor UO_748 (O_748,N_24865,N_24939);
nand UO_749 (O_749,N_24847,N_24823);
and UO_750 (O_750,N_24986,N_24827);
or UO_751 (O_751,N_24986,N_24990);
and UO_752 (O_752,N_24913,N_24884);
or UO_753 (O_753,N_24840,N_24937);
or UO_754 (O_754,N_24870,N_24816);
nor UO_755 (O_755,N_24990,N_24932);
or UO_756 (O_756,N_24928,N_24910);
and UO_757 (O_757,N_24839,N_24985);
nand UO_758 (O_758,N_24901,N_24951);
or UO_759 (O_759,N_24897,N_24874);
nor UO_760 (O_760,N_24810,N_24883);
xor UO_761 (O_761,N_24876,N_24845);
or UO_762 (O_762,N_24803,N_24895);
nand UO_763 (O_763,N_24823,N_24914);
nand UO_764 (O_764,N_24851,N_24933);
xnor UO_765 (O_765,N_24812,N_24815);
nand UO_766 (O_766,N_24848,N_24952);
nand UO_767 (O_767,N_24809,N_24952);
xor UO_768 (O_768,N_24954,N_24956);
nor UO_769 (O_769,N_24916,N_24953);
or UO_770 (O_770,N_24880,N_24962);
or UO_771 (O_771,N_24852,N_24880);
and UO_772 (O_772,N_24811,N_24937);
xnor UO_773 (O_773,N_24888,N_24812);
nor UO_774 (O_774,N_24977,N_24972);
nand UO_775 (O_775,N_24930,N_24962);
or UO_776 (O_776,N_24998,N_24823);
and UO_777 (O_777,N_24987,N_24899);
or UO_778 (O_778,N_24844,N_24972);
xnor UO_779 (O_779,N_24813,N_24882);
nor UO_780 (O_780,N_24969,N_24839);
nor UO_781 (O_781,N_24818,N_24811);
and UO_782 (O_782,N_24899,N_24922);
xnor UO_783 (O_783,N_24994,N_24905);
nor UO_784 (O_784,N_24928,N_24867);
xnor UO_785 (O_785,N_24908,N_24934);
xor UO_786 (O_786,N_24842,N_24819);
or UO_787 (O_787,N_24984,N_24853);
nand UO_788 (O_788,N_24925,N_24808);
or UO_789 (O_789,N_24816,N_24867);
xnor UO_790 (O_790,N_24818,N_24886);
xor UO_791 (O_791,N_24924,N_24941);
or UO_792 (O_792,N_24982,N_24978);
xor UO_793 (O_793,N_24912,N_24909);
and UO_794 (O_794,N_24809,N_24859);
xnor UO_795 (O_795,N_24924,N_24852);
nand UO_796 (O_796,N_24977,N_24856);
or UO_797 (O_797,N_24858,N_24972);
xnor UO_798 (O_798,N_24911,N_24876);
and UO_799 (O_799,N_24877,N_24916);
nand UO_800 (O_800,N_24972,N_24876);
xnor UO_801 (O_801,N_24827,N_24996);
xnor UO_802 (O_802,N_24973,N_24919);
nor UO_803 (O_803,N_24897,N_24811);
nor UO_804 (O_804,N_24879,N_24970);
or UO_805 (O_805,N_24946,N_24807);
xnor UO_806 (O_806,N_24933,N_24902);
nand UO_807 (O_807,N_24963,N_24909);
or UO_808 (O_808,N_24909,N_24997);
or UO_809 (O_809,N_24838,N_24810);
nand UO_810 (O_810,N_24877,N_24997);
or UO_811 (O_811,N_24899,N_24825);
nor UO_812 (O_812,N_24964,N_24887);
and UO_813 (O_813,N_24804,N_24805);
nand UO_814 (O_814,N_24817,N_24892);
nand UO_815 (O_815,N_24934,N_24990);
nor UO_816 (O_816,N_24964,N_24985);
nand UO_817 (O_817,N_24976,N_24868);
and UO_818 (O_818,N_24897,N_24908);
nor UO_819 (O_819,N_24842,N_24868);
nand UO_820 (O_820,N_24972,N_24942);
nor UO_821 (O_821,N_24851,N_24829);
nand UO_822 (O_822,N_24836,N_24960);
nor UO_823 (O_823,N_24909,N_24870);
or UO_824 (O_824,N_24804,N_24932);
or UO_825 (O_825,N_24836,N_24984);
nor UO_826 (O_826,N_24964,N_24855);
nand UO_827 (O_827,N_24994,N_24802);
nor UO_828 (O_828,N_24997,N_24933);
nor UO_829 (O_829,N_24924,N_24829);
nor UO_830 (O_830,N_24875,N_24896);
and UO_831 (O_831,N_24970,N_24801);
and UO_832 (O_832,N_24926,N_24921);
or UO_833 (O_833,N_24962,N_24960);
or UO_834 (O_834,N_24908,N_24858);
or UO_835 (O_835,N_24906,N_24953);
nand UO_836 (O_836,N_24980,N_24928);
nor UO_837 (O_837,N_24890,N_24976);
nor UO_838 (O_838,N_24882,N_24866);
nand UO_839 (O_839,N_24824,N_24878);
nand UO_840 (O_840,N_24887,N_24851);
xor UO_841 (O_841,N_24931,N_24951);
or UO_842 (O_842,N_24843,N_24860);
or UO_843 (O_843,N_24824,N_24812);
and UO_844 (O_844,N_24911,N_24902);
nand UO_845 (O_845,N_24859,N_24941);
or UO_846 (O_846,N_24809,N_24931);
nor UO_847 (O_847,N_24925,N_24905);
or UO_848 (O_848,N_24967,N_24946);
and UO_849 (O_849,N_24962,N_24969);
xor UO_850 (O_850,N_24992,N_24927);
nand UO_851 (O_851,N_24876,N_24844);
nor UO_852 (O_852,N_24933,N_24908);
and UO_853 (O_853,N_24806,N_24879);
and UO_854 (O_854,N_24984,N_24919);
nor UO_855 (O_855,N_24902,N_24884);
nand UO_856 (O_856,N_24868,N_24869);
xnor UO_857 (O_857,N_24864,N_24897);
or UO_858 (O_858,N_24894,N_24936);
and UO_859 (O_859,N_24948,N_24902);
xnor UO_860 (O_860,N_24890,N_24917);
xor UO_861 (O_861,N_24961,N_24923);
nor UO_862 (O_862,N_24923,N_24896);
nand UO_863 (O_863,N_24902,N_24859);
nand UO_864 (O_864,N_24916,N_24859);
nor UO_865 (O_865,N_24939,N_24836);
and UO_866 (O_866,N_24932,N_24976);
and UO_867 (O_867,N_24945,N_24882);
or UO_868 (O_868,N_24954,N_24976);
and UO_869 (O_869,N_24892,N_24984);
and UO_870 (O_870,N_24953,N_24904);
xnor UO_871 (O_871,N_24926,N_24923);
nand UO_872 (O_872,N_24923,N_24808);
or UO_873 (O_873,N_24857,N_24884);
or UO_874 (O_874,N_24811,N_24828);
nor UO_875 (O_875,N_24988,N_24857);
xnor UO_876 (O_876,N_24911,N_24923);
nand UO_877 (O_877,N_24945,N_24981);
or UO_878 (O_878,N_24977,N_24823);
or UO_879 (O_879,N_24806,N_24881);
and UO_880 (O_880,N_24848,N_24843);
nand UO_881 (O_881,N_24888,N_24892);
and UO_882 (O_882,N_24968,N_24924);
nand UO_883 (O_883,N_24923,N_24884);
xor UO_884 (O_884,N_24854,N_24983);
or UO_885 (O_885,N_24915,N_24983);
and UO_886 (O_886,N_24818,N_24979);
or UO_887 (O_887,N_24916,N_24963);
xnor UO_888 (O_888,N_24853,N_24974);
and UO_889 (O_889,N_24906,N_24900);
and UO_890 (O_890,N_24957,N_24840);
and UO_891 (O_891,N_24945,N_24934);
nor UO_892 (O_892,N_24803,N_24806);
and UO_893 (O_893,N_24944,N_24892);
xor UO_894 (O_894,N_24860,N_24917);
or UO_895 (O_895,N_24948,N_24822);
xnor UO_896 (O_896,N_24895,N_24911);
nand UO_897 (O_897,N_24955,N_24870);
xor UO_898 (O_898,N_24822,N_24843);
nand UO_899 (O_899,N_24944,N_24999);
and UO_900 (O_900,N_24823,N_24889);
or UO_901 (O_901,N_24901,N_24800);
nor UO_902 (O_902,N_24861,N_24924);
nor UO_903 (O_903,N_24880,N_24845);
or UO_904 (O_904,N_24995,N_24896);
xnor UO_905 (O_905,N_24907,N_24888);
nor UO_906 (O_906,N_24971,N_24834);
nand UO_907 (O_907,N_24912,N_24977);
or UO_908 (O_908,N_24895,N_24850);
or UO_909 (O_909,N_24837,N_24977);
and UO_910 (O_910,N_24848,N_24908);
nand UO_911 (O_911,N_24950,N_24944);
nand UO_912 (O_912,N_24807,N_24966);
xnor UO_913 (O_913,N_24973,N_24902);
and UO_914 (O_914,N_24903,N_24957);
or UO_915 (O_915,N_24835,N_24964);
nand UO_916 (O_916,N_24961,N_24920);
nand UO_917 (O_917,N_24955,N_24893);
xor UO_918 (O_918,N_24919,N_24825);
nand UO_919 (O_919,N_24931,N_24890);
nor UO_920 (O_920,N_24802,N_24997);
nor UO_921 (O_921,N_24857,N_24838);
and UO_922 (O_922,N_24965,N_24891);
or UO_923 (O_923,N_24931,N_24969);
xor UO_924 (O_924,N_24885,N_24950);
and UO_925 (O_925,N_24937,N_24843);
and UO_926 (O_926,N_24979,N_24985);
or UO_927 (O_927,N_24929,N_24927);
nand UO_928 (O_928,N_24802,N_24810);
or UO_929 (O_929,N_24942,N_24817);
or UO_930 (O_930,N_24868,N_24864);
or UO_931 (O_931,N_24903,N_24808);
and UO_932 (O_932,N_24985,N_24977);
and UO_933 (O_933,N_24901,N_24881);
and UO_934 (O_934,N_24918,N_24973);
nor UO_935 (O_935,N_24979,N_24808);
nand UO_936 (O_936,N_24877,N_24876);
or UO_937 (O_937,N_24930,N_24918);
xor UO_938 (O_938,N_24998,N_24844);
nand UO_939 (O_939,N_24906,N_24902);
xor UO_940 (O_940,N_24892,N_24921);
and UO_941 (O_941,N_24974,N_24972);
and UO_942 (O_942,N_24866,N_24885);
and UO_943 (O_943,N_24949,N_24897);
nand UO_944 (O_944,N_24923,N_24800);
or UO_945 (O_945,N_24983,N_24893);
or UO_946 (O_946,N_24806,N_24906);
nand UO_947 (O_947,N_24986,N_24861);
and UO_948 (O_948,N_24945,N_24839);
or UO_949 (O_949,N_24837,N_24801);
or UO_950 (O_950,N_24849,N_24823);
nor UO_951 (O_951,N_24866,N_24998);
nand UO_952 (O_952,N_24845,N_24965);
xnor UO_953 (O_953,N_24955,N_24882);
nand UO_954 (O_954,N_24956,N_24934);
and UO_955 (O_955,N_24962,N_24914);
or UO_956 (O_956,N_24876,N_24823);
or UO_957 (O_957,N_24871,N_24961);
nor UO_958 (O_958,N_24877,N_24938);
nand UO_959 (O_959,N_24923,N_24858);
or UO_960 (O_960,N_24812,N_24956);
nand UO_961 (O_961,N_24865,N_24944);
and UO_962 (O_962,N_24806,N_24825);
or UO_963 (O_963,N_24989,N_24840);
nand UO_964 (O_964,N_24852,N_24863);
xor UO_965 (O_965,N_24917,N_24925);
and UO_966 (O_966,N_24809,N_24933);
nor UO_967 (O_967,N_24995,N_24839);
nor UO_968 (O_968,N_24843,N_24839);
nand UO_969 (O_969,N_24982,N_24920);
nand UO_970 (O_970,N_24948,N_24845);
xor UO_971 (O_971,N_24849,N_24892);
xor UO_972 (O_972,N_24863,N_24812);
nor UO_973 (O_973,N_24868,N_24899);
xnor UO_974 (O_974,N_24848,N_24906);
nand UO_975 (O_975,N_24916,N_24973);
nor UO_976 (O_976,N_24866,N_24964);
xor UO_977 (O_977,N_24982,N_24910);
or UO_978 (O_978,N_24858,N_24873);
xor UO_979 (O_979,N_24929,N_24839);
nand UO_980 (O_980,N_24879,N_24871);
or UO_981 (O_981,N_24958,N_24803);
nand UO_982 (O_982,N_24804,N_24840);
or UO_983 (O_983,N_24824,N_24938);
or UO_984 (O_984,N_24925,N_24869);
or UO_985 (O_985,N_24973,N_24847);
nand UO_986 (O_986,N_24934,N_24868);
or UO_987 (O_987,N_24900,N_24976);
and UO_988 (O_988,N_24957,N_24930);
nor UO_989 (O_989,N_24956,N_24967);
and UO_990 (O_990,N_24898,N_24955);
nor UO_991 (O_991,N_24866,N_24933);
xor UO_992 (O_992,N_24950,N_24945);
nor UO_993 (O_993,N_24821,N_24901);
xnor UO_994 (O_994,N_24946,N_24977);
or UO_995 (O_995,N_24857,N_24902);
xnor UO_996 (O_996,N_24927,N_24990);
nand UO_997 (O_997,N_24855,N_24914);
nand UO_998 (O_998,N_24971,N_24842);
xnor UO_999 (O_999,N_24945,N_24812);
nand UO_1000 (O_1000,N_24870,N_24988);
or UO_1001 (O_1001,N_24997,N_24948);
nor UO_1002 (O_1002,N_24843,N_24945);
nor UO_1003 (O_1003,N_24991,N_24929);
nor UO_1004 (O_1004,N_24833,N_24855);
nor UO_1005 (O_1005,N_24873,N_24921);
xor UO_1006 (O_1006,N_24850,N_24877);
nor UO_1007 (O_1007,N_24830,N_24879);
nand UO_1008 (O_1008,N_24996,N_24975);
nor UO_1009 (O_1009,N_24869,N_24900);
xnor UO_1010 (O_1010,N_24976,N_24822);
xor UO_1011 (O_1011,N_24806,N_24988);
and UO_1012 (O_1012,N_24972,N_24955);
nand UO_1013 (O_1013,N_24899,N_24915);
or UO_1014 (O_1014,N_24889,N_24985);
or UO_1015 (O_1015,N_24846,N_24926);
nand UO_1016 (O_1016,N_24803,N_24983);
nand UO_1017 (O_1017,N_24927,N_24832);
nand UO_1018 (O_1018,N_24821,N_24952);
or UO_1019 (O_1019,N_24800,N_24908);
xor UO_1020 (O_1020,N_24870,N_24970);
and UO_1021 (O_1021,N_24878,N_24800);
or UO_1022 (O_1022,N_24859,N_24849);
nand UO_1023 (O_1023,N_24965,N_24949);
and UO_1024 (O_1024,N_24888,N_24891);
nand UO_1025 (O_1025,N_24825,N_24812);
or UO_1026 (O_1026,N_24945,N_24887);
and UO_1027 (O_1027,N_24961,N_24841);
nand UO_1028 (O_1028,N_24872,N_24978);
or UO_1029 (O_1029,N_24881,N_24987);
xnor UO_1030 (O_1030,N_24969,N_24836);
and UO_1031 (O_1031,N_24832,N_24973);
nand UO_1032 (O_1032,N_24800,N_24954);
or UO_1033 (O_1033,N_24833,N_24842);
nor UO_1034 (O_1034,N_24920,N_24964);
or UO_1035 (O_1035,N_24834,N_24898);
nand UO_1036 (O_1036,N_24984,N_24832);
xnor UO_1037 (O_1037,N_24988,N_24813);
and UO_1038 (O_1038,N_24871,N_24884);
and UO_1039 (O_1039,N_24805,N_24893);
nor UO_1040 (O_1040,N_24861,N_24949);
and UO_1041 (O_1041,N_24950,N_24861);
nand UO_1042 (O_1042,N_24804,N_24957);
and UO_1043 (O_1043,N_24946,N_24877);
or UO_1044 (O_1044,N_24898,N_24886);
or UO_1045 (O_1045,N_24880,N_24984);
xor UO_1046 (O_1046,N_24981,N_24854);
and UO_1047 (O_1047,N_24838,N_24917);
nor UO_1048 (O_1048,N_24848,N_24969);
nand UO_1049 (O_1049,N_24852,N_24957);
nand UO_1050 (O_1050,N_24821,N_24935);
xnor UO_1051 (O_1051,N_24825,N_24828);
or UO_1052 (O_1052,N_24943,N_24834);
or UO_1053 (O_1053,N_24897,N_24872);
nand UO_1054 (O_1054,N_24919,N_24923);
xnor UO_1055 (O_1055,N_24887,N_24957);
nor UO_1056 (O_1056,N_24856,N_24859);
xnor UO_1057 (O_1057,N_24857,N_24877);
and UO_1058 (O_1058,N_24859,N_24890);
or UO_1059 (O_1059,N_24933,N_24833);
nor UO_1060 (O_1060,N_24974,N_24823);
xor UO_1061 (O_1061,N_24971,N_24802);
nand UO_1062 (O_1062,N_24983,N_24903);
xnor UO_1063 (O_1063,N_24989,N_24923);
or UO_1064 (O_1064,N_24956,N_24882);
xnor UO_1065 (O_1065,N_24991,N_24987);
nor UO_1066 (O_1066,N_24806,N_24949);
and UO_1067 (O_1067,N_24812,N_24879);
nor UO_1068 (O_1068,N_24896,N_24846);
xor UO_1069 (O_1069,N_24895,N_24890);
nor UO_1070 (O_1070,N_24886,N_24968);
and UO_1071 (O_1071,N_24884,N_24905);
xnor UO_1072 (O_1072,N_24867,N_24926);
xor UO_1073 (O_1073,N_24987,N_24821);
xnor UO_1074 (O_1074,N_24974,N_24818);
or UO_1075 (O_1075,N_24967,N_24917);
nor UO_1076 (O_1076,N_24961,N_24873);
nor UO_1077 (O_1077,N_24954,N_24929);
xor UO_1078 (O_1078,N_24803,N_24960);
and UO_1079 (O_1079,N_24919,N_24998);
nand UO_1080 (O_1080,N_24928,N_24890);
and UO_1081 (O_1081,N_24942,N_24864);
nand UO_1082 (O_1082,N_24856,N_24952);
or UO_1083 (O_1083,N_24838,N_24881);
or UO_1084 (O_1084,N_24823,N_24856);
nor UO_1085 (O_1085,N_24983,N_24808);
nand UO_1086 (O_1086,N_24841,N_24987);
or UO_1087 (O_1087,N_24944,N_24929);
or UO_1088 (O_1088,N_24951,N_24918);
nand UO_1089 (O_1089,N_24860,N_24911);
or UO_1090 (O_1090,N_24915,N_24804);
or UO_1091 (O_1091,N_24934,N_24916);
or UO_1092 (O_1092,N_24886,N_24858);
nor UO_1093 (O_1093,N_24828,N_24930);
and UO_1094 (O_1094,N_24909,N_24861);
nor UO_1095 (O_1095,N_24996,N_24891);
or UO_1096 (O_1096,N_24805,N_24977);
nand UO_1097 (O_1097,N_24984,N_24823);
and UO_1098 (O_1098,N_24980,N_24821);
xor UO_1099 (O_1099,N_24985,N_24969);
xor UO_1100 (O_1100,N_24869,N_24871);
nand UO_1101 (O_1101,N_24961,N_24830);
xnor UO_1102 (O_1102,N_24879,N_24883);
and UO_1103 (O_1103,N_24838,N_24960);
nand UO_1104 (O_1104,N_24890,N_24955);
xnor UO_1105 (O_1105,N_24896,N_24812);
xnor UO_1106 (O_1106,N_24817,N_24837);
or UO_1107 (O_1107,N_24937,N_24866);
and UO_1108 (O_1108,N_24844,N_24908);
or UO_1109 (O_1109,N_24841,N_24898);
nor UO_1110 (O_1110,N_24803,N_24957);
nor UO_1111 (O_1111,N_24826,N_24879);
and UO_1112 (O_1112,N_24962,N_24994);
xor UO_1113 (O_1113,N_24835,N_24958);
nor UO_1114 (O_1114,N_24883,N_24935);
and UO_1115 (O_1115,N_24909,N_24886);
and UO_1116 (O_1116,N_24873,N_24943);
xnor UO_1117 (O_1117,N_24914,N_24906);
nor UO_1118 (O_1118,N_24993,N_24928);
xor UO_1119 (O_1119,N_24953,N_24972);
nand UO_1120 (O_1120,N_24874,N_24887);
nand UO_1121 (O_1121,N_24816,N_24979);
nor UO_1122 (O_1122,N_24866,N_24856);
nand UO_1123 (O_1123,N_24802,N_24846);
or UO_1124 (O_1124,N_24933,N_24856);
nor UO_1125 (O_1125,N_24883,N_24964);
or UO_1126 (O_1126,N_24942,N_24810);
xnor UO_1127 (O_1127,N_24855,N_24953);
xnor UO_1128 (O_1128,N_24918,N_24819);
nor UO_1129 (O_1129,N_24939,N_24979);
nand UO_1130 (O_1130,N_24970,N_24873);
xnor UO_1131 (O_1131,N_24809,N_24930);
nor UO_1132 (O_1132,N_24876,N_24917);
and UO_1133 (O_1133,N_24908,N_24949);
nand UO_1134 (O_1134,N_24874,N_24917);
nand UO_1135 (O_1135,N_24814,N_24864);
or UO_1136 (O_1136,N_24975,N_24899);
xor UO_1137 (O_1137,N_24923,N_24904);
xor UO_1138 (O_1138,N_24829,N_24910);
nand UO_1139 (O_1139,N_24947,N_24892);
or UO_1140 (O_1140,N_24813,N_24922);
nand UO_1141 (O_1141,N_24968,N_24861);
nand UO_1142 (O_1142,N_24802,N_24959);
nand UO_1143 (O_1143,N_24988,N_24833);
nor UO_1144 (O_1144,N_24941,N_24880);
and UO_1145 (O_1145,N_24844,N_24801);
nor UO_1146 (O_1146,N_24873,N_24854);
nand UO_1147 (O_1147,N_24920,N_24882);
nand UO_1148 (O_1148,N_24911,N_24913);
nor UO_1149 (O_1149,N_24901,N_24840);
xor UO_1150 (O_1150,N_24882,N_24907);
nand UO_1151 (O_1151,N_24950,N_24948);
or UO_1152 (O_1152,N_24810,N_24878);
xnor UO_1153 (O_1153,N_24867,N_24968);
or UO_1154 (O_1154,N_24825,N_24962);
and UO_1155 (O_1155,N_24915,N_24815);
xor UO_1156 (O_1156,N_24846,N_24847);
and UO_1157 (O_1157,N_24937,N_24833);
and UO_1158 (O_1158,N_24831,N_24835);
and UO_1159 (O_1159,N_24892,N_24902);
and UO_1160 (O_1160,N_24859,N_24982);
or UO_1161 (O_1161,N_24891,N_24948);
or UO_1162 (O_1162,N_24995,N_24836);
nand UO_1163 (O_1163,N_24835,N_24869);
xor UO_1164 (O_1164,N_24804,N_24833);
and UO_1165 (O_1165,N_24977,N_24920);
or UO_1166 (O_1166,N_24975,N_24925);
xnor UO_1167 (O_1167,N_24935,N_24967);
nor UO_1168 (O_1168,N_24896,N_24956);
and UO_1169 (O_1169,N_24974,N_24828);
or UO_1170 (O_1170,N_24905,N_24954);
nand UO_1171 (O_1171,N_24930,N_24897);
nand UO_1172 (O_1172,N_24967,N_24997);
or UO_1173 (O_1173,N_24828,N_24847);
xnor UO_1174 (O_1174,N_24839,N_24916);
and UO_1175 (O_1175,N_24814,N_24911);
nor UO_1176 (O_1176,N_24984,N_24986);
and UO_1177 (O_1177,N_24962,N_24956);
xnor UO_1178 (O_1178,N_24969,N_24886);
and UO_1179 (O_1179,N_24887,N_24856);
and UO_1180 (O_1180,N_24851,N_24892);
or UO_1181 (O_1181,N_24988,N_24981);
and UO_1182 (O_1182,N_24952,N_24887);
and UO_1183 (O_1183,N_24975,N_24945);
nor UO_1184 (O_1184,N_24875,N_24921);
nand UO_1185 (O_1185,N_24917,N_24957);
or UO_1186 (O_1186,N_24805,N_24960);
or UO_1187 (O_1187,N_24943,N_24888);
and UO_1188 (O_1188,N_24888,N_24868);
xnor UO_1189 (O_1189,N_24936,N_24838);
xnor UO_1190 (O_1190,N_24969,N_24832);
xnor UO_1191 (O_1191,N_24843,N_24970);
and UO_1192 (O_1192,N_24974,N_24888);
nand UO_1193 (O_1193,N_24926,N_24939);
nor UO_1194 (O_1194,N_24959,N_24978);
and UO_1195 (O_1195,N_24833,N_24897);
or UO_1196 (O_1196,N_24949,N_24870);
and UO_1197 (O_1197,N_24874,N_24830);
nor UO_1198 (O_1198,N_24992,N_24919);
xor UO_1199 (O_1199,N_24905,N_24893);
or UO_1200 (O_1200,N_24819,N_24866);
nand UO_1201 (O_1201,N_24991,N_24961);
and UO_1202 (O_1202,N_24941,N_24999);
xor UO_1203 (O_1203,N_24925,N_24980);
nand UO_1204 (O_1204,N_24853,N_24943);
nand UO_1205 (O_1205,N_24887,N_24965);
nand UO_1206 (O_1206,N_24955,N_24942);
and UO_1207 (O_1207,N_24909,N_24840);
and UO_1208 (O_1208,N_24902,N_24944);
and UO_1209 (O_1209,N_24913,N_24820);
nor UO_1210 (O_1210,N_24946,N_24956);
or UO_1211 (O_1211,N_24981,N_24826);
xnor UO_1212 (O_1212,N_24836,N_24991);
nand UO_1213 (O_1213,N_24828,N_24946);
nand UO_1214 (O_1214,N_24990,N_24837);
xnor UO_1215 (O_1215,N_24809,N_24969);
xor UO_1216 (O_1216,N_24936,N_24818);
nand UO_1217 (O_1217,N_24845,N_24954);
or UO_1218 (O_1218,N_24960,N_24801);
nand UO_1219 (O_1219,N_24836,N_24844);
and UO_1220 (O_1220,N_24859,N_24891);
or UO_1221 (O_1221,N_24842,N_24924);
or UO_1222 (O_1222,N_24811,N_24984);
or UO_1223 (O_1223,N_24983,N_24815);
nor UO_1224 (O_1224,N_24955,N_24938);
and UO_1225 (O_1225,N_24899,N_24824);
and UO_1226 (O_1226,N_24851,N_24852);
xnor UO_1227 (O_1227,N_24828,N_24954);
xnor UO_1228 (O_1228,N_24957,N_24940);
nand UO_1229 (O_1229,N_24810,N_24982);
nor UO_1230 (O_1230,N_24860,N_24985);
nand UO_1231 (O_1231,N_24974,N_24822);
nor UO_1232 (O_1232,N_24889,N_24987);
nor UO_1233 (O_1233,N_24853,N_24918);
xor UO_1234 (O_1234,N_24872,N_24850);
and UO_1235 (O_1235,N_24883,N_24928);
nor UO_1236 (O_1236,N_24921,N_24944);
nor UO_1237 (O_1237,N_24812,N_24912);
xnor UO_1238 (O_1238,N_24933,N_24981);
or UO_1239 (O_1239,N_24841,N_24844);
and UO_1240 (O_1240,N_24862,N_24801);
and UO_1241 (O_1241,N_24952,N_24857);
nand UO_1242 (O_1242,N_24969,N_24823);
and UO_1243 (O_1243,N_24881,N_24976);
or UO_1244 (O_1244,N_24960,N_24907);
or UO_1245 (O_1245,N_24937,N_24987);
xor UO_1246 (O_1246,N_24993,N_24949);
xnor UO_1247 (O_1247,N_24823,N_24858);
nor UO_1248 (O_1248,N_24801,N_24956);
nor UO_1249 (O_1249,N_24993,N_24978);
or UO_1250 (O_1250,N_24974,N_24986);
and UO_1251 (O_1251,N_24838,N_24907);
nor UO_1252 (O_1252,N_24953,N_24974);
or UO_1253 (O_1253,N_24826,N_24947);
or UO_1254 (O_1254,N_24870,N_24942);
nand UO_1255 (O_1255,N_24959,N_24905);
nand UO_1256 (O_1256,N_24967,N_24970);
nor UO_1257 (O_1257,N_24829,N_24964);
xnor UO_1258 (O_1258,N_24949,N_24956);
and UO_1259 (O_1259,N_24820,N_24849);
xnor UO_1260 (O_1260,N_24994,N_24963);
or UO_1261 (O_1261,N_24870,N_24913);
nor UO_1262 (O_1262,N_24808,N_24825);
or UO_1263 (O_1263,N_24829,N_24902);
and UO_1264 (O_1264,N_24893,N_24819);
nand UO_1265 (O_1265,N_24904,N_24928);
xnor UO_1266 (O_1266,N_24983,N_24961);
or UO_1267 (O_1267,N_24809,N_24830);
nand UO_1268 (O_1268,N_24956,N_24838);
or UO_1269 (O_1269,N_24958,N_24911);
and UO_1270 (O_1270,N_24976,N_24926);
and UO_1271 (O_1271,N_24838,N_24818);
xnor UO_1272 (O_1272,N_24940,N_24832);
nand UO_1273 (O_1273,N_24986,N_24806);
and UO_1274 (O_1274,N_24988,N_24895);
nor UO_1275 (O_1275,N_24907,N_24852);
nor UO_1276 (O_1276,N_24869,N_24895);
nand UO_1277 (O_1277,N_24983,N_24879);
nand UO_1278 (O_1278,N_24995,N_24917);
nand UO_1279 (O_1279,N_24810,N_24828);
nand UO_1280 (O_1280,N_24893,N_24888);
or UO_1281 (O_1281,N_24803,N_24926);
or UO_1282 (O_1282,N_24947,N_24810);
and UO_1283 (O_1283,N_24858,N_24891);
nor UO_1284 (O_1284,N_24952,N_24910);
nand UO_1285 (O_1285,N_24962,N_24924);
nor UO_1286 (O_1286,N_24885,N_24844);
nand UO_1287 (O_1287,N_24835,N_24969);
or UO_1288 (O_1288,N_24833,N_24993);
or UO_1289 (O_1289,N_24859,N_24892);
nand UO_1290 (O_1290,N_24836,N_24864);
xnor UO_1291 (O_1291,N_24980,N_24971);
xor UO_1292 (O_1292,N_24962,N_24944);
nor UO_1293 (O_1293,N_24933,N_24826);
nand UO_1294 (O_1294,N_24924,N_24815);
xnor UO_1295 (O_1295,N_24832,N_24837);
nand UO_1296 (O_1296,N_24843,N_24941);
and UO_1297 (O_1297,N_24980,N_24824);
and UO_1298 (O_1298,N_24818,N_24898);
and UO_1299 (O_1299,N_24805,N_24894);
xor UO_1300 (O_1300,N_24934,N_24857);
and UO_1301 (O_1301,N_24824,N_24978);
nand UO_1302 (O_1302,N_24942,N_24820);
and UO_1303 (O_1303,N_24829,N_24854);
xor UO_1304 (O_1304,N_24957,N_24904);
nand UO_1305 (O_1305,N_24931,N_24919);
or UO_1306 (O_1306,N_24995,N_24909);
nor UO_1307 (O_1307,N_24911,N_24903);
xor UO_1308 (O_1308,N_24972,N_24878);
and UO_1309 (O_1309,N_24943,N_24955);
nand UO_1310 (O_1310,N_24843,N_24993);
and UO_1311 (O_1311,N_24828,N_24949);
nand UO_1312 (O_1312,N_24814,N_24895);
nor UO_1313 (O_1313,N_24948,N_24869);
or UO_1314 (O_1314,N_24937,N_24855);
nand UO_1315 (O_1315,N_24888,N_24980);
xnor UO_1316 (O_1316,N_24926,N_24938);
nand UO_1317 (O_1317,N_24861,N_24911);
or UO_1318 (O_1318,N_24897,N_24824);
nor UO_1319 (O_1319,N_24837,N_24970);
nand UO_1320 (O_1320,N_24823,N_24888);
xnor UO_1321 (O_1321,N_24870,N_24804);
xor UO_1322 (O_1322,N_24855,N_24897);
and UO_1323 (O_1323,N_24935,N_24915);
or UO_1324 (O_1324,N_24856,N_24907);
xor UO_1325 (O_1325,N_24817,N_24832);
or UO_1326 (O_1326,N_24818,N_24861);
xnor UO_1327 (O_1327,N_24955,N_24855);
and UO_1328 (O_1328,N_24854,N_24986);
nor UO_1329 (O_1329,N_24863,N_24878);
nand UO_1330 (O_1330,N_24968,N_24928);
nor UO_1331 (O_1331,N_24948,N_24817);
xor UO_1332 (O_1332,N_24809,N_24977);
xor UO_1333 (O_1333,N_24942,N_24858);
xnor UO_1334 (O_1334,N_24844,N_24884);
nor UO_1335 (O_1335,N_24892,N_24874);
or UO_1336 (O_1336,N_24946,N_24840);
nor UO_1337 (O_1337,N_24935,N_24894);
xor UO_1338 (O_1338,N_24876,N_24841);
xor UO_1339 (O_1339,N_24932,N_24884);
nor UO_1340 (O_1340,N_24987,N_24940);
or UO_1341 (O_1341,N_24931,N_24859);
xor UO_1342 (O_1342,N_24976,N_24989);
and UO_1343 (O_1343,N_24857,N_24987);
nor UO_1344 (O_1344,N_24904,N_24981);
and UO_1345 (O_1345,N_24827,N_24911);
or UO_1346 (O_1346,N_24911,N_24893);
nor UO_1347 (O_1347,N_24800,N_24900);
and UO_1348 (O_1348,N_24872,N_24868);
nor UO_1349 (O_1349,N_24872,N_24919);
or UO_1350 (O_1350,N_24866,N_24852);
and UO_1351 (O_1351,N_24862,N_24904);
and UO_1352 (O_1352,N_24825,N_24987);
or UO_1353 (O_1353,N_24901,N_24898);
or UO_1354 (O_1354,N_24840,N_24954);
nor UO_1355 (O_1355,N_24986,N_24826);
xor UO_1356 (O_1356,N_24845,N_24999);
xor UO_1357 (O_1357,N_24803,N_24823);
nor UO_1358 (O_1358,N_24824,N_24834);
and UO_1359 (O_1359,N_24858,N_24845);
and UO_1360 (O_1360,N_24907,N_24869);
or UO_1361 (O_1361,N_24831,N_24830);
xor UO_1362 (O_1362,N_24991,N_24906);
nand UO_1363 (O_1363,N_24999,N_24968);
and UO_1364 (O_1364,N_24992,N_24831);
xnor UO_1365 (O_1365,N_24981,N_24916);
and UO_1366 (O_1366,N_24957,N_24869);
xnor UO_1367 (O_1367,N_24860,N_24926);
nor UO_1368 (O_1368,N_24856,N_24828);
and UO_1369 (O_1369,N_24897,N_24968);
or UO_1370 (O_1370,N_24941,N_24940);
or UO_1371 (O_1371,N_24811,N_24813);
or UO_1372 (O_1372,N_24993,N_24871);
nand UO_1373 (O_1373,N_24864,N_24820);
and UO_1374 (O_1374,N_24923,N_24928);
nand UO_1375 (O_1375,N_24985,N_24974);
nor UO_1376 (O_1376,N_24801,N_24950);
nand UO_1377 (O_1377,N_24829,N_24928);
and UO_1378 (O_1378,N_24986,N_24889);
and UO_1379 (O_1379,N_24843,N_24960);
and UO_1380 (O_1380,N_24800,N_24836);
or UO_1381 (O_1381,N_24804,N_24940);
xnor UO_1382 (O_1382,N_24946,N_24900);
xnor UO_1383 (O_1383,N_24961,N_24933);
or UO_1384 (O_1384,N_24894,N_24843);
xnor UO_1385 (O_1385,N_24960,N_24813);
and UO_1386 (O_1386,N_24961,N_24886);
nand UO_1387 (O_1387,N_24955,N_24916);
nand UO_1388 (O_1388,N_24905,N_24806);
nand UO_1389 (O_1389,N_24830,N_24848);
and UO_1390 (O_1390,N_24941,N_24865);
xor UO_1391 (O_1391,N_24874,N_24828);
nand UO_1392 (O_1392,N_24906,N_24801);
xor UO_1393 (O_1393,N_24844,N_24871);
or UO_1394 (O_1394,N_24893,N_24818);
nand UO_1395 (O_1395,N_24972,N_24909);
or UO_1396 (O_1396,N_24937,N_24923);
nor UO_1397 (O_1397,N_24936,N_24949);
nand UO_1398 (O_1398,N_24951,N_24957);
nor UO_1399 (O_1399,N_24801,N_24849);
or UO_1400 (O_1400,N_24879,N_24926);
or UO_1401 (O_1401,N_24993,N_24838);
xor UO_1402 (O_1402,N_24958,N_24817);
nor UO_1403 (O_1403,N_24948,N_24846);
nor UO_1404 (O_1404,N_24901,N_24910);
nand UO_1405 (O_1405,N_24836,N_24988);
or UO_1406 (O_1406,N_24990,N_24865);
and UO_1407 (O_1407,N_24991,N_24878);
xnor UO_1408 (O_1408,N_24981,N_24925);
nand UO_1409 (O_1409,N_24933,N_24819);
and UO_1410 (O_1410,N_24886,N_24948);
and UO_1411 (O_1411,N_24893,N_24866);
nor UO_1412 (O_1412,N_24845,N_24812);
and UO_1413 (O_1413,N_24868,N_24821);
or UO_1414 (O_1414,N_24943,N_24942);
and UO_1415 (O_1415,N_24974,N_24839);
nor UO_1416 (O_1416,N_24887,N_24873);
nand UO_1417 (O_1417,N_24889,N_24925);
nor UO_1418 (O_1418,N_24955,N_24853);
nand UO_1419 (O_1419,N_24909,N_24859);
nand UO_1420 (O_1420,N_24910,N_24994);
nand UO_1421 (O_1421,N_24832,N_24999);
xnor UO_1422 (O_1422,N_24885,N_24880);
xnor UO_1423 (O_1423,N_24868,N_24964);
or UO_1424 (O_1424,N_24963,N_24836);
nor UO_1425 (O_1425,N_24955,N_24878);
or UO_1426 (O_1426,N_24819,N_24875);
nand UO_1427 (O_1427,N_24876,N_24950);
xor UO_1428 (O_1428,N_24943,N_24805);
nand UO_1429 (O_1429,N_24858,N_24890);
xor UO_1430 (O_1430,N_24851,N_24909);
and UO_1431 (O_1431,N_24958,N_24959);
and UO_1432 (O_1432,N_24878,N_24852);
and UO_1433 (O_1433,N_24869,N_24963);
nor UO_1434 (O_1434,N_24857,N_24998);
and UO_1435 (O_1435,N_24829,N_24947);
nand UO_1436 (O_1436,N_24825,N_24844);
xnor UO_1437 (O_1437,N_24855,N_24907);
and UO_1438 (O_1438,N_24832,N_24953);
xor UO_1439 (O_1439,N_24989,N_24802);
and UO_1440 (O_1440,N_24817,N_24927);
or UO_1441 (O_1441,N_24915,N_24986);
or UO_1442 (O_1442,N_24961,N_24953);
and UO_1443 (O_1443,N_24983,N_24801);
xnor UO_1444 (O_1444,N_24969,N_24841);
nor UO_1445 (O_1445,N_24945,N_24880);
nor UO_1446 (O_1446,N_24972,N_24961);
or UO_1447 (O_1447,N_24949,N_24903);
xnor UO_1448 (O_1448,N_24879,N_24901);
nand UO_1449 (O_1449,N_24999,N_24816);
xor UO_1450 (O_1450,N_24952,N_24840);
nand UO_1451 (O_1451,N_24869,N_24844);
xor UO_1452 (O_1452,N_24859,N_24811);
nor UO_1453 (O_1453,N_24988,N_24959);
nand UO_1454 (O_1454,N_24988,N_24812);
and UO_1455 (O_1455,N_24861,N_24804);
and UO_1456 (O_1456,N_24996,N_24981);
and UO_1457 (O_1457,N_24966,N_24852);
nor UO_1458 (O_1458,N_24900,N_24873);
nand UO_1459 (O_1459,N_24978,N_24946);
or UO_1460 (O_1460,N_24877,N_24892);
xnor UO_1461 (O_1461,N_24993,N_24954);
and UO_1462 (O_1462,N_24981,N_24984);
nor UO_1463 (O_1463,N_24864,N_24956);
nand UO_1464 (O_1464,N_24848,N_24884);
and UO_1465 (O_1465,N_24968,N_24915);
or UO_1466 (O_1466,N_24817,N_24896);
nor UO_1467 (O_1467,N_24916,N_24937);
nand UO_1468 (O_1468,N_24995,N_24849);
and UO_1469 (O_1469,N_24976,N_24927);
and UO_1470 (O_1470,N_24951,N_24820);
or UO_1471 (O_1471,N_24939,N_24995);
nor UO_1472 (O_1472,N_24893,N_24986);
and UO_1473 (O_1473,N_24966,N_24874);
and UO_1474 (O_1474,N_24801,N_24843);
and UO_1475 (O_1475,N_24871,N_24880);
nand UO_1476 (O_1476,N_24833,N_24968);
nor UO_1477 (O_1477,N_24845,N_24873);
nor UO_1478 (O_1478,N_24901,N_24926);
or UO_1479 (O_1479,N_24838,N_24919);
and UO_1480 (O_1480,N_24818,N_24953);
xor UO_1481 (O_1481,N_24806,N_24885);
nor UO_1482 (O_1482,N_24871,N_24975);
nor UO_1483 (O_1483,N_24814,N_24996);
nor UO_1484 (O_1484,N_24901,N_24920);
nand UO_1485 (O_1485,N_24903,N_24896);
nand UO_1486 (O_1486,N_24896,N_24873);
nand UO_1487 (O_1487,N_24962,N_24997);
xor UO_1488 (O_1488,N_24962,N_24826);
xnor UO_1489 (O_1489,N_24800,N_24966);
xor UO_1490 (O_1490,N_24891,N_24846);
nand UO_1491 (O_1491,N_24966,N_24850);
xor UO_1492 (O_1492,N_24806,N_24880);
nor UO_1493 (O_1493,N_24893,N_24870);
nand UO_1494 (O_1494,N_24899,N_24985);
xor UO_1495 (O_1495,N_24861,N_24830);
xnor UO_1496 (O_1496,N_24836,N_24898);
nor UO_1497 (O_1497,N_24918,N_24985);
xor UO_1498 (O_1498,N_24876,N_24920);
nor UO_1499 (O_1499,N_24952,N_24962);
or UO_1500 (O_1500,N_24946,N_24959);
or UO_1501 (O_1501,N_24958,N_24985);
xnor UO_1502 (O_1502,N_24996,N_24965);
nand UO_1503 (O_1503,N_24984,N_24833);
nor UO_1504 (O_1504,N_24977,N_24910);
nor UO_1505 (O_1505,N_24949,N_24973);
xor UO_1506 (O_1506,N_24832,N_24988);
or UO_1507 (O_1507,N_24978,N_24980);
nor UO_1508 (O_1508,N_24981,N_24803);
nand UO_1509 (O_1509,N_24891,N_24842);
or UO_1510 (O_1510,N_24986,N_24821);
or UO_1511 (O_1511,N_24891,N_24986);
and UO_1512 (O_1512,N_24805,N_24973);
xnor UO_1513 (O_1513,N_24924,N_24867);
nand UO_1514 (O_1514,N_24810,N_24831);
nand UO_1515 (O_1515,N_24975,N_24877);
nor UO_1516 (O_1516,N_24935,N_24833);
nor UO_1517 (O_1517,N_24958,N_24858);
nor UO_1518 (O_1518,N_24809,N_24807);
or UO_1519 (O_1519,N_24840,N_24843);
nor UO_1520 (O_1520,N_24903,N_24809);
or UO_1521 (O_1521,N_24959,N_24981);
nand UO_1522 (O_1522,N_24830,N_24878);
nor UO_1523 (O_1523,N_24928,N_24868);
xor UO_1524 (O_1524,N_24848,N_24821);
nand UO_1525 (O_1525,N_24823,N_24820);
or UO_1526 (O_1526,N_24804,N_24855);
nand UO_1527 (O_1527,N_24979,N_24912);
xor UO_1528 (O_1528,N_24946,N_24922);
and UO_1529 (O_1529,N_24947,N_24896);
nand UO_1530 (O_1530,N_24823,N_24859);
xor UO_1531 (O_1531,N_24802,N_24890);
xor UO_1532 (O_1532,N_24919,N_24990);
nor UO_1533 (O_1533,N_24962,N_24820);
or UO_1534 (O_1534,N_24955,N_24950);
and UO_1535 (O_1535,N_24930,N_24819);
nand UO_1536 (O_1536,N_24833,N_24805);
xor UO_1537 (O_1537,N_24838,N_24940);
nor UO_1538 (O_1538,N_24940,N_24835);
xor UO_1539 (O_1539,N_24994,N_24805);
nand UO_1540 (O_1540,N_24967,N_24941);
nand UO_1541 (O_1541,N_24824,N_24896);
and UO_1542 (O_1542,N_24969,N_24860);
nor UO_1543 (O_1543,N_24956,N_24885);
nand UO_1544 (O_1544,N_24827,N_24952);
nand UO_1545 (O_1545,N_24931,N_24865);
nand UO_1546 (O_1546,N_24873,N_24912);
or UO_1547 (O_1547,N_24912,N_24910);
xor UO_1548 (O_1548,N_24866,N_24876);
xnor UO_1549 (O_1549,N_24992,N_24913);
and UO_1550 (O_1550,N_24848,N_24873);
or UO_1551 (O_1551,N_24948,N_24862);
nor UO_1552 (O_1552,N_24917,N_24946);
nand UO_1553 (O_1553,N_24915,N_24832);
and UO_1554 (O_1554,N_24921,N_24977);
nand UO_1555 (O_1555,N_24825,N_24993);
nand UO_1556 (O_1556,N_24953,N_24884);
nand UO_1557 (O_1557,N_24840,N_24962);
nand UO_1558 (O_1558,N_24815,N_24948);
nand UO_1559 (O_1559,N_24945,N_24956);
xor UO_1560 (O_1560,N_24948,N_24802);
or UO_1561 (O_1561,N_24986,N_24914);
nor UO_1562 (O_1562,N_24889,N_24909);
or UO_1563 (O_1563,N_24808,N_24902);
xnor UO_1564 (O_1564,N_24882,N_24865);
or UO_1565 (O_1565,N_24974,N_24806);
nand UO_1566 (O_1566,N_24922,N_24861);
and UO_1567 (O_1567,N_24944,N_24946);
xnor UO_1568 (O_1568,N_24989,N_24846);
and UO_1569 (O_1569,N_24962,N_24957);
and UO_1570 (O_1570,N_24952,N_24942);
or UO_1571 (O_1571,N_24960,N_24950);
nand UO_1572 (O_1572,N_24845,N_24996);
nand UO_1573 (O_1573,N_24857,N_24999);
xor UO_1574 (O_1574,N_24909,N_24957);
nor UO_1575 (O_1575,N_24829,N_24804);
nand UO_1576 (O_1576,N_24975,N_24872);
nand UO_1577 (O_1577,N_24901,N_24963);
nor UO_1578 (O_1578,N_24932,N_24862);
nor UO_1579 (O_1579,N_24940,N_24939);
nor UO_1580 (O_1580,N_24985,N_24870);
or UO_1581 (O_1581,N_24902,N_24803);
or UO_1582 (O_1582,N_24993,N_24847);
nor UO_1583 (O_1583,N_24994,N_24839);
xor UO_1584 (O_1584,N_24935,N_24827);
or UO_1585 (O_1585,N_24816,N_24971);
or UO_1586 (O_1586,N_24990,N_24980);
nand UO_1587 (O_1587,N_24893,N_24875);
or UO_1588 (O_1588,N_24997,N_24924);
nor UO_1589 (O_1589,N_24903,N_24901);
nand UO_1590 (O_1590,N_24874,N_24834);
nand UO_1591 (O_1591,N_24801,N_24914);
nand UO_1592 (O_1592,N_24937,N_24821);
or UO_1593 (O_1593,N_24989,N_24905);
nand UO_1594 (O_1594,N_24893,N_24936);
or UO_1595 (O_1595,N_24970,N_24819);
xnor UO_1596 (O_1596,N_24957,N_24967);
nand UO_1597 (O_1597,N_24967,N_24888);
nor UO_1598 (O_1598,N_24841,N_24836);
nor UO_1599 (O_1599,N_24861,N_24851);
xor UO_1600 (O_1600,N_24936,N_24901);
nand UO_1601 (O_1601,N_24910,N_24824);
xnor UO_1602 (O_1602,N_24984,N_24995);
and UO_1603 (O_1603,N_24973,N_24886);
or UO_1604 (O_1604,N_24857,N_24852);
and UO_1605 (O_1605,N_24890,N_24847);
nand UO_1606 (O_1606,N_24820,N_24895);
nand UO_1607 (O_1607,N_24869,N_24946);
xnor UO_1608 (O_1608,N_24951,N_24851);
nor UO_1609 (O_1609,N_24949,N_24859);
nor UO_1610 (O_1610,N_24837,N_24877);
xnor UO_1611 (O_1611,N_24924,N_24870);
or UO_1612 (O_1612,N_24975,N_24954);
and UO_1613 (O_1613,N_24874,N_24981);
xor UO_1614 (O_1614,N_24892,N_24957);
nor UO_1615 (O_1615,N_24948,N_24974);
xnor UO_1616 (O_1616,N_24831,N_24806);
nand UO_1617 (O_1617,N_24926,N_24931);
and UO_1618 (O_1618,N_24900,N_24818);
or UO_1619 (O_1619,N_24933,N_24832);
or UO_1620 (O_1620,N_24831,N_24909);
or UO_1621 (O_1621,N_24897,N_24837);
nand UO_1622 (O_1622,N_24908,N_24974);
nand UO_1623 (O_1623,N_24801,N_24812);
nor UO_1624 (O_1624,N_24859,N_24991);
or UO_1625 (O_1625,N_24895,N_24839);
nor UO_1626 (O_1626,N_24809,N_24961);
nor UO_1627 (O_1627,N_24863,N_24876);
nor UO_1628 (O_1628,N_24982,N_24822);
xnor UO_1629 (O_1629,N_24857,N_24906);
nand UO_1630 (O_1630,N_24907,N_24993);
and UO_1631 (O_1631,N_24904,N_24814);
nand UO_1632 (O_1632,N_24935,N_24921);
and UO_1633 (O_1633,N_24851,N_24832);
nor UO_1634 (O_1634,N_24929,N_24937);
nor UO_1635 (O_1635,N_24969,N_24972);
nand UO_1636 (O_1636,N_24897,N_24878);
nor UO_1637 (O_1637,N_24860,N_24885);
xnor UO_1638 (O_1638,N_24853,N_24980);
nand UO_1639 (O_1639,N_24944,N_24854);
or UO_1640 (O_1640,N_24935,N_24900);
or UO_1641 (O_1641,N_24884,N_24931);
and UO_1642 (O_1642,N_24839,N_24850);
or UO_1643 (O_1643,N_24854,N_24927);
xnor UO_1644 (O_1644,N_24967,N_24975);
and UO_1645 (O_1645,N_24963,N_24827);
xor UO_1646 (O_1646,N_24955,N_24883);
or UO_1647 (O_1647,N_24915,N_24954);
xor UO_1648 (O_1648,N_24805,N_24832);
nand UO_1649 (O_1649,N_24972,N_24952);
xnor UO_1650 (O_1650,N_24934,N_24935);
xnor UO_1651 (O_1651,N_24951,N_24965);
or UO_1652 (O_1652,N_24825,N_24902);
or UO_1653 (O_1653,N_24952,N_24990);
and UO_1654 (O_1654,N_24832,N_24947);
and UO_1655 (O_1655,N_24930,N_24991);
nor UO_1656 (O_1656,N_24879,N_24851);
or UO_1657 (O_1657,N_24815,N_24943);
and UO_1658 (O_1658,N_24804,N_24800);
or UO_1659 (O_1659,N_24964,N_24932);
and UO_1660 (O_1660,N_24920,N_24857);
nor UO_1661 (O_1661,N_24956,N_24859);
nand UO_1662 (O_1662,N_24871,N_24874);
and UO_1663 (O_1663,N_24992,N_24822);
nand UO_1664 (O_1664,N_24886,N_24997);
xnor UO_1665 (O_1665,N_24821,N_24966);
or UO_1666 (O_1666,N_24922,N_24880);
nor UO_1667 (O_1667,N_24880,N_24929);
and UO_1668 (O_1668,N_24836,N_24974);
and UO_1669 (O_1669,N_24916,N_24886);
or UO_1670 (O_1670,N_24818,N_24810);
xnor UO_1671 (O_1671,N_24880,N_24866);
nor UO_1672 (O_1672,N_24810,N_24885);
xnor UO_1673 (O_1673,N_24884,N_24945);
nor UO_1674 (O_1674,N_24896,N_24803);
nand UO_1675 (O_1675,N_24901,N_24804);
and UO_1676 (O_1676,N_24805,N_24904);
nand UO_1677 (O_1677,N_24917,N_24891);
nand UO_1678 (O_1678,N_24973,N_24859);
and UO_1679 (O_1679,N_24942,N_24805);
nor UO_1680 (O_1680,N_24938,N_24931);
nor UO_1681 (O_1681,N_24941,N_24831);
nor UO_1682 (O_1682,N_24802,N_24977);
and UO_1683 (O_1683,N_24818,N_24879);
or UO_1684 (O_1684,N_24991,N_24945);
and UO_1685 (O_1685,N_24908,N_24873);
or UO_1686 (O_1686,N_24895,N_24859);
and UO_1687 (O_1687,N_24849,N_24994);
xnor UO_1688 (O_1688,N_24957,N_24941);
nand UO_1689 (O_1689,N_24884,N_24994);
nor UO_1690 (O_1690,N_24955,N_24885);
nor UO_1691 (O_1691,N_24901,N_24956);
or UO_1692 (O_1692,N_24821,N_24981);
nand UO_1693 (O_1693,N_24954,N_24815);
nand UO_1694 (O_1694,N_24974,N_24962);
xnor UO_1695 (O_1695,N_24834,N_24946);
xnor UO_1696 (O_1696,N_24842,N_24961);
xnor UO_1697 (O_1697,N_24816,N_24988);
nand UO_1698 (O_1698,N_24927,N_24839);
nor UO_1699 (O_1699,N_24971,N_24961);
nor UO_1700 (O_1700,N_24881,N_24893);
xnor UO_1701 (O_1701,N_24841,N_24881);
and UO_1702 (O_1702,N_24891,N_24931);
nand UO_1703 (O_1703,N_24824,N_24823);
and UO_1704 (O_1704,N_24916,N_24936);
and UO_1705 (O_1705,N_24968,N_24817);
nor UO_1706 (O_1706,N_24867,N_24936);
or UO_1707 (O_1707,N_24858,N_24805);
and UO_1708 (O_1708,N_24963,N_24805);
and UO_1709 (O_1709,N_24995,N_24998);
xor UO_1710 (O_1710,N_24986,N_24811);
or UO_1711 (O_1711,N_24848,N_24864);
or UO_1712 (O_1712,N_24967,N_24902);
xor UO_1713 (O_1713,N_24892,N_24819);
and UO_1714 (O_1714,N_24903,N_24892);
xor UO_1715 (O_1715,N_24891,N_24860);
and UO_1716 (O_1716,N_24835,N_24943);
nor UO_1717 (O_1717,N_24849,N_24834);
nor UO_1718 (O_1718,N_24968,N_24879);
nand UO_1719 (O_1719,N_24895,N_24914);
and UO_1720 (O_1720,N_24850,N_24893);
or UO_1721 (O_1721,N_24993,N_24917);
nand UO_1722 (O_1722,N_24853,N_24847);
xor UO_1723 (O_1723,N_24836,N_24847);
nor UO_1724 (O_1724,N_24928,N_24853);
or UO_1725 (O_1725,N_24811,N_24827);
and UO_1726 (O_1726,N_24830,N_24915);
xor UO_1727 (O_1727,N_24897,N_24957);
or UO_1728 (O_1728,N_24925,N_24984);
xnor UO_1729 (O_1729,N_24828,N_24926);
nor UO_1730 (O_1730,N_24849,N_24920);
xnor UO_1731 (O_1731,N_24890,N_24866);
or UO_1732 (O_1732,N_24873,N_24825);
or UO_1733 (O_1733,N_24819,N_24983);
nand UO_1734 (O_1734,N_24944,N_24937);
nand UO_1735 (O_1735,N_24815,N_24932);
nand UO_1736 (O_1736,N_24854,N_24891);
or UO_1737 (O_1737,N_24805,N_24952);
nand UO_1738 (O_1738,N_24962,N_24827);
xnor UO_1739 (O_1739,N_24869,N_24896);
or UO_1740 (O_1740,N_24829,N_24898);
nor UO_1741 (O_1741,N_24986,N_24831);
nand UO_1742 (O_1742,N_24807,N_24974);
xnor UO_1743 (O_1743,N_24835,N_24913);
nor UO_1744 (O_1744,N_24800,N_24963);
or UO_1745 (O_1745,N_24976,N_24929);
xnor UO_1746 (O_1746,N_24900,N_24825);
and UO_1747 (O_1747,N_24945,N_24960);
or UO_1748 (O_1748,N_24921,N_24832);
and UO_1749 (O_1749,N_24926,N_24864);
xnor UO_1750 (O_1750,N_24805,N_24844);
or UO_1751 (O_1751,N_24947,N_24863);
xnor UO_1752 (O_1752,N_24854,N_24925);
and UO_1753 (O_1753,N_24961,N_24893);
nor UO_1754 (O_1754,N_24930,N_24844);
nand UO_1755 (O_1755,N_24975,N_24939);
nor UO_1756 (O_1756,N_24909,N_24892);
nand UO_1757 (O_1757,N_24965,N_24830);
and UO_1758 (O_1758,N_24908,N_24871);
nand UO_1759 (O_1759,N_24929,N_24819);
nor UO_1760 (O_1760,N_24865,N_24857);
or UO_1761 (O_1761,N_24981,N_24847);
nand UO_1762 (O_1762,N_24859,N_24934);
nor UO_1763 (O_1763,N_24957,N_24943);
nand UO_1764 (O_1764,N_24999,N_24834);
and UO_1765 (O_1765,N_24937,N_24897);
or UO_1766 (O_1766,N_24994,N_24827);
nor UO_1767 (O_1767,N_24984,N_24863);
or UO_1768 (O_1768,N_24995,N_24934);
nor UO_1769 (O_1769,N_24888,N_24889);
xnor UO_1770 (O_1770,N_24817,N_24889);
or UO_1771 (O_1771,N_24892,N_24936);
nor UO_1772 (O_1772,N_24995,N_24844);
nor UO_1773 (O_1773,N_24973,N_24893);
or UO_1774 (O_1774,N_24967,N_24931);
or UO_1775 (O_1775,N_24972,N_24915);
or UO_1776 (O_1776,N_24868,N_24967);
or UO_1777 (O_1777,N_24872,N_24961);
or UO_1778 (O_1778,N_24945,N_24890);
xnor UO_1779 (O_1779,N_24831,N_24821);
nor UO_1780 (O_1780,N_24892,N_24960);
nor UO_1781 (O_1781,N_24863,N_24829);
nor UO_1782 (O_1782,N_24893,N_24827);
nand UO_1783 (O_1783,N_24913,N_24842);
nor UO_1784 (O_1784,N_24914,N_24956);
nand UO_1785 (O_1785,N_24819,N_24853);
and UO_1786 (O_1786,N_24931,N_24918);
or UO_1787 (O_1787,N_24874,N_24852);
nand UO_1788 (O_1788,N_24953,N_24895);
or UO_1789 (O_1789,N_24976,N_24952);
xnor UO_1790 (O_1790,N_24920,N_24998);
nor UO_1791 (O_1791,N_24866,N_24945);
and UO_1792 (O_1792,N_24902,N_24867);
and UO_1793 (O_1793,N_24934,N_24892);
and UO_1794 (O_1794,N_24844,N_24873);
nand UO_1795 (O_1795,N_24830,N_24910);
nand UO_1796 (O_1796,N_24840,N_24922);
xor UO_1797 (O_1797,N_24928,N_24938);
or UO_1798 (O_1798,N_24964,N_24923);
nand UO_1799 (O_1799,N_24820,N_24803);
and UO_1800 (O_1800,N_24871,N_24862);
and UO_1801 (O_1801,N_24967,N_24831);
nor UO_1802 (O_1802,N_24803,N_24999);
nand UO_1803 (O_1803,N_24897,N_24871);
xnor UO_1804 (O_1804,N_24998,N_24902);
nand UO_1805 (O_1805,N_24888,N_24821);
xnor UO_1806 (O_1806,N_24820,N_24813);
and UO_1807 (O_1807,N_24990,N_24987);
nor UO_1808 (O_1808,N_24883,N_24895);
or UO_1809 (O_1809,N_24842,N_24992);
nor UO_1810 (O_1810,N_24907,N_24805);
nand UO_1811 (O_1811,N_24941,N_24930);
or UO_1812 (O_1812,N_24898,N_24919);
or UO_1813 (O_1813,N_24803,N_24998);
nand UO_1814 (O_1814,N_24860,N_24973);
nand UO_1815 (O_1815,N_24913,N_24909);
or UO_1816 (O_1816,N_24905,N_24979);
and UO_1817 (O_1817,N_24815,N_24867);
xnor UO_1818 (O_1818,N_24887,N_24857);
nor UO_1819 (O_1819,N_24973,N_24922);
or UO_1820 (O_1820,N_24980,N_24875);
nand UO_1821 (O_1821,N_24874,N_24811);
or UO_1822 (O_1822,N_24842,N_24920);
nor UO_1823 (O_1823,N_24880,N_24837);
and UO_1824 (O_1824,N_24886,N_24803);
nand UO_1825 (O_1825,N_24826,N_24922);
nor UO_1826 (O_1826,N_24912,N_24894);
or UO_1827 (O_1827,N_24878,N_24909);
or UO_1828 (O_1828,N_24995,N_24936);
nor UO_1829 (O_1829,N_24882,N_24830);
nor UO_1830 (O_1830,N_24955,N_24976);
and UO_1831 (O_1831,N_24988,N_24825);
or UO_1832 (O_1832,N_24932,N_24869);
xnor UO_1833 (O_1833,N_24846,N_24863);
and UO_1834 (O_1834,N_24968,N_24826);
nor UO_1835 (O_1835,N_24863,N_24975);
nor UO_1836 (O_1836,N_24915,N_24812);
or UO_1837 (O_1837,N_24963,N_24894);
nand UO_1838 (O_1838,N_24850,N_24924);
xor UO_1839 (O_1839,N_24825,N_24938);
and UO_1840 (O_1840,N_24999,N_24947);
nand UO_1841 (O_1841,N_24842,N_24813);
xnor UO_1842 (O_1842,N_24937,N_24993);
xor UO_1843 (O_1843,N_24937,N_24826);
or UO_1844 (O_1844,N_24994,N_24970);
or UO_1845 (O_1845,N_24863,N_24819);
nand UO_1846 (O_1846,N_24903,N_24840);
xor UO_1847 (O_1847,N_24976,N_24964);
and UO_1848 (O_1848,N_24826,N_24824);
or UO_1849 (O_1849,N_24922,N_24901);
and UO_1850 (O_1850,N_24934,N_24926);
xor UO_1851 (O_1851,N_24836,N_24907);
nor UO_1852 (O_1852,N_24801,N_24869);
xor UO_1853 (O_1853,N_24935,N_24872);
nor UO_1854 (O_1854,N_24955,N_24860);
and UO_1855 (O_1855,N_24821,N_24931);
and UO_1856 (O_1856,N_24868,N_24867);
nor UO_1857 (O_1857,N_24885,N_24854);
or UO_1858 (O_1858,N_24882,N_24924);
nand UO_1859 (O_1859,N_24905,N_24964);
and UO_1860 (O_1860,N_24917,N_24828);
nand UO_1861 (O_1861,N_24901,N_24937);
nand UO_1862 (O_1862,N_24859,N_24881);
xnor UO_1863 (O_1863,N_24904,N_24806);
nand UO_1864 (O_1864,N_24893,N_24886);
or UO_1865 (O_1865,N_24884,N_24919);
and UO_1866 (O_1866,N_24932,N_24813);
xnor UO_1867 (O_1867,N_24992,N_24961);
or UO_1868 (O_1868,N_24818,N_24867);
and UO_1869 (O_1869,N_24823,N_24935);
nand UO_1870 (O_1870,N_24855,N_24841);
nand UO_1871 (O_1871,N_24874,N_24858);
nor UO_1872 (O_1872,N_24816,N_24974);
or UO_1873 (O_1873,N_24875,N_24833);
xnor UO_1874 (O_1874,N_24939,N_24955);
nor UO_1875 (O_1875,N_24974,N_24802);
nand UO_1876 (O_1876,N_24854,N_24910);
xnor UO_1877 (O_1877,N_24833,N_24802);
or UO_1878 (O_1878,N_24884,N_24854);
and UO_1879 (O_1879,N_24939,N_24946);
nor UO_1880 (O_1880,N_24805,N_24912);
xnor UO_1881 (O_1881,N_24877,N_24973);
nor UO_1882 (O_1882,N_24917,N_24983);
nand UO_1883 (O_1883,N_24833,N_24979);
and UO_1884 (O_1884,N_24854,N_24907);
nor UO_1885 (O_1885,N_24823,N_24850);
nor UO_1886 (O_1886,N_24951,N_24831);
nand UO_1887 (O_1887,N_24949,N_24827);
or UO_1888 (O_1888,N_24959,N_24996);
nor UO_1889 (O_1889,N_24976,N_24918);
or UO_1890 (O_1890,N_24830,N_24912);
nand UO_1891 (O_1891,N_24970,N_24968);
xnor UO_1892 (O_1892,N_24867,N_24852);
nor UO_1893 (O_1893,N_24933,N_24978);
nor UO_1894 (O_1894,N_24899,N_24838);
nand UO_1895 (O_1895,N_24989,N_24934);
xnor UO_1896 (O_1896,N_24934,N_24946);
nor UO_1897 (O_1897,N_24897,N_24919);
xor UO_1898 (O_1898,N_24926,N_24968);
or UO_1899 (O_1899,N_24997,N_24908);
nand UO_1900 (O_1900,N_24917,N_24831);
xnor UO_1901 (O_1901,N_24942,N_24915);
xnor UO_1902 (O_1902,N_24990,N_24886);
nand UO_1903 (O_1903,N_24883,N_24977);
nand UO_1904 (O_1904,N_24943,N_24885);
xnor UO_1905 (O_1905,N_24973,N_24926);
or UO_1906 (O_1906,N_24963,N_24937);
nor UO_1907 (O_1907,N_24987,N_24927);
nor UO_1908 (O_1908,N_24952,N_24855);
xor UO_1909 (O_1909,N_24814,N_24979);
nor UO_1910 (O_1910,N_24954,N_24804);
nand UO_1911 (O_1911,N_24820,N_24995);
or UO_1912 (O_1912,N_24853,N_24906);
and UO_1913 (O_1913,N_24961,N_24844);
nand UO_1914 (O_1914,N_24901,N_24934);
nor UO_1915 (O_1915,N_24952,N_24882);
and UO_1916 (O_1916,N_24897,N_24804);
nand UO_1917 (O_1917,N_24827,N_24946);
nand UO_1918 (O_1918,N_24829,N_24823);
or UO_1919 (O_1919,N_24852,N_24849);
xor UO_1920 (O_1920,N_24821,N_24924);
or UO_1921 (O_1921,N_24977,N_24978);
nor UO_1922 (O_1922,N_24883,N_24939);
xor UO_1923 (O_1923,N_24861,N_24869);
and UO_1924 (O_1924,N_24900,N_24887);
or UO_1925 (O_1925,N_24814,N_24830);
or UO_1926 (O_1926,N_24947,N_24937);
xor UO_1927 (O_1927,N_24949,N_24909);
xor UO_1928 (O_1928,N_24950,N_24893);
nor UO_1929 (O_1929,N_24889,N_24996);
or UO_1930 (O_1930,N_24918,N_24889);
nor UO_1931 (O_1931,N_24855,N_24809);
nand UO_1932 (O_1932,N_24910,N_24873);
or UO_1933 (O_1933,N_24849,N_24929);
nor UO_1934 (O_1934,N_24925,N_24993);
and UO_1935 (O_1935,N_24939,N_24922);
nor UO_1936 (O_1936,N_24952,N_24919);
and UO_1937 (O_1937,N_24821,N_24900);
xnor UO_1938 (O_1938,N_24837,N_24932);
xnor UO_1939 (O_1939,N_24973,N_24853);
nand UO_1940 (O_1940,N_24922,N_24888);
nand UO_1941 (O_1941,N_24866,N_24901);
nor UO_1942 (O_1942,N_24825,N_24837);
and UO_1943 (O_1943,N_24992,N_24911);
or UO_1944 (O_1944,N_24912,N_24998);
and UO_1945 (O_1945,N_24965,N_24905);
nor UO_1946 (O_1946,N_24957,N_24997);
or UO_1947 (O_1947,N_24856,N_24899);
or UO_1948 (O_1948,N_24854,N_24844);
nor UO_1949 (O_1949,N_24873,N_24934);
or UO_1950 (O_1950,N_24944,N_24804);
or UO_1951 (O_1951,N_24828,N_24969);
or UO_1952 (O_1952,N_24995,N_24804);
nand UO_1953 (O_1953,N_24808,N_24864);
xnor UO_1954 (O_1954,N_24934,N_24869);
xnor UO_1955 (O_1955,N_24928,N_24931);
nor UO_1956 (O_1956,N_24872,N_24906);
xnor UO_1957 (O_1957,N_24830,N_24907);
nor UO_1958 (O_1958,N_24940,N_24870);
nor UO_1959 (O_1959,N_24892,N_24928);
and UO_1960 (O_1960,N_24953,N_24973);
xor UO_1961 (O_1961,N_24877,N_24871);
xnor UO_1962 (O_1962,N_24855,N_24913);
xnor UO_1963 (O_1963,N_24890,N_24848);
nor UO_1964 (O_1964,N_24815,N_24951);
and UO_1965 (O_1965,N_24806,N_24851);
xor UO_1966 (O_1966,N_24872,N_24802);
nand UO_1967 (O_1967,N_24854,N_24896);
and UO_1968 (O_1968,N_24989,N_24841);
and UO_1969 (O_1969,N_24999,N_24838);
or UO_1970 (O_1970,N_24905,N_24911);
nor UO_1971 (O_1971,N_24917,N_24968);
nand UO_1972 (O_1972,N_24905,N_24892);
nand UO_1973 (O_1973,N_24987,N_24999);
nand UO_1974 (O_1974,N_24873,N_24836);
nand UO_1975 (O_1975,N_24970,N_24824);
or UO_1976 (O_1976,N_24836,N_24965);
nand UO_1977 (O_1977,N_24970,N_24912);
xnor UO_1978 (O_1978,N_24890,N_24982);
or UO_1979 (O_1979,N_24834,N_24901);
or UO_1980 (O_1980,N_24838,N_24805);
and UO_1981 (O_1981,N_24806,N_24898);
or UO_1982 (O_1982,N_24900,N_24846);
nor UO_1983 (O_1983,N_24973,N_24856);
nor UO_1984 (O_1984,N_24878,N_24969);
xnor UO_1985 (O_1985,N_24850,N_24939);
nand UO_1986 (O_1986,N_24914,N_24832);
nand UO_1987 (O_1987,N_24913,N_24955);
nand UO_1988 (O_1988,N_24835,N_24892);
nand UO_1989 (O_1989,N_24903,N_24850);
and UO_1990 (O_1990,N_24808,N_24910);
nor UO_1991 (O_1991,N_24829,N_24815);
or UO_1992 (O_1992,N_24904,N_24886);
or UO_1993 (O_1993,N_24803,N_24948);
nand UO_1994 (O_1994,N_24826,N_24939);
nor UO_1995 (O_1995,N_24921,N_24846);
or UO_1996 (O_1996,N_24987,N_24960);
nor UO_1997 (O_1997,N_24824,N_24825);
xnor UO_1998 (O_1998,N_24881,N_24821);
and UO_1999 (O_1999,N_24887,N_24906);
nand UO_2000 (O_2000,N_24973,N_24981);
and UO_2001 (O_2001,N_24841,N_24996);
nand UO_2002 (O_2002,N_24868,N_24830);
and UO_2003 (O_2003,N_24987,N_24954);
nand UO_2004 (O_2004,N_24903,N_24889);
nand UO_2005 (O_2005,N_24838,N_24800);
or UO_2006 (O_2006,N_24889,N_24994);
xnor UO_2007 (O_2007,N_24809,N_24941);
or UO_2008 (O_2008,N_24971,N_24926);
or UO_2009 (O_2009,N_24966,N_24826);
nor UO_2010 (O_2010,N_24895,N_24874);
xor UO_2011 (O_2011,N_24983,N_24935);
nand UO_2012 (O_2012,N_24808,N_24973);
nand UO_2013 (O_2013,N_24811,N_24803);
and UO_2014 (O_2014,N_24914,N_24881);
and UO_2015 (O_2015,N_24802,N_24902);
xor UO_2016 (O_2016,N_24995,N_24899);
and UO_2017 (O_2017,N_24843,N_24892);
and UO_2018 (O_2018,N_24994,N_24811);
or UO_2019 (O_2019,N_24859,N_24804);
and UO_2020 (O_2020,N_24809,N_24874);
nand UO_2021 (O_2021,N_24917,N_24963);
nand UO_2022 (O_2022,N_24805,N_24877);
xnor UO_2023 (O_2023,N_24956,N_24891);
nand UO_2024 (O_2024,N_24819,N_24960);
xnor UO_2025 (O_2025,N_24816,N_24935);
nor UO_2026 (O_2026,N_24908,N_24899);
xnor UO_2027 (O_2027,N_24830,N_24898);
or UO_2028 (O_2028,N_24873,N_24865);
nand UO_2029 (O_2029,N_24964,N_24806);
nor UO_2030 (O_2030,N_24964,N_24823);
nor UO_2031 (O_2031,N_24913,N_24828);
and UO_2032 (O_2032,N_24963,N_24958);
nor UO_2033 (O_2033,N_24952,N_24886);
nand UO_2034 (O_2034,N_24984,N_24911);
nor UO_2035 (O_2035,N_24831,N_24813);
and UO_2036 (O_2036,N_24974,N_24861);
nand UO_2037 (O_2037,N_24948,N_24897);
and UO_2038 (O_2038,N_24933,N_24853);
and UO_2039 (O_2039,N_24934,N_24960);
or UO_2040 (O_2040,N_24937,N_24875);
xnor UO_2041 (O_2041,N_24807,N_24950);
or UO_2042 (O_2042,N_24865,N_24936);
xor UO_2043 (O_2043,N_24943,N_24934);
or UO_2044 (O_2044,N_24998,N_24874);
nor UO_2045 (O_2045,N_24913,N_24887);
and UO_2046 (O_2046,N_24878,N_24999);
xor UO_2047 (O_2047,N_24821,N_24943);
nand UO_2048 (O_2048,N_24908,N_24944);
xor UO_2049 (O_2049,N_24915,N_24843);
or UO_2050 (O_2050,N_24935,N_24913);
nor UO_2051 (O_2051,N_24958,N_24892);
xor UO_2052 (O_2052,N_24819,N_24837);
and UO_2053 (O_2053,N_24954,N_24906);
nor UO_2054 (O_2054,N_24869,N_24949);
nand UO_2055 (O_2055,N_24981,N_24924);
nor UO_2056 (O_2056,N_24814,N_24891);
xor UO_2057 (O_2057,N_24802,N_24961);
nand UO_2058 (O_2058,N_24892,N_24971);
and UO_2059 (O_2059,N_24893,N_24857);
or UO_2060 (O_2060,N_24832,N_24831);
or UO_2061 (O_2061,N_24974,N_24981);
or UO_2062 (O_2062,N_24881,N_24952);
nand UO_2063 (O_2063,N_24931,N_24813);
and UO_2064 (O_2064,N_24820,N_24998);
or UO_2065 (O_2065,N_24915,N_24847);
nand UO_2066 (O_2066,N_24889,N_24942);
xnor UO_2067 (O_2067,N_24960,N_24826);
xor UO_2068 (O_2068,N_24990,N_24959);
or UO_2069 (O_2069,N_24981,N_24882);
or UO_2070 (O_2070,N_24985,N_24802);
or UO_2071 (O_2071,N_24807,N_24909);
nor UO_2072 (O_2072,N_24907,N_24980);
nor UO_2073 (O_2073,N_24947,N_24989);
or UO_2074 (O_2074,N_24918,N_24956);
and UO_2075 (O_2075,N_24846,N_24800);
and UO_2076 (O_2076,N_24808,N_24919);
nand UO_2077 (O_2077,N_24864,N_24806);
nand UO_2078 (O_2078,N_24943,N_24803);
nand UO_2079 (O_2079,N_24819,N_24820);
nand UO_2080 (O_2080,N_24960,N_24895);
or UO_2081 (O_2081,N_24950,N_24847);
or UO_2082 (O_2082,N_24906,N_24810);
nor UO_2083 (O_2083,N_24967,N_24988);
and UO_2084 (O_2084,N_24899,N_24891);
xor UO_2085 (O_2085,N_24896,N_24880);
or UO_2086 (O_2086,N_24899,N_24811);
xnor UO_2087 (O_2087,N_24890,N_24821);
nor UO_2088 (O_2088,N_24863,N_24986);
and UO_2089 (O_2089,N_24998,N_24812);
nand UO_2090 (O_2090,N_24973,N_24845);
and UO_2091 (O_2091,N_24920,N_24804);
or UO_2092 (O_2092,N_24910,N_24801);
xnor UO_2093 (O_2093,N_24892,N_24895);
nor UO_2094 (O_2094,N_24856,N_24822);
nor UO_2095 (O_2095,N_24950,N_24886);
nand UO_2096 (O_2096,N_24954,N_24817);
xnor UO_2097 (O_2097,N_24965,N_24838);
nand UO_2098 (O_2098,N_24874,N_24800);
and UO_2099 (O_2099,N_24847,N_24863);
nand UO_2100 (O_2100,N_24889,N_24924);
nor UO_2101 (O_2101,N_24981,N_24877);
or UO_2102 (O_2102,N_24949,N_24819);
or UO_2103 (O_2103,N_24809,N_24848);
xor UO_2104 (O_2104,N_24977,N_24810);
nand UO_2105 (O_2105,N_24891,N_24971);
and UO_2106 (O_2106,N_24897,N_24953);
or UO_2107 (O_2107,N_24986,N_24847);
nand UO_2108 (O_2108,N_24886,N_24894);
nor UO_2109 (O_2109,N_24999,N_24901);
and UO_2110 (O_2110,N_24946,N_24819);
xor UO_2111 (O_2111,N_24938,N_24845);
nand UO_2112 (O_2112,N_24950,N_24833);
nand UO_2113 (O_2113,N_24895,N_24834);
nor UO_2114 (O_2114,N_24908,N_24982);
xor UO_2115 (O_2115,N_24871,N_24854);
or UO_2116 (O_2116,N_24922,N_24987);
xor UO_2117 (O_2117,N_24964,N_24970);
nand UO_2118 (O_2118,N_24987,N_24961);
nor UO_2119 (O_2119,N_24907,N_24952);
nor UO_2120 (O_2120,N_24855,N_24888);
xnor UO_2121 (O_2121,N_24912,N_24927);
nand UO_2122 (O_2122,N_24900,N_24867);
nand UO_2123 (O_2123,N_24937,N_24932);
nand UO_2124 (O_2124,N_24974,N_24833);
and UO_2125 (O_2125,N_24835,N_24979);
and UO_2126 (O_2126,N_24865,N_24949);
xnor UO_2127 (O_2127,N_24872,N_24999);
xnor UO_2128 (O_2128,N_24921,N_24868);
nor UO_2129 (O_2129,N_24940,N_24862);
nor UO_2130 (O_2130,N_24937,N_24825);
xnor UO_2131 (O_2131,N_24979,N_24874);
nand UO_2132 (O_2132,N_24897,N_24989);
xnor UO_2133 (O_2133,N_24960,N_24816);
or UO_2134 (O_2134,N_24953,N_24940);
nand UO_2135 (O_2135,N_24913,N_24924);
nand UO_2136 (O_2136,N_24984,N_24901);
and UO_2137 (O_2137,N_24946,N_24999);
and UO_2138 (O_2138,N_24985,N_24897);
nor UO_2139 (O_2139,N_24917,N_24887);
nand UO_2140 (O_2140,N_24969,N_24928);
and UO_2141 (O_2141,N_24944,N_24807);
nand UO_2142 (O_2142,N_24917,N_24875);
nor UO_2143 (O_2143,N_24994,N_24808);
nand UO_2144 (O_2144,N_24852,N_24889);
nand UO_2145 (O_2145,N_24894,N_24929);
nand UO_2146 (O_2146,N_24865,N_24859);
and UO_2147 (O_2147,N_24887,N_24842);
and UO_2148 (O_2148,N_24860,N_24974);
nand UO_2149 (O_2149,N_24968,N_24969);
and UO_2150 (O_2150,N_24890,N_24816);
xor UO_2151 (O_2151,N_24911,N_24801);
and UO_2152 (O_2152,N_24814,N_24811);
nor UO_2153 (O_2153,N_24964,N_24951);
or UO_2154 (O_2154,N_24821,N_24851);
xnor UO_2155 (O_2155,N_24957,N_24949);
nand UO_2156 (O_2156,N_24891,N_24822);
xnor UO_2157 (O_2157,N_24885,N_24919);
xnor UO_2158 (O_2158,N_24956,N_24951);
or UO_2159 (O_2159,N_24987,N_24988);
nor UO_2160 (O_2160,N_24922,N_24924);
xor UO_2161 (O_2161,N_24996,N_24866);
nor UO_2162 (O_2162,N_24859,N_24924);
nand UO_2163 (O_2163,N_24994,N_24904);
or UO_2164 (O_2164,N_24946,N_24893);
xnor UO_2165 (O_2165,N_24902,N_24993);
and UO_2166 (O_2166,N_24940,N_24974);
xnor UO_2167 (O_2167,N_24828,N_24800);
nand UO_2168 (O_2168,N_24945,N_24829);
and UO_2169 (O_2169,N_24942,N_24880);
and UO_2170 (O_2170,N_24818,N_24912);
nand UO_2171 (O_2171,N_24872,N_24831);
nand UO_2172 (O_2172,N_24899,N_24892);
nor UO_2173 (O_2173,N_24832,N_24815);
and UO_2174 (O_2174,N_24841,N_24806);
or UO_2175 (O_2175,N_24919,N_24971);
or UO_2176 (O_2176,N_24851,N_24820);
nand UO_2177 (O_2177,N_24840,N_24812);
nor UO_2178 (O_2178,N_24939,N_24866);
nand UO_2179 (O_2179,N_24994,N_24836);
nand UO_2180 (O_2180,N_24859,N_24874);
and UO_2181 (O_2181,N_24926,N_24826);
nand UO_2182 (O_2182,N_24804,N_24858);
nor UO_2183 (O_2183,N_24837,N_24864);
and UO_2184 (O_2184,N_24868,N_24908);
and UO_2185 (O_2185,N_24813,N_24802);
nor UO_2186 (O_2186,N_24984,N_24992);
xnor UO_2187 (O_2187,N_24926,N_24897);
xor UO_2188 (O_2188,N_24983,N_24837);
nand UO_2189 (O_2189,N_24825,N_24820);
nand UO_2190 (O_2190,N_24880,N_24873);
nor UO_2191 (O_2191,N_24818,N_24864);
nand UO_2192 (O_2192,N_24964,N_24957);
or UO_2193 (O_2193,N_24978,N_24905);
xnor UO_2194 (O_2194,N_24892,N_24940);
nor UO_2195 (O_2195,N_24823,N_24805);
xnor UO_2196 (O_2196,N_24916,N_24850);
nor UO_2197 (O_2197,N_24839,N_24830);
xnor UO_2198 (O_2198,N_24913,N_24810);
xnor UO_2199 (O_2199,N_24970,N_24990);
and UO_2200 (O_2200,N_24962,N_24897);
and UO_2201 (O_2201,N_24949,N_24901);
nor UO_2202 (O_2202,N_24985,N_24945);
nand UO_2203 (O_2203,N_24885,N_24966);
xor UO_2204 (O_2204,N_24962,N_24892);
nand UO_2205 (O_2205,N_24833,N_24848);
xnor UO_2206 (O_2206,N_24999,N_24939);
nand UO_2207 (O_2207,N_24810,N_24994);
nand UO_2208 (O_2208,N_24947,N_24992);
nand UO_2209 (O_2209,N_24861,N_24948);
nand UO_2210 (O_2210,N_24848,N_24991);
nand UO_2211 (O_2211,N_24843,N_24837);
or UO_2212 (O_2212,N_24997,N_24983);
or UO_2213 (O_2213,N_24813,N_24901);
or UO_2214 (O_2214,N_24832,N_24905);
xor UO_2215 (O_2215,N_24985,N_24924);
and UO_2216 (O_2216,N_24930,N_24801);
nor UO_2217 (O_2217,N_24820,N_24876);
nand UO_2218 (O_2218,N_24875,N_24816);
or UO_2219 (O_2219,N_24850,N_24962);
nand UO_2220 (O_2220,N_24800,N_24885);
nand UO_2221 (O_2221,N_24939,N_24934);
or UO_2222 (O_2222,N_24867,N_24996);
or UO_2223 (O_2223,N_24842,N_24923);
nor UO_2224 (O_2224,N_24966,N_24898);
xnor UO_2225 (O_2225,N_24965,N_24895);
nand UO_2226 (O_2226,N_24922,N_24910);
and UO_2227 (O_2227,N_24900,N_24924);
nand UO_2228 (O_2228,N_24812,N_24804);
nor UO_2229 (O_2229,N_24928,N_24981);
xor UO_2230 (O_2230,N_24983,N_24929);
nand UO_2231 (O_2231,N_24935,N_24926);
xnor UO_2232 (O_2232,N_24811,N_24888);
xnor UO_2233 (O_2233,N_24811,N_24871);
nand UO_2234 (O_2234,N_24959,N_24880);
and UO_2235 (O_2235,N_24812,N_24921);
nand UO_2236 (O_2236,N_24889,N_24897);
and UO_2237 (O_2237,N_24978,N_24818);
nand UO_2238 (O_2238,N_24839,N_24835);
and UO_2239 (O_2239,N_24980,N_24908);
xor UO_2240 (O_2240,N_24868,N_24906);
and UO_2241 (O_2241,N_24803,N_24993);
and UO_2242 (O_2242,N_24855,N_24836);
xor UO_2243 (O_2243,N_24919,N_24929);
and UO_2244 (O_2244,N_24940,N_24972);
xor UO_2245 (O_2245,N_24929,N_24995);
or UO_2246 (O_2246,N_24999,N_24841);
and UO_2247 (O_2247,N_24892,N_24967);
nor UO_2248 (O_2248,N_24889,N_24952);
and UO_2249 (O_2249,N_24878,N_24929);
and UO_2250 (O_2250,N_24969,N_24948);
or UO_2251 (O_2251,N_24853,N_24814);
or UO_2252 (O_2252,N_24885,N_24952);
nand UO_2253 (O_2253,N_24826,N_24976);
or UO_2254 (O_2254,N_24831,N_24898);
xnor UO_2255 (O_2255,N_24832,N_24813);
nor UO_2256 (O_2256,N_24995,N_24878);
and UO_2257 (O_2257,N_24917,N_24908);
and UO_2258 (O_2258,N_24974,N_24846);
xor UO_2259 (O_2259,N_24931,N_24989);
and UO_2260 (O_2260,N_24967,N_24981);
nor UO_2261 (O_2261,N_24910,N_24887);
and UO_2262 (O_2262,N_24919,N_24836);
or UO_2263 (O_2263,N_24998,N_24849);
xnor UO_2264 (O_2264,N_24800,N_24883);
or UO_2265 (O_2265,N_24933,N_24803);
or UO_2266 (O_2266,N_24810,N_24931);
or UO_2267 (O_2267,N_24870,N_24972);
or UO_2268 (O_2268,N_24905,N_24969);
and UO_2269 (O_2269,N_24956,N_24974);
xnor UO_2270 (O_2270,N_24998,N_24951);
nand UO_2271 (O_2271,N_24890,N_24830);
xnor UO_2272 (O_2272,N_24958,N_24899);
or UO_2273 (O_2273,N_24958,N_24914);
or UO_2274 (O_2274,N_24903,N_24828);
nor UO_2275 (O_2275,N_24976,N_24917);
or UO_2276 (O_2276,N_24961,N_24950);
or UO_2277 (O_2277,N_24846,N_24933);
xnor UO_2278 (O_2278,N_24873,N_24871);
or UO_2279 (O_2279,N_24926,N_24963);
or UO_2280 (O_2280,N_24866,N_24895);
and UO_2281 (O_2281,N_24976,N_24992);
or UO_2282 (O_2282,N_24829,N_24830);
and UO_2283 (O_2283,N_24997,N_24851);
and UO_2284 (O_2284,N_24874,N_24849);
and UO_2285 (O_2285,N_24982,N_24981);
xor UO_2286 (O_2286,N_24980,N_24815);
nand UO_2287 (O_2287,N_24876,N_24944);
xnor UO_2288 (O_2288,N_24840,N_24967);
nor UO_2289 (O_2289,N_24834,N_24980);
nor UO_2290 (O_2290,N_24937,N_24995);
nor UO_2291 (O_2291,N_24810,N_24920);
xnor UO_2292 (O_2292,N_24817,N_24988);
nor UO_2293 (O_2293,N_24862,N_24929);
or UO_2294 (O_2294,N_24812,N_24961);
nand UO_2295 (O_2295,N_24939,N_24882);
nor UO_2296 (O_2296,N_24882,N_24853);
xnor UO_2297 (O_2297,N_24807,N_24880);
or UO_2298 (O_2298,N_24998,N_24868);
nor UO_2299 (O_2299,N_24918,N_24905);
xor UO_2300 (O_2300,N_24974,N_24992);
nand UO_2301 (O_2301,N_24900,N_24891);
xnor UO_2302 (O_2302,N_24995,N_24843);
or UO_2303 (O_2303,N_24835,N_24916);
nor UO_2304 (O_2304,N_24978,N_24840);
nor UO_2305 (O_2305,N_24976,N_24873);
nand UO_2306 (O_2306,N_24841,N_24865);
nand UO_2307 (O_2307,N_24829,N_24878);
nor UO_2308 (O_2308,N_24984,N_24856);
or UO_2309 (O_2309,N_24974,N_24873);
or UO_2310 (O_2310,N_24832,N_24840);
xnor UO_2311 (O_2311,N_24852,N_24879);
nor UO_2312 (O_2312,N_24866,N_24948);
nor UO_2313 (O_2313,N_24859,N_24901);
nor UO_2314 (O_2314,N_24858,N_24895);
xor UO_2315 (O_2315,N_24968,N_24907);
and UO_2316 (O_2316,N_24988,N_24889);
or UO_2317 (O_2317,N_24877,N_24897);
or UO_2318 (O_2318,N_24930,N_24811);
and UO_2319 (O_2319,N_24887,N_24908);
nor UO_2320 (O_2320,N_24878,N_24937);
nor UO_2321 (O_2321,N_24996,N_24802);
nand UO_2322 (O_2322,N_24920,N_24846);
and UO_2323 (O_2323,N_24953,N_24901);
nor UO_2324 (O_2324,N_24908,N_24966);
xor UO_2325 (O_2325,N_24884,N_24810);
xor UO_2326 (O_2326,N_24960,N_24992);
nor UO_2327 (O_2327,N_24919,N_24880);
xor UO_2328 (O_2328,N_24928,N_24974);
or UO_2329 (O_2329,N_24926,N_24887);
and UO_2330 (O_2330,N_24946,N_24874);
nand UO_2331 (O_2331,N_24809,N_24813);
nor UO_2332 (O_2332,N_24982,N_24845);
nand UO_2333 (O_2333,N_24933,N_24806);
nand UO_2334 (O_2334,N_24804,N_24931);
xor UO_2335 (O_2335,N_24950,N_24873);
or UO_2336 (O_2336,N_24875,N_24981);
nand UO_2337 (O_2337,N_24892,N_24875);
nand UO_2338 (O_2338,N_24824,N_24993);
nand UO_2339 (O_2339,N_24940,N_24833);
nand UO_2340 (O_2340,N_24968,N_24831);
xor UO_2341 (O_2341,N_24909,N_24979);
or UO_2342 (O_2342,N_24807,N_24806);
or UO_2343 (O_2343,N_24835,N_24982);
xnor UO_2344 (O_2344,N_24838,N_24853);
xnor UO_2345 (O_2345,N_24989,N_24999);
xnor UO_2346 (O_2346,N_24891,N_24803);
or UO_2347 (O_2347,N_24837,N_24830);
xor UO_2348 (O_2348,N_24809,N_24995);
xnor UO_2349 (O_2349,N_24991,N_24955);
or UO_2350 (O_2350,N_24989,N_24820);
and UO_2351 (O_2351,N_24951,N_24813);
or UO_2352 (O_2352,N_24968,N_24805);
and UO_2353 (O_2353,N_24918,N_24856);
xor UO_2354 (O_2354,N_24893,N_24929);
nor UO_2355 (O_2355,N_24866,N_24915);
nor UO_2356 (O_2356,N_24838,N_24985);
nor UO_2357 (O_2357,N_24850,N_24860);
or UO_2358 (O_2358,N_24810,N_24858);
xor UO_2359 (O_2359,N_24803,N_24913);
xor UO_2360 (O_2360,N_24890,N_24832);
nand UO_2361 (O_2361,N_24900,N_24965);
or UO_2362 (O_2362,N_24915,N_24973);
xnor UO_2363 (O_2363,N_24842,N_24867);
xnor UO_2364 (O_2364,N_24852,N_24805);
nor UO_2365 (O_2365,N_24919,N_24826);
nand UO_2366 (O_2366,N_24914,N_24810);
xor UO_2367 (O_2367,N_24854,N_24950);
xor UO_2368 (O_2368,N_24918,N_24924);
nor UO_2369 (O_2369,N_24910,N_24865);
or UO_2370 (O_2370,N_24964,N_24988);
or UO_2371 (O_2371,N_24865,N_24946);
and UO_2372 (O_2372,N_24862,N_24931);
and UO_2373 (O_2373,N_24898,N_24939);
nand UO_2374 (O_2374,N_24902,N_24828);
nor UO_2375 (O_2375,N_24907,N_24971);
xnor UO_2376 (O_2376,N_24967,N_24870);
nor UO_2377 (O_2377,N_24975,N_24875);
nand UO_2378 (O_2378,N_24917,N_24834);
nand UO_2379 (O_2379,N_24816,N_24892);
xor UO_2380 (O_2380,N_24989,N_24877);
xnor UO_2381 (O_2381,N_24914,N_24928);
nand UO_2382 (O_2382,N_24825,N_24948);
xnor UO_2383 (O_2383,N_24893,N_24891);
nor UO_2384 (O_2384,N_24953,N_24965);
nand UO_2385 (O_2385,N_24877,N_24921);
and UO_2386 (O_2386,N_24970,N_24849);
xnor UO_2387 (O_2387,N_24993,N_24835);
xnor UO_2388 (O_2388,N_24865,N_24872);
or UO_2389 (O_2389,N_24924,N_24917);
nand UO_2390 (O_2390,N_24822,N_24914);
xnor UO_2391 (O_2391,N_24842,N_24979);
and UO_2392 (O_2392,N_24992,N_24890);
nor UO_2393 (O_2393,N_24909,N_24965);
nor UO_2394 (O_2394,N_24839,N_24900);
nor UO_2395 (O_2395,N_24873,N_24824);
nand UO_2396 (O_2396,N_24835,N_24870);
nand UO_2397 (O_2397,N_24963,N_24883);
nand UO_2398 (O_2398,N_24822,N_24917);
xor UO_2399 (O_2399,N_24829,N_24921);
xnor UO_2400 (O_2400,N_24883,N_24867);
xor UO_2401 (O_2401,N_24933,N_24932);
nor UO_2402 (O_2402,N_24925,N_24910);
xor UO_2403 (O_2403,N_24803,N_24964);
nor UO_2404 (O_2404,N_24920,N_24971);
nand UO_2405 (O_2405,N_24840,N_24985);
and UO_2406 (O_2406,N_24991,N_24956);
nor UO_2407 (O_2407,N_24873,N_24810);
xnor UO_2408 (O_2408,N_24804,N_24984);
xnor UO_2409 (O_2409,N_24805,N_24931);
nand UO_2410 (O_2410,N_24862,N_24983);
xor UO_2411 (O_2411,N_24981,N_24900);
and UO_2412 (O_2412,N_24972,N_24951);
nor UO_2413 (O_2413,N_24911,N_24936);
nor UO_2414 (O_2414,N_24898,N_24839);
and UO_2415 (O_2415,N_24880,N_24955);
nand UO_2416 (O_2416,N_24855,N_24957);
and UO_2417 (O_2417,N_24816,N_24852);
nand UO_2418 (O_2418,N_24922,N_24966);
or UO_2419 (O_2419,N_24829,N_24967);
or UO_2420 (O_2420,N_24822,N_24996);
and UO_2421 (O_2421,N_24901,N_24997);
nor UO_2422 (O_2422,N_24852,N_24998);
nor UO_2423 (O_2423,N_24845,N_24994);
xnor UO_2424 (O_2424,N_24998,N_24905);
xnor UO_2425 (O_2425,N_24804,N_24819);
nand UO_2426 (O_2426,N_24899,N_24988);
or UO_2427 (O_2427,N_24991,N_24903);
xor UO_2428 (O_2428,N_24832,N_24873);
xor UO_2429 (O_2429,N_24924,N_24826);
or UO_2430 (O_2430,N_24987,N_24917);
nor UO_2431 (O_2431,N_24875,N_24900);
and UO_2432 (O_2432,N_24829,N_24996);
or UO_2433 (O_2433,N_24925,N_24806);
and UO_2434 (O_2434,N_24967,N_24880);
xnor UO_2435 (O_2435,N_24942,N_24844);
and UO_2436 (O_2436,N_24894,N_24930);
nand UO_2437 (O_2437,N_24879,N_24894);
xor UO_2438 (O_2438,N_24800,N_24875);
nor UO_2439 (O_2439,N_24820,N_24892);
or UO_2440 (O_2440,N_24984,N_24897);
nand UO_2441 (O_2441,N_24973,N_24848);
nor UO_2442 (O_2442,N_24990,N_24859);
and UO_2443 (O_2443,N_24973,N_24972);
nor UO_2444 (O_2444,N_24842,N_24987);
or UO_2445 (O_2445,N_24966,N_24980);
or UO_2446 (O_2446,N_24938,N_24894);
or UO_2447 (O_2447,N_24960,N_24917);
nand UO_2448 (O_2448,N_24813,N_24841);
nand UO_2449 (O_2449,N_24850,N_24955);
nor UO_2450 (O_2450,N_24858,N_24999);
and UO_2451 (O_2451,N_24935,N_24892);
nand UO_2452 (O_2452,N_24927,N_24851);
or UO_2453 (O_2453,N_24972,N_24824);
nor UO_2454 (O_2454,N_24966,N_24854);
xnor UO_2455 (O_2455,N_24821,N_24876);
or UO_2456 (O_2456,N_24991,N_24938);
xnor UO_2457 (O_2457,N_24805,N_24851);
or UO_2458 (O_2458,N_24992,N_24939);
xor UO_2459 (O_2459,N_24815,N_24979);
nand UO_2460 (O_2460,N_24964,N_24853);
nor UO_2461 (O_2461,N_24933,N_24889);
xor UO_2462 (O_2462,N_24819,N_24921);
xnor UO_2463 (O_2463,N_24828,N_24819);
nor UO_2464 (O_2464,N_24867,N_24965);
and UO_2465 (O_2465,N_24957,N_24876);
nor UO_2466 (O_2466,N_24816,N_24902);
and UO_2467 (O_2467,N_24933,N_24918);
nand UO_2468 (O_2468,N_24860,N_24930);
or UO_2469 (O_2469,N_24947,N_24852);
xnor UO_2470 (O_2470,N_24999,N_24933);
xnor UO_2471 (O_2471,N_24969,N_24961);
or UO_2472 (O_2472,N_24966,N_24910);
or UO_2473 (O_2473,N_24874,N_24907);
nand UO_2474 (O_2474,N_24904,N_24836);
nor UO_2475 (O_2475,N_24990,N_24882);
nor UO_2476 (O_2476,N_24855,N_24988);
xor UO_2477 (O_2477,N_24971,N_24811);
xnor UO_2478 (O_2478,N_24820,N_24805);
nand UO_2479 (O_2479,N_24849,N_24923);
xnor UO_2480 (O_2480,N_24993,N_24896);
and UO_2481 (O_2481,N_24950,N_24947);
and UO_2482 (O_2482,N_24944,N_24956);
xor UO_2483 (O_2483,N_24884,N_24838);
and UO_2484 (O_2484,N_24959,N_24977);
nor UO_2485 (O_2485,N_24882,N_24902);
and UO_2486 (O_2486,N_24956,N_24852);
nand UO_2487 (O_2487,N_24945,N_24891);
or UO_2488 (O_2488,N_24810,N_24972);
and UO_2489 (O_2489,N_24856,N_24900);
xnor UO_2490 (O_2490,N_24870,N_24815);
or UO_2491 (O_2491,N_24814,N_24992);
nand UO_2492 (O_2492,N_24879,N_24932);
nor UO_2493 (O_2493,N_24876,N_24800);
and UO_2494 (O_2494,N_24934,N_24863);
nand UO_2495 (O_2495,N_24947,N_24924);
and UO_2496 (O_2496,N_24890,N_24921);
or UO_2497 (O_2497,N_24938,N_24853);
xnor UO_2498 (O_2498,N_24804,N_24811);
nor UO_2499 (O_2499,N_24953,N_24921);
xor UO_2500 (O_2500,N_24929,N_24863);
nor UO_2501 (O_2501,N_24832,N_24811);
xor UO_2502 (O_2502,N_24901,N_24875);
xor UO_2503 (O_2503,N_24830,N_24889);
nand UO_2504 (O_2504,N_24858,N_24863);
nor UO_2505 (O_2505,N_24860,N_24938);
xor UO_2506 (O_2506,N_24927,N_24846);
nand UO_2507 (O_2507,N_24964,N_24940);
and UO_2508 (O_2508,N_24915,N_24873);
xnor UO_2509 (O_2509,N_24866,N_24990);
nor UO_2510 (O_2510,N_24998,N_24860);
nand UO_2511 (O_2511,N_24893,N_24902);
nand UO_2512 (O_2512,N_24935,N_24867);
and UO_2513 (O_2513,N_24866,N_24807);
and UO_2514 (O_2514,N_24877,N_24910);
and UO_2515 (O_2515,N_24911,N_24887);
nand UO_2516 (O_2516,N_24849,N_24824);
and UO_2517 (O_2517,N_24898,N_24937);
nor UO_2518 (O_2518,N_24810,N_24825);
xnor UO_2519 (O_2519,N_24842,N_24834);
and UO_2520 (O_2520,N_24812,N_24829);
nor UO_2521 (O_2521,N_24937,N_24941);
xor UO_2522 (O_2522,N_24809,N_24864);
xor UO_2523 (O_2523,N_24897,N_24831);
or UO_2524 (O_2524,N_24900,N_24909);
and UO_2525 (O_2525,N_24972,N_24872);
or UO_2526 (O_2526,N_24999,N_24882);
and UO_2527 (O_2527,N_24966,N_24985);
and UO_2528 (O_2528,N_24915,N_24869);
nand UO_2529 (O_2529,N_24899,N_24826);
nor UO_2530 (O_2530,N_24895,N_24921);
and UO_2531 (O_2531,N_24801,N_24981);
xnor UO_2532 (O_2532,N_24969,N_24958);
nand UO_2533 (O_2533,N_24800,N_24865);
and UO_2534 (O_2534,N_24879,N_24939);
xnor UO_2535 (O_2535,N_24878,N_24811);
or UO_2536 (O_2536,N_24985,N_24999);
and UO_2537 (O_2537,N_24910,N_24911);
nand UO_2538 (O_2538,N_24882,N_24940);
nand UO_2539 (O_2539,N_24905,N_24910);
xnor UO_2540 (O_2540,N_24939,N_24810);
and UO_2541 (O_2541,N_24826,N_24928);
and UO_2542 (O_2542,N_24929,N_24808);
nor UO_2543 (O_2543,N_24910,N_24979);
nor UO_2544 (O_2544,N_24876,N_24974);
nand UO_2545 (O_2545,N_24863,N_24932);
nand UO_2546 (O_2546,N_24809,N_24901);
xor UO_2547 (O_2547,N_24882,N_24808);
xnor UO_2548 (O_2548,N_24956,N_24890);
and UO_2549 (O_2549,N_24917,N_24892);
or UO_2550 (O_2550,N_24857,N_24907);
nor UO_2551 (O_2551,N_24802,N_24862);
and UO_2552 (O_2552,N_24995,N_24963);
or UO_2553 (O_2553,N_24819,N_24841);
xnor UO_2554 (O_2554,N_24800,N_24891);
and UO_2555 (O_2555,N_24810,N_24988);
or UO_2556 (O_2556,N_24868,N_24851);
or UO_2557 (O_2557,N_24992,N_24990);
xor UO_2558 (O_2558,N_24867,N_24885);
and UO_2559 (O_2559,N_24884,N_24903);
nor UO_2560 (O_2560,N_24890,N_24950);
nand UO_2561 (O_2561,N_24879,N_24933);
nor UO_2562 (O_2562,N_24807,N_24805);
nor UO_2563 (O_2563,N_24861,N_24942);
xor UO_2564 (O_2564,N_24924,N_24915);
xnor UO_2565 (O_2565,N_24886,N_24902);
or UO_2566 (O_2566,N_24896,N_24897);
nand UO_2567 (O_2567,N_24937,N_24913);
nand UO_2568 (O_2568,N_24838,N_24825);
nand UO_2569 (O_2569,N_24859,N_24979);
nand UO_2570 (O_2570,N_24853,N_24930);
and UO_2571 (O_2571,N_24895,N_24977);
or UO_2572 (O_2572,N_24833,N_24915);
xnor UO_2573 (O_2573,N_24880,N_24985);
nand UO_2574 (O_2574,N_24990,N_24968);
or UO_2575 (O_2575,N_24832,N_24853);
and UO_2576 (O_2576,N_24840,N_24902);
or UO_2577 (O_2577,N_24926,N_24902);
and UO_2578 (O_2578,N_24901,N_24905);
nand UO_2579 (O_2579,N_24836,N_24850);
nand UO_2580 (O_2580,N_24836,N_24911);
or UO_2581 (O_2581,N_24866,N_24868);
or UO_2582 (O_2582,N_24837,N_24966);
and UO_2583 (O_2583,N_24804,N_24843);
or UO_2584 (O_2584,N_24941,N_24825);
or UO_2585 (O_2585,N_24897,N_24857);
xor UO_2586 (O_2586,N_24925,N_24976);
or UO_2587 (O_2587,N_24828,N_24955);
xor UO_2588 (O_2588,N_24836,N_24881);
nand UO_2589 (O_2589,N_24960,N_24925);
xor UO_2590 (O_2590,N_24911,N_24829);
or UO_2591 (O_2591,N_24833,N_24914);
xnor UO_2592 (O_2592,N_24989,N_24828);
and UO_2593 (O_2593,N_24907,N_24933);
or UO_2594 (O_2594,N_24891,N_24922);
or UO_2595 (O_2595,N_24994,N_24869);
or UO_2596 (O_2596,N_24919,N_24932);
nor UO_2597 (O_2597,N_24993,N_24880);
or UO_2598 (O_2598,N_24852,N_24981);
nand UO_2599 (O_2599,N_24894,N_24872);
or UO_2600 (O_2600,N_24856,N_24976);
xor UO_2601 (O_2601,N_24964,N_24944);
nand UO_2602 (O_2602,N_24982,N_24975);
xor UO_2603 (O_2603,N_24822,N_24821);
nand UO_2604 (O_2604,N_24864,N_24901);
nor UO_2605 (O_2605,N_24816,N_24815);
xor UO_2606 (O_2606,N_24837,N_24855);
or UO_2607 (O_2607,N_24970,N_24859);
or UO_2608 (O_2608,N_24988,N_24898);
or UO_2609 (O_2609,N_24805,N_24800);
nor UO_2610 (O_2610,N_24806,N_24991);
nand UO_2611 (O_2611,N_24996,N_24871);
or UO_2612 (O_2612,N_24972,N_24827);
or UO_2613 (O_2613,N_24986,N_24972);
nor UO_2614 (O_2614,N_24845,N_24940);
nand UO_2615 (O_2615,N_24846,N_24893);
nand UO_2616 (O_2616,N_24923,N_24815);
xnor UO_2617 (O_2617,N_24846,N_24978);
nor UO_2618 (O_2618,N_24859,N_24958);
nor UO_2619 (O_2619,N_24936,N_24841);
nor UO_2620 (O_2620,N_24851,N_24921);
nor UO_2621 (O_2621,N_24809,N_24870);
or UO_2622 (O_2622,N_24836,N_24938);
xnor UO_2623 (O_2623,N_24854,N_24803);
nand UO_2624 (O_2624,N_24855,N_24832);
xor UO_2625 (O_2625,N_24861,N_24979);
and UO_2626 (O_2626,N_24851,N_24916);
nor UO_2627 (O_2627,N_24959,N_24842);
xnor UO_2628 (O_2628,N_24936,N_24876);
and UO_2629 (O_2629,N_24853,N_24924);
xor UO_2630 (O_2630,N_24946,N_24942);
nand UO_2631 (O_2631,N_24870,N_24847);
xnor UO_2632 (O_2632,N_24869,N_24849);
and UO_2633 (O_2633,N_24944,N_24934);
xor UO_2634 (O_2634,N_24840,N_24849);
and UO_2635 (O_2635,N_24894,N_24917);
or UO_2636 (O_2636,N_24915,N_24880);
xnor UO_2637 (O_2637,N_24921,N_24842);
and UO_2638 (O_2638,N_24866,N_24884);
or UO_2639 (O_2639,N_24965,N_24890);
xor UO_2640 (O_2640,N_24831,N_24893);
or UO_2641 (O_2641,N_24995,N_24858);
and UO_2642 (O_2642,N_24962,N_24908);
xor UO_2643 (O_2643,N_24809,N_24937);
and UO_2644 (O_2644,N_24844,N_24849);
nand UO_2645 (O_2645,N_24807,N_24877);
and UO_2646 (O_2646,N_24928,N_24802);
nor UO_2647 (O_2647,N_24848,N_24920);
nand UO_2648 (O_2648,N_24889,N_24803);
and UO_2649 (O_2649,N_24924,N_24872);
or UO_2650 (O_2650,N_24871,N_24856);
nand UO_2651 (O_2651,N_24851,N_24890);
and UO_2652 (O_2652,N_24909,N_24810);
xnor UO_2653 (O_2653,N_24945,N_24824);
and UO_2654 (O_2654,N_24822,N_24804);
nor UO_2655 (O_2655,N_24895,N_24804);
nor UO_2656 (O_2656,N_24873,N_24994);
nor UO_2657 (O_2657,N_24991,N_24843);
xor UO_2658 (O_2658,N_24953,N_24984);
nor UO_2659 (O_2659,N_24809,N_24898);
nor UO_2660 (O_2660,N_24873,N_24941);
and UO_2661 (O_2661,N_24953,N_24950);
and UO_2662 (O_2662,N_24869,N_24964);
nor UO_2663 (O_2663,N_24857,N_24855);
nor UO_2664 (O_2664,N_24854,N_24980);
or UO_2665 (O_2665,N_24883,N_24920);
xnor UO_2666 (O_2666,N_24908,N_24914);
or UO_2667 (O_2667,N_24981,N_24804);
or UO_2668 (O_2668,N_24957,N_24929);
nor UO_2669 (O_2669,N_24980,N_24900);
nor UO_2670 (O_2670,N_24977,N_24909);
and UO_2671 (O_2671,N_24832,N_24986);
xor UO_2672 (O_2672,N_24860,N_24835);
nand UO_2673 (O_2673,N_24993,N_24853);
and UO_2674 (O_2674,N_24928,N_24885);
or UO_2675 (O_2675,N_24874,N_24835);
or UO_2676 (O_2676,N_24944,N_24900);
and UO_2677 (O_2677,N_24980,N_24848);
xnor UO_2678 (O_2678,N_24983,N_24844);
or UO_2679 (O_2679,N_24829,N_24923);
nand UO_2680 (O_2680,N_24953,N_24814);
and UO_2681 (O_2681,N_24960,N_24832);
xnor UO_2682 (O_2682,N_24844,N_24842);
nand UO_2683 (O_2683,N_24895,N_24976);
nor UO_2684 (O_2684,N_24931,N_24877);
and UO_2685 (O_2685,N_24900,N_24804);
and UO_2686 (O_2686,N_24810,N_24803);
nor UO_2687 (O_2687,N_24840,N_24809);
and UO_2688 (O_2688,N_24997,N_24860);
nor UO_2689 (O_2689,N_24928,N_24936);
xor UO_2690 (O_2690,N_24965,N_24852);
or UO_2691 (O_2691,N_24893,N_24828);
nor UO_2692 (O_2692,N_24936,N_24866);
or UO_2693 (O_2693,N_24965,N_24903);
and UO_2694 (O_2694,N_24941,N_24819);
xor UO_2695 (O_2695,N_24952,N_24967);
nor UO_2696 (O_2696,N_24903,N_24912);
nand UO_2697 (O_2697,N_24823,N_24827);
xor UO_2698 (O_2698,N_24847,N_24839);
nor UO_2699 (O_2699,N_24859,N_24974);
nand UO_2700 (O_2700,N_24860,N_24975);
nand UO_2701 (O_2701,N_24864,N_24953);
or UO_2702 (O_2702,N_24993,N_24991);
nand UO_2703 (O_2703,N_24891,N_24828);
nor UO_2704 (O_2704,N_24913,N_24961);
nand UO_2705 (O_2705,N_24903,N_24868);
xnor UO_2706 (O_2706,N_24902,N_24992);
xor UO_2707 (O_2707,N_24992,N_24998);
nor UO_2708 (O_2708,N_24811,N_24933);
nor UO_2709 (O_2709,N_24865,N_24884);
nand UO_2710 (O_2710,N_24989,N_24843);
nand UO_2711 (O_2711,N_24912,N_24908);
or UO_2712 (O_2712,N_24898,N_24814);
or UO_2713 (O_2713,N_24878,N_24957);
nand UO_2714 (O_2714,N_24807,N_24999);
xnor UO_2715 (O_2715,N_24883,N_24983);
nand UO_2716 (O_2716,N_24813,N_24955);
nand UO_2717 (O_2717,N_24826,N_24896);
nor UO_2718 (O_2718,N_24959,N_24815);
xor UO_2719 (O_2719,N_24819,N_24957);
xnor UO_2720 (O_2720,N_24992,N_24819);
nor UO_2721 (O_2721,N_24874,N_24899);
and UO_2722 (O_2722,N_24846,N_24869);
xnor UO_2723 (O_2723,N_24982,N_24865);
xnor UO_2724 (O_2724,N_24873,N_24967);
xor UO_2725 (O_2725,N_24836,N_24803);
nor UO_2726 (O_2726,N_24933,N_24882);
and UO_2727 (O_2727,N_24925,N_24894);
nand UO_2728 (O_2728,N_24964,N_24864);
or UO_2729 (O_2729,N_24829,N_24932);
xor UO_2730 (O_2730,N_24973,N_24829);
nor UO_2731 (O_2731,N_24897,N_24839);
or UO_2732 (O_2732,N_24925,N_24907);
or UO_2733 (O_2733,N_24975,N_24965);
and UO_2734 (O_2734,N_24846,N_24907);
and UO_2735 (O_2735,N_24903,N_24981);
xor UO_2736 (O_2736,N_24873,N_24842);
nor UO_2737 (O_2737,N_24868,N_24933);
or UO_2738 (O_2738,N_24830,N_24832);
nor UO_2739 (O_2739,N_24835,N_24833);
xnor UO_2740 (O_2740,N_24859,N_24935);
xnor UO_2741 (O_2741,N_24886,N_24816);
xnor UO_2742 (O_2742,N_24952,N_24995);
nor UO_2743 (O_2743,N_24950,N_24919);
xor UO_2744 (O_2744,N_24931,N_24842);
and UO_2745 (O_2745,N_24958,N_24915);
nor UO_2746 (O_2746,N_24977,N_24822);
or UO_2747 (O_2747,N_24969,N_24953);
or UO_2748 (O_2748,N_24930,N_24952);
nand UO_2749 (O_2749,N_24959,N_24828);
or UO_2750 (O_2750,N_24847,N_24895);
nand UO_2751 (O_2751,N_24928,N_24860);
or UO_2752 (O_2752,N_24864,N_24825);
nor UO_2753 (O_2753,N_24910,N_24973);
nand UO_2754 (O_2754,N_24828,N_24899);
nor UO_2755 (O_2755,N_24928,N_24915);
nor UO_2756 (O_2756,N_24997,N_24817);
or UO_2757 (O_2757,N_24947,N_24964);
and UO_2758 (O_2758,N_24931,N_24883);
nor UO_2759 (O_2759,N_24892,N_24951);
xor UO_2760 (O_2760,N_24838,N_24860);
and UO_2761 (O_2761,N_24864,N_24945);
and UO_2762 (O_2762,N_24928,N_24987);
nor UO_2763 (O_2763,N_24960,N_24909);
nor UO_2764 (O_2764,N_24884,N_24874);
nand UO_2765 (O_2765,N_24874,N_24819);
and UO_2766 (O_2766,N_24850,N_24885);
and UO_2767 (O_2767,N_24923,N_24956);
nand UO_2768 (O_2768,N_24812,N_24924);
and UO_2769 (O_2769,N_24823,N_24928);
or UO_2770 (O_2770,N_24900,N_24910);
nand UO_2771 (O_2771,N_24921,N_24960);
xnor UO_2772 (O_2772,N_24992,N_24978);
or UO_2773 (O_2773,N_24837,N_24967);
nor UO_2774 (O_2774,N_24835,N_24915);
and UO_2775 (O_2775,N_24984,N_24851);
and UO_2776 (O_2776,N_24948,N_24851);
nand UO_2777 (O_2777,N_24914,N_24896);
xor UO_2778 (O_2778,N_24876,N_24953);
and UO_2779 (O_2779,N_24865,N_24816);
nand UO_2780 (O_2780,N_24912,N_24808);
nor UO_2781 (O_2781,N_24889,N_24990);
xor UO_2782 (O_2782,N_24881,N_24813);
xnor UO_2783 (O_2783,N_24980,N_24915);
nand UO_2784 (O_2784,N_24820,N_24835);
xnor UO_2785 (O_2785,N_24827,N_24836);
xor UO_2786 (O_2786,N_24897,N_24835);
or UO_2787 (O_2787,N_24827,N_24906);
nand UO_2788 (O_2788,N_24976,N_24978);
and UO_2789 (O_2789,N_24880,N_24887);
and UO_2790 (O_2790,N_24918,N_24997);
nor UO_2791 (O_2791,N_24926,N_24843);
or UO_2792 (O_2792,N_24942,N_24879);
xnor UO_2793 (O_2793,N_24813,N_24939);
or UO_2794 (O_2794,N_24970,N_24950);
and UO_2795 (O_2795,N_24901,N_24941);
nor UO_2796 (O_2796,N_24812,N_24914);
xor UO_2797 (O_2797,N_24952,N_24874);
nand UO_2798 (O_2798,N_24843,N_24818);
nand UO_2799 (O_2799,N_24887,N_24996);
or UO_2800 (O_2800,N_24828,N_24879);
nand UO_2801 (O_2801,N_24879,N_24966);
nand UO_2802 (O_2802,N_24851,N_24998);
and UO_2803 (O_2803,N_24867,N_24843);
xor UO_2804 (O_2804,N_24853,N_24935);
or UO_2805 (O_2805,N_24851,N_24869);
and UO_2806 (O_2806,N_24810,N_24958);
or UO_2807 (O_2807,N_24983,N_24896);
or UO_2808 (O_2808,N_24953,N_24914);
nand UO_2809 (O_2809,N_24934,N_24826);
nor UO_2810 (O_2810,N_24988,N_24896);
and UO_2811 (O_2811,N_24878,N_24905);
nor UO_2812 (O_2812,N_24885,N_24863);
or UO_2813 (O_2813,N_24981,N_24870);
xnor UO_2814 (O_2814,N_24866,N_24839);
nand UO_2815 (O_2815,N_24883,N_24865);
and UO_2816 (O_2816,N_24985,N_24987);
or UO_2817 (O_2817,N_24954,N_24881);
or UO_2818 (O_2818,N_24888,N_24951);
nand UO_2819 (O_2819,N_24822,N_24965);
or UO_2820 (O_2820,N_24977,N_24979);
nand UO_2821 (O_2821,N_24988,N_24978);
xor UO_2822 (O_2822,N_24909,N_24955);
xnor UO_2823 (O_2823,N_24955,N_24848);
nand UO_2824 (O_2824,N_24930,N_24872);
and UO_2825 (O_2825,N_24815,N_24952);
or UO_2826 (O_2826,N_24838,N_24939);
nand UO_2827 (O_2827,N_24987,N_24976);
or UO_2828 (O_2828,N_24972,N_24851);
nand UO_2829 (O_2829,N_24917,N_24818);
nand UO_2830 (O_2830,N_24893,N_24835);
and UO_2831 (O_2831,N_24889,N_24845);
and UO_2832 (O_2832,N_24866,N_24837);
nand UO_2833 (O_2833,N_24999,N_24885);
or UO_2834 (O_2834,N_24842,N_24988);
nor UO_2835 (O_2835,N_24819,N_24806);
xor UO_2836 (O_2836,N_24949,N_24836);
nand UO_2837 (O_2837,N_24858,N_24920);
xor UO_2838 (O_2838,N_24822,N_24806);
and UO_2839 (O_2839,N_24958,N_24839);
xor UO_2840 (O_2840,N_24846,N_24854);
nand UO_2841 (O_2841,N_24941,N_24938);
or UO_2842 (O_2842,N_24835,N_24828);
and UO_2843 (O_2843,N_24959,N_24937);
or UO_2844 (O_2844,N_24989,N_24919);
xnor UO_2845 (O_2845,N_24981,N_24937);
xnor UO_2846 (O_2846,N_24828,N_24905);
and UO_2847 (O_2847,N_24938,N_24905);
or UO_2848 (O_2848,N_24986,N_24962);
and UO_2849 (O_2849,N_24941,N_24844);
xnor UO_2850 (O_2850,N_24827,N_24832);
xnor UO_2851 (O_2851,N_24852,N_24990);
or UO_2852 (O_2852,N_24903,N_24880);
or UO_2853 (O_2853,N_24894,N_24895);
and UO_2854 (O_2854,N_24815,N_24852);
and UO_2855 (O_2855,N_24841,N_24888);
or UO_2856 (O_2856,N_24809,N_24972);
xor UO_2857 (O_2857,N_24872,N_24925);
nand UO_2858 (O_2858,N_24987,N_24977);
or UO_2859 (O_2859,N_24996,N_24947);
or UO_2860 (O_2860,N_24851,N_24826);
or UO_2861 (O_2861,N_24889,N_24863);
xnor UO_2862 (O_2862,N_24977,N_24873);
nand UO_2863 (O_2863,N_24881,N_24883);
xnor UO_2864 (O_2864,N_24871,N_24839);
and UO_2865 (O_2865,N_24955,N_24812);
nand UO_2866 (O_2866,N_24951,N_24992);
xnor UO_2867 (O_2867,N_24971,N_24969);
nand UO_2868 (O_2868,N_24954,N_24967);
or UO_2869 (O_2869,N_24851,N_24915);
nor UO_2870 (O_2870,N_24915,N_24839);
and UO_2871 (O_2871,N_24888,N_24818);
or UO_2872 (O_2872,N_24869,N_24987);
xnor UO_2873 (O_2873,N_24967,N_24901);
xnor UO_2874 (O_2874,N_24818,N_24971);
xor UO_2875 (O_2875,N_24827,N_24913);
nor UO_2876 (O_2876,N_24862,N_24816);
and UO_2877 (O_2877,N_24923,N_24844);
xor UO_2878 (O_2878,N_24988,N_24977);
nand UO_2879 (O_2879,N_24876,N_24946);
or UO_2880 (O_2880,N_24817,N_24823);
or UO_2881 (O_2881,N_24868,N_24881);
and UO_2882 (O_2882,N_24853,N_24937);
nand UO_2883 (O_2883,N_24970,N_24831);
xor UO_2884 (O_2884,N_24938,N_24875);
xnor UO_2885 (O_2885,N_24979,N_24891);
and UO_2886 (O_2886,N_24901,N_24857);
xnor UO_2887 (O_2887,N_24920,N_24843);
or UO_2888 (O_2888,N_24825,N_24800);
nor UO_2889 (O_2889,N_24942,N_24941);
or UO_2890 (O_2890,N_24876,N_24812);
nor UO_2891 (O_2891,N_24894,N_24868);
xor UO_2892 (O_2892,N_24867,N_24903);
or UO_2893 (O_2893,N_24887,N_24899);
nor UO_2894 (O_2894,N_24940,N_24899);
nor UO_2895 (O_2895,N_24867,N_24980);
nor UO_2896 (O_2896,N_24996,N_24932);
nand UO_2897 (O_2897,N_24852,N_24903);
and UO_2898 (O_2898,N_24824,N_24887);
nor UO_2899 (O_2899,N_24990,N_24855);
xor UO_2900 (O_2900,N_24831,N_24978);
or UO_2901 (O_2901,N_24993,N_24882);
or UO_2902 (O_2902,N_24946,N_24842);
xnor UO_2903 (O_2903,N_24904,N_24955);
or UO_2904 (O_2904,N_24862,N_24861);
xnor UO_2905 (O_2905,N_24859,N_24928);
and UO_2906 (O_2906,N_24923,N_24965);
or UO_2907 (O_2907,N_24906,N_24967);
nand UO_2908 (O_2908,N_24824,N_24937);
xor UO_2909 (O_2909,N_24999,N_24921);
nand UO_2910 (O_2910,N_24952,N_24826);
xor UO_2911 (O_2911,N_24907,N_24931);
or UO_2912 (O_2912,N_24911,N_24918);
nand UO_2913 (O_2913,N_24826,N_24855);
or UO_2914 (O_2914,N_24834,N_24885);
xnor UO_2915 (O_2915,N_24938,N_24886);
nand UO_2916 (O_2916,N_24895,N_24980);
or UO_2917 (O_2917,N_24847,N_24924);
xnor UO_2918 (O_2918,N_24911,N_24944);
nor UO_2919 (O_2919,N_24919,N_24841);
xnor UO_2920 (O_2920,N_24838,N_24814);
or UO_2921 (O_2921,N_24826,N_24804);
xor UO_2922 (O_2922,N_24846,N_24956);
nand UO_2923 (O_2923,N_24853,N_24835);
and UO_2924 (O_2924,N_24956,N_24971);
and UO_2925 (O_2925,N_24809,N_24819);
nor UO_2926 (O_2926,N_24950,N_24915);
or UO_2927 (O_2927,N_24803,N_24830);
xnor UO_2928 (O_2928,N_24905,N_24974);
and UO_2929 (O_2929,N_24843,N_24939);
nor UO_2930 (O_2930,N_24952,N_24931);
and UO_2931 (O_2931,N_24837,N_24928);
nand UO_2932 (O_2932,N_24993,N_24870);
xor UO_2933 (O_2933,N_24820,N_24889);
nand UO_2934 (O_2934,N_24828,N_24871);
xor UO_2935 (O_2935,N_24855,N_24912);
xnor UO_2936 (O_2936,N_24923,N_24929);
and UO_2937 (O_2937,N_24974,N_24961);
nor UO_2938 (O_2938,N_24815,N_24857);
and UO_2939 (O_2939,N_24954,N_24829);
nor UO_2940 (O_2940,N_24994,N_24876);
nand UO_2941 (O_2941,N_24839,N_24811);
nand UO_2942 (O_2942,N_24940,N_24993);
nor UO_2943 (O_2943,N_24904,N_24880);
or UO_2944 (O_2944,N_24981,N_24811);
nor UO_2945 (O_2945,N_24912,N_24913);
nand UO_2946 (O_2946,N_24835,N_24990);
and UO_2947 (O_2947,N_24958,N_24995);
and UO_2948 (O_2948,N_24998,N_24827);
or UO_2949 (O_2949,N_24886,N_24977);
xnor UO_2950 (O_2950,N_24878,N_24846);
xnor UO_2951 (O_2951,N_24862,N_24874);
or UO_2952 (O_2952,N_24999,N_24980);
and UO_2953 (O_2953,N_24808,N_24818);
xnor UO_2954 (O_2954,N_24815,N_24842);
nand UO_2955 (O_2955,N_24897,N_24963);
nand UO_2956 (O_2956,N_24881,N_24906);
and UO_2957 (O_2957,N_24833,N_24894);
nor UO_2958 (O_2958,N_24867,N_24870);
xor UO_2959 (O_2959,N_24960,N_24811);
and UO_2960 (O_2960,N_24962,N_24871);
xnor UO_2961 (O_2961,N_24872,N_24866);
or UO_2962 (O_2962,N_24894,N_24900);
and UO_2963 (O_2963,N_24861,N_24958);
and UO_2964 (O_2964,N_24982,N_24870);
xnor UO_2965 (O_2965,N_24908,N_24877);
or UO_2966 (O_2966,N_24838,N_24878);
or UO_2967 (O_2967,N_24969,N_24947);
nor UO_2968 (O_2968,N_24970,N_24828);
or UO_2969 (O_2969,N_24837,N_24961);
or UO_2970 (O_2970,N_24984,N_24874);
or UO_2971 (O_2971,N_24985,N_24993);
xor UO_2972 (O_2972,N_24803,N_24914);
nand UO_2973 (O_2973,N_24831,N_24847);
nor UO_2974 (O_2974,N_24968,N_24868);
xor UO_2975 (O_2975,N_24827,N_24990);
xnor UO_2976 (O_2976,N_24966,N_24804);
nor UO_2977 (O_2977,N_24812,N_24980);
nand UO_2978 (O_2978,N_24880,N_24949);
and UO_2979 (O_2979,N_24914,N_24931);
nor UO_2980 (O_2980,N_24897,N_24817);
or UO_2981 (O_2981,N_24815,N_24941);
nand UO_2982 (O_2982,N_24801,N_24845);
nand UO_2983 (O_2983,N_24858,N_24993);
and UO_2984 (O_2984,N_24817,N_24814);
nand UO_2985 (O_2985,N_24993,N_24911);
xor UO_2986 (O_2986,N_24852,N_24881);
or UO_2987 (O_2987,N_24804,N_24922);
nor UO_2988 (O_2988,N_24900,N_24971);
xnor UO_2989 (O_2989,N_24982,N_24823);
nand UO_2990 (O_2990,N_24903,N_24817);
and UO_2991 (O_2991,N_24901,N_24882);
xnor UO_2992 (O_2992,N_24805,N_24970);
or UO_2993 (O_2993,N_24802,N_24888);
or UO_2994 (O_2994,N_24915,N_24995);
nand UO_2995 (O_2995,N_24815,N_24927);
or UO_2996 (O_2996,N_24844,N_24855);
xnor UO_2997 (O_2997,N_24806,N_24817);
or UO_2998 (O_2998,N_24913,N_24846);
xnor UO_2999 (O_2999,N_24857,N_24847);
endmodule