module basic_2500_25000_3000_20_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_137,In_1322);
nand U1 (N_1,In_425,In_1718);
nor U2 (N_2,In_742,In_988);
xnor U3 (N_3,In_284,In_1871);
and U4 (N_4,In_915,In_2248);
and U5 (N_5,In_1558,In_153);
or U6 (N_6,In_737,In_264);
nor U7 (N_7,In_1764,In_1228);
nand U8 (N_8,In_1373,In_1496);
nand U9 (N_9,In_2051,In_99);
and U10 (N_10,In_50,In_1732);
nor U11 (N_11,In_1946,In_777);
and U12 (N_12,In_75,In_40);
xor U13 (N_13,In_1502,In_2155);
nand U14 (N_14,In_1619,In_1746);
or U15 (N_15,In_800,In_1484);
nand U16 (N_16,In_2181,In_1021);
nor U17 (N_17,In_1741,In_2230);
nand U18 (N_18,In_1109,In_1375);
and U19 (N_19,In_1638,In_353);
or U20 (N_20,In_1213,In_1684);
and U21 (N_21,In_205,In_1955);
nand U22 (N_22,In_2396,In_799);
nand U23 (N_23,In_1574,In_1167);
and U24 (N_24,In_1550,In_1782);
nor U25 (N_25,In_2351,In_2428);
xnor U26 (N_26,In_1355,In_2385);
and U27 (N_27,In_758,In_1399);
and U28 (N_28,In_2427,In_1145);
nand U29 (N_29,In_190,In_1847);
and U30 (N_30,In_1194,In_1664);
or U31 (N_31,In_1873,In_2370);
and U32 (N_32,In_2134,In_1293);
nand U33 (N_33,In_1261,In_1328);
or U34 (N_34,In_885,In_1263);
nor U35 (N_35,In_1757,In_1608);
and U36 (N_36,In_862,In_1295);
nand U37 (N_37,In_453,In_790);
and U38 (N_38,In_1111,In_2380);
nand U39 (N_39,In_1158,In_402);
and U40 (N_40,In_2093,In_8);
nor U41 (N_41,In_2465,In_388);
xnor U42 (N_42,In_407,In_797);
nor U43 (N_43,In_439,In_1609);
nor U44 (N_44,In_1846,In_950);
or U45 (N_45,In_516,In_2384);
or U46 (N_46,In_1792,In_1233);
nand U47 (N_47,In_2106,In_376);
xnor U48 (N_48,In_1205,In_2116);
nand U49 (N_49,In_1105,In_1093);
nor U50 (N_50,In_766,In_1660);
and U51 (N_51,In_515,In_1441);
and U52 (N_52,In_2124,In_440);
nor U53 (N_53,In_1788,In_1505);
xnor U54 (N_54,In_47,In_1382);
and U55 (N_55,In_1709,In_143);
nand U56 (N_56,In_1379,In_1269);
nor U57 (N_57,In_37,In_2392);
xnor U58 (N_58,In_1602,In_1273);
and U59 (N_59,In_1420,In_612);
xnor U60 (N_60,In_106,In_1138);
nand U61 (N_61,In_1125,In_923);
or U62 (N_62,In_1942,In_2343);
and U63 (N_63,In_1738,In_2444);
or U64 (N_64,In_2300,In_2405);
and U65 (N_65,In_1115,In_452);
or U66 (N_66,In_17,In_1945);
xor U67 (N_67,In_698,In_282);
and U68 (N_68,In_1665,In_1548);
or U69 (N_69,In_1011,In_88);
xor U70 (N_70,In_151,In_545);
or U71 (N_71,In_1223,In_464);
and U72 (N_72,In_721,In_2252);
or U73 (N_73,In_1606,In_405);
xnor U74 (N_74,In_1041,In_20);
and U75 (N_75,In_1249,In_581);
xor U76 (N_76,In_1311,In_932);
xor U77 (N_77,In_2060,In_2157);
and U78 (N_78,In_100,In_551);
xor U79 (N_79,In_772,In_798);
xnor U80 (N_80,In_2467,In_1837);
nand U81 (N_81,In_2306,In_842);
and U82 (N_82,In_1830,In_716);
xor U83 (N_83,In_2057,In_1381);
and U84 (N_84,In_292,In_171);
xor U85 (N_85,In_29,In_658);
nand U86 (N_86,In_2175,In_1226);
or U87 (N_87,In_2113,In_1380);
nand U88 (N_88,In_1095,In_277);
or U89 (N_89,In_228,In_528);
nand U90 (N_90,In_2286,In_1767);
nand U91 (N_91,In_1467,In_96);
xnor U92 (N_92,In_2218,In_601);
xor U93 (N_93,In_470,In_1979);
nor U94 (N_94,In_499,In_1482);
nor U95 (N_95,In_2091,In_332);
and U96 (N_96,In_2419,In_1691);
or U97 (N_97,In_557,In_2043);
nand U98 (N_98,In_1928,In_141);
nor U99 (N_99,In_2247,In_1722);
nand U100 (N_100,In_616,In_2037);
nor U101 (N_101,In_2455,In_1985);
nor U102 (N_102,In_1214,In_669);
nand U103 (N_103,In_638,In_1986);
xnor U104 (N_104,In_403,In_1279);
nor U105 (N_105,In_1806,In_1840);
and U106 (N_106,In_1219,In_261);
xor U107 (N_107,In_496,In_1939);
xor U108 (N_108,In_2470,In_2110);
and U109 (N_109,In_1057,In_87);
nand U110 (N_110,In_2180,In_1156);
xnor U111 (N_111,In_1256,In_1298);
and U112 (N_112,In_1912,In_314);
or U113 (N_113,In_2259,In_1737);
xor U114 (N_114,In_1045,In_1504);
or U115 (N_115,In_1130,In_2479);
nand U116 (N_116,In_34,In_1875);
nand U117 (N_117,In_637,In_1013);
nand U118 (N_118,In_1824,In_2459);
xnor U119 (N_119,In_1934,In_2061);
xnor U120 (N_120,In_172,In_691);
and U121 (N_121,In_209,In_286);
xnor U122 (N_122,In_629,In_1405);
xor U123 (N_123,In_523,In_1348);
and U124 (N_124,In_1758,In_849);
nor U125 (N_125,In_163,In_665);
nand U126 (N_126,In_446,In_935);
and U127 (N_127,In_572,In_1462);
or U128 (N_128,In_1176,In_2219);
or U129 (N_129,In_155,In_1769);
or U130 (N_130,In_2012,In_2242);
and U131 (N_131,In_2152,In_2194);
nand U132 (N_132,In_1535,In_951);
nand U133 (N_133,In_2197,In_834);
xnor U134 (N_134,In_1828,In_483);
nand U135 (N_135,In_929,In_2413);
xor U136 (N_136,In_53,In_1687);
or U137 (N_137,In_2112,In_1612);
and U138 (N_138,In_904,In_1804);
xor U139 (N_139,In_1181,In_1644);
nor U140 (N_140,In_1007,In_896);
and U141 (N_141,In_1540,In_160);
or U142 (N_142,In_2067,In_1353);
xor U143 (N_143,In_1489,In_2289);
and U144 (N_144,In_1345,In_2406);
nor U145 (N_145,In_450,In_2096);
xor U146 (N_146,In_1523,In_2222);
and U147 (N_147,In_9,In_1452);
xnor U148 (N_148,In_433,In_1493);
xor U149 (N_149,In_1440,In_2358);
and U150 (N_150,In_1090,In_1036);
nand U151 (N_151,In_1605,In_760);
or U152 (N_152,In_956,In_930);
nor U153 (N_153,In_2034,In_1186);
nand U154 (N_154,In_829,In_838);
and U155 (N_155,In_1437,In_130);
or U156 (N_156,In_1162,In_193);
or U157 (N_157,In_1259,In_1067);
xor U158 (N_158,In_1598,In_1336);
xor U159 (N_159,In_2210,In_2365);
nor U160 (N_160,In_181,In_1062);
or U161 (N_161,In_1187,In_1189);
and U162 (N_162,In_531,In_196);
and U163 (N_163,In_1142,In_2065);
nor U164 (N_164,In_1997,In_2327);
xor U165 (N_165,In_2402,In_1981);
or U166 (N_166,In_1819,In_1394);
nor U167 (N_167,In_497,In_2310);
xnor U168 (N_168,In_2308,In_1087);
and U169 (N_169,In_444,In_2466);
or U170 (N_170,In_1246,In_1335);
and U171 (N_171,In_1887,In_1675);
xor U172 (N_172,In_1290,In_438);
and U173 (N_173,In_415,In_273);
and U174 (N_174,In_1584,In_586);
xnor U175 (N_175,In_482,In_848);
and U176 (N_176,In_2480,In_13);
or U177 (N_177,In_199,In_189);
nor U178 (N_178,In_1422,In_2148);
or U179 (N_179,In_1610,In_2364);
or U180 (N_180,In_1049,In_379);
nand U181 (N_181,In_1628,In_754);
or U182 (N_182,In_1747,In_875);
nand U183 (N_183,In_469,In_2332);
or U184 (N_184,In_2042,In_856);
nand U185 (N_185,In_119,In_1245);
nor U186 (N_186,In_890,In_471);
and U187 (N_187,In_144,In_1427);
or U188 (N_188,In_2225,In_145);
or U189 (N_189,In_931,In_2277);
nand U190 (N_190,In_413,In_1351);
nor U191 (N_191,In_1250,In_2378);
and U192 (N_192,In_2131,In_1369);
nand U193 (N_193,In_169,In_957);
nand U194 (N_194,In_27,In_533);
nand U195 (N_195,In_1106,In_818);
and U196 (N_196,In_136,In_1310);
nor U197 (N_197,In_301,In_142);
nor U198 (N_198,In_1877,In_1292);
nor U199 (N_199,In_1640,In_1302);
xnor U200 (N_200,In_632,In_969);
or U201 (N_201,In_934,In_2062);
nor U202 (N_202,In_973,In_2135);
nor U203 (N_203,In_1796,In_580);
nand U204 (N_204,In_435,In_2346);
and U205 (N_205,In_2064,In_2420);
nor U206 (N_206,In_1148,In_1719);
nand U207 (N_207,In_63,In_1658);
nor U208 (N_208,In_1038,In_788);
or U209 (N_209,In_2321,In_1274);
or U210 (N_210,In_786,In_1066);
and U211 (N_211,In_2301,In_692);
nand U212 (N_212,In_204,In_2019);
nand U213 (N_213,In_1135,In_1994);
or U214 (N_214,In_317,In_426);
or U215 (N_215,In_1697,In_318);
and U216 (N_216,In_600,In_1593);
nand U217 (N_217,In_245,In_307);
nor U218 (N_218,In_1305,In_1672);
nor U219 (N_219,In_1413,In_1973);
nand U220 (N_220,In_1688,In_152);
or U221 (N_221,In_1490,In_903);
xor U222 (N_222,In_720,In_908);
and U223 (N_223,In_2080,In_2446);
nor U224 (N_224,In_837,In_819);
or U225 (N_225,In_2342,In_1461);
or U226 (N_226,In_1825,In_1933);
xnor U227 (N_227,In_1026,In_762);
nor U228 (N_228,In_510,In_2071);
xnor U229 (N_229,In_14,In_752);
nand U230 (N_230,In_2324,In_101);
xnor U231 (N_231,In_1770,In_1277);
or U232 (N_232,In_1588,In_2212);
nor U233 (N_233,In_219,In_239);
xor U234 (N_234,In_1431,In_399);
nand U235 (N_235,In_701,In_1108);
and U236 (N_236,In_371,In_1040);
xnor U237 (N_237,In_955,In_465);
nand U238 (N_238,In_2460,In_2174);
and U239 (N_239,In_1065,In_1301);
nor U240 (N_240,In_1848,In_2383);
xnor U241 (N_241,In_1060,In_1607);
nand U242 (N_242,In_962,In_275);
nor U243 (N_243,In_2429,In_650);
and U244 (N_244,In_2153,In_1029);
nor U245 (N_245,In_1211,In_1362);
and U246 (N_246,In_33,In_180);
nor U247 (N_247,In_2442,In_2317);
nor U248 (N_248,In_356,In_1486);
xnor U249 (N_249,In_237,In_1019);
xnor U250 (N_250,In_197,In_1491);
nor U251 (N_251,In_389,In_125);
nor U252 (N_252,In_921,In_1294);
and U253 (N_253,In_1773,In_1168);
nand U254 (N_254,In_133,In_769);
and U255 (N_255,In_2244,In_2389);
nor U256 (N_256,In_2490,In_1208);
nor U257 (N_257,In_1297,In_649);
or U258 (N_258,In_576,In_984);
nand U259 (N_259,In_128,In_1161);
xnor U260 (N_260,In_392,In_1433);
or U261 (N_261,In_534,In_2350);
nand U262 (N_262,In_2297,In_1350);
nand U263 (N_263,In_467,In_1790);
or U264 (N_264,In_945,In_571);
or U265 (N_265,In_906,In_1339);
and U266 (N_266,In_147,In_1417);
or U267 (N_267,In_1633,In_547);
xnor U268 (N_268,In_2101,In_1567);
and U269 (N_269,In_1701,In_173);
nor U270 (N_270,In_1009,In_905);
nor U271 (N_271,In_2319,In_1935);
nand U272 (N_272,In_595,In_1749);
nand U273 (N_273,In_1814,In_1519);
and U274 (N_274,In_1635,In_607);
nor U275 (N_275,In_1177,In_2224);
nor U276 (N_276,In_2109,In_964);
or U277 (N_277,In_2407,In_641);
and U278 (N_278,In_2246,In_1079);
nand U279 (N_279,In_526,In_1199);
nor U280 (N_280,In_1786,In_1561);
and U281 (N_281,In_2495,In_319);
nand U282 (N_282,In_1833,In_370);
and U283 (N_283,In_430,In_1055);
nand U284 (N_284,In_1894,In_2268);
and U285 (N_285,In_1349,In_2331);
and U286 (N_286,In_946,In_1596);
or U287 (N_287,In_731,In_1240);
xnor U288 (N_288,In_1838,In_1384);
or U289 (N_289,In_1444,In_1175);
or U290 (N_290,In_312,In_993);
xor U291 (N_291,In_1185,In_343);
nand U292 (N_292,In_457,In_1844);
nor U293 (N_293,In_2424,In_605);
nor U294 (N_294,In_1510,In_288);
nor U295 (N_295,In_211,In_1116);
and U296 (N_296,In_363,In_1891);
nand U297 (N_297,In_2438,In_2015);
or U298 (N_298,In_1202,In_255);
nor U299 (N_299,In_191,In_2036);
xor U300 (N_300,In_591,In_1378);
or U301 (N_301,In_566,In_1107);
or U302 (N_302,In_304,In_1617);
nor U303 (N_303,In_1260,In_892);
nand U304 (N_304,In_1153,In_1562);
or U305 (N_305,In_2081,In_1178);
or U306 (N_306,In_744,In_1423);
nor U307 (N_307,In_718,In_7);
nand U308 (N_308,In_556,In_1851);
xnor U309 (N_309,In_1627,In_901);
or U310 (N_310,In_1377,In_2401);
and U311 (N_311,In_1827,In_1793);
nor U312 (N_312,In_1666,In_1603);
or U313 (N_313,In_909,In_1064);
or U314 (N_314,In_778,In_1458);
or U315 (N_315,In_539,In_588);
nor U316 (N_316,In_1629,In_162);
nor U317 (N_317,In_705,In_809);
xnor U318 (N_318,In_2395,In_1892);
and U319 (N_319,In_920,In_2399);
xnor U320 (N_320,In_306,In_815);
xor U321 (N_321,In_1412,In_2341);
nand U322 (N_322,In_1283,In_410);
or U323 (N_323,In_1650,In_1655);
or U324 (N_324,In_958,In_336);
xnor U325 (N_325,In_982,In_661);
xnor U326 (N_326,In_479,In_1266);
xnor U327 (N_327,In_1165,In_573);
nand U328 (N_328,In_224,In_2216);
and U329 (N_329,In_530,In_1795);
xnor U330 (N_330,In_618,In_1716);
or U331 (N_331,In_1210,In_148);
and U332 (N_332,In_1849,In_1959);
xnor U333 (N_333,In_2333,In_400);
or U334 (N_334,In_643,In_1768);
nand U335 (N_335,In_337,In_2262);
or U336 (N_336,In_2498,In_2117);
nand U337 (N_337,In_559,In_996);
xnor U338 (N_338,In_759,In_226);
or U339 (N_339,In_709,In_2323);
nor U340 (N_340,In_899,In_229);
nor U341 (N_341,In_2241,In_803);
and U342 (N_342,In_1068,In_1587);
and U343 (N_343,In_719,In_2398);
and U344 (N_344,In_1906,In_1455);
xor U345 (N_345,In_670,In_1772);
xor U346 (N_346,In_1128,In_2345);
xnor U347 (N_347,In_1112,In_1654);
nor U348 (N_348,In_553,In_1248);
and U349 (N_349,In_188,In_2291);
or U350 (N_350,In_300,In_1204);
and U351 (N_351,In_1229,In_2376);
nand U352 (N_352,In_2488,In_1779);
xnor U353 (N_353,In_1438,In_1101);
or U354 (N_354,In_2257,In_107);
or U355 (N_355,In_478,In_2184);
and U356 (N_356,In_19,In_208);
xnor U357 (N_357,In_913,In_463);
nand U358 (N_358,In_1469,In_174);
or U359 (N_359,In_11,In_1543);
xor U360 (N_360,In_912,In_1957);
and U361 (N_361,In_1341,In_2126);
and U362 (N_362,In_1984,In_1966);
and U363 (N_363,In_1876,In_2469);
and U364 (N_364,In_2176,In_1797);
nor U365 (N_365,In_1626,In_1434);
and U366 (N_366,In_568,In_1308);
xnor U367 (N_367,In_924,In_1418);
nor U368 (N_368,In_1252,In_2140);
xor U369 (N_369,In_10,In_688);
and U370 (N_370,In_213,In_1657);
and U371 (N_371,In_714,In_1338);
nand U372 (N_372,In_1733,In_2235);
nor U373 (N_373,In_1443,In_1542);
nor U374 (N_374,In_1898,In_390);
or U375 (N_375,In_883,In_1332);
or U376 (N_376,In_833,In_2170);
or U377 (N_377,In_1251,In_877);
or U378 (N_378,In_266,In_503);
xnor U379 (N_379,In_960,In_2169);
nand U380 (N_380,In_575,In_717);
nand U381 (N_381,In_448,In_222);
or U382 (N_382,In_2464,In_1030);
xor U383 (N_383,In_2120,In_1344);
or U384 (N_384,In_2136,In_801);
and U385 (N_385,In_990,In_2097);
and U386 (N_386,In_1926,In_6);
xor U387 (N_387,In_2437,In_689);
nor U388 (N_388,In_910,In_216);
xnor U389 (N_389,In_606,In_2021);
nor U390 (N_390,In_1998,In_62);
and U391 (N_391,In_2027,In_747);
and U392 (N_392,In_347,In_477);
nand U393 (N_393,In_585,In_210);
or U394 (N_394,In_512,In_699);
xnor U395 (N_395,In_2154,In_1520);
and U396 (N_396,In_1474,In_646);
and U397 (N_397,In_1053,In_1669);
xor U398 (N_398,In_2183,In_344);
nand U399 (N_399,In_1200,In_79);
and U400 (N_400,In_2294,In_1268);
and U401 (N_401,In_51,In_1693);
xor U402 (N_402,In_808,In_897);
or U403 (N_403,In_1487,In_919);
xor U404 (N_404,In_1620,In_1385);
nor U405 (N_405,In_1989,In_1777);
nand U406 (N_406,In_1100,In_881);
xnor U407 (N_407,In_2312,In_2171);
or U408 (N_408,In_1439,In_253);
or U409 (N_409,In_623,In_1803);
or U410 (N_410,In_880,In_305);
nor U411 (N_411,In_406,In_1730);
or U412 (N_412,In_678,In_1763);
xor U413 (N_413,In_2434,In_1193);
xnor U414 (N_414,In_1300,In_1645);
xnor U415 (N_415,In_122,In_1149);
or U416 (N_416,In_167,In_1734);
or U417 (N_417,In_680,In_230);
or U418 (N_418,In_1319,In_2476);
and U419 (N_419,In_673,In_2099);
and U420 (N_420,In_2379,In_865);
xnor U421 (N_421,In_1564,In_290);
xnor U422 (N_422,In_84,In_2160);
or U423 (N_423,In_2223,In_490);
nand U424 (N_424,In_1872,In_1206);
nor U425 (N_425,In_1503,In_81);
nor U426 (N_426,In_1868,In_628);
xnor U427 (N_427,In_2400,In_653);
and U428 (N_428,In_291,In_1088);
and U429 (N_429,In_1356,In_1901);
and U430 (N_430,In_1247,In_2288);
or U431 (N_431,In_489,In_583);
and U432 (N_432,In_682,In_1695);
xnor U433 (N_433,In_1987,In_2198);
nand U434 (N_434,In_2177,In_339);
xnor U435 (N_435,In_2001,In_1537);
or U436 (N_436,In_52,In_1671);
and U437 (N_437,In_2292,In_1878);
or U438 (N_438,In_380,In_2334);
nand U439 (N_439,In_1020,In_460);
xnor U440 (N_440,In_1329,In_30);
nand U441 (N_441,In_240,In_394);
and U442 (N_442,In_247,In_1435);
nor U443 (N_443,In_1334,In_2011);
xor U444 (N_444,In_1033,In_1024);
nand U445 (N_445,In_1575,In_335);
and U446 (N_446,In_527,In_1034);
and U447 (N_447,In_455,In_1970);
or U448 (N_448,In_97,In_1517);
nand U449 (N_449,In_544,In_111);
or U450 (N_450,In_2128,In_810);
nor U451 (N_451,In_104,In_804);
and U452 (N_452,In_2484,In_1059);
and U453 (N_453,In_1585,In_1164);
nor U454 (N_454,In_743,In_108);
or U455 (N_455,In_2044,In_110);
nor U456 (N_456,In_1190,In_1299);
or U457 (N_457,In_114,In_640);
and U458 (N_458,In_728,In_333);
nand U459 (N_459,In_1000,In_1126);
nor U460 (N_460,In_1706,In_1996);
and U461 (N_461,In_419,In_31);
and U462 (N_462,In_321,In_46);
nand U463 (N_463,In_847,In_2255);
nor U464 (N_464,In_361,In_773);
nand U465 (N_465,In_164,In_475);
or U466 (N_466,In_416,In_2276);
nor U467 (N_467,In_608,In_262);
nor U468 (N_468,In_963,In_1147);
nand U469 (N_469,In_289,In_409);
nand U470 (N_470,In_386,In_131);
or U471 (N_471,In_2228,In_2403);
nand U472 (N_472,In_651,In_1639);
or U473 (N_473,In_664,In_1180);
and U474 (N_474,In_1980,In_1974);
xnor U475 (N_475,In_666,In_140);
nor U476 (N_476,In_1541,In_1513);
and U477 (N_477,In_1929,In_15);
xor U478 (N_478,In_979,In_2443);
or U479 (N_479,In_1395,In_2371);
or U480 (N_480,In_2143,In_611);
and U481 (N_481,In_1726,In_1573);
nand U482 (N_482,In_418,In_352);
xnor U483 (N_483,In_659,In_2014);
nor U484 (N_484,In_1649,In_2220);
nand U485 (N_485,In_1656,In_270);
and U486 (N_486,In_1236,In_2387);
nand U487 (N_487,In_2486,In_1621);
xor U488 (N_488,In_985,In_434);
or U489 (N_489,In_398,In_1529);
nor U490 (N_490,In_1631,In_195);
xnor U491 (N_491,In_1216,In_1318);
and U492 (N_492,In_2471,In_1778);
nand U493 (N_493,In_1374,In_2431);
nor U494 (N_494,In_840,In_168);
nand U495 (N_495,In_1965,In_831);
or U496 (N_496,In_146,In_1171);
nand U497 (N_497,In_2447,In_1563);
xnor U498 (N_498,In_393,In_1725);
xor U499 (N_499,In_2372,In_1531);
nand U500 (N_500,In_1634,In_1625);
or U501 (N_501,In_1595,In_2283);
or U502 (N_502,In_238,In_2325);
nor U503 (N_503,In_1993,In_615);
and U504 (N_504,In_2272,In_297);
xnor U505 (N_505,In_540,In_889);
and U506 (N_506,In_845,In_2133);
nor U507 (N_507,In_1044,In_1137);
or U508 (N_508,In_421,In_42);
and U509 (N_509,In_2487,In_1477);
nor U510 (N_510,In_1744,In_980);
or U511 (N_511,In_2404,In_488);
nand U512 (N_512,In_2226,In_1330);
or U513 (N_513,In_676,In_2296);
or U514 (N_514,In_2054,In_671);
or U515 (N_515,In_200,In_1920);
and U516 (N_516,In_590,In_1522);
or U517 (N_517,In_1546,In_1081);
nor U518 (N_518,In_2344,In_1556);
xor U519 (N_519,In_1342,In_1663);
and U520 (N_520,In_741,In_91);
xnor U521 (N_521,In_1022,In_918);
xnor U522 (N_522,In_2200,In_1651);
nand U523 (N_523,In_821,In_2132);
nor U524 (N_524,In_1727,In_552);
and U525 (N_525,In_535,In_1209);
nand U526 (N_526,In_5,In_2440);
or U527 (N_527,In_1398,In_1416);
nor U528 (N_528,In_3,In_2284);
and U529 (N_529,In_1999,In_2489);
and U530 (N_530,In_2251,In_1512);
nor U531 (N_531,In_2164,In_1832);
xnor U532 (N_532,In_926,In_2204);
nand U533 (N_533,In_736,In_328);
and U534 (N_534,In_26,In_445);
nor U535 (N_535,In_1525,In_1415);
or U536 (N_536,In_298,In_2295);
or U537 (N_537,In_675,In_2040);
and U538 (N_538,In_871,In_1811);
or U539 (N_539,In_1157,In_1717);
and U540 (N_540,In_1370,In_1028);
xor U541 (N_541,In_408,In_1705);
nor U542 (N_542,In_227,In_1073);
nor U543 (N_543,In_2115,In_2360);
or U544 (N_544,In_250,In_2016);
or U545 (N_545,In_185,In_696);
xnor U546 (N_546,In_2273,In_733);
nor U547 (N_547,In_2441,In_851);
nand U548 (N_548,In_437,In_1475);
nor U549 (N_549,In_480,In_345);
xor U550 (N_550,In_2059,In_2274);
nand U551 (N_551,In_1821,In_1861);
nor U552 (N_552,In_2477,In_1670);
or U553 (N_553,In_462,In_992);
or U554 (N_554,In_366,In_1070);
xor U555 (N_555,In_1750,In_1536);
nand U556 (N_556,In_299,In_1903);
or U557 (N_557,In_898,In_72);
xor U558 (N_558,In_1812,In_2281);
and U559 (N_559,In_814,In_1258);
nand U560 (N_560,In_911,In_894);
and U561 (N_561,In_1050,In_1842);
and U562 (N_562,In_1285,In_2330);
nor U563 (N_563,In_2264,In_414);
or U564 (N_564,In_1284,In_135);
xor U565 (N_565,In_2139,In_767);
and U566 (N_566,In_2074,In_2010);
and U567 (N_567,In_1781,In_2008);
and U568 (N_568,In_502,In_2326);
nand U569 (N_569,In_2339,In_1566);
nor U570 (N_570,In_1220,In_916);
or U571 (N_571,In_1276,In_2349);
and U572 (N_572,In_1755,In_184);
nand U573 (N_573,In_761,In_1241);
nand U574 (N_574,In_1459,In_1083);
nor U575 (N_575,In_1127,In_2024);
xor U576 (N_576,In_2382,In_2009);
nand U577 (N_577,In_1198,In_60);
xnor U578 (N_578,In_1850,In_2202);
nor U579 (N_579,In_619,In_1908);
nand U580 (N_580,In_1560,In_257);
nor U581 (N_581,In_679,In_983);
nor U582 (N_582,In_2100,In_1937);
xor U583 (N_583,In_2086,In_782);
nor U584 (N_584,In_1315,In_451);
or U585 (N_585,In_2494,In_157);
and U586 (N_586,In_1466,In_2493);
nor U587 (N_587,In_166,In_1472);
nor U588 (N_588,In_2474,In_1841);
or U589 (N_589,In_220,In_431);
nor U590 (N_590,In_182,In_966);
nand U591 (N_591,In_41,In_1321);
xor U592 (N_592,In_1479,In_2215);
or U593 (N_593,In_165,In_2430);
and U594 (N_594,In_1839,In_707);
nor U595 (N_595,In_85,In_2144);
nand U596 (N_596,In_1463,In_2092);
nand U597 (N_597,In_1900,In_604);
and U598 (N_598,In_1860,In_1275);
nor U599 (N_599,In_1085,In_2196);
and U600 (N_600,In_1636,In_780);
nand U601 (N_601,In_233,In_127);
and U602 (N_602,In_597,In_1949);
and U603 (N_603,In_360,In_1756);
xor U604 (N_604,In_1235,In_1854);
xnor U605 (N_605,In_2004,In_1751);
and U606 (N_606,In_1387,In_473);
xnor U607 (N_607,In_1401,In_1940);
xnor U608 (N_608,In_315,In_2266);
or U609 (N_609,In_493,In_2263);
xor U610 (N_610,In_2393,In_1554);
nand U611 (N_611,In_1309,In_2227);
nand U612 (N_612,In_1291,In_2108);
and U613 (N_613,In_1201,In_1499);
xnor U614 (N_614,In_592,In_827);
or U615 (N_615,In_355,In_690);
nand U616 (N_616,In_975,In_21);
nor U617 (N_617,In_971,In_2119);
or U618 (N_618,In_2315,In_2445);
or U619 (N_619,In_1951,In_1048);
and U620 (N_620,In_458,In_2293);
nor U621 (N_621,In_1386,In_1436);
and U622 (N_622,In_64,In_2022);
nor U623 (N_623,In_853,In_796);
xnor U624 (N_624,In_598,In_2408);
xor U625 (N_625,In_436,In_443);
xor U626 (N_626,In_1170,In_2391);
and U627 (N_627,In_322,In_1911);
nor U628 (N_628,In_2411,In_1402);
xor U629 (N_629,In_636,In_879);
nand U630 (N_630,In_2278,In_1155);
xor U631 (N_631,In_1885,In_2085);
nor U632 (N_632,In_2122,In_214);
xnor U633 (N_633,In_750,In_1927);
and U634 (N_634,In_1904,In_1953);
nand U635 (N_635,In_521,In_1971);
xnor U636 (N_636,In_1312,In_2063);
nand U637 (N_637,In_1473,In_466);
or U638 (N_638,In_620,In_1922);
nand U639 (N_639,In_1497,In_2007);
nor U640 (N_640,In_1015,In_1724);
nor U641 (N_641,In_246,In_1692);
xnor U642 (N_642,In_1110,In_23);
nor U643 (N_643,In_2491,In_1333);
or U644 (N_644,In_67,In_2167);
and U645 (N_645,In_1253,In_1432);
or U646 (N_646,In_1464,In_2245);
and U647 (N_647,In_234,In_1326);
and U648 (N_648,In_2313,In_350);
xor U649 (N_649,In_1410,In_1451);
nor U650 (N_650,In_2436,In_1184);
nor U651 (N_651,In_1218,In_71);
nor U652 (N_652,In_1449,In_965);
and U653 (N_653,In_1715,In_65);
or U654 (N_654,In_2193,In_2492);
nand U655 (N_655,In_32,In_850);
and U656 (N_656,In_357,In_192);
nand U657 (N_657,In_1761,In_2121);
and U658 (N_658,In_2254,In_456);
nand U659 (N_659,In_1549,In_1010);
xnor U660 (N_660,In_1591,In_278);
and U661 (N_661,In_866,In_732);
xor U662 (N_662,In_1454,In_1921);
nor U663 (N_663,In_627,In_1017);
or U664 (N_664,In_359,In_1207);
xor U665 (N_665,In_872,In_259);
and U666 (N_666,In_656,In_1409);
and U667 (N_667,In_1714,In_1331);
nand U668 (N_668,In_1414,In_1592);
nor U669 (N_669,In_2458,In_1151);
nand U670 (N_670,In_2013,In_1859);
nand U671 (N_671,In_187,In_1943);
and U672 (N_672,In_1450,In_642);
xnor U673 (N_673,In_441,In_812);
or U674 (N_674,In_1278,In_2039);
nand U675 (N_675,In_0,In_978);
or U676 (N_676,In_1144,In_887);
or U677 (N_677,In_1659,In_1882);
and U678 (N_678,In_863,In_873);
or U679 (N_679,In_1578,In_442);
or U680 (N_680,In_1146,In_38);
nor U681 (N_681,In_1637,In_1089);
nor U682 (N_682,In_260,In_1853);
or U683 (N_683,In_2410,In_1884);
or U684 (N_684,In_1470,In_501);
nand U685 (N_685,In_631,In_1287);
nor U686 (N_686,In_2423,In_1035);
or U687 (N_687,In_2418,In_1323);
nor U688 (N_688,In_522,In_327);
nor U689 (N_689,In_1836,In_1314);
nand U690 (N_690,In_2473,In_1411);
nand U691 (N_691,In_2433,In_2229);
and U692 (N_692,In_271,In_1270);
nand U693 (N_693,In_1320,In_2314);
or U694 (N_694,In_212,In_2416);
nand U695 (N_695,In_1016,In_223);
or U696 (N_696,In_1265,In_2361);
or U697 (N_697,In_1879,In_693);
nor U698 (N_698,In_1257,In_579);
nor U699 (N_699,In_476,In_293);
nand U700 (N_700,In_2137,In_625);
nand U701 (N_701,In_1720,In_970);
nor U702 (N_702,In_555,In_1509);
and U703 (N_703,In_1390,In_56);
or U704 (N_704,In_2355,In_1886);
nand U705 (N_705,In_922,In_2147);
xor U706 (N_706,In_2322,In_541);
or U707 (N_707,In_1975,In_358);
nand U708 (N_708,In_1511,In_217);
xnor U709 (N_709,In_1611,In_868);
nand U710 (N_710,In_1712,In_2485);
or U711 (N_711,In_2397,In_974);
nor U712 (N_712,In_420,In_567);
and U713 (N_713,In_1092,In_396);
or U714 (N_714,In_685,In_1383);
nand U715 (N_715,In_706,In_449);
nand U716 (N_716,In_2002,In_1430);
or U717 (N_717,In_285,In_1869);
nor U718 (N_718,In_80,In_424);
nand U719 (N_719,In_243,In_596);
xnor U720 (N_720,In_115,In_1080);
nand U721 (N_721,In_684,In_2461);
nor U722 (N_722,In_1961,In_1174);
nor U723 (N_723,In_2499,In_1972);
xnor U724 (N_724,In_2421,In_2045);
nor U725 (N_725,In_948,In_1913);
and U726 (N_726,In_1570,In_2279);
or U727 (N_727,In_123,In_504);
and U728 (N_728,In_2145,In_1518);
nand U729 (N_729,In_813,In_944);
and U730 (N_730,In_1084,In_1507);
nor U731 (N_731,In_2201,In_1255);
nand U732 (N_732,In_2000,In_570);
xnor U733 (N_733,In_28,In_835);
xnor U734 (N_734,In_385,In_206);
or U735 (N_735,In_1932,In_2151);
xor U736 (N_736,In_1124,In_2187);
xor U737 (N_737,In_1881,In_1944);
nor U738 (N_738,In_2090,In_546);
and U739 (N_739,In_565,In_381);
nor U740 (N_740,In_2454,In_2149);
xor U741 (N_741,In_2207,In_2138);
nand U742 (N_742,In_697,In_1071);
xnor U743 (N_743,In_2320,In_1916);
nand U744 (N_744,In_2269,In_776);
nand U745 (N_745,In_55,In_1004);
xor U746 (N_746,In_2353,In_202);
xor U747 (N_747,In_427,In_1368);
nor U748 (N_748,In_117,In_383);
or U749 (N_749,In_295,In_593);
nor U750 (N_750,In_1569,In_511);
or U751 (N_751,In_411,In_129);
nand U752 (N_752,In_1618,In_296);
and U753 (N_753,In_1703,In_806);
nor U754 (N_754,In_1704,In_2260);
nand U755 (N_755,In_1023,In_2282);
nor U756 (N_756,In_1646,In_1766);
xnor U757 (N_757,In_1969,In_1391);
and U758 (N_758,In_149,In_346);
nand U759 (N_759,In_2462,In_2192);
and U760 (N_760,In_1682,In_73);
and U761 (N_761,In_1357,In_323);
and U762 (N_762,In_1771,In_2415);
nand U763 (N_763,In_2127,In_1624);
nor U764 (N_764,In_1232,In_1058);
and U765 (N_765,In_1604,In_1215);
xnor U766 (N_766,In_154,In_2456);
nand U767 (N_767,In_279,In_1739);
nor U768 (N_768,In_1515,In_2261);
xor U769 (N_769,In_487,In_686);
and U770 (N_770,In_554,In_89);
xor U771 (N_771,In_1580,In_1930);
nand U772 (N_772,In_1267,In_1271);
nor U773 (N_773,In_1552,In_1752);
and U774 (N_774,In_2478,In_609);
and U775 (N_775,In_235,In_1888);
or U776 (N_776,In_48,In_2072);
nor U777 (N_777,In_1586,In_77);
or U778 (N_778,In_2304,In_1785);
nand U779 (N_779,In_221,In_1690);
xor U780 (N_780,In_1077,In_232);
nand U781 (N_781,In_751,In_1534);
xor U782 (N_782,In_2190,In_1069);
nand U783 (N_783,In_859,In_2199);
and U784 (N_784,In_1123,In_1447);
nand U785 (N_785,In_1242,In_1818);
nand U786 (N_786,In_1217,In_1681);
or U787 (N_787,In_558,In_2191);
nand U788 (N_788,In_765,In_1363);
nor U789 (N_789,In_900,In_1043);
nand U790 (N_790,In_1834,In_1160);
nor U791 (N_791,In_485,In_2359);
nor U792 (N_792,In_1532,In_1074);
xor U793 (N_793,In_1866,In_1551);
nand U794 (N_794,In_76,In_708);
and U795 (N_795,In_1992,In_45);
and U796 (N_796,In_711,In_2270);
nand U797 (N_797,In_1889,In_2107);
nor U798 (N_798,In_613,In_2450);
nand U799 (N_799,In_324,In_158);
and U800 (N_800,In_2449,In_429);
nand U801 (N_801,In_1012,In_1113);
or U802 (N_802,In_1909,In_822);
nor U803 (N_803,In_513,In_69);
nand U804 (N_804,In_2475,In_367);
or U805 (N_805,In_1143,In_1131);
nand U806 (N_806,In_93,In_1865);
or U807 (N_807,In_771,In_2352);
nor U808 (N_808,In_1005,In_139);
xnor U809 (N_809,In_805,In_893);
and U810 (N_810,In_2305,In_61);
and U811 (N_811,In_302,In_2050);
and U812 (N_812,In_1641,In_348);
or U813 (N_813,In_739,In_1962);
or U814 (N_814,In_660,In_1702);
nand U815 (N_815,In_1533,In_839);
nand U816 (N_816,In_2066,In_2237);
nor U817 (N_817,In_1794,In_823);
nand U818 (N_818,In_1630,In_2068);
xnor U819 (N_819,In_1555,In_703);
or U820 (N_820,In_1858,In_78);
nand U821 (N_821,In_610,In_1129);
nand U822 (N_822,In_1428,In_2285);
nor U823 (N_823,In_820,In_1192);
and U824 (N_824,In_313,In_529);
or U825 (N_825,In_225,In_795);
xnor U826 (N_826,In_362,In_617);
xnor U827 (N_827,In_2088,In_794);
nand U828 (N_828,In_2203,In_198);
xnor U829 (N_829,In_126,In_1027);
or U830 (N_830,In_940,In_1288);
and U831 (N_831,In_1306,In_1742);
xnor U832 (N_832,In_1899,In_268);
or U833 (N_833,In_1713,In_1590);
xor U834 (N_834,In_498,In_2468);
xor U835 (N_835,In_118,In_537);
nand U836 (N_836,In_1918,In_713);
and U837 (N_837,In_44,In_159);
nand U838 (N_838,In_54,In_263);
or U839 (N_839,In_1905,In_2275);
nor U840 (N_840,In_179,In_2414);
xor U841 (N_841,In_1352,In_1307);
xnor U842 (N_842,In_2056,In_1728);
nor U843 (N_843,In_2298,In_991);
nand U844 (N_844,In_2243,In_517);
and U845 (N_845,In_2047,In_652);
and U846 (N_846,In_2166,In_1103);
or U847 (N_847,In_92,In_1354);
xor U848 (N_848,In_177,In_1392);
or U849 (N_849,In_1855,In_1787);
nand U850 (N_850,In_1735,In_287);
or U851 (N_851,In_1662,In_2409);
xnor U852 (N_852,In_635,In_2189);
nand U853 (N_853,In_730,In_2287);
and U854 (N_854,In_1197,In_961);
or U855 (N_855,In_2041,In_2094);
nand U856 (N_856,In_639,In_589);
or U857 (N_857,In_231,In_329);
nor U858 (N_858,In_1173,In_2347);
nand U859 (N_859,In_1364,In_888);
or U860 (N_860,In_2388,In_68);
xnor U861 (N_861,In_2018,In_2448);
and U862 (N_862,In_24,In_644);
or U863 (N_863,In_542,In_369);
nor U864 (N_864,In_1445,In_1991);
xnor U865 (N_865,In_621,In_326);
nand U866 (N_866,In_1182,In_1694);
xor U867 (N_867,In_1408,In_2231);
xnor U868 (N_868,In_2058,In_1063);
nand U869 (N_869,In_2374,In_2250);
or U870 (N_870,In_1317,In_1446);
and U871 (N_871,In_1008,In_1122);
nor U872 (N_872,In_495,In_1893);
nor U873 (N_873,In_325,In_112);
nand U874 (N_874,In_672,In_1325);
nand U875 (N_875,In_2186,In_2084);
nand U876 (N_876,In_1805,In_936);
nand U877 (N_877,In_365,In_109);
and U878 (N_878,In_525,In_506);
nor U879 (N_879,In_1480,In_1516);
xnor U880 (N_880,In_378,In_316);
nand U881 (N_881,In_624,In_1667);
and U882 (N_882,In_1990,In_1938);
and U883 (N_883,In_1647,In_86);
xor U884 (N_884,In_2497,In_569);
or U885 (N_885,In_1568,In_1919);
or U886 (N_886,In_928,In_1039);
and U887 (N_887,In_1003,In_1483);
nor U888 (N_888,In_1802,In_156);
and U889 (N_889,In_2214,In_397);
nor U890 (N_890,In_1388,In_2335);
nor U891 (N_891,In_1018,In_1327);
and U892 (N_892,In_1711,In_508);
nand U893 (N_893,In_134,In_1539);
xor U894 (N_894,In_1615,In_1163);
or U895 (N_895,In_102,In_1583);
xnor U896 (N_896,In_2369,In_1597);
nand U897 (N_897,In_1492,In_283);
or U898 (N_898,In_994,In_401);
nand U899 (N_899,In_830,In_1280);
or U900 (N_900,In_494,In_998);
nor U901 (N_901,In_518,In_1051);
nor U902 (N_902,In_633,In_1810);
and U903 (N_903,In_201,In_2114);
nand U904 (N_904,In_1988,In_36);
nand U905 (N_905,In_2029,In_1500);
and U906 (N_906,In_2053,In_12);
xor U907 (N_907,In_103,In_1589);
xnor U908 (N_908,In_560,In_1576);
and U909 (N_909,In_252,In_857);
nor U910 (N_910,In_858,In_2354);
xnor U911 (N_911,In_1910,In_2318);
and U912 (N_912,In_207,In_340);
nor U913 (N_913,In_933,In_2104);
nor U914 (N_914,In_1133,In_2098);
nand U915 (N_915,In_1678,In_738);
and U916 (N_916,In_1632,In_1856);
nor U917 (N_917,In_1407,In_663);
xnor U918 (N_918,In_987,In_1001);
nand U919 (N_919,In_947,In_2221);
nor U920 (N_920,In_447,In_2129);
xor U921 (N_921,In_373,In_2457);
xor U922 (N_922,In_1801,In_1765);
nand U923 (N_923,In_2087,In_1091);
nand U924 (N_924,In_1075,In_1862);
nor U925 (N_925,In_543,In_1286);
and U926 (N_926,In_520,In_2141);
nor U927 (N_927,In_972,In_310);
and U928 (N_928,In_1272,In_384);
xnor U929 (N_929,In_1478,In_1599);
and U930 (N_930,In_2463,In_1396);
nand U931 (N_931,In_1426,In_334);
and U932 (N_932,In_1572,In_1150);
and U933 (N_933,In_734,In_2432);
nand U934 (N_934,In_2102,In_550);
and U935 (N_935,In_953,In_952);
or U936 (N_936,In_895,In_1506);
nor U937 (N_937,In_681,In_2142);
or U938 (N_938,In_1400,In_740);
nor U939 (N_939,In_1376,In_25);
nor U940 (N_940,In_841,In_265);
or U941 (N_941,In_116,In_2105);
nand U942 (N_942,In_1680,In_1225);
nand U943 (N_943,In_1668,In_1037);
or U944 (N_944,In_294,In_1042);
xor U945 (N_945,In_942,In_1097);
and U946 (N_946,In_1941,In_1488);
xor U947 (N_947,In_2168,In_377);
or U948 (N_948,In_2020,In_662);
and U949 (N_949,In_1102,In_1457);
xnor U950 (N_950,In_967,In_2390);
or U951 (N_951,In_341,In_997);
and U952 (N_952,In_1304,In_1553);
nor U953 (N_953,In_1754,In_132);
and U954 (N_954,In_1296,In_1817);
xnor U955 (N_955,In_2481,In_2033);
nor U956 (N_956,In_1188,In_532);
or U957 (N_957,In_1195,In_1798);
and U958 (N_958,In_602,In_2316);
xor U959 (N_959,In_1471,In_1653);
or U960 (N_960,In_1978,In_1465);
xnor U961 (N_961,In_269,In_1234);
nor U962 (N_962,In_1915,In_1581);
or U963 (N_963,In_756,In_867);
or U964 (N_964,In_1343,In_2267);
nor U965 (N_965,In_791,In_949);
nor U966 (N_966,In_1826,In_320);
xnor U967 (N_967,In_519,In_1460);
xnor U968 (N_968,In_1952,In_1203);
nand U969 (N_969,In_1600,In_655);
and U970 (N_970,In_2052,In_375);
nor U971 (N_971,In_1963,In_1191);
xor U972 (N_972,In_176,In_1056);
nor U973 (N_973,In_178,In_1337);
or U974 (N_974,In_1835,In_1372);
or U975 (N_975,In_981,In_2069);
nand U976 (N_976,In_1132,In_500);
or U977 (N_977,In_505,In_712);
or U978 (N_978,In_2234,In_2205);
and U979 (N_979,In_884,In_562);
and U980 (N_980,In_2280,In_1843);
nor U981 (N_981,In_654,In_1547);
or U982 (N_982,In_1776,In_1964);
xnor U983 (N_983,In_2146,In_787);
nor U984 (N_984,In_2005,In_1614);
nand U985 (N_985,In_1864,In_1076);
nand U986 (N_986,In_1616,In_789);
and U987 (N_987,In_861,In_74);
xor U988 (N_988,In_2363,In_1896);
nand U989 (N_989,In_1880,In_1579);
xnor U990 (N_990,In_704,In_1601);
and U991 (N_991,In_836,In_886);
xnor U992 (N_992,In_989,In_2206);
xor U993 (N_993,In_937,In_764);
or U994 (N_994,In_2453,In_1025);
nor U995 (N_995,In_1179,In_674);
nand U996 (N_996,In_687,In_39);
and U997 (N_997,In_2162,In_1565);
nand U998 (N_998,In_2338,In_753);
or U999 (N_999,In_203,In_1498);
and U1000 (N_1000,In_1052,In_1172);
or U1001 (N_1001,In_727,In_1950);
nand U1002 (N_1002,In_2159,In_999);
xor U1003 (N_1003,In_1104,In_1571);
and U1004 (N_1004,In_1442,In_2336);
or U1005 (N_1005,In_2028,In_1237);
nand U1006 (N_1006,In_968,In_2172);
xor U1007 (N_1007,In_2239,In_914);
and U1008 (N_1008,In_2362,In_2211);
xor U1009 (N_1009,In_1700,In_391);
nand U1010 (N_1010,In_1774,In_258);
nor U1011 (N_1011,In_1134,In_1524);
xnor U1012 (N_1012,In_215,In_105);
or U1013 (N_1013,In_700,In_412);
and U1014 (N_1014,In_1262,In_1784);
and U1015 (N_1015,In_2233,In_1468);
and U1016 (N_1016,In_459,In_1424);
and U1017 (N_1017,In_1281,In_2150);
nor U1018 (N_1018,In_2111,In_1141);
xnor U1019 (N_1019,In_461,In_468);
or U1020 (N_1020,In_2046,In_1577);
and U1021 (N_1021,In_622,In_1907);
nor U1022 (N_1022,In_1982,In_1683);
and U1023 (N_1023,In_1393,In_1397);
nand U1024 (N_1024,In_16,In_2256);
xor U1025 (N_1025,In_2017,In_1448);
nor U1026 (N_1026,In_2035,In_2079);
xnor U1027 (N_1027,In_783,In_121);
xnor U1028 (N_1028,In_582,In_1119);
xnor U1029 (N_1029,In_514,In_161);
and U1030 (N_1030,In_1594,In_594);
and U1031 (N_1031,In_1366,In_1983);
nand U1032 (N_1032,In_248,In_763);
and U1033 (N_1033,In_770,In_2125);
and U1034 (N_1034,In_2208,In_2123);
nand U1035 (N_1035,In_150,In_1222);
or U1036 (N_1036,In_83,In_2156);
nor U1037 (N_1037,In_417,In_2367);
nand U1038 (N_1038,In_1613,In_577);
or U1039 (N_1039,In_1006,In_792);
or U1040 (N_1040,In_1481,In_1117);
nand U1041 (N_1041,In_303,In_1925);
and U1042 (N_1042,In_1421,In_1118);
nor U1043 (N_1043,In_2195,In_855);
and U1044 (N_1044,In_1967,In_2161);
or U1045 (N_1045,In_1923,In_2265);
xor U1046 (N_1046,In_138,In_2377);
nor U1047 (N_1047,In_2173,In_2356);
xor U1048 (N_1048,In_524,In_2049);
xor U1049 (N_1049,In_1783,In_668);
nor U1050 (N_1050,In_2422,In_423);
or U1051 (N_1051,In_1002,In_1406);
xor U1052 (N_1052,In_1508,In_2340);
nor U1053 (N_1053,In_1313,In_2083);
xor U1054 (N_1054,In_1622,In_1429);
nor U1055 (N_1055,In_256,In_846);
and U1056 (N_1056,In_2103,In_2426);
nand U1057 (N_1057,In_2217,In_349);
xor U1058 (N_1058,In_374,In_614);
nor U1059 (N_1059,In_82,In_2118);
or U1060 (N_1060,In_2329,In_860);
and U1061 (N_1061,In_1707,In_1371);
or U1062 (N_1062,In_657,In_387);
nand U1063 (N_1063,In_722,In_351);
nand U1064 (N_1064,In_587,In_66);
and U1065 (N_1065,In_702,In_98);
nor U1066 (N_1066,In_2031,In_2078);
xnor U1067 (N_1067,In_1582,In_274);
xor U1068 (N_1068,In_1780,In_907);
and U1069 (N_1069,In_1968,In_1897);
and U1070 (N_1070,In_1404,In_1453);
xor U1071 (N_1071,In_864,In_1815);
xor U1072 (N_1072,In_977,In_59);
nor U1073 (N_1073,In_1948,In_729);
nor U1074 (N_1074,In_1139,In_647);
or U1075 (N_1075,In_749,In_626);
and U1076 (N_1076,In_1324,In_254);
and U1077 (N_1077,In_677,In_1748);
nor U1078 (N_1078,In_1419,In_2299);
and U1079 (N_1079,In_1238,In_486);
nand U1080 (N_1080,In_1227,In_1183);
and U1081 (N_1081,In_1403,In_927);
or U1082 (N_1082,In_1829,In_825);
xor U1083 (N_1083,In_308,In_1082);
or U1084 (N_1084,In_1947,In_891);
and U1085 (N_1085,In_2249,In_1528);
nand U1086 (N_1086,In_1867,In_120);
nor U1087 (N_1087,In_2130,In_1358);
or U1088 (N_1088,In_1365,In_509);
nor U1089 (N_1089,In_1890,In_1816);
and U1090 (N_1090,In_1120,In_2472);
or U1091 (N_1091,In_2,In_354);
and U1092 (N_1092,In_1699,In_2075);
and U1093 (N_1093,In_1046,In_1514);
nand U1094 (N_1094,In_1775,In_1347);
or U1095 (N_1095,In_1096,In_1883);
xnor U1096 (N_1096,In_1014,In_941);
nand U1097 (N_1097,In_1282,In_986);
nor U1098 (N_1098,In_1852,In_2030);
nor U1099 (N_1099,In_694,In_1264);
nor U1100 (N_1100,In_2025,In_2165);
xnor U1101 (N_1101,In_785,In_549);
nand U1102 (N_1102,In_1661,In_2213);
nor U1103 (N_1103,In_2082,In_1740);
xor U1104 (N_1104,In_683,In_1674);
nand U1105 (N_1105,In_1072,In_1538);
nand U1106 (N_1106,In_2366,In_1729);
xnor U1107 (N_1107,In_2375,In_824);
xnor U1108 (N_1108,In_630,In_1902);
xor U1109 (N_1109,In_1289,In_1094);
nand U1110 (N_1110,In_311,In_368);
and U1111 (N_1111,In_2055,In_244);
and U1112 (N_1112,In_1895,In_276);
nor U1113 (N_1113,In_723,In_43);
xnor U1114 (N_1114,In_2003,In_1917);
nor U1115 (N_1115,In_1823,In_1736);
nand U1116 (N_1116,In_342,In_1845);
or U1117 (N_1117,In_372,In_1425);
or U1118 (N_1118,In_563,In_1791);
nor U1119 (N_1119,In_784,In_2185);
nand U1120 (N_1120,In_793,In_802);
nand U1121 (N_1121,In_1530,In_938);
xor U1122 (N_1122,In_251,In_1521);
nor U1123 (N_1123,In_816,In_331);
and U1124 (N_1124,In_1544,In_2439);
nor U1125 (N_1125,In_746,In_491);
and U1126 (N_1126,In_175,In_432);
nand U1127 (N_1127,In_852,In_2328);
nand U1128 (N_1128,In_781,In_1648);
and U1129 (N_1129,In_1710,In_272);
or U1130 (N_1130,In_2309,In_1822);
nand U1131 (N_1131,In_2236,In_1976);
nand U1132 (N_1132,In_725,In_603);
xor U1133 (N_1133,In_1874,In_2412);
nor U1134 (N_1134,In_2048,In_1230);
nand U1135 (N_1135,In_1924,In_472);
nor U1136 (N_1136,In_1367,In_1954);
or U1137 (N_1137,In_745,In_35);
nand U1138 (N_1138,In_811,In_925);
or U1139 (N_1139,In_280,In_194);
or U1140 (N_1140,In_715,In_1526);
and U1141 (N_1141,In_1224,In_4);
and U1142 (N_1142,In_2386,In_1054);
nor U1143 (N_1143,In_667,In_1495);
xnor U1144 (N_1144,In_22,In_1152);
or U1145 (N_1145,In_854,In_1494);
or U1146 (N_1146,In_1799,In_976);
nand U1147 (N_1147,In_1808,In_1723);
and U1148 (N_1148,In_94,In_1244);
xor U1149 (N_1149,In_2258,In_2311);
or U1150 (N_1150,In_1914,In_1673);
xor U1151 (N_1151,In_2381,In_1557);
nand U1152 (N_1152,In_775,In_1685);
and U1153 (N_1153,In_1527,In_2032);
nand U1154 (N_1154,In_695,In_170);
nor U1155 (N_1155,In_1078,In_1958);
nand U1156 (N_1156,In_2290,In_564);
xor U1157 (N_1157,In_2209,In_330);
nand U1158 (N_1158,In_2073,In_1652);
nand U1159 (N_1159,In_1212,In_2182);
nor U1160 (N_1160,In_578,In_1679);
or U1161 (N_1161,In_2089,In_1140);
nand U1162 (N_1162,In_1456,In_1820);
xnor U1163 (N_1163,In_1977,In_828);
xnor U1164 (N_1164,In_1114,In_2302);
and U1165 (N_1165,In_2070,In_1031);
xor U1166 (N_1166,In_1476,In_395);
or U1167 (N_1167,In_281,In_2452);
nor U1168 (N_1168,In_1169,In_70);
or U1169 (N_1169,In_364,In_1485);
nor U1170 (N_1170,In_1154,In_2076);
nor U1171 (N_1171,In_2179,In_186);
or U1172 (N_1172,In_1676,In_807);
or U1173 (N_1173,In_1857,In_1762);
or U1174 (N_1174,In_2026,In_2394);
or U1175 (N_1175,In_1831,In_538);
nor U1176 (N_1176,In_57,In_2417);
nand U1177 (N_1177,In_1863,In_832);
or U1178 (N_1178,In_49,In_939);
or U1179 (N_1179,In_1760,In_2240);
nand U1180 (N_1180,In_574,In_748);
xor U1181 (N_1181,In_1316,In_474);
xnor U1182 (N_1182,In_1642,In_826);
and U1183 (N_1183,In_236,In_2435);
xnor U1184 (N_1184,In_2095,In_124);
xnor U1185 (N_1185,In_2368,In_1);
xor U1186 (N_1186,In_2232,In_870);
and U1187 (N_1187,In_309,In_1708);
and U1188 (N_1188,In_2451,In_548);
and U1189 (N_1189,In_648,In_1956);
and U1190 (N_1190,In_2348,In_2357);
xor U1191 (N_1191,In_1731,In_634);
or U1192 (N_1192,In_959,In_2483);
or U1193 (N_1193,In_382,In_2178);
nand U1194 (N_1194,In_1545,In_507);
or U1195 (N_1195,In_1166,In_484);
and U1196 (N_1196,In_1689,In_492);
and U1197 (N_1197,In_878,In_1086);
xor U1198 (N_1198,In_1809,In_2307);
or U1199 (N_1199,In_954,In_1032);
and U1200 (N_1200,In_561,In_2006);
nand U1201 (N_1201,In_1239,In_757);
xor U1202 (N_1202,In_1696,In_1800);
and U1203 (N_1203,In_1061,In_726);
nor U1204 (N_1204,In_249,In_242);
nor U1205 (N_1205,In_774,In_995);
or U1206 (N_1206,In_454,In_1931);
nand U1207 (N_1207,In_768,In_1159);
or U1208 (N_1208,In_536,In_1813);
xor U1209 (N_1209,In_1136,In_2163);
xnor U1210 (N_1210,In_1254,In_2038);
or U1211 (N_1211,In_422,In_917);
nor U1212 (N_1212,In_1196,In_1686);
nor U1213 (N_1213,In_1360,In_1047);
xor U1214 (N_1214,In_1231,In_2188);
nand U1215 (N_1215,In_844,In_2373);
nor U1216 (N_1216,In_869,In_1623);
nor U1217 (N_1217,In_843,In_1643);
xnor U1218 (N_1218,In_338,In_1745);
nor U1219 (N_1219,In_1698,In_817);
nand U1220 (N_1220,In_1099,In_1121);
and U1221 (N_1221,In_599,In_1807);
and U1222 (N_1222,In_2303,In_2238);
and U1223 (N_1223,In_2253,In_1340);
or U1224 (N_1224,In_267,In_1789);
or U1225 (N_1225,In_1346,In_876);
and U1226 (N_1226,In_1677,In_2337);
and U1227 (N_1227,In_2158,In_874);
nand U1228 (N_1228,In_1559,In_1960);
nand U1229 (N_1229,In_1870,In_1501);
and U1230 (N_1230,In_241,In_1359);
and U1231 (N_1231,In_779,In_1721);
xnor U1232 (N_1232,In_1389,In_584);
or U1233 (N_1233,In_902,In_1743);
nor U1234 (N_1234,In_90,In_710);
xnor U1235 (N_1235,In_1936,In_755);
and U1236 (N_1236,In_2077,In_1753);
or U1237 (N_1237,In_1243,In_428);
xor U1238 (N_1238,In_481,In_1759);
nor U1239 (N_1239,In_943,In_1303);
nor U1240 (N_1240,In_1098,In_18);
xnor U1241 (N_1241,In_2496,In_2271);
nand U1242 (N_1242,In_1995,In_735);
and U1243 (N_1243,In_183,In_2425);
xor U1244 (N_1244,In_645,In_2023);
nor U1245 (N_1245,In_404,In_58);
and U1246 (N_1246,In_95,In_724);
and U1247 (N_1247,In_2482,In_218);
and U1248 (N_1248,In_1221,In_1361);
nor U1249 (N_1249,In_882,In_113);
or U1250 (N_1250,N_628,N_770);
nor U1251 (N_1251,N_736,N_553);
nand U1252 (N_1252,N_964,N_230);
or U1253 (N_1253,N_669,N_386);
and U1254 (N_1254,N_1186,N_985);
nor U1255 (N_1255,N_449,N_176);
and U1256 (N_1256,N_5,N_746);
nand U1257 (N_1257,N_760,N_854);
nor U1258 (N_1258,N_896,N_956);
or U1259 (N_1259,N_247,N_693);
nor U1260 (N_1260,N_440,N_659);
xnor U1261 (N_1261,N_175,N_1139);
xor U1262 (N_1262,N_77,N_552);
nand U1263 (N_1263,N_150,N_315);
and U1264 (N_1264,N_439,N_713);
and U1265 (N_1265,N_1027,N_255);
nor U1266 (N_1266,N_246,N_194);
nand U1267 (N_1267,N_1215,N_573);
xor U1268 (N_1268,N_568,N_660);
and U1269 (N_1269,N_723,N_860);
nor U1270 (N_1270,N_144,N_1100);
or U1271 (N_1271,N_771,N_847);
nand U1272 (N_1272,N_498,N_1158);
or U1273 (N_1273,N_634,N_33);
nand U1274 (N_1274,N_735,N_438);
or U1275 (N_1275,N_1221,N_221);
nand U1276 (N_1276,N_614,N_138);
or U1277 (N_1277,N_49,N_548);
and U1278 (N_1278,N_502,N_578);
nand U1279 (N_1279,N_782,N_859);
xor U1280 (N_1280,N_139,N_218);
nand U1281 (N_1281,N_288,N_848);
or U1282 (N_1282,N_402,N_1137);
nor U1283 (N_1283,N_711,N_467);
nor U1284 (N_1284,N_201,N_397);
and U1285 (N_1285,N_401,N_67);
nand U1286 (N_1286,N_480,N_346);
or U1287 (N_1287,N_1169,N_967);
xor U1288 (N_1288,N_649,N_793);
nor U1289 (N_1289,N_1068,N_163);
nor U1290 (N_1290,N_581,N_24);
xnor U1291 (N_1291,N_489,N_753);
nor U1292 (N_1292,N_1083,N_441);
or U1293 (N_1293,N_1131,N_281);
and U1294 (N_1294,N_507,N_668);
and U1295 (N_1295,N_1220,N_792);
nand U1296 (N_1296,N_1004,N_17);
and U1297 (N_1297,N_991,N_470);
or U1298 (N_1298,N_1026,N_481);
nand U1299 (N_1299,N_118,N_688);
or U1300 (N_1300,N_635,N_172);
xnor U1301 (N_1301,N_1223,N_50);
or U1302 (N_1302,N_8,N_811);
nor U1303 (N_1303,N_1007,N_360);
nand U1304 (N_1304,N_1151,N_143);
nand U1305 (N_1305,N_119,N_667);
and U1306 (N_1306,N_1086,N_174);
or U1307 (N_1307,N_199,N_432);
nand U1308 (N_1308,N_14,N_237);
and U1309 (N_1309,N_1226,N_975);
xor U1310 (N_1310,N_679,N_1211);
nand U1311 (N_1311,N_1230,N_947);
nor U1312 (N_1312,N_475,N_1070);
and U1313 (N_1313,N_133,N_1097);
and U1314 (N_1314,N_1037,N_823);
xnor U1315 (N_1315,N_727,N_126);
or U1316 (N_1316,N_328,N_365);
or U1317 (N_1317,N_541,N_153);
and U1318 (N_1318,N_377,N_1062);
xnor U1319 (N_1319,N_640,N_580);
or U1320 (N_1320,N_617,N_238);
nor U1321 (N_1321,N_708,N_1154);
and U1322 (N_1322,N_652,N_897);
nor U1323 (N_1323,N_290,N_40);
xnor U1324 (N_1324,N_883,N_531);
nor U1325 (N_1325,N_534,N_493);
and U1326 (N_1326,N_239,N_84);
nor U1327 (N_1327,N_1020,N_382);
and U1328 (N_1328,N_719,N_2);
nor U1329 (N_1329,N_524,N_1059);
xnor U1330 (N_1330,N_390,N_666);
and U1331 (N_1331,N_876,N_979);
nor U1332 (N_1332,N_11,N_41);
or U1333 (N_1333,N_1051,N_453);
nand U1334 (N_1334,N_1144,N_343);
and U1335 (N_1335,N_393,N_943);
nor U1336 (N_1336,N_79,N_1034);
and U1337 (N_1337,N_1089,N_81);
nand U1338 (N_1338,N_62,N_105);
nand U1339 (N_1339,N_162,N_104);
xnor U1340 (N_1340,N_654,N_58);
and U1341 (N_1341,N_1016,N_880);
xor U1342 (N_1342,N_795,N_1061);
nor U1343 (N_1343,N_932,N_148);
or U1344 (N_1344,N_10,N_827);
xor U1345 (N_1345,N_384,N_38);
nor U1346 (N_1346,N_535,N_560);
nand U1347 (N_1347,N_1066,N_82);
or U1348 (N_1348,N_774,N_836);
nor U1349 (N_1349,N_170,N_1244);
nor U1350 (N_1350,N_137,N_706);
nand U1351 (N_1351,N_969,N_814);
nor U1352 (N_1352,N_1105,N_805);
nor U1353 (N_1353,N_1110,N_1035);
nand U1354 (N_1354,N_55,N_1145);
or U1355 (N_1355,N_444,N_100);
xnor U1356 (N_1356,N_630,N_1071);
nand U1357 (N_1357,N_341,N_1063);
or U1358 (N_1358,N_408,N_1127);
and U1359 (N_1359,N_1079,N_355);
or U1360 (N_1360,N_182,N_696);
or U1361 (N_1361,N_167,N_110);
nor U1362 (N_1362,N_1067,N_988);
or U1363 (N_1363,N_561,N_683);
nand U1364 (N_1364,N_491,N_973);
xor U1365 (N_1365,N_222,N_955);
nand U1366 (N_1366,N_734,N_154);
or U1367 (N_1367,N_677,N_737);
and U1368 (N_1368,N_92,N_1200);
or U1369 (N_1369,N_922,N_921);
or U1370 (N_1370,N_788,N_538);
nand U1371 (N_1371,N_752,N_487);
or U1372 (N_1372,N_161,N_692);
xor U1373 (N_1373,N_837,N_1210);
nand U1374 (N_1374,N_852,N_1231);
and U1375 (N_1375,N_1011,N_958);
nor U1376 (N_1376,N_845,N_252);
nor U1377 (N_1377,N_690,N_1164);
xnor U1378 (N_1378,N_46,N_822);
nand U1379 (N_1379,N_326,N_270);
or U1380 (N_1380,N_336,N_849);
nand U1381 (N_1381,N_933,N_1040);
or U1382 (N_1382,N_603,N_812);
xor U1383 (N_1383,N_1224,N_1195);
nor U1384 (N_1384,N_961,N_572);
nand U1385 (N_1385,N_1232,N_678);
and U1386 (N_1386,N_323,N_1045);
nor U1387 (N_1387,N_413,N_717);
nand U1388 (N_1388,N_530,N_1172);
nand U1389 (N_1389,N_529,N_1138);
xor U1390 (N_1390,N_145,N_865);
nand U1391 (N_1391,N_1123,N_591);
and U1392 (N_1392,N_395,N_807);
nand U1393 (N_1393,N_940,N_231);
nand U1394 (N_1394,N_160,N_851);
xor U1395 (N_1395,N_43,N_637);
nand U1396 (N_1396,N_482,N_1052);
nand U1397 (N_1397,N_1214,N_1111);
or U1398 (N_1398,N_405,N_949);
xnor U1399 (N_1399,N_796,N_398);
nor U1400 (N_1400,N_1208,N_935);
nor U1401 (N_1401,N_368,N_499);
nand U1402 (N_1402,N_1057,N_178);
or U1403 (N_1403,N_54,N_579);
or U1404 (N_1404,N_1162,N_773);
and U1405 (N_1405,N_98,N_798);
nor U1406 (N_1406,N_334,N_602);
or U1407 (N_1407,N_998,N_1133);
nand U1408 (N_1408,N_982,N_305);
nor U1409 (N_1409,N_1125,N_186);
and U1410 (N_1410,N_569,N_682);
or U1411 (N_1411,N_1174,N_89);
nand U1412 (N_1412,N_989,N_636);
and U1413 (N_1413,N_210,N_70);
xor U1414 (N_1414,N_117,N_1121);
and U1415 (N_1415,N_1190,N_1217);
xnor U1416 (N_1416,N_1192,N_516);
nand U1417 (N_1417,N_404,N_582);
nor U1418 (N_1418,N_604,N_939);
and U1419 (N_1419,N_846,N_1194);
xnor U1420 (N_1420,N_416,N_1113);
xnor U1421 (N_1421,N_1130,N_892);
xnor U1422 (N_1422,N_806,N_37);
nand U1423 (N_1423,N_942,N_644);
xor U1424 (N_1424,N_515,N_372);
xnor U1425 (N_1425,N_517,N_1202);
xor U1426 (N_1426,N_1042,N_26);
xnor U1427 (N_1427,N_362,N_1168);
or U1428 (N_1428,N_303,N_598);
nor U1429 (N_1429,N_1228,N_1116);
nor U1430 (N_1430,N_878,N_297);
nor U1431 (N_1431,N_592,N_913);
xor U1432 (N_1432,N_820,N_166);
nor U1433 (N_1433,N_1118,N_31);
nor U1434 (N_1434,N_891,N_45);
nand U1435 (N_1435,N_731,N_208);
nor U1436 (N_1436,N_226,N_586);
nor U1437 (N_1437,N_533,N_309);
nand U1438 (N_1438,N_631,N_695);
nand U1439 (N_1439,N_1247,N_1096);
or U1440 (N_1440,N_945,N_120);
nor U1441 (N_1441,N_433,N_1191);
nor U1442 (N_1442,N_465,N_25);
nand U1443 (N_1443,N_127,N_1104);
xor U1444 (N_1444,N_779,N_285);
nor U1445 (N_1445,N_224,N_742);
nand U1446 (N_1446,N_351,N_1126);
and U1447 (N_1447,N_220,N_358);
nand U1448 (N_1448,N_34,N_1182);
and U1449 (N_1449,N_278,N_471);
xnor U1450 (N_1450,N_1015,N_911);
xnor U1451 (N_1451,N_310,N_313);
xnor U1452 (N_1452,N_1108,N_387);
nand U1453 (N_1453,N_4,N_1073);
nor U1454 (N_1454,N_1044,N_71);
and U1455 (N_1455,N_862,N_1193);
nand U1456 (N_1456,N_214,N_1031);
xor U1457 (N_1457,N_497,N_1077);
and U1458 (N_1458,N_298,N_778);
nand U1459 (N_1459,N_35,N_920);
xnor U1460 (N_1460,N_1082,N_329);
xnor U1461 (N_1461,N_403,N_959);
nor U1462 (N_1462,N_1094,N_352);
nor U1463 (N_1463,N_767,N_96);
or U1464 (N_1464,N_687,N_686);
xnor U1465 (N_1465,N_27,N_195);
and U1466 (N_1466,N_374,N_267);
xor U1467 (N_1467,N_960,N_312);
nand U1468 (N_1468,N_757,N_898);
or U1469 (N_1469,N_664,N_809);
nand U1470 (N_1470,N_321,N_919);
nand U1471 (N_1471,N_207,N_1021);
xnor U1472 (N_1472,N_508,N_1084);
xnor U1473 (N_1473,N_112,N_775);
and U1474 (N_1474,N_269,N_1114);
xnor U1475 (N_1475,N_714,N_1024);
nand U1476 (N_1476,N_295,N_259);
nor U1477 (N_1477,N_463,N_681);
and U1478 (N_1478,N_129,N_625);
nand U1479 (N_1479,N_347,N_835);
xor U1480 (N_1480,N_394,N_544);
nand U1481 (N_1481,N_367,N_928);
nor U1482 (N_1482,N_789,N_462);
xor U1483 (N_1483,N_86,N_615);
nor U1484 (N_1484,N_981,N_1141);
nor U1485 (N_1485,N_1204,N_699);
xnor U1486 (N_1486,N_509,N_1205);
nor U1487 (N_1487,N_318,N_506);
xnor U1488 (N_1488,N_272,N_164);
nor U1489 (N_1489,N_16,N_997);
or U1490 (N_1490,N_483,N_545);
and U1491 (N_1491,N_769,N_103);
nand U1492 (N_1492,N_234,N_751);
nand U1493 (N_1493,N_294,N_818);
xnor U1494 (N_1494,N_1209,N_364);
nor U1495 (N_1495,N_136,N_142);
xor U1496 (N_1496,N_32,N_638);
nor U1497 (N_1497,N_510,N_146);
and U1498 (N_1498,N_749,N_722);
nand U1499 (N_1499,N_324,N_319);
nand U1500 (N_1500,N_1180,N_202);
and U1501 (N_1501,N_747,N_356);
nand U1502 (N_1502,N_1019,N_765);
nand U1503 (N_1503,N_206,N_426);
xor U1504 (N_1504,N_721,N_417);
and U1505 (N_1505,N_1201,N_768);
xnor U1506 (N_1506,N_1041,N_1239);
nor U1507 (N_1507,N_881,N_1003);
or U1508 (N_1508,N_607,N_791);
nand U1509 (N_1509,N_824,N_832);
and U1510 (N_1510,N_1,N_488);
xor U1511 (N_1511,N_950,N_915);
nand U1512 (N_1512,N_446,N_720);
nand U1513 (N_1513,N_523,N_1155);
nor U1514 (N_1514,N_442,N_155);
nor U1515 (N_1515,N_264,N_375);
nor U1516 (N_1516,N_597,N_263);
xor U1517 (N_1517,N_424,N_1122);
and U1518 (N_1518,N_858,N_813);
nand U1519 (N_1519,N_694,N_842);
or U1520 (N_1520,N_66,N_957);
nor U1521 (N_1521,N_1064,N_831);
xor U1522 (N_1522,N_741,N_1128);
or U1523 (N_1523,N_63,N_1008);
xor U1524 (N_1524,N_948,N_513);
xnor U1525 (N_1525,N_665,N_331);
and U1526 (N_1526,N_562,N_235);
or U1527 (N_1527,N_414,N_20);
and U1528 (N_1528,N_861,N_672);
and U1529 (N_1529,N_520,N_703);
or U1530 (N_1530,N_1075,N_583);
nor U1531 (N_1531,N_227,N_275);
nand U1532 (N_1532,N_1179,N_1119);
xnor U1533 (N_1533,N_1053,N_826);
and U1534 (N_1534,N_74,N_430);
and U1535 (N_1535,N_728,N_68);
nor U1536 (N_1536,N_726,N_134);
xnor U1537 (N_1537,N_1048,N_203);
nand U1538 (N_1538,N_626,N_787);
nand U1539 (N_1539,N_828,N_109);
or U1540 (N_1540,N_458,N_926);
nand U1541 (N_1541,N_344,N_1129);
xnor U1542 (N_1542,N_777,N_1022);
nand U1543 (N_1543,N_473,N_419);
or U1544 (N_1544,N_790,N_349);
nand U1545 (N_1545,N_622,N_1178);
xor U1546 (N_1546,N_140,N_1207);
xor U1547 (N_1547,N_657,N_1227);
nand U1548 (N_1548,N_299,N_1240);
nand U1549 (N_1549,N_115,N_627);
xnor U1550 (N_1550,N_645,N_786);
and U1551 (N_1551,N_443,N_191);
and U1552 (N_1552,N_585,N_1233);
nand U1553 (N_1553,N_1234,N_633);
xor U1554 (N_1554,N_917,N_400);
xor U1555 (N_1555,N_147,N_1103);
and U1556 (N_1556,N_527,N_707);
xnor U1557 (N_1557,N_528,N_188);
or U1558 (N_1558,N_781,N_213);
or U1559 (N_1559,N_1142,N_415);
nand U1560 (N_1560,N_361,N_550);
nor U1561 (N_1561,N_564,N_1199);
or U1562 (N_1562,N_342,N_141);
nand U1563 (N_1563,N_445,N_196);
nor U1564 (N_1564,N_651,N_850);
or U1565 (N_1565,N_1197,N_611);
xnor U1566 (N_1566,N_674,N_1124);
and U1567 (N_1567,N_761,N_165);
or U1568 (N_1568,N_965,N_1005);
xor U1569 (N_1569,N_745,N_1076);
nor U1570 (N_1570,N_558,N_407);
nand U1571 (N_1571,N_6,N_434);
nor U1572 (N_1572,N_1189,N_376);
and U1573 (N_1573,N_1173,N_1092);
xor U1574 (N_1574,N_451,N_983);
nand U1575 (N_1575,N_28,N_385);
nand U1576 (N_1576,N_9,N_325);
and U1577 (N_1577,N_610,N_431);
nand U1578 (N_1578,N_701,N_893);
or U1579 (N_1579,N_514,N_423);
and U1580 (N_1580,N_882,N_1198);
xor U1581 (N_1581,N_800,N_976);
xnor U1582 (N_1582,N_494,N_1159);
nand U1583 (N_1583,N_648,N_563);
and U1584 (N_1584,N_923,N_168);
and U1585 (N_1585,N_258,N_511);
or U1586 (N_1586,N_418,N_875);
xor U1587 (N_1587,N_301,N_931);
and U1588 (N_1588,N_1049,N_912);
and U1589 (N_1589,N_1212,N_1038);
and U1590 (N_1590,N_1036,N_539);
xor U1591 (N_1591,N_748,N_543);
or U1592 (N_1592,N_1032,N_241);
nor U1593 (N_1593,N_1000,N_816);
and U1594 (N_1594,N_383,N_829);
xnor U1595 (N_1595,N_565,N_3);
and U1596 (N_1596,N_877,N_780);
nor U1597 (N_1597,N_570,N_1033);
xnor U1598 (N_1598,N_113,N_276);
nor U1599 (N_1599,N_1243,N_1177);
or U1600 (N_1600,N_551,N_1136);
xor U1601 (N_1601,N_606,N_698);
or U1602 (N_1602,N_1181,N_863);
nor U1603 (N_1603,N_316,N_420);
or U1604 (N_1604,N_292,N_867);
or U1605 (N_1605,N_952,N_1196);
and U1606 (N_1606,N_559,N_1135);
xnor U1607 (N_1607,N_293,N_691);
and U1608 (N_1608,N_87,N_53);
xor U1609 (N_1609,N_459,N_966);
or U1610 (N_1610,N_843,N_799);
and U1611 (N_1611,N_750,N_608);
xor U1612 (N_1612,N_306,N_639);
or U1613 (N_1613,N_464,N_890);
or U1614 (N_1614,N_135,N_1107);
xor U1615 (N_1615,N_587,N_19);
nand U1616 (N_1616,N_277,N_609);
nor U1617 (N_1617,N_158,N_1153);
nor U1618 (N_1618,N_675,N_804);
or U1619 (N_1619,N_1120,N_518);
and U1620 (N_1620,N_980,N_461);
xnor U1621 (N_1621,N_48,N_599);
and U1622 (N_1622,N_1229,N_744);
and U1623 (N_1623,N_1009,N_759);
or U1624 (N_1624,N_57,N_962);
and U1625 (N_1625,N_557,N_83);
nand U1626 (N_1626,N_874,N_280);
nand U1627 (N_1627,N_522,N_712);
and U1628 (N_1628,N_339,N_332);
xnor U1629 (N_1629,N_994,N_974);
or U1630 (N_1630,N_457,N_85);
xor U1631 (N_1631,N_856,N_547);
or U1632 (N_1632,N_1170,N_479);
nor U1633 (N_1633,N_840,N_245);
nor U1634 (N_1634,N_205,N_1058);
xor U1635 (N_1635,N_918,N_121);
nand U1636 (N_1636,N_1056,N_1219);
nand U1637 (N_1637,N_266,N_260);
xnor U1638 (N_1638,N_906,N_571);
xor U1639 (N_1639,N_179,N_593);
nor U1640 (N_1640,N_619,N_743);
and U1641 (N_1641,N_577,N_653);
or U1642 (N_1642,N_111,N_501);
nor U1643 (N_1643,N_159,N_102);
and U1644 (N_1644,N_90,N_1157);
xnor U1645 (N_1645,N_624,N_1043);
or U1646 (N_1646,N_389,N_185);
nor U1647 (N_1647,N_594,N_1109);
xor U1648 (N_1648,N_819,N_307);
nor U1649 (N_1649,N_171,N_838);
and U1650 (N_1650,N_1095,N_283);
and U1651 (N_1651,N_1081,N_320);
xor U1652 (N_1652,N_184,N_888);
nor U1653 (N_1653,N_725,N_702);
xor U1654 (N_1654,N_51,N_732);
nand U1655 (N_1655,N_1017,N_546);
nor U1656 (N_1656,N_886,N_337);
and U1657 (N_1657,N_80,N_1088);
or U1658 (N_1658,N_485,N_1206);
nor U1659 (N_1659,N_618,N_392);
or U1660 (N_1660,N_810,N_934);
nand U1661 (N_1661,N_658,N_212);
xnor U1662 (N_1662,N_486,N_1091);
nor U1663 (N_1663,N_902,N_1241);
nand U1664 (N_1664,N_916,N_373);
xor U1665 (N_1665,N_1012,N_173);
xor U1666 (N_1666,N_1163,N_869);
nand U1667 (N_1667,N_1087,N_1047);
and U1668 (N_1668,N_478,N_549);
xor U1669 (N_1669,N_183,N_422);
or U1670 (N_1670,N_1167,N_60);
or U1671 (N_1671,N_951,N_525);
xnor U1672 (N_1672,N_925,N_1099);
nor U1673 (N_1673,N_370,N_335);
nor U1674 (N_1674,N_783,N_894);
or U1675 (N_1675,N_1188,N_899);
xnor U1676 (N_1676,N_595,N_21);
or U1677 (N_1677,N_938,N_1237);
xor U1678 (N_1678,N_1249,N_996);
nor U1679 (N_1679,N_42,N_354);
or U1680 (N_1680,N_632,N_215);
or U1681 (N_1681,N_620,N_588);
and U1682 (N_1682,N_521,N_1085);
xnor U1683 (N_1683,N_1117,N_399);
xnor U1684 (N_1684,N_287,N_492);
and U1685 (N_1685,N_904,N_302);
nor U1686 (N_1686,N_1161,N_772);
nor U1687 (N_1687,N_410,N_455);
or U1688 (N_1688,N_794,N_872);
and U1689 (N_1689,N_99,N_350);
xnor U1690 (N_1690,N_785,N_642);
and U1691 (N_1691,N_1246,N_1023);
or U1692 (N_1692,N_1150,N_1245);
or U1693 (N_1693,N_1065,N_1213);
nand U1694 (N_1694,N_512,N_271);
xor U1695 (N_1695,N_977,N_39);
nand U1696 (N_1696,N_406,N_460);
xor U1697 (N_1697,N_177,N_866);
nand U1698 (N_1698,N_596,N_327);
nand U1699 (N_1699,N_908,N_1149);
nand U1700 (N_1700,N_1175,N_661);
nand U1701 (N_1701,N_36,N_412);
xnor U1702 (N_1702,N_766,N_447);
nand U1703 (N_1703,N_1132,N_64);
xnor U1704 (N_1704,N_825,N_130);
or U1705 (N_1705,N_454,N_1112);
nor U1706 (N_1706,N_466,N_1074);
xor U1707 (N_1707,N_44,N_123);
or U1708 (N_1708,N_590,N_738);
xnor U1709 (N_1709,N_605,N_724);
and U1710 (N_1710,N_187,N_116);
xnor U1711 (N_1711,N_540,N_61);
xnor U1712 (N_1712,N_889,N_429);
and U1713 (N_1713,N_348,N_1055);
and U1714 (N_1714,N_248,N_914);
nor U1715 (N_1715,N_411,N_984);
or U1716 (N_1716,N_233,N_1236);
nor U1717 (N_1717,N_474,N_378);
xor U1718 (N_1718,N_643,N_1225);
and U1719 (N_1719,N_23,N_296);
and U1720 (N_1720,N_803,N_1046);
nor U1721 (N_1721,N_391,N_1183);
xor U1722 (N_1722,N_1025,N_114);
xnor U1723 (N_1723,N_671,N_1106);
and U1724 (N_1724,N_536,N_901);
and U1725 (N_1725,N_970,N_223);
xnor U1726 (N_1726,N_1060,N_225);
or U1727 (N_1727,N_1203,N_1160);
xnor U1728 (N_1728,N_261,N_219);
xor U1729 (N_1729,N_986,N_268);
xor U1730 (N_1730,N_733,N_314);
and U1731 (N_1731,N_601,N_556);
xor U1732 (N_1732,N_198,N_504);
nor U1733 (N_1733,N_476,N_169);
and U1734 (N_1734,N_282,N_197);
xor U1735 (N_1735,N_930,N_436);
nand U1736 (N_1736,N_340,N_1093);
or U1737 (N_1737,N_503,N_243);
xor U1738 (N_1738,N_937,N_262);
nor U1739 (N_1739,N_240,N_868);
xor U1740 (N_1740,N_953,N_662);
and U1741 (N_1741,N_125,N_363);
or U1742 (N_1742,N_670,N_448);
xor U1743 (N_1743,N_435,N_873);
or U1744 (N_1744,N_566,N_500);
or U1745 (N_1745,N_784,N_1222);
nand U1746 (N_1746,N_623,N_870);
xnor U1747 (N_1747,N_229,N_274);
and U1748 (N_1748,N_1002,N_1242);
nand U1749 (N_1749,N_380,N_963);
nand U1750 (N_1750,N_716,N_232);
or U1751 (N_1751,N_1146,N_1187);
and U1752 (N_1752,N_817,N_496);
xnor U1753 (N_1753,N_802,N_317);
nand U1754 (N_1754,N_1238,N_249);
and U1755 (N_1755,N_7,N_833);
or U1756 (N_1756,N_621,N_1152);
or U1757 (N_1757,N_519,N_600);
xor U1758 (N_1758,N_484,N_758);
nor U1759 (N_1759,N_1166,N_1148);
and U1760 (N_1760,N_575,N_576);
xnor U1761 (N_1761,N_844,N_685);
or U1762 (N_1762,N_30,N_655);
xor U1763 (N_1763,N_47,N_700);
or U1764 (N_1764,N_189,N_279);
nor U1765 (N_1765,N_75,N_1050);
and U1766 (N_1766,N_59,N_1134);
nand U1767 (N_1767,N_830,N_242);
xor U1768 (N_1768,N_106,N_353);
and U1769 (N_1769,N_542,N_124);
or U1770 (N_1770,N_801,N_855);
and U1771 (N_1771,N_18,N_1147);
and U1772 (N_1772,N_900,N_656);
and U1773 (N_1773,N_456,N_157);
nand U1774 (N_1774,N_756,N_990);
xnor U1775 (N_1775,N_616,N_15);
or U1776 (N_1776,N_650,N_663);
nand U1777 (N_1777,N_291,N_73);
xor U1778 (N_1778,N_477,N_180);
and U1779 (N_1779,N_1143,N_257);
xnor U1780 (N_1780,N_762,N_396);
xor U1781 (N_1781,N_1054,N_946);
and U1782 (N_1782,N_971,N_345);
nor U1783 (N_1783,N_537,N_428);
nor U1784 (N_1784,N_300,N_684);
xnor U1785 (N_1785,N_1078,N_371);
xor U1786 (N_1786,N_204,N_927);
nand U1787 (N_1787,N_76,N_265);
and U1788 (N_1788,N_612,N_1069);
xnor U1789 (N_1789,N_273,N_647);
xor U1790 (N_1790,N_244,N_1102);
xnor U1791 (N_1791,N_311,N_91);
nor U1792 (N_1792,N_156,N_495);
and U1793 (N_1793,N_108,N_1165);
and U1794 (N_1794,N_322,N_107);
xnor U1795 (N_1795,N_330,N_452);
nor U1796 (N_1796,N_56,N_641);
or U1797 (N_1797,N_821,N_629);
or U1798 (N_1798,N_1216,N_589);
or U1799 (N_1799,N_1171,N_0);
or U1800 (N_1800,N_211,N_381);
or U1801 (N_1801,N_730,N_236);
nor U1802 (N_1802,N_88,N_705);
and U1803 (N_1803,N_132,N_192);
nor U1804 (N_1804,N_879,N_193);
nand U1805 (N_1805,N_884,N_409);
nor U1806 (N_1806,N_1218,N_94);
and U1807 (N_1807,N_763,N_673);
xor U1808 (N_1808,N_1010,N_567);
nor U1809 (N_1809,N_999,N_887);
or U1810 (N_1810,N_490,N_697);
or U1811 (N_1811,N_1098,N_755);
nor U1812 (N_1812,N_993,N_200);
xor U1813 (N_1813,N_101,N_808);
and U1814 (N_1814,N_905,N_217);
and U1815 (N_1815,N_308,N_613);
nand U1816 (N_1816,N_776,N_379);
or U1817 (N_1817,N_1018,N_228);
and U1818 (N_1818,N_65,N_941);
xnor U1819 (N_1819,N_574,N_680);
nor U1820 (N_1820,N_357,N_388);
xor U1821 (N_1821,N_1101,N_944);
nor U1822 (N_1822,N_52,N_554);
and U1823 (N_1823,N_72,N_437);
nand U1824 (N_1824,N_715,N_505);
nor U1825 (N_1825,N_333,N_472);
and U1826 (N_1826,N_1014,N_834);
or U1827 (N_1827,N_1156,N_450);
nor U1828 (N_1828,N_936,N_1176);
xnor U1829 (N_1829,N_190,N_338);
or U1830 (N_1830,N_253,N_995);
xor U1831 (N_1831,N_1080,N_359);
or U1832 (N_1832,N_704,N_1090);
and U1833 (N_1833,N_929,N_181);
xnor U1834 (N_1834,N_1013,N_97);
xnor U1835 (N_1835,N_427,N_815);
xnor U1836 (N_1836,N_853,N_1001);
and U1837 (N_1837,N_1115,N_584);
and U1838 (N_1838,N_968,N_304);
and U1839 (N_1839,N_251,N_954);
nor U1840 (N_1840,N_1248,N_128);
xnor U1841 (N_1841,N_152,N_78);
nor U1842 (N_1842,N_739,N_366);
or U1843 (N_1843,N_909,N_885);
and U1844 (N_1844,N_841,N_1185);
nor U1845 (N_1845,N_1140,N_689);
nand U1846 (N_1846,N_903,N_709);
nand U1847 (N_1847,N_1028,N_69);
nand U1848 (N_1848,N_93,N_22);
nand U1849 (N_1849,N_924,N_425);
or U1850 (N_1850,N_421,N_839);
xor U1851 (N_1851,N_676,N_987);
or U1852 (N_1852,N_978,N_12);
nor U1853 (N_1853,N_532,N_149);
xnor U1854 (N_1854,N_122,N_871);
and U1855 (N_1855,N_369,N_151);
and U1856 (N_1856,N_764,N_710);
or U1857 (N_1857,N_646,N_555);
nand U1858 (N_1858,N_1235,N_1030);
nand U1859 (N_1859,N_526,N_284);
xnor U1860 (N_1860,N_797,N_972);
nor U1861 (N_1861,N_254,N_256);
xnor U1862 (N_1862,N_289,N_131);
nor U1863 (N_1863,N_29,N_216);
nand U1864 (N_1864,N_209,N_469);
xor U1865 (N_1865,N_907,N_718);
and U1866 (N_1866,N_250,N_857);
nor U1867 (N_1867,N_286,N_13);
nor U1868 (N_1868,N_895,N_1029);
nor U1869 (N_1869,N_864,N_95);
or U1870 (N_1870,N_468,N_992);
nor U1871 (N_1871,N_910,N_1072);
and U1872 (N_1872,N_1184,N_1006);
or U1873 (N_1873,N_1039,N_754);
and U1874 (N_1874,N_740,N_729);
or U1875 (N_1875,N_346,N_427);
nand U1876 (N_1876,N_1054,N_838);
and U1877 (N_1877,N_858,N_503);
nor U1878 (N_1878,N_1018,N_991);
and U1879 (N_1879,N_518,N_918);
xnor U1880 (N_1880,N_135,N_219);
or U1881 (N_1881,N_1185,N_290);
or U1882 (N_1882,N_25,N_1105);
xnor U1883 (N_1883,N_801,N_363);
xnor U1884 (N_1884,N_912,N_1225);
nand U1885 (N_1885,N_197,N_971);
nor U1886 (N_1886,N_1011,N_9);
xor U1887 (N_1887,N_632,N_604);
nor U1888 (N_1888,N_424,N_271);
and U1889 (N_1889,N_1098,N_362);
and U1890 (N_1890,N_114,N_67);
nand U1891 (N_1891,N_741,N_312);
and U1892 (N_1892,N_216,N_928);
nor U1893 (N_1893,N_449,N_477);
and U1894 (N_1894,N_366,N_1173);
xor U1895 (N_1895,N_334,N_417);
nand U1896 (N_1896,N_330,N_510);
nand U1897 (N_1897,N_839,N_273);
and U1898 (N_1898,N_168,N_719);
nand U1899 (N_1899,N_185,N_999);
and U1900 (N_1900,N_39,N_866);
nand U1901 (N_1901,N_283,N_267);
nor U1902 (N_1902,N_150,N_832);
or U1903 (N_1903,N_1166,N_971);
nor U1904 (N_1904,N_339,N_888);
xor U1905 (N_1905,N_281,N_191);
nor U1906 (N_1906,N_144,N_1189);
and U1907 (N_1907,N_277,N_650);
nand U1908 (N_1908,N_1047,N_1215);
xnor U1909 (N_1909,N_583,N_692);
nor U1910 (N_1910,N_629,N_857);
or U1911 (N_1911,N_787,N_614);
nor U1912 (N_1912,N_977,N_602);
and U1913 (N_1913,N_635,N_447);
or U1914 (N_1914,N_876,N_1138);
xor U1915 (N_1915,N_203,N_747);
nand U1916 (N_1916,N_1146,N_1066);
and U1917 (N_1917,N_1087,N_1221);
or U1918 (N_1918,N_729,N_1033);
xor U1919 (N_1919,N_1224,N_902);
xor U1920 (N_1920,N_532,N_862);
nand U1921 (N_1921,N_370,N_581);
xnor U1922 (N_1922,N_935,N_898);
nor U1923 (N_1923,N_338,N_332);
and U1924 (N_1924,N_398,N_222);
nand U1925 (N_1925,N_1229,N_819);
xor U1926 (N_1926,N_1049,N_838);
nand U1927 (N_1927,N_543,N_1222);
nand U1928 (N_1928,N_240,N_144);
or U1929 (N_1929,N_104,N_946);
and U1930 (N_1930,N_591,N_645);
or U1931 (N_1931,N_378,N_767);
nor U1932 (N_1932,N_654,N_1201);
nand U1933 (N_1933,N_55,N_677);
and U1934 (N_1934,N_372,N_504);
nor U1935 (N_1935,N_1222,N_444);
xnor U1936 (N_1936,N_802,N_332);
xor U1937 (N_1937,N_896,N_199);
and U1938 (N_1938,N_1084,N_390);
or U1939 (N_1939,N_1198,N_399);
and U1940 (N_1940,N_685,N_893);
and U1941 (N_1941,N_3,N_1020);
and U1942 (N_1942,N_579,N_231);
or U1943 (N_1943,N_747,N_649);
nor U1944 (N_1944,N_48,N_596);
nand U1945 (N_1945,N_438,N_875);
xor U1946 (N_1946,N_1060,N_630);
or U1947 (N_1947,N_1055,N_71);
and U1948 (N_1948,N_275,N_594);
or U1949 (N_1949,N_459,N_784);
and U1950 (N_1950,N_101,N_1227);
nand U1951 (N_1951,N_69,N_1047);
or U1952 (N_1952,N_741,N_985);
xor U1953 (N_1953,N_1130,N_236);
or U1954 (N_1954,N_401,N_213);
nand U1955 (N_1955,N_1247,N_154);
xor U1956 (N_1956,N_748,N_624);
xnor U1957 (N_1957,N_833,N_819);
nand U1958 (N_1958,N_712,N_1247);
xnor U1959 (N_1959,N_398,N_1138);
xnor U1960 (N_1960,N_359,N_250);
or U1961 (N_1961,N_719,N_562);
or U1962 (N_1962,N_906,N_1042);
or U1963 (N_1963,N_777,N_625);
xnor U1964 (N_1964,N_52,N_664);
or U1965 (N_1965,N_1206,N_1006);
and U1966 (N_1966,N_1041,N_475);
nand U1967 (N_1967,N_401,N_123);
nor U1968 (N_1968,N_79,N_1128);
or U1969 (N_1969,N_331,N_155);
nand U1970 (N_1970,N_952,N_310);
and U1971 (N_1971,N_454,N_881);
and U1972 (N_1972,N_351,N_988);
xor U1973 (N_1973,N_677,N_217);
or U1974 (N_1974,N_907,N_531);
nor U1975 (N_1975,N_95,N_149);
or U1976 (N_1976,N_1023,N_206);
xnor U1977 (N_1977,N_611,N_607);
nand U1978 (N_1978,N_770,N_1181);
or U1979 (N_1979,N_978,N_306);
nand U1980 (N_1980,N_39,N_1168);
or U1981 (N_1981,N_766,N_149);
nor U1982 (N_1982,N_295,N_534);
xor U1983 (N_1983,N_627,N_734);
and U1984 (N_1984,N_12,N_158);
xor U1985 (N_1985,N_320,N_166);
xnor U1986 (N_1986,N_863,N_922);
nand U1987 (N_1987,N_163,N_1229);
nand U1988 (N_1988,N_745,N_640);
or U1989 (N_1989,N_668,N_416);
nand U1990 (N_1990,N_97,N_473);
or U1991 (N_1991,N_254,N_614);
nor U1992 (N_1992,N_1212,N_837);
or U1993 (N_1993,N_1091,N_182);
or U1994 (N_1994,N_25,N_62);
nor U1995 (N_1995,N_1058,N_984);
xnor U1996 (N_1996,N_626,N_465);
xor U1997 (N_1997,N_594,N_824);
nand U1998 (N_1998,N_511,N_998);
or U1999 (N_1999,N_1019,N_134);
nand U2000 (N_2000,N_859,N_322);
xnor U2001 (N_2001,N_1052,N_1200);
and U2002 (N_2002,N_1242,N_424);
nand U2003 (N_2003,N_724,N_1071);
xor U2004 (N_2004,N_1054,N_869);
xnor U2005 (N_2005,N_361,N_172);
nor U2006 (N_2006,N_1103,N_197);
or U2007 (N_2007,N_834,N_1186);
or U2008 (N_2008,N_628,N_576);
nor U2009 (N_2009,N_77,N_703);
nand U2010 (N_2010,N_1100,N_175);
xor U2011 (N_2011,N_688,N_254);
and U2012 (N_2012,N_1012,N_965);
nor U2013 (N_2013,N_341,N_1009);
xnor U2014 (N_2014,N_1132,N_492);
nand U2015 (N_2015,N_952,N_917);
nor U2016 (N_2016,N_92,N_45);
nor U2017 (N_2017,N_872,N_538);
nand U2018 (N_2018,N_686,N_103);
and U2019 (N_2019,N_124,N_688);
and U2020 (N_2020,N_159,N_339);
xnor U2021 (N_2021,N_650,N_496);
xor U2022 (N_2022,N_885,N_65);
and U2023 (N_2023,N_1233,N_382);
nand U2024 (N_2024,N_1116,N_223);
xnor U2025 (N_2025,N_625,N_548);
nand U2026 (N_2026,N_9,N_104);
and U2027 (N_2027,N_368,N_196);
xnor U2028 (N_2028,N_445,N_153);
nand U2029 (N_2029,N_14,N_1246);
nand U2030 (N_2030,N_501,N_996);
and U2031 (N_2031,N_397,N_345);
xnor U2032 (N_2032,N_863,N_134);
and U2033 (N_2033,N_585,N_13);
and U2034 (N_2034,N_399,N_879);
and U2035 (N_2035,N_470,N_287);
and U2036 (N_2036,N_1186,N_260);
nand U2037 (N_2037,N_1224,N_622);
xor U2038 (N_2038,N_561,N_961);
xnor U2039 (N_2039,N_546,N_1192);
nor U2040 (N_2040,N_512,N_949);
xnor U2041 (N_2041,N_326,N_1198);
and U2042 (N_2042,N_5,N_174);
or U2043 (N_2043,N_960,N_317);
or U2044 (N_2044,N_899,N_489);
xor U2045 (N_2045,N_239,N_171);
nor U2046 (N_2046,N_1132,N_1086);
nor U2047 (N_2047,N_987,N_392);
or U2048 (N_2048,N_897,N_659);
nor U2049 (N_2049,N_1013,N_225);
nor U2050 (N_2050,N_786,N_321);
nand U2051 (N_2051,N_524,N_822);
nand U2052 (N_2052,N_418,N_853);
nor U2053 (N_2053,N_866,N_1227);
and U2054 (N_2054,N_443,N_477);
nand U2055 (N_2055,N_333,N_502);
or U2056 (N_2056,N_1079,N_735);
xnor U2057 (N_2057,N_208,N_885);
nor U2058 (N_2058,N_367,N_1162);
nand U2059 (N_2059,N_1019,N_469);
nand U2060 (N_2060,N_912,N_1092);
xnor U2061 (N_2061,N_823,N_731);
nand U2062 (N_2062,N_387,N_38);
nand U2063 (N_2063,N_1008,N_382);
or U2064 (N_2064,N_812,N_456);
nor U2065 (N_2065,N_1083,N_780);
nor U2066 (N_2066,N_193,N_929);
nor U2067 (N_2067,N_596,N_423);
xnor U2068 (N_2068,N_885,N_327);
or U2069 (N_2069,N_624,N_315);
or U2070 (N_2070,N_489,N_1178);
xnor U2071 (N_2071,N_424,N_433);
xor U2072 (N_2072,N_757,N_67);
nand U2073 (N_2073,N_1101,N_749);
and U2074 (N_2074,N_286,N_574);
or U2075 (N_2075,N_1119,N_48);
xor U2076 (N_2076,N_502,N_511);
nand U2077 (N_2077,N_336,N_1182);
and U2078 (N_2078,N_346,N_997);
nor U2079 (N_2079,N_98,N_840);
or U2080 (N_2080,N_835,N_1209);
xnor U2081 (N_2081,N_448,N_871);
xor U2082 (N_2082,N_477,N_1194);
nor U2083 (N_2083,N_415,N_1238);
and U2084 (N_2084,N_971,N_353);
nand U2085 (N_2085,N_1083,N_481);
nor U2086 (N_2086,N_1122,N_148);
or U2087 (N_2087,N_806,N_358);
nand U2088 (N_2088,N_323,N_594);
and U2089 (N_2089,N_487,N_966);
xnor U2090 (N_2090,N_437,N_215);
nand U2091 (N_2091,N_621,N_1172);
nand U2092 (N_2092,N_517,N_288);
nand U2093 (N_2093,N_993,N_387);
or U2094 (N_2094,N_562,N_557);
and U2095 (N_2095,N_742,N_355);
nand U2096 (N_2096,N_652,N_1083);
or U2097 (N_2097,N_860,N_537);
nand U2098 (N_2098,N_49,N_955);
nor U2099 (N_2099,N_1073,N_464);
xor U2100 (N_2100,N_278,N_873);
nand U2101 (N_2101,N_148,N_623);
xnor U2102 (N_2102,N_1143,N_488);
and U2103 (N_2103,N_1000,N_834);
nor U2104 (N_2104,N_442,N_648);
xnor U2105 (N_2105,N_618,N_445);
or U2106 (N_2106,N_794,N_1079);
xor U2107 (N_2107,N_275,N_687);
and U2108 (N_2108,N_250,N_726);
and U2109 (N_2109,N_32,N_1166);
nor U2110 (N_2110,N_323,N_948);
and U2111 (N_2111,N_512,N_788);
nor U2112 (N_2112,N_976,N_576);
nand U2113 (N_2113,N_1208,N_997);
xnor U2114 (N_2114,N_1034,N_2);
nor U2115 (N_2115,N_94,N_481);
or U2116 (N_2116,N_1081,N_403);
nand U2117 (N_2117,N_85,N_256);
xor U2118 (N_2118,N_17,N_782);
nand U2119 (N_2119,N_153,N_1012);
and U2120 (N_2120,N_244,N_1104);
nor U2121 (N_2121,N_862,N_1136);
nand U2122 (N_2122,N_1178,N_909);
and U2123 (N_2123,N_424,N_305);
xnor U2124 (N_2124,N_1223,N_710);
nand U2125 (N_2125,N_579,N_748);
and U2126 (N_2126,N_846,N_244);
and U2127 (N_2127,N_1240,N_840);
nor U2128 (N_2128,N_353,N_960);
xor U2129 (N_2129,N_101,N_431);
xor U2130 (N_2130,N_389,N_377);
nand U2131 (N_2131,N_52,N_174);
nand U2132 (N_2132,N_586,N_204);
xor U2133 (N_2133,N_1188,N_747);
xor U2134 (N_2134,N_476,N_1048);
xnor U2135 (N_2135,N_471,N_422);
xnor U2136 (N_2136,N_307,N_234);
nor U2137 (N_2137,N_1175,N_349);
or U2138 (N_2138,N_586,N_1136);
xor U2139 (N_2139,N_815,N_174);
xor U2140 (N_2140,N_1206,N_465);
nor U2141 (N_2141,N_890,N_235);
nand U2142 (N_2142,N_1056,N_1145);
or U2143 (N_2143,N_738,N_230);
nor U2144 (N_2144,N_294,N_648);
xor U2145 (N_2145,N_969,N_1102);
nand U2146 (N_2146,N_518,N_1010);
nand U2147 (N_2147,N_785,N_52);
nor U2148 (N_2148,N_450,N_162);
xnor U2149 (N_2149,N_71,N_1024);
and U2150 (N_2150,N_456,N_849);
nor U2151 (N_2151,N_27,N_603);
nor U2152 (N_2152,N_471,N_377);
nor U2153 (N_2153,N_864,N_1233);
and U2154 (N_2154,N_924,N_1214);
or U2155 (N_2155,N_1223,N_470);
nor U2156 (N_2156,N_18,N_540);
and U2157 (N_2157,N_403,N_1047);
and U2158 (N_2158,N_261,N_213);
or U2159 (N_2159,N_608,N_958);
nor U2160 (N_2160,N_92,N_122);
and U2161 (N_2161,N_502,N_1002);
nor U2162 (N_2162,N_1039,N_65);
and U2163 (N_2163,N_141,N_1137);
nand U2164 (N_2164,N_1218,N_531);
or U2165 (N_2165,N_1106,N_771);
and U2166 (N_2166,N_882,N_585);
nor U2167 (N_2167,N_258,N_651);
nor U2168 (N_2168,N_307,N_1231);
or U2169 (N_2169,N_60,N_1055);
nor U2170 (N_2170,N_707,N_1236);
and U2171 (N_2171,N_520,N_1108);
or U2172 (N_2172,N_630,N_334);
nor U2173 (N_2173,N_351,N_777);
xor U2174 (N_2174,N_805,N_60);
nand U2175 (N_2175,N_308,N_15);
xor U2176 (N_2176,N_889,N_906);
xnor U2177 (N_2177,N_943,N_45);
xor U2178 (N_2178,N_61,N_1058);
nor U2179 (N_2179,N_497,N_112);
nand U2180 (N_2180,N_537,N_567);
and U2181 (N_2181,N_25,N_170);
and U2182 (N_2182,N_667,N_198);
nand U2183 (N_2183,N_463,N_529);
and U2184 (N_2184,N_288,N_890);
nor U2185 (N_2185,N_8,N_154);
nor U2186 (N_2186,N_1195,N_628);
nor U2187 (N_2187,N_485,N_33);
nand U2188 (N_2188,N_616,N_979);
xnor U2189 (N_2189,N_200,N_669);
or U2190 (N_2190,N_987,N_99);
nor U2191 (N_2191,N_259,N_3);
nor U2192 (N_2192,N_1072,N_128);
nor U2193 (N_2193,N_778,N_898);
nand U2194 (N_2194,N_1172,N_967);
and U2195 (N_2195,N_1043,N_288);
xor U2196 (N_2196,N_22,N_989);
and U2197 (N_2197,N_607,N_60);
nand U2198 (N_2198,N_5,N_648);
or U2199 (N_2199,N_218,N_594);
nor U2200 (N_2200,N_432,N_392);
nand U2201 (N_2201,N_272,N_128);
or U2202 (N_2202,N_182,N_932);
and U2203 (N_2203,N_1010,N_476);
and U2204 (N_2204,N_399,N_428);
xor U2205 (N_2205,N_1081,N_511);
and U2206 (N_2206,N_144,N_1164);
xnor U2207 (N_2207,N_675,N_3);
or U2208 (N_2208,N_417,N_379);
and U2209 (N_2209,N_418,N_180);
nand U2210 (N_2210,N_722,N_230);
nand U2211 (N_2211,N_1180,N_785);
or U2212 (N_2212,N_1202,N_419);
or U2213 (N_2213,N_764,N_762);
nor U2214 (N_2214,N_833,N_473);
xnor U2215 (N_2215,N_1009,N_1035);
and U2216 (N_2216,N_255,N_540);
xnor U2217 (N_2217,N_229,N_684);
nor U2218 (N_2218,N_48,N_342);
nor U2219 (N_2219,N_644,N_960);
nand U2220 (N_2220,N_1077,N_480);
or U2221 (N_2221,N_108,N_206);
and U2222 (N_2222,N_469,N_873);
nand U2223 (N_2223,N_143,N_123);
xor U2224 (N_2224,N_956,N_301);
nor U2225 (N_2225,N_613,N_251);
nand U2226 (N_2226,N_96,N_1170);
nor U2227 (N_2227,N_231,N_528);
and U2228 (N_2228,N_105,N_977);
nor U2229 (N_2229,N_1106,N_1045);
nor U2230 (N_2230,N_491,N_257);
and U2231 (N_2231,N_785,N_499);
nand U2232 (N_2232,N_266,N_265);
nand U2233 (N_2233,N_880,N_593);
nor U2234 (N_2234,N_773,N_137);
nor U2235 (N_2235,N_961,N_496);
nand U2236 (N_2236,N_44,N_633);
nor U2237 (N_2237,N_94,N_681);
and U2238 (N_2238,N_21,N_406);
xnor U2239 (N_2239,N_486,N_814);
nor U2240 (N_2240,N_982,N_209);
or U2241 (N_2241,N_1166,N_298);
xor U2242 (N_2242,N_481,N_676);
or U2243 (N_2243,N_1170,N_109);
nor U2244 (N_2244,N_273,N_994);
or U2245 (N_2245,N_494,N_32);
xnor U2246 (N_2246,N_183,N_467);
or U2247 (N_2247,N_822,N_1177);
nor U2248 (N_2248,N_937,N_949);
or U2249 (N_2249,N_1054,N_803);
or U2250 (N_2250,N_222,N_1016);
and U2251 (N_2251,N_1188,N_923);
nand U2252 (N_2252,N_704,N_430);
xnor U2253 (N_2253,N_512,N_457);
nor U2254 (N_2254,N_775,N_747);
nor U2255 (N_2255,N_687,N_155);
nand U2256 (N_2256,N_1192,N_624);
and U2257 (N_2257,N_55,N_557);
nor U2258 (N_2258,N_873,N_1123);
or U2259 (N_2259,N_1165,N_1206);
nand U2260 (N_2260,N_404,N_208);
xor U2261 (N_2261,N_541,N_945);
or U2262 (N_2262,N_249,N_491);
and U2263 (N_2263,N_582,N_34);
or U2264 (N_2264,N_103,N_1160);
xor U2265 (N_2265,N_437,N_963);
nor U2266 (N_2266,N_44,N_700);
and U2267 (N_2267,N_1134,N_197);
or U2268 (N_2268,N_63,N_599);
nand U2269 (N_2269,N_1045,N_407);
nand U2270 (N_2270,N_1224,N_1040);
nand U2271 (N_2271,N_1121,N_1108);
or U2272 (N_2272,N_647,N_833);
nor U2273 (N_2273,N_738,N_1040);
nor U2274 (N_2274,N_809,N_415);
nor U2275 (N_2275,N_187,N_994);
xnor U2276 (N_2276,N_984,N_591);
xnor U2277 (N_2277,N_823,N_553);
and U2278 (N_2278,N_252,N_178);
nand U2279 (N_2279,N_475,N_77);
xor U2280 (N_2280,N_263,N_626);
and U2281 (N_2281,N_1178,N_66);
nand U2282 (N_2282,N_13,N_688);
nand U2283 (N_2283,N_580,N_1120);
nand U2284 (N_2284,N_239,N_837);
and U2285 (N_2285,N_1234,N_702);
nor U2286 (N_2286,N_1124,N_403);
and U2287 (N_2287,N_292,N_684);
nand U2288 (N_2288,N_1216,N_1217);
and U2289 (N_2289,N_1194,N_658);
nand U2290 (N_2290,N_967,N_557);
xnor U2291 (N_2291,N_646,N_526);
nor U2292 (N_2292,N_911,N_1134);
nand U2293 (N_2293,N_691,N_525);
xnor U2294 (N_2294,N_892,N_756);
nand U2295 (N_2295,N_737,N_500);
xor U2296 (N_2296,N_364,N_373);
nand U2297 (N_2297,N_295,N_339);
xnor U2298 (N_2298,N_521,N_821);
and U2299 (N_2299,N_1147,N_97);
nor U2300 (N_2300,N_299,N_916);
and U2301 (N_2301,N_947,N_647);
xor U2302 (N_2302,N_1248,N_215);
and U2303 (N_2303,N_157,N_16);
or U2304 (N_2304,N_1076,N_541);
xnor U2305 (N_2305,N_768,N_974);
and U2306 (N_2306,N_985,N_272);
or U2307 (N_2307,N_1017,N_527);
xor U2308 (N_2308,N_716,N_743);
or U2309 (N_2309,N_937,N_818);
nor U2310 (N_2310,N_0,N_743);
or U2311 (N_2311,N_843,N_765);
nand U2312 (N_2312,N_927,N_573);
nor U2313 (N_2313,N_571,N_590);
nor U2314 (N_2314,N_1099,N_1);
nand U2315 (N_2315,N_747,N_586);
nor U2316 (N_2316,N_733,N_206);
or U2317 (N_2317,N_636,N_981);
and U2318 (N_2318,N_638,N_1190);
or U2319 (N_2319,N_406,N_985);
xnor U2320 (N_2320,N_514,N_222);
and U2321 (N_2321,N_987,N_1149);
xnor U2322 (N_2322,N_1001,N_439);
nor U2323 (N_2323,N_138,N_104);
or U2324 (N_2324,N_758,N_1183);
xor U2325 (N_2325,N_809,N_896);
and U2326 (N_2326,N_127,N_996);
nor U2327 (N_2327,N_686,N_1008);
nor U2328 (N_2328,N_1058,N_41);
nor U2329 (N_2329,N_267,N_1209);
nor U2330 (N_2330,N_262,N_399);
xor U2331 (N_2331,N_382,N_939);
nor U2332 (N_2332,N_671,N_885);
nor U2333 (N_2333,N_390,N_176);
nor U2334 (N_2334,N_432,N_939);
nand U2335 (N_2335,N_1085,N_529);
nor U2336 (N_2336,N_1137,N_642);
and U2337 (N_2337,N_622,N_1199);
nand U2338 (N_2338,N_1113,N_928);
nand U2339 (N_2339,N_355,N_713);
or U2340 (N_2340,N_1002,N_415);
or U2341 (N_2341,N_946,N_1019);
or U2342 (N_2342,N_341,N_1064);
nor U2343 (N_2343,N_1075,N_1035);
and U2344 (N_2344,N_5,N_146);
or U2345 (N_2345,N_729,N_779);
and U2346 (N_2346,N_111,N_1004);
and U2347 (N_2347,N_417,N_20);
and U2348 (N_2348,N_68,N_62);
or U2349 (N_2349,N_1173,N_168);
xor U2350 (N_2350,N_1009,N_79);
xnor U2351 (N_2351,N_635,N_1109);
xnor U2352 (N_2352,N_576,N_306);
or U2353 (N_2353,N_321,N_946);
nor U2354 (N_2354,N_1023,N_892);
or U2355 (N_2355,N_337,N_1227);
or U2356 (N_2356,N_55,N_20);
nor U2357 (N_2357,N_850,N_1241);
and U2358 (N_2358,N_378,N_301);
nand U2359 (N_2359,N_1132,N_1119);
and U2360 (N_2360,N_521,N_922);
nor U2361 (N_2361,N_674,N_22);
and U2362 (N_2362,N_1162,N_311);
xor U2363 (N_2363,N_1080,N_198);
or U2364 (N_2364,N_364,N_631);
xor U2365 (N_2365,N_1140,N_42);
xnor U2366 (N_2366,N_167,N_530);
and U2367 (N_2367,N_510,N_1093);
xor U2368 (N_2368,N_806,N_995);
nor U2369 (N_2369,N_896,N_58);
xnor U2370 (N_2370,N_614,N_1131);
nand U2371 (N_2371,N_797,N_860);
nor U2372 (N_2372,N_652,N_281);
xor U2373 (N_2373,N_471,N_476);
and U2374 (N_2374,N_1094,N_1111);
nand U2375 (N_2375,N_961,N_774);
and U2376 (N_2376,N_133,N_83);
nand U2377 (N_2377,N_939,N_143);
xor U2378 (N_2378,N_832,N_1056);
or U2379 (N_2379,N_1022,N_331);
and U2380 (N_2380,N_681,N_123);
and U2381 (N_2381,N_774,N_736);
nand U2382 (N_2382,N_1100,N_525);
xnor U2383 (N_2383,N_1057,N_834);
nand U2384 (N_2384,N_811,N_380);
or U2385 (N_2385,N_1123,N_562);
nand U2386 (N_2386,N_1128,N_973);
xor U2387 (N_2387,N_81,N_166);
nand U2388 (N_2388,N_158,N_168);
xnor U2389 (N_2389,N_1130,N_114);
nand U2390 (N_2390,N_626,N_439);
or U2391 (N_2391,N_1077,N_333);
and U2392 (N_2392,N_446,N_807);
nor U2393 (N_2393,N_895,N_1101);
nor U2394 (N_2394,N_575,N_1233);
and U2395 (N_2395,N_1094,N_478);
and U2396 (N_2396,N_474,N_585);
or U2397 (N_2397,N_107,N_150);
xnor U2398 (N_2398,N_954,N_485);
nor U2399 (N_2399,N_984,N_352);
nand U2400 (N_2400,N_803,N_548);
or U2401 (N_2401,N_315,N_676);
nor U2402 (N_2402,N_835,N_253);
nor U2403 (N_2403,N_15,N_394);
xor U2404 (N_2404,N_1110,N_848);
xnor U2405 (N_2405,N_478,N_491);
and U2406 (N_2406,N_427,N_805);
or U2407 (N_2407,N_168,N_1084);
or U2408 (N_2408,N_1139,N_928);
or U2409 (N_2409,N_611,N_721);
or U2410 (N_2410,N_858,N_851);
and U2411 (N_2411,N_780,N_1167);
xnor U2412 (N_2412,N_223,N_205);
or U2413 (N_2413,N_147,N_746);
or U2414 (N_2414,N_692,N_186);
nand U2415 (N_2415,N_1129,N_912);
or U2416 (N_2416,N_6,N_1213);
nand U2417 (N_2417,N_550,N_970);
and U2418 (N_2418,N_1132,N_717);
xnor U2419 (N_2419,N_631,N_620);
nand U2420 (N_2420,N_822,N_708);
or U2421 (N_2421,N_1188,N_1036);
nand U2422 (N_2422,N_31,N_662);
xnor U2423 (N_2423,N_798,N_208);
and U2424 (N_2424,N_1012,N_541);
nand U2425 (N_2425,N_562,N_413);
nor U2426 (N_2426,N_886,N_1081);
and U2427 (N_2427,N_596,N_403);
or U2428 (N_2428,N_923,N_17);
nand U2429 (N_2429,N_1153,N_679);
nand U2430 (N_2430,N_932,N_415);
and U2431 (N_2431,N_520,N_937);
nor U2432 (N_2432,N_22,N_718);
nor U2433 (N_2433,N_400,N_284);
xnor U2434 (N_2434,N_705,N_231);
and U2435 (N_2435,N_982,N_108);
nor U2436 (N_2436,N_1080,N_756);
and U2437 (N_2437,N_952,N_185);
nand U2438 (N_2438,N_1154,N_378);
nor U2439 (N_2439,N_487,N_669);
nand U2440 (N_2440,N_651,N_1239);
nor U2441 (N_2441,N_313,N_1123);
nand U2442 (N_2442,N_360,N_1008);
xor U2443 (N_2443,N_840,N_918);
nand U2444 (N_2444,N_1220,N_1007);
nand U2445 (N_2445,N_712,N_299);
and U2446 (N_2446,N_561,N_742);
and U2447 (N_2447,N_673,N_759);
nand U2448 (N_2448,N_843,N_583);
nand U2449 (N_2449,N_427,N_1117);
xnor U2450 (N_2450,N_841,N_41);
or U2451 (N_2451,N_658,N_239);
nor U2452 (N_2452,N_442,N_1193);
or U2453 (N_2453,N_226,N_849);
or U2454 (N_2454,N_942,N_380);
and U2455 (N_2455,N_223,N_1122);
nor U2456 (N_2456,N_392,N_339);
xor U2457 (N_2457,N_798,N_802);
nor U2458 (N_2458,N_766,N_951);
and U2459 (N_2459,N_1170,N_246);
xor U2460 (N_2460,N_7,N_408);
nand U2461 (N_2461,N_364,N_1219);
nor U2462 (N_2462,N_993,N_330);
and U2463 (N_2463,N_101,N_1004);
and U2464 (N_2464,N_627,N_317);
or U2465 (N_2465,N_217,N_567);
and U2466 (N_2466,N_830,N_725);
xor U2467 (N_2467,N_99,N_799);
xnor U2468 (N_2468,N_333,N_250);
nand U2469 (N_2469,N_1192,N_1129);
nor U2470 (N_2470,N_260,N_489);
nor U2471 (N_2471,N_1209,N_691);
nor U2472 (N_2472,N_1185,N_1132);
or U2473 (N_2473,N_718,N_788);
and U2474 (N_2474,N_520,N_823);
nor U2475 (N_2475,N_478,N_950);
nor U2476 (N_2476,N_686,N_804);
or U2477 (N_2477,N_1055,N_254);
nor U2478 (N_2478,N_728,N_619);
xor U2479 (N_2479,N_820,N_495);
nand U2480 (N_2480,N_58,N_705);
nand U2481 (N_2481,N_553,N_357);
and U2482 (N_2482,N_1055,N_924);
and U2483 (N_2483,N_1227,N_310);
xor U2484 (N_2484,N_823,N_697);
nor U2485 (N_2485,N_657,N_738);
nor U2486 (N_2486,N_670,N_52);
and U2487 (N_2487,N_554,N_340);
nor U2488 (N_2488,N_74,N_418);
or U2489 (N_2489,N_937,N_960);
nand U2490 (N_2490,N_518,N_117);
or U2491 (N_2491,N_71,N_128);
or U2492 (N_2492,N_969,N_740);
or U2493 (N_2493,N_260,N_66);
nor U2494 (N_2494,N_400,N_1041);
nor U2495 (N_2495,N_272,N_919);
nor U2496 (N_2496,N_539,N_1077);
and U2497 (N_2497,N_1106,N_82);
or U2498 (N_2498,N_774,N_177);
and U2499 (N_2499,N_426,N_1110);
xor U2500 (N_2500,N_2377,N_1419);
nor U2501 (N_2501,N_1856,N_2100);
nor U2502 (N_2502,N_1936,N_2246);
xor U2503 (N_2503,N_1942,N_2494);
nor U2504 (N_2504,N_1945,N_2256);
xnor U2505 (N_2505,N_1576,N_1747);
xnor U2506 (N_2506,N_2031,N_1263);
or U2507 (N_2507,N_1264,N_1486);
xnor U2508 (N_2508,N_1331,N_1421);
nand U2509 (N_2509,N_1451,N_2417);
and U2510 (N_2510,N_1581,N_2185);
and U2511 (N_2511,N_1535,N_2002);
xor U2512 (N_2512,N_1575,N_2281);
nor U2513 (N_2513,N_2141,N_1358);
nand U2514 (N_2514,N_1333,N_1403);
nor U2515 (N_2515,N_1366,N_2387);
nand U2516 (N_2516,N_2467,N_1391);
nand U2517 (N_2517,N_1834,N_1422);
xnor U2518 (N_2518,N_1554,N_2403);
nand U2519 (N_2519,N_1696,N_2086);
or U2520 (N_2520,N_2145,N_2419);
nor U2521 (N_2521,N_1356,N_1322);
xor U2522 (N_2522,N_1935,N_1347);
and U2523 (N_2523,N_1296,N_1888);
or U2524 (N_2524,N_2139,N_1976);
nor U2525 (N_2525,N_1710,N_1843);
or U2526 (N_2526,N_2429,N_2069);
nor U2527 (N_2527,N_2395,N_1655);
nor U2528 (N_2528,N_2216,N_1519);
or U2529 (N_2529,N_1574,N_2340);
xnor U2530 (N_2530,N_2114,N_1932);
and U2531 (N_2531,N_2226,N_1266);
nor U2532 (N_2532,N_1878,N_1408);
nor U2533 (N_2533,N_2346,N_1648);
or U2534 (N_2534,N_2336,N_1405);
xnor U2535 (N_2535,N_2365,N_1619);
xor U2536 (N_2536,N_1795,N_2268);
nor U2537 (N_2537,N_1534,N_2455);
or U2538 (N_2538,N_1427,N_1555);
nand U2539 (N_2539,N_1917,N_2280);
or U2540 (N_2540,N_1773,N_2442);
nand U2541 (N_2541,N_2112,N_2271);
nor U2542 (N_2542,N_1270,N_1305);
nor U2543 (N_2543,N_1780,N_1662);
nand U2544 (N_2544,N_2229,N_2394);
or U2545 (N_2545,N_2083,N_1991);
nand U2546 (N_2546,N_2287,N_2372);
nand U2547 (N_2547,N_2208,N_1384);
and U2548 (N_2548,N_2016,N_2361);
nor U2549 (N_2549,N_1453,N_1595);
and U2550 (N_2550,N_1349,N_1560);
and U2551 (N_2551,N_1415,N_2279);
nand U2552 (N_2552,N_1321,N_1869);
or U2553 (N_2553,N_2151,N_2286);
nand U2554 (N_2554,N_1596,N_1489);
and U2555 (N_2555,N_2096,N_2276);
xor U2556 (N_2556,N_2113,N_2356);
nand U2557 (N_2557,N_2202,N_2483);
or U2558 (N_2558,N_1533,N_1964);
nor U2559 (N_2559,N_1372,N_1731);
xnor U2560 (N_2560,N_1685,N_1737);
nor U2561 (N_2561,N_1549,N_1606);
nand U2562 (N_2562,N_2485,N_2265);
xnor U2563 (N_2563,N_1804,N_1918);
nor U2564 (N_2564,N_1371,N_2027);
xnor U2565 (N_2565,N_1440,N_1849);
and U2566 (N_2566,N_2009,N_2349);
nor U2567 (N_2567,N_1874,N_2401);
or U2568 (N_2568,N_2073,N_1610);
and U2569 (N_2569,N_2160,N_2149);
nand U2570 (N_2570,N_1317,N_2228);
nand U2571 (N_2571,N_1570,N_1407);
or U2572 (N_2572,N_1944,N_1703);
nand U2573 (N_2573,N_2253,N_1877);
or U2574 (N_2574,N_2457,N_1414);
and U2575 (N_2575,N_1520,N_1452);
and U2576 (N_2576,N_1522,N_2317);
or U2577 (N_2577,N_2423,N_1857);
xor U2578 (N_2578,N_1307,N_1251);
nand U2579 (N_2579,N_1492,N_1390);
xnor U2580 (N_2580,N_2306,N_1341);
nor U2581 (N_2581,N_1736,N_2464);
and U2582 (N_2582,N_1751,N_2375);
and U2583 (N_2583,N_1272,N_2488);
and U2584 (N_2584,N_1679,N_2410);
and U2585 (N_2585,N_1521,N_2045);
or U2586 (N_2586,N_2376,N_2320);
or U2587 (N_2587,N_1608,N_1280);
or U2588 (N_2588,N_2043,N_2050);
xor U2589 (N_2589,N_1496,N_1503);
nand U2590 (N_2590,N_1873,N_2334);
or U2591 (N_2591,N_1424,N_2000);
or U2592 (N_2592,N_2180,N_2108);
xor U2593 (N_2593,N_1962,N_1882);
nand U2594 (N_2594,N_2104,N_1892);
nand U2595 (N_2595,N_1512,N_1690);
or U2596 (N_2596,N_2332,N_1338);
and U2597 (N_2597,N_2269,N_1664);
xnor U2598 (N_2598,N_2218,N_1768);
and U2599 (N_2599,N_1707,N_1536);
nand U2600 (N_2600,N_1926,N_1631);
nand U2601 (N_2601,N_1837,N_2299);
xor U2602 (N_2602,N_1516,N_2267);
nand U2603 (N_2603,N_2446,N_2222);
nand U2604 (N_2604,N_2352,N_1661);
nor U2605 (N_2605,N_2040,N_1819);
or U2606 (N_2606,N_1865,N_2188);
xnor U2607 (N_2607,N_2278,N_1671);
nor U2608 (N_2608,N_1968,N_1459);
nor U2609 (N_2609,N_1404,N_2316);
or U2610 (N_2610,N_2437,N_1430);
nor U2611 (N_2611,N_1981,N_1934);
nor U2612 (N_2612,N_1916,N_2155);
nand U2613 (N_2613,N_2059,N_1590);
or U2614 (N_2614,N_1276,N_2170);
and U2615 (N_2615,N_1584,N_2262);
and U2616 (N_2616,N_1941,N_1591);
or U2617 (N_2617,N_1268,N_2416);
nand U2618 (N_2618,N_2243,N_2017);
and U2619 (N_2619,N_2033,N_1914);
nor U2620 (N_2620,N_1250,N_2138);
and U2621 (N_2621,N_1547,N_1624);
nor U2622 (N_2622,N_1706,N_1855);
nand U2623 (N_2623,N_1365,N_1497);
xnor U2624 (N_2624,N_1684,N_2065);
nor U2625 (N_2625,N_2072,N_1744);
and U2626 (N_2626,N_1670,N_2301);
nor U2627 (N_2627,N_2178,N_1495);
and U2628 (N_2628,N_1604,N_2110);
or U2629 (N_2629,N_1899,N_1688);
xor U2630 (N_2630,N_1472,N_2198);
nand U2631 (N_2631,N_2289,N_2475);
nand U2632 (N_2632,N_2004,N_2470);
and U2633 (N_2633,N_2166,N_2194);
xnor U2634 (N_2634,N_1695,N_2380);
nand U2635 (N_2635,N_1359,N_2184);
nand U2636 (N_2636,N_1805,N_1894);
xor U2637 (N_2637,N_1312,N_1548);
or U2638 (N_2638,N_1434,N_2205);
xor U2639 (N_2639,N_1638,N_2121);
nand U2640 (N_2640,N_1327,N_1694);
xor U2641 (N_2641,N_1676,N_2117);
or U2642 (N_2642,N_1513,N_1388);
xnor U2643 (N_2643,N_1600,N_1309);
xnor U2644 (N_2644,N_1754,N_1642);
or U2645 (N_2645,N_1890,N_2408);
or U2646 (N_2646,N_1789,N_2133);
and U2647 (N_2647,N_2374,N_1902);
and U2648 (N_2648,N_1973,N_1858);
and U2649 (N_2649,N_2235,N_1637);
or U2650 (N_2650,N_1514,N_1314);
xor U2651 (N_2651,N_1719,N_1546);
xor U2652 (N_2652,N_2263,N_1470);
nor U2653 (N_2653,N_1720,N_1779);
nor U2654 (N_2654,N_1903,N_1368);
or U2655 (N_2655,N_1727,N_2313);
and U2656 (N_2656,N_2127,N_2061);
nand U2657 (N_2657,N_1807,N_2319);
nand U2658 (N_2658,N_1313,N_1846);
xor U2659 (N_2659,N_1871,N_2252);
nor U2660 (N_2660,N_2146,N_2163);
nor U2661 (N_2661,N_2456,N_1675);
or U2662 (N_2662,N_2438,N_1836);
xnor U2663 (N_2663,N_1303,N_2147);
and U2664 (N_2664,N_2323,N_2026);
or U2665 (N_2665,N_2199,N_1788);
nand U2666 (N_2666,N_1911,N_1850);
and U2667 (N_2667,N_1288,N_1258);
nand U2668 (N_2668,N_2118,N_1699);
nand U2669 (N_2669,N_2079,N_1545);
and U2670 (N_2670,N_1940,N_1443);
nand U2671 (N_2671,N_2052,N_1448);
nand U2672 (N_2672,N_1929,N_1820);
nand U2673 (N_2673,N_1983,N_1401);
xor U2674 (N_2674,N_2240,N_1515);
xor U2675 (N_2675,N_1588,N_2122);
nand U2676 (N_2676,N_1783,N_1668);
nand U2677 (N_2677,N_1647,N_1646);
nand U2678 (N_2678,N_1881,N_2115);
nand U2679 (N_2679,N_1801,N_1396);
nand U2680 (N_2680,N_2157,N_1697);
nand U2681 (N_2681,N_1848,N_1884);
nor U2682 (N_2682,N_1798,N_2030);
and U2683 (N_2683,N_1989,N_2035);
nor U2684 (N_2684,N_2053,N_1580);
nor U2685 (N_2685,N_1920,N_1399);
xnor U2686 (N_2686,N_1665,N_1825);
nor U2687 (N_2687,N_2359,N_2249);
nor U2688 (N_2688,N_1910,N_2328);
xor U2689 (N_2689,N_1666,N_1813);
or U2690 (N_2690,N_2099,N_1550);
nor U2691 (N_2691,N_1445,N_1352);
or U2692 (N_2692,N_1998,N_1502);
xnor U2693 (N_2693,N_1474,N_2389);
nor U2694 (N_2694,N_1669,N_1763);
and U2695 (N_2695,N_1660,N_2024);
nand U2696 (N_2696,N_1538,N_1335);
nor U2697 (N_2697,N_1708,N_1473);
or U2698 (N_2698,N_1650,N_2101);
xor U2699 (N_2699,N_2131,N_2036);
nand U2700 (N_2700,N_1378,N_2075);
or U2701 (N_2701,N_2368,N_2430);
or U2702 (N_2702,N_1829,N_1880);
nor U2703 (N_2703,N_1449,N_2493);
or U2704 (N_2704,N_2421,N_2227);
or U2705 (N_2705,N_2436,N_1735);
nor U2706 (N_2706,N_2225,N_1557);
nor U2707 (N_2707,N_1300,N_1394);
xnor U2708 (N_2708,N_1304,N_2007);
or U2709 (N_2709,N_2441,N_1893);
and U2710 (N_2710,N_1827,N_1283);
nand U2711 (N_2711,N_2171,N_1921);
and U2712 (N_2712,N_2070,N_2062);
or U2713 (N_2713,N_2080,N_1504);
and U2714 (N_2714,N_2324,N_2314);
nor U2715 (N_2715,N_2047,N_1809);
nand U2716 (N_2716,N_1797,N_1901);
or U2717 (N_2717,N_1839,N_1682);
and U2718 (N_2718,N_2244,N_2220);
and U2719 (N_2719,N_2284,N_2221);
nor U2720 (N_2720,N_2496,N_2382);
or U2721 (N_2721,N_1782,N_1762);
and U2722 (N_2722,N_1255,N_1528);
nand U2723 (N_2723,N_1386,N_2028);
or U2724 (N_2724,N_1506,N_2291);
nand U2725 (N_2725,N_1475,N_1566);
or U2726 (N_2726,N_2405,N_2452);
or U2727 (N_2727,N_2048,N_1992);
xnor U2728 (N_2728,N_1367,N_1308);
nor U2729 (N_2729,N_1537,N_2200);
nor U2730 (N_2730,N_1814,N_1416);
nor U2731 (N_2731,N_1994,N_1639);
nand U2732 (N_2732,N_1441,N_1320);
xor U2733 (N_2733,N_1274,N_2261);
xnor U2734 (N_2734,N_2169,N_1806);
or U2735 (N_2735,N_2362,N_1979);
and U2736 (N_2736,N_1818,N_1835);
nor U2737 (N_2737,N_1672,N_1567);
or U2738 (N_2738,N_2189,N_2137);
nor U2739 (N_2739,N_2272,N_2107);
nand U2740 (N_2740,N_1975,N_2491);
nand U2741 (N_2741,N_1879,N_2136);
xor U2742 (N_2742,N_1769,N_1479);
or U2743 (N_2743,N_2095,N_1716);
nand U2744 (N_2744,N_1598,N_2106);
or U2745 (N_2745,N_2415,N_2019);
xnor U2746 (N_2746,N_1812,N_1931);
xor U2747 (N_2747,N_2091,N_2130);
xor U2748 (N_2748,N_1776,N_2266);
or U2749 (N_2749,N_2449,N_2239);
xnor U2750 (N_2750,N_1722,N_1306);
nor U2751 (N_2751,N_2116,N_2119);
nand U2752 (N_2752,N_1411,N_1544);
and U2753 (N_2753,N_2302,N_2466);
nor U2754 (N_2754,N_2288,N_2411);
or U2755 (N_2755,N_2018,N_2105);
nand U2756 (N_2756,N_1483,N_1426);
xor U2757 (N_2757,N_1628,N_1420);
and U2758 (N_2758,N_1970,N_1718);
nor U2759 (N_2759,N_1605,N_2183);
nor U2760 (N_2760,N_1791,N_1558);
or U2761 (N_2761,N_1742,N_1490);
or U2762 (N_2762,N_1630,N_1252);
or U2763 (N_2763,N_2124,N_2078);
nor U2764 (N_2764,N_2495,N_1900);
xnor U2765 (N_2765,N_1949,N_1946);
or U2766 (N_2766,N_2233,N_2203);
xnor U2767 (N_2767,N_1374,N_1505);
nand U2768 (N_2768,N_2406,N_1915);
xnor U2769 (N_2769,N_1644,N_1864);
nor U2770 (N_2770,N_1692,N_1480);
nand U2771 (N_2771,N_2103,N_1589);
and U2772 (N_2772,N_1417,N_2303);
or U2773 (N_2773,N_1267,N_2486);
or U2774 (N_2774,N_1875,N_1725);
xnor U2775 (N_2775,N_1568,N_2013);
nand U2776 (N_2776,N_1436,N_1923);
nor U2777 (N_2777,N_1913,N_1380);
nand U2778 (N_2778,N_2392,N_2335);
nand U2779 (N_2779,N_2168,N_1299);
nand U2780 (N_2780,N_1438,N_2498);
xor U2781 (N_2781,N_1621,N_2247);
xnor U2782 (N_2782,N_1767,N_2418);
nand U2783 (N_2783,N_2089,N_1641);
nand U2784 (N_2784,N_2309,N_2177);
nand U2785 (N_2785,N_1579,N_1526);
and U2786 (N_2786,N_1643,N_1543);
and U2787 (N_2787,N_2478,N_1799);
or U2788 (N_2788,N_1463,N_1966);
nor U2789 (N_2789,N_1289,N_2029);
and U2790 (N_2790,N_2399,N_2172);
nor U2791 (N_2791,N_2192,N_1573);
xnor U2792 (N_2792,N_1344,N_2046);
and U2793 (N_2793,N_1615,N_2426);
or U2794 (N_2794,N_2167,N_2162);
and U2795 (N_2795,N_1632,N_1393);
nand U2796 (N_2796,N_2329,N_2242);
nand U2797 (N_2797,N_1518,N_1285);
nand U2798 (N_2798,N_1753,N_1410);
xnor U2799 (N_2799,N_1866,N_2164);
or U2800 (N_2800,N_1260,N_2210);
xor U2801 (N_2801,N_1571,N_2125);
xnor U2802 (N_2802,N_1955,N_2409);
or U2803 (N_2803,N_1540,N_2388);
xnor U2804 (N_2804,N_2297,N_1928);
nor U2805 (N_2805,N_1948,N_1997);
nor U2806 (N_2806,N_2321,N_2427);
xnor U2807 (N_2807,N_1377,N_1723);
and U2808 (N_2808,N_1318,N_2412);
xnor U2809 (N_2809,N_2481,N_1265);
or U2810 (N_2810,N_2477,N_1823);
and U2811 (N_2811,N_1387,N_1721);
nor U2812 (N_2812,N_1509,N_1402);
xnor U2813 (N_2813,N_2443,N_2010);
nand U2814 (N_2814,N_2071,N_1468);
xnor U2815 (N_2815,N_1332,N_1481);
nand U2816 (N_2816,N_1974,N_2195);
xnor U2817 (N_2817,N_2087,N_1887);
nor U2818 (N_2818,N_1986,N_1634);
or U2819 (N_2819,N_1862,N_1397);
or U2820 (N_2820,N_1350,N_1587);
xor U2821 (N_2821,N_2311,N_2369);
and U2822 (N_2822,N_1833,N_2129);
nand U2823 (N_2823,N_1585,N_1398);
xnor U2824 (N_2824,N_1578,N_1821);
xor U2825 (N_2825,N_2090,N_1339);
xnor U2826 (N_2826,N_2230,N_1599);
or U2827 (N_2827,N_2021,N_1293);
or U2828 (N_2828,N_2003,N_1379);
and U2829 (N_2829,N_2440,N_2450);
and U2830 (N_2830,N_1277,N_1455);
nor U2831 (N_2831,N_1689,N_2219);
nor U2832 (N_2832,N_1746,N_1362);
or U2833 (N_2833,N_2039,N_2379);
xor U2834 (N_2834,N_1508,N_1625);
or U2835 (N_2835,N_1898,N_1532);
nand U2836 (N_2836,N_1654,N_1851);
nor U2837 (N_2837,N_1269,N_2055);
or U2838 (N_2838,N_2236,N_2420);
xnor U2839 (N_2839,N_1891,N_2092);
and U2840 (N_2840,N_2304,N_1925);
and U2841 (N_2841,N_2424,N_1466);
xor U2842 (N_2842,N_1844,N_2447);
and U2843 (N_2843,N_1781,N_1761);
or U2844 (N_2844,N_1256,N_2295);
xor U2845 (N_2845,N_1824,N_2294);
xnor U2846 (N_2846,N_1469,N_1556);
or U2847 (N_2847,N_1457,N_2479);
and U2848 (N_2848,N_2407,N_1413);
nand U2849 (N_2849,N_1484,N_2217);
or U2850 (N_2850,N_1343,N_2123);
nor U2851 (N_2851,N_2402,N_1889);
nand U2852 (N_2852,N_2468,N_1954);
and U2853 (N_2853,N_1253,N_1956);
nand U2854 (N_2854,N_2326,N_2474);
or U2855 (N_2855,N_2414,N_1450);
xnor U2856 (N_2856,N_2161,N_1467);
or U2857 (N_2857,N_1409,N_1896);
and U2858 (N_2858,N_2094,N_2081);
nor U2859 (N_2859,N_1461,N_1860);
or U2860 (N_2860,N_2153,N_1930);
or U2861 (N_2861,N_1883,N_1700);
nand U2862 (N_2862,N_2214,N_1802);
nand U2863 (N_2863,N_1912,N_1325);
xor U2864 (N_2864,N_2383,N_1524);
xor U2865 (N_2865,N_2197,N_2175);
and U2866 (N_2866,N_2282,N_2234);
nand U2867 (N_2867,N_1609,N_2384);
and U2868 (N_2868,N_1561,N_1577);
nor U2869 (N_2869,N_1478,N_2337);
xor U2870 (N_2870,N_1471,N_2260);
and U2871 (N_2871,N_2308,N_2032);
nand U2872 (N_2872,N_1678,N_2142);
nor U2873 (N_2873,N_2011,N_1686);
xor U2874 (N_2874,N_1297,N_1603);
or U2875 (N_2875,N_1510,N_2283);
nand U2876 (N_2876,N_1724,N_1759);
nand U2877 (N_2877,N_1740,N_2413);
and U2878 (N_2878,N_2355,N_2490);
or U2879 (N_2879,N_1563,N_2298);
nand U2880 (N_2880,N_1953,N_2274);
xnor U2881 (N_2881,N_1919,N_2255);
or U2882 (N_2882,N_2135,N_2425);
nor U2883 (N_2883,N_1456,N_2159);
and U2884 (N_2884,N_1831,N_2223);
nand U2885 (N_2885,N_2148,N_2093);
xor U2886 (N_2886,N_1950,N_1826);
or U2887 (N_2887,N_1363,N_2422);
nor U2888 (N_2888,N_1261,N_1464);
nand U2889 (N_2889,N_1663,N_2005);
or U2890 (N_2890,N_2275,N_1340);
nand U2891 (N_2891,N_1815,N_2499);
nand U2892 (N_2892,N_2128,N_2154);
and U2893 (N_2893,N_1760,N_1683);
or U2894 (N_2894,N_1967,N_1792);
or U2895 (N_2895,N_2034,N_2463);
xnor U2896 (N_2896,N_1730,N_1729);
xnor U2897 (N_2897,N_1704,N_2237);
xnor U2898 (N_2898,N_2398,N_2174);
xnor U2899 (N_2899,N_1987,N_2325);
and U2900 (N_2900,N_1922,N_1709);
or U2901 (N_2901,N_1476,N_1487);
or U2902 (N_2902,N_1658,N_2315);
nand U2903 (N_2903,N_1832,N_2434);
xnor U2904 (N_2904,N_2056,N_1257);
and U2905 (N_2905,N_2432,N_1418);
nor U2906 (N_2906,N_1488,N_1732);
nor U2907 (N_2907,N_1395,N_2396);
or U2908 (N_2908,N_1651,N_2182);
or U2909 (N_2909,N_1500,N_1342);
nand U2910 (N_2910,N_1381,N_1301);
nand U2911 (N_2911,N_1785,N_1714);
nand U2912 (N_2912,N_2391,N_1817);
nor U2913 (N_2913,N_2015,N_1254);
nor U2914 (N_2914,N_1771,N_1593);
nor U2915 (N_2915,N_1530,N_2001);
or U2916 (N_2916,N_2371,N_2085);
or U2917 (N_2917,N_1758,N_1959);
nand U2918 (N_2918,N_2204,N_2357);
nor U2919 (N_2919,N_2254,N_2473);
nand U2920 (N_2920,N_2097,N_1870);
and U2921 (N_2921,N_1961,N_1601);
nand U2922 (N_2922,N_1446,N_2126);
or U2923 (N_2923,N_2064,N_1906);
nand U2924 (N_2924,N_2454,N_1262);
nor U2925 (N_2925,N_2270,N_2067);
nor U2926 (N_2926,N_1863,N_1659);
xnor U2927 (N_2927,N_2179,N_2176);
or U2928 (N_2928,N_1310,N_2259);
nand U2929 (N_2929,N_1995,N_1373);
xor U2930 (N_2930,N_1745,N_2331);
nand U2931 (N_2931,N_2076,N_1947);
nand U2932 (N_2932,N_1594,N_1969);
xor U2933 (N_2933,N_2480,N_2385);
xor U2934 (N_2934,N_1636,N_1432);
nand U2935 (N_2935,N_1757,N_2386);
nand U2936 (N_2936,N_1282,N_1793);
and U2937 (N_2937,N_1938,N_1984);
and U2938 (N_2938,N_2196,N_1551);
nor U2939 (N_2939,N_2292,N_1431);
nor U2940 (N_2940,N_2111,N_2333);
nand U2941 (N_2941,N_1626,N_1868);
nand U2942 (N_2942,N_1750,N_1529);
or U2943 (N_2943,N_2381,N_2134);
or U2944 (N_2944,N_2150,N_2460);
xor U2945 (N_2945,N_1400,N_1982);
and U2946 (N_2946,N_2343,N_1978);
nand U2947 (N_2947,N_1354,N_2212);
nand U2948 (N_2948,N_1677,N_2211);
nor U2949 (N_2949,N_1392,N_1988);
nor U2950 (N_2950,N_2393,N_1645);
and U2951 (N_2951,N_1369,N_1774);
nor U2952 (N_2952,N_1351,N_1927);
nand U2953 (N_2953,N_1957,N_1298);
or U2954 (N_2954,N_1749,N_1437);
nor U2955 (N_2955,N_1712,N_2193);
and U2956 (N_2956,N_1733,N_2458);
nand U2957 (N_2957,N_2140,N_2354);
and U2958 (N_2958,N_1958,N_2042);
and U2959 (N_2959,N_2310,N_2060);
nor U2960 (N_2960,N_1796,N_2238);
xor U2961 (N_2961,N_2305,N_2487);
xor U2962 (N_2962,N_2472,N_1383);
nor U2963 (N_2963,N_1433,N_1853);
and U2964 (N_2964,N_1360,N_1429);
or U2965 (N_2965,N_1370,N_1702);
nor U2966 (N_2966,N_2264,N_1943);
or U2967 (N_2967,N_2186,N_1275);
nand U2968 (N_2968,N_1681,N_1498);
and U2969 (N_2969,N_2348,N_1290);
xnor U2970 (N_2970,N_2300,N_1653);
nor U2971 (N_2971,N_1965,N_2257);
and U2972 (N_2972,N_2444,N_2258);
nand U2973 (N_2973,N_2435,N_1353);
and U2974 (N_2974,N_1477,N_2058);
nor U2975 (N_2975,N_1786,N_1511);
xor U2976 (N_2976,N_1302,N_1259);
and U2977 (N_2977,N_1627,N_1346);
and U2978 (N_2978,N_2373,N_2025);
nor U2979 (N_2979,N_1273,N_1617);
or U2980 (N_2980,N_1939,N_2431);
nand U2981 (N_2981,N_2339,N_1531);
nor U2982 (N_2982,N_2277,N_2482);
nand U2983 (N_2983,N_1523,N_1442);
nand U2984 (N_2984,N_1784,N_1385);
nand U2985 (N_2985,N_2489,N_1990);
nand U2986 (N_2986,N_1582,N_1465);
nor U2987 (N_2987,N_1854,N_1326);
nor U2988 (N_2988,N_1376,N_1772);
nor U2989 (N_2989,N_1541,N_1775);
xnor U2990 (N_2990,N_1717,N_1838);
xor U2991 (N_2991,N_1425,N_2345);
and U2992 (N_2992,N_2063,N_2181);
or U2993 (N_2993,N_1607,N_1565);
and U2994 (N_2994,N_2293,N_2158);
nor U2995 (N_2995,N_2492,N_1808);
nor U2996 (N_2996,N_2451,N_2465);
xor U2997 (N_2997,N_1324,N_1960);
and U2998 (N_2998,N_1357,N_2132);
nand U2999 (N_2999,N_1454,N_2173);
xnor U3000 (N_3000,N_1375,N_2037);
and U3001 (N_3001,N_1527,N_2307);
nor U3002 (N_3002,N_2088,N_1909);
nor U3003 (N_3003,N_1328,N_1897);
xnor U3004 (N_3004,N_1423,N_1777);
and U3005 (N_3005,N_2344,N_1564);
and U3006 (N_3006,N_1618,N_2459);
or U3007 (N_3007,N_1462,N_1382);
nand U3008 (N_3008,N_1652,N_2312);
and U3009 (N_3009,N_1355,N_1972);
nand U3010 (N_3010,N_1755,N_2044);
and U3011 (N_3011,N_1766,N_1840);
nor U3012 (N_3012,N_2120,N_1583);
nand U3013 (N_3013,N_2008,N_1623);
nor U3014 (N_3014,N_1517,N_1345);
or U3015 (N_3015,N_1287,N_1491);
nor U3016 (N_3016,N_2360,N_2250);
xnor U3017 (N_3017,N_1592,N_1715);
nand U3018 (N_3018,N_2453,N_1810);
xor U3019 (N_3019,N_2012,N_2342);
xnor U3020 (N_3020,N_2206,N_2248);
nor U3021 (N_3021,N_1364,N_1905);
xor U3022 (N_3022,N_2209,N_1572);
xnor U3023 (N_3023,N_2351,N_1842);
or U3024 (N_3024,N_1734,N_1933);
nor U3025 (N_3025,N_2006,N_2051);
or U3026 (N_3026,N_1728,N_1635);
nand U3027 (N_3027,N_1691,N_2400);
or U3028 (N_3028,N_1811,N_2187);
and U3029 (N_3029,N_1867,N_1616);
xnor U3030 (N_3030,N_1316,N_1698);
or U3031 (N_3031,N_1447,N_1501);
and U3032 (N_3032,N_1389,N_1971);
and U3033 (N_3033,N_1952,N_1284);
and U3034 (N_3034,N_1999,N_1907);
nor U3035 (N_3035,N_1680,N_1713);
nand U3036 (N_3036,N_1552,N_1741);
and U3037 (N_3037,N_2367,N_1859);
xor U3038 (N_3038,N_1886,N_2366);
and U3039 (N_3039,N_1794,N_2433);
or U3040 (N_3040,N_1361,N_1336);
or U3041 (N_3041,N_1752,N_1649);
xor U3042 (N_3042,N_2165,N_1611);
xnor U3043 (N_3043,N_2448,N_2143);
or U3044 (N_3044,N_2102,N_1319);
and U3045 (N_3045,N_1569,N_1330);
or U3046 (N_3046,N_2190,N_1493);
xor U3047 (N_3047,N_1485,N_1701);
nor U3048 (N_3048,N_1444,N_1861);
nand U3049 (N_3049,N_2077,N_1525);
nand U3050 (N_3050,N_1673,N_2144);
nand U3051 (N_3051,N_1559,N_1311);
or U3052 (N_3052,N_1281,N_2338);
xnor U3053 (N_3053,N_2341,N_2327);
xor U3054 (N_3054,N_2484,N_2378);
or U3055 (N_3055,N_1993,N_2404);
nor U3056 (N_3056,N_2156,N_2390);
xor U3057 (N_3057,N_1597,N_1904);
xnor U3058 (N_3058,N_1586,N_1937);
and U3059 (N_3059,N_1406,N_1614);
nand U3060 (N_3060,N_1800,N_1951);
xnor U3061 (N_3061,N_1778,N_1841);
nand U3062 (N_3062,N_1705,N_1602);
nand U3063 (N_3063,N_2022,N_1499);
xor U3064 (N_3064,N_1726,N_1790);
and U3065 (N_3065,N_1507,N_2370);
and U3066 (N_3066,N_1412,N_1674);
xor U3067 (N_3067,N_1872,N_1315);
xor U3068 (N_3068,N_2231,N_1553);
nor U3069 (N_3069,N_2353,N_2347);
nand U3070 (N_3070,N_1764,N_1739);
and U3071 (N_3071,N_1816,N_2014);
or U3072 (N_3072,N_2469,N_1787);
nand U3073 (N_3073,N_2215,N_2224);
xnor U3074 (N_3074,N_1985,N_1629);
nor U3075 (N_3075,N_2363,N_2038);
and U3076 (N_3076,N_1756,N_1458);
xor U3077 (N_3077,N_1830,N_2057);
or U3078 (N_3078,N_2241,N_2462);
xor U3079 (N_3079,N_1980,N_2068);
or U3080 (N_3080,N_1803,N_2054);
nand U3081 (N_3081,N_1852,N_2245);
nand U3082 (N_3082,N_1656,N_2066);
nand U3083 (N_3083,N_1908,N_1770);
xnor U3084 (N_3084,N_1334,N_2296);
xnor U3085 (N_3085,N_2476,N_1667);
nand U3086 (N_3086,N_2213,N_2207);
xor U3087 (N_3087,N_2497,N_1613);
nor U3088 (N_3088,N_1292,N_1828);
or U3089 (N_3089,N_2439,N_2471);
or U3090 (N_3090,N_1657,N_1885);
and U3091 (N_3091,N_2082,N_2041);
or U3092 (N_3092,N_2109,N_2251);
or U3093 (N_3093,N_2461,N_1977);
nor U3094 (N_3094,N_1748,N_2074);
xnor U3095 (N_3095,N_1963,N_1847);
xor U3096 (N_3096,N_1435,N_1765);
and U3097 (N_3097,N_1924,N_1822);
xnor U3098 (N_3098,N_1337,N_1460);
nor U3099 (N_3099,N_1539,N_1895);
nor U3100 (N_3100,N_2232,N_1542);
nor U3101 (N_3101,N_2428,N_2364);
nand U3102 (N_3102,N_1291,N_1294);
xnor U3103 (N_3103,N_2191,N_1348);
nor U3104 (N_3104,N_2358,N_2318);
nand U3105 (N_3105,N_1876,N_2020);
xnor U3106 (N_3106,N_1428,N_2445);
nor U3107 (N_3107,N_2098,N_2322);
and U3108 (N_3108,N_1279,N_2397);
xnor U3109 (N_3109,N_1612,N_1845);
nor U3110 (N_3110,N_2152,N_2330);
and U3111 (N_3111,N_1278,N_1693);
xnor U3112 (N_3112,N_2273,N_1633);
xnor U3113 (N_3113,N_2049,N_1439);
xor U3114 (N_3114,N_1738,N_1329);
nand U3115 (N_3115,N_1482,N_2285);
nand U3116 (N_3116,N_1494,N_1323);
nand U3117 (N_3117,N_1286,N_1295);
and U3118 (N_3118,N_1640,N_1620);
nand U3119 (N_3119,N_2290,N_1271);
or U3120 (N_3120,N_1711,N_2350);
nor U3121 (N_3121,N_1743,N_1996);
xnor U3122 (N_3122,N_2201,N_1687);
xnor U3123 (N_3123,N_1622,N_2084);
nor U3124 (N_3124,N_2023,N_1562);
nand U3125 (N_3125,N_1430,N_1397);
and U3126 (N_3126,N_2103,N_1651);
xnor U3127 (N_3127,N_1781,N_2192);
nor U3128 (N_3128,N_2078,N_1849);
nand U3129 (N_3129,N_1962,N_2034);
or U3130 (N_3130,N_2264,N_1915);
nand U3131 (N_3131,N_1696,N_1880);
and U3132 (N_3132,N_1943,N_1311);
and U3133 (N_3133,N_1774,N_1438);
and U3134 (N_3134,N_1343,N_1279);
nand U3135 (N_3135,N_1607,N_1971);
nor U3136 (N_3136,N_2268,N_2338);
nand U3137 (N_3137,N_2116,N_1444);
and U3138 (N_3138,N_2168,N_2289);
or U3139 (N_3139,N_1698,N_2307);
nor U3140 (N_3140,N_1914,N_2312);
nor U3141 (N_3141,N_1620,N_1572);
nor U3142 (N_3142,N_1609,N_2409);
nand U3143 (N_3143,N_1975,N_1844);
xnor U3144 (N_3144,N_1907,N_1631);
nand U3145 (N_3145,N_2259,N_1925);
nor U3146 (N_3146,N_2078,N_1795);
nor U3147 (N_3147,N_2431,N_2115);
nor U3148 (N_3148,N_1375,N_1508);
nor U3149 (N_3149,N_1277,N_2100);
and U3150 (N_3150,N_1926,N_1872);
or U3151 (N_3151,N_2101,N_1328);
and U3152 (N_3152,N_1791,N_1434);
and U3153 (N_3153,N_1679,N_1302);
xnor U3154 (N_3154,N_1447,N_1270);
xnor U3155 (N_3155,N_1409,N_2248);
and U3156 (N_3156,N_2422,N_1379);
xnor U3157 (N_3157,N_1631,N_1664);
xnor U3158 (N_3158,N_2076,N_2087);
nor U3159 (N_3159,N_2273,N_1660);
or U3160 (N_3160,N_1990,N_1523);
nand U3161 (N_3161,N_2086,N_1811);
nor U3162 (N_3162,N_2315,N_1891);
nand U3163 (N_3163,N_2148,N_2315);
and U3164 (N_3164,N_2488,N_1675);
nand U3165 (N_3165,N_1937,N_2220);
or U3166 (N_3166,N_2221,N_2085);
nand U3167 (N_3167,N_2251,N_1448);
xor U3168 (N_3168,N_2031,N_2426);
nor U3169 (N_3169,N_1453,N_2399);
nor U3170 (N_3170,N_1946,N_2354);
or U3171 (N_3171,N_1358,N_2029);
xnor U3172 (N_3172,N_1443,N_1551);
nor U3173 (N_3173,N_2051,N_1981);
nor U3174 (N_3174,N_2169,N_1258);
nand U3175 (N_3175,N_1911,N_2040);
nand U3176 (N_3176,N_1294,N_2117);
and U3177 (N_3177,N_1596,N_2065);
and U3178 (N_3178,N_1986,N_2070);
or U3179 (N_3179,N_2306,N_2416);
nand U3180 (N_3180,N_1926,N_1742);
nand U3181 (N_3181,N_1732,N_2017);
nand U3182 (N_3182,N_2117,N_2205);
nand U3183 (N_3183,N_2072,N_2343);
nor U3184 (N_3184,N_2418,N_2148);
and U3185 (N_3185,N_1714,N_2253);
nor U3186 (N_3186,N_1323,N_1970);
xnor U3187 (N_3187,N_2373,N_2161);
nand U3188 (N_3188,N_1429,N_2446);
and U3189 (N_3189,N_1913,N_2272);
xnor U3190 (N_3190,N_2078,N_1400);
nand U3191 (N_3191,N_2458,N_1975);
xor U3192 (N_3192,N_1530,N_2121);
or U3193 (N_3193,N_1552,N_2075);
nor U3194 (N_3194,N_2441,N_1486);
or U3195 (N_3195,N_1508,N_1565);
or U3196 (N_3196,N_1502,N_2244);
xor U3197 (N_3197,N_1340,N_2132);
nand U3198 (N_3198,N_1495,N_1831);
or U3199 (N_3199,N_1777,N_1753);
and U3200 (N_3200,N_2315,N_1780);
nor U3201 (N_3201,N_1988,N_1805);
xor U3202 (N_3202,N_1558,N_2278);
and U3203 (N_3203,N_2228,N_1662);
or U3204 (N_3204,N_2448,N_1345);
nand U3205 (N_3205,N_2057,N_1567);
or U3206 (N_3206,N_1391,N_1832);
xor U3207 (N_3207,N_1800,N_2057);
and U3208 (N_3208,N_1683,N_2218);
nand U3209 (N_3209,N_1575,N_2489);
or U3210 (N_3210,N_1843,N_1542);
xnor U3211 (N_3211,N_1672,N_2316);
nand U3212 (N_3212,N_1629,N_1979);
nand U3213 (N_3213,N_1739,N_1844);
and U3214 (N_3214,N_2201,N_1393);
xnor U3215 (N_3215,N_1622,N_2004);
and U3216 (N_3216,N_2407,N_1593);
nand U3217 (N_3217,N_2123,N_2373);
xnor U3218 (N_3218,N_2467,N_2412);
and U3219 (N_3219,N_1306,N_2188);
or U3220 (N_3220,N_2254,N_2343);
nor U3221 (N_3221,N_1698,N_1350);
and U3222 (N_3222,N_1697,N_1782);
or U3223 (N_3223,N_1578,N_2270);
xor U3224 (N_3224,N_1992,N_1842);
nor U3225 (N_3225,N_2328,N_2235);
and U3226 (N_3226,N_1479,N_1893);
xor U3227 (N_3227,N_2249,N_1344);
or U3228 (N_3228,N_1821,N_1651);
nand U3229 (N_3229,N_2467,N_2017);
xnor U3230 (N_3230,N_1423,N_2427);
xor U3231 (N_3231,N_1330,N_1718);
nand U3232 (N_3232,N_2378,N_1364);
nand U3233 (N_3233,N_1400,N_1755);
or U3234 (N_3234,N_1492,N_2415);
nand U3235 (N_3235,N_1695,N_1857);
or U3236 (N_3236,N_2468,N_2032);
and U3237 (N_3237,N_2025,N_1398);
xor U3238 (N_3238,N_2224,N_1525);
or U3239 (N_3239,N_1906,N_1287);
and U3240 (N_3240,N_2062,N_1250);
xor U3241 (N_3241,N_1443,N_2199);
or U3242 (N_3242,N_1507,N_2355);
nor U3243 (N_3243,N_2104,N_1940);
and U3244 (N_3244,N_2010,N_1774);
xor U3245 (N_3245,N_2238,N_2283);
nor U3246 (N_3246,N_1397,N_1769);
or U3247 (N_3247,N_1819,N_1503);
or U3248 (N_3248,N_1518,N_1757);
and U3249 (N_3249,N_2005,N_2202);
xnor U3250 (N_3250,N_2106,N_1288);
nor U3251 (N_3251,N_1801,N_1951);
xor U3252 (N_3252,N_2273,N_2020);
and U3253 (N_3253,N_2006,N_2133);
or U3254 (N_3254,N_2037,N_1381);
nor U3255 (N_3255,N_2219,N_2294);
nor U3256 (N_3256,N_1331,N_1608);
nand U3257 (N_3257,N_1508,N_1269);
or U3258 (N_3258,N_2064,N_2243);
or U3259 (N_3259,N_2265,N_1453);
xor U3260 (N_3260,N_1974,N_2037);
or U3261 (N_3261,N_2342,N_1722);
xor U3262 (N_3262,N_1549,N_1573);
or U3263 (N_3263,N_1631,N_1996);
and U3264 (N_3264,N_2461,N_1860);
nor U3265 (N_3265,N_2061,N_1792);
and U3266 (N_3266,N_1368,N_1593);
or U3267 (N_3267,N_1583,N_2216);
and U3268 (N_3268,N_1773,N_1542);
or U3269 (N_3269,N_2139,N_1773);
xnor U3270 (N_3270,N_2183,N_2073);
and U3271 (N_3271,N_1879,N_1371);
xor U3272 (N_3272,N_1672,N_2477);
and U3273 (N_3273,N_2297,N_1264);
or U3274 (N_3274,N_1560,N_1301);
and U3275 (N_3275,N_1513,N_1622);
and U3276 (N_3276,N_2047,N_1347);
xor U3277 (N_3277,N_2201,N_2220);
or U3278 (N_3278,N_1302,N_1514);
or U3279 (N_3279,N_1932,N_1281);
and U3280 (N_3280,N_2073,N_2259);
nand U3281 (N_3281,N_1856,N_1547);
and U3282 (N_3282,N_2441,N_1654);
xor U3283 (N_3283,N_2097,N_2476);
nor U3284 (N_3284,N_1576,N_2090);
nor U3285 (N_3285,N_1340,N_1572);
or U3286 (N_3286,N_2462,N_1808);
or U3287 (N_3287,N_2034,N_2115);
nand U3288 (N_3288,N_1645,N_2252);
nand U3289 (N_3289,N_1979,N_1635);
and U3290 (N_3290,N_2202,N_2077);
xor U3291 (N_3291,N_2261,N_2383);
and U3292 (N_3292,N_2136,N_1739);
xnor U3293 (N_3293,N_1580,N_2066);
or U3294 (N_3294,N_2209,N_1914);
xor U3295 (N_3295,N_1972,N_2216);
nand U3296 (N_3296,N_1250,N_2368);
xor U3297 (N_3297,N_1748,N_1255);
xor U3298 (N_3298,N_1601,N_2164);
nand U3299 (N_3299,N_2459,N_1544);
or U3300 (N_3300,N_1934,N_2124);
nor U3301 (N_3301,N_1325,N_1691);
or U3302 (N_3302,N_1761,N_2071);
nor U3303 (N_3303,N_1705,N_1786);
or U3304 (N_3304,N_2285,N_1831);
xor U3305 (N_3305,N_1933,N_1508);
nor U3306 (N_3306,N_1604,N_1832);
nand U3307 (N_3307,N_1899,N_2206);
and U3308 (N_3308,N_1637,N_2437);
or U3309 (N_3309,N_2265,N_1396);
nor U3310 (N_3310,N_2164,N_1480);
nor U3311 (N_3311,N_2188,N_1423);
and U3312 (N_3312,N_2092,N_1449);
and U3313 (N_3313,N_1730,N_2362);
and U3314 (N_3314,N_2019,N_1551);
nand U3315 (N_3315,N_1807,N_1689);
or U3316 (N_3316,N_1999,N_2123);
and U3317 (N_3317,N_2354,N_1783);
or U3318 (N_3318,N_2285,N_1900);
and U3319 (N_3319,N_2392,N_1314);
or U3320 (N_3320,N_2339,N_2299);
nand U3321 (N_3321,N_2412,N_1326);
xnor U3322 (N_3322,N_1384,N_1460);
nand U3323 (N_3323,N_2273,N_1976);
xnor U3324 (N_3324,N_1804,N_2285);
or U3325 (N_3325,N_1924,N_1514);
and U3326 (N_3326,N_1489,N_2154);
or U3327 (N_3327,N_1620,N_1292);
and U3328 (N_3328,N_1552,N_1821);
xnor U3329 (N_3329,N_1390,N_2252);
or U3330 (N_3330,N_1649,N_2242);
nor U3331 (N_3331,N_1342,N_2346);
and U3332 (N_3332,N_2196,N_2100);
nand U3333 (N_3333,N_2150,N_1900);
and U3334 (N_3334,N_1607,N_1277);
xnor U3335 (N_3335,N_1620,N_1706);
and U3336 (N_3336,N_2303,N_1344);
or U3337 (N_3337,N_1721,N_1298);
xor U3338 (N_3338,N_1638,N_1258);
xnor U3339 (N_3339,N_1802,N_1904);
nand U3340 (N_3340,N_1513,N_1718);
nor U3341 (N_3341,N_1393,N_1641);
nand U3342 (N_3342,N_1836,N_1826);
and U3343 (N_3343,N_2172,N_2211);
nand U3344 (N_3344,N_2471,N_2293);
xnor U3345 (N_3345,N_1633,N_2185);
xnor U3346 (N_3346,N_2011,N_1495);
and U3347 (N_3347,N_2146,N_1532);
and U3348 (N_3348,N_1691,N_2466);
and U3349 (N_3349,N_1575,N_1788);
nand U3350 (N_3350,N_2305,N_1796);
and U3351 (N_3351,N_1555,N_2265);
nand U3352 (N_3352,N_1466,N_1269);
xor U3353 (N_3353,N_1881,N_2496);
or U3354 (N_3354,N_1868,N_1743);
nor U3355 (N_3355,N_1981,N_2014);
and U3356 (N_3356,N_2063,N_1512);
and U3357 (N_3357,N_1583,N_1543);
nor U3358 (N_3358,N_2339,N_1564);
nand U3359 (N_3359,N_1667,N_2359);
or U3360 (N_3360,N_1408,N_2256);
and U3361 (N_3361,N_2073,N_1320);
or U3362 (N_3362,N_1428,N_1503);
nand U3363 (N_3363,N_2291,N_1661);
and U3364 (N_3364,N_1881,N_2405);
nand U3365 (N_3365,N_1729,N_1288);
or U3366 (N_3366,N_2043,N_2264);
or U3367 (N_3367,N_1918,N_2373);
nor U3368 (N_3368,N_2498,N_1816);
or U3369 (N_3369,N_1782,N_1530);
nor U3370 (N_3370,N_1837,N_2305);
and U3371 (N_3371,N_1736,N_2002);
and U3372 (N_3372,N_2175,N_1645);
xnor U3373 (N_3373,N_1672,N_2076);
and U3374 (N_3374,N_1434,N_1471);
or U3375 (N_3375,N_2083,N_2402);
and U3376 (N_3376,N_1820,N_1275);
and U3377 (N_3377,N_2439,N_1428);
or U3378 (N_3378,N_1424,N_2409);
or U3379 (N_3379,N_2221,N_2029);
xnor U3380 (N_3380,N_1713,N_1491);
nor U3381 (N_3381,N_2094,N_2082);
nand U3382 (N_3382,N_2420,N_1500);
nand U3383 (N_3383,N_1791,N_1501);
xnor U3384 (N_3384,N_1447,N_2409);
nand U3385 (N_3385,N_1917,N_1392);
nor U3386 (N_3386,N_1824,N_2368);
nor U3387 (N_3387,N_1863,N_2066);
and U3388 (N_3388,N_2098,N_1895);
nor U3389 (N_3389,N_1478,N_2100);
and U3390 (N_3390,N_1988,N_1839);
nor U3391 (N_3391,N_1436,N_1391);
or U3392 (N_3392,N_1456,N_2461);
and U3393 (N_3393,N_1468,N_1828);
nor U3394 (N_3394,N_1718,N_1656);
xor U3395 (N_3395,N_1743,N_2074);
and U3396 (N_3396,N_2023,N_1344);
nand U3397 (N_3397,N_1288,N_2448);
and U3398 (N_3398,N_1725,N_1685);
nor U3399 (N_3399,N_2497,N_1421);
and U3400 (N_3400,N_1660,N_1629);
or U3401 (N_3401,N_1857,N_2030);
xnor U3402 (N_3402,N_1368,N_1825);
nand U3403 (N_3403,N_2300,N_1976);
nand U3404 (N_3404,N_1621,N_1838);
and U3405 (N_3405,N_1407,N_1636);
xor U3406 (N_3406,N_1445,N_1432);
and U3407 (N_3407,N_1882,N_2044);
and U3408 (N_3408,N_2200,N_2218);
nor U3409 (N_3409,N_1646,N_1798);
nand U3410 (N_3410,N_1669,N_2069);
or U3411 (N_3411,N_1418,N_1978);
nand U3412 (N_3412,N_1811,N_1871);
or U3413 (N_3413,N_2335,N_1877);
and U3414 (N_3414,N_1963,N_1635);
and U3415 (N_3415,N_1982,N_1403);
or U3416 (N_3416,N_2103,N_2385);
or U3417 (N_3417,N_2010,N_2002);
xor U3418 (N_3418,N_1286,N_1721);
or U3419 (N_3419,N_1587,N_2428);
and U3420 (N_3420,N_2021,N_1554);
nand U3421 (N_3421,N_2141,N_1288);
nor U3422 (N_3422,N_1785,N_2190);
nor U3423 (N_3423,N_1908,N_1309);
or U3424 (N_3424,N_2095,N_2119);
nand U3425 (N_3425,N_2068,N_2198);
or U3426 (N_3426,N_2469,N_1878);
or U3427 (N_3427,N_1959,N_1906);
and U3428 (N_3428,N_1474,N_1821);
nor U3429 (N_3429,N_1295,N_1353);
or U3430 (N_3430,N_2134,N_1561);
or U3431 (N_3431,N_1642,N_2132);
nor U3432 (N_3432,N_2255,N_1431);
nand U3433 (N_3433,N_1946,N_2353);
nor U3434 (N_3434,N_1612,N_1379);
xnor U3435 (N_3435,N_2059,N_2232);
nor U3436 (N_3436,N_2346,N_2253);
or U3437 (N_3437,N_1808,N_2223);
xnor U3438 (N_3438,N_1521,N_2039);
nand U3439 (N_3439,N_1685,N_2497);
nor U3440 (N_3440,N_2406,N_2402);
or U3441 (N_3441,N_2056,N_1473);
xor U3442 (N_3442,N_1953,N_1880);
xnor U3443 (N_3443,N_1595,N_1765);
nand U3444 (N_3444,N_2299,N_2420);
nand U3445 (N_3445,N_2294,N_1299);
or U3446 (N_3446,N_1471,N_1503);
xnor U3447 (N_3447,N_1493,N_1611);
nand U3448 (N_3448,N_1618,N_2421);
nand U3449 (N_3449,N_2248,N_2234);
nand U3450 (N_3450,N_2381,N_1850);
nand U3451 (N_3451,N_1335,N_1871);
or U3452 (N_3452,N_1297,N_2322);
nor U3453 (N_3453,N_1520,N_2371);
nand U3454 (N_3454,N_1337,N_1970);
nor U3455 (N_3455,N_1844,N_1919);
nor U3456 (N_3456,N_2380,N_1755);
nor U3457 (N_3457,N_1714,N_1363);
nand U3458 (N_3458,N_1885,N_1731);
or U3459 (N_3459,N_2469,N_1732);
nor U3460 (N_3460,N_1913,N_2289);
xnor U3461 (N_3461,N_1404,N_1569);
or U3462 (N_3462,N_2136,N_2312);
and U3463 (N_3463,N_1508,N_2361);
or U3464 (N_3464,N_2071,N_2070);
or U3465 (N_3465,N_1958,N_2252);
xor U3466 (N_3466,N_1330,N_1428);
xnor U3467 (N_3467,N_1392,N_2059);
nor U3468 (N_3468,N_2377,N_1380);
and U3469 (N_3469,N_2488,N_2485);
xnor U3470 (N_3470,N_1670,N_2178);
or U3471 (N_3471,N_1422,N_1673);
or U3472 (N_3472,N_1650,N_1868);
nor U3473 (N_3473,N_2013,N_1902);
nor U3474 (N_3474,N_2024,N_1465);
nand U3475 (N_3475,N_1650,N_2084);
nor U3476 (N_3476,N_1592,N_1402);
and U3477 (N_3477,N_1506,N_1422);
nand U3478 (N_3478,N_1859,N_1837);
and U3479 (N_3479,N_2209,N_2419);
and U3480 (N_3480,N_2115,N_2085);
or U3481 (N_3481,N_1690,N_2195);
and U3482 (N_3482,N_1986,N_2158);
nand U3483 (N_3483,N_1981,N_1288);
nor U3484 (N_3484,N_1946,N_2171);
nor U3485 (N_3485,N_2255,N_2112);
nand U3486 (N_3486,N_1318,N_1718);
xnor U3487 (N_3487,N_1253,N_2123);
nand U3488 (N_3488,N_1821,N_1440);
and U3489 (N_3489,N_1570,N_1744);
nand U3490 (N_3490,N_1601,N_1401);
and U3491 (N_3491,N_1624,N_2046);
or U3492 (N_3492,N_1381,N_1609);
xor U3493 (N_3493,N_2195,N_1674);
and U3494 (N_3494,N_2386,N_1535);
xnor U3495 (N_3495,N_1591,N_1985);
nand U3496 (N_3496,N_1447,N_1872);
xor U3497 (N_3497,N_1431,N_2439);
or U3498 (N_3498,N_1688,N_2440);
xnor U3499 (N_3499,N_1436,N_1687);
nand U3500 (N_3500,N_1581,N_2422);
or U3501 (N_3501,N_1759,N_2404);
xor U3502 (N_3502,N_2242,N_1663);
nor U3503 (N_3503,N_2058,N_1758);
or U3504 (N_3504,N_1685,N_1463);
and U3505 (N_3505,N_1929,N_1446);
nand U3506 (N_3506,N_2160,N_1967);
and U3507 (N_3507,N_1317,N_2127);
nor U3508 (N_3508,N_2481,N_2348);
or U3509 (N_3509,N_2044,N_1792);
xnor U3510 (N_3510,N_2493,N_1606);
or U3511 (N_3511,N_1865,N_2364);
xor U3512 (N_3512,N_2418,N_2279);
and U3513 (N_3513,N_2092,N_2444);
or U3514 (N_3514,N_2490,N_2185);
and U3515 (N_3515,N_2260,N_1842);
xnor U3516 (N_3516,N_1594,N_1367);
and U3517 (N_3517,N_1353,N_1316);
nor U3518 (N_3518,N_2435,N_1762);
and U3519 (N_3519,N_1391,N_1427);
or U3520 (N_3520,N_1281,N_1832);
xor U3521 (N_3521,N_1537,N_1989);
or U3522 (N_3522,N_1551,N_2121);
or U3523 (N_3523,N_1845,N_1973);
xnor U3524 (N_3524,N_1255,N_1666);
and U3525 (N_3525,N_1908,N_2141);
nor U3526 (N_3526,N_1597,N_1454);
xnor U3527 (N_3527,N_1656,N_1860);
and U3528 (N_3528,N_1893,N_2034);
and U3529 (N_3529,N_1806,N_1370);
and U3530 (N_3530,N_1534,N_1275);
nand U3531 (N_3531,N_2259,N_1492);
and U3532 (N_3532,N_1647,N_2109);
nor U3533 (N_3533,N_1308,N_1452);
or U3534 (N_3534,N_1625,N_1895);
or U3535 (N_3535,N_2037,N_1481);
and U3536 (N_3536,N_1470,N_2072);
nor U3537 (N_3537,N_1472,N_2169);
xnor U3538 (N_3538,N_1833,N_1649);
nor U3539 (N_3539,N_1858,N_1507);
nand U3540 (N_3540,N_1875,N_1389);
nor U3541 (N_3541,N_2171,N_1496);
nand U3542 (N_3542,N_2356,N_1720);
xnor U3543 (N_3543,N_1336,N_1725);
or U3544 (N_3544,N_2342,N_2042);
xor U3545 (N_3545,N_2059,N_2098);
or U3546 (N_3546,N_2160,N_2209);
nor U3547 (N_3547,N_1958,N_1587);
nor U3548 (N_3548,N_1793,N_1967);
and U3549 (N_3549,N_1439,N_1883);
or U3550 (N_3550,N_1987,N_1652);
and U3551 (N_3551,N_2151,N_1603);
nand U3552 (N_3552,N_1706,N_2264);
nor U3553 (N_3553,N_1892,N_2454);
xnor U3554 (N_3554,N_2093,N_1562);
nand U3555 (N_3555,N_1814,N_2015);
and U3556 (N_3556,N_2357,N_1420);
nand U3557 (N_3557,N_2072,N_1833);
or U3558 (N_3558,N_1872,N_1999);
nor U3559 (N_3559,N_1914,N_2458);
nor U3560 (N_3560,N_1646,N_1642);
or U3561 (N_3561,N_1426,N_1920);
xnor U3562 (N_3562,N_1609,N_1451);
nand U3563 (N_3563,N_1881,N_1981);
nand U3564 (N_3564,N_1732,N_2468);
or U3565 (N_3565,N_1992,N_2358);
nor U3566 (N_3566,N_2323,N_1653);
nor U3567 (N_3567,N_1953,N_2316);
nand U3568 (N_3568,N_1961,N_2273);
nand U3569 (N_3569,N_2355,N_1312);
xnor U3570 (N_3570,N_2286,N_1661);
nor U3571 (N_3571,N_2414,N_2135);
or U3572 (N_3572,N_1695,N_2119);
and U3573 (N_3573,N_1902,N_1561);
nand U3574 (N_3574,N_2232,N_1830);
xor U3575 (N_3575,N_2477,N_1349);
nand U3576 (N_3576,N_2053,N_2100);
and U3577 (N_3577,N_2376,N_2378);
xor U3578 (N_3578,N_2145,N_2138);
xor U3579 (N_3579,N_1656,N_1763);
and U3580 (N_3580,N_1622,N_1767);
or U3581 (N_3581,N_1346,N_2391);
and U3582 (N_3582,N_2106,N_1959);
and U3583 (N_3583,N_1947,N_2296);
nand U3584 (N_3584,N_1714,N_1923);
or U3585 (N_3585,N_1875,N_2454);
xor U3586 (N_3586,N_1494,N_2271);
xor U3587 (N_3587,N_1705,N_1960);
xor U3588 (N_3588,N_1312,N_1822);
nand U3589 (N_3589,N_1920,N_2259);
or U3590 (N_3590,N_1537,N_1464);
nand U3591 (N_3591,N_2333,N_1909);
nand U3592 (N_3592,N_1474,N_1360);
nor U3593 (N_3593,N_1424,N_2020);
or U3594 (N_3594,N_2234,N_2428);
and U3595 (N_3595,N_1502,N_2190);
and U3596 (N_3596,N_1728,N_1792);
or U3597 (N_3597,N_2342,N_1534);
xor U3598 (N_3598,N_1927,N_1919);
and U3599 (N_3599,N_1316,N_2080);
and U3600 (N_3600,N_1938,N_1729);
and U3601 (N_3601,N_1880,N_2049);
or U3602 (N_3602,N_1488,N_1288);
xnor U3603 (N_3603,N_1351,N_2265);
and U3604 (N_3604,N_1915,N_2341);
or U3605 (N_3605,N_1665,N_1606);
nor U3606 (N_3606,N_1784,N_2216);
or U3607 (N_3607,N_2481,N_1691);
and U3608 (N_3608,N_1314,N_2039);
nand U3609 (N_3609,N_2155,N_1796);
xor U3610 (N_3610,N_1521,N_1647);
and U3611 (N_3611,N_1303,N_1651);
and U3612 (N_3612,N_1774,N_2325);
xnor U3613 (N_3613,N_1451,N_1450);
nor U3614 (N_3614,N_2123,N_2026);
nor U3615 (N_3615,N_2413,N_2023);
xor U3616 (N_3616,N_1325,N_1606);
or U3617 (N_3617,N_1436,N_1704);
or U3618 (N_3618,N_2071,N_1469);
and U3619 (N_3619,N_2014,N_1644);
and U3620 (N_3620,N_1481,N_1619);
or U3621 (N_3621,N_1536,N_1417);
xor U3622 (N_3622,N_2373,N_2003);
nor U3623 (N_3623,N_1503,N_1294);
nor U3624 (N_3624,N_1753,N_1759);
nand U3625 (N_3625,N_1361,N_1320);
nand U3626 (N_3626,N_1333,N_2059);
or U3627 (N_3627,N_1963,N_1801);
nor U3628 (N_3628,N_1752,N_2121);
nand U3629 (N_3629,N_2098,N_1558);
or U3630 (N_3630,N_1348,N_1797);
or U3631 (N_3631,N_2466,N_1473);
nor U3632 (N_3632,N_1850,N_1754);
or U3633 (N_3633,N_2445,N_1323);
and U3634 (N_3634,N_1961,N_2020);
or U3635 (N_3635,N_1809,N_1834);
nand U3636 (N_3636,N_2299,N_2235);
nand U3637 (N_3637,N_1578,N_1966);
and U3638 (N_3638,N_1470,N_2409);
or U3639 (N_3639,N_2213,N_2335);
nand U3640 (N_3640,N_2289,N_2269);
nand U3641 (N_3641,N_1378,N_2025);
nand U3642 (N_3642,N_2339,N_1817);
xnor U3643 (N_3643,N_1342,N_2372);
and U3644 (N_3644,N_2442,N_1405);
or U3645 (N_3645,N_1940,N_2198);
nand U3646 (N_3646,N_1412,N_2318);
nor U3647 (N_3647,N_1995,N_1361);
xor U3648 (N_3648,N_2055,N_2016);
xnor U3649 (N_3649,N_2214,N_1736);
nand U3650 (N_3650,N_2160,N_1859);
nor U3651 (N_3651,N_1507,N_1907);
or U3652 (N_3652,N_2355,N_1764);
and U3653 (N_3653,N_1381,N_1483);
xor U3654 (N_3654,N_1802,N_1900);
or U3655 (N_3655,N_2234,N_2215);
and U3656 (N_3656,N_1422,N_1827);
and U3657 (N_3657,N_2474,N_1945);
and U3658 (N_3658,N_1322,N_1580);
or U3659 (N_3659,N_1910,N_2057);
nand U3660 (N_3660,N_1788,N_2414);
or U3661 (N_3661,N_1588,N_1545);
xnor U3662 (N_3662,N_2492,N_1685);
xnor U3663 (N_3663,N_1369,N_1823);
xnor U3664 (N_3664,N_2487,N_1764);
or U3665 (N_3665,N_1302,N_2453);
nor U3666 (N_3666,N_1513,N_1658);
or U3667 (N_3667,N_1619,N_2053);
nor U3668 (N_3668,N_1390,N_1324);
or U3669 (N_3669,N_2127,N_2156);
or U3670 (N_3670,N_2227,N_1312);
or U3671 (N_3671,N_1787,N_1943);
nand U3672 (N_3672,N_2190,N_1364);
nand U3673 (N_3673,N_2304,N_1659);
xnor U3674 (N_3674,N_2342,N_1324);
xnor U3675 (N_3675,N_1296,N_2453);
and U3676 (N_3676,N_1643,N_1511);
nand U3677 (N_3677,N_1333,N_1536);
nand U3678 (N_3678,N_2003,N_1721);
nand U3679 (N_3679,N_1391,N_1506);
and U3680 (N_3680,N_2420,N_1278);
xnor U3681 (N_3681,N_1666,N_2019);
nand U3682 (N_3682,N_1884,N_1637);
and U3683 (N_3683,N_1576,N_2289);
nand U3684 (N_3684,N_2264,N_2218);
and U3685 (N_3685,N_2311,N_1267);
nor U3686 (N_3686,N_1309,N_1360);
xnor U3687 (N_3687,N_1857,N_1346);
and U3688 (N_3688,N_1635,N_1843);
nand U3689 (N_3689,N_2303,N_2081);
nor U3690 (N_3690,N_1556,N_2028);
nor U3691 (N_3691,N_1829,N_2353);
nor U3692 (N_3692,N_1357,N_2397);
nand U3693 (N_3693,N_2195,N_2186);
or U3694 (N_3694,N_2332,N_2214);
or U3695 (N_3695,N_2497,N_1802);
or U3696 (N_3696,N_1593,N_2365);
nand U3697 (N_3697,N_1869,N_1775);
or U3698 (N_3698,N_1604,N_2302);
nor U3699 (N_3699,N_1443,N_2193);
and U3700 (N_3700,N_2111,N_1872);
xnor U3701 (N_3701,N_2041,N_2493);
or U3702 (N_3702,N_2297,N_2394);
and U3703 (N_3703,N_1880,N_1608);
nand U3704 (N_3704,N_2269,N_1468);
xnor U3705 (N_3705,N_2076,N_1697);
nor U3706 (N_3706,N_1331,N_1510);
xnor U3707 (N_3707,N_1289,N_2204);
nor U3708 (N_3708,N_1738,N_2000);
nor U3709 (N_3709,N_1877,N_1653);
xor U3710 (N_3710,N_1459,N_2420);
and U3711 (N_3711,N_1320,N_1604);
and U3712 (N_3712,N_1826,N_2057);
nand U3713 (N_3713,N_2300,N_1636);
and U3714 (N_3714,N_2241,N_1759);
xor U3715 (N_3715,N_2224,N_2265);
xor U3716 (N_3716,N_1618,N_1629);
nand U3717 (N_3717,N_1412,N_1634);
nand U3718 (N_3718,N_1755,N_2383);
xnor U3719 (N_3719,N_1902,N_1514);
nor U3720 (N_3720,N_1521,N_2000);
xor U3721 (N_3721,N_1790,N_1881);
or U3722 (N_3722,N_2077,N_1827);
nand U3723 (N_3723,N_2113,N_1776);
or U3724 (N_3724,N_1982,N_1541);
or U3725 (N_3725,N_2403,N_1625);
nand U3726 (N_3726,N_2422,N_2316);
xnor U3727 (N_3727,N_1967,N_2297);
nand U3728 (N_3728,N_2432,N_2087);
and U3729 (N_3729,N_1897,N_2053);
nand U3730 (N_3730,N_1311,N_2048);
nor U3731 (N_3731,N_1599,N_1294);
xor U3732 (N_3732,N_2329,N_1537);
xor U3733 (N_3733,N_1680,N_2263);
or U3734 (N_3734,N_1878,N_1730);
xnor U3735 (N_3735,N_2091,N_2050);
nand U3736 (N_3736,N_1484,N_1689);
nand U3737 (N_3737,N_1761,N_1381);
nor U3738 (N_3738,N_1927,N_1517);
xnor U3739 (N_3739,N_2033,N_2385);
and U3740 (N_3740,N_1773,N_2390);
and U3741 (N_3741,N_2449,N_1265);
nor U3742 (N_3742,N_2376,N_1941);
nor U3743 (N_3743,N_1332,N_1269);
nand U3744 (N_3744,N_1453,N_2175);
xor U3745 (N_3745,N_2375,N_2158);
nor U3746 (N_3746,N_2123,N_2164);
and U3747 (N_3747,N_2348,N_2147);
nand U3748 (N_3748,N_1306,N_2154);
or U3749 (N_3749,N_1440,N_2253);
xor U3750 (N_3750,N_3661,N_2709);
and U3751 (N_3751,N_3527,N_3403);
or U3752 (N_3752,N_3524,N_3178);
xnor U3753 (N_3753,N_2983,N_3351);
nand U3754 (N_3754,N_3481,N_2680);
or U3755 (N_3755,N_2631,N_3457);
or U3756 (N_3756,N_2538,N_2947);
nor U3757 (N_3757,N_3017,N_2771);
nor U3758 (N_3758,N_3005,N_3747);
and U3759 (N_3759,N_2896,N_2634);
and U3760 (N_3760,N_3504,N_3271);
or U3761 (N_3761,N_2853,N_3036);
xnor U3762 (N_3762,N_3620,N_2550);
xnor U3763 (N_3763,N_2872,N_2751);
nand U3764 (N_3764,N_2991,N_3255);
nand U3765 (N_3765,N_2944,N_2578);
and U3766 (N_3766,N_2980,N_2621);
nor U3767 (N_3767,N_2523,N_3023);
nor U3768 (N_3768,N_3229,N_3076);
xnor U3769 (N_3769,N_2607,N_2598);
nor U3770 (N_3770,N_2839,N_2881);
xnor U3771 (N_3771,N_3226,N_2987);
or U3772 (N_3772,N_2614,N_3369);
or U3773 (N_3773,N_2951,N_3198);
xnor U3774 (N_3774,N_2545,N_2911);
xnor U3775 (N_3775,N_2752,N_3409);
or U3776 (N_3776,N_3621,N_2804);
xnor U3777 (N_3777,N_3328,N_3103);
nor U3778 (N_3778,N_3040,N_3566);
nand U3779 (N_3779,N_3066,N_2518);
nand U3780 (N_3780,N_2921,N_2585);
nor U3781 (N_3781,N_3435,N_3533);
nor U3782 (N_3782,N_2852,N_3074);
nor U3783 (N_3783,N_3570,N_3393);
and U3784 (N_3784,N_3394,N_3249);
nand U3785 (N_3785,N_3565,N_3118);
and U3786 (N_3786,N_3731,N_3625);
or U3787 (N_3787,N_3618,N_3519);
nor U3788 (N_3788,N_3711,N_3647);
xor U3789 (N_3789,N_3237,N_2899);
or U3790 (N_3790,N_2889,N_2652);
or U3791 (N_3791,N_3173,N_3218);
nand U3792 (N_3792,N_2761,N_3186);
xnor U3793 (N_3793,N_2686,N_3551);
nand U3794 (N_3794,N_2711,N_2782);
xor U3795 (N_3795,N_3438,N_2836);
or U3796 (N_3796,N_3538,N_3289);
and U3797 (N_3797,N_3601,N_3706);
nor U3798 (N_3798,N_3308,N_3384);
xor U3799 (N_3799,N_3658,N_3248);
and U3800 (N_3800,N_3117,N_3631);
xnor U3801 (N_3801,N_3130,N_3689);
and U3802 (N_3802,N_3137,N_3267);
nand U3803 (N_3803,N_3395,N_2920);
nand U3804 (N_3804,N_2883,N_3217);
nand U3805 (N_3805,N_3743,N_2575);
nor U3806 (N_3806,N_2620,N_3145);
nand U3807 (N_3807,N_3682,N_2644);
xor U3808 (N_3808,N_2582,N_3083);
nand U3809 (N_3809,N_3167,N_2741);
and U3810 (N_3810,N_3113,N_3441);
or U3811 (N_3811,N_3468,N_3474);
nand U3812 (N_3812,N_2616,N_3192);
nor U3813 (N_3813,N_2970,N_3526);
or U3814 (N_3814,N_2641,N_3509);
nand U3815 (N_3815,N_3084,N_3303);
xnor U3816 (N_3816,N_3253,N_2733);
nand U3817 (N_3817,N_3588,N_2873);
nand U3818 (N_3818,N_3556,N_3344);
nand U3819 (N_3819,N_2957,N_3685);
and U3820 (N_3820,N_2848,N_3413);
or U3821 (N_3821,N_3710,N_3039);
or U3822 (N_3822,N_2871,N_3397);
or U3823 (N_3823,N_3189,N_3626);
xnor U3824 (N_3824,N_2508,N_3326);
nand U3825 (N_3825,N_3325,N_3247);
xnor U3826 (N_3826,N_3460,N_2603);
and U3827 (N_3827,N_3168,N_3242);
xnor U3828 (N_3828,N_2812,N_3211);
nor U3829 (N_3829,N_3494,N_3108);
nor U3830 (N_3830,N_3748,N_3321);
nand U3831 (N_3831,N_2758,N_2723);
and U3832 (N_3832,N_3518,N_3312);
nor U3833 (N_3833,N_3613,N_2588);
nand U3834 (N_3834,N_3085,N_2901);
or U3835 (N_3835,N_2590,N_3480);
and U3836 (N_3836,N_3560,N_2805);
xor U3837 (N_3837,N_2560,N_3387);
or U3838 (N_3838,N_2994,N_3490);
nor U3839 (N_3839,N_3204,N_2981);
and U3840 (N_3840,N_2956,N_3109);
nand U3841 (N_3841,N_3707,N_2638);
xor U3842 (N_3842,N_3745,N_3712);
nor U3843 (N_3843,N_3641,N_3236);
or U3844 (N_3844,N_2551,N_3425);
nand U3845 (N_3845,N_3071,N_3715);
or U3846 (N_3846,N_3699,N_3734);
or U3847 (N_3847,N_2689,N_2724);
or U3848 (N_3848,N_3529,N_2697);
or U3849 (N_3849,N_2504,N_3127);
or U3850 (N_3850,N_3170,N_2824);
nand U3851 (N_3851,N_3210,N_3119);
nand U3852 (N_3852,N_3452,N_2613);
and U3853 (N_3853,N_3503,N_2690);
nand U3854 (N_3854,N_2938,N_2636);
xor U3855 (N_3855,N_2831,N_2977);
xnor U3856 (N_3856,N_2735,N_3616);
and U3857 (N_3857,N_2754,N_2894);
xnor U3858 (N_3858,N_3042,N_3528);
or U3859 (N_3859,N_2778,N_2919);
nand U3860 (N_3860,N_2978,N_3680);
nand U3861 (N_3861,N_3738,N_2567);
or U3862 (N_3862,N_3391,N_3022);
nand U3863 (N_3863,N_3670,N_2584);
and U3864 (N_3864,N_3521,N_2583);
xnor U3865 (N_3865,N_2505,N_3287);
nor U3866 (N_3866,N_2639,N_2882);
nand U3867 (N_3867,N_2655,N_2840);
and U3868 (N_3868,N_3027,N_3431);
nor U3869 (N_3869,N_3506,N_3059);
and U3870 (N_3870,N_2602,N_3428);
and U3871 (N_3871,N_2605,N_3098);
and U3872 (N_3872,N_3619,N_3422);
and U3873 (N_3873,N_2997,N_3306);
or U3874 (N_3874,N_3335,N_2816);
xor U3875 (N_3875,N_3291,N_2838);
nor U3876 (N_3876,N_3692,N_3047);
or U3877 (N_3877,N_3583,N_3479);
nand U3878 (N_3878,N_3385,N_2945);
nand U3879 (N_3879,N_3199,N_2884);
xor U3880 (N_3880,N_2826,N_2813);
or U3881 (N_3881,N_3125,N_3446);
nor U3882 (N_3882,N_3116,N_2666);
and U3883 (N_3883,N_3106,N_3194);
nor U3884 (N_3884,N_2799,N_3544);
xnor U3885 (N_3885,N_2541,N_3193);
nand U3886 (N_3886,N_2592,N_2695);
nand U3887 (N_3887,N_3184,N_3592);
or U3888 (N_3888,N_3426,N_3639);
nor U3889 (N_3889,N_2513,N_3644);
or U3890 (N_3890,N_3231,N_3126);
xor U3891 (N_3891,N_3548,N_3095);
nand U3892 (N_3892,N_3594,N_3164);
or U3893 (N_3893,N_2609,N_3187);
xnor U3894 (N_3894,N_3695,N_3448);
or U3895 (N_3895,N_3300,N_3667);
nor U3896 (N_3896,N_3553,N_3128);
or U3897 (N_3897,N_3359,N_3094);
nand U3898 (N_3898,N_3493,N_3461);
nand U3899 (N_3899,N_3342,N_3096);
or U3900 (N_3900,N_2669,N_3634);
or U3901 (N_3901,N_3681,N_3181);
and U3902 (N_3902,N_2687,N_3102);
xor U3903 (N_3903,N_2738,N_3546);
xor U3904 (N_3904,N_2903,N_3587);
or U3905 (N_3905,N_2877,N_2516);
xnor U3906 (N_3906,N_3139,N_2861);
or U3907 (N_3907,N_3294,N_3251);
and U3908 (N_3908,N_3659,N_2912);
nand U3909 (N_3909,N_2581,N_3576);
xnor U3910 (N_3910,N_2880,N_2930);
xnor U3911 (N_3911,N_2918,N_3402);
nand U3912 (N_3912,N_2924,N_3572);
or U3913 (N_3913,N_2942,N_3179);
nor U3914 (N_3914,N_2793,N_3188);
xor U3915 (N_3915,N_2952,N_3323);
and U3916 (N_3916,N_3286,N_3174);
and U3917 (N_3917,N_2536,N_3324);
nor U3918 (N_3918,N_2643,N_3223);
and U3919 (N_3919,N_3606,N_3112);
nor U3920 (N_3920,N_3270,N_3221);
or U3921 (N_3921,N_3314,N_3258);
or U3922 (N_3922,N_3668,N_3605);
nor U3923 (N_3923,N_2657,N_2966);
or U3924 (N_3924,N_3020,N_3728);
and U3925 (N_3925,N_2719,N_3632);
and U3926 (N_3926,N_3408,N_3157);
and U3927 (N_3927,N_2969,N_3687);
and U3928 (N_3928,N_3197,N_3175);
and U3929 (N_3929,N_3702,N_3311);
nor U3930 (N_3930,N_2502,N_2961);
and U3931 (N_3931,N_2500,N_3586);
nand U3932 (N_3932,N_3567,N_2787);
nor U3933 (N_3933,N_3058,N_3648);
nor U3934 (N_3934,N_3531,N_2954);
and U3935 (N_3935,N_2628,N_2841);
or U3936 (N_3936,N_2715,N_3055);
and U3937 (N_3937,N_3052,N_2718);
nand U3938 (N_3938,N_2774,N_3115);
xor U3939 (N_3939,N_2801,N_2594);
or U3940 (N_3940,N_3001,N_3742);
nand U3941 (N_3941,N_3361,N_3357);
nor U3942 (N_3942,N_3337,N_3640);
nor U3943 (N_3943,N_3144,N_3230);
or U3944 (N_3944,N_3726,N_2955);
and U3945 (N_3945,N_2768,N_2985);
or U3946 (N_3946,N_3444,N_2731);
xor U3947 (N_3947,N_3464,N_3612);
or U3948 (N_3948,N_2726,N_2535);
nor U3949 (N_3949,N_2658,N_3675);
and U3950 (N_3950,N_2902,N_3525);
and U3951 (N_3951,N_3575,N_2928);
nor U3952 (N_3952,N_2950,N_3327);
and U3953 (N_3953,N_3716,N_3578);
and U3954 (N_3954,N_3346,N_2650);
xor U3955 (N_3955,N_3028,N_3688);
nor U3956 (N_3956,N_3362,N_2822);
and U3957 (N_3957,N_3590,N_3744);
and U3958 (N_3958,N_3741,N_3407);
and U3959 (N_3959,N_2790,N_2984);
xor U3960 (N_3960,N_3355,N_2637);
or U3961 (N_3961,N_2916,N_2737);
nor U3962 (N_3962,N_3298,N_3339);
nor U3963 (N_3963,N_3637,N_3260);
nand U3964 (N_3964,N_2597,N_3135);
xor U3965 (N_3965,N_3338,N_3649);
or U3966 (N_3966,N_3693,N_2716);
nor U3967 (N_3967,N_2781,N_3041);
or U3968 (N_3968,N_2962,N_2647);
and U3969 (N_3969,N_3523,N_2789);
and U3970 (N_3970,N_3165,N_3269);
nor U3971 (N_3971,N_3482,N_2815);
xor U3972 (N_3972,N_2850,N_2743);
nand U3973 (N_3973,N_3622,N_2688);
nand U3974 (N_3974,N_2832,N_3495);
or U3975 (N_3975,N_3153,N_3347);
and U3976 (N_3976,N_2553,N_2755);
xnor U3977 (N_3977,N_3740,N_3143);
nor U3978 (N_3978,N_2648,N_3305);
nor U3979 (N_3979,N_3598,N_3176);
xnor U3980 (N_3980,N_3088,N_2829);
nand U3981 (N_3981,N_3379,N_2979);
nand U3982 (N_3982,N_2777,N_3000);
nor U3983 (N_3983,N_2514,N_2512);
xnor U3984 (N_3984,N_2725,N_3498);
xnor U3985 (N_3985,N_3172,N_2624);
or U3986 (N_3986,N_3050,N_2593);
nor U3987 (N_3987,N_2606,N_3054);
nand U3988 (N_3988,N_3301,N_2915);
or U3989 (N_3989,N_3019,N_2557);
or U3990 (N_3990,N_2527,N_2975);
nand U3991 (N_3991,N_3320,N_2661);
xnor U3992 (N_3992,N_3439,N_3206);
or U3993 (N_3993,N_2646,N_2909);
and U3994 (N_3994,N_2530,N_3233);
xnor U3995 (N_3995,N_3180,N_2810);
xor U3996 (N_3996,N_3541,N_3016);
nor U3997 (N_3997,N_2507,N_2868);
and U3998 (N_3998,N_3063,N_3558);
xor U3999 (N_3999,N_3540,N_3595);
or U4000 (N_4000,N_3124,N_3638);
and U4001 (N_4001,N_3358,N_3150);
xor U4002 (N_4002,N_3122,N_3073);
xor U4003 (N_4003,N_3442,N_2904);
nor U4004 (N_4004,N_2651,N_3319);
xnor U4005 (N_4005,N_3486,N_3110);
xor U4006 (N_4006,N_3132,N_3013);
nand U4007 (N_4007,N_2803,N_2501);
and U4008 (N_4008,N_2948,N_3161);
nand U4009 (N_4009,N_3543,N_2722);
nand U4010 (N_4010,N_2933,N_3026);
and U4011 (N_4011,N_3352,N_3065);
xnor U4012 (N_4012,N_3010,N_2859);
and U4013 (N_4013,N_3256,N_3735);
or U4014 (N_4014,N_2668,N_2862);
nor U4015 (N_4015,N_3365,N_2760);
or U4016 (N_4016,N_3274,N_3536);
or U4017 (N_4017,N_2765,N_3239);
or U4018 (N_4018,N_3212,N_3507);
nand U4019 (N_4019,N_3263,N_3080);
xor U4020 (N_4020,N_2897,N_3183);
or U4021 (N_4021,N_3629,N_2586);
nand U4022 (N_4022,N_3310,N_3445);
xor U4023 (N_4023,N_3225,N_2905);
xnor U4024 (N_4024,N_3645,N_2802);
xnor U4025 (N_4025,N_3581,N_3471);
nor U4026 (N_4026,N_3709,N_3732);
nor U4027 (N_4027,N_3254,N_3404);
nand U4028 (N_4028,N_3003,N_2554);
xor U4029 (N_4029,N_2509,N_2696);
xor U4030 (N_4030,N_3101,N_3686);
nor U4031 (N_4031,N_3375,N_2958);
nand U4032 (N_4032,N_2833,N_3033);
or U4033 (N_4033,N_3141,N_2746);
nand U4034 (N_4034,N_2866,N_2684);
xor U4035 (N_4035,N_3160,N_3288);
nor U4036 (N_4036,N_2779,N_3257);
nand U4037 (N_4037,N_2845,N_3151);
or U4038 (N_4038,N_3304,N_3694);
nor U4039 (N_4039,N_3348,N_3148);
nand U4040 (N_4040,N_3008,N_3099);
and U4041 (N_4041,N_2764,N_3636);
nor U4042 (N_4042,N_2665,N_3049);
nor U4043 (N_4043,N_3500,N_2849);
xor U4044 (N_4044,N_3025,N_3714);
xnor U4045 (N_4045,N_3559,N_2574);
xor U4046 (N_4046,N_2934,N_3154);
and U4047 (N_4047,N_2807,N_3574);
or U4048 (N_4048,N_3579,N_2681);
nor U4049 (N_4049,N_3350,N_2797);
nand U4050 (N_4050,N_2775,N_3561);
xor U4051 (N_4051,N_3545,N_2670);
nor U4052 (N_4052,N_3573,N_2562);
nor U4053 (N_4053,N_3353,N_2784);
or U4054 (N_4054,N_2732,N_3070);
and U4055 (N_4055,N_2965,N_3004);
nor U4056 (N_4056,N_2710,N_3276);
nand U4057 (N_4057,N_2964,N_3203);
or U4058 (N_4058,N_3653,N_2855);
and U4059 (N_4059,N_3190,N_3302);
nor U4060 (N_4060,N_3380,N_3429);
xor U4061 (N_4061,N_2908,N_2534);
or U4062 (N_4062,N_2503,N_2580);
xor U4063 (N_4063,N_2885,N_3749);
nor U4064 (N_4064,N_3234,N_2608);
nor U4065 (N_4065,N_3664,N_2730);
nor U4066 (N_4066,N_3081,N_3259);
nor U4067 (N_4067,N_3163,N_3185);
and U4068 (N_4068,N_3666,N_3158);
nand U4069 (N_4069,N_3508,N_2863);
and U4070 (N_4070,N_3723,N_3371);
nor U4071 (N_4071,N_3502,N_3275);
xnor U4072 (N_4072,N_2568,N_3034);
nor U4073 (N_4073,N_3698,N_3496);
or U4074 (N_4074,N_3532,N_3162);
and U4075 (N_4075,N_3549,N_3313);
xnor U4076 (N_4076,N_3285,N_3295);
xor U4077 (N_4077,N_2703,N_2932);
nand U4078 (N_4078,N_3297,N_3440);
nand U4079 (N_4079,N_2993,N_3662);
or U4080 (N_4080,N_2679,N_3458);
nor U4081 (N_4081,N_2576,N_3031);
and U4082 (N_4082,N_3671,N_3673);
nor U4083 (N_4083,N_3089,N_2900);
nand U4084 (N_4084,N_3463,N_2796);
xor U4085 (N_4085,N_2806,N_2522);
nand U4086 (N_4086,N_3720,N_3552);
and U4087 (N_4087,N_2992,N_3038);
nand U4088 (N_4088,N_2618,N_2707);
nand U4089 (N_4089,N_2706,N_3411);
nand U4090 (N_4090,N_3195,N_2600);
and U4091 (N_4091,N_3398,N_2629);
nor U4092 (N_4092,N_3562,N_3542);
and U4093 (N_4093,N_3657,N_2895);
or U4094 (N_4094,N_2943,N_3227);
nor U4095 (N_4095,N_3554,N_3123);
or U4096 (N_4096,N_2867,N_3571);
xor U4097 (N_4097,N_3410,N_3418);
and U4098 (N_4098,N_3246,N_2677);
and U4099 (N_4099,N_2663,N_3512);
nand U4100 (N_4100,N_3278,N_2940);
nor U4101 (N_4101,N_3539,N_3420);
nand U4102 (N_4102,N_3608,N_2972);
and U4103 (N_4103,N_2525,N_3417);
or U4104 (N_4104,N_3356,N_2558);
and U4105 (N_4105,N_3060,N_3651);
or U4106 (N_4106,N_2556,N_3120);
xnor U4107 (N_4107,N_3390,N_2570);
nor U4108 (N_4108,N_2869,N_2898);
nor U4109 (N_4109,N_3679,N_3330);
and U4110 (N_4110,N_2999,N_2546);
nor U4111 (N_4111,N_2886,N_3736);
or U4112 (N_4112,N_2893,N_3208);
and U4113 (N_4113,N_2772,N_2704);
and U4114 (N_4114,N_3207,N_3633);
and U4115 (N_4115,N_3467,N_3196);
nor U4116 (N_4116,N_2596,N_3603);
and U4117 (N_4117,N_3273,N_3419);
and U4118 (N_4118,N_2623,N_3577);
nor U4119 (N_4119,N_3696,N_2595);
and U4120 (N_4120,N_3243,N_2907);
and U4121 (N_4121,N_3427,N_3635);
xnor U4122 (N_4122,N_3491,N_2653);
xnor U4123 (N_4123,N_2734,N_3349);
xor U4124 (N_4124,N_3456,N_2701);
and U4125 (N_4125,N_2892,N_2783);
nand U4126 (N_4126,N_2630,N_2820);
or U4127 (N_4127,N_2953,N_2524);
xor U4128 (N_4128,N_3465,N_2828);
and U4129 (N_4129,N_2720,N_3580);
xnor U4130 (N_4130,N_3284,N_3091);
xnor U4131 (N_4131,N_3149,N_2672);
nor U4132 (N_4132,N_3614,N_3092);
nor U4133 (N_4133,N_3470,N_3447);
or U4134 (N_4134,N_3615,N_3607);
nor U4135 (N_4135,N_3245,N_2808);
and U4136 (N_4136,N_3436,N_3600);
or U4137 (N_4137,N_3191,N_2537);
nor U4138 (N_4138,N_3006,N_2561);
or U4139 (N_4139,N_3730,N_2971);
nand U4140 (N_4140,N_3555,N_2742);
xor U4141 (N_4141,N_3568,N_2973);
xnor U4142 (N_4142,N_2963,N_3364);
or U4143 (N_4143,N_2740,N_3146);
or U4144 (N_4144,N_3376,N_2798);
and U4145 (N_4145,N_2599,N_3663);
nor U4146 (N_4146,N_2531,N_2721);
or U4147 (N_4147,N_2968,N_3655);
and U4148 (N_4148,N_2995,N_2520);
nor U4149 (N_4149,N_2996,N_2569);
or U4150 (N_4150,N_3389,N_2564);
nand U4151 (N_4151,N_2511,N_3046);
nand U4152 (N_4152,N_3282,N_2864);
or U4153 (N_4153,N_3104,N_3437);
or U4154 (N_4154,N_3497,N_2814);
xnor U4155 (N_4155,N_3534,N_2671);
and U4156 (N_4156,N_2788,N_3515);
xnor U4157 (N_4157,N_2601,N_2632);
xor U4158 (N_4158,N_3216,N_3318);
nor U4159 (N_4159,N_2976,N_2949);
and U4160 (N_4160,N_3235,N_3232);
xnor U4161 (N_4161,N_2865,N_3697);
nand U4162 (N_4162,N_2759,N_2766);
and U4163 (N_4163,N_2891,N_3416);
nand U4164 (N_4164,N_3377,N_2674);
or U4165 (N_4165,N_3138,N_3370);
nand U4166 (N_4166,N_3087,N_3704);
nand U4167 (N_4167,N_2929,N_2876);
nor U4168 (N_4168,N_3646,N_3093);
or U4169 (N_4169,N_3727,N_2573);
xnor U4170 (N_4170,N_2837,N_3433);
nand U4171 (N_4171,N_3037,N_3002);
nand U4172 (N_4172,N_3746,N_3228);
xor U4173 (N_4173,N_3374,N_3478);
nor U4174 (N_4174,N_3224,N_3265);
xor U4175 (N_4175,N_3596,N_3563);
and U4176 (N_4176,N_2611,N_2811);
or U4177 (N_4177,N_3341,N_3133);
and U4178 (N_4178,N_3719,N_3244);
and U4179 (N_4179,N_2517,N_3522);
xor U4180 (N_4180,N_2555,N_3281);
and U4181 (N_4181,N_3378,N_2913);
xnor U4182 (N_4182,N_2756,N_3501);
nor U4183 (N_4183,N_2773,N_3477);
or U4184 (N_4184,N_3056,N_3209);
xor U4185 (N_4185,N_3678,N_3064);
or U4186 (N_4186,N_3317,N_2540);
nand U4187 (N_4187,N_3530,N_3547);
xnor U4188 (N_4188,N_3643,N_3381);
or U4189 (N_4189,N_2809,N_2959);
and U4190 (N_4190,N_3068,N_3086);
nand U4191 (N_4191,N_2923,N_3261);
nand U4192 (N_4192,N_2619,N_3299);
nand U4193 (N_4193,N_3483,N_3617);
xnor U4194 (N_4194,N_2664,N_3372);
xor U4195 (N_4195,N_3061,N_3090);
nand U4196 (N_4196,N_2547,N_2794);
nand U4197 (N_4197,N_2510,N_2888);
and U4198 (N_4198,N_2800,N_2589);
xnor U4199 (N_4199,N_2542,N_2625);
nor U4200 (N_4200,N_2577,N_2579);
nand U4201 (N_4201,N_3107,N_3309);
nor U4202 (N_4202,N_2544,N_3032);
or U4203 (N_4203,N_2615,N_2700);
or U4204 (N_4204,N_2563,N_3513);
xnor U4205 (N_4205,N_2914,N_3564);
nor U4206 (N_4206,N_2656,N_3283);
or U4207 (N_4207,N_2649,N_3690);
nor U4208 (N_4208,N_3669,N_3343);
nor U4209 (N_4209,N_2572,N_2827);
or U4210 (N_4210,N_2559,N_3602);
nor U4211 (N_4211,N_2587,N_3296);
nor U4212 (N_4212,N_3652,N_2693);
nor U4213 (N_4213,N_3292,N_2926);
nand U4214 (N_4214,N_2591,N_3213);
and U4215 (N_4215,N_3492,N_2705);
xnor U4216 (N_4216,N_2515,N_2937);
nor U4217 (N_4217,N_2612,N_3654);
nand U4218 (N_4218,N_2708,N_3535);
nor U4219 (N_4219,N_2714,N_3051);
xor U4220 (N_4220,N_3166,N_3582);
nor U4221 (N_4221,N_2792,N_2526);
or U4222 (N_4222,N_3069,N_2757);
and U4223 (N_4223,N_2887,N_3363);
nor U4224 (N_4224,N_3100,N_3708);
or U4225 (N_4225,N_3067,N_2786);
or U4226 (N_4226,N_3214,N_2642);
nand U4227 (N_4227,N_3131,N_3450);
nand U4228 (N_4228,N_3114,N_3520);
and U4229 (N_4229,N_3434,N_3140);
nand U4230 (N_4230,N_2842,N_3367);
or U4231 (N_4231,N_3366,N_2830);
and U4232 (N_4232,N_3683,N_3424);
xnor U4233 (N_4233,N_3293,N_2890);
xor U4234 (N_4234,N_3705,N_2982);
and U4235 (N_4235,N_3737,N_3459);
xor U4236 (N_4236,N_3676,N_2694);
and U4237 (N_4237,N_2633,N_3266);
nand U4238 (N_4238,N_3268,N_3642);
xnor U4239 (N_4239,N_3584,N_3333);
nor U4240 (N_4240,N_3322,N_2640);
xor U4241 (N_4241,N_3215,N_2854);
and U4242 (N_4242,N_2662,N_3156);
nor U4243 (N_4243,N_3142,N_3057);
nand U4244 (N_4244,N_3200,N_3627);
nor U4245 (N_4245,N_3485,N_3475);
and U4246 (N_4246,N_3220,N_3550);
or U4247 (N_4247,N_2660,N_3511);
and U4248 (N_4248,N_3121,N_3340);
or U4249 (N_4249,N_2654,N_3078);
nand U4250 (N_4250,N_3048,N_2750);
xnor U4251 (N_4251,N_3171,N_3472);
nor U4252 (N_4252,N_3722,N_3399);
nor U4253 (N_4253,N_3514,N_3250);
xor U4254 (N_4254,N_3430,N_3725);
and U4255 (N_4255,N_2604,N_3077);
and U4256 (N_4256,N_3334,N_2879);
xor U4257 (N_4257,N_3386,N_2989);
or U4258 (N_4258,N_3272,N_3589);
xor U4259 (N_4259,N_2747,N_2533);
nand U4260 (N_4260,N_2673,N_2770);
and U4261 (N_4261,N_3159,N_3280);
xnor U4262 (N_4262,N_2795,N_2860);
nand U4263 (N_4263,N_2667,N_2565);
and U4264 (N_4264,N_3373,N_3354);
xor U4265 (N_4265,N_3012,N_3405);
xor U4266 (N_4266,N_3219,N_3015);
xnor U4267 (N_4267,N_2532,N_2878);
or U4268 (N_4268,N_3097,N_3691);
nand U4269 (N_4269,N_2762,N_3400);
and U4270 (N_4270,N_3018,N_2906);
nor U4271 (N_4271,N_3488,N_2847);
nand U4272 (N_4272,N_2834,N_2571);
xor U4273 (N_4273,N_3473,N_3316);
nand U4274 (N_4274,N_2974,N_3593);
and U4275 (N_4275,N_2931,N_2729);
or U4276 (N_4276,N_2925,N_2698);
or U4277 (N_4277,N_3451,N_2529);
nand U4278 (N_4278,N_2506,N_2817);
nor U4279 (N_4279,N_3277,N_2851);
or U4280 (N_4280,N_2936,N_2818);
nand U4281 (N_4281,N_2835,N_2960);
or U4282 (N_4282,N_3569,N_2702);
xnor U4283 (N_4283,N_3462,N_3201);
or U4284 (N_4284,N_2728,N_2988);
xor U4285 (N_4285,N_3599,N_3035);
xor U4286 (N_4286,N_3129,N_3043);
nor U4287 (N_4287,N_2659,N_2610);
nand U4288 (N_4288,N_3252,N_2691);
nand U4289 (N_4289,N_3388,N_2699);
or U4290 (N_4290,N_3406,N_3505);
xnor U4291 (N_4291,N_3336,N_3510);
xnor U4292 (N_4292,N_2986,N_3238);
xnor U4293 (N_4293,N_3489,N_3672);
or U4294 (N_4294,N_2519,N_3345);
xnor U4295 (N_4295,N_3007,N_2990);
nor U4296 (N_4296,N_2749,N_3677);
nand U4297 (N_4297,N_3072,N_2617);
nand U4298 (N_4298,N_3700,N_3262);
xnor U4299 (N_4299,N_3045,N_3591);
or U4300 (N_4300,N_3454,N_3703);
nand U4301 (N_4301,N_2675,N_2910);
nor U4302 (N_4302,N_3152,N_2736);
nor U4303 (N_4303,N_3656,N_2844);
nor U4304 (N_4304,N_2626,N_2870);
nor U4305 (N_4305,N_2552,N_2543);
and U4306 (N_4306,N_2857,N_2683);
nand U4307 (N_4307,N_3701,N_2712);
and U4308 (N_4308,N_2927,N_3182);
nor U4309 (N_4309,N_3610,N_2819);
xor U4310 (N_4310,N_2823,N_3733);
and U4311 (N_4311,N_2791,N_3401);
xnor U4312 (N_4312,N_2769,N_3134);
nor U4313 (N_4313,N_3155,N_3739);
xor U4314 (N_4314,N_2622,N_3516);
or U4315 (N_4315,N_2548,N_3222);
or U4316 (N_4316,N_3014,N_2846);
nor U4317 (N_4317,N_3674,N_2917);
nor U4318 (N_4318,N_3044,N_2767);
xor U4319 (N_4319,N_3383,N_2676);
nand U4320 (N_4320,N_3290,N_3368);
and U4321 (N_4321,N_3030,N_3021);
nor U4322 (N_4322,N_3053,N_3315);
xor U4323 (N_4323,N_3476,N_2776);
and U4324 (N_4324,N_3202,N_3630);
or U4325 (N_4325,N_3466,N_3029);
and U4326 (N_4326,N_3718,N_3136);
nor U4327 (N_4327,N_3412,N_3279);
or U4328 (N_4328,N_2946,N_3062);
or U4329 (N_4329,N_2566,N_3075);
nand U4330 (N_4330,N_3517,N_3147);
nor U4331 (N_4331,N_3724,N_3329);
and U4332 (N_4332,N_2875,N_3499);
xor U4333 (N_4333,N_3487,N_2967);
nand U4334 (N_4334,N_3011,N_3609);
nand U4335 (N_4335,N_3240,N_3332);
nand U4336 (N_4336,N_2825,N_2739);
or U4337 (N_4337,N_3585,N_3382);
or U4338 (N_4338,N_3423,N_2780);
xor U4339 (N_4339,N_3484,N_2785);
xnor U4340 (N_4340,N_2528,N_2821);
nand U4341 (N_4341,N_2748,N_3453);
nand U4342 (N_4342,N_2678,N_3611);
xnor U4343 (N_4343,N_2539,N_3264);
or U4344 (N_4344,N_3628,N_3241);
nor U4345 (N_4345,N_3169,N_3111);
or U4346 (N_4346,N_2935,N_2753);
nand U4347 (N_4347,N_2521,N_3331);
nand U4348 (N_4348,N_2763,N_3665);
and U4349 (N_4349,N_3449,N_2682);
and U4350 (N_4350,N_3469,N_3557);
or U4351 (N_4351,N_2635,N_3624);
nor U4352 (N_4352,N_2627,N_2645);
and U4353 (N_4353,N_3455,N_3537);
and U4354 (N_4354,N_3082,N_3713);
nor U4355 (N_4355,N_3307,N_3079);
xor U4356 (N_4356,N_3729,N_3604);
nor U4357 (N_4357,N_2858,N_2744);
nor U4358 (N_4358,N_2939,N_2922);
xor U4359 (N_4359,N_3443,N_2998);
nor U4360 (N_4360,N_2685,N_3024);
nor U4361 (N_4361,N_3432,N_3205);
nand U4362 (N_4362,N_2549,N_3392);
xnor U4363 (N_4363,N_2717,N_3360);
nor U4364 (N_4364,N_2856,N_2713);
and U4365 (N_4365,N_2745,N_3717);
or U4366 (N_4366,N_2843,N_3396);
and U4367 (N_4367,N_2941,N_3105);
or U4368 (N_4368,N_3421,N_3623);
xor U4369 (N_4369,N_2874,N_3684);
nor U4370 (N_4370,N_3660,N_2727);
nand U4371 (N_4371,N_3177,N_3415);
nor U4372 (N_4372,N_3650,N_3721);
nand U4373 (N_4373,N_3414,N_2692);
nand U4374 (N_4374,N_3597,N_3009);
or U4375 (N_4375,N_3239,N_3253);
xor U4376 (N_4376,N_2623,N_3243);
nor U4377 (N_4377,N_2503,N_2569);
xor U4378 (N_4378,N_3709,N_2541);
or U4379 (N_4379,N_3437,N_3250);
nand U4380 (N_4380,N_2753,N_3109);
nand U4381 (N_4381,N_2652,N_3564);
nor U4382 (N_4382,N_2929,N_3343);
or U4383 (N_4383,N_3537,N_3422);
xnor U4384 (N_4384,N_3314,N_3200);
nor U4385 (N_4385,N_2600,N_3022);
and U4386 (N_4386,N_3092,N_2738);
or U4387 (N_4387,N_3438,N_3521);
or U4388 (N_4388,N_2939,N_3355);
nor U4389 (N_4389,N_2699,N_3491);
or U4390 (N_4390,N_2858,N_2930);
nand U4391 (N_4391,N_3021,N_3392);
or U4392 (N_4392,N_2972,N_3361);
xnor U4393 (N_4393,N_3495,N_3368);
or U4394 (N_4394,N_2914,N_2899);
nor U4395 (N_4395,N_2758,N_2891);
nor U4396 (N_4396,N_3411,N_3554);
nor U4397 (N_4397,N_3662,N_3133);
nor U4398 (N_4398,N_2662,N_3744);
nand U4399 (N_4399,N_2895,N_3605);
or U4400 (N_4400,N_3554,N_2624);
and U4401 (N_4401,N_2988,N_2870);
or U4402 (N_4402,N_2746,N_2760);
or U4403 (N_4403,N_3311,N_2820);
nand U4404 (N_4404,N_2640,N_3109);
nor U4405 (N_4405,N_2845,N_3147);
or U4406 (N_4406,N_3612,N_3031);
or U4407 (N_4407,N_2810,N_3014);
nand U4408 (N_4408,N_3191,N_2901);
xor U4409 (N_4409,N_2919,N_2575);
xnor U4410 (N_4410,N_3586,N_3420);
nand U4411 (N_4411,N_2593,N_2933);
nand U4412 (N_4412,N_3590,N_2657);
nand U4413 (N_4413,N_3290,N_3512);
nand U4414 (N_4414,N_2605,N_3037);
xor U4415 (N_4415,N_2812,N_3528);
or U4416 (N_4416,N_2728,N_3702);
and U4417 (N_4417,N_3346,N_3515);
or U4418 (N_4418,N_2572,N_3130);
xor U4419 (N_4419,N_3533,N_2627);
or U4420 (N_4420,N_2876,N_2910);
or U4421 (N_4421,N_2604,N_2912);
xor U4422 (N_4422,N_3223,N_2782);
nand U4423 (N_4423,N_2543,N_3635);
and U4424 (N_4424,N_3041,N_2646);
nand U4425 (N_4425,N_3562,N_3749);
nand U4426 (N_4426,N_3106,N_2846);
nor U4427 (N_4427,N_2770,N_3136);
xnor U4428 (N_4428,N_2715,N_2585);
or U4429 (N_4429,N_3021,N_2969);
nand U4430 (N_4430,N_3157,N_3487);
xnor U4431 (N_4431,N_2598,N_3500);
nor U4432 (N_4432,N_3543,N_2520);
or U4433 (N_4433,N_3357,N_3035);
nand U4434 (N_4434,N_3087,N_2857);
or U4435 (N_4435,N_3082,N_3080);
nand U4436 (N_4436,N_2680,N_2655);
or U4437 (N_4437,N_2682,N_2823);
or U4438 (N_4438,N_3740,N_3318);
or U4439 (N_4439,N_3445,N_2902);
and U4440 (N_4440,N_3749,N_3683);
xor U4441 (N_4441,N_2989,N_2687);
nor U4442 (N_4442,N_3164,N_3314);
nor U4443 (N_4443,N_2581,N_2706);
nand U4444 (N_4444,N_3548,N_3283);
nor U4445 (N_4445,N_3590,N_3350);
xnor U4446 (N_4446,N_2857,N_2610);
nand U4447 (N_4447,N_3599,N_2834);
nand U4448 (N_4448,N_2591,N_3262);
nor U4449 (N_4449,N_3486,N_3403);
and U4450 (N_4450,N_3297,N_2823);
or U4451 (N_4451,N_3220,N_2528);
or U4452 (N_4452,N_2917,N_3380);
nand U4453 (N_4453,N_2896,N_3118);
or U4454 (N_4454,N_3202,N_2730);
or U4455 (N_4455,N_3152,N_3714);
xor U4456 (N_4456,N_3617,N_3426);
xnor U4457 (N_4457,N_3319,N_2898);
or U4458 (N_4458,N_3482,N_3547);
nor U4459 (N_4459,N_3265,N_2550);
nor U4460 (N_4460,N_2703,N_2785);
nand U4461 (N_4461,N_3139,N_2688);
or U4462 (N_4462,N_3676,N_3385);
or U4463 (N_4463,N_2872,N_3280);
nand U4464 (N_4464,N_2892,N_3288);
xor U4465 (N_4465,N_2923,N_3594);
nor U4466 (N_4466,N_2610,N_2920);
nand U4467 (N_4467,N_3264,N_3357);
and U4468 (N_4468,N_3038,N_3343);
xor U4469 (N_4469,N_3733,N_3168);
or U4470 (N_4470,N_3414,N_3052);
and U4471 (N_4471,N_3569,N_2850);
or U4472 (N_4472,N_2941,N_2756);
xor U4473 (N_4473,N_3569,N_2979);
nand U4474 (N_4474,N_3576,N_3298);
xor U4475 (N_4475,N_2643,N_3348);
xnor U4476 (N_4476,N_3455,N_3674);
xor U4477 (N_4477,N_2789,N_2779);
nor U4478 (N_4478,N_3349,N_2691);
or U4479 (N_4479,N_2607,N_2840);
and U4480 (N_4480,N_3129,N_3337);
or U4481 (N_4481,N_3202,N_2527);
nor U4482 (N_4482,N_2615,N_3263);
and U4483 (N_4483,N_2709,N_3012);
or U4484 (N_4484,N_2951,N_3064);
and U4485 (N_4485,N_3285,N_3521);
and U4486 (N_4486,N_3636,N_2957);
and U4487 (N_4487,N_3577,N_2894);
and U4488 (N_4488,N_2540,N_2547);
xor U4489 (N_4489,N_2523,N_2741);
nand U4490 (N_4490,N_3561,N_3305);
or U4491 (N_4491,N_3113,N_3318);
xnor U4492 (N_4492,N_3702,N_3365);
or U4493 (N_4493,N_2803,N_3105);
and U4494 (N_4494,N_2508,N_3019);
and U4495 (N_4495,N_2763,N_3141);
nand U4496 (N_4496,N_2813,N_3687);
nor U4497 (N_4497,N_3559,N_2727);
nor U4498 (N_4498,N_2698,N_3387);
nand U4499 (N_4499,N_3280,N_2907);
and U4500 (N_4500,N_2824,N_3054);
nor U4501 (N_4501,N_3385,N_3606);
and U4502 (N_4502,N_2795,N_2759);
or U4503 (N_4503,N_2604,N_2774);
nor U4504 (N_4504,N_2815,N_2666);
and U4505 (N_4505,N_3322,N_2839);
or U4506 (N_4506,N_2608,N_3122);
nand U4507 (N_4507,N_3732,N_2781);
nor U4508 (N_4508,N_3127,N_2772);
or U4509 (N_4509,N_2998,N_2579);
nand U4510 (N_4510,N_3396,N_2795);
nand U4511 (N_4511,N_3316,N_3354);
or U4512 (N_4512,N_2564,N_3104);
xnor U4513 (N_4513,N_2628,N_3423);
nand U4514 (N_4514,N_3385,N_3128);
xnor U4515 (N_4515,N_2673,N_2536);
and U4516 (N_4516,N_2701,N_3141);
nand U4517 (N_4517,N_3547,N_3107);
or U4518 (N_4518,N_3024,N_2603);
and U4519 (N_4519,N_3154,N_2615);
xor U4520 (N_4520,N_2663,N_3658);
nand U4521 (N_4521,N_2852,N_3255);
nor U4522 (N_4522,N_2908,N_3083);
or U4523 (N_4523,N_2627,N_2621);
or U4524 (N_4524,N_3354,N_2547);
or U4525 (N_4525,N_3651,N_2776);
nand U4526 (N_4526,N_3223,N_3125);
nand U4527 (N_4527,N_2844,N_2726);
xnor U4528 (N_4528,N_3141,N_3182);
and U4529 (N_4529,N_2925,N_2950);
or U4530 (N_4530,N_3322,N_2921);
or U4531 (N_4531,N_3456,N_2633);
nor U4532 (N_4532,N_2748,N_3143);
nor U4533 (N_4533,N_3313,N_2581);
xnor U4534 (N_4534,N_3428,N_3476);
xor U4535 (N_4535,N_3023,N_3093);
xor U4536 (N_4536,N_2831,N_2943);
nand U4537 (N_4537,N_3738,N_2571);
nor U4538 (N_4538,N_3620,N_3541);
or U4539 (N_4539,N_2550,N_3384);
xnor U4540 (N_4540,N_2686,N_2515);
xor U4541 (N_4541,N_3425,N_3562);
and U4542 (N_4542,N_3321,N_3143);
nor U4543 (N_4543,N_3253,N_2763);
nand U4544 (N_4544,N_3158,N_2807);
nor U4545 (N_4545,N_3354,N_2983);
and U4546 (N_4546,N_3257,N_3172);
nand U4547 (N_4547,N_2671,N_3571);
nand U4548 (N_4548,N_2895,N_3639);
or U4549 (N_4549,N_3735,N_2990);
xnor U4550 (N_4550,N_2639,N_2555);
xor U4551 (N_4551,N_2728,N_3687);
or U4552 (N_4552,N_3271,N_3683);
nand U4553 (N_4553,N_3604,N_2694);
nand U4554 (N_4554,N_3349,N_3230);
nor U4555 (N_4555,N_3667,N_2757);
nor U4556 (N_4556,N_3544,N_3489);
xnor U4557 (N_4557,N_3292,N_3326);
nand U4558 (N_4558,N_2541,N_3046);
or U4559 (N_4559,N_2872,N_3655);
xor U4560 (N_4560,N_2998,N_2839);
and U4561 (N_4561,N_2653,N_3636);
or U4562 (N_4562,N_3455,N_3516);
or U4563 (N_4563,N_2917,N_3122);
nor U4564 (N_4564,N_3040,N_3299);
and U4565 (N_4565,N_3130,N_3575);
or U4566 (N_4566,N_2882,N_2993);
nand U4567 (N_4567,N_2886,N_2503);
nand U4568 (N_4568,N_3008,N_3267);
and U4569 (N_4569,N_2935,N_2930);
or U4570 (N_4570,N_3025,N_3268);
nor U4571 (N_4571,N_2547,N_2837);
xor U4572 (N_4572,N_3258,N_3637);
xor U4573 (N_4573,N_2673,N_3737);
xnor U4574 (N_4574,N_2864,N_3232);
xor U4575 (N_4575,N_3290,N_3385);
and U4576 (N_4576,N_3078,N_3460);
xor U4577 (N_4577,N_3024,N_2650);
nand U4578 (N_4578,N_3663,N_3449);
nand U4579 (N_4579,N_3661,N_2939);
nor U4580 (N_4580,N_2694,N_2730);
and U4581 (N_4581,N_2952,N_2751);
nor U4582 (N_4582,N_3585,N_3642);
and U4583 (N_4583,N_3274,N_3719);
xor U4584 (N_4584,N_3462,N_2861);
and U4585 (N_4585,N_2738,N_2838);
nand U4586 (N_4586,N_2878,N_3725);
nor U4587 (N_4587,N_2658,N_3609);
nand U4588 (N_4588,N_3459,N_3149);
nor U4589 (N_4589,N_3117,N_3717);
nor U4590 (N_4590,N_2748,N_2566);
and U4591 (N_4591,N_3280,N_3127);
and U4592 (N_4592,N_2568,N_3088);
and U4593 (N_4593,N_2585,N_3340);
or U4594 (N_4594,N_2975,N_3651);
nor U4595 (N_4595,N_3679,N_2523);
nand U4596 (N_4596,N_2590,N_3273);
nand U4597 (N_4597,N_2833,N_2503);
or U4598 (N_4598,N_2647,N_2932);
and U4599 (N_4599,N_2523,N_3576);
or U4600 (N_4600,N_3186,N_3500);
nor U4601 (N_4601,N_3291,N_2645);
nor U4602 (N_4602,N_2547,N_2887);
nor U4603 (N_4603,N_3364,N_3579);
nor U4604 (N_4604,N_3659,N_2978);
or U4605 (N_4605,N_3620,N_3176);
xnor U4606 (N_4606,N_2638,N_3105);
and U4607 (N_4607,N_2947,N_3652);
nand U4608 (N_4608,N_2871,N_3040);
or U4609 (N_4609,N_3465,N_3432);
xor U4610 (N_4610,N_2878,N_2990);
xor U4611 (N_4611,N_3588,N_3660);
and U4612 (N_4612,N_3502,N_2902);
xnor U4613 (N_4613,N_3113,N_2914);
xor U4614 (N_4614,N_3717,N_3426);
nor U4615 (N_4615,N_3188,N_3714);
nand U4616 (N_4616,N_3149,N_2845);
or U4617 (N_4617,N_3659,N_2980);
nand U4618 (N_4618,N_3030,N_3564);
and U4619 (N_4619,N_3027,N_3149);
or U4620 (N_4620,N_3451,N_3483);
xor U4621 (N_4621,N_2982,N_3457);
or U4622 (N_4622,N_3552,N_2561);
nor U4623 (N_4623,N_3035,N_3602);
nor U4624 (N_4624,N_3258,N_3165);
nor U4625 (N_4625,N_3269,N_3604);
xnor U4626 (N_4626,N_3638,N_3103);
xor U4627 (N_4627,N_3413,N_3484);
or U4628 (N_4628,N_3313,N_3447);
nor U4629 (N_4629,N_3700,N_3337);
and U4630 (N_4630,N_2685,N_2766);
or U4631 (N_4631,N_2723,N_3526);
nor U4632 (N_4632,N_3411,N_2831);
or U4633 (N_4633,N_2671,N_3704);
nand U4634 (N_4634,N_3195,N_3521);
nand U4635 (N_4635,N_2888,N_2968);
nand U4636 (N_4636,N_3676,N_2715);
or U4637 (N_4637,N_2986,N_2790);
xnor U4638 (N_4638,N_3407,N_3500);
and U4639 (N_4639,N_3180,N_3717);
nor U4640 (N_4640,N_3220,N_3187);
nor U4641 (N_4641,N_3106,N_3219);
nor U4642 (N_4642,N_3331,N_2807);
nand U4643 (N_4643,N_3286,N_2673);
nor U4644 (N_4644,N_3197,N_2897);
nand U4645 (N_4645,N_3543,N_3734);
nand U4646 (N_4646,N_3177,N_3473);
xnor U4647 (N_4647,N_3357,N_2880);
and U4648 (N_4648,N_2869,N_2997);
and U4649 (N_4649,N_3501,N_3527);
xor U4650 (N_4650,N_3235,N_3219);
or U4651 (N_4651,N_2820,N_3289);
xnor U4652 (N_4652,N_3255,N_3222);
nand U4653 (N_4653,N_3695,N_3540);
xnor U4654 (N_4654,N_3299,N_3276);
xor U4655 (N_4655,N_2806,N_3318);
nand U4656 (N_4656,N_2522,N_3743);
nor U4657 (N_4657,N_3706,N_3313);
and U4658 (N_4658,N_3175,N_2776);
and U4659 (N_4659,N_2620,N_3529);
xor U4660 (N_4660,N_2897,N_2797);
nor U4661 (N_4661,N_3611,N_3016);
xor U4662 (N_4662,N_2514,N_3402);
nand U4663 (N_4663,N_2627,N_3598);
xor U4664 (N_4664,N_3006,N_3738);
or U4665 (N_4665,N_3458,N_3195);
and U4666 (N_4666,N_3297,N_3161);
and U4667 (N_4667,N_3635,N_3306);
xnor U4668 (N_4668,N_2890,N_3254);
nand U4669 (N_4669,N_3464,N_3385);
xnor U4670 (N_4670,N_2603,N_2719);
and U4671 (N_4671,N_3432,N_3643);
nor U4672 (N_4672,N_2783,N_2711);
nor U4673 (N_4673,N_2932,N_2993);
nor U4674 (N_4674,N_3589,N_2823);
or U4675 (N_4675,N_3055,N_3640);
or U4676 (N_4676,N_2865,N_3278);
nor U4677 (N_4677,N_2986,N_3168);
and U4678 (N_4678,N_3726,N_2763);
or U4679 (N_4679,N_2876,N_3491);
and U4680 (N_4680,N_3159,N_2982);
nand U4681 (N_4681,N_3742,N_3127);
nand U4682 (N_4682,N_3237,N_3537);
or U4683 (N_4683,N_3385,N_3312);
or U4684 (N_4684,N_2972,N_3551);
xor U4685 (N_4685,N_2871,N_3329);
nand U4686 (N_4686,N_3484,N_3702);
and U4687 (N_4687,N_3741,N_3133);
xnor U4688 (N_4688,N_3545,N_3571);
nor U4689 (N_4689,N_3540,N_2669);
or U4690 (N_4690,N_2798,N_3158);
nor U4691 (N_4691,N_2602,N_2714);
or U4692 (N_4692,N_3122,N_3333);
xor U4693 (N_4693,N_3120,N_2763);
or U4694 (N_4694,N_3172,N_3082);
xor U4695 (N_4695,N_3068,N_3151);
xor U4696 (N_4696,N_2780,N_3136);
nand U4697 (N_4697,N_3355,N_3443);
and U4698 (N_4698,N_3241,N_2605);
nor U4699 (N_4699,N_3470,N_3676);
nor U4700 (N_4700,N_2973,N_2507);
and U4701 (N_4701,N_3676,N_3002);
or U4702 (N_4702,N_2837,N_2555);
or U4703 (N_4703,N_3147,N_3146);
and U4704 (N_4704,N_3081,N_3108);
or U4705 (N_4705,N_3462,N_2590);
nand U4706 (N_4706,N_3662,N_3329);
or U4707 (N_4707,N_2534,N_2847);
xor U4708 (N_4708,N_3063,N_3102);
xnor U4709 (N_4709,N_3097,N_2542);
xor U4710 (N_4710,N_3583,N_3051);
nand U4711 (N_4711,N_3150,N_2963);
xor U4712 (N_4712,N_3656,N_3621);
nand U4713 (N_4713,N_3257,N_2676);
nand U4714 (N_4714,N_3397,N_2835);
and U4715 (N_4715,N_2805,N_2856);
nor U4716 (N_4716,N_3188,N_2837);
or U4717 (N_4717,N_3307,N_3356);
nor U4718 (N_4718,N_3425,N_2529);
nor U4719 (N_4719,N_2793,N_3667);
or U4720 (N_4720,N_3409,N_3391);
nand U4721 (N_4721,N_3027,N_3698);
or U4722 (N_4722,N_2940,N_3399);
nor U4723 (N_4723,N_3511,N_3252);
nor U4724 (N_4724,N_2761,N_2911);
and U4725 (N_4725,N_3099,N_3186);
nor U4726 (N_4726,N_2856,N_3506);
and U4727 (N_4727,N_3638,N_2614);
or U4728 (N_4728,N_2555,N_3068);
nand U4729 (N_4729,N_3275,N_2680);
or U4730 (N_4730,N_3604,N_3741);
xnor U4731 (N_4731,N_2837,N_3649);
nor U4732 (N_4732,N_2602,N_3456);
and U4733 (N_4733,N_2660,N_3425);
xor U4734 (N_4734,N_3193,N_2771);
xor U4735 (N_4735,N_2801,N_3572);
nand U4736 (N_4736,N_3123,N_2733);
nand U4737 (N_4737,N_3348,N_2843);
nand U4738 (N_4738,N_2719,N_2818);
or U4739 (N_4739,N_2696,N_3135);
xor U4740 (N_4740,N_3710,N_3324);
nor U4741 (N_4741,N_2989,N_2500);
and U4742 (N_4742,N_2601,N_3008);
and U4743 (N_4743,N_2525,N_3416);
nand U4744 (N_4744,N_3408,N_3185);
or U4745 (N_4745,N_3024,N_3406);
nand U4746 (N_4746,N_3436,N_2865);
xnor U4747 (N_4747,N_2809,N_3047);
nand U4748 (N_4748,N_2618,N_3323);
or U4749 (N_4749,N_3012,N_2912);
nand U4750 (N_4750,N_3619,N_2736);
nand U4751 (N_4751,N_3614,N_2516);
nand U4752 (N_4752,N_3389,N_2865);
nor U4753 (N_4753,N_2848,N_3318);
xnor U4754 (N_4754,N_2746,N_3410);
or U4755 (N_4755,N_3520,N_2538);
and U4756 (N_4756,N_2784,N_3549);
or U4757 (N_4757,N_2571,N_3332);
xor U4758 (N_4758,N_3673,N_3613);
nand U4759 (N_4759,N_3241,N_3123);
or U4760 (N_4760,N_3455,N_3195);
and U4761 (N_4761,N_2625,N_3016);
or U4762 (N_4762,N_3049,N_2894);
or U4763 (N_4763,N_3695,N_2528);
nor U4764 (N_4764,N_3713,N_2935);
xor U4765 (N_4765,N_3677,N_2887);
nor U4766 (N_4766,N_2576,N_3436);
or U4767 (N_4767,N_3526,N_3353);
nor U4768 (N_4768,N_3076,N_2514);
or U4769 (N_4769,N_3116,N_3517);
or U4770 (N_4770,N_3614,N_2965);
nand U4771 (N_4771,N_3531,N_3652);
nor U4772 (N_4772,N_3087,N_3268);
xor U4773 (N_4773,N_3234,N_2766);
xor U4774 (N_4774,N_2839,N_3718);
xor U4775 (N_4775,N_3072,N_3521);
xor U4776 (N_4776,N_3119,N_3570);
nand U4777 (N_4777,N_3230,N_3189);
and U4778 (N_4778,N_3596,N_2715);
and U4779 (N_4779,N_2906,N_3198);
nor U4780 (N_4780,N_3420,N_3471);
and U4781 (N_4781,N_3690,N_2590);
and U4782 (N_4782,N_3466,N_2716);
xnor U4783 (N_4783,N_3132,N_3452);
nor U4784 (N_4784,N_3026,N_3098);
and U4785 (N_4785,N_3724,N_3288);
nand U4786 (N_4786,N_3746,N_3486);
nand U4787 (N_4787,N_3493,N_2960);
or U4788 (N_4788,N_2560,N_2588);
or U4789 (N_4789,N_3502,N_3033);
or U4790 (N_4790,N_2527,N_3217);
and U4791 (N_4791,N_2944,N_2507);
nand U4792 (N_4792,N_3177,N_3574);
nor U4793 (N_4793,N_3722,N_2542);
and U4794 (N_4794,N_2748,N_2755);
nand U4795 (N_4795,N_3635,N_3545);
nand U4796 (N_4796,N_3267,N_3236);
nor U4797 (N_4797,N_3245,N_2814);
and U4798 (N_4798,N_2526,N_2756);
xnor U4799 (N_4799,N_3596,N_3592);
xor U4800 (N_4800,N_3659,N_3186);
nor U4801 (N_4801,N_3558,N_2677);
or U4802 (N_4802,N_3698,N_3113);
and U4803 (N_4803,N_2922,N_2759);
and U4804 (N_4804,N_3242,N_3093);
nand U4805 (N_4805,N_3241,N_2750);
or U4806 (N_4806,N_3126,N_3190);
and U4807 (N_4807,N_3104,N_3652);
nand U4808 (N_4808,N_2689,N_3411);
and U4809 (N_4809,N_3152,N_2663);
and U4810 (N_4810,N_3650,N_3131);
xnor U4811 (N_4811,N_3321,N_2997);
xnor U4812 (N_4812,N_3567,N_3307);
and U4813 (N_4813,N_3717,N_3490);
nand U4814 (N_4814,N_3558,N_3352);
or U4815 (N_4815,N_2887,N_2728);
xor U4816 (N_4816,N_2791,N_3275);
and U4817 (N_4817,N_3157,N_3090);
nand U4818 (N_4818,N_3593,N_3650);
xor U4819 (N_4819,N_2580,N_3720);
xor U4820 (N_4820,N_2656,N_2788);
and U4821 (N_4821,N_2572,N_3539);
or U4822 (N_4822,N_3160,N_3061);
and U4823 (N_4823,N_3023,N_2659);
and U4824 (N_4824,N_3430,N_3613);
nor U4825 (N_4825,N_2951,N_2542);
or U4826 (N_4826,N_2893,N_2904);
nand U4827 (N_4827,N_2580,N_3732);
xnor U4828 (N_4828,N_3254,N_2945);
and U4829 (N_4829,N_2779,N_2513);
xor U4830 (N_4830,N_3488,N_3724);
or U4831 (N_4831,N_2577,N_3310);
or U4832 (N_4832,N_3407,N_2973);
and U4833 (N_4833,N_3369,N_3156);
xor U4834 (N_4834,N_3016,N_3496);
xor U4835 (N_4835,N_2633,N_2948);
or U4836 (N_4836,N_3715,N_2526);
or U4837 (N_4837,N_2655,N_2820);
nor U4838 (N_4838,N_3727,N_3154);
and U4839 (N_4839,N_3155,N_3215);
nand U4840 (N_4840,N_2617,N_2673);
nand U4841 (N_4841,N_3418,N_3555);
nor U4842 (N_4842,N_3473,N_3675);
nor U4843 (N_4843,N_2815,N_3716);
nand U4844 (N_4844,N_2687,N_3067);
and U4845 (N_4845,N_3134,N_3048);
nand U4846 (N_4846,N_2527,N_3634);
and U4847 (N_4847,N_3025,N_3545);
nor U4848 (N_4848,N_2563,N_3710);
and U4849 (N_4849,N_3426,N_3723);
xor U4850 (N_4850,N_2736,N_2815);
xnor U4851 (N_4851,N_3720,N_2912);
nor U4852 (N_4852,N_2683,N_3459);
nand U4853 (N_4853,N_3634,N_3296);
nor U4854 (N_4854,N_2841,N_2943);
xnor U4855 (N_4855,N_3299,N_3332);
and U4856 (N_4856,N_2635,N_3377);
or U4857 (N_4857,N_3471,N_3500);
and U4858 (N_4858,N_3650,N_2569);
nor U4859 (N_4859,N_3334,N_3615);
and U4860 (N_4860,N_3184,N_2578);
and U4861 (N_4861,N_3174,N_2622);
xor U4862 (N_4862,N_2930,N_2953);
nand U4863 (N_4863,N_3175,N_2606);
xnor U4864 (N_4864,N_2597,N_3328);
nor U4865 (N_4865,N_3627,N_2782);
nor U4866 (N_4866,N_3308,N_2953);
nand U4867 (N_4867,N_3311,N_2953);
and U4868 (N_4868,N_3006,N_3704);
or U4869 (N_4869,N_3063,N_3484);
and U4870 (N_4870,N_2754,N_3611);
nor U4871 (N_4871,N_3378,N_3696);
and U4872 (N_4872,N_2849,N_2697);
or U4873 (N_4873,N_3370,N_2662);
or U4874 (N_4874,N_3690,N_3379);
xor U4875 (N_4875,N_3462,N_3697);
nor U4876 (N_4876,N_3257,N_3161);
and U4877 (N_4877,N_3370,N_2959);
nor U4878 (N_4878,N_2983,N_2755);
and U4879 (N_4879,N_3574,N_3065);
or U4880 (N_4880,N_2605,N_3393);
or U4881 (N_4881,N_2608,N_2882);
nor U4882 (N_4882,N_2930,N_3235);
xor U4883 (N_4883,N_3392,N_3617);
and U4884 (N_4884,N_2596,N_3393);
xnor U4885 (N_4885,N_3424,N_2837);
and U4886 (N_4886,N_3281,N_2899);
nand U4887 (N_4887,N_3140,N_2740);
or U4888 (N_4888,N_3435,N_3044);
nor U4889 (N_4889,N_2719,N_3682);
or U4890 (N_4890,N_3671,N_3257);
xnor U4891 (N_4891,N_3180,N_3068);
nor U4892 (N_4892,N_3172,N_2977);
nor U4893 (N_4893,N_2517,N_3554);
or U4894 (N_4894,N_2866,N_2966);
or U4895 (N_4895,N_3483,N_3560);
and U4896 (N_4896,N_3433,N_3424);
and U4897 (N_4897,N_2850,N_3561);
nor U4898 (N_4898,N_3547,N_3253);
and U4899 (N_4899,N_2984,N_3512);
or U4900 (N_4900,N_2850,N_3455);
nand U4901 (N_4901,N_3491,N_3513);
xor U4902 (N_4902,N_3142,N_3116);
xnor U4903 (N_4903,N_2918,N_3641);
or U4904 (N_4904,N_3632,N_3443);
nand U4905 (N_4905,N_3749,N_2856);
nor U4906 (N_4906,N_3060,N_3551);
xor U4907 (N_4907,N_3680,N_3354);
nor U4908 (N_4908,N_3315,N_2896);
xor U4909 (N_4909,N_3103,N_3483);
and U4910 (N_4910,N_3192,N_2718);
and U4911 (N_4911,N_2934,N_3027);
or U4912 (N_4912,N_2945,N_3411);
and U4913 (N_4913,N_3193,N_2647);
and U4914 (N_4914,N_3552,N_3585);
nor U4915 (N_4915,N_2797,N_3632);
nand U4916 (N_4916,N_2631,N_3153);
xor U4917 (N_4917,N_3055,N_3402);
nor U4918 (N_4918,N_3431,N_3631);
and U4919 (N_4919,N_2985,N_2645);
and U4920 (N_4920,N_3556,N_3189);
nor U4921 (N_4921,N_2722,N_2575);
or U4922 (N_4922,N_2863,N_3390);
or U4923 (N_4923,N_2843,N_2799);
nand U4924 (N_4924,N_3344,N_3525);
nand U4925 (N_4925,N_3312,N_2537);
nor U4926 (N_4926,N_3502,N_3189);
or U4927 (N_4927,N_3023,N_2838);
and U4928 (N_4928,N_3476,N_2749);
xnor U4929 (N_4929,N_2859,N_3622);
or U4930 (N_4930,N_3329,N_3139);
nand U4931 (N_4931,N_3114,N_3477);
and U4932 (N_4932,N_2838,N_2936);
xor U4933 (N_4933,N_3151,N_2528);
or U4934 (N_4934,N_3568,N_3217);
xnor U4935 (N_4935,N_2703,N_3146);
nand U4936 (N_4936,N_3272,N_2548);
nand U4937 (N_4937,N_2562,N_3365);
or U4938 (N_4938,N_3251,N_3190);
nor U4939 (N_4939,N_3564,N_3436);
nor U4940 (N_4940,N_3489,N_3029);
or U4941 (N_4941,N_3066,N_2792);
nand U4942 (N_4942,N_2805,N_2949);
xor U4943 (N_4943,N_3280,N_3701);
and U4944 (N_4944,N_3220,N_2915);
and U4945 (N_4945,N_3073,N_3714);
or U4946 (N_4946,N_3167,N_3465);
nand U4947 (N_4947,N_3576,N_3488);
nor U4948 (N_4948,N_2719,N_3175);
xnor U4949 (N_4949,N_2980,N_3247);
xor U4950 (N_4950,N_3285,N_3704);
or U4951 (N_4951,N_3157,N_3511);
nand U4952 (N_4952,N_3617,N_3257);
xnor U4953 (N_4953,N_2832,N_2988);
nor U4954 (N_4954,N_2666,N_3104);
and U4955 (N_4955,N_2860,N_2907);
and U4956 (N_4956,N_3682,N_2579);
and U4957 (N_4957,N_2653,N_2761);
nand U4958 (N_4958,N_2899,N_2812);
nand U4959 (N_4959,N_3097,N_3448);
xor U4960 (N_4960,N_3090,N_2988);
and U4961 (N_4961,N_2855,N_2766);
nor U4962 (N_4962,N_2668,N_2907);
nor U4963 (N_4963,N_3032,N_3260);
nand U4964 (N_4964,N_3194,N_2883);
or U4965 (N_4965,N_2586,N_3515);
xnor U4966 (N_4966,N_3309,N_2615);
nand U4967 (N_4967,N_2906,N_3119);
nand U4968 (N_4968,N_2916,N_3231);
nor U4969 (N_4969,N_3235,N_2570);
and U4970 (N_4970,N_3247,N_2738);
nor U4971 (N_4971,N_2853,N_3745);
and U4972 (N_4972,N_2948,N_3630);
nor U4973 (N_4973,N_2925,N_3376);
nand U4974 (N_4974,N_2550,N_3530);
nand U4975 (N_4975,N_3634,N_2898);
xor U4976 (N_4976,N_3499,N_2853);
nor U4977 (N_4977,N_2526,N_2825);
nor U4978 (N_4978,N_2657,N_3155);
nand U4979 (N_4979,N_3173,N_3220);
or U4980 (N_4980,N_2706,N_3237);
xor U4981 (N_4981,N_3394,N_3033);
and U4982 (N_4982,N_2867,N_2866);
xor U4983 (N_4983,N_2956,N_2611);
nand U4984 (N_4984,N_3364,N_3519);
xor U4985 (N_4985,N_2892,N_2604);
and U4986 (N_4986,N_2658,N_2655);
or U4987 (N_4987,N_3105,N_3277);
nand U4988 (N_4988,N_2986,N_3640);
nor U4989 (N_4989,N_2794,N_3559);
or U4990 (N_4990,N_3645,N_2583);
nand U4991 (N_4991,N_2543,N_2608);
nor U4992 (N_4992,N_2976,N_3281);
and U4993 (N_4993,N_2902,N_3085);
nand U4994 (N_4994,N_3408,N_3113);
nand U4995 (N_4995,N_2959,N_3268);
xnor U4996 (N_4996,N_2586,N_3136);
and U4997 (N_4997,N_3524,N_2542);
nand U4998 (N_4998,N_3077,N_3428);
nor U4999 (N_4999,N_3271,N_3356);
nand U5000 (N_5000,N_4719,N_4053);
nor U5001 (N_5001,N_4656,N_3839);
xor U5002 (N_5002,N_3838,N_3875);
nor U5003 (N_5003,N_4153,N_4019);
or U5004 (N_5004,N_3889,N_3771);
and U5005 (N_5005,N_4471,N_4553);
nor U5006 (N_5006,N_4340,N_4700);
or U5007 (N_5007,N_4076,N_4268);
xor U5008 (N_5008,N_3803,N_4399);
and U5009 (N_5009,N_4087,N_4410);
or U5010 (N_5010,N_4004,N_4417);
or U5011 (N_5011,N_4458,N_4002);
nor U5012 (N_5012,N_4708,N_4689);
nand U5013 (N_5013,N_4431,N_4230);
nor U5014 (N_5014,N_3904,N_4822);
xnor U5015 (N_5015,N_4829,N_3952);
xor U5016 (N_5016,N_4008,N_4118);
or U5017 (N_5017,N_3978,N_4762);
nand U5018 (N_5018,N_4786,N_4723);
xor U5019 (N_5019,N_4720,N_4824);
nor U5020 (N_5020,N_4047,N_4804);
xor U5021 (N_5021,N_4180,N_4310);
and U5022 (N_5022,N_4859,N_4332);
nand U5023 (N_5023,N_4074,N_4358);
xnor U5024 (N_5024,N_4551,N_4009);
nand U5025 (N_5025,N_4263,N_4450);
nand U5026 (N_5026,N_3821,N_4576);
xor U5027 (N_5027,N_4059,N_4351);
nand U5028 (N_5028,N_4269,N_4120);
nor U5029 (N_5029,N_3774,N_3807);
and U5030 (N_5030,N_3766,N_4368);
nand U5031 (N_5031,N_4667,N_3897);
nor U5032 (N_5032,N_3895,N_4549);
nor U5033 (N_5033,N_4906,N_4404);
nand U5034 (N_5034,N_4513,N_4803);
or U5035 (N_5035,N_4608,N_4485);
nor U5036 (N_5036,N_4344,N_4045);
xor U5037 (N_5037,N_4209,N_4609);
nor U5038 (N_5038,N_4502,N_4743);
and U5039 (N_5039,N_3922,N_4562);
and U5040 (N_5040,N_4379,N_4636);
nor U5041 (N_5041,N_4459,N_3997);
nand U5042 (N_5042,N_4691,N_3805);
xor U5043 (N_5043,N_4878,N_4833);
nand U5044 (N_5044,N_4106,N_4383);
and U5045 (N_5045,N_3806,N_4790);
nand U5046 (N_5046,N_4542,N_4797);
nor U5047 (N_5047,N_4114,N_4515);
nor U5048 (N_5048,N_4628,N_4623);
nand U5049 (N_5049,N_4799,N_4242);
nor U5050 (N_5050,N_3896,N_4999);
nor U5051 (N_5051,N_4684,N_4634);
nor U5052 (N_5052,N_3906,N_4967);
nand U5053 (N_5053,N_4856,N_4854);
xnor U5054 (N_5054,N_4082,N_4579);
or U5055 (N_5055,N_4674,N_4078);
and U5056 (N_5056,N_4255,N_4845);
xor U5057 (N_5057,N_4238,N_4001);
nor U5058 (N_5058,N_4452,N_4058);
xor U5059 (N_5059,N_3844,N_3768);
or U5060 (N_5060,N_4875,N_4131);
or U5061 (N_5061,N_4624,N_4936);
or U5062 (N_5062,N_4718,N_4466);
nand U5063 (N_5063,N_4121,N_4325);
or U5064 (N_5064,N_4827,N_4658);
and U5065 (N_5065,N_4503,N_4963);
or U5066 (N_5066,N_4319,N_4013);
or U5067 (N_5067,N_4802,N_4895);
nand U5068 (N_5068,N_4297,N_3798);
or U5069 (N_5069,N_4384,N_4166);
nand U5070 (N_5070,N_3886,N_4687);
nand U5071 (N_5071,N_4961,N_4470);
nor U5072 (N_5072,N_4710,N_4327);
xnor U5073 (N_5073,N_4888,N_4834);
nor U5074 (N_5074,N_4488,N_4475);
nor U5075 (N_5075,N_3971,N_4704);
nor U5076 (N_5076,N_3977,N_4188);
or U5077 (N_5077,N_4267,N_4215);
and U5078 (N_5078,N_4776,N_4205);
and U5079 (N_5079,N_4127,N_4218);
nand U5080 (N_5080,N_4148,N_4499);
nor U5081 (N_5081,N_4232,N_4398);
and U5082 (N_5082,N_4334,N_4435);
and U5083 (N_5083,N_4552,N_4280);
xor U5084 (N_5084,N_4200,N_4326);
nor U5085 (N_5085,N_4530,N_3877);
and U5086 (N_5086,N_4449,N_3827);
nand U5087 (N_5087,N_4742,N_3953);
nand U5088 (N_5088,N_4876,N_4807);
nand U5089 (N_5089,N_4525,N_4671);
nor U5090 (N_5090,N_3857,N_4226);
xor U5091 (N_5091,N_4300,N_3975);
nor U5092 (N_5092,N_4993,N_3939);
xor U5093 (N_5093,N_3752,N_3927);
and U5094 (N_5094,N_4025,N_4357);
and U5095 (N_5095,N_4080,N_3817);
nand U5096 (N_5096,N_4977,N_4314);
nand U5097 (N_5097,N_4543,N_4679);
nor U5098 (N_5098,N_4428,N_4778);
xnor U5099 (N_5099,N_4362,N_4491);
xnor U5100 (N_5100,N_4100,N_4145);
nor U5101 (N_5101,N_3945,N_4860);
nor U5102 (N_5102,N_4196,N_4464);
xnor U5103 (N_5103,N_3882,N_4261);
nor U5104 (N_5104,N_3826,N_3760);
or U5105 (N_5105,N_4213,N_4649);
and U5106 (N_5106,N_4590,N_4302);
nand U5107 (N_5107,N_4930,N_3893);
xor U5108 (N_5108,N_4821,N_4976);
xnor U5109 (N_5109,N_4840,N_4673);
nor U5110 (N_5110,N_3790,N_4770);
or U5111 (N_5111,N_4216,N_4482);
or U5112 (N_5112,N_4281,N_4190);
xor U5113 (N_5113,N_3993,N_4007);
nor U5114 (N_5114,N_4274,N_4419);
and U5115 (N_5115,N_4457,N_4165);
xor U5116 (N_5116,N_4725,N_4923);
xnor U5117 (N_5117,N_4746,N_4915);
and U5118 (N_5118,N_4254,N_3796);
and U5119 (N_5119,N_4713,N_4851);
nand U5120 (N_5120,N_4406,N_4387);
nor U5121 (N_5121,N_4638,N_4757);
nand U5122 (N_5122,N_4496,N_3932);
nand U5123 (N_5123,N_4115,N_4548);
and U5124 (N_5124,N_3923,N_3991);
nor U5125 (N_5125,N_3958,N_4338);
or U5126 (N_5126,N_3980,N_3900);
nand U5127 (N_5127,N_3847,N_4388);
and U5128 (N_5128,N_4819,N_4805);
and U5129 (N_5129,N_4555,N_4264);
nor U5130 (N_5130,N_4138,N_4451);
xnor U5131 (N_5131,N_4441,N_4093);
xor U5132 (N_5132,N_4554,N_4568);
xor U5133 (N_5133,N_3845,N_4390);
nand U5134 (N_5134,N_4806,N_4198);
and U5135 (N_5135,N_4126,N_4817);
and U5136 (N_5136,N_4577,N_4760);
nor U5137 (N_5137,N_4015,N_4316);
nand U5138 (N_5138,N_3959,N_4685);
and U5139 (N_5139,N_4333,N_4810);
xnor U5140 (N_5140,N_4887,N_4077);
xnor U5141 (N_5141,N_3884,N_4146);
or U5142 (N_5142,N_4686,N_4937);
and U5143 (N_5143,N_3899,N_4291);
xnor U5144 (N_5144,N_4092,N_4716);
and U5145 (N_5145,N_4486,N_4273);
nor U5146 (N_5146,N_3800,N_4905);
xor U5147 (N_5147,N_4779,N_3814);
or U5148 (N_5148,N_4174,N_4397);
xnor U5149 (N_5149,N_4870,N_4607);
xnor U5150 (N_5150,N_4473,N_4520);
nor U5151 (N_5151,N_4309,N_3762);
nand U5152 (N_5152,N_4260,N_4643);
or U5153 (N_5153,N_4155,N_4403);
or U5154 (N_5154,N_3957,N_4133);
xor U5155 (N_5155,N_4814,N_4957);
nand U5156 (N_5156,N_4071,N_3797);
nand U5157 (N_5157,N_4016,N_4423);
and U5158 (N_5158,N_4698,N_4563);
or U5159 (N_5159,N_3892,N_4154);
xnor U5160 (N_5160,N_4434,N_4212);
xnor U5161 (N_5161,N_4699,N_4282);
nand U5162 (N_5162,N_4633,N_3829);
or U5163 (N_5163,N_4992,N_4996);
or U5164 (N_5164,N_4935,N_4991);
and U5165 (N_5165,N_4376,N_3984);
and U5166 (N_5166,N_4510,N_3972);
nor U5167 (N_5167,N_4920,N_4601);
and U5168 (N_5168,N_3910,N_4744);
xnor U5169 (N_5169,N_4617,N_4170);
xor U5170 (N_5170,N_3960,N_4695);
xnor U5171 (N_5171,N_4570,N_4277);
and U5172 (N_5172,N_3843,N_4306);
xor U5173 (N_5173,N_4149,N_4670);
xor U5174 (N_5174,N_3990,N_4882);
nand U5175 (N_5175,N_4066,N_4248);
nor U5176 (N_5176,N_4613,N_4838);
nand U5177 (N_5177,N_4446,N_4245);
nor U5178 (N_5178,N_4831,N_4644);
and U5179 (N_5179,N_4561,N_4429);
nor U5180 (N_5180,N_4538,N_4857);
and U5181 (N_5181,N_4900,N_4861);
nor U5182 (N_5182,N_3954,N_4849);
xnor U5183 (N_5183,N_3869,N_4257);
or U5184 (N_5184,N_3824,N_4581);
nor U5185 (N_5185,N_3874,N_4067);
nor U5186 (N_5186,N_4756,N_3890);
nand U5187 (N_5187,N_4249,N_4294);
xnor U5188 (N_5188,N_4873,N_4328);
xor U5189 (N_5189,N_4924,N_4356);
nor U5190 (N_5190,N_4753,N_4278);
nand U5191 (N_5191,N_4727,N_4908);
xor U5192 (N_5192,N_4195,N_3983);
nand U5193 (N_5193,N_3795,N_3947);
nand U5194 (N_5194,N_4694,N_4521);
xor U5195 (N_5195,N_4023,N_4184);
or U5196 (N_5196,N_4081,N_4690);
or U5197 (N_5197,N_3979,N_3823);
xor U5198 (N_5198,N_4545,N_4096);
and U5199 (N_5199,N_3849,N_4569);
nand U5200 (N_5200,N_3846,N_4186);
or U5201 (N_5201,N_4233,N_3761);
nor U5202 (N_5202,N_3915,N_4970);
and U5203 (N_5203,N_4104,N_4841);
and U5204 (N_5204,N_4020,N_4714);
or U5205 (N_5205,N_3966,N_4626);
xnor U5206 (N_5206,N_4794,N_4764);
nor U5207 (N_5207,N_4490,N_4639);
xnor U5208 (N_5208,N_4741,N_4185);
xnor U5209 (N_5209,N_4947,N_4954);
or U5210 (N_5210,N_3940,N_4672);
or U5211 (N_5211,N_4311,N_4614);
and U5212 (N_5212,N_4536,N_4701);
nand U5213 (N_5213,N_4479,N_4228);
nor U5214 (N_5214,N_4495,N_4848);
and U5215 (N_5215,N_4172,N_4089);
nand U5216 (N_5216,N_4424,N_4842);
and U5217 (N_5217,N_4921,N_4312);
nand U5218 (N_5218,N_4645,N_3825);
and U5219 (N_5219,N_4094,N_4903);
xnor U5220 (N_5220,N_4504,N_4413);
nor U5221 (N_5221,N_3982,N_4012);
or U5222 (N_5222,N_4811,N_3773);
nor U5223 (N_5223,N_4589,N_3902);
xor U5224 (N_5224,N_4173,N_3986);
nor U5225 (N_5225,N_3763,N_4880);
and U5226 (N_5226,N_4051,N_4669);
nor U5227 (N_5227,N_3969,N_3935);
nand U5228 (N_5228,N_4181,N_4355);
nor U5229 (N_5229,N_4182,N_4111);
nor U5230 (N_5230,N_4474,N_4049);
or U5231 (N_5231,N_4550,N_3867);
nor U5232 (N_5232,N_4702,N_4892);
nor U5233 (N_5233,N_4421,N_4335);
nor U5234 (N_5234,N_4330,N_4011);
and U5235 (N_5235,N_4974,N_4914);
nand U5236 (N_5236,N_4763,N_4402);
xnor U5237 (N_5237,N_3819,N_4337);
nand U5238 (N_5238,N_4559,N_4780);
xor U5239 (N_5239,N_4734,N_3913);
nand U5240 (N_5240,N_4295,N_4313);
xnor U5241 (N_5241,N_3999,N_4984);
or U5242 (N_5242,N_4136,N_4864);
xnor U5243 (N_5243,N_3905,N_4140);
nor U5244 (N_5244,N_4632,N_4095);
or U5245 (N_5245,N_4444,N_4972);
and U5246 (N_5246,N_4604,N_3770);
nor U5247 (N_5247,N_4630,N_4083);
or U5248 (N_5248,N_4766,N_4505);
nor U5249 (N_5249,N_4676,N_3868);
nor U5250 (N_5250,N_3802,N_4792);
nand U5251 (N_5251,N_4073,N_3944);
nor U5252 (N_5252,N_4863,N_4054);
and U5253 (N_5253,N_3785,N_3961);
nand U5254 (N_5254,N_3811,N_4808);
and U5255 (N_5255,N_4729,N_4733);
nor U5256 (N_5256,N_4986,N_4227);
and U5257 (N_5257,N_4640,N_4442);
and U5258 (N_5258,N_4730,N_4637);
nand U5259 (N_5259,N_4363,N_4151);
or U5260 (N_5260,N_4222,N_4925);
and U5261 (N_5261,N_4517,N_4026);
nand U5262 (N_5262,N_3920,N_3938);
nand U5263 (N_5263,N_4949,N_4266);
or U5264 (N_5264,N_3791,N_4751);
nand U5265 (N_5265,N_4711,N_4271);
or U5266 (N_5266,N_4582,N_4005);
nand U5267 (N_5267,N_4580,N_4109);
or U5268 (N_5268,N_4422,N_4946);
xor U5269 (N_5269,N_4044,N_4270);
and U5270 (N_5270,N_4303,N_4783);
and U5271 (N_5271,N_4728,N_3888);
xor U5272 (N_5272,N_4627,N_4605);
xor U5273 (N_5273,N_4901,N_3778);
or U5274 (N_5274,N_4789,N_4646);
nor U5275 (N_5275,N_4324,N_4108);
nor U5276 (N_5276,N_4385,N_4307);
nand U5277 (N_5277,N_4341,N_4995);
or U5278 (N_5278,N_4354,N_4498);
xnor U5279 (N_5279,N_4688,N_4202);
xor U5280 (N_5280,N_4132,N_3912);
and U5281 (N_5281,N_4346,N_3842);
nand U5282 (N_5282,N_4463,N_4392);
or U5283 (N_5283,N_4465,N_4732);
and U5284 (N_5284,N_4612,N_3925);
nand U5285 (N_5285,N_4443,N_4339);
xor U5286 (N_5286,N_4506,N_4787);
or U5287 (N_5287,N_4349,N_4738);
or U5288 (N_5288,N_3767,N_4938);
or U5289 (N_5289,N_4668,N_4844);
and U5290 (N_5290,N_4225,N_4210);
xor U5291 (N_5291,N_4377,N_4365);
or U5292 (N_5292,N_4130,N_3883);
or U5293 (N_5293,N_4414,N_4231);
and U5294 (N_5294,N_4692,N_4918);
nand U5295 (N_5295,N_3914,N_4758);
nor U5296 (N_5296,N_4982,N_3919);
or U5297 (N_5297,N_4454,N_4801);
nand U5298 (N_5298,N_4476,N_4566);
or U5299 (N_5299,N_4142,N_4110);
xor U5300 (N_5300,N_4024,N_4010);
and U5301 (N_5301,N_4411,N_4620);
nand U5302 (N_5302,N_4603,N_3758);
xnor U5303 (N_5303,N_4572,N_4825);
nand U5304 (N_5304,N_4987,N_4176);
xor U5305 (N_5305,N_4765,N_4955);
nor U5306 (N_5306,N_4158,N_3908);
or U5307 (N_5307,N_4818,N_3786);
and U5308 (N_5308,N_3864,N_4430);
nor U5309 (N_5309,N_3981,N_4724);
and U5310 (N_5310,N_4432,N_3853);
nor U5311 (N_5311,N_4535,N_4735);
nor U5312 (N_5312,N_4754,N_4677);
nor U5313 (N_5313,N_4544,N_4843);
nand U5314 (N_5314,N_3815,N_4129);
nand U5315 (N_5315,N_4039,N_4380);
nor U5316 (N_5316,N_4438,N_4445);
xor U5317 (N_5317,N_4360,N_4740);
xnor U5318 (N_5318,N_3941,N_4647);
and U5319 (N_5319,N_4652,N_4796);
and U5320 (N_5320,N_4037,N_4512);
nand U5321 (N_5321,N_4769,N_4336);
and U5322 (N_5322,N_4602,N_3926);
and U5323 (N_5323,N_3873,N_4899);
or U5324 (N_5324,N_3759,N_4929);
or U5325 (N_5325,N_4983,N_4006);
xnor U5326 (N_5326,N_4211,N_4102);
or U5327 (N_5327,N_4033,N_4064);
and U5328 (N_5328,N_4162,N_4125);
or U5329 (N_5329,N_3801,N_4703);
nor U5330 (N_5330,N_3764,N_4469);
xor U5331 (N_5331,N_3934,N_4161);
xor U5332 (N_5332,N_4537,N_4409);
nor U5333 (N_5333,N_3929,N_4660);
nand U5334 (N_5334,N_4866,N_3784);
or U5335 (N_5335,N_4119,N_4830);
and U5336 (N_5336,N_4401,N_4235);
and U5337 (N_5337,N_3777,N_4298);
nor U5338 (N_5338,N_4862,N_4084);
xor U5339 (N_5339,N_4029,N_4147);
xor U5340 (N_5340,N_4017,N_4556);
nand U5341 (N_5341,N_4871,N_4284);
or U5342 (N_5342,N_4150,N_3994);
nor U5343 (N_5343,N_4042,N_4361);
nand U5344 (N_5344,N_3757,N_4426);
xor U5345 (N_5345,N_4846,N_4697);
or U5346 (N_5346,N_4560,N_4917);
nor U5347 (N_5347,N_4000,N_3996);
or U5348 (N_5348,N_4031,N_4460);
or U5349 (N_5349,N_3871,N_4169);
and U5350 (N_5350,N_3831,N_4412);
or U5351 (N_5351,N_4289,N_4893);
nor U5352 (N_5352,N_4919,N_3928);
or U5353 (N_5353,N_4781,N_4522);
nor U5354 (N_5354,N_4812,N_4139);
nor U5355 (N_5355,N_4113,N_3756);
xnor U5356 (N_5356,N_4301,N_4192);
xor U5357 (N_5357,N_4969,N_3963);
and U5358 (N_5358,N_4507,N_4706);
or U5359 (N_5359,N_3943,N_4199);
nor U5360 (N_5360,N_4400,N_4086);
nor U5361 (N_5361,N_3787,N_4985);
nor U5362 (N_5362,N_4953,N_3862);
and U5363 (N_5363,N_3809,N_4487);
or U5364 (N_5364,N_3917,N_4731);
nand U5365 (N_5365,N_4027,N_4912);
xnor U5366 (N_5366,N_4350,N_4839);
or U5367 (N_5367,N_4964,N_4558);
or U5368 (N_5368,N_4099,N_3985);
nor U5369 (N_5369,N_4610,N_4323);
xor U5370 (N_5370,N_4378,N_4853);
or U5371 (N_5371,N_4524,N_4041);
nand U5372 (N_5372,N_3863,N_3876);
and U5373 (N_5373,N_4911,N_4394);
xor U5374 (N_5374,N_4867,N_3813);
nor U5375 (N_5375,N_4540,N_4641);
xor U5376 (N_5376,N_4493,N_4107);
or U5377 (N_5377,N_4461,N_3832);
nor U5378 (N_5378,N_3841,N_4123);
nor U5379 (N_5379,N_4622,N_4455);
nand U5380 (N_5380,N_4193,N_4523);
nand U5381 (N_5381,N_4366,N_3789);
xor U5382 (N_5382,N_3881,N_3754);
or U5383 (N_5383,N_3916,N_4014);
or U5384 (N_5384,N_4299,N_4978);
nor U5385 (N_5385,N_4981,N_4865);
nor U5386 (N_5386,N_4234,N_4246);
nor U5387 (N_5387,N_3782,N_4030);
xnor U5388 (N_5388,N_3955,N_4791);
nand U5389 (N_5389,N_3860,N_4304);
and U5390 (N_5390,N_4948,N_4395);
xnor U5391 (N_5391,N_4533,N_4343);
nor U5392 (N_5392,N_3755,N_4747);
nand U5393 (N_5393,N_4886,N_4179);
nor U5394 (N_5394,N_4877,N_4879);
nor U5395 (N_5395,N_3967,N_3772);
and U5396 (N_5396,N_3851,N_3870);
xor U5397 (N_5397,N_3810,N_3992);
and U5398 (N_5398,N_4835,N_4750);
xor U5399 (N_5399,N_4960,N_4418);
and U5400 (N_5400,N_4069,N_3866);
nor U5401 (N_5401,N_4191,N_3834);
xnor U5402 (N_5402,N_4826,N_3780);
xor U5403 (N_5403,N_4897,N_4171);
nor U5404 (N_5404,N_4236,N_4480);
xor U5405 (N_5405,N_4910,N_4966);
nand U5406 (N_5406,N_4823,N_4056);
xnor U5407 (N_5407,N_4591,N_4492);
and U5408 (N_5408,N_4331,N_4881);
and U5409 (N_5409,N_4352,N_3924);
nand U5410 (N_5410,N_4253,N_4290);
xnor U5411 (N_5411,N_4945,N_4478);
nor U5412 (N_5412,N_4721,N_4600);
nand U5413 (N_5413,N_4160,N_4795);
xor U5414 (N_5414,N_4793,N_4588);
or U5415 (N_5415,N_4575,N_4275);
xnor U5416 (N_5416,N_4250,N_4828);
nand U5417 (N_5417,N_4484,N_4439);
nand U5418 (N_5418,N_4251,N_3995);
xnor U5419 (N_5419,N_4079,N_4128);
nand U5420 (N_5420,N_4229,N_4527);
and U5421 (N_5421,N_4813,N_4518);
nand U5422 (N_5422,N_3799,N_4836);
nor U5423 (N_5423,N_4772,N_3970);
nor U5424 (N_5424,N_4272,N_4050);
xor U5425 (N_5425,N_4497,N_4519);
nand U5426 (N_5426,N_3976,N_4705);
nor U5427 (N_5427,N_4364,N_4468);
xnor U5428 (N_5428,N_4292,N_4777);
and U5429 (N_5429,N_4574,N_4565);
xnor U5430 (N_5430,N_4666,N_4143);
xnor U5431 (N_5431,N_4869,N_4663);
nor U5432 (N_5432,N_4022,N_3854);
and U5433 (N_5433,N_4913,N_4427);
and U5434 (N_5434,N_4737,N_4405);
nand U5435 (N_5435,N_3885,N_4152);
and U5436 (N_5436,N_4648,N_4068);
xnor U5437 (N_5437,N_4683,N_4244);
nand U5438 (N_5438,N_4573,N_3769);
and U5439 (N_5439,N_3918,N_4767);
and U5440 (N_5440,N_4070,N_4951);
xnor U5441 (N_5441,N_3865,N_4651);
or U5442 (N_5442,N_4531,N_4768);
xor U5443 (N_5443,N_4407,N_4816);
xnor U5444 (N_5444,N_3948,N_3775);
xnor U5445 (N_5445,N_4509,N_4197);
and U5446 (N_5446,N_4852,N_4375);
nor U5447 (N_5447,N_4564,N_3901);
nor U5448 (N_5448,N_4965,N_4883);
xnor U5449 (N_5449,N_4595,N_3804);
and U5450 (N_5450,N_4578,N_3907);
nand U5451 (N_5451,N_3988,N_4489);
nand U5452 (N_5452,N_4534,N_3909);
nand U5453 (N_5453,N_3776,N_3818);
nand U5454 (N_5454,N_4980,N_4359);
nand U5455 (N_5455,N_4712,N_4103);
or U5456 (N_5456,N_4501,N_4782);
xor U5457 (N_5457,N_4771,N_3998);
or U5458 (N_5458,N_4526,N_4943);
xor U5459 (N_5459,N_4243,N_3987);
and U5460 (N_5460,N_4124,N_4884);
xor U5461 (N_5461,N_4722,N_4973);
nor U5462 (N_5462,N_4183,N_4208);
nor U5463 (N_5463,N_4137,N_4618);
or U5464 (N_5464,N_4276,N_4625);
and U5465 (N_5465,N_4085,N_4279);
nand U5466 (N_5466,N_4293,N_4097);
nand U5467 (N_5467,N_3812,N_4157);
nand U5468 (N_5468,N_4329,N_4653);
nand U5469 (N_5469,N_4988,N_4717);
and U5470 (N_5470,N_4707,N_4858);
nand U5471 (N_5471,N_4516,N_4063);
or U5472 (N_5472,N_4141,N_4396);
nand U5473 (N_5473,N_4511,N_3781);
nand U5474 (N_5474,N_3779,N_3879);
or U5475 (N_5475,N_4606,N_4483);
nand U5476 (N_5476,N_4745,N_4371);
and U5477 (N_5477,N_4416,N_4239);
nand U5478 (N_5478,N_4447,N_4597);
nor U5479 (N_5479,N_4353,N_4437);
or U5480 (N_5480,N_4933,N_3835);
or U5481 (N_5481,N_4664,N_4940);
xnor U5482 (N_5482,N_3792,N_4837);
and U5483 (N_5483,N_3751,N_4348);
nand U5484 (N_5484,N_4288,N_4386);
or U5485 (N_5485,N_3949,N_4749);
nand U5486 (N_5486,N_4959,N_3820);
or U5487 (N_5487,N_3933,N_3833);
and U5488 (N_5488,N_4621,N_4736);
nand U5489 (N_5489,N_4372,N_4391);
xnor U5490 (N_5490,N_4178,N_4305);
or U5491 (N_5491,N_4462,N_3837);
nor U5492 (N_5492,N_4583,N_4420);
and U5493 (N_5493,N_4134,N_4221);
or U5494 (N_5494,N_4979,N_4453);
or U5495 (N_5495,N_4798,N_4204);
nand U5496 (N_5496,N_4922,N_4481);
nor U5497 (N_5497,N_4320,N_4696);
or U5498 (N_5498,N_4532,N_3956);
and U5499 (N_5499,N_4164,N_4774);
and U5500 (N_5500,N_3968,N_4726);
or U5501 (N_5501,N_4994,N_4629);
and U5502 (N_5502,N_4259,N_4872);
or U5503 (N_5503,N_4809,N_4286);
nand U5504 (N_5504,N_4642,N_4389);
or U5505 (N_5505,N_4715,N_3930);
or U5506 (N_5506,N_3942,N_4370);
and U5507 (N_5507,N_4847,N_4885);
and U5508 (N_5508,N_4528,N_4832);
and U5509 (N_5509,N_4322,N_4262);
nor U5510 (N_5510,N_4675,N_4927);
and U5511 (N_5511,N_4285,N_4514);
nand U5512 (N_5512,N_4773,N_4003);
nand U5513 (N_5513,N_4784,N_4156);
nor U5514 (N_5514,N_4203,N_4367);
or U5515 (N_5515,N_4163,N_4956);
nor U5516 (N_5516,N_4587,N_4654);
xnor U5517 (N_5517,N_4105,N_4631);
nand U5518 (N_5518,N_3855,N_3964);
or U5519 (N_5519,N_3856,N_4962);
nor U5520 (N_5520,N_4214,N_3783);
nand U5521 (N_5521,N_4219,N_4678);
xor U5522 (N_5522,N_3848,N_4971);
and U5523 (N_5523,N_4494,N_4611);
nor U5524 (N_5524,N_3936,N_3816);
and U5525 (N_5525,N_3891,N_4061);
and U5526 (N_5526,N_3965,N_4998);
nor U5527 (N_5527,N_4062,N_4693);
and U5528 (N_5528,N_4223,N_4060);
nor U5529 (N_5529,N_3793,N_4159);
nor U5530 (N_5530,N_4187,N_4855);
xnor U5531 (N_5531,N_4018,N_3950);
and U5532 (N_5532,N_4889,N_3894);
nand U5533 (N_5533,N_4775,N_4529);
nor U5534 (N_5534,N_4932,N_3937);
nand U5535 (N_5535,N_3903,N_4373);
nand U5536 (N_5536,N_4101,N_4759);
or U5537 (N_5537,N_4425,N_4315);
xor U5538 (N_5538,N_3765,N_4065);
and U5539 (N_5539,N_4217,N_3872);
and U5540 (N_5540,N_4472,N_4036);
or U5541 (N_5541,N_4241,N_3852);
and U5542 (N_5542,N_4456,N_3946);
or U5543 (N_5543,N_4237,N_4944);
nor U5544 (N_5544,N_4584,N_4598);
xnor U5545 (N_5545,N_3911,N_4122);
nand U5546 (N_5546,N_4571,N_4308);
nor U5547 (N_5547,N_4616,N_4135);
or U5548 (N_5548,N_3962,N_4941);
or U5549 (N_5549,N_4500,N_4415);
nand U5550 (N_5550,N_4206,N_4934);
nor U5551 (N_5551,N_4755,N_4038);
or U5552 (N_5552,N_4896,N_3822);
xnor U5553 (N_5553,N_4931,N_3898);
xnor U5554 (N_5554,N_4635,N_4448);
and U5555 (N_5555,N_4318,N_4035);
nand U5556 (N_5556,N_4321,N_4477);
or U5557 (N_5557,N_4990,N_4592);
and U5558 (N_5558,N_4467,N_3753);
nand U5559 (N_5559,N_4393,N_4907);
and U5560 (N_5560,N_4252,N_4890);
xor U5561 (N_5561,N_4508,N_4599);
nand U5562 (N_5562,N_4369,N_4116);
nor U5563 (N_5563,N_4342,N_4317);
nor U5564 (N_5564,N_4098,N_4939);
xor U5565 (N_5565,N_4661,N_4258);
xnor U5566 (N_5566,N_4942,N_3794);
and U5567 (N_5567,N_4567,N_3861);
and U5568 (N_5568,N_4220,N_4247);
or U5569 (N_5569,N_4619,N_4975);
nor U5570 (N_5570,N_4032,N_4752);
xor U5571 (N_5571,N_4874,N_3750);
nor U5572 (N_5572,N_4546,N_4052);
or U5573 (N_5573,N_4168,N_4117);
nand U5574 (N_5574,N_4739,N_4194);
and U5575 (N_5575,N_4958,N_4594);
nor U5576 (N_5576,N_4057,N_4952);
nor U5577 (N_5577,N_4585,N_4904);
and U5578 (N_5578,N_4167,N_4680);
or U5579 (N_5579,N_4596,N_3973);
or U5580 (N_5580,N_3887,N_4655);
or U5581 (N_5581,N_4201,N_4997);
nand U5582 (N_5582,N_4382,N_4265);
nor U5583 (N_5583,N_3974,N_4224);
and U5584 (N_5584,N_4072,N_3931);
nand U5585 (N_5585,N_4021,N_4586);
nand U5586 (N_5586,N_4928,N_4709);
or U5587 (N_5587,N_4539,N_4968);
nor U5588 (N_5588,N_4761,N_4748);
and U5589 (N_5589,N_4894,N_4055);
nand U5590 (N_5590,N_4091,N_4433);
nor U5591 (N_5591,N_3840,N_4541);
xnor U5592 (N_5592,N_4815,N_3878);
xnor U5593 (N_5593,N_4650,N_4381);
and U5594 (N_5594,N_4909,N_4088);
or U5595 (N_5595,N_4090,N_3880);
nand U5596 (N_5596,N_4950,N_4665);
or U5597 (N_5597,N_4868,N_4046);
nand U5598 (N_5598,N_4593,N_4989);
or U5599 (N_5599,N_4785,N_3808);
nand U5600 (N_5600,N_4891,N_4615);
or U5601 (N_5601,N_4347,N_3921);
nor U5602 (N_5602,N_4408,N_3859);
xor U5603 (N_5603,N_4043,N_4283);
nor U5604 (N_5604,N_3836,N_4189);
nor U5605 (N_5605,N_4926,N_4800);
xnor U5606 (N_5606,N_4547,N_3858);
nand U5607 (N_5607,N_3788,N_4256);
xor U5608 (N_5608,N_4207,N_4902);
nor U5609 (N_5609,N_4557,N_4112);
and U5610 (N_5610,N_4681,N_4175);
and U5611 (N_5611,N_3989,N_4075);
xor U5612 (N_5612,N_4287,N_4659);
nand U5613 (N_5613,N_4048,N_3828);
nor U5614 (N_5614,N_4040,N_4436);
and U5615 (N_5615,N_4682,N_4374);
nor U5616 (N_5616,N_3951,N_4916);
xor U5617 (N_5617,N_4296,N_4034);
and U5618 (N_5618,N_4788,N_3850);
nand U5619 (N_5619,N_4850,N_4820);
nand U5620 (N_5620,N_4898,N_4662);
nor U5621 (N_5621,N_3830,N_4657);
or U5622 (N_5622,N_4028,N_4345);
or U5623 (N_5623,N_4440,N_4177);
nand U5624 (N_5624,N_4240,N_4144);
nand U5625 (N_5625,N_4941,N_3830);
and U5626 (N_5626,N_3911,N_4405);
or U5627 (N_5627,N_4164,N_4884);
and U5628 (N_5628,N_3808,N_3957);
xor U5629 (N_5629,N_4504,N_4930);
nor U5630 (N_5630,N_4748,N_4564);
or U5631 (N_5631,N_4391,N_4338);
or U5632 (N_5632,N_4219,N_4358);
or U5633 (N_5633,N_4046,N_4523);
or U5634 (N_5634,N_4273,N_4268);
and U5635 (N_5635,N_3952,N_4591);
nor U5636 (N_5636,N_4071,N_4159);
nand U5637 (N_5637,N_4112,N_3797);
xnor U5638 (N_5638,N_4988,N_4369);
xnor U5639 (N_5639,N_4212,N_4991);
and U5640 (N_5640,N_4919,N_4082);
nor U5641 (N_5641,N_4022,N_4816);
xnor U5642 (N_5642,N_3851,N_4967);
or U5643 (N_5643,N_3808,N_4686);
nor U5644 (N_5644,N_4214,N_4042);
nor U5645 (N_5645,N_4340,N_3762);
xnor U5646 (N_5646,N_4677,N_3943);
nor U5647 (N_5647,N_4794,N_3756);
xnor U5648 (N_5648,N_4864,N_4026);
and U5649 (N_5649,N_3777,N_4924);
nor U5650 (N_5650,N_4943,N_4704);
nand U5651 (N_5651,N_4671,N_3825);
and U5652 (N_5652,N_4447,N_3901);
and U5653 (N_5653,N_4620,N_4400);
nor U5654 (N_5654,N_4241,N_4998);
nor U5655 (N_5655,N_4913,N_4219);
or U5656 (N_5656,N_3938,N_4948);
or U5657 (N_5657,N_4262,N_4190);
and U5658 (N_5658,N_4177,N_4295);
xnor U5659 (N_5659,N_4062,N_4776);
or U5660 (N_5660,N_4146,N_3863);
and U5661 (N_5661,N_4910,N_4759);
nor U5662 (N_5662,N_4945,N_4938);
xor U5663 (N_5663,N_3789,N_4867);
or U5664 (N_5664,N_4865,N_3875);
xnor U5665 (N_5665,N_4903,N_4317);
nand U5666 (N_5666,N_4876,N_4862);
nor U5667 (N_5667,N_4549,N_4323);
and U5668 (N_5668,N_4629,N_4423);
nand U5669 (N_5669,N_4495,N_4779);
xor U5670 (N_5670,N_4859,N_4078);
xnor U5671 (N_5671,N_3963,N_3839);
xnor U5672 (N_5672,N_4178,N_4409);
or U5673 (N_5673,N_4300,N_4584);
or U5674 (N_5674,N_3763,N_4966);
or U5675 (N_5675,N_4647,N_4892);
xnor U5676 (N_5676,N_4286,N_4626);
xnor U5677 (N_5677,N_4943,N_4931);
and U5678 (N_5678,N_3958,N_4152);
nor U5679 (N_5679,N_4921,N_4306);
nand U5680 (N_5680,N_4072,N_3837);
or U5681 (N_5681,N_4661,N_4259);
and U5682 (N_5682,N_4726,N_4905);
nand U5683 (N_5683,N_3808,N_4983);
nand U5684 (N_5684,N_3980,N_4415);
xor U5685 (N_5685,N_4487,N_4735);
xnor U5686 (N_5686,N_4755,N_4402);
nand U5687 (N_5687,N_4061,N_4911);
nor U5688 (N_5688,N_4104,N_4776);
nor U5689 (N_5689,N_4751,N_4212);
xor U5690 (N_5690,N_4262,N_4921);
or U5691 (N_5691,N_4094,N_4258);
nor U5692 (N_5692,N_4561,N_4461);
nor U5693 (N_5693,N_4687,N_4810);
xnor U5694 (N_5694,N_4659,N_3923);
nand U5695 (N_5695,N_4993,N_4632);
xnor U5696 (N_5696,N_4910,N_4546);
xor U5697 (N_5697,N_3900,N_4993);
or U5698 (N_5698,N_4844,N_4480);
and U5699 (N_5699,N_3865,N_4306);
nor U5700 (N_5700,N_3880,N_4324);
xnor U5701 (N_5701,N_4055,N_4509);
nor U5702 (N_5702,N_4528,N_4857);
nand U5703 (N_5703,N_4655,N_4650);
xnor U5704 (N_5704,N_4591,N_4714);
nand U5705 (N_5705,N_4765,N_4807);
and U5706 (N_5706,N_4305,N_4917);
xor U5707 (N_5707,N_4482,N_4149);
and U5708 (N_5708,N_4063,N_4376);
nor U5709 (N_5709,N_4692,N_4385);
and U5710 (N_5710,N_4126,N_4042);
xnor U5711 (N_5711,N_4113,N_4525);
xnor U5712 (N_5712,N_4242,N_4659);
or U5713 (N_5713,N_4627,N_4048);
xor U5714 (N_5714,N_4178,N_4821);
xnor U5715 (N_5715,N_3922,N_4350);
or U5716 (N_5716,N_4610,N_4902);
or U5717 (N_5717,N_4784,N_4877);
nor U5718 (N_5718,N_4644,N_3753);
or U5719 (N_5719,N_4972,N_4685);
nor U5720 (N_5720,N_4369,N_4987);
xor U5721 (N_5721,N_3906,N_3783);
nand U5722 (N_5722,N_4053,N_4802);
xnor U5723 (N_5723,N_4725,N_4232);
or U5724 (N_5724,N_4460,N_4125);
or U5725 (N_5725,N_4509,N_4498);
or U5726 (N_5726,N_4031,N_4847);
and U5727 (N_5727,N_3761,N_4995);
xor U5728 (N_5728,N_4820,N_4849);
nor U5729 (N_5729,N_4751,N_4424);
nand U5730 (N_5730,N_4693,N_4399);
or U5731 (N_5731,N_3994,N_3973);
or U5732 (N_5732,N_4608,N_4348);
xnor U5733 (N_5733,N_3890,N_4337);
or U5734 (N_5734,N_4805,N_4973);
or U5735 (N_5735,N_4812,N_4381);
and U5736 (N_5736,N_4419,N_3967);
nand U5737 (N_5737,N_4081,N_4214);
and U5738 (N_5738,N_4409,N_3958);
or U5739 (N_5739,N_4753,N_3775);
and U5740 (N_5740,N_4547,N_4198);
nor U5741 (N_5741,N_3908,N_4605);
nand U5742 (N_5742,N_4072,N_4310);
nand U5743 (N_5743,N_4555,N_4010);
nand U5744 (N_5744,N_4772,N_4362);
xor U5745 (N_5745,N_4090,N_4730);
or U5746 (N_5746,N_4586,N_4731);
xnor U5747 (N_5747,N_4381,N_4019);
and U5748 (N_5748,N_4544,N_4072);
nand U5749 (N_5749,N_4773,N_4220);
nor U5750 (N_5750,N_4664,N_3864);
or U5751 (N_5751,N_4206,N_4488);
and U5752 (N_5752,N_4274,N_4895);
or U5753 (N_5753,N_4667,N_4072);
nand U5754 (N_5754,N_4653,N_4974);
and U5755 (N_5755,N_4664,N_4896);
nand U5756 (N_5756,N_4155,N_4629);
and U5757 (N_5757,N_4729,N_4297);
xnor U5758 (N_5758,N_4621,N_3954);
xnor U5759 (N_5759,N_4141,N_4286);
nand U5760 (N_5760,N_4136,N_4782);
or U5761 (N_5761,N_4188,N_4636);
nor U5762 (N_5762,N_4522,N_4721);
and U5763 (N_5763,N_4878,N_3812);
and U5764 (N_5764,N_3979,N_4944);
and U5765 (N_5765,N_4746,N_4725);
or U5766 (N_5766,N_4554,N_4906);
xnor U5767 (N_5767,N_4362,N_4834);
xnor U5768 (N_5768,N_4854,N_4456);
and U5769 (N_5769,N_3816,N_4388);
and U5770 (N_5770,N_4728,N_4029);
xor U5771 (N_5771,N_4219,N_4352);
nor U5772 (N_5772,N_4945,N_4261);
or U5773 (N_5773,N_4134,N_3925);
and U5774 (N_5774,N_3806,N_4162);
or U5775 (N_5775,N_4012,N_4062);
nor U5776 (N_5776,N_4902,N_4141);
or U5777 (N_5777,N_4293,N_4088);
nor U5778 (N_5778,N_3789,N_3816);
nor U5779 (N_5779,N_4768,N_4180);
nand U5780 (N_5780,N_4782,N_4045);
nand U5781 (N_5781,N_4251,N_4032);
or U5782 (N_5782,N_4614,N_4978);
nand U5783 (N_5783,N_4851,N_4172);
xnor U5784 (N_5784,N_4282,N_4513);
nand U5785 (N_5785,N_4817,N_3976);
or U5786 (N_5786,N_4696,N_3999);
or U5787 (N_5787,N_4990,N_4734);
or U5788 (N_5788,N_4089,N_3947);
or U5789 (N_5789,N_4705,N_3864);
nor U5790 (N_5790,N_4197,N_4085);
xnor U5791 (N_5791,N_4532,N_4767);
xnor U5792 (N_5792,N_4520,N_4334);
xor U5793 (N_5793,N_4365,N_4271);
xor U5794 (N_5794,N_4221,N_3904);
xor U5795 (N_5795,N_4886,N_4723);
nand U5796 (N_5796,N_4501,N_4230);
and U5797 (N_5797,N_4021,N_4118);
nor U5798 (N_5798,N_4552,N_4257);
and U5799 (N_5799,N_4611,N_4655);
nand U5800 (N_5800,N_4743,N_4731);
and U5801 (N_5801,N_4670,N_4796);
and U5802 (N_5802,N_4822,N_4929);
nor U5803 (N_5803,N_4245,N_4233);
xnor U5804 (N_5804,N_4122,N_4663);
nor U5805 (N_5805,N_4656,N_4659);
nand U5806 (N_5806,N_4363,N_4195);
and U5807 (N_5807,N_4386,N_4273);
nand U5808 (N_5808,N_4197,N_4347);
and U5809 (N_5809,N_4009,N_3957);
and U5810 (N_5810,N_4190,N_4181);
nand U5811 (N_5811,N_3989,N_4458);
nand U5812 (N_5812,N_3955,N_4572);
nand U5813 (N_5813,N_4379,N_4246);
and U5814 (N_5814,N_4576,N_4066);
nor U5815 (N_5815,N_4714,N_4563);
and U5816 (N_5816,N_4770,N_4797);
and U5817 (N_5817,N_3892,N_4542);
and U5818 (N_5818,N_4327,N_3869);
nand U5819 (N_5819,N_4335,N_4774);
and U5820 (N_5820,N_4449,N_4118);
nor U5821 (N_5821,N_4658,N_4960);
xor U5822 (N_5822,N_4857,N_3955);
nor U5823 (N_5823,N_3803,N_3941);
nand U5824 (N_5824,N_3996,N_4284);
or U5825 (N_5825,N_3995,N_4703);
xor U5826 (N_5826,N_4613,N_3970);
xor U5827 (N_5827,N_4511,N_4562);
or U5828 (N_5828,N_4158,N_3776);
xnor U5829 (N_5829,N_4047,N_4475);
and U5830 (N_5830,N_4387,N_4130);
or U5831 (N_5831,N_4777,N_4608);
xnor U5832 (N_5832,N_4329,N_4298);
xnor U5833 (N_5833,N_4212,N_4378);
nor U5834 (N_5834,N_4414,N_4012);
nand U5835 (N_5835,N_4321,N_4935);
or U5836 (N_5836,N_4772,N_4753);
nor U5837 (N_5837,N_4200,N_4983);
or U5838 (N_5838,N_4443,N_4224);
nand U5839 (N_5839,N_3796,N_4680);
nand U5840 (N_5840,N_4437,N_3954);
nor U5841 (N_5841,N_3765,N_4317);
and U5842 (N_5842,N_4133,N_3915);
or U5843 (N_5843,N_4843,N_4566);
xnor U5844 (N_5844,N_4510,N_4283);
nor U5845 (N_5845,N_4304,N_4323);
nor U5846 (N_5846,N_4657,N_3804);
xor U5847 (N_5847,N_4695,N_4752);
nand U5848 (N_5848,N_4864,N_3898);
xnor U5849 (N_5849,N_3814,N_4411);
nand U5850 (N_5850,N_4634,N_4549);
nand U5851 (N_5851,N_4765,N_4359);
or U5852 (N_5852,N_3753,N_4780);
or U5853 (N_5853,N_4165,N_4239);
nand U5854 (N_5854,N_4683,N_3875);
nor U5855 (N_5855,N_4350,N_3923);
xor U5856 (N_5856,N_4742,N_4912);
xor U5857 (N_5857,N_3865,N_3791);
or U5858 (N_5858,N_4782,N_4932);
or U5859 (N_5859,N_4342,N_4761);
nand U5860 (N_5860,N_4711,N_4799);
nand U5861 (N_5861,N_4587,N_4964);
xor U5862 (N_5862,N_3922,N_4175);
and U5863 (N_5863,N_4899,N_4319);
and U5864 (N_5864,N_4392,N_4635);
and U5865 (N_5865,N_4893,N_4360);
nor U5866 (N_5866,N_4336,N_4720);
xor U5867 (N_5867,N_3882,N_4315);
xnor U5868 (N_5868,N_4827,N_4193);
or U5869 (N_5869,N_4700,N_4994);
nor U5870 (N_5870,N_3861,N_3883);
nor U5871 (N_5871,N_4752,N_4533);
nor U5872 (N_5872,N_4895,N_4177);
or U5873 (N_5873,N_3881,N_4071);
xnor U5874 (N_5874,N_3809,N_4173);
and U5875 (N_5875,N_4821,N_4738);
xor U5876 (N_5876,N_4752,N_4028);
nor U5877 (N_5877,N_4398,N_4526);
nand U5878 (N_5878,N_4891,N_4243);
xor U5879 (N_5879,N_3837,N_4577);
and U5880 (N_5880,N_4468,N_4611);
and U5881 (N_5881,N_4620,N_3870);
nor U5882 (N_5882,N_4141,N_4038);
or U5883 (N_5883,N_4528,N_4072);
and U5884 (N_5884,N_3935,N_4644);
and U5885 (N_5885,N_4718,N_4418);
xnor U5886 (N_5886,N_4225,N_3789);
nand U5887 (N_5887,N_4232,N_4328);
nand U5888 (N_5888,N_4602,N_4784);
nor U5889 (N_5889,N_4891,N_3765);
nand U5890 (N_5890,N_3970,N_4678);
and U5891 (N_5891,N_3851,N_3824);
and U5892 (N_5892,N_4323,N_4983);
and U5893 (N_5893,N_4129,N_4399);
nor U5894 (N_5894,N_4806,N_4746);
and U5895 (N_5895,N_3981,N_3792);
xor U5896 (N_5896,N_4305,N_4182);
or U5897 (N_5897,N_4543,N_4860);
or U5898 (N_5898,N_4520,N_4725);
or U5899 (N_5899,N_4047,N_4675);
nand U5900 (N_5900,N_3880,N_4876);
xnor U5901 (N_5901,N_3773,N_3975);
nand U5902 (N_5902,N_3785,N_4667);
and U5903 (N_5903,N_4065,N_4616);
or U5904 (N_5904,N_4090,N_3936);
xor U5905 (N_5905,N_4473,N_3760);
nand U5906 (N_5906,N_3836,N_4233);
or U5907 (N_5907,N_3948,N_4442);
and U5908 (N_5908,N_3842,N_4250);
or U5909 (N_5909,N_3868,N_4284);
or U5910 (N_5910,N_4992,N_4276);
or U5911 (N_5911,N_4297,N_4232);
xor U5912 (N_5912,N_4796,N_4264);
xnor U5913 (N_5913,N_4896,N_4778);
nor U5914 (N_5914,N_4419,N_4281);
and U5915 (N_5915,N_4082,N_4332);
nor U5916 (N_5916,N_4690,N_4790);
xor U5917 (N_5917,N_3838,N_3964);
xnor U5918 (N_5918,N_3768,N_4577);
xnor U5919 (N_5919,N_4034,N_4039);
xor U5920 (N_5920,N_4757,N_4963);
or U5921 (N_5921,N_4580,N_4673);
nand U5922 (N_5922,N_4689,N_3968);
and U5923 (N_5923,N_4078,N_4297);
and U5924 (N_5924,N_4206,N_4128);
nand U5925 (N_5925,N_4594,N_4569);
nor U5926 (N_5926,N_4030,N_4333);
and U5927 (N_5927,N_4566,N_4041);
xnor U5928 (N_5928,N_4273,N_3813);
and U5929 (N_5929,N_4115,N_3879);
xnor U5930 (N_5930,N_4829,N_4312);
nand U5931 (N_5931,N_4021,N_4547);
nor U5932 (N_5932,N_4982,N_3896);
nand U5933 (N_5933,N_3964,N_4964);
nor U5934 (N_5934,N_4753,N_4911);
or U5935 (N_5935,N_4234,N_4668);
and U5936 (N_5936,N_4507,N_4482);
nor U5937 (N_5937,N_4504,N_3904);
and U5938 (N_5938,N_4316,N_4531);
nand U5939 (N_5939,N_4530,N_4613);
xor U5940 (N_5940,N_4804,N_4566);
xor U5941 (N_5941,N_4118,N_4047);
xor U5942 (N_5942,N_4858,N_4643);
and U5943 (N_5943,N_4430,N_3961);
or U5944 (N_5944,N_4868,N_4623);
xor U5945 (N_5945,N_4328,N_4754);
nand U5946 (N_5946,N_3924,N_3858);
nand U5947 (N_5947,N_3905,N_4504);
nand U5948 (N_5948,N_4305,N_4470);
nor U5949 (N_5949,N_4664,N_4007);
nor U5950 (N_5950,N_4040,N_4467);
and U5951 (N_5951,N_4188,N_4709);
nor U5952 (N_5952,N_4520,N_4901);
xnor U5953 (N_5953,N_4665,N_4562);
and U5954 (N_5954,N_3845,N_4288);
and U5955 (N_5955,N_4034,N_4546);
and U5956 (N_5956,N_4293,N_4680);
nor U5957 (N_5957,N_4375,N_3819);
nand U5958 (N_5958,N_3914,N_4797);
and U5959 (N_5959,N_3860,N_3966);
or U5960 (N_5960,N_4433,N_3755);
and U5961 (N_5961,N_4719,N_4571);
nand U5962 (N_5962,N_4699,N_3966);
nand U5963 (N_5963,N_4379,N_3875);
xnor U5964 (N_5964,N_4185,N_3956);
or U5965 (N_5965,N_4177,N_4199);
xor U5966 (N_5966,N_4933,N_4739);
xnor U5967 (N_5967,N_4998,N_4260);
xnor U5968 (N_5968,N_4134,N_4189);
nand U5969 (N_5969,N_4589,N_4744);
nand U5970 (N_5970,N_4272,N_3925);
nand U5971 (N_5971,N_4354,N_4178);
and U5972 (N_5972,N_4367,N_4047);
and U5973 (N_5973,N_4515,N_4294);
nor U5974 (N_5974,N_4915,N_4886);
or U5975 (N_5975,N_4436,N_4995);
nand U5976 (N_5976,N_4939,N_4571);
and U5977 (N_5977,N_4070,N_4725);
nor U5978 (N_5978,N_4738,N_3762);
nor U5979 (N_5979,N_4594,N_4983);
or U5980 (N_5980,N_3905,N_4512);
nor U5981 (N_5981,N_4405,N_4830);
and U5982 (N_5982,N_3966,N_4039);
and U5983 (N_5983,N_4876,N_4770);
nor U5984 (N_5984,N_3898,N_3862);
nand U5985 (N_5985,N_4412,N_4770);
or U5986 (N_5986,N_4516,N_4985);
xnor U5987 (N_5987,N_4351,N_4221);
and U5988 (N_5988,N_4646,N_4975);
nor U5989 (N_5989,N_4822,N_4118);
nand U5990 (N_5990,N_4491,N_4987);
and U5991 (N_5991,N_4130,N_4183);
xor U5992 (N_5992,N_4325,N_4905);
nand U5993 (N_5993,N_3838,N_4954);
nand U5994 (N_5994,N_4409,N_4018);
nand U5995 (N_5995,N_4079,N_4923);
and U5996 (N_5996,N_4548,N_3871);
xnor U5997 (N_5997,N_4031,N_3901);
nor U5998 (N_5998,N_3859,N_4679);
or U5999 (N_5999,N_4101,N_4238);
nor U6000 (N_6000,N_4045,N_4975);
xnor U6001 (N_6001,N_4173,N_4953);
or U6002 (N_6002,N_4545,N_3884);
xnor U6003 (N_6003,N_4661,N_4678);
and U6004 (N_6004,N_4203,N_4835);
and U6005 (N_6005,N_3961,N_4575);
nand U6006 (N_6006,N_4836,N_4357);
and U6007 (N_6007,N_4114,N_3796);
and U6008 (N_6008,N_4210,N_3804);
and U6009 (N_6009,N_4554,N_4308);
and U6010 (N_6010,N_4936,N_4551);
nor U6011 (N_6011,N_4937,N_4448);
and U6012 (N_6012,N_4966,N_3963);
or U6013 (N_6013,N_3784,N_4666);
and U6014 (N_6014,N_4751,N_3973);
nor U6015 (N_6015,N_4221,N_4633);
nor U6016 (N_6016,N_4303,N_4760);
nor U6017 (N_6017,N_4986,N_4085);
xor U6018 (N_6018,N_4040,N_4951);
xor U6019 (N_6019,N_4198,N_3860);
nor U6020 (N_6020,N_4722,N_4250);
and U6021 (N_6021,N_4693,N_4568);
or U6022 (N_6022,N_3780,N_4470);
nand U6023 (N_6023,N_4396,N_4733);
and U6024 (N_6024,N_4537,N_4704);
or U6025 (N_6025,N_4683,N_4674);
nand U6026 (N_6026,N_3870,N_4595);
nor U6027 (N_6027,N_4782,N_4731);
nor U6028 (N_6028,N_4561,N_4909);
nor U6029 (N_6029,N_4741,N_4213);
and U6030 (N_6030,N_4704,N_4104);
and U6031 (N_6031,N_4025,N_3860);
nor U6032 (N_6032,N_3880,N_4823);
xnor U6033 (N_6033,N_4397,N_4389);
nor U6034 (N_6034,N_4236,N_4330);
xnor U6035 (N_6035,N_4035,N_4736);
nor U6036 (N_6036,N_4181,N_4602);
nor U6037 (N_6037,N_4222,N_4950);
nand U6038 (N_6038,N_4677,N_3845);
nand U6039 (N_6039,N_4284,N_4472);
nand U6040 (N_6040,N_4335,N_4527);
and U6041 (N_6041,N_4804,N_4598);
xnor U6042 (N_6042,N_4238,N_4643);
and U6043 (N_6043,N_4335,N_4831);
xor U6044 (N_6044,N_4663,N_4319);
or U6045 (N_6045,N_3771,N_4830);
or U6046 (N_6046,N_3886,N_4621);
and U6047 (N_6047,N_4813,N_4848);
xnor U6048 (N_6048,N_4884,N_4485);
nand U6049 (N_6049,N_4014,N_4531);
and U6050 (N_6050,N_3841,N_4797);
nor U6051 (N_6051,N_3779,N_4061);
or U6052 (N_6052,N_4738,N_4720);
nand U6053 (N_6053,N_4673,N_4563);
and U6054 (N_6054,N_4991,N_4853);
nor U6055 (N_6055,N_4473,N_3877);
xnor U6056 (N_6056,N_4807,N_4771);
or U6057 (N_6057,N_3796,N_3809);
and U6058 (N_6058,N_4046,N_3830);
nor U6059 (N_6059,N_4058,N_4194);
nand U6060 (N_6060,N_4750,N_4663);
nor U6061 (N_6061,N_3829,N_4309);
xnor U6062 (N_6062,N_4170,N_4353);
xnor U6063 (N_6063,N_4303,N_4192);
nand U6064 (N_6064,N_4905,N_4753);
or U6065 (N_6065,N_3865,N_4022);
xor U6066 (N_6066,N_4573,N_4439);
or U6067 (N_6067,N_4391,N_4200);
nor U6068 (N_6068,N_4823,N_4460);
and U6069 (N_6069,N_4543,N_4769);
or U6070 (N_6070,N_3847,N_4445);
nand U6071 (N_6071,N_4588,N_4423);
and U6072 (N_6072,N_3862,N_3884);
xnor U6073 (N_6073,N_4582,N_3945);
and U6074 (N_6074,N_3845,N_3966);
nor U6075 (N_6075,N_4536,N_4670);
nand U6076 (N_6076,N_4293,N_3925);
nor U6077 (N_6077,N_4715,N_4068);
nand U6078 (N_6078,N_4440,N_4621);
xnor U6079 (N_6079,N_4031,N_4912);
nor U6080 (N_6080,N_4251,N_4853);
xnor U6081 (N_6081,N_4859,N_3760);
xor U6082 (N_6082,N_4665,N_3917);
and U6083 (N_6083,N_4793,N_3996);
nand U6084 (N_6084,N_4046,N_4288);
or U6085 (N_6085,N_4354,N_4798);
and U6086 (N_6086,N_3831,N_3821);
xor U6087 (N_6087,N_4944,N_4859);
or U6088 (N_6088,N_4698,N_4384);
or U6089 (N_6089,N_4296,N_4395);
nor U6090 (N_6090,N_4278,N_4696);
xor U6091 (N_6091,N_4849,N_4701);
xnor U6092 (N_6092,N_4682,N_4970);
nand U6093 (N_6093,N_4134,N_4861);
xnor U6094 (N_6094,N_4466,N_4378);
nand U6095 (N_6095,N_4966,N_4057);
and U6096 (N_6096,N_3784,N_4263);
nand U6097 (N_6097,N_4584,N_3878);
or U6098 (N_6098,N_3988,N_4728);
nand U6099 (N_6099,N_4361,N_4525);
nor U6100 (N_6100,N_4232,N_4283);
or U6101 (N_6101,N_4525,N_4226);
xor U6102 (N_6102,N_4240,N_3875);
nand U6103 (N_6103,N_4192,N_4460);
nand U6104 (N_6104,N_3777,N_4724);
nand U6105 (N_6105,N_4842,N_4102);
and U6106 (N_6106,N_4386,N_4322);
nand U6107 (N_6107,N_4659,N_4144);
nand U6108 (N_6108,N_3998,N_3959);
or U6109 (N_6109,N_4734,N_3957);
nand U6110 (N_6110,N_3826,N_4890);
xor U6111 (N_6111,N_4317,N_4356);
nor U6112 (N_6112,N_4881,N_3950);
or U6113 (N_6113,N_4932,N_4967);
or U6114 (N_6114,N_4976,N_4607);
nor U6115 (N_6115,N_4902,N_4357);
nor U6116 (N_6116,N_3843,N_4363);
xor U6117 (N_6117,N_4799,N_4216);
and U6118 (N_6118,N_4301,N_4508);
nor U6119 (N_6119,N_3856,N_3971);
and U6120 (N_6120,N_4447,N_4412);
and U6121 (N_6121,N_4332,N_4498);
xnor U6122 (N_6122,N_3882,N_4722);
or U6123 (N_6123,N_3971,N_4907);
or U6124 (N_6124,N_3766,N_4898);
or U6125 (N_6125,N_4556,N_3811);
nor U6126 (N_6126,N_4250,N_4513);
and U6127 (N_6127,N_4182,N_3874);
and U6128 (N_6128,N_4402,N_4167);
and U6129 (N_6129,N_4048,N_4290);
nand U6130 (N_6130,N_4595,N_4169);
nand U6131 (N_6131,N_4755,N_4342);
or U6132 (N_6132,N_4226,N_4622);
nand U6133 (N_6133,N_4166,N_4503);
nand U6134 (N_6134,N_4104,N_4365);
or U6135 (N_6135,N_4783,N_4043);
xor U6136 (N_6136,N_4819,N_4420);
or U6137 (N_6137,N_4222,N_4228);
xnor U6138 (N_6138,N_4282,N_4649);
xnor U6139 (N_6139,N_4468,N_4911);
xor U6140 (N_6140,N_4346,N_4201);
nor U6141 (N_6141,N_3765,N_4192);
nor U6142 (N_6142,N_3986,N_4587);
nor U6143 (N_6143,N_4457,N_3820);
or U6144 (N_6144,N_4349,N_4538);
xor U6145 (N_6145,N_4162,N_4025);
and U6146 (N_6146,N_4364,N_4415);
and U6147 (N_6147,N_4015,N_4469);
xor U6148 (N_6148,N_4418,N_4158);
or U6149 (N_6149,N_4639,N_4054);
nor U6150 (N_6150,N_4242,N_4704);
or U6151 (N_6151,N_3963,N_4828);
nand U6152 (N_6152,N_4972,N_4486);
nor U6153 (N_6153,N_4575,N_3775);
or U6154 (N_6154,N_3837,N_4730);
nand U6155 (N_6155,N_4986,N_4909);
nor U6156 (N_6156,N_4685,N_4791);
xnor U6157 (N_6157,N_4966,N_4406);
xnor U6158 (N_6158,N_4959,N_4638);
xnor U6159 (N_6159,N_4508,N_4655);
and U6160 (N_6160,N_3794,N_4529);
and U6161 (N_6161,N_3756,N_4095);
nor U6162 (N_6162,N_4314,N_4394);
or U6163 (N_6163,N_4826,N_4604);
xor U6164 (N_6164,N_4099,N_4624);
and U6165 (N_6165,N_4611,N_4851);
or U6166 (N_6166,N_4122,N_4861);
nand U6167 (N_6167,N_3754,N_4899);
and U6168 (N_6168,N_3859,N_4971);
nor U6169 (N_6169,N_4442,N_4004);
xor U6170 (N_6170,N_4837,N_4222);
or U6171 (N_6171,N_4958,N_4415);
nor U6172 (N_6172,N_4170,N_4862);
nand U6173 (N_6173,N_4632,N_3765);
nor U6174 (N_6174,N_3766,N_4320);
nand U6175 (N_6175,N_3931,N_4963);
xor U6176 (N_6176,N_4562,N_4557);
and U6177 (N_6177,N_4915,N_4544);
or U6178 (N_6178,N_4472,N_4626);
xnor U6179 (N_6179,N_4871,N_4018);
or U6180 (N_6180,N_4014,N_4280);
nand U6181 (N_6181,N_3842,N_4097);
xor U6182 (N_6182,N_4005,N_4154);
nand U6183 (N_6183,N_4981,N_4619);
and U6184 (N_6184,N_4451,N_4155);
and U6185 (N_6185,N_4601,N_4854);
nand U6186 (N_6186,N_4074,N_4549);
nand U6187 (N_6187,N_4852,N_4933);
or U6188 (N_6188,N_4643,N_4219);
and U6189 (N_6189,N_4462,N_4256);
and U6190 (N_6190,N_3975,N_3767);
or U6191 (N_6191,N_3860,N_4218);
nand U6192 (N_6192,N_4354,N_3789);
and U6193 (N_6193,N_3888,N_4387);
xor U6194 (N_6194,N_4838,N_4298);
nor U6195 (N_6195,N_4651,N_4252);
and U6196 (N_6196,N_4577,N_4543);
and U6197 (N_6197,N_4050,N_4175);
nor U6198 (N_6198,N_4743,N_4033);
and U6199 (N_6199,N_4306,N_4293);
and U6200 (N_6200,N_4458,N_4356);
xnor U6201 (N_6201,N_4094,N_4367);
or U6202 (N_6202,N_4002,N_3996);
nand U6203 (N_6203,N_4684,N_4306);
nand U6204 (N_6204,N_4794,N_4470);
nand U6205 (N_6205,N_4510,N_4177);
and U6206 (N_6206,N_3821,N_4934);
nand U6207 (N_6207,N_4738,N_4848);
and U6208 (N_6208,N_3853,N_4120);
nor U6209 (N_6209,N_4455,N_4409);
xnor U6210 (N_6210,N_4913,N_4798);
and U6211 (N_6211,N_4354,N_4118);
xnor U6212 (N_6212,N_3840,N_4039);
or U6213 (N_6213,N_4406,N_4196);
xor U6214 (N_6214,N_4799,N_4295);
xnor U6215 (N_6215,N_4654,N_4505);
nor U6216 (N_6216,N_4801,N_3987);
nand U6217 (N_6217,N_4257,N_3950);
nand U6218 (N_6218,N_4970,N_4475);
nand U6219 (N_6219,N_4096,N_4787);
nor U6220 (N_6220,N_4012,N_3774);
nor U6221 (N_6221,N_3804,N_3756);
xnor U6222 (N_6222,N_4535,N_4137);
or U6223 (N_6223,N_4853,N_4657);
or U6224 (N_6224,N_4720,N_4345);
or U6225 (N_6225,N_4532,N_4259);
nand U6226 (N_6226,N_3994,N_3775);
and U6227 (N_6227,N_4035,N_4641);
nor U6228 (N_6228,N_4360,N_3775);
and U6229 (N_6229,N_4611,N_3889);
nor U6230 (N_6230,N_4183,N_4601);
nor U6231 (N_6231,N_4580,N_4962);
or U6232 (N_6232,N_4917,N_4807);
xor U6233 (N_6233,N_4384,N_4245);
xnor U6234 (N_6234,N_3935,N_4877);
nor U6235 (N_6235,N_4843,N_4414);
xnor U6236 (N_6236,N_4255,N_4222);
xor U6237 (N_6237,N_4149,N_4982);
or U6238 (N_6238,N_4489,N_3959);
nand U6239 (N_6239,N_3801,N_4238);
and U6240 (N_6240,N_4281,N_4880);
or U6241 (N_6241,N_3958,N_3932);
xor U6242 (N_6242,N_4131,N_4129);
xor U6243 (N_6243,N_4761,N_4993);
nand U6244 (N_6244,N_4091,N_4274);
or U6245 (N_6245,N_4315,N_3954);
nor U6246 (N_6246,N_4993,N_4653);
xnor U6247 (N_6247,N_3869,N_4992);
and U6248 (N_6248,N_4745,N_3823);
or U6249 (N_6249,N_4066,N_4655);
xor U6250 (N_6250,N_5510,N_6061);
nor U6251 (N_6251,N_5305,N_5969);
and U6252 (N_6252,N_5046,N_5007);
nor U6253 (N_6253,N_5430,N_5115);
and U6254 (N_6254,N_5754,N_5935);
and U6255 (N_6255,N_5348,N_5696);
xor U6256 (N_6256,N_5050,N_5592);
and U6257 (N_6257,N_5474,N_6175);
nor U6258 (N_6258,N_6108,N_5763);
nor U6259 (N_6259,N_5166,N_5365);
or U6260 (N_6260,N_6031,N_5715);
nand U6261 (N_6261,N_5039,N_5880);
nor U6262 (N_6262,N_5630,N_5083);
and U6263 (N_6263,N_5746,N_5629);
nand U6264 (N_6264,N_5383,N_5875);
nor U6265 (N_6265,N_5570,N_6132);
nor U6266 (N_6266,N_6066,N_6243);
xor U6267 (N_6267,N_5994,N_5183);
xnor U6268 (N_6268,N_6159,N_5025);
nand U6269 (N_6269,N_5056,N_5834);
xnor U6270 (N_6270,N_6103,N_6017);
xor U6271 (N_6271,N_5968,N_6086);
nand U6272 (N_6272,N_6021,N_5739);
and U6273 (N_6273,N_5605,N_5463);
nor U6274 (N_6274,N_5472,N_6213);
nor U6275 (N_6275,N_5084,N_5883);
or U6276 (N_6276,N_5732,N_5977);
nor U6277 (N_6277,N_6200,N_5077);
or U6278 (N_6278,N_5061,N_6166);
and U6279 (N_6279,N_5639,N_6116);
xor U6280 (N_6280,N_5210,N_5176);
nor U6281 (N_6281,N_5721,N_6208);
or U6282 (N_6282,N_5281,N_5042);
or U6283 (N_6283,N_5964,N_5819);
nor U6284 (N_6284,N_6245,N_5030);
nor U6285 (N_6285,N_5989,N_6045);
xor U6286 (N_6286,N_5979,N_5691);
or U6287 (N_6287,N_5829,N_5925);
and U6288 (N_6288,N_5847,N_6240);
or U6289 (N_6289,N_5349,N_5985);
xor U6290 (N_6290,N_5566,N_5098);
nand U6291 (N_6291,N_5535,N_5613);
xnor U6292 (N_6292,N_5826,N_5102);
or U6293 (N_6293,N_5353,N_5646);
and U6294 (N_6294,N_5720,N_5653);
nor U6295 (N_6295,N_5218,N_6225);
nor U6296 (N_6296,N_5800,N_5422);
and U6297 (N_6297,N_5869,N_5892);
nor U6298 (N_6298,N_5788,N_5745);
or U6299 (N_6299,N_5725,N_6034);
nor U6300 (N_6300,N_6207,N_6079);
xor U6301 (N_6301,N_5101,N_5870);
nand U6302 (N_6302,N_5648,N_5481);
nand U6303 (N_6303,N_5297,N_5329);
and U6304 (N_6304,N_5433,N_5685);
nand U6305 (N_6305,N_6222,N_5934);
or U6306 (N_6306,N_5560,N_5151);
nand U6307 (N_6307,N_5505,N_5719);
or U6308 (N_6308,N_6075,N_6076);
nor U6309 (N_6309,N_5947,N_5212);
nor U6310 (N_6310,N_5354,N_5769);
nor U6311 (N_6311,N_5864,N_5246);
xor U6312 (N_6312,N_5206,N_5181);
or U6313 (N_6313,N_5375,N_5073);
or U6314 (N_6314,N_5108,N_6133);
or U6315 (N_6315,N_6105,N_5028);
or U6316 (N_6316,N_5758,N_5309);
nor U6317 (N_6317,N_5252,N_5086);
xor U6318 (N_6318,N_5737,N_5120);
and U6319 (N_6319,N_6053,N_5448);
or U6320 (N_6320,N_6134,N_5960);
nor U6321 (N_6321,N_6101,N_6139);
and U6322 (N_6322,N_5052,N_5397);
nor U6323 (N_6323,N_5045,N_6118);
and U6324 (N_6324,N_5043,N_5150);
and U6325 (N_6325,N_6064,N_5274);
or U6326 (N_6326,N_5138,N_5285);
or U6327 (N_6327,N_5756,N_5453);
nand U6328 (N_6328,N_6135,N_6177);
and U6329 (N_6329,N_5584,N_5621);
nor U6330 (N_6330,N_6089,N_5014);
and U6331 (N_6331,N_5016,N_5018);
and U6332 (N_6332,N_5517,N_5438);
nand U6333 (N_6333,N_5263,N_5440);
nand U6334 (N_6334,N_5807,N_5502);
or U6335 (N_6335,N_5233,N_5713);
xnor U6336 (N_6336,N_5228,N_5187);
nor U6337 (N_6337,N_5011,N_6220);
or U6338 (N_6338,N_6150,N_5953);
and U6339 (N_6339,N_5997,N_5972);
and U6340 (N_6340,N_5905,N_5067);
nand U6341 (N_6341,N_5147,N_5189);
and U6342 (N_6342,N_5109,N_5303);
and U6343 (N_6343,N_6148,N_6239);
nand U6344 (N_6344,N_5603,N_5919);
or U6345 (N_6345,N_5716,N_5874);
xor U6346 (N_6346,N_5160,N_5265);
and U6347 (N_6347,N_5678,N_5139);
and U6348 (N_6348,N_5550,N_5359);
or U6349 (N_6349,N_5226,N_5373);
nor U6350 (N_6350,N_5565,N_6221);
xnor U6351 (N_6351,N_5827,N_5385);
or U6352 (N_6352,N_5786,N_5457);
and U6353 (N_6353,N_6090,N_5488);
or U6354 (N_6354,N_5848,N_6039);
and U6355 (N_6355,N_5902,N_5232);
xor U6356 (N_6356,N_5024,N_5482);
nand U6357 (N_6357,N_5624,N_5171);
nor U6358 (N_6358,N_5106,N_5300);
xnor U6359 (N_6359,N_5227,N_5573);
or U6360 (N_6360,N_5751,N_5406);
or U6361 (N_6361,N_6110,N_5749);
nand U6362 (N_6362,N_5319,N_6165);
or U6363 (N_6363,N_5454,N_5118);
xor U6364 (N_6364,N_5296,N_6085);
nor U6365 (N_6365,N_5292,N_6181);
xnor U6366 (N_6366,N_6044,N_5220);
or U6367 (N_6367,N_5930,N_5967);
xor U6368 (N_6368,N_5248,N_5586);
nor U6369 (N_6369,N_6130,N_6215);
or U6370 (N_6370,N_5891,N_5242);
and U6371 (N_6371,N_5814,N_5623);
xor U6372 (N_6372,N_5524,N_6151);
nand U6373 (N_6373,N_5669,N_6125);
or U6374 (N_6374,N_5954,N_5062);
or U6375 (N_6375,N_6174,N_5950);
nand U6376 (N_6376,N_5031,N_5003);
or U6377 (N_6377,N_5583,N_5983);
nor U6378 (N_6378,N_5620,N_5127);
or U6379 (N_6379,N_5339,N_6147);
nor U6380 (N_6380,N_5866,N_5331);
and U6381 (N_6381,N_5378,N_5790);
nor U6382 (N_6382,N_6160,N_5033);
and U6383 (N_6383,N_5146,N_6205);
nand U6384 (N_6384,N_5889,N_5497);
nor U6385 (N_6385,N_5679,N_5940);
and U6386 (N_6386,N_5165,N_5390);
nand U6387 (N_6387,N_5890,N_5149);
nor U6388 (N_6388,N_5405,N_6106);
nor U6389 (N_6389,N_5501,N_6069);
nor U6390 (N_6390,N_5671,N_5134);
or U6391 (N_6391,N_5254,N_5662);
nand U6392 (N_6392,N_6102,N_5652);
nor U6393 (N_6393,N_6027,N_5230);
and U6394 (N_6394,N_5010,N_5901);
nor U6395 (N_6395,N_6009,N_5267);
nand U6396 (N_6396,N_5626,N_6236);
or U6397 (N_6397,N_5882,N_5424);
xor U6398 (N_6398,N_5765,N_5377);
or U6399 (N_6399,N_5304,N_5493);
and U6400 (N_6400,N_5207,N_5002);
or U6401 (N_6401,N_5247,N_5355);
xnor U6402 (N_6402,N_6188,N_6144);
and U6403 (N_6403,N_5873,N_5104);
xnor U6404 (N_6404,N_5742,N_5490);
or U6405 (N_6405,N_5116,N_6008);
nand U6406 (N_6406,N_5724,N_6248);
xnor U6407 (N_6407,N_6104,N_5794);
or U6408 (N_6408,N_6016,N_5809);
nor U6409 (N_6409,N_5484,N_5789);
nor U6410 (N_6410,N_6227,N_5468);
xnor U6411 (N_6411,N_5401,N_5216);
and U6412 (N_6412,N_5854,N_6001);
xnor U6413 (N_6413,N_5782,N_5687);
xnor U6414 (N_6414,N_5625,N_5519);
or U6415 (N_6415,N_5633,N_5852);
xnor U6416 (N_6416,N_5838,N_5879);
or U6417 (N_6417,N_5812,N_5193);
nand U6418 (N_6418,N_6117,N_5973);
or U6419 (N_6419,N_5436,N_5069);
or U6420 (N_6420,N_6142,N_5649);
and U6421 (N_6421,N_5221,N_5013);
nor U6422 (N_6422,N_6242,N_5409);
nor U6423 (N_6423,N_5970,N_6238);
or U6424 (N_6424,N_6019,N_5429);
or U6425 (N_6425,N_5412,N_5148);
or U6426 (N_6426,N_6022,N_5860);
xor U6427 (N_6427,N_5072,N_5551);
nor U6428 (N_6428,N_5418,N_5461);
xor U6429 (N_6429,N_5956,N_5264);
xor U6430 (N_6430,N_5037,N_5078);
and U6431 (N_6431,N_5403,N_5740);
or U6432 (N_6432,N_5437,N_6097);
and U6433 (N_6433,N_5387,N_5998);
or U6434 (N_6434,N_5219,N_5175);
nand U6435 (N_6435,N_6137,N_5236);
xnor U6436 (N_6436,N_5100,N_5299);
and U6437 (N_6437,N_5689,N_5546);
xor U6438 (N_6438,N_5734,N_5656);
nor U6439 (N_6439,N_6155,N_5755);
and U6440 (N_6440,N_5993,N_6235);
and U6441 (N_6441,N_5558,N_5974);
nand U6442 (N_6442,N_5709,N_5244);
nor U6443 (N_6443,N_6011,N_5702);
nand U6444 (N_6444,N_5926,N_5540);
and U6445 (N_6445,N_5295,N_5795);
nand U6446 (N_6446,N_5032,N_5130);
and U6447 (N_6447,N_5810,N_5371);
nor U6448 (N_6448,N_5898,N_5347);
nand U6449 (N_6449,N_5664,N_5279);
and U6450 (N_6450,N_5076,N_5728);
nand U6451 (N_6451,N_6083,N_5167);
xnor U6452 (N_6452,N_5817,N_5133);
nand U6453 (N_6453,N_6184,N_5632);
and U6454 (N_6454,N_5180,N_6054);
nor U6455 (N_6455,N_5485,N_5744);
or U6456 (N_6456,N_5526,N_5512);
nor U6457 (N_6457,N_5094,N_5628);
nor U6458 (N_6458,N_5562,N_5311);
nand U6459 (N_6459,N_5743,N_6120);
nor U6460 (N_6460,N_5420,N_5272);
nor U6461 (N_6461,N_5386,N_5017);
nand U6462 (N_6462,N_5352,N_5301);
nand U6463 (N_6463,N_6041,N_5867);
nand U6464 (N_6464,N_5486,N_5912);
xor U6465 (N_6465,N_6247,N_5853);
nand U6466 (N_6466,N_5465,N_5174);
nor U6467 (N_6467,N_6096,N_5491);
xnor U6468 (N_6468,N_5792,N_6173);
nand U6469 (N_6469,N_6206,N_5785);
nand U6470 (N_6470,N_5021,N_5381);
nor U6471 (N_6471,N_5239,N_5340);
nand U6472 (N_6472,N_5700,N_5135);
nor U6473 (N_6473,N_6229,N_5277);
and U6474 (N_6474,N_5258,N_5774);
and U6475 (N_6475,N_5389,N_5394);
nand U6476 (N_6476,N_5757,N_5326);
xor U6477 (N_6477,N_5170,N_6036);
nor U6478 (N_6478,N_5040,N_5241);
or U6479 (N_6479,N_6025,N_5576);
nor U6480 (N_6480,N_5411,N_5255);
or U6481 (N_6481,N_5999,N_5136);
and U6482 (N_6482,N_5775,N_6124);
nor U6483 (N_6483,N_5975,N_5538);
and U6484 (N_6484,N_5356,N_6187);
or U6485 (N_6485,N_5959,N_5446);
or U6486 (N_6486,N_6024,N_5152);
nor U6487 (N_6487,N_6204,N_5943);
or U6488 (N_6488,N_5640,N_5682);
or U6489 (N_6489,N_5182,N_5107);
xnor U6490 (N_6490,N_5521,N_5958);
nand U6491 (N_6491,N_5419,N_5191);
and U6492 (N_6492,N_5609,N_5222);
nand U6493 (N_6493,N_5396,N_6051);
nor U6494 (N_6494,N_5400,N_5198);
or U6495 (N_6495,N_5055,N_6199);
nand U6496 (N_6496,N_6163,N_5618);
nand U6497 (N_6497,N_5747,N_5859);
and U6498 (N_6498,N_5172,N_5990);
nand U6499 (N_6499,N_6091,N_5851);
nand U6500 (N_6500,N_5726,N_5336);
and U6501 (N_6501,N_5752,N_5657);
xor U6502 (N_6502,N_5494,N_5200);
or U6503 (N_6503,N_5766,N_6129);
and U6504 (N_6504,N_5784,N_5284);
or U6505 (N_6505,N_5345,N_5578);
xnor U6506 (N_6506,N_5350,N_5850);
nand U6507 (N_6507,N_6058,N_5435);
nand U6508 (N_6508,N_5112,N_5333);
nand U6509 (N_6509,N_5840,N_6088);
xor U6510 (N_6510,N_5856,N_5557);
or U6511 (N_6511,N_5690,N_5423);
nor U6512 (N_6512,N_5861,N_5748);
xor U6513 (N_6513,N_6186,N_6111);
nand U6514 (N_6514,N_6196,N_6094);
and U6515 (N_6515,N_5450,N_5213);
nor U6516 (N_6516,N_5986,N_5780);
and U6517 (N_6517,N_5799,N_5910);
xor U6518 (N_6518,N_5103,N_6081);
nor U6519 (N_6519,N_5545,N_5665);
xnor U6520 (N_6520,N_5129,N_5820);
nor U6521 (N_6521,N_6212,N_5644);
or U6522 (N_6522,N_5132,N_5320);
and U6523 (N_6523,N_5384,N_5289);
or U6524 (N_6524,N_5572,N_5865);
nor U6525 (N_6525,N_6140,N_5527);
nand U6526 (N_6526,N_5821,N_5314);
or U6527 (N_6527,N_6152,N_5862);
or U6528 (N_6528,N_5514,N_5057);
or U6529 (N_6529,N_5642,N_5666);
xnor U6530 (N_6530,N_5949,N_5523);
and U6531 (N_6531,N_5895,N_6010);
and U6532 (N_6532,N_5868,N_6000);
or U6533 (N_6533,N_6068,N_5416);
nand U6534 (N_6534,N_6003,N_5730);
or U6535 (N_6535,N_5179,N_5262);
nor U6536 (N_6536,N_5932,N_5841);
nand U6537 (N_6537,N_5273,N_6168);
or U6538 (N_6538,N_5580,N_5503);
nand U6539 (N_6539,N_5399,N_5981);
or U6540 (N_6540,N_5564,N_5637);
nand U6541 (N_6541,N_5119,N_5325);
xnor U6542 (N_6542,N_5881,N_5855);
nand U6543 (N_6543,N_5466,N_5563);
and U6544 (N_6544,N_6107,N_6219);
or U6545 (N_6545,N_5068,N_5845);
and U6546 (N_6546,N_5005,N_5408);
and U6547 (N_6547,N_5995,N_5020);
nand U6548 (N_6548,N_5802,N_5761);
or U6549 (N_6549,N_5708,N_5894);
nor U6550 (N_6550,N_5773,N_5522);
or U6551 (N_6551,N_5579,N_5434);
nor U6552 (N_6552,N_5729,N_6121);
nand U6553 (N_6553,N_5805,N_5590);
or U6554 (N_6554,N_5245,N_5984);
or U6555 (N_6555,N_5278,N_5909);
xor U6556 (N_6556,N_5695,N_5250);
and U6557 (N_6557,N_6141,N_5796);
xor U6558 (N_6558,N_5920,N_5508);
xor U6559 (N_6559,N_5287,N_5951);
xnor U6560 (N_6560,N_5798,N_5651);
and U6561 (N_6561,N_5914,N_5158);
nand U6562 (N_6562,N_5587,N_5929);
nor U6563 (N_6563,N_5699,N_5019);
xnor U6564 (N_6564,N_5051,N_5924);
or U6565 (N_6565,N_6015,N_5323);
nor U6566 (N_6566,N_5759,N_6071);
nor U6567 (N_6567,N_5598,N_6042);
or U6568 (N_6568,N_5904,N_6194);
xnor U6569 (N_6569,N_6100,N_6072);
and U6570 (N_6570,N_5617,N_6007);
nand U6571 (N_6571,N_5878,N_5647);
or U6572 (N_6572,N_5568,N_5338);
xnor U6573 (N_6573,N_5459,N_5760);
or U6574 (N_6574,N_6084,N_5684);
and U6575 (N_6575,N_5770,N_6059);
nand U6576 (N_6576,N_5328,N_5513);
nor U6577 (N_6577,N_5066,N_5082);
and U6578 (N_6578,N_5631,N_5477);
or U6579 (N_6579,N_5487,N_5828);
nand U6580 (N_6580,N_5034,N_5074);
or U6581 (N_6581,N_5741,N_5122);
or U6582 (N_6582,N_6033,N_6078);
or U6583 (N_6583,N_5916,N_6123);
or U6584 (N_6584,N_5393,N_6180);
nand U6585 (N_6585,N_5458,N_5507);
or U6586 (N_6586,N_5164,N_5608);
and U6587 (N_6587,N_5818,N_5395);
or U6588 (N_6588,N_6195,N_6037);
xor U6589 (N_6589,N_5806,N_5388);
xnor U6590 (N_6590,N_5616,N_5288);
or U6591 (N_6591,N_5768,N_6127);
or U6592 (N_6592,N_5332,N_6190);
or U6593 (N_6593,N_6201,N_5543);
nor U6594 (N_6594,N_5196,N_5641);
nor U6595 (N_6595,N_5065,N_5987);
xor U6596 (N_6596,N_5214,N_6126);
or U6597 (N_6597,N_6035,N_5643);
nor U6598 (N_6598,N_5306,N_5871);
nor U6599 (N_6599,N_5302,N_6246);
and U6600 (N_6600,N_5079,N_5939);
nor U6601 (N_6601,N_5425,N_5224);
or U6602 (N_6602,N_5936,N_5442);
nand U6603 (N_6603,N_5893,N_6014);
nor U6604 (N_6604,N_5075,N_5733);
xnor U6605 (N_6605,N_5683,N_5750);
nand U6606 (N_6606,N_6136,N_5091);
and U6607 (N_6607,N_5900,N_5211);
and U6608 (N_6608,N_5815,N_5313);
and U6609 (N_6609,N_5908,N_5374);
and U6610 (N_6610,N_6145,N_5597);
and U6611 (N_6611,N_5753,N_5645);
or U6612 (N_6612,N_6029,N_5449);
and U6613 (N_6613,N_6048,N_5811);
nor U6614 (N_6614,N_5469,N_5735);
or U6615 (N_6615,N_5764,N_5452);
nor U6616 (N_6616,N_6149,N_5367);
nor U6617 (N_6617,N_5884,N_5711);
nor U6618 (N_6618,N_5499,N_5823);
nor U6619 (N_6619,N_5363,N_5334);
nor U6620 (N_6620,N_6032,N_5492);
nor U6621 (N_6621,N_5439,N_5677);
or U6622 (N_6622,N_5121,N_6223);
xor U6623 (N_6623,N_5697,N_5942);
xnor U6624 (N_6624,N_5161,N_5188);
and U6625 (N_6625,N_5053,N_5813);
nor U6626 (N_6626,N_5269,N_5154);
nand U6627 (N_6627,N_5567,N_5366);
nor U6628 (N_6628,N_5081,N_5516);
nor U6629 (N_6629,N_5532,N_5594);
nand U6630 (N_6630,N_5688,N_5447);
xor U6631 (N_6631,N_5324,N_5364);
and U6632 (N_6632,N_5803,N_5346);
and U6633 (N_6633,N_5208,N_5614);
nor U6634 (N_6634,N_6154,N_5680);
nor U6635 (N_6635,N_5585,N_5173);
xor U6636 (N_6636,N_5602,N_6046);
nand U6637 (N_6637,N_5610,N_6018);
or U6638 (N_6638,N_5681,N_6230);
nor U6639 (N_6639,N_5982,N_5322);
xor U6640 (N_6640,N_5351,N_6237);
nand U6641 (N_6641,N_5703,N_5293);
nor U6642 (N_6642,N_5080,N_5791);
nor U6643 (N_6643,N_5256,N_5515);
nand U6644 (N_6644,N_6119,N_5004);
or U6645 (N_6645,N_6002,N_5635);
nor U6646 (N_6646,N_5125,N_5506);
nor U6647 (N_6647,N_5670,N_5298);
or U6648 (N_6648,N_5674,N_5470);
nor U6649 (N_6649,N_5195,N_5822);
xor U6650 (N_6650,N_5548,N_5672);
or U6651 (N_6651,N_5111,N_5661);
nand U6652 (N_6652,N_5842,N_5243);
nor U6653 (N_6653,N_5554,N_5237);
or U6654 (N_6654,N_6052,N_5321);
nor U6655 (N_6655,N_5738,N_5952);
nand U6656 (N_6656,N_6170,N_5382);
nor U6657 (N_6657,N_5194,N_5599);
or U6658 (N_6658,N_5318,N_5344);
and U6659 (N_6659,N_5559,N_5271);
nor U6660 (N_6660,N_6060,N_5105);
and U6661 (N_6661,N_5140,N_6115);
or U6662 (N_6662,N_5876,N_5783);
and U6663 (N_6663,N_6198,N_5342);
or U6664 (N_6664,N_5906,N_5145);
and U6665 (N_6665,N_5204,N_5962);
nor U6666 (N_6666,N_6030,N_5574);
xnor U6667 (N_6667,N_5225,N_5824);
and U6668 (N_6668,N_6210,N_5676);
nand U6669 (N_6669,N_5996,N_6109);
nand U6670 (N_6670,N_6006,N_5009);
xor U6671 (N_6671,N_5312,N_6211);
nand U6672 (N_6672,N_5965,N_5542);
and U6673 (N_6673,N_6241,N_5938);
or U6674 (N_6674,N_5736,N_6162);
nand U6675 (N_6675,N_5727,N_5992);
nor U6676 (N_6676,N_5192,N_5456);
nor U6677 (N_6677,N_5015,N_5831);
and U6678 (N_6678,N_6047,N_5928);
and U6679 (N_6679,N_5663,N_5622);
xnor U6680 (N_6680,N_5261,N_6249);
xnor U6681 (N_6681,N_5555,N_5008);
nor U6682 (N_6682,N_6050,N_5012);
nor U6683 (N_6683,N_5327,N_6114);
nor U6684 (N_6684,N_5706,N_5591);
or U6685 (N_6685,N_5520,N_6073);
and U6686 (N_6686,N_5832,N_6112);
nand U6687 (N_6687,N_5054,N_5308);
and U6688 (N_6688,N_5128,N_5923);
xnor U6689 (N_6689,N_5144,N_5064);
or U6690 (N_6690,N_5899,N_5601);
nor U6691 (N_6691,N_5153,N_5070);
xor U6692 (N_6692,N_5544,N_6028);
and U6693 (N_6693,N_5337,N_5692);
nor U6694 (N_6694,N_5185,N_5911);
xnor U6695 (N_6695,N_6005,N_5650);
nand U6696 (N_6696,N_5445,N_6067);
nand U6697 (N_6697,N_5071,N_6138);
xnor U6698 (N_6698,N_5718,N_5604);
and U6699 (N_6699,N_5240,N_5537);
nor U6700 (N_6700,N_5223,N_6233);
nor U6701 (N_6701,N_6234,N_5529);
xnor U6702 (N_6702,N_5467,N_5931);
xnor U6703 (N_6703,N_5460,N_5229);
and U6704 (N_6704,N_6063,N_5606);
and U6705 (N_6705,N_5443,N_6156);
xnor U6706 (N_6706,N_5260,N_6128);
or U6707 (N_6707,N_5159,N_6077);
xnor U6708 (N_6708,N_5897,N_6146);
or U6709 (N_6709,N_5498,N_5777);
and U6710 (N_6710,N_5957,N_5552);
nand U6711 (N_6711,N_5169,N_5801);
nand U6712 (N_6712,N_6228,N_6043);
and U6713 (N_6713,N_5413,N_5097);
nor U6714 (N_6714,N_5843,N_5376);
xnor U6715 (N_6715,N_5705,N_5907);
or U6716 (N_6716,N_5571,N_5858);
nand U6717 (N_6717,N_5533,N_5600);
nor U6718 (N_6718,N_5280,N_5509);
nand U6719 (N_6719,N_5582,N_5634);
xor U6720 (N_6720,N_5528,N_6070);
nor U6721 (N_6721,N_5414,N_5142);
and U6722 (N_6722,N_6012,N_5155);
and U6723 (N_6723,N_5534,N_6191);
nor U6724 (N_6724,N_6062,N_5536);
or U6725 (N_6725,N_5589,N_5668);
nor U6726 (N_6726,N_5036,N_5872);
nand U6727 (N_6727,N_5451,N_5955);
or U6728 (N_6728,N_5686,N_5844);
and U6729 (N_6729,N_5978,N_5483);
and U6730 (N_6730,N_5698,N_6218);
xor U6731 (N_6731,N_5804,N_5561);
nand U6732 (N_6732,N_5933,N_5787);
nor U6733 (N_6733,N_5063,N_6157);
xor U6734 (N_6734,N_5693,N_6158);
or U6735 (N_6735,N_6065,N_5123);
xor U6736 (N_6736,N_5569,N_5205);
and U6737 (N_6737,N_6182,N_5944);
nor U6738 (N_6738,N_6057,N_6171);
nand U6739 (N_6739,N_6153,N_5235);
nor U6740 (N_6740,N_5178,N_5886);
nand U6741 (N_6741,N_5547,N_5275);
nor U6742 (N_6742,N_5163,N_6176);
nor U6743 (N_6743,N_5310,N_5588);
xnor U6744 (N_6744,N_5945,N_5918);
xnor U6745 (N_6745,N_6082,N_6202);
xnor U6746 (N_6746,N_5156,N_5251);
or U6747 (N_6747,N_5088,N_5391);
xor U6748 (N_6748,N_5941,N_5023);
nand U6749 (N_6749,N_5917,N_5575);
xnor U6750 (N_6750,N_5026,N_6214);
nor U6751 (N_6751,N_5887,N_5511);
nor U6752 (N_6752,N_5636,N_5476);
nor U6753 (N_6753,N_5421,N_5471);
or U6754 (N_6754,N_5863,N_5549);
and U6755 (N_6755,N_5479,N_5291);
or U6756 (N_6756,N_5504,N_5707);
or U6757 (N_6757,N_5369,N_5480);
nor U6758 (N_6758,N_5410,N_5141);
and U6759 (N_6759,N_6164,N_5307);
nand U6760 (N_6760,N_5268,N_6193);
xnor U6761 (N_6761,N_5215,N_5849);
nor U6762 (N_6762,N_5593,N_5963);
nor U6763 (N_6763,N_5722,N_5095);
or U6764 (N_6764,N_6095,N_5290);
and U6765 (N_6765,N_5489,N_5714);
nand U6766 (N_6766,N_6040,N_5627);
nor U6767 (N_6767,N_5238,N_5276);
nor U6768 (N_6768,N_5922,N_5462);
or U6769 (N_6769,N_5475,N_5317);
xor U6770 (N_6770,N_5360,N_5368);
nand U6771 (N_6771,N_5335,N_5673);
nor U6772 (N_6772,N_5444,N_5048);
xnor U6773 (N_6773,N_5379,N_5157);
nand U6774 (N_6774,N_6161,N_5776);
nand U6775 (N_6775,N_5991,N_5234);
xor U6776 (N_6776,N_6172,N_6023);
xor U6777 (N_6777,N_5044,N_6131);
nor U6778 (N_6778,N_5049,N_5294);
and U6779 (N_6779,N_5370,N_5797);
nand U6780 (N_6780,N_6185,N_5190);
nand U6781 (N_6781,N_5595,N_5358);
xnor U6782 (N_6782,N_5553,N_5428);
nor U6783 (N_6783,N_5427,N_6092);
nor U6784 (N_6784,N_6178,N_5833);
nand U6785 (N_6785,N_6049,N_6197);
nand U6786 (N_6786,N_5638,N_5404);
nor U6787 (N_6787,N_5779,N_5825);
xnor U6788 (N_6788,N_5846,N_5808);
nand U6789 (N_6789,N_5201,N_5837);
and U6790 (N_6790,N_5885,N_5704);
and U6791 (N_6791,N_5000,N_5060);
nand U6792 (N_6792,N_5341,N_5380);
and U6793 (N_6793,N_6203,N_6179);
or U6794 (N_6794,N_5114,N_5432);
or U6795 (N_6795,N_5525,N_5092);
or U6796 (N_6796,N_5249,N_5266);
or U6797 (N_6797,N_5431,N_5658);
nand U6798 (N_6798,N_5772,N_5316);
xnor U6799 (N_6799,N_5168,N_5927);
xnor U6800 (N_6800,N_5980,N_5330);
xor U6801 (N_6801,N_5857,N_5362);
nor U6802 (N_6802,N_5209,N_5966);
nor U6803 (N_6803,N_6093,N_5717);
xnor U6804 (N_6804,N_5282,N_5946);
and U6805 (N_6805,N_5202,N_5478);
nand U6806 (N_6806,N_5830,N_5162);
xnor U6807 (N_6807,N_5143,N_5217);
or U6808 (N_6808,N_5441,N_6143);
nand U6809 (N_6809,N_6244,N_6224);
xor U6810 (N_6810,N_5022,N_5001);
or U6811 (N_6811,N_5539,N_5113);
nor U6812 (N_6812,N_6169,N_5701);
nand U6813 (N_6813,N_5398,N_6113);
or U6814 (N_6814,N_6080,N_6026);
nor U6815 (N_6815,N_5315,N_5654);
and U6816 (N_6816,N_5619,N_5793);
nor U6817 (N_6817,N_5877,N_6231);
or U6818 (N_6818,N_6074,N_5402);
xor U6819 (N_6819,N_5581,N_6004);
or U6820 (N_6820,N_5126,N_5027);
nand U6821 (N_6821,N_5518,N_5577);
xor U6822 (N_6822,N_5203,N_5231);
xor U6823 (N_6823,N_5464,N_5976);
nand U6824 (N_6824,N_5655,N_5710);
nand U6825 (N_6825,N_5343,N_6055);
nor U6826 (N_6826,N_5357,N_5035);
nor U6827 (N_6827,N_5415,N_5948);
nor U6828 (N_6828,N_6209,N_5530);
or U6829 (N_6829,N_5731,N_5455);
nor U6830 (N_6830,N_6013,N_5372);
and U6831 (N_6831,N_5270,N_6216);
or U6832 (N_6832,N_5607,N_5835);
and U6833 (N_6833,N_5058,N_5903);
nand U6834 (N_6834,N_5778,N_5541);
nor U6835 (N_6835,N_6189,N_5417);
xnor U6836 (N_6836,N_5762,N_5667);
nor U6837 (N_6837,N_5177,N_6038);
xor U6838 (N_6838,N_5093,N_5283);
xor U6839 (N_6839,N_5781,N_5186);
nor U6840 (N_6840,N_5771,N_5767);
xnor U6841 (N_6841,N_5988,N_5712);
and U6842 (N_6842,N_5059,N_5047);
nand U6843 (N_6843,N_5500,N_5836);
nor U6844 (N_6844,N_5694,N_5921);
or U6845 (N_6845,N_5257,N_6098);
and U6846 (N_6846,N_5723,N_5426);
xor U6847 (N_6847,N_6122,N_5896);
nor U6848 (N_6848,N_5041,N_5615);
or U6849 (N_6849,N_6232,N_5816);
xor U6850 (N_6850,N_5888,N_6020);
and U6851 (N_6851,N_5184,N_5496);
xor U6852 (N_6852,N_5937,N_5473);
or U6853 (N_6853,N_6087,N_5556);
xnor U6854 (N_6854,N_5096,N_5839);
and U6855 (N_6855,N_5006,N_6183);
xor U6856 (N_6856,N_5961,N_5913);
or U6857 (N_6857,N_5611,N_5253);
nor U6858 (N_6858,N_5971,N_5087);
nand U6859 (N_6859,N_5392,N_5259);
and U6860 (N_6860,N_5124,N_6192);
and U6861 (N_6861,N_5137,N_5531);
xor U6862 (N_6862,N_6056,N_5596);
or U6863 (N_6863,N_6099,N_5612);
nor U6864 (N_6864,N_5089,N_5199);
and U6865 (N_6865,N_5131,N_5407);
nand U6866 (N_6866,N_6167,N_5286);
and U6867 (N_6867,N_5110,N_5659);
and U6868 (N_6868,N_5495,N_5197);
xnor U6869 (N_6869,N_5660,N_5915);
and U6870 (N_6870,N_5361,N_6217);
nand U6871 (N_6871,N_5090,N_5117);
xor U6872 (N_6872,N_6226,N_5099);
nor U6873 (N_6873,N_5029,N_5038);
nor U6874 (N_6874,N_5085,N_5675);
and U6875 (N_6875,N_5513,N_5002);
nor U6876 (N_6876,N_6048,N_5523);
and U6877 (N_6877,N_5637,N_5773);
or U6878 (N_6878,N_5902,N_5708);
nand U6879 (N_6879,N_5125,N_5992);
or U6880 (N_6880,N_5610,N_5091);
or U6881 (N_6881,N_5334,N_5056);
nand U6882 (N_6882,N_5768,N_5646);
nand U6883 (N_6883,N_5647,N_5332);
nand U6884 (N_6884,N_5806,N_5668);
nor U6885 (N_6885,N_6130,N_5020);
nand U6886 (N_6886,N_5592,N_5086);
nand U6887 (N_6887,N_5048,N_5416);
or U6888 (N_6888,N_5401,N_5485);
xor U6889 (N_6889,N_5001,N_5198);
nand U6890 (N_6890,N_5876,N_5433);
xor U6891 (N_6891,N_5487,N_5787);
or U6892 (N_6892,N_5211,N_6042);
or U6893 (N_6893,N_5859,N_6042);
nand U6894 (N_6894,N_5479,N_5175);
nand U6895 (N_6895,N_5905,N_5646);
or U6896 (N_6896,N_5017,N_5828);
or U6897 (N_6897,N_5165,N_5554);
or U6898 (N_6898,N_6175,N_5255);
and U6899 (N_6899,N_5991,N_6146);
or U6900 (N_6900,N_5228,N_5706);
xor U6901 (N_6901,N_5183,N_6160);
and U6902 (N_6902,N_5260,N_5688);
or U6903 (N_6903,N_5730,N_5004);
nor U6904 (N_6904,N_6138,N_5262);
xor U6905 (N_6905,N_6196,N_5700);
and U6906 (N_6906,N_5660,N_6110);
nand U6907 (N_6907,N_5915,N_5824);
and U6908 (N_6908,N_6063,N_5758);
xor U6909 (N_6909,N_5215,N_5320);
or U6910 (N_6910,N_5750,N_5345);
xor U6911 (N_6911,N_5989,N_5030);
nor U6912 (N_6912,N_5615,N_6203);
xor U6913 (N_6913,N_5418,N_5023);
xnor U6914 (N_6914,N_5485,N_5361);
xnor U6915 (N_6915,N_5207,N_5930);
and U6916 (N_6916,N_5768,N_5639);
or U6917 (N_6917,N_6134,N_5787);
xnor U6918 (N_6918,N_5309,N_5722);
and U6919 (N_6919,N_5388,N_6145);
and U6920 (N_6920,N_6227,N_5576);
nor U6921 (N_6921,N_6056,N_6065);
or U6922 (N_6922,N_5994,N_5339);
nor U6923 (N_6923,N_5462,N_5553);
and U6924 (N_6924,N_5962,N_5504);
or U6925 (N_6925,N_5357,N_5072);
xor U6926 (N_6926,N_5185,N_6177);
and U6927 (N_6927,N_5691,N_5950);
and U6928 (N_6928,N_6165,N_5821);
or U6929 (N_6929,N_5628,N_5450);
or U6930 (N_6930,N_5902,N_5115);
nor U6931 (N_6931,N_5345,N_6193);
nand U6932 (N_6932,N_5577,N_5650);
or U6933 (N_6933,N_5533,N_5708);
xor U6934 (N_6934,N_5410,N_6236);
nor U6935 (N_6935,N_6132,N_5144);
nor U6936 (N_6936,N_5834,N_5725);
nor U6937 (N_6937,N_5534,N_5091);
nand U6938 (N_6938,N_5340,N_5640);
nand U6939 (N_6939,N_5056,N_5108);
and U6940 (N_6940,N_5145,N_5300);
or U6941 (N_6941,N_5556,N_6211);
or U6942 (N_6942,N_6154,N_5032);
nor U6943 (N_6943,N_6138,N_5640);
xor U6944 (N_6944,N_5533,N_6224);
nand U6945 (N_6945,N_5004,N_5014);
xor U6946 (N_6946,N_5805,N_5473);
or U6947 (N_6947,N_5151,N_6162);
nand U6948 (N_6948,N_5811,N_5741);
nand U6949 (N_6949,N_6207,N_5104);
xnor U6950 (N_6950,N_5352,N_5003);
or U6951 (N_6951,N_5008,N_6054);
nor U6952 (N_6952,N_5403,N_5286);
nor U6953 (N_6953,N_6020,N_5236);
xnor U6954 (N_6954,N_6181,N_5551);
nand U6955 (N_6955,N_5020,N_5056);
or U6956 (N_6956,N_5662,N_5055);
or U6957 (N_6957,N_5445,N_5459);
nor U6958 (N_6958,N_5900,N_5282);
xor U6959 (N_6959,N_5557,N_5533);
or U6960 (N_6960,N_5263,N_5748);
or U6961 (N_6961,N_5298,N_5809);
nor U6962 (N_6962,N_5983,N_5699);
nor U6963 (N_6963,N_5309,N_5976);
and U6964 (N_6964,N_5312,N_5756);
nor U6965 (N_6965,N_5993,N_5707);
nand U6966 (N_6966,N_5042,N_5654);
xor U6967 (N_6967,N_5004,N_5994);
nand U6968 (N_6968,N_5527,N_5925);
nand U6969 (N_6969,N_5140,N_5358);
xor U6970 (N_6970,N_5111,N_6076);
nor U6971 (N_6971,N_5864,N_6007);
and U6972 (N_6972,N_5410,N_5322);
nor U6973 (N_6973,N_5617,N_5770);
nor U6974 (N_6974,N_6071,N_5735);
nand U6975 (N_6975,N_5607,N_5190);
and U6976 (N_6976,N_5449,N_5231);
nor U6977 (N_6977,N_5846,N_5537);
xor U6978 (N_6978,N_5301,N_5441);
nand U6979 (N_6979,N_5182,N_5020);
nand U6980 (N_6980,N_5389,N_5902);
and U6981 (N_6981,N_5507,N_5081);
xnor U6982 (N_6982,N_5529,N_5703);
nand U6983 (N_6983,N_6187,N_6049);
or U6984 (N_6984,N_5995,N_5635);
or U6985 (N_6985,N_6107,N_6113);
nor U6986 (N_6986,N_5001,N_5853);
nand U6987 (N_6987,N_5007,N_6029);
nor U6988 (N_6988,N_6086,N_5083);
or U6989 (N_6989,N_6125,N_5945);
and U6990 (N_6990,N_6238,N_6010);
nand U6991 (N_6991,N_5040,N_5601);
xor U6992 (N_6992,N_6201,N_5846);
xnor U6993 (N_6993,N_5631,N_5185);
nor U6994 (N_6994,N_5499,N_5261);
and U6995 (N_6995,N_5483,N_5154);
and U6996 (N_6996,N_5006,N_5658);
xor U6997 (N_6997,N_5636,N_5970);
and U6998 (N_6998,N_5210,N_6111);
or U6999 (N_6999,N_6037,N_5910);
and U7000 (N_7000,N_5488,N_5376);
or U7001 (N_7001,N_6144,N_6100);
nor U7002 (N_7002,N_5860,N_5706);
and U7003 (N_7003,N_5697,N_6049);
and U7004 (N_7004,N_5181,N_5494);
and U7005 (N_7005,N_5845,N_5576);
nor U7006 (N_7006,N_5972,N_5926);
nor U7007 (N_7007,N_5333,N_5659);
and U7008 (N_7008,N_5951,N_5657);
xor U7009 (N_7009,N_5822,N_5369);
or U7010 (N_7010,N_5366,N_5997);
or U7011 (N_7011,N_6170,N_5909);
and U7012 (N_7012,N_6042,N_5922);
nor U7013 (N_7013,N_5722,N_5834);
and U7014 (N_7014,N_5924,N_5262);
nand U7015 (N_7015,N_5121,N_5031);
nor U7016 (N_7016,N_5049,N_5513);
or U7017 (N_7017,N_5000,N_5937);
nor U7018 (N_7018,N_5662,N_5711);
nor U7019 (N_7019,N_5615,N_6218);
or U7020 (N_7020,N_5785,N_6148);
xor U7021 (N_7021,N_5613,N_6200);
nand U7022 (N_7022,N_5871,N_5576);
nor U7023 (N_7023,N_6151,N_5533);
xor U7024 (N_7024,N_5170,N_6186);
xor U7025 (N_7025,N_5720,N_5870);
nor U7026 (N_7026,N_5298,N_5093);
xnor U7027 (N_7027,N_5998,N_6039);
xnor U7028 (N_7028,N_6231,N_5674);
xor U7029 (N_7029,N_6014,N_5873);
xor U7030 (N_7030,N_5172,N_5435);
xor U7031 (N_7031,N_5693,N_5432);
or U7032 (N_7032,N_6063,N_5825);
or U7033 (N_7033,N_5001,N_5698);
and U7034 (N_7034,N_5416,N_5357);
or U7035 (N_7035,N_6175,N_6237);
nor U7036 (N_7036,N_5419,N_5661);
xor U7037 (N_7037,N_5865,N_5822);
nand U7038 (N_7038,N_5576,N_5637);
nor U7039 (N_7039,N_5245,N_5146);
or U7040 (N_7040,N_6151,N_5973);
or U7041 (N_7041,N_5966,N_5113);
nor U7042 (N_7042,N_5721,N_5533);
and U7043 (N_7043,N_5646,N_5462);
or U7044 (N_7044,N_5888,N_5915);
nor U7045 (N_7045,N_5166,N_5359);
and U7046 (N_7046,N_6215,N_5753);
and U7047 (N_7047,N_5817,N_6020);
or U7048 (N_7048,N_5169,N_5516);
nor U7049 (N_7049,N_5165,N_5693);
xor U7050 (N_7050,N_5275,N_5932);
or U7051 (N_7051,N_6146,N_5374);
nand U7052 (N_7052,N_5211,N_6203);
nand U7053 (N_7053,N_5125,N_5977);
and U7054 (N_7054,N_5155,N_5710);
xnor U7055 (N_7055,N_5747,N_6071);
nor U7056 (N_7056,N_6225,N_5741);
and U7057 (N_7057,N_5710,N_5369);
nor U7058 (N_7058,N_5635,N_5262);
nor U7059 (N_7059,N_5854,N_5162);
xnor U7060 (N_7060,N_5623,N_5492);
or U7061 (N_7061,N_5822,N_5109);
nor U7062 (N_7062,N_5557,N_5875);
xnor U7063 (N_7063,N_5637,N_5122);
xor U7064 (N_7064,N_5848,N_5612);
nor U7065 (N_7065,N_5779,N_5159);
or U7066 (N_7066,N_5886,N_5225);
xor U7067 (N_7067,N_6055,N_6231);
and U7068 (N_7068,N_6221,N_5190);
xnor U7069 (N_7069,N_5287,N_5345);
nand U7070 (N_7070,N_5960,N_5906);
nor U7071 (N_7071,N_6100,N_5681);
xor U7072 (N_7072,N_5872,N_5250);
nand U7073 (N_7073,N_5987,N_5609);
xor U7074 (N_7074,N_5519,N_6052);
nand U7075 (N_7075,N_5283,N_6119);
or U7076 (N_7076,N_6225,N_5926);
or U7077 (N_7077,N_5740,N_5491);
nor U7078 (N_7078,N_5017,N_5528);
or U7079 (N_7079,N_5953,N_5716);
nor U7080 (N_7080,N_5463,N_5900);
nor U7081 (N_7081,N_5722,N_5471);
nor U7082 (N_7082,N_5279,N_5190);
and U7083 (N_7083,N_5220,N_5722);
or U7084 (N_7084,N_5795,N_5041);
or U7085 (N_7085,N_5288,N_6130);
and U7086 (N_7086,N_6084,N_5445);
or U7087 (N_7087,N_6011,N_5817);
or U7088 (N_7088,N_5273,N_5956);
or U7089 (N_7089,N_5701,N_6077);
or U7090 (N_7090,N_5708,N_5218);
or U7091 (N_7091,N_5218,N_5395);
and U7092 (N_7092,N_5318,N_5937);
nor U7093 (N_7093,N_5543,N_6161);
or U7094 (N_7094,N_6128,N_6023);
and U7095 (N_7095,N_5857,N_5871);
nor U7096 (N_7096,N_6129,N_5321);
and U7097 (N_7097,N_5509,N_6180);
nor U7098 (N_7098,N_5314,N_5176);
and U7099 (N_7099,N_5810,N_5576);
or U7100 (N_7100,N_5136,N_6079);
or U7101 (N_7101,N_5542,N_5789);
xor U7102 (N_7102,N_5962,N_5798);
and U7103 (N_7103,N_5996,N_6180);
nand U7104 (N_7104,N_5951,N_5965);
nor U7105 (N_7105,N_5321,N_5797);
and U7106 (N_7106,N_5327,N_5239);
or U7107 (N_7107,N_5056,N_5405);
xor U7108 (N_7108,N_5546,N_5583);
or U7109 (N_7109,N_5411,N_5784);
or U7110 (N_7110,N_5449,N_5911);
nor U7111 (N_7111,N_6087,N_5115);
nor U7112 (N_7112,N_5459,N_5954);
or U7113 (N_7113,N_5316,N_5466);
nand U7114 (N_7114,N_5685,N_5463);
xor U7115 (N_7115,N_5059,N_5580);
and U7116 (N_7116,N_5773,N_5649);
and U7117 (N_7117,N_6075,N_5923);
or U7118 (N_7118,N_5058,N_6043);
nand U7119 (N_7119,N_6074,N_5192);
and U7120 (N_7120,N_6072,N_5557);
xnor U7121 (N_7121,N_5370,N_5364);
xnor U7122 (N_7122,N_6090,N_6111);
or U7123 (N_7123,N_5869,N_6056);
nand U7124 (N_7124,N_5812,N_5372);
and U7125 (N_7125,N_5564,N_5318);
nor U7126 (N_7126,N_5676,N_5888);
nor U7127 (N_7127,N_5270,N_5322);
xnor U7128 (N_7128,N_5398,N_5472);
nor U7129 (N_7129,N_5449,N_5300);
nand U7130 (N_7130,N_5340,N_6208);
nand U7131 (N_7131,N_5699,N_5681);
and U7132 (N_7132,N_5448,N_5464);
and U7133 (N_7133,N_5667,N_5026);
nor U7134 (N_7134,N_5064,N_5929);
xnor U7135 (N_7135,N_5559,N_5082);
or U7136 (N_7136,N_5377,N_5027);
nor U7137 (N_7137,N_5547,N_5532);
xor U7138 (N_7138,N_5983,N_5341);
xnor U7139 (N_7139,N_5230,N_5331);
or U7140 (N_7140,N_5737,N_5431);
xor U7141 (N_7141,N_5853,N_5462);
nand U7142 (N_7142,N_5900,N_5185);
nand U7143 (N_7143,N_5932,N_5871);
nor U7144 (N_7144,N_5768,N_5545);
nor U7145 (N_7145,N_5521,N_6145);
nand U7146 (N_7146,N_5383,N_5850);
nand U7147 (N_7147,N_5470,N_6042);
nand U7148 (N_7148,N_5569,N_5494);
or U7149 (N_7149,N_5660,N_6247);
nand U7150 (N_7150,N_5826,N_5551);
or U7151 (N_7151,N_5492,N_5319);
nand U7152 (N_7152,N_5930,N_5812);
xor U7153 (N_7153,N_5070,N_5501);
and U7154 (N_7154,N_5520,N_5938);
and U7155 (N_7155,N_6167,N_5680);
xnor U7156 (N_7156,N_5992,N_6054);
nand U7157 (N_7157,N_5475,N_5672);
nor U7158 (N_7158,N_5114,N_5448);
and U7159 (N_7159,N_6186,N_5853);
nor U7160 (N_7160,N_5573,N_5154);
xor U7161 (N_7161,N_5386,N_5824);
nor U7162 (N_7162,N_5422,N_5307);
xor U7163 (N_7163,N_5986,N_5219);
or U7164 (N_7164,N_6040,N_5239);
and U7165 (N_7165,N_6107,N_5976);
nand U7166 (N_7166,N_5557,N_5735);
nand U7167 (N_7167,N_5664,N_5332);
nand U7168 (N_7168,N_5539,N_5492);
xor U7169 (N_7169,N_5764,N_5163);
or U7170 (N_7170,N_5818,N_5063);
and U7171 (N_7171,N_5587,N_5257);
or U7172 (N_7172,N_5294,N_5283);
nor U7173 (N_7173,N_6012,N_5024);
or U7174 (N_7174,N_5217,N_6107);
nand U7175 (N_7175,N_5614,N_5917);
or U7176 (N_7176,N_6208,N_5579);
and U7177 (N_7177,N_5876,N_5794);
and U7178 (N_7178,N_5245,N_6107);
or U7179 (N_7179,N_5090,N_5988);
or U7180 (N_7180,N_5736,N_5325);
xnor U7181 (N_7181,N_5577,N_5730);
xnor U7182 (N_7182,N_5248,N_5986);
nand U7183 (N_7183,N_5188,N_6025);
or U7184 (N_7184,N_5075,N_5268);
xor U7185 (N_7185,N_5828,N_6097);
or U7186 (N_7186,N_5942,N_5192);
xor U7187 (N_7187,N_5436,N_5589);
nand U7188 (N_7188,N_6146,N_5619);
xnor U7189 (N_7189,N_5699,N_5152);
nand U7190 (N_7190,N_6177,N_5393);
xnor U7191 (N_7191,N_5206,N_5689);
nand U7192 (N_7192,N_5535,N_5956);
xnor U7193 (N_7193,N_6227,N_5546);
nand U7194 (N_7194,N_5517,N_5422);
nand U7195 (N_7195,N_5089,N_6117);
nand U7196 (N_7196,N_5677,N_5529);
or U7197 (N_7197,N_6238,N_6206);
or U7198 (N_7198,N_5478,N_5911);
or U7199 (N_7199,N_6210,N_5527);
nand U7200 (N_7200,N_5126,N_5585);
xor U7201 (N_7201,N_5198,N_5310);
nand U7202 (N_7202,N_6103,N_5499);
nand U7203 (N_7203,N_6060,N_5771);
or U7204 (N_7204,N_5642,N_5961);
xnor U7205 (N_7205,N_5701,N_5813);
xnor U7206 (N_7206,N_5416,N_5508);
nand U7207 (N_7207,N_5732,N_5517);
nand U7208 (N_7208,N_5462,N_6233);
and U7209 (N_7209,N_5961,N_5010);
or U7210 (N_7210,N_5716,N_6236);
or U7211 (N_7211,N_5207,N_5403);
nor U7212 (N_7212,N_6231,N_5283);
nand U7213 (N_7213,N_5556,N_5538);
xor U7214 (N_7214,N_6208,N_6110);
and U7215 (N_7215,N_5585,N_5277);
and U7216 (N_7216,N_5776,N_5698);
nand U7217 (N_7217,N_5419,N_6103);
and U7218 (N_7218,N_6120,N_5974);
and U7219 (N_7219,N_5120,N_5671);
nand U7220 (N_7220,N_5892,N_5354);
nand U7221 (N_7221,N_6181,N_6120);
xor U7222 (N_7222,N_5096,N_5012);
and U7223 (N_7223,N_5552,N_5345);
and U7224 (N_7224,N_5299,N_6209);
xnor U7225 (N_7225,N_5137,N_5067);
nand U7226 (N_7226,N_5550,N_5545);
xnor U7227 (N_7227,N_5070,N_5759);
nor U7228 (N_7228,N_5599,N_5610);
and U7229 (N_7229,N_5949,N_5934);
nand U7230 (N_7230,N_5690,N_5317);
and U7231 (N_7231,N_5014,N_6047);
or U7232 (N_7232,N_5190,N_5178);
and U7233 (N_7233,N_6106,N_5803);
nand U7234 (N_7234,N_5630,N_6087);
or U7235 (N_7235,N_5723,N_5194);
nor U7236 (N_7236,N_6111,N_5413);
or U7237 (N_7237,N_6078,N_5391);
or U7238 (N_7238,N_5418,N_5455);
and U7239 (N_7239,N_5153,N_5751);
or U7240 (N_7240,N_5773,N_6038);
or U7241 (N_7241,N_5056,N_5396);
nor U7242 (N_7242,N_5117,N_6231);
nand U7243 (N_7243,N_6069,N_5042);
nand U7244 (N_7244,N_5758,N_5911);
or U7245 (N_7245,N_5774,N_5130);
or U7246 (N_7246,N_6234,N_5147);
and U7247 (N_7247,N_5821,N_5765);
and U7248 (N_7248,N_5522,N_5494);
nand U7249 (N_7249,N_6135,N_5035);
xnor U7250 (N_7250,N_6179,N_5282);
and U7251 (N_7251,N_5774,N_5342);
nor U7252 (N_7252,N_5318,N_5501);
nor U7253 (N_7253,N_5276,N_5990);
nor U7254 (N_7254,N_6141,N_5321);
nor U7255 (N_7255,N_6187,N_6139);
or U7256 (N_7256,N_6067,N_5673);
nor U7257 (N_7257,N_5626,N_6091);
nor U7258 (N_7258,N_6098,N_5189);
nor U7259 (N_7259,N_6044,N_5867);
and U7260 (N_7260,N_5405,N_5579);
or U7261 (N_7261,N_5218,N_5745);
nor U7262 (N_7262,N_5659,N_6170);
nor U7263 (N_7263,N_5404,N_5166);
nor U7264 (N_7264,N_5445,N_5020);
or U7265 (N_7265,N_5674,N_5227);
nand U7266 (N_7266,N_5476,N_5514);
nor U7267 (N_7267,N_5251,N_6118);
or U7268 (N_7268,N_5649,N_5093);
and U7269 (N_7269,N_5107,N_5642);
or U7270 (N_7270,N_5848,N_5960);
xnor U7271 (N_7271,N_5322,N_5739);
and U7272 (N_7272,N_5758,N_6090);
xor U7273 (N_7273,N_5286,N_5732);
xnor U7274 (N_7274,N_5924,N_5171);
nand U7275 (N_7275,N_5352,N_5323);
nor U7276 (N_7276,N_5692,N_6137);
xnor U7277 (N_7277,N_5346,N_5132);
nand U7278 (N_7278,N_5337,N_5132);
nor U7279 (N_7279,N_5412,N_5836);
xnor U7280 (N_7280,N_6168,N_6076);
nor U7281 (N_7281,N_5478,N_5143);
nand U7282 (N_7282,N_5422,N_6235);
nor U7283 (N_7283,N_5606,N_6000);
nand U7284 (N_7284,N_5469,N_5909);
nor U7285 (N_7285,N_6047,N_5898);
xnor U7286 (N_7286,N_5750,N_5615);
nor U7287 (N_7287,N_5589,N_5654);
and U7288 (N_7288,N_5833,N_5050);
or U7289 (N_7289,N_6143,N_5841);
nor U7290 (N_7290,N_5106,N_5067);
nand U7291 (N_7291,N_5902,N_6120);
nor U7292 (N_7292,N_5180,N_5656);
or U7293 (N_7293,N_6065,N_5174);
and U7294 (N_7294,N_5145,N_5117);
and U7295 (N_7295,N_5810,N_5592);
or U7296 (N_7296,N_6050,N_5954);
nor U7297 (N_7297,N_5869,N_6132);
or U7298 (N_7298,N_5242,N_5235);
or U7299 (N_7299,N_5665,N_5760);
nand U7300 (N_7300,N_5166,N_5152);
nand U7301 (N_7301,N_6206,N_5877);
xor U7302 (N_7302,N_5468,N_5262);
nor U7303 (N_7303,N_5337,N_5357);
or U7304 (N_7304,N_5351,N_5512);
or U7305 (N_7305,N_5734,N_5913);
xnor U7306 (N_7306,N_5550,N_5293);
nor U7307 (N_7307,N_5761,N_6116);
nand U7308 (N_7308,N_6212,N_5123);
nor U7309 (N_7309,N_5796,N_6130);
or U7310 (N_7310,N_5005,N_5230);
xnor U7311 (N_7311,N_5645,N_5315);
nor U7312 (N_7312,N_5653,N_5825);
or U7313 (N_7313,N_5014,N_6008);
and U7314 (N_7314,N_5549,N_5031);
xor U7315 (N_7315,N_5752,N_6063);
nand U7316 (N_7316,N_5232,N_5498);
xnor U7317 (N_7317,N_6195,N_5465);
xnor U7318 (N_7318,N_5627,N_5892);
or U7319 (N_7319,N_5150,N_5998);
xnor U7320 (N_7320,N_5910,N_6051);
nor U7321 (N_7321,N_5964,N_5721);
or U7322 (N_7322,N_5904,N_5670);
nand U7323 (N_7323,N_5898,N_6160);
xor U7324 (N_7324,N_6009,N_5611);
nand U7325 (N_7325,N_5502,N_6026);
nor U7326 (N_7326,N_5728,N_5794);
or U7327 (N_7327,N_6163,N_5222);
nor U7328 (N_7328,N_5626,N_5629);
nand U7329 (N_7329,N_6111,N_5282);
nand U7330 (N_7330,N_6083,N_5813);
and U7331 (N_7331,N_5899,N_6067);
nor U7332 (N_7332,N_5228,N_5657);
xor U7333 (N_7333,N_6076,N_6104);
xor U7334 (N_7334,N_6056,N_6028);
or U7335 (N_7335,N_5638,N_5598);
xnor U7336 (N_7336,N_5100,N_5357);
or U7337 (N_7337,N_5065,N_5602);
or U7338 (N_7338,N_5500,N_6168);
and U7339 (N_7339,N_5453,N_5522);
xnor U7340 (N_7340,N_5150,N_5436);
xor U7341 (N_7341,N_6023,N_5617);
nand U7342 (N_7342,N_5132,N_5911);
nand U7343 (N_7343,N_5923,N_5042);
nor U7344 (N_7344,N_5372,N_6128);
nor U7345 (N_7345,N_6113,N_5867);
nand U7346 (N_7346,N_5261,N_5345);
nand U7347 (N_7347,N_6051,N_5228);
nor U7348 (N_7348,N_6011,N_5710);
and U7349 (N_7349,N_6210,N_5581);
nand U7350 (N_7350,N_6187,N_5296);
nor U7351 (N_7351,N_5543,N_5020);
or U7352 (N_7352,N_6137,N_5370);
or U7353 (N_7353,N_6114,N_5810);
nand U7354 (N_7354,N_5126,N_6088);
nor U7355 (N_7355,N_5779,N_5432);
nor U7356 (N_7356,N_5569,N_5639);
xnor U7357 (N_7357,N_5763,N_6098);
or U7358 (N_7358,N_5838,N_5790);
nand U7359 (N_7359,N_5659,N_6164);
nor U7360 (N_7360,N_5445,N_6224);
or U7361 (N_7361,N_5573,N_5717);
nor U7362 (N_7362,N_5256,N_5627);
nor U7363 (N_7363,N_5258,N_5996);
or U7364 (N_7364,N_5989,N_5497);
xor U7365 (N_7365,N_5781,N_5701);
nand U7366 (N_7366,N_5865,N_6000);
nand U7367 (N_7367,N_5096,N_5500);
nor U7368 (N_7368,N_5599,N_6094);
or U7369 (N_7369,N_5122,N_5835);
or U7370 (N_7370,N_5068,N_5183);
nand U7371 (N_7371,N_5990,N_6179);
or U7372 (N_7372,N_5530,N_6051);
or U7373 (N_7373,N_6132,N_5560);
nor U7374 (N_7374,N_5586,N_6245);
nor U7375 (N_7375,N_5421,N_5192);
or U7376 (N_7376,N_5762,N_5707);
or U7377 (N_7377,N_5423,N_6039);
or U7378 (N_7378,N_5547,N_5220);
or U7379 (N_7379,N_5060,N_6144);
xor U7380 (N_7380,N_5438,N_5164);
xor U7381 (N_7381,N_5846,N_5954);
xnor U7382 (N_7382,N_5143,N_5923);
xor U7383 (N_7383,N_5405,N_6178);
nand U7384 (N_7384,N_5006,N_5504);
nor U7385 (N_7385,N_5843,N_6154);
xnor U7386 (N_7386,N_5479,N_5594);
nor U7387 (N_7387,N_5176,N_6160);
xnor U7388 (N_7388,N_5255,N_5127);
nand U7389 (N_7389,N_5919,N_5536);
or U7390 (N_7390,N_5705,N_5436);
and U7391 (N_7391,N_6063,N_5834);
or U7392 (N_7392,N_6070,N_5670);
nor U7393 (N_7393,N_5546,N_5769);
nor U7394 (N_7394,N_6113,N_5529);
nand U7395 (N_7395,N_5295,N_6058);
or U7396 (N_7396,N_5752,N_5722);
nor U7397 (N_7397,N_5661,N_5601);
or U7398 (N_7398,N_5695,N_5896);
or U7399 (N_7399,N_5144,N_5656);
nand U7400 (N_7400,N_5291,N_5064);
xor U7401 (N_7401,N_5884,N_5517);
nor U7402 (N_7402,N_5813,N_5780);
xor U7403 (N_7403,N_5805,N_5458);
nand U7404 (N_7404,N_5582,N_5708);
and U7405 (N_7405,N_5663,N_6213);
or U7406 (N_7406,N_5210,N_6238);
nand U7407 (N_7407,N_6242,N_5817);
xor U7408 (N_7408,N_6082,N_5308);
nand U7409 (N_7409,N_6104,N_5233);
and U7410 (N_7410,N_5164,N_5858);
nand U7411 (N_7411,N_5637,N_6061);
and U7412 (N_7412,N_5016,N_5783);
and U7413 (N_7413,N_6216,N_6023);
nor U7414 (N_7414,N_6173,N_5645);
or U7415 (N_7415,N_5096,N_5395);
nor U7416 (N_7416,N_6043,N_5755);
nor U7417 (N_7417,N_5991,N_6123);
nor U7418 (N_7418,N_5195,N_5747);
nand U7419 (N_7419,N_5524,N_5280);
or U7420 (N_7420,N_5149,N_5109);
nand U7421 (N_7421,N_5561,N_5952);
and U7422 (N_7422,N_5625,N_5641);
xor U7423 (N_7423,N_5813,N_5738);
or U7424 (N_7424,N_5931,N_5426);
xnor U7425 (N_7425,N_5469,N_5797);
xor U7426 (N_7426,N_5651,N_5714);
nor U7427 (N_7427,N_5154,N_5461);
xor U7428 (N_7428,N_5843,N_5900);
nor U7429 (N_7429,N_5737,N_5934);
nor U7430 (N_7430,N_5658,N_5433);
nand U7431 (N_7431,N_5936,N_6203);
xor U7432 (N_7432,N_5912,N_6120);
or U7433 (N_7433,N_5306,N_5167);
or U7434 (N_7434,N_5199,N_5628);
nor U7435 (N_7435,N_5679,N_5498);
and U7436 (N_7436,N_5286,N_5304);
nor U7437 (N_7437,N_6210,N_5134);
and U7438 (N_7438,N_6070,N_5661);
nand U7439 (N_7439,N_6078,N_5110);
or U7440 (N_7440,N_5251,N_6091);
xor U7441 (N_7441,N_5809,N_5021);
or U7442 (N_7442,N_5717,N_5949);
nand U7443 (N_7443,N_5211,N_6235);
and U7444 (N_7444,N_5945,N_5489);
nand U7445 (N_7445,N_5155,N_5898);
nor U7446 (N_7446,N_5545,N_5248);
xnor U7447 (N_7447,N_5371,N_6198);
xnor U7448 (N_7448,N_5749,N_5555);
and U7449 (N_7449,N_5496,N_5088);
nand U7450 (N_7450,N_6195,N_6248);
nand U7451 (N_7451,N_5403,N_5418);
xnor U7452 (N_7452,N_6011,N_5503);
xor U7453 (N_7453,N_5723,N_5685);
nand U7454 (N_7454,N_5256,N_5177);
nand U7455 (N_7455,N_5399,N_5537);
or U7456 (N_7456,N_5938,N_5925);
xnor U7457 (N_7457,N_5591,N_6188);
xnor U7458 (N_7458,N_5474,N_6226);
xor U7459 (N_7459,N_5725,N_5547);
and U7460 (N_7460,N_5841,N_6115);
nor U7461 (N_7461,N_6036,N_6098);
and U7462 (N_7462,N_5978,N_5190);
or U7463 (N_7463,N_6137,N_5799);
or U7464 (N_7464,N_5928,N_5464);
nor U7465 (N_7465,N_5480,N_6201);
and U7466 (N_7466,N_5215,N_5696);
xor U7467 (N_7467,N_6060,N_5782);
or U7468 (N_7468,N_5952,N_5808);
or U7469 (N_7469,N_6132,N_5794);
or U7470 (N_7470,N_5214,N_5434);
xnor U7471 (N_7471,N_6055,N_5442);
and U7472 (N_7472,N_5701,N_5320);
and U7473 (N_7473,N_6162,N_5973);
or U7474 (N_7474,N_5460,N_5500);
nor U7475 (N_7475,N_5436,N_6044);
or U7476 (N_7476,N_5041,N_5089);
nor U7477 (N_7477,N_5293,N_5187);
xnor U7478 (N_7478,N_6097,N_5897);
xor U7479 (N_7479,N_5299,N_5754);
nand U7480 (N_7480,N_6122,N_5032);
nor U7481 (N_7481,N_6230,N_5845);
nand U7482 (N_7482,N_5856,N_6247);
xnor U7483 (N_7483,N_6070,N_5499);
and U7484 (N_7484,N_5327,N_6247);
and U7485 (N_7485,N_6073,N_5342);
xor U7486 (N_7486,N_5895,N_6020);
nand U7487 (N_7487,N_5398,N_5531);
nor U7488 (N_7488,N_5503,N_5488);
or U7489 (N_7489,N_5246,N_5776);
nand U7490 (N_7490,N_5262,N_5651);
nor U7491 (N_7491,N_5509,N_5768);
nor U7492 (N_7492,N_5481,N_5173);
nor U7493 (N_7493,N_5147,N_5677);
nand U7494 (N_7494,N_5578,N_6172);
xnor U7495 (N_7495,N_5313,N_6038);
or U7496 (N_7496,N_5180,N_5482);
xnor U7497 (N_7497,N_6108,N_5965);
nor U7498 (N_7498,N_6245,N_5792);
or U7499 (N_7499,N_6187,N_5434);
nor U7500 (N_7500,N_7013,N_6685);
xnor U7501 (N_7501,N_6341,N_6864);
nand U7502 (N_7502,N_6834,N_7221);
nor U7503 (N_7503,N_6682,N_7193);
or U7504 (N_7504,N_6468,N_6478);
and U7505 (N_7505,N_6824,N_7340);
xnor U7506 (N_7506,N_6585,N_6916);
or U7507 (N_7507,N_6778,N_6790);
xnor U7508 (N_7508,N_6499,N_7407);
and U7509 (N_7509,N_6562,N_7307);
xnor U7510 (N_7510,N_7256,N_6513);
and U7511 (N_7511,N_6668,N_6607);
xnor U7512 (N_7512,N_6703,N_7198);
xnor U7513 (N_7513,N_6310,N_7481);
xor U7514 (N_7514,N_6748,N_7357);
xnor U7515 (N_7515,N_7254,N_7294);
or U7516 (N_7516,N_7384,N_7067);
or U7517 (N_7517,N_6299,N_6776);
nor U7518 (N_7518,N_7313,N_6613);
nor U7519 (N_7519,N_6892,N_6351);
xnor U7520 (N_7520,N_7204,N_6352);
or U7521 (N_7521,N_7385,N_6569);
or U7522 (N_7522,N_7114,N_6886);
or U7523 (N_7523,N_7282,N_6885);
nand U7524 (N_7524,N_7015,N_6984);
nand U7525 (N_7525,N_7241,N_7485);
and U7526 (N_7526,N_6554,N_7492);
and U7527 (N_7527,N_6413,N_7170);
nor U7528 (N_7528,N_6485,N_6952);
xor U7529 (N_7529,N_6833,N_6504);
nor U7530 (N_7530,N_6838,N_7332);
xnor U7531 (N_7531,N_6666,N_6939);
nor U7532 (N_7532,N_6662,N_6909);
and U7533 (N_7533,N_7480,N_6544);
nor U7534 (N_7534,N_6684,N_7352);
nand U7535 (N_7535,N_7094,N_6798);
and U7536 (N_7536,N_6805,N_6789);
or U7537 (N_7537,N_6292,N_6837);
nor U7538 (N_7538,N_6333,N_6626);
nor U7539 (N_7539,N_6720,N_6603);
xnor U7540 (N_7540,N_7199,N_7403);
or U7541 (N_7541,N_7267,N_7300);
xnor U7542 (N_7542,N_7440,N_7315);
xnor U7543 (N_7543,N_6592,N_7494);
nand U7544 (N_7544,N_7394,N_6469);
nor U7545 (N_7545,N_6525,N_7181);
nand U7546 (N_7546,N_6825,N_6871);
nand U7547 (N_7547,N_6364,N_6880);
and U7548 (N_7548,N_7323,N_7257);
or U7549 (N_7549,N_7118,N_6815);
nor U7550 (N_7550,N_6502,N_7248);
or U7551 (N_7551,N_6318,N_7262);
and U7552 (N_7552,N_6641,N_6987);
nor U7553 (N_7553,N_7209,N_6579);
nor U7554 (N_7554,N_7308,N_7116);
nor U7555 (N_7555,N_7306,N_6814);
nor U7556 (N_7556,N_6313,N_6900);
xnor U7557 (N_7557,N_6951,N_7123);
or U7558 (N_7558,N_6770,N_6575);
nand U7559 (N_7559,N_7400,N_7318);
nand U7560 (N_7560,N_6922,N_6663);
nand U7561 (N_7561,N_6865,N_6978);
nand U7562 (N_7562,N_6873,N_6368);
xor U7563 (N_7563,N_7219,N_6994);
and U7564 (N_7564,N_7174,N_6411);
nor U7565 (N_7565,N_6854,N_6383);
or U7566 (N_7566,N_6869,N_6968);
xnor U7567 (N_7567,N_6903,N_6379);
and U7568 (N_7568,N_6424,N_6561);
or U7569 (N_7569,N_6983,N_6938);
or U7570 (N_7570,N_6336,N_6301);
xnor U7571 (N_7571,N_6881,N_6345);
xnor U7572 (N_7572,N_7197,N_7053);
nor U7573 (N_7573,N_6919,N_7185);
nor U7574 (N_7574,N_7234,N_7005);
and U7575 (N_7575,N_6332,N_7032);
and U7576 (N_7576,N_6761,N_7218);
or U7577 (N_7577,N_7047,N_6680);
nor U7578 (N_7578,N_7152,N_6971);
and U7579 (N_7579,N_6698,N_6969);
and U7580 (N_7580,N_6508,N_7497);
and U7581 (N_7581,N_6724,N_6399);
xor U7582 (N_7582,N_6997,N_6889);
nor U7583 (N_7583,N_7115,N_7406);
xor U7584 (N_7584,N_6564,N_6774);
nand U7585 (N_7585,N_7206,N_6599);
and U7586 (N_7586,N_7127,N_7455);
and U7587 (N_7587,N_7371,N_7432);
nand U7588 (N_7588,N_6705,N_7413);
nand U7589 (N_7589,N_7243,N_6709);
or U7590 (N_7590,N_7078,N_6557);
nor U7591 (N_7591,N_6665,N_6386);
xnor U7592 (N_7592,N_7430,N_7097);
nand U7593 (N_7593,N_6573,N_7088);
or U7594 (N_7594,N_7498,N_7040);
nor U7595 (N_7595,N_6325,N_7454);
nor U7596 (N_7596,N_7309,N_6960);
xnor U7597 (N_7597,N_7439,N_7145);
nor U7598 (N_7598,N_7264,N_6921);
nor U7599 (N_7599,N_6850,N_6539);
nand U7600 (N_7600,N_7423,N_6392);
xor U7601 (N_7601,N_7141,N_6286);
and U7602 (N_7602,N_6689,N_7251);
or U7603 (N_7603,N_6500,N_6631);
and U7604 (N_7604,N_7249,N_6363);
and U7605 (N_7605,N_6330,N_6782);
nor U7606 (N_7606,N_6962,N_7082);
nand U7607 (N_7607,N_6745,N_6870);
or U7608 (N_7608,N_7111,N_7240);
nand U7609 (N_7609,N_6560,N_6576);
and U7610 (N_7610,N_7464,N_6786);
and U7611 (N_7611,N_6675,N_6718);
nor U7612 (N_7612,N_7212,N_7024);
or U7613 (N_7613,N_6595,N_6635);
nand U7614 (N_7614,N_6660,N_7071);
nor U7615 (N_7615,N_6862,N_7232);
nor U7616 (N_7616,N_6510,N_7333);
and U7617 (N_7617,N_6722,N_7102);
nand U7618 (N_7618,N_6326,N_6337);
xor U7619 (N_7619,N_7390,N_6540);
xor U7620 (N_7620,N_6591,N_6811);
nor U7621 (N_7621,N_7069,N_6929);
or U7622 (N_7622,N_6739,N_6849);
xnor U7623 (N_7623,N_6781,N_7353);
nor U7624 (N_7624,N_6537,N_7148);
and U7625 (N_7625,N_6656,N_6602);
xor U7626 (N_7626,N_6910,N_7250);
nor U7627 (N_7627,N_6260,N_6580);
or U7628 (N_7628,N_6650,N_7054);
or U7629 (N_7629,N_7428,N_6498);
or U7630 (N_7630,N_7006,N_7038);
and U7631 (N_7631,N_7190,N_6767);
xnor U7632 (N_7632,N_6528,N_7136);
and U7633 (N_7633,N_6694,N_7211);
nor U7634 (N_7634,N_7237,N_6716);
or U7635 (N_7635,N_6412,N_6877);
nand U7636 (N_7636,N_6421,N_6594);
and U7637 (N_7637,N_7387,N_6477);
xnor U7638 (N_7638,N_7335,N_6842);
and U7639 (N_7639,N_7161,N_6653);
or U7640 (N_7640,N_7466,N_7443);
nor U7641 (N_7641,N_6358,N_6691);
nand U7642 (N_7642,N_7080,N_7397);
xnor U7643 (N_7643,N_6747,N_7052);
xor U7644 (N_7644,N_7475,N_6643);
nor U7645 (N_7645,N_7220,N_6494);
nand U7646 (N_7646,N_6751,N_6290);
and U7647 (N_7647,N_6863,N_6566);
xnor U7648 (N_7648,N_6911,N_7336);
nand U7649 (N_7649,N_6415,N_6568);
xnor U7650 (N_7650,N_7496,N_7391);
xnor U7651 (N_7651,N_7245,N_6453);
nand U7652 (N_7652,N_6993,N_7351);
nor U7653 (N_7653,N_7096,N_6484);
nor U7654 (N_7654,N_6674,N_6407);
nor U7655 (N_7655,N_7280,N_7091);
and U7656 (N_7656,N_6901,N_7459);
nor U7657 (N_7657,N_6376,N_7292);
nand U7658 (N_7658,N_6306,N_6370);
nand U7659 (N_7659,N_6622,N_6460);
nand U7660 (N_7660,N_7229,N_6394);
xor U7661 (N_7661,N_6257,N_6533);
and U7662 (N_7662,N_6746,N_7304);
nor U7663 (N_7663,N_6466,N_6479);
xnor U7664 (N_7664,N_6645,N_7214);
nand U7665 (N_7665,N_7416,N_7062);
and U7666 (N_7666,N_7298,N_7195);
and U7667 (N_7667,N_6324,N_7408);
or U7668 (N_7668,N_6866,N_7470);
nor U7669 (N_7669,N_6604,N_6446);
or U7670 (N_7670,N_6536,N_6273);
nor U7671 (N_7671,N_7489,N_6395);
and U7672 (N_7672,N_7433,N_6841);
nand U7673 (N_7673,N_6282,N_6719);
xnor U7674 (N_7674,N_6744,N_6859);
nand U7675 (N_7675,N_6483,N_6338);
xor U7676 (N_7676,N_7020,N_7007);
nor U7677 (N_7677,N_6633,N_6311);
xnor U7678 (N_7678,N_6893,N_6343);
xor U7679 (N_7679,N_6549,N_7027);
and U7680 (N_7680,N_6879,N_6760);
and U7681 (N_7681,N_6270,N_7399);
nand U7682 (N_7682,N_6924,N_6572);
or U7683 (N_7683,N_6927,N_7187);
or U7684 (N_7684,N_7499,N_6753);
nor U7685 (N_7685,N_7339,N_6287);
and U7686 (N_7686,N_6342,N_6737);
or U7687 (N_7687,N_6953,N_6616);
or U7688 (N_7688,N_6956,N_6868);
or U7689 (N_7689,N_6456,N_7177);
and U7690 (N_7690,N_6496,N_6339);
and U7691 (N_7691,N_7401,N_6743);
and U7692 (N_7692,N_6371,N_6923);
or U7693 (N_7693,N_7004,N_7441);
and U7694 (N_7694,N_6957,N_7448);
or U7695 (N_7695,N_6894,N_6891);
xor U7696 (N_7696,N_7119,N_6804);
xor U7697 (N_7697,N_6320,N_7365);
and U7698 (N_7698,N_7429,N_7488);
xor U7699 (N_7699,N_7477,N_7095);
nor U7700 (N_7700,N_6813,N_7044);
nor U7701 (N_7701,N_7216,N_6296);
nor U7702 (N_7702,N_6571,N_7479);
or U7703 (N_7703,N_6522,N_7246);
xnor U7704 (N_7704,N_6312,N_6915);
and U7705 (N_7705,N_6808,N_6601);
and U7706 (N_7706,N_6816,N_7056);
or U7707 (N_7707,N_6552,N_7143);
nand U7708 (N_7708,N_6696,N_6988);
nor U7709 (N_7709,N_6940,N_6433);
nor U7710 (N_7710,N_6692,N_6657);
nand U7711 (N_7711,N_6418,N_7350);
nor U7712 (N_7712,N_7129,N_7085);
or U7713 (N_7713,N_6711,N_7046);
or U7714 (N_7714,N_7151,N_6373);
xnor U7715 (N_7715,N_7073,N_6729);
xnor U7716 (N_7716,N_6832,N_6487);
and U7717 (N_7717,N_6520,N_7182);
or U7718 (N_7718,N_6807,N_7048);
xor U7719 (N_7719,N_6565,N_7421);
nor U7720 (N_7720,N_6905,N_6791);
and U7721 (N_7721,N_7079,N_7301);
nand U7722 (N_7722,N_7456,N_7184);
nor U7723 (N_7723,N_7355,N_6925);
or U7724 (N_7724,N_6389,N_7453);
nand U7725 (N_7725,N_7382,N_7128);
nand U7726 (N_7726,N_6545,N_7173);
xnor U7727 (N_7727,N_6829,N_6878);
or U7728 (N_7728,N_6426,N_7144);
and U7729 (N_7729,N_7370,N_7068);
xor U7730 (N_7730,N_6272,N_6884);
xnor U7731 (N_7731,N_6252,N_6627);
xnor U7732 (N_7732,N_7369,N_6796);
or U7733 (N_7733,N_6405,N_6876);
xnor U7734 (N_7734,N_7472,N_6624);
or U7735 (N_7735,N_6874,N_7230);
or U7736 (N_7736,N_7233,N_6896);
or U7737 (N_7737,N_7157,N_6372);
or U7738 (N_7738,N_7140,N_6276);
and U7739 (N_7739,N_6442,N_6895);
or U7740 (N_7740,N_6797,N_6348);
and U7741 (N_7741,N_6681,N_6269);
xor U7742 (N_7742,N_6608,N_7081);
nand U7743 (N_7743,N_6979,N_6470);
or U7744 (N_7744,N_6844,N_7106);
nand U7745 (N_7745,N_6687,N_6949);
and U7746 (N_7746,N_6437,N_6340);
or U7747 (N_7747,N_7099,N_7021);
nor U7748 (N_7748,N_7154,N_6490);
nor U7749 (N_7749,N_6511,N_7261);
nand U7750 (N_7750,N_6697,N_7389);
and U7751 (N_7751,N_6861,N_7050);
xor U7752 (N_7752,N_6611,N_7431);
nand U7753 (N_7753,N_6596,N_6731);
nand U7754 (N_7754,N_6904,N_6823);
and U7755 (N_7755,N_6985,N_7271);
nor U7756 (N_7756,N_6977,N_6738);
xnor U7757 (N_7757,N_7137,N_7314);
and U7758 (N_7758,N_7328,N_7058);
nand U7759 (N_7759,N_7124,N_6839);
or U7760 (N_7760,N_6678,N_7017);
or U7761 (N_7761,N_6817,N_6550);
or U7762 (N_7762,N_7077,N_7166);
and U7763 (N_7763,N_6365,N_7295);
nor U7764 (N_7764,N_6941,N_7253);
nand U7765 (N_7765,N_7192,N_6652);
nor U7766 (N_7766,N_6582,N_6523);
or U7767 (N_7767,N_7200,N_6621);
or U7768 (N_7768,N_6827,N_6414);
nor U7769 (N_7769,N_6427,N_6473);
xnor U7770 (N_7770,N_6639,N_6907);
nand U7771 (N_7771,N_6733,N_7134);
or U7772 (N_7772,N_7034,N_6913);
nand U7773 (N_7773,N_7378,N_6360);
xnor U7774 (N_7774,N_6688,N_6806);
nand U7775 (N_7775,N_6600,N_7434);
xnor U7776 (N_7776,N_6930,N_6742);
nand U7777 (N_7777,N_6809,N_6712);
nor U7778 (N_7778,N_6515,N_7270);
nand U7779 (N_7779,N_6589,N_7213);
xnor U7780 (N_7780,N_6771,N_6958);
nand U7781 (N_7781,N_6556,N_6261);
and U7782 (N_7782,N_6636,N_7409);
xnor U7783 (N_7783,N_7338,N_6555);
nand U7784 (N_7784,N_6779,N_7277);
and U7785 (N_7785,N_7093,N_6417);
nor U7786 (N_7786,N_6353,N_7347);
and U7787 (N_7787,N_7359,N_7083);
and U7788 (N_7788,N_6534,N_6448);
and U7789 (N_7789,N_6543,N_7285);
nand U7790 (N_7790,N_6449,N_6787);
nor U7791 (N_7791,N_6435,N_6375);
nand U7792 (N_7792,N_6707,N_6777);
xor U7793 (N_7793,N_7417,N_7325);
nor U7794 (N_7794,N_7284,N_6784);
nor U7795 (N_7795,N_7147,N_7103);
nor U7796 (N_7796,N_7450,N_7022);
xnor U7797 (N_7797,N_7263,N_6480);
and U7798 (N_7798,N_6769,N_7225);
xnor U7799 (N_7799,N_6259,N_7065);
and U7800 (N_7800,N_7405,N_6492);
or U7801 (N_7801,N_6950,N_6380);
and U7802 (N_7802,N_6975,N_6506);
or U7803 (N_7803,N_7210,N_7286);
or U7804 (N_7804,N_6420,N_7364);
nand U7805 (N_7805,N_7160,N_6553);
or U7806 (N_7806,N_7414,N_6683);
xor U7807 (N_7807,N_6423,N_6967);
nor U7808 (N_7808,N_7312,N_7373);
xor U7809 (N_7809,N_7003,N_6799);
nor U7810 (N_7810,N_7425,N_7076);
or U7811 (N_7811,N_6846,N_7037);
nand U7812 (N_7812,N_6280,N_7162);
and U7813 (N_7813,N_6455,N_6519);
nand U7814 (N_7814,N_6759,N_6998);
xor U7815 (N_7815,N_6443,N_7363);
xor U7816 (N_7816,N_7383,N_6476);
nand U7817 (N_7817,N_6377,N_6640);
nand U7818 (N_7818,N_6757,N_7420);
xor U7819 (N_7819,N_7461,N_7009);
or U7820 (N_7820,N_6538,N_7183);
nand U7821 (N_7821,N_6676,N_7109);
or U7822 (N_7822,N_6514,N_6830);
xor U7823 (N_7823,N_6278,N_7484);
and U7824 (N_7824,N_6762,N_6357);
xnor U7825 (N_7825,N_7012,N_6404);
or U7826 (N_7826,N_6465,N_7236);
nor U7827 (N_7827,N_6917,N_7061);
nor U7828 (N_7828,N_7419,N_7337);
and U7829 (N_7829,N_6574,N_7331);
or U7830 (N_7830,N_7036,N_7223);
nor U7831 (N_7831,N_6661,N_7486);
nor U7832 (N_7832,N_6634,N_6847);
and U7833 (N_7833,N_6942,N_6704);
xor U7834 (N_7834,N_7011,N_7155);
xnor U7835 (N_7835,N_6463,N_7194);
and U7836 (N_7836,N_6819,N_6385);
or U7837 (N_7837,N_6964,N_6361);
nand U7838 (N_7838,N_6587,N_6647);
or U7839 (N_7839,N_6717,N_6867);
and U7840 (N_7840,N_6321,N_6546);
nand U7841 (N_7841,N_7089,N_6788);
nand U7842 (N_7842,N_7168,N_7342);
or U7843 (N_7843,N_6772,N_7458);
or U7844 (N_7844,N_7474,N_7287);
or U7845 (N_7845,N_7327,N_6251);
nor U7846 (N_7846,N_6851,N_7231);
nand U7847 (N_7847,N_6831,N_7202);
and U7848 (N_7848,N_6531,N_6700);
or U7849 (N_7849,N_6714,N_7074);
nand U7850 (N_7850,N_7296,N_7031);
or U7851 (N_7851,N_6763,N_7469);
nand U7852 (N_7852,N_7297,N_7483);
or U7853 (N_7853,N_6670,N_6721);
and U7854 (N_7854,N_7275,N_6464);
or U7855 (N_7855,N_6529,N_7468);
xnor U7856 (N_7856,N_6298,N_7100);
xnor U7857 (N_7857,N_6995,N_6532);
and U7858 (N_7858,N_7130,N_6605);
and U7859 (N_7859,N_7139,N_7276);
nand U7860 (N_7860,N_6293,N_6673);
nand U7861 (N_7861,N_6996,N_7110);
or U7862 (N_7862,N_7279,N_6517);
nand U7863 (N_7863,N_7217,N_6277);
and U7864 (N_7864,N_6570,N_7438);
and U7865 (N_7865,N_6725,N_6547);
and U7866 (N_7866,N_7422,N_6936);
nand U7867 (N_7867,N_6436,N_6501);
xnor U7868 (N_7868,N_7346,N_6822);
xor U7869 (N_7869,N_7164,N_7235);
nor U7870 (N_7870,N_6530,N_7228);
xor U7871 (N_7871,N_6651,N_6902);
or U7872 (N_7872,N_6398,N_6431);
and U7873 (N_7873,N_6860,N_7321);
and U7874 (N_7874,N_7478,N_7060);
or U7875 (N_7875,N_7238,N_6335);
nor U7876 (N_7876,N_6820,N_6541);
xor U7877 (N_7877,N_7258,N_6291);
nor U7878 (N_7878,N_6265,N_6275);
or U7879 (N_7879,N_6669,N_6344);
nand U7880 (N_7880,N_7268,N_6381);
or U7881 (N_7881,N_7135,N_6754);
or U7882 (N_7882,N_6734,N_7092);
or U7883 (N_7883,N_7188,N_6255);
nand U7884 (N_7884,N_7150,N_6526);
and U7885 (N_7885,N_7437,N_7226);
or U7886 (N_7886,N_7142,N_7377);
xnor U7887 (N_7887,N_6391,N_7462);
or U7888 (N_7888,N_6999,N_6388);
xor U7889 (N_7889,N_7395,N_6920);
xnor U7890 (N_7890,N_7293,N_7444);
nand U7891 (N_7891,N_6471,N_7205);
and U7892 (N_7892,N_7146,N_6946);
xnor U7893 (N_7893,N_6323,N_6440);
nor U7894 (N_7894,N_6706,N_6852);
nand U7895 (N_7895,N_7386,N_7348);
nor U7896 (N_7896,N_6783,N_6558);
xnor U7897 (N_7897,N_6677,N_6349);
or U7898 (N_7898,N_6285,N_6367);
and U7899 (N_7899,N_6409,N_6818);
and U7900 (N_7900,N_6289,N_7112);
xnor U7901 (N_7901,N_6434,N_7222);
nand U7902 (N_7902,N_6853,N_6785);
xor U7903 (N_7903,N_6690,N_7344);
nand U7904 (N_7904,N_7426,N_6664);
or U7905 (N_7905,N_6752,N_6482);
xnor U7906 (N_7906,N_6315,N_7467);
nand U7907 (N_7907,N_7418,N_7288);
nand U7908 (N_7908,N_7104,N_6593);
xor U7909 (N_7909,N_7122,N_7179);
and U7910 (N_7910,N_6974,N_6359);
nor U7911 (N_7911,N_7379,N_6396);
nand U7912 (N_7912,N_6474,N_6933);
nor U7913 (N_7913,N_7266,N_6328);
nand U7914 (N_7914,N_7404,N_6989);
xnor U7915 (N_7915,N_6935,N_6812);
xor U7916 (N_7916,N_7084,N_7274);
and U7917 (N_7917,N_7131,N_7107);
nor U7918 (N_7918,N_6267,N_6966);
or U7919 (N_7919,N_6708,N_7402);
nor U7920 (N_7920,N_7070,N_6932);
nor U7921 (N_7921,N_6948,N_7039);
xnor U7922 (N_7922,N_6872,N_6459);
xnor U7923 (N_7923,N_7473,N_6931);
or U7924 (N_7924,N_6727,N_7030);
or U7925 (N_7925,N_7343,N_7023);
or U7926 (N_7926,N_6659,N_6644);
xnor U7927 (N_7927,N_6461,N_6350);
and U7928 (N_7928,N_7349,N_7055);
xnor U7929 (N_7929,N_6256,N_6454);
and U7930 (N_7930,N_6356,N_6524);
and U7931 (N_7931,N_6495,N_6726);
nor U7932 (N_7932,N_6535,N_7334);
or U7933 (N_7933,N_6638,N_6620);
nand U7934 (N_7934,N_7354,N_6567);
xnor U7935 (N_7935,N_6281,N_7172);
and U7936 (N_7936,N_6374,N_6992);
xor U7937 (N_7937,N_6382,N_6390);
xnor U7938 (N_7938,N_6491,N_6715);
and U7939 (N_7939,N_6625,N_6457);
xor U7940 (N_7940,N_6710,N_7010);
nand U7941 (N_7941,N_7303,N_6648);
nand U7942 (N_7942,N_6283,N_6982);
xnor U7943 (N_7943,N_6462,N_7396);
nor U7944 (N_7944,N_7043,N_6497);
and U7945 (N_7945,N_6583,N_7330);
nand U7946 (N_7946,N_6548,N_6410);
xnor U7947 (N_7947,N_7283,N_7113);
nand U7948 (N_7948,N_7487,N_6322);
nor U7949 (N_7949,N_7059,N_7117);
xor U7950 (N_7950,N_7465,N_6944);
xor U7951 (N_7951,N_6947,N_6912);
and U7952 (N_7952,N_7072,N_6972);
nor U7953 (N_7953,N_6990,N_6764);
or U7954 (N_7954,N_6581,N_6756);
nor U7955 (N_7955,N_7042,N_6749);
and U7956 (N_7956,N_7196,N_6821);
or U7957 (N_7957,N_6793,N_6632);
xnor U7958 (N_7958,N_6472,N_6327);
nand U7959 (N_7959,N_6897,N_6493);
or U7960 (N_7960,N_6890,N_7490);
and U7961 (N_7961,N_6578,N_6887);
nand U7962 (N_7962,N_7326,N_6354);
and U7963 (N_7963,N_6981,N_7493);
xor U7964 (N_7964,N_6505,N_7090);
nor U7965 (N_7965,N_6918,N_6857);
nor U7966 (N_7966,N_7026,N_6305);
nand U7967 (N_7967,N_7272,N_6836);
nor U7968 (N_7968,N_7311,N_7302);
and U7969 (N_7969,N_6654,N_7362);
and U7970 (N_7970,N_6963,N_6735);
or U7971 (N_7971,N_6402,N_7075);
xor U7972 (N_7972,N_6355,N_6598);
xnor U7973 (N_7973,N_7086,N_6810);
xor U7974 (N_7974,N_7033,N_6615);
and U7975 (N_7975,N_7446,N_6628);
xor U7976 (N_7976,N_7310,N_6646);
and U7977 (N_7977,N_6792,N_6362);
and U7978 (N_7978,N_7153,N_6955);
nor U7979 (N_7979,N_7415,N_7452);
nor U7980 (N_7980,N_6366,N_6250);
xor U7981 (N_7981,N_7203,N_6845);
and U7982 (N_7982,N_6618,N_7000);
nand U7983 (N_7983,N_6408,N_6467);
nand U7984 (N_7984,N_6403,N_7063);
nor U7985 (N_7985,N_6658,N_7175);
and U7986 (N_7986,N_7201,N_6794);
nor U7987 (N_7987,N_6450,N_6630);
nand U7988 (N_7988,N_7041,N_6503);
nor U7989 (N_7989,N_7299,N_6268);
or U7990 (N_7990,N_6303,N_6898);
nor U7991 (N_7991,N_6765,N_6264);
or U7992 (N_7992,N_6279,N_6610);
nand U7993 (N_7993,N_6667,N_6439);
xnor U7994 (N_7994,N_7322,N_7014);
nand U7995 (N_7995,N_6518,N_6750);
nand U7996 (N_7996,N_6295,N_6856);
xor U7997 (N_7997,N_6489,N_7372);
nor U7998 (N_7998,N_7361,N_6713);
xnor U7999 (N_7999,N_7002,N_7329);
xnor U8000 (N_8000,N_6438,N_6429);
and U8001 (N_8001,N_6945,N_6773);
nand U8002 (N_8002,N_7163,N_6649);
nor U8003 (N_8003,N_7045,N_7207);
or U8004 (N_8004,N_7451,N_6699);
and U8005 (N_8005,N_6258,N_6314);
nand U8006 (N_8006,N_7066,N_7289);
nand U8007 (N_8007,N_7049,N_6447);
and U8008 (N_8008,N_6802,N_7411);
nor U8009 (N_8009,N_7178,N_6430);
and U8010 (N_8010,N_6284,N_7035);
xnor U8011 (N_8011,N_7412,N_6766);
or U8012 (N_8012,N_7180,N_6686);
nand U8013 (N_8013,N_6384,N_6954);
xor U8014 (N_8014,N_6521,N_6906);
xor U8015 (N_8015,N_7016,N_7018);
xnor U8016 (N_8016,N_6693,N_7224);
nor U8017 (N_8017,N_6271,N_6609);
or U8018 (N_8018,N_6393,N_6980);
nand U8019 (N_8019,N_6481,N_7368);
or U8020 (N_8020,N_6588,N_7227);
and U8021 (N_8021,N_7239,N_6253);
xnor U8022 (N_8022,N_6262,N_6614);
nand U8023 (N_8023,N_6316,N_7374);
nand U8024 (N_8024,N_6319,N_6826);
xor U8025 (N_8025,N_7132,N_6551);
or U8026 (N_8026,N_7491,N_6527);
and U8027 (N_8027,N_7269,N_7133);
and U8028 (N_8028,N_7247,N_7410);
and U8029 (N_8029,N_6347,N_6451);
and U8030 (N_8030,N_7156,N_6679);
nand U8031 (N_8031,N_7019,N_6835);
nand U8032 (N_8032,N_7457,N_6309);
nand U8033 (N_8033,N_6655,N_7424);
nand U8034 (N_8034,N_6458,N_7358);
xor U8035 (N_8035,N_7149,N_6507);
or U8036 (N_8036,N_6559,N_7189);
xor U8037 (N_8037,N_6976,N_6848);
and U8038 (N_8038,N_7290,N_7176);
nor U8039 (N_8039,N_7165,N_6425);
xor U8040 (N_8040,N_6755,N_6800);
xor U8041 (N_8041,N_7215,N_6914);
nor U8042 (N_8042,N_7393,N_6973);
nor U8043 (N_8043,N_7375,N_6331);
xor U8044 (N_8044,N_6937,N_7392);
and U8045 (N_8045,N_6855,N_7125);
or U8046 (N_8046,N_7460,N_6888);
or U8047 (N_8047,N_6263,N_7259);
or U8048 (N_8048,N_6803,N_6516);
nor U8049 (N_8049,N_7381,N_6961);
xnor U8050 (N_8050,N_6934,N_6828);
nor U8051 (N_8051,N_7447,N_6444);
xor U8052 (N_8052,N_6758,N_7445);
nor U8053 (N_8053,N_6586,N_6991);
xnor U8054 (N_8054,N_6304,N_7367);
or U8055 (N_8055,N_7121,N_7341);
and U8056 (N_8056,N_6775,N_6612);
and U8057 (N_8057,N_7471,N_6346);
nand U8058 (N_8058,N_7191,N_6928);
and U8059 (N_8059,N_7305,N_6619);
nand U8060 (N_8060,N_7495,N_7138);
or U8061 (N_8061,N_6701,N_6736);
and U8062 (N_8062,N_7126,N_6406);
nand U8063 (N_8063,N_7320,N_7098);
nand U8064 (N_8064,N_7345,N_6419);
nor U8065 (N_8065,N_6266,N_6882);
nor U8066 (N_8066,N_6629,N_6740);
nand U8067 (N_8067,N_6965,N_6445);
xor U8068 (N_8068,N_7281,N_7105);
and U8069 (N_8069,N_6617,N_7316);
or U8070 (N_8070,N_6432,N_7265);
and U8071 (N_8071,N_7029,N_7087);
and U8072 (N_8072,N_7319,N_6422);
nand U8073 (N_8073,N_6441,N_6702);
nor U8074 (N_8074,N_6730,N_7167);
xor U8075 (N_8075,N_7252,N_7008);
or U8076 (N_8076,N_6563,N_7278);
nand U8077 (N_8077,N_6843,N_6307);
nor U8078 (N_8078,N_6584,N_6475);
or U8079 (N_8079,N_7158,N_6986);
or U8080 (N_8080,N_6488,N_7366);
or U8081 (N_8081,N_6695,N_7101);
or U8082 (N_8082,N_6329,N_7317);
and U8083 (N_8083,N_6334,N_7064);
nand U8084 (N_8084,N_7051,N_7108);
and U8085 (N_8085,N_7025,N_6671);
nand U8086 (N_8086,N_6590,N_6512);
xnor U8087 (N_8087,N_6732,N_7120);
or U8088 (N_8088,N_7376,N_7171);
nand U8089 (N_8089,N_7427,N_6959);
or U8090 (N_8090,N_7436,N_6428);
or U8091 (N_8091,N_6943,N_7360);
and U8092 (N_8092,N_6387,N_7255);
or U8093 (N_8093,N_7356,N_6254);
and U8094 (N_8094,N_6401,N_6741);
xnor U8095 (N_8095,N_6397,N_6378);
xor U8096 (N_8096,N_7244,N_7398);
and U8097 (N_8097,N_6840,N_6970);
and U8098 (N_8098,N_7449,N_6597);
nor U8099 (N_8099,N_6768,N_6899);
and U8100 (N_8100,N_6577,N_6780);
or U8101 (N_8101,N_6300,N_7208);
xor U8102 (N_8102,N_7186,N_7001);
nor U8103 (N_8103,N_7028,N_6400);
nor U8104 (N_8104,N_6606,N_6416);
or U8105 (N_8105,N_6274,N_7482);
nor U8106 (N_8106,N_6623,N_6637);
or U8107 (N_8107,N_6926,N_6308);
nor U8108 (N_8108,N_7435,N_6728);
xor U8109 (N_8109,N_6875,N_6452);
nand U8110 (N_8110,N_7388,N_6672);
xor U8111 (N_8111,N_7169,N_6908);
or U8112 (N_8112,N_7324,N_6723);
nor U8113 (N_8113,N_7476,N_7463);
or U8114 (N_8114,N_6486,N_7159);
and U8115 (N_8115,N_7260,N_7442);
nand U8116 (N_8116,N_6288,N_6883);
or U8117 (N_8117,N_7057,N_6801);
and U8118 (N_8118,N_6302,N_6795);
nor U8119 (N_8119,N_6317,N_7380);
xor U8120 (N_8120,N_6858,N_6369);
and U8121 (N_8121,N_6642,N_7273);
and U8122 (N_8122,N_6297,N_6294);
and U8123 (N_8123,N_6509,N_7291);
or U8124 (N_8124,N_6542,N_7242);
nor U8125 (N_8125,N_7150,N_7144);
xnor U8126 (N_8126,N_6843,N_6314);
or U8127 (N_8127,N_7117,N_6776);
nand U8128 (N_8128,N_7375,N_7075);
nand U8129 (N_8129,N_6647,N_6518);
or U8130 (N_8130,N_7184,N_7337);
or U8131 (N_8131,N_6987,N_7079);
nand U8132 (N_8132,N_7421,N_7385);
xor U8133 (N_8133,N_7035,N_7196);
xor U8134 (N_8134,N_7355,N_6421);
xnor U8135 (N_8135,N_7337,N_6770);
xor U8136 (N_8136,N_6431,N_6409);
xor U8137 (N_8137,N_7305,N_6728);
or U8138 (N_8138,N_6928,N_7210);
nand U8139 (N_8139,N_6273,N_6603);
nand U8140 (N_8140,N_6397,N_6366);
nand U8141 (N_8141,N_6489,N_6765);
or U8142 (N_8142,N_6399,N_6974);
nor U8143 (N_8143,N_6836,N_6551);
and U8144 (N_8144,N_6861,N_6846);
nand U8145 (N_8145,N_7210,N_6545);
or U8146 (N_8146,N_7483,N_7287);
and U8147 (N_8147,N_6847,N_7185);
nand U8148 (N_8148,N_7487,N_6533);
and U8149 (N_8149,N_7104,N_6414);
or U8150 (N_8150,N_6506,N_6690);
and U8151 (N_8151,N_7044,N_6799);
nand U8152 (N_8152,N_6979,N_6958);
nand U8153 (N_8153,N_6430,N_6310);
xor U8154 (N_8154,N_6605,N_6600);
xnor U8155 (N_8155,N_6255,N_6817);
or U8156 (N_8156,N_7231,N_7410);
xnor U8157 (N_8157,N_7233,N_6847);
nor U8158 (N_8158,N_6920,N_6502);
and U8159 (N_8159,N_7044,N_7132);
nand U8160 (N_8160,N_7483,N_7081);
xor U8161 (N_8161,N_7032,N_6591);
nand U8162 (N_8162,N_7428,N_7169);
nand U8163 (N_8163,N_7343,N_6658);
xnor U8164 (N_8164,N_7140,N_7225);
xor U8165 (N_8165,N_6796,N_6497);
xor U8166 (N_8166,N_7212,N_6851);
and U8167 (N_8167,N_7096,N_6563);
xnor U8168 (N_8168,N_6274,N_6897);
and U8169 (N_8169,N_6349,N_6656);
or U8170 (N_8170,N_6530,N_7342);
or U8171 (N_8171,N_6919,N_7331);
xnor U8172 (N_8172,N_6638,N_6701);
xnor U8173 (N_8173,N_6769,N_6841);
and U8174 (N_8174,N_6950,N_7104);
nand U8175 (N_8175,N_7456,N_6368);
and U8176 (N_8176,N_6458,N_6500);
and U8177 (N_8177,N_6567,N_6690);
or U8178 (N_8178,N_7126,N_7059);
or U8179 (N_8179,N_7269,N_7400);
nor U8180 (N_8180,N_6674,N_6648);
nor U8181 (N_8181,N_7009,N_7412);
or U8182 (N_8182,N_7032,N_6536);
or U8183 (N_8183,N_6383,N_6785);
or U8184 (N_8184,N_7102,N_7476);
nor U8185 (N_8185,N_6974,N_6429);
and U8186 (N_8186,N_6484,N_6926);
nand U8187 (N_8187,N_6821,N_7142);
or U8188 (N_8188,N_7316,N_6632);
nor U8189 (N_8189,N_7290,N_6728);
xnor U8190 (N_8190,N_6268,N_6795);
nand U8191 (N_8191,N_6864,N_6402);
nor U8192 (N_8192,N_7190,N_6339);
nand U8193 (N_8193,N_7254,N_7103);
and U8194 (N_8194,N_7261,N_6408);
nand U8195 (N_8195,N_7343,N_6510);
nor U8196 (N_8196,N_6339,N_7119);
xnor U8197 (N_8197,N_6689,N_7018);
or U8198 (N_8198,N_6801,N_6624);
nor U8199 (N_8199,N_6838,N_7484);
nand U8200 (N_8200,N_6921,N_6896);
xnor U8201 (N_8201,N_7071,N_7403);
nand U8202 (N_8202,N_6892,N_6562);
xor U8203 (N_8203,N_7373,N_6910);
and U8204 (N_8204,N_6716,N_7088);
nand U8205 (N_8205,N_7184,N_7336);
nor U8206 (N_8206,N_7200,N_7438);
nor U8207 (N_8207,N_6423,N_6420);
and U8208 (N_8208,N_6554,N_6516);
or U8209 (N_8209,N_6872,N_6562);
nand U8210 (N_8210,N_6399,N_6804);
and U8211 (N_8211,N_6965,N_6954);
xnor U8212 (N_8212,N_7018,N_6306);
or U8213 (N_8213,N_7381,N_7443);
and U8214 (N_8214,N_7321,N_7352);
or U8215 (N_8215,N_6907,N_6662);
nor U8216 (N_8216,N_7305,N_6559);
nand U8217 (N_8217,N_6854,N_7281);
or U8218 (N_8218,N_7020,N_6687);
or U8219 (N_8219,N_6955,N_7011);
xnor U8220 (N_8220,N_7051,N_7194);
nand U8221 (N_8221,N_7168,N_6515);
nand U8222 (N_8222,N_7109,N_6407);
xnor U8223 (N_8223,N_6532,N_6828);
and U8224 (N_8224,N_6534,N_6761);
nand U8225 (N_8225,N_6770,N_6682);
nor U8226 (N_8226,N_7277,N_6413);
and U8227 (N_8227,N_7243,N_6982);
or U8228 (N_8228,N_6870,N_6625);
xor U8229 (N_8229,N_6544,N_6528);
nand U8230 (N_8230,N_6890,N_6835);
xnor U8231 (N_8231,N_6310,N_6959);
or U8232 (N_8232,N_7276,N_7273);
nand U8233 (N_8233,N_6530,N_7390);
nand U8234 (N_8234,N_7282,N_6895);
nor U8235 (N_8235,N_6582,N_7437);
xnor U8236 (N_8236,N_7425,N_6318);
nand U8237 (N_8237,N_7324,N_6272);
and U8238 (N_8238,N_6315,N_7169);
or U8239 (N_8239,N_6693,N_6362);
nand U8240 (N_8240,N_7061,N_6739);
or U8241 (N_8241,N_6272,N_6975);
nand U8242 (N_8242,N_6516,N_6402);
or U8243 (N_8243,N_6854,N_7181);
and U8244 (N_8244,N_6357,N_7130);
or U8245 (N_8245,N_6343,N_6775);
xor U8246 (N_8246,N_7297,N_7410);
nor U8247 (N_8247,N_7378,N_6273);
or U8248 (N_8248,N_6438,N_7210);
nand U8249 (N_8249,N_6360,N_7431);
xnor U8250 (N_8250,N_6309,N_6431);
and U8251 (N_8251,N_7159,N_6565);
nand U8252 (N_8252,N_7387,N_7041);
nor U8253 (N_8253,N_6796,N_6623);
or U8254 (N_8254,N_7483,N_6591);
or U8255 (N_8255,N_7100,N_6602);
and U8256 (N_8256,N_7252,N_7025);
xor U8257 (N_8257,N_6494,N_7040);
nand U8258 (N_8258,N_6920,N_6640);
nor U8259 (N_8259,N_6964,N_7081);
nor U8260 (N_8260,N_7090,N_6551);
nand U8261 (N_8261,N_6881,N_7447);
nand U8262 (N_8262,N_7068,N_6826);
nor U8263 (N_8263,N_6767,N_6739);
or U8264 (N_8264,N_6682,N_6627);
xnor U8265 (N_8265,N_6495,N_6652);
nor U8266 (N_8266,N_7076,N_6781);
or U8267 (N_8267,N_7049,N_6839);
or U8268 (N_8268,N_6747,N_6529);
nor U8269 (N_8269,N_6268,N_7429);
nand U8270 (N_8270,N_6278,N_6651);
xor U8271 (N_8271,N_7447,N_6269);
nor U8272 (N_8272,N_6368,N_6993);
xor U8273 (N_8273,N_7008,N_6977);
nand U8274 (N_8274,N_7087,N_6854);
nand U8275 (N_8275,N_7272,N_6677);
and U8276 (N_8276,N_7406,N_7395);
nor U8277 (N_8277,N_7367,N_7369);
nand U8278 (N_8278,N_6542,N_6895);
nor U8279 (N_8279,N_6394,N_7050);
or U8280 (N_8280,N_6289,N_6682);
nand U8281 (N_8281,N_7136,N_7467);
or U8282 (N_8282,N_6727,N_6574);
nand U8283 (N_8283,N_6444,N_7400);
nor U8284 (N_8284,N_6653,N_7215);
and U8285 (N_8285,N_6672,N_6308);
xnor U8286 (N_8286,N_6255,N_7168);
and U8287 (N_8287,N_7428,N_6671);
or U8288 (N_8288,N_6642,N_6369);
xnor U8289 (N_8289,N_7361,N_6521);
xnor U8290 (N_8290,N_6546,N_6326);
xnor U8291 (N_8291,N_7294,N_7018);
and U8292 (N_8292,N_7263,N_6872);
xnor U8293 (N_8293,N_6852,N_6751);
and U8294 (N_8294,N_7145,N_7031);
or U8295 (N_8295,N_6593,N_6524);
and U8296 (N_8296,N_7414,N_6567);
nand U8297 (N_8297,N_7101,N_7168);
or U8298 (N_8298,N_6429,N_6783);
and U8299 (N_8299,N_6998,N_7168);
and U8300 (N_8300,N_6965,N_7447);
nand U8301 (N_8301,N_6980,N_6414);
nor U8302 (N_8302,N_6290,N_6413);
or U8303 (N_8303,N_7423,N_6822);
nor U8304 (N_8304,N_6458,N_6794);
nor U8305 (N_8305,N_6467,N_6411);
or U8306 (N_8306,N_7029,N_7066);
nand U8307 (N_8307,N_6679,N_7047);
nand U8308 (N_8308,N_7085,N_6995);
nand U8309 (N_8309,N_7369,N_6408);
nor U8310 (N_8310,N_6588,N_7287);
nor U8311 (N_8311,N_6638,N_7181);
nand U8312 (N_8312,N_6506,N_7457);
and U8313 (N_8313,N_7428,N_7191);
nand U8314 (N_8314,N_6821,N_7050);
nor U8315 (N_8315,N_7120,N_6341);
nand U8316 (N_8316,N_6471,N_6658);
xnor U8317 (N_8317,N_7479,N_6521);
or U8318 (N_8318,N_7301,N_7392);
or U8319 (N_8319,N_7049,N_6516);
xor U8320 (N_8320,N_7054,N_6682);
nor U8321 (N_8321,N_7385,N_6703);
nand U8322 (N_8322,N_6970,N_7155);
or U8323 (N_8323,N_7400,N_7265);
and U8324 (N_8324,N_6824,N_6503);
nand U8325 (N_8325,N_7120,N_6340);
nand U8326 (N_8326,N_6553,N_7000);
and U8327 (N_8327,N_6838,N_7248);
or U8328 (N_8328,N_6260,N_6881);
xor U8329 (N_8329,N_6663,N_6912);
and U8330 (N_8330,N_7203,N_6904);
nand U8331 (N_8331,N_6828,N_6331);
and U8332 (N_8332,N_7413,N_7337);
nand U8333 (N_8333,N_7228,N_6690);
xnor U8334 (N_8334,N_6841,N_6388);
nand U8335 (N_8335,N_6823,N_6794);
nor U8336 (N_8336,N_6828,N_6276);
xor U8337 (N_8337,N_6474,N_6664);
nand U8338 (N_8338,N_7434,N_6297);
nor U8339 (N_8339,N_6458,N_6682);
nand U8340 (N_8340,N_7016,N_7329);
nor U8341 (N_8341,N_6488,N_7021);
xnor U8342 (N_8342,N_6524,N_7172);
nand U8343 (N_8343,N_7479,N_7109);
xnor U8344 (N_8344,N_7189,N_7383);
nand U8345 (N_8345,N_6813,N_6531);
or U8346 (N_8346,N_7110,N_6731);
xnor U8347 (N_8347,N_7117,N_7086);
nor U8348 (N_8348,N_7055,N_7461);
nor U8349 (N_8349,N_7099,N_6709);
nor U8350 (N_8350,N_7014,N_6571);
xor U8351 (N_8351,N_7295,N_7253);
and U8352 (N_8352,N_6957,N_6546);
or U8353 (N_8353,N_6764,N_6285);
xnor U8354 (N_8354,N_6927,N_6618);
xor U8355 (N_8355,N_7461,N_7486);
or U8356 (N_8356,N_7415,N_7450);
nand U8357 (N_8357,N_6510,N_6742);
nor U8358 (N_8358,N_7483,N_7484);
xor U8359 (N_8359,N_6994,N_7430);
xor U8360 (N_8360,N_6601,N_7401);
nor U8361 (N_8361,N_6502,N_6815);
or U8362 (N_8362,N_7062,N_7367);
xnor U8363 (N_8363,N_7441,N_7211);
xor U8364 (N_8364,N_6493,N_6787);
nor U8365 (N_8365,N_6551,N_6878);
and U8366 (N_8366,N_6524,N_6340);
nor U8367 (N_8367,N_6921,N_7329);
nand U8368 (N_8368,N_7096,N_6627);
xnor U8369 (N_8369,N_7022,N_6952);
xor U8370 (N_8370,N_6597,N_6992);
and U8371 (N_8371,N_6402,N_6802);
and U8372 (N_8372,N_6274,N_7223);
xnor U8373 (N_8373,N_6639,N_6597);
nand U8374 (N_8374,N_6910,N_7110);
nand U8375 (N_8375,N_7471,N_6704);
and U8376 (N_8376,N_6263,N_7210);
nor U8377 (N_8377,N_6884,N_6672);
and U8378 (N_8378,N_7254,N_6428);
and U8379 (N_8379,N_7400,N_6505);
nor U8380 (N_8380,N_7153,N_6701);
xnor U8381 (N_8381,N_7058,N_7437);
xnor U8382 (N_8382,N_7001,N_7348);
and U8383 (N_8383,N_7314,N_7150);
or U8384 (N_8384,N_6510,N_7360);
nand U8385 (N_8385,N_6275,N_6282);
nor U8386 (N_8386,N_7333,N_6832);
nor U8387 (N_8387,N_7025,N_6982);
and U8388 (N_8388,N_7461,N_6799);
xnor U8389 (N_8389,N_6297,N_6664);
or U8390 (N_8390,N_6598,N_7110);
nand U8391 (N_8391,N_6502,N_6735);
and U8392 (N_8392,N_7293,N_6674);
xor U8393 (N_8393,N_6956,N_6365);
nor U8394 (N_8394,N_6768,N_7034);
nand U8395 (N_8395,N_7376,N_6946);
or U8396 (N_8396,N_7302,N_6308);
nand U8397 (N_8397,N_6904,N_7488);
nand U8398 (N_8398,N_6620,N_7116);
xor U8399 (N_8399,N_7392,N_7426);
nand U8400 (N_8400,N_6450,N_6984);
xnor U8401 (N_8401,N_6655,N_6925);
or U8402 (N_8402,N_7238,N_6359);
and U8403 (N_8403,N_7280,N_6708);
xnor U8404 (N_8404,N_7374,N_6394);
or U8405 (N_8405,N_6351,N_7491);
nand U8406 (N_8406,N_7019,N_6309);
or U8407 (N_8407,N_7406,N_7011);
or U8408 (N_8408,N_6427,N_7277);
xor U8409 (N_8409,N_7471,N_6368);
nand U8410 (N_8410,N_7439,N_6500);
or U8411 (N_8411,N_6433,N_6913);
and U8412 (N_8412,N_6826,N_7462);
and U8413 (N_8413,N_6498,N_6447);
nor U8414 (N_8414,N_7094,N_6568);
or U8415 (N_8415,N_7211,N_6708);
and U8416 (N_8416,N_6441,N_7119);
and U8417 (N_8417,N_6986,N_7155);
nor U8418 (N_8418,N_7390,N_6766);
and U8419 (N_8419,N_6952,N_6830);
and U8420 (N_8420,N_6831,N_6826);
and U8421 (N_8421,N_7018,N_7108);
xnor U8422 (N_8422,N_7179,N_6953);
nor U8423 (N_8423,N_7094,N_7114);
xor U8424 (N_8424,N_6295,N_7435);
xor U8425 (N_8425,N_6599,N_6283);
nor U8426 (N_8426,N_6812,N_7308);
xor U8427 (N_8427,N_7414,N_6983);
or U8428 (N_8428,N_7206,N_6460);
and U8429 (N_8429,N_6453,N_6713);
and U8430 (N_8430,N_6622,N_7413);
and U8431 (N_8431,N_7295,N_7474);
or U8432 (N_8432,N_6333,N_6914);
nor U8433 (N_8433,N_6941,N_6960);
xor U8434 (N_8434,N_6311,N_7286);
xor U8435 (N_8435,N_6858,N_6592);
xor U8436 (N_8436,N_7062,N_6498);
nand U8437 (N_8437,N_7493,N_6370);
or U8438 (N_8438,N_6442,N_6783);
and U8439 (N_8439,N_7328,N_7136);
nor U8440 (N_8440,N_6636,N_6725);
xor U8441 (N_8441,N_7078,N_7101);
and U8442 (N_8442,N_7181,N_6904);
nor U8443 (N_8443,N_6894,N_6581);
nor U8444 (N_8444,N_7399,N_6829);
nor U8445 (N_8445,N_6791,N_6902);
xnor U8446 (N_8446,N_6426,N_7022);
and U8447 (N_8447,N_7261,N_6288);
or U8448 (N_8448,N_7176,N_6924);
or U8449 (N_8449,N_6447,N_7265);
nand U8450 (N_8450,N_6904,N_7447);
nor U8451 (N_8451,N_6746,N_6324);
or U8452 (N_8452,N_7290,N_6606);
and U8453 (N_8453,N_7378,N_6806);
nor U8454 (N_8454,N_6454,N_7195);
or U8455 (N_8455,N_6917,N_6566);
nor U8456 (N_8456,N_6425,N_7345);
and U8457 (N_8457,N_6633,N_6997);
nor U8458 (N_8458,N_7392,N_6818);
or U8459 (N_8459,N_6857,N_6364);
and U8460 (N_8460,N_7200,N_7362);
or U8461 (N_8461,N_7274,N_7309);
nand U8462 (N_8462,N_7281,N_7009);
and U8463 (N_8463,N_7246,N_7073);
nor U8464 (N_8464,N_7066,N_6292);
and U8465 (N_8465,N_6343,N_6342);
or U8466 (N_8466,N_7387,N_6799);
and U8467 (N_8467,N_6269,N_6968);
or U8468 (N_8468,N_7302,N_6301);
nand U8469 (N_8469,N_7223,N_6565);
xor U8470 (N_8470,N_6805,N_6386);
xnor U8471 (N_8471,N_7473,N_6551);
or U8472 (N_8472,N_6945,N_7460);
nor U8473 (N_8473,N_7229,N_6382);
nand U8474 (N_8474,N_6264,N_6905);
or U8475 (N_8475,N_7034,N_6328);
and U8476 (N_8476,N_6251,N_7242);
or U8477 (N_8477,N_6370,N_6865);
and U8478 (N_8478,N_6767,N_6814);
and U8479 (N_8479,N_7093,N_6977);
and U8480 (N_8480,N_7421,N_6387);
and U8481 (N_8481,N_7054,N_6970);
or U8482 (N_8482,N_6406,N_6366);
nand U8483 (N_8483,N_7108,N_6466);
xnor U8484 (N_8484,N_6273,N_7343);
nand U8485 (N_8485,N_6314,N_6470);
nor U8486 (N_8486,N_7046,N_6402);
or U8487 (N_8487,N_7332,N_7091);
nand U8488 (N_8488,N_6892,N_6598);
xnor U8489 (N_8489,N_6884,N_7172);
xor U8490 (N_8490,N_6533,N_7326);
nand U8491 (N_8491,N_6809,N_6705);
or U8492 (N_8492,N_7250,N_6480);
xor U8493 (N_8493,N_6829,N_6957);
or U8494 (N_8494,N_6433,N_6879);
xnor U8495 (N_8495,N_6654,N_6857);
and U8496 (N_8496,N_7103,N_6731);
nand U8497 (N_8497,N_7033,N_6642);
nand U8498 (N_8498,N_6907,N_7487);
nor U8499 (N_8499,N_7137,N_6406);
and U8500 (N_8500,N_7345,N_7014);
or U8501 (N_8501,N_6542,N_6448);
or U8502 (N_8502,N_6285,N_7015);
and U8503 (N_8503,N_6423,N_6338);
or U8504 (N_8504,N_6382,N_6812);
xor U8505 (N_8505,N_7139,N_6938);
xor U8506 (N_8506,N_7220,N_6875);
or U8507 (N_8507,N_7052,N_7088);
or U8508 (N_8508,N_6936,N_7133);
nand U8509 (N_8509,N_6948,N_6286);
nor U8510 (N_8510,N_6393,N_6685);
and U8511 (N_8511,N_7434,N_6728);
and U8512 (N_8512,N_6292,N_6273);
nand U8513 (N_8513,N_6381,N_6537);
nor U8514 (N_8514,N_6280,N_6344);
xor U8515 (N_8515,N_6441,N_7253);
nand U8516 (N_8516,N_6928,N_6805);
and U8517 (N_8517,N_6709,N_7386);
nor U8518 (N_8518,N_6614,N_7154);
xor U8519 (N_8519,N_7061,N_6885);
nor U8520 (N_8520,N_7099,N_6861);
or U8521 (N_8521,N_7412,N_7357);
nand U8522 (N_8522,N_7480,N_7164);
nor U8523 (N_8523,N_6559,N_7149);
or U8524 (N_8524,N_6359,N_7013);
nand U8525 (N_8525,N_6724,N_6978);
nand U8526 (N_8526,N_6808,N_6448);
or U8527 (N_8527,N_7315,N_6932);
or U8528 (N_8528,N_6869,N_6966);
xor U8529 (N_8529,N_7086,N_7223);
or U8530 (N_8530,N_7349,N_7316);
nand U8531 (N_8531,N_6272,N_6732);
nor U8532 (N_8532,N_6809,N_6670);
nor U8533 (N_8533,N_7273,N_6256);
nor U8534 (N_8534,N_6565,N_7303);
xnor U8535 (N_8535,N_6890,N_6317);
xnor U8536 (N_8536,N_6397,N_6721);
xnor U8537 (N_8537,N_6569,N_6768);
nand U8538 (N_8538,N_6501,N_6607);
and U8539 (N_8539,N_6844,N_7028);
and U8540 (N_8540,N_7131,N_7002);
or U8541 (N_8541,N_6918,N_7336);
or U8542 (N_8542,N_7040,N_6686);
nor U8543 (N_8543,N_6537,N_7041);
nand U8544 (N_8544,N_7317,N_6349);
nor U8545 (N_8545,N_7351,N_7120);
and U8546 (N_8546,N_7169,N_6998);
nor U8547 (N_8547,N_7334,N_6996);
and U8548 (N_8548,N_7051,N_6679);
and U8549 (N_8549,N_6828,N_6754);
nor U8550 (N_8550,N_7147,N_6938);
or U8551 (N_8551,N_6580,N_7462);
nand U8552 (N_8552,N_6724,N_6778);
xor U8553 (N_8553,N_7491,N_6825);
nor U8554 (N_8554,N_6444,N_6538);
xor U8555 (N_8555,N_6917,N_6342);
or U8556 (N_8556,N_6985,N_6649);
xnor U8557 (N_8557,N_6333,N_6465);
nand U8558 (N_8558,N_6736,N_7087);
and U8559 (N_8559,N_7326,N_6406);
xor U8560 (N_8560,N_7355,N_6258);
xnor U8561 (N_8561,N_7088,N_6930);
nor U8562 (N_8562,N_7423,N_6606);
or U8563 (N_8563,N_7399,N_6387);
xor U8564 (N_8564,N_6919,N_7171);
and U8565 (N_8565,N_6951,N_6485);
nand U8566 (N_8566,N_6470,N_7392);
or U8567 (N_8567,N_6645,N_7391);
and U8568 (N_8568,N_6452,N_7491);
or U8569 (N_8569,N_6853,N_7485);
nor U8570 (N_8570,N_6674,N_7054);
nand U8571 (N_8571,N_6945,N_7421);
nand U8572 (N_8572,N_7058,N_7184);
nand U8573 (N_8573,N_6790,N_6798);
or U8574 (N_8574,N_6291,N_6968);
and U8575 (N_8575,N_6444,N_6335);
or U8576 (N_8576,N_7110,N_7004);
or U8577 (N_8577,N_6325,N_7062);
and U8578 (N_8578,N_6965,N_6583);
nor U8579 (N_8579,N_7274,N_6265);
or U8580 (N_8580,N_6448,N_7334);
nand U8581 (N_8581,N_7407,N_6802);
xor U8582 (N_8582,N_7054,N_7289);
or U8583 (N_8583,N_6527,N_6719);
or U8584 (N_8584,N_7248,N_6972);
or U8585 (N_8585,N_6806,N_6410);
or U8586 (N_8586,N_6387,N_7265);
nand U8587 (N_8587,N_7088,N_6659);
nand U8588 (N_8588,N_6929,N_7126);
nand U8589 (N_8589,N_7458,N_6980);
nor U8590 (N_8590,N_7449,N_6819);
nand U8591 (N_8591,N_7217,N_7027);
nor U8592 (N_8592,N_6901,N_7026);
or U8593 (N_8593,N_7491,N_6544);
xnor U8594 (N_8594,N_6465,N_7150);
or U8595 (N_8595,N_7296,N_7221);
nor U8596 (N_8596,N_6980,N_6552);
and U8597 (N_8597,N_6841,N_7086);
and U8598 (N_8598,N_7075,N_6325);
nand U8599 (N_8599,N_7161,N_6612);
and U8600 (N_8600,N_6773,N_6648);
or U8601 (N_8601,N_7442,N_6849);
xnor U8602 (N_8602,N_7128,N_6502);
nand U8603 (N_8603,N_7449,N_7103);
nand U8604 (N_8604,N_7265,N_6702);
xor U8605 (N_8605,N_6978,N_6635);
or U8606 (N_8606,N_6904,N_7258);
xor U8607 (N_8607,N_7018,N_7335);
nand U8608 (N_8608,N_6867,N_7081);
or U8609 (N_8609,N_6574,N_7377);
or U8610 (N_8610,N_6740,N_6256);
xor U8611 (N_8611,N_6869,N_6505);
and U8612 (N_8612,N_6765,N_6529);
xor U8613 (N_8613,N_6821,N_6951);
xor U8614 (N_8614,N_7350,N_6323);
xor U8615 (N_8615,N_7377,N_6748);
nand U8616 (N_8616,N_6656,N_7279);
nor U8617 (N_8617,N_6808,N_6764);
nor U8618 (N_8618,N_6839,N_6301);
or U8619 (N_8619,N_7425,N_6365);
nor U8620 (N_8620,N_7244,N_7466);
nand U8621 (N_8621,N_6993,N_6929);
nor U8622 (N_8622,N_6476,N_7264);
and U8623 (N_8623,N_7085,N_7187);
nand U8624 (N_8624,N_6509,N_7214);
or U8625 (N_8625,N_6539,N_6465);
xor U8626 (N_8626,N_7439,N_6485);
nor U8627 (N_8627,N_6412,N_6813);
nand U8628 (N_8628,N_6584,N_6694);
or U8629 (N_8629,N_6335,N_6341);
or U8630 (N_8630,N_6273,N_6877);
xor U8631 (N_8631,N_6979,N_6788);
nor U8632 (N_8632,N_6311,N_7013);
or U8633 (N_8633,N_7329,N_6879);
and U8634 (N_8634,N_6684,N_7233);
nand U8635 (N_8635,N_6884,N_7274);
xor U8636 (N_8636,N_7343,N_6750);
or U8637 (N_8637,N_6778,N_6502);
nand U8638 (N_8638,N_7463,N_6255);
nor U8639 (N_8639,N_7440,N_6273);
and U8640 (N_8640,N_7045,N_6587);
xnor U8641 (N_8641,N_7465,N_7166);
nand U8642 (N_8642,N_7140,N_7079);
nor U8643 (N_8643,N_6582,N_7242);
and U8644 (N_8644,N_7428,N_7433);
nand U8645 (N_8645,N_6350,N_6760);
or U8646 (N_8646,N_6406,N_7360);
or U8647 (N_8647,N_7250,N_6584);
nand U8648 (N_8648,N_7328,N_6996);
or U8649 (N_8649,N_7109,N_6345);
or U8650 (N_8650,N_6405,N_7266);
or U8651 (N_8651,N_7228,N_6926);
xor U8652 (N_8652,N_6474,N_6692);
and U8653 (N_8653,N_6256,N_6416);
nand U8654 (N_8654,N_7372,N_7297);
and U8655 (N_8655,N_6421,N_6692);
nor U8656 (N_8656,N_7393,N_7046);
nand U8657 (N_8657,N_7065,N_6781);
and U8658 (N_8658,N_7114,N_7188);
or U8659 (N_8659,N_6339,N_6640);
nor U8660 (N_8660,N_7344,N_7273);
xnor U8661 (N_8661,N_6803,N_6556);
and U8662 (N_8662,N_6513,N_6905);
nand U8663 (N_8663,N_6653,N_6819);
nand U8664 (N_8664,N_6329,N_7322);
or U8665 (N_8665,N_6920,N_6500);
or U8666 (N_8666,N_6288,N_6860);
or U8667 (N_8667,N_6843,N_6433);
or U8668 (N_8668,N_6425,N_7389);
nor U8669 (N_8669,N_7147,N_6820);
nor U8670 (N_8670,N_6611,N_6423);
nor U8671 (N_8671,N_6838,N_6549);
nand U8672 (N_8672,N_7243,N_6962);
nor U8673 (N_8673,N_7483,N_7108);
nand U8674 (N_8674,N_7028,N_7353);
and U8675 (N_8675,N_7182,N_6568);
or U8676 (N_8676,N_6322,N_7386);
or U8677 (N_8677,N_6280,N_7248);
nor U8678 (N_8678,N_7323,N_6844);
nor U8679 (N_8679,N_6841,N_7302);
nand U8680 (N_8680,N_7253,N_7380);
nand U8681 (N_8681,N_7159,N_7331);
nor U8682 (N_8682,N_6320,N_7337);
nand U8683 (N_8683,N_7043,N_7205);
or U8684 (N_8684,N_6808,N_7350);
nor U8685 (N_8685,N_6444,N_6500);
xnor U8686 (N_8686,N_6482,N_6463);
nor U8687 (N_8687,N_6295,N_6321);
and U8688 (N_8688,N_6377,N_7480);
nand U8689 (N_8689,N_6864,N_6743);
nor U8690 (N_8690,N_6717,N_7253);
nor U8691 (N_8691,N_7066,N_7181);
or U8692 (N_8692,N_6617,N_6535);
xnor U8693 (N_8693,N_6648,N_6590);
xor U8694 (N_8694,N_6458,N_7236);
and U8695 (N_8695,N_6570,N_7489);
or U8696 (N_8696,N_6587,N_7347);
xnor U8697 (N_8697,N_6759,N_7440);
and U8698 (N_8698,N_6871,N_6501);
nand U8699 (N_8699,N_6734,N_7494);
xor U8700 (N_8700,N_6975,N_7289);
nor U8701 (N_8701,N_6296,N_7494);
or U8702 (N_8702,N_7192,N_6980);
nand U8703 (N_8703,N_7384,N_6670);
nand U8704 (N_8704,N_6974,N_6290);
nor U8705 (N_8705,N_6771,N_7453);
and U8706 (N_8706,N_6779,N_7376);
xnor U8707 (N_8707,N_6401,N_7452);
or U8708 (N_8708,N_7026,N_7223);
and U8709 (N_8709,N_6482,N_6428);
or U8710 (N_8710,N_7152,N_7407);
nand U8711 (N_8711,N_7410,N_6458);
and U8712 (N_8712,N_7238,N_6515);
nand U8713 (N_8713,N_6364,N_7385);
nor U8714 (N_8714,N_6405,N_6353);
and U8715 (N_8715,N_6806,N_6984);
nor U8716 (N_8716,N_7054,N_6381);
and U8717 (N_8717,N_6621,N_7257);
nand U8718 (N_8718,N_6811,N_6795);
nor U8719 (N_8719,N_7346,N_6720);
and U8720 (N_8720,N_7266,N_6319);
and U8721 (N_8721,N_6964,N_7086);
xnor U8722 (N_8722,N_6268,N_6705);
xor U8723 (N_8723,N_7243,N_6620);
nor U8724 (N_8724,N_6981,N_7180);
nor U8725 (N_8725,N_6986,N_7457);
or U8726 (N_8726,N_7422,N_6707);
xor U8727 (N_8727,N_6304,N_7481);
nor U8728 (N_8728,N_7316,N_6563);
nand U8729 (N_8729,N_6950,N_7009);
nand U8730 (N_8730,N_6868,N_7067);
xor U8731 (N_8731,N_7006,N_7381);
and U8732 (N_8732,N_7474,N_6293);
and U8733 (N_8733,N_6677,N_6799);
or U8734 (N_8734,N_6330,N_7137);
or U8735 (N_8735,N_6561,N_6261);
nand U8736 (N_8736,N_6467,N_7405);
or U8737 (N_8737,N_6997,N_6412);
or U8738 (N_8738,N_7140,N_7134);
and U8739 (N_8739,N_6729,N_6431);
and U8740 (N_8740,N_7346,N_6420);
or U8741 (N_8741,N_6474,N_7375);
xnor U8742 (N_8742,N_6659,N_6682);
and U8743 (N_8743,N_6807,N_7002);
nor U8744 (N_8744,N_7279,N_6980);
xnor U8745 (N_8745,N_6674,N_6652);
nor U8746 (N_8746,N_7455,N_6835);
and U8747 (N_8747,N_6548,N_7298);
and U8748 (N_8748,N_7435,N_7454);
nor U8749 (N_8749,N_7146,N_7342);
xor U8750 (N_8750,N_7978,N_8528);
nor U8751 (N_8751,N_8048,N_8044);
xnor U8752 (N_8752,N_8713,N_8588);
and U8753 (N_8753,N_8018,N_8672);
or U8754 (N_8754,N_8057,N_8236);
or U8755 (N_8755,N_7993,N_8223);
xor U8756 (N_8756,N_7576,N_8167);
or U8757 (N_8757,N_8724,N_8093);
and U8758 (N_8758,N_8301,N_7778);
nand U8759 (N_8759,N_8158,N_7785);
nor U8760 (N_8760,N_8164,N_8328);
xnor U8761 (N_8761,N_7983,N_8388);
nand U8762 (N_8762,N_8368,N_8186);
nand U8763 (N_8763,N_8137,N_8337);
and U8764 (N_8764,N_8051,N_8639);
and U8765 (N_8765,N_8210,N_7768);
or U8766 (N_8766,N_7554,N_7617);
and U8767 (N_8767,N_8042,N_8105);
and U8768 (N_8768,N_8361,N_8670);
or U8769 (N_8769,N_7527,N_7774);
xnor U8770 (N_8770,N_8172,N_8159);
xor U8771 (N_8771,N_8017,N_7919);
and U8772 (N_8772,N_7917,N_8094);
nor U8773 (N_8773,N_7505,N_8088);
xnor U8774 (N_8774,N_8671,N_8596);
or U8775 (N_8775,N_7786,N_8128);
nand U8776 (N_8776,N_7870,N_8099);
nand U8777 (N_8777,N_7562,N_8590);
and U8778 (N_8778,N_8379,N_7784);
nor U8779 (N_8779,N_8106,N_7904);
and U8780 (N_8780,N_7963,N_8631);
or U8781 (N_8781,N_8216,N_8552);
nand U8782 (N_8782,N_8119,N_8173);
nand U8783 (N_8783,N_7747,N_8634);
and U8784 (N_8784,N_7691,N_7654);
nor U8785 (N_8785,N_7821,N_8605);
nor U8786 (N_8786,N_8180,N_8476);
nor U8787 (N_8787,N_7560,N_7994);
nand U8788 (N_8788,N_8657,N_8129);
nor U8789 (N_8789,N_7912,N_7638);
or U8790 (N_8790,N_7659,N_8225);
nor U8791 (N_8791,N_8649,N_8263);
nand U8792 (N_8792,N_7507,N_8356);
nor U8793 (N_8793,N_7591,N_7825);
nor U8794 (N_8794,N_7893,N_7865);
or U8795 (N_8795,N_7707,N_8147);
xnor U8796 (N_8796,N_7552,N_7502);
and U8797 (N_8797,N_8743,N_8660);
nand U8798 (N_8798,N_7705,N_8015);
xnor U8799 (N_8799,N_8347,N_7824);
or U8800 (N_8800,N_8206,N_8747);
xor U8801 (N_8801,N_8011,N_8560);
xnor U8802 (N_8802,N_8456,N_8124);
nand U8803 (N_8803,N_7811,N_7672);
and U8804 (N_8804,N_8086,N_8358);
nor U8805 (N_8805,N_7814,N_8055);
xnor U8806 (N_8806,N_8187,N_8679);
xnor U8807 (N_8807,N_8324,N_7533);
or U8808 (N_8808,N_7548,N_8498);
nand U8809 (N_8809,N_8647,N_8281);
or U8810 (N_8810,N_8344,N_8242);
nand U8811 (N_8811,N_7667,N_8694);
and U8812 (N_8812,N_8544,N_7750);
xor U8813 (N_8813,N_8475,N_8635);
or U8814 (N_8814,N_7823,N_8697);
or U8815 (N_8815,N_8633,N_8268);
nand U8816 (N_8816,N_8563,N_8643);
or U8817 (N_8817,N_7635,N_8036);
nor U8818 (N_8818,N_7520,N_7905);
xor U8819 (N_8819,N_8529,N_8097);
or U8820 (N_8820,N_8653,N_7506);
nor U8821 (N_8821,N_8708,N_7839);
nand U8822 (N_8822,N_7655,N_8402);
or U8823 (N_8823,N_8580,N_8079);
and U8824 (N_8824,N_7696,N_8480);
or U8825 (N_8825,N_7923,N_8355);
nor U8826 (N_8826,N_8722,N_7595);
nor U8827 (N_8827,N_7868,N_8441);
xnor U8828 (N_8828,N_8006,N_8212);
or U8829 (N_8829,N_7967,N_8168);
nor U8830 (N_8830,N_8244,N_8618);
xor U8831 (N_8831,N_8197,N_7982);
nand U8832 (N_8832,N_8686,N_8472);
nor U8833 (N_8833,N_8235,N_8690);
or U8834 (N_8834,N_8515,N_8287);
and U8835 (N_8835,N_8485,N_8295);
xnor U8836 (N_8836,N_8698,N_7657);
nor U8837 (N_8837,N_7561,N_7932);
and U8838 (N_8838,N_8246,N_7934);
xor U8839 (N_8839,N_8422,N_8658);
nor U8840 (N_8840,N_8196,N_8502);
xor U8841 (N_8841,N_8539,N_7519);
and U8842 (N_8842,N_8360,N_7801);
nand U8843 (N_8843,N_7602,N_8313);
or U8844 (N_8844,N_7564,N_8117);
and U8845 (N_8845,N_8334,N_8192);
or U8846 (N_8846,N_7544,N_8260);
nand U8847 (N_8847,N_7951,N_8642);
or U8848 (N_8848,N_8102,N_8004);
nand U8849 (N_8849,N_8150,N_8156);
and U8850 (N_8850,N_8655,N_8453);
xnor U8851 (N_8851,N_7847,N_8477);
and U8852 (N_8852,N_8030,N_7566);
nand U8853 (N_8853,N_8659,N_8711);
or U8854 (N_8854,N_7930,N_8449);
nand U8855 (N_8855,N_7517,N_7709);
nor U8856 (N_8856,N_7733,N_8134);
xnor U8857 (N_8857,N_7626,N_7619);
and U8858 (N_8858,N_7641,N_8406);
nor U8859 (N_8859,N_7515,N_7933);
and U8860 (N_8860,N_8250,N_8296);
nor U8861 (N_8861,N_8194,N_7920);
nor U8862 (N_8862,N_7910,N_7628);
or U8863 (N_8863,N_8740,N_7601);
nand U8864 (N_8864,N_7568,N_8614);
nand U8865 (N_8865,N_8325,N_8511);
xor U8866 (N_8866,N_7528,N_8022);
nand U8867 (N_8867,N_7632,N_8569);
xnor U8868 (N_8868,N_8601,N_8567);
xnor U8869 (N_8869,N_8664,N_8510);
xor U8870 (N_8870,N_7772,N_7926);
and U8871 (N_8871,N_8503,N_8182);
xnor U8872 (N_8872,N_8043,N_8056);
nand U8873 (N_8873,N_8509,N_7715);
xor U8874 (N_8874,N_8507,N_8157);
nor U8875 (N_8875,N_8024,N_7556);
xnor U8876 (N_8876,N_8416,N_7902);
nand U8877 (N_8877,N_7749,N_8508);
xnor U8878 (N_8878,N_7866,N_7843);
nand U8879 (N_8879,N_7583,N_8204);
xnor U8880 (N_8880,N_8597,N_8673);
xor U8881 (N_8881,N_7804,N_8426);
nand U8882 (N_8882,N_8266,N_7985);
xor U8883 (N_8883,N_8491,N_8166);
nor U8884 (N_8884,N_7521,N_7991);
xnor U8885 (N_8885,N_8745,N_8321);
and U8886 (N_8886,N_8153,N_8237);
and U8887 (N_8887,N_7639,N_7625);
nand U8888 (N_8888,N_7692,N_7661);
xnor U8889 (N_8889,N_8543,N_7935);
and U8890 (N_8890,N_7722,N_7634);
xor U8891 (N_8891,N_8059,N_7553);
nor U8892 (N_8892,N_8314,N_8098);
xnor U8893 (N_8893,N_8683,N_8726);
nor U8894 (N_8894,N_8365,N_8691);
or U8895 (N_8895,N_7597,N_8739);
nor U8896 (N_8896,N_8113,N_7909);
and U8897 (N_8897,N_7802,N_8568);
nand U8898 (N_8898,N_8359,N_8371);
and U8899 (N_8899,N_8702,N_8257);
nor U8900 (N_8900,N_7777,N_8570);
and U8901 (N_8901,N_7612,N_7914);
or U8902 (N_8902,N_7673,N_8464);
and U8903 (N_8903,N_7752,N_8104);
and U8904 (N_8904,N_8482,N_8737);
xnor U8905 (N_8905,N_7927,N_8514);
and U8906 (N_8906,N_8541,N_8294);
and U8907 (N_8907,N_7813,N_7600);
or U8908 (N_8908,N_8000,N_8499);
and U8909 (N_8909,N_8351,N_8233);
nand U8910 (N_8910,N_7833,N_7587);
nand U8911 (N_8911,N_7588,N_8027);
nand U8912 (N_8912,N_8530,N_7854);
xnor U8913 (N_8913,N_7850,N_7862);
xnor U8914 (N_8914,N_7557,N_7737);
nand U8915 (N_8915,N_7846,N_8318);
and U8916 (N_8916,N_8049,N_8363);
nor U8917 (N_8917,N_7864,N_8034);
and U8918 (N_8918,N_8200,N_7646);
and U8919 (N_8919,N_8165,N_8558);
xnor U8920 (N_8920,N_7944,N_7828);
and U8921 (N_8921,N_8073,N_7637);
nand U8922 (N_8922,N_7649,N_8252);
or U8923 (N_8923,N_8305,N_8185);
nor U8924 (N_8924,N_8526,N_7762);
xor U8925 (N_8925,N_8218,N_8442);
nand U8926 (N_8926,N_7915,N_8193);
nand U8927 (N_8927,N_7732,N_8396);
nor U8928 (N_8928,N_8705,N_8427);
nor U8929 (N_8929,N_8523,N_7816);
and U8930 (N_8930,N_8444,N_7995);
or U8931 (N_8931,N_7878,N_7793);
and U8932 (N_8932,N_7852,N_8584);
and U8933 (N_8933,N_7542,N_7798);
or U8934 (N_8934,N_8145,N_8610);
xnor U8935 (N_8935,N_8282,N_7578);
xnor U8936 (N_8936,N_7900,N_8710);
and U8937 (N_8937,N_8688,N_8343);
nand U8938 (N_8938,N_8557,N_8001);
and U8939 (N_8939,N_8741,N_7976);
nor U8940 (N_8940,N_7742,N_7681);
nand U8941 (N_8941,N_8339,N_7781);
nor U8942 (N_8942,N_8322,N_7730);
xor U8943 (N_8943,N_8468,N_7647);
or U8944 (N_8944,N_8332,N_8219);
nand U8945 (N_8945,N_7514,N_7650);
nor U8946 (N_8946,N_8127,N_8581);
nand U8947 (N_8947,N_7782,N_8341);
nor U8948 (N_8948,N_8021,N_8395);
or U8949 (N_8949,N_7663,N_8392);
nand U8950 (N_8950,N_7535,N_7541);
or U8951 (N_8951,N_8357,N_8035);
nand U8952 (N_8952,N_7805,N_8249);
nand U8953 (N_8953,N_8687,N_8254);
and U8954 (N_8954,N_8651,N_8524);
nand U8955 (N_8955,N_8700,N_7872);
nand U8956 (N_8956,N_7998,N_7669);
nor U8957 (N_8957,N_8394,N_8559);
and U8958 (N_8958,N_8364,N_8555);
xnor U8959 (N_8959,N_8604,N_7939);
and U8960 (N_8960,N_7518,N_7690);
or U8961 (N_8961,N_7894,N_8646);
nand U8962 (N_8962,N_8668,N_7799);
nand U8963 (N_8963,N_8023,N_8130);
xor U8964 (N_8964,N_7567,N_8730);
nand U8965 (N_8965,N_8376,N_8594);
xnor U8966 (N_8966,N_8654,N_8008);
xnor U8967 (N_8967,N_7728,N_8116);
nand U8968 (N_8968,N_8652,N_7841);
or U8969 (N_8969,N_7710,N_8207);
and U8970 (N_8970,N_8208,N_8629);
and U8971 (N_8971,N_7524,N_8488);
xnor U8972 (N_8972,N_8215,N_7792);
or U8973 (N_8973,N_8211,N_7529);
xnor U8974 (N_8974,N_7599,N_8238);
nand U8975 (N_8975,N_7558,N_7656);
nor U8976 (N_8976,N_8072,N_7563);
nor U8977 (N_8977,N_7744,N_8744);
nand U8978 (N_8978,N_8005,N_8420);
nor U8979 (N_8979,N_7537,N_7877);
nor U8980 (N_8980,N_8714,N_8685);
nand U8981 (N_8981,N_7636,N_8076);
nand U8982 (N_8982,N_7565,N_8010);
nor U8983 (N_8983,N_8537,N_8565);
or U8984 (N_8984,N_8280,N_7718);
nor U8985 (N_8985,N_7968,N_8434);
nor U8986 (N_8986,N_7598,N_8626);
nor U8987 (N_8987,N_8566,N_8576);
and U8988 (N_8988,N_8289,N_8029);
nand U8989 (N_8989,N_8495,N_7511);
nand U8990 (N_8990,N_8198,N_8431);
xnor U8991 (N_8991,N_8648,N_8175);
nor U8992 (N_8992,N_8707,N_8184);
xnor U8993 (N_8993,N_8133,N_8733);
nor U8994 (N_8994,N_8411,N_7604);
nor U8995 (N_8995,N_8292,N_7789);
or U8996 (N_8996,N_8384,N_7820);
and U8997 (N_8997,N_7648,N_8053);
nor U8998 (N_8998,N_7571,N_8715);
or U8999 (N_8999,N_7855,N_7779);
or U9000 (N_9000,N_8403,N_8675);
and U9001 (N_9001,N_7662,N_8556);
and U9002 (N_9002,N_8622,N_8163);
or U9003 (N_9003,N_8662,N_7908);
and U9004 (N_9004,N_8333,N_7848);
nand U9005 (N_9005,N_8738,N_7879);
xnor U9006 (N_9006,N_8330,N_7840);
nand U9007 (N_9007,N_7640,N_8540);
nor U9008 (N_9008,N_8108,N_8288);
and U9009 (N_9009,N_8032,N_8577);
or U9010 (N_9010,N_8573,N_7590);
or U9011 (N_9011,N_7702,N_7684);
nand U9012 (N_9012,N_8650,N_8418);
xor U9013 (N_9013,N_8704,N_8720);
nor U9014 (N_9014,N_8349,N_7538);
xor U9015 (N_9015,N_8645,N_8272);
or U9016 (N_9016,N_8479,N_8013);
xnor U9017 (N_9017,N_7947,N_8123);
nor U9018 (N_9018,N_7513,N_8436);
and U9019 (N_9019,N_8387,N_8276);
nor U9020 (N_9020,N_8169,N_7961);
and U9021 (N_9021,N_7895,N_7838);
xor U9022 (N_9022,N_8362,N_8014);
or U9023 (N_9023,N_8255,N_7666);
nor U9024 (N_9024,N_8177,N_8382);
and U9025 (N_9025,N_7579,N_7745);
nor U9026 (N_9026,N_8439,N_8107);
and U9027 (N_9027,N_7753,N_7959);
and U9028 (N_9028,N_8593,N_7664);
nor U9029 (N_9029,N_7965,N_7523);
and U9030 (N_9030,N_8082,N_7929);
nor U9031 (N_9031,N_7996,N_8217);
nand U9032 (N_9032,N_7853,N_7791);
or U9033 (N_9033,N_7950,N_7508);
nand U9034 (N_9034,N_8025,N_8309);
and U9035 (N_9035,N_8518,N_8081);
or U9036 (N_9036,N_7531,N_8636);
or U9037 (N_9037,N_8727,N_8078);
or U9038 (N_9038,N_7500,N_8619);
nor U9039 (N_9039,N_8452,N_7644);
xnor U9040 (N_9040,N_8297,N_7689);
nor U9041 (N_9041,N_8732,N_8112);
and U9042 (N_9042,N_7577,N_8621);
and U9043 (N_9043,N_8342,N_8669);
nor U9044 (N_9044,N_8348,N_8549);
nor U9045 (N_9045,N_8703,N_7891);
and U9046 (N_9046,N_8447,N_8111);
and U9047 (N_9047,N_7629,N_8609);
nor U9048 (N_9048,N_8269,N_7780);
xor U9049 (N_9049,N_7901,N_7703);
nand U9050 (N_9050,N_8571,N_8587);
or U9051 (N_9051,N_8397,N_7992);
nand U9052 (N_9052,N_8500,N_8400);
and U9053 (N_9053,N_7633,N_7871);
nand U9054 (N_9054,N_8624,N_7921);
xor U9055 (N_9055,N_7540,N_8519);
and U9056 (N_9056,N_7607,N_8151);
xor U9057 (N_9057,N_8031,N_7860);
nand U9058 (N_9058,N_7760,N_8299);
or U9059 (N_9059,N_7835,N_8132);
or U9060 (N_9060,N_7694,N_8389);
nor U9061 (N_9061,N_7621,N_8298);
xnor U9062 (N_9062,N_7999,N_8421);
or U9063 (N_9063,N_7711,N_7594);
nor U9064 (N_9064,N_8140,N_7988);
nor U9065 (N_9065,N_8574,N_7688);
nand U9066 (N_9066,N_7569,N_8709);
and U9067 (N_9067,N_7888,N_8632);
nor U9068 (N_9068,N_8125,N_8459);
xor U9069 (N_9069,N_8152,N_7979);
xnor U9070 (N_9070,N_7706,N_7546);
nor U9071 (N_9071,N_8228,N_8290);
nand U9072 (N_9072,N_8399,N_7516);
nor U9073 (N_9073,N_8103,N_8516);
or U9074 (N_9074,N_7503,N_7754);
xor U9075 (N_9075,N_8696,N_7676);
or U9076 (N_9076,N_7949,N_7570);
xnor U9077 (N_9077,N_8037,N_7970);
or U9078 (N_9078,N_8188,N_7660);
nand U9079 (N_9079,N_8248,N_7620);
or U9080 (N_9080,N_8285,N_8390);
nand U9081 (N_9081,N_8644,N_8612);
or U9082 (N_9082,N_7708,N_7832);
xor U9083 (N_9083,N_8603,N_8409);
and U9084 (N_9084,N_8028,N_8096);
nand U9085 (N_9085,N_8458,N_8007);
nor U9086 (N_9086,N_7997,N_8678);
nor U9087 (N_9087,N_8578,N_8087);
or U9088 (N_9088,N_8267,N_8623);
or U9089 (N_9089,N_8692,N_8701);
nand U9090 (N_9090,N_8278,N_7756);
or U9091 (N_9091,N_7882,N_8437);
nor U9092 (N_9092,N_8582,N_8546);
xnor U9093 (N_9093,N_8615,N_8162);
nand U9094 (N_9094,N_8554,N_7960);
or U9095 (N_9095,N_7671,N_7551);
nor U9096 (N_9096,N_8012,N_8120);
nor U9097 (N_9097,N_8367,N_7683);
nand U9098 (N_9098,N_8039,N_8706);
and U9099 (N_9099,N_8115,N_7759);
or U9100 (N_9100,N_8474,N_8572);
or U9101 (N_9101,N_8160,N_8545);
and U9102 (N_9102,N_7721,N_7719);
nand U9103 (N_9103,N_8265,N_7734);
nand U9104 (N_9104,N_7844,N_7896);
nor U9105 (N_9105,N_7631,N_8469);
xnor U9106 (N_9106,N_8234,N_8243);
nor U9107 (N_9107,N_7555,N_7716);
nand U9108 (N_9108,N_7962,N_8095);
or U9109 (N_9109,N_7643,N_8617);
or U9110 (N_9110,N_8717,N_7547);
or U9111 (N_9111,N_8492,N_8063);
and U9112 (N_9112,N_7790,N_8251);
xnor U9113 (N_9113,N_8083,N_7758);
or U9114 (N_9114,N_8728,N_7972);
nor U9115 (N_9115,N_7769,N_8521);
xor U9116 (N_9116,N_7738,N_8202);
nor U9117 (N_9117,N_7755,N_7966);
nand U9118 (N_9118,N_7739,N_7642);
or U9119 (N_9119,N_7586,N_8637);
nand U9120 (N_9120,N_8203,N_8536);
nor U9121 (N_9121,N_7810,N_7724);
or U9122 (N_9122,N_7881,N_8199);
or U9123 (N_9123,N_8126,N_7956);
nor U9124 (N_9124,N_8630,N_8110);
nor U9125 (N_9125,N_7899,N_8429);
or U9126 (N_9126,N_7943,N_8293);
and U9127 (N_9127,N_7559,N_7796);
xnor U9128 (N_9128,N_7830,N_8273);
xor U9129 (N_9129,N_8378,N_7770);
nand U9130 (N_9130,N_8311,N_7971);
xnor U9131 (N_9131,N_8494,N_7526);
or U9132 (N_9132,N_7543,N_8602);
nand U9133 (N_9133,N_8258,N_8391);
nor U9134 (N_9134,N_7767,N_8398);
nor U9135 (N_9135,N_7928,N_7861);
nand U9136 (N_9136,N_7618,N_7748);
nor U9137 (N_9137,N_8676,N_8075);
or U9138 (N_9138,N_8561,N_8695);
or U9139 (N_9139,N_7685,N_8122);
xnor U9140 (N_9140,N_8625,N_8412);
nand U9141 (N_9141,N_7603,N_7534);
nand U9142 (N_9142,N_8262,N_7836);
or U9143 (N_9143,N_7585,N_8061);
or U9144 (N_9144,N_7977,N_8641);
nor U9145 (N_9145,N_7624,N_7580);
xor U9146 (N_9146,N_7857,N_8253);
and U9147 (N_9147,N_8047,N_8227);
or U9148 (N_9148,N_7686,N_8408);
or U9149 (N_9149,N_7677,N_8174);
xor U9150 (N_9150,N_8331,N_8699);
or U9151 (N_9151,N_7700,N_8307);
or U9152 (N_9152,N_8139,N_8501);
nand U9153 (N_9153,N_8170,N_8749);
nand U9154 (N_9154,N_8306,N_8746);
nor U9155 (N_9155,N_7613,N_7775);
and U9156 (N_9156,N_7794,N_8279);
or U9157 (N_9157,N_8440,N_8338);
nand U9158 (N_9158,N_8532,N_8680);
nand U9159 (N_9159,N_8080,N_8689);
xor U9160 (N_9160,N_7615,N_8547);
xnor U9161 (N_9161,N_7574,N_7890);
and U9162 (N_9162,N_7913,N_7668);
or U9163 (N_9163,N_7948,N_8731);
or U9164 (N_9164,N_8542,N_8489);
or U9165 (N_9165,N_8534,N_8522);
nand U9166 (N_9166,N_8329,N_7863);
xnor U9167 (N_9167,N_8304,N_8229);
nor U9168 (N_9168,N_8209,N_7815);
nor U9169 (N_9169,N_7581,N_8481);
xor U9170 (N_9170,N_8383,N_8283);
and U9171 (N_9171,N_8473,N_7610);
or U9172 (N_9172,N_7842,N_8484);
xnor U9173 (N_9173,N_7937,N_7773);
xnor U9174 (N_9174,N_7936,N_7889);
or U9175 (N_9175,N_7990,N_8423);
nand U9176 (N_9176,N_8375,N_7898);
nor U9177 (N_9177,N_7741,N_8564);
nor U9178 (N_9178,N_7757,N_7884);
nor U9179 (N_9179,N_8598,N_8016);
nor U9180 (N_9180,N_7674,N_8600);
nand U9181 (N_9181,N_7817,N_8220);
or U9182 (N_9182,N_7892,N_8487);
or U9183 (N_9183,N_7873,N_8109);
nand U9184 (N_9184,N_8608,N_8144);
or U9185 (N_9185,N_8443,N_7504);
or U9186 (N_9186,N_7679,N_8681);
xnor U9187 (N_9187,N_8060,N_8121);
nand U9188 (N_9188,N_8084,N_7918);
and U9189 (N_9189,N_8386,N_7682);
xnor U9190 (N_9190,N_8413,N_8141);
nor U9191 (N_9191,N_8045,N_8527);
nand U9192 (N_9192,N_8496,N_8451);
and U9193 (N_9193,N_8354,N_7731);
xnor U9194 (N_9194,N_8401,N_7945);
xor U9195 (N_9195,N_7788,N_8454);
or U9196 (N_9196,N_7729,N_7614);
and U9197 (N_9197,N_7787,N_8221);
xnor U9198 (N_9198,N_8377,N_8725);
nor U9199 (N_9199,N_7942,N_7726);
nand U9200 (N_9200,N_8665,N_7818);
nor U9201 (N_9201,N_7911,N_7764);
nand U9202 (N_9202,N_8070,N_8435);
and U9203 (N_9203,N_7725,N_8734);
nand U9204 (N_9204,N_7974,N_8224);
nor U9205 (N_9205,N_8667,N_7522);
and U9206 (N_9206,N_8414,N_8191);
and U9207 (N_9207,N_7678,N_8531);
nand U9208 (N_9208,N_7776,N_8052);
nor U9209 (N_9209,N_8131,N_8467);
and U9210 (N_9210,N_8077,N_7783);
nor U9211 (N_9211,N_8589,N_8241);
nor U9212 (N_9212,N_8729,N_7530);
and U9213 (N_9213,N_8684,N_7827);
and U9214 (N_9214,N_8009,N_7938);
nand U9215 (N_9215,N_8068,N_7606);
and U9216 (N_9216,N_7897,N_8101);
nor U9217 (N_9217,N_8407,N_8230);
nor U9218 (N_9218,N_7975,N_8090);
xnor U9219 (N_9219,N_7797,N_7589);
xnor U9220 (N_9220,N_8419,N_7957);
and U9221 (N_9221,N_8065,N_8712);
or U9222 (N_9222,N_8171,N_8446);
nand U9223 (N_9223,N_7876,N_8226);
xor U9224 (N_9224,N_7867,N_7986);
nor U9225 (N_9225,N_8448,N_8661);
nand U9226 (N_9226,N_7973,N_8716);
nand U9227 (N_9227,N_8189,N_8033);
or U9228 (N_9228,N_8195,N_7596);
and U9229 (N_9229,N_7701,N_8312);
or U9230 (N_9230,N_7653,N_8483);
nand U9231 (N_9231,N_8179,N_8300);
xor U9232 (N_9232,N_8415,N_7727);
and U9233 (N_9233,N_8369,N_8585);
nor U9234 (N_9234,N_7627,N_7593);
nor U9235 (N_9235,N_7532,N_8327);
nand U9236 (N_9236,N_8091,N_8410);
nand U9237 (N_9237,N_7964,N_8026);
nand U9238 (N_9238,N_8430,N_7687);
or U9239 (N_9239,N_7622,N_8583);
or U9240 (N_9240,N_7925,N_8682);
nor U9241 (N_9241,N_7693,N_8424);
or U9242 (N_9242,N_8457,N_8019);
and U9243 (N_9243,N_8595,N_7766);
xor U9244 (N_9244,N_8240,N_7695);
or U9245 (N_9245,N_8404,N_8261);
nand U9246 (N_9246,N_7723,N_8310);
nor U9247 (N_9247,N_7761,N_7717);
nor U9248 (N_9248,N_8493,N_7849);
and U9249 (N_9249,N_8317,N_7808);
or U9250 (N_9250,N_7575,N_8352);
nand U9251 (N_9251,N_8149,N_8486);
nor U9252 (N_9252,N_8148,N_8345);
and U9253 (N_9253,N_7958,N_7819);
and U9254 (N_9254,N_8478,N_8136);
or U9255 (N_9255,N_7980,N_7907);
nor U9256 (N_9256,N_8640,N_7605);
and U9257 (N_9257,N_7670,N_7856);
xnor U9258 (N_9258,N_8620,N_7883);
nand U9259 (N_9259,N_7984,N_8461);
xnor U9260 (N_9260,N_7906,N_8286);
and U9261 (N_9261,N_8385,N_7525);
nand U9262 (N_9262,N_8092,N_7875);
nor U9263 (N_9263,N_8591,N_7652);
nand U9264 (N_9264,N_8463,N_7981);
or U9265 (N_9265,N_7584,N_7549);
xnor U9266 (N_9266,N_8592,N_8393);
nand U9267 (N_9267,N_8142,N_8058);
nand U9268 (N_9268,N_8050,N_8748);
nor U9269 (N_9269,N_8613,N_7765);
nor U9270 (N_9270,N_8155,N_8271);
nand U9271 (N_9271,N_8041,N_7946);
or U9272 (N_9272,N_8340,N_8214);
nor U9273 (N_9273,N_7916,N_8181);
and U9274 (N_9274,N_8353,N_8579);
xnor U9275 (N_9275,N_7582,N_7807);
nor U9276 (N_9276,N_8506,N_7829);
xor U9277 (N_9277,N_7851,N_8054);
xor U9278 (N_9278,N_8239,N_7714);
or U9279 (N_9279,N_8062,N_8548);
or U9280 (N_9280,N_8462,N_8606);
nand U9281 (N_9281,N_8512,N_8663);
nor U9282 (N_9282,N_8405,N_8046);
xor U9283 (N_9283,N_7989,N_8143);
nor U9284 (N_9284,N_8693,N_8003);
nand U9285 (N_9285,N_7512,N_8302);
or U9286 (N_9286,N_7812,N_7763);
or U9287 (N_9287,N_8736,N_7845);
or U9288 (N_9288,N_8551,N_8315);
and U9289 (N_9289,N_7698,N_8161);
or U9290 (N_9290,N_7539,N_8465);
xor U9291 (N_9291,N_8335,N_7651);
and U9292 (N_9292,N_7987,N_7697);
xnor U9293 (N_9293,N_7886,N_8277);
and U9294 (N_9294,N_7887,N_8183);
and U9295 (N_9295,N_8513,N_8525);
or U9296 (N_9296,N_7751,N_7931);
nand U9297 (N_9297,N_8274,N_7573);
and U9298 (N_9298,N_8264,N_8154);
nand U9299 (N_9299,N_7885,N_8718);
xor U9300 (N_9300,N_8231,N_7501);
nand U9301 (N_9301,N_8432,N_7924);
xor U9302 (N_9302,N_8504,N_7955);
xnor U9303 (N_9303,N_8428,N_8067);
nor U9304 (N_9304,N_8085,N_7940);
nor U9305 (N_9305,N_8259,N_8002);
xnor U9306 (N_9306,N_8319,N_8505);
nand U9307 (N_9307,N_8138,N_7665);
nand U9308 (N_9308,N_8316,N_8599);
nand U9309 (N_9309,N_7869,N_8350);
nand U9310 (N_9310,N_7509,N_8497);
nor U9311 (N_9311,N_8071,N_8284);
and U9312 (N_9312,N_8586,N_7837);
nor U9313 (N_9313,N_8666,N_8245);
xor U9314 (N_9314,N_8517,N_8303);
xnor U9315 (N_9315,N_8346,N_7922);
or U9316 (N_9316,N_8323,N_8222);
or U9317 (N_9317,N_8460,N_8114);
nand U9318 (N_9318,N_7630,N_8373);
xor U9319 (N_9319,N_8256,N_8638);
nor U9320 (N_9320,N_8201,N_8066);
xor U9321 (N_9321,N_8433,N_8372);
xor U9322 (N_9322,N_7536,N_7611);
nand U9323 (N_9323,N_7740,N_8466);
and U9324 (N_9324,N_7675,N_8677);
and U9325 (N_9325,N_8719,N_8291);
or U9326 (N_9326,N_8425,N_7510);
or U9327 (N_9327,N_7550,N_8038);
xnor U9328 (N_9328,N_8721,N_8520);
or U9329 (N_9329,N_8723,N_8135);
xnor U9330 (N_9330,N_8146,N_7720);
and U9331 (N_9331,N_8178,N_8450);
or U9332 (N_9332,N_7953,N_7616);
and U9333 (N_9333,N_8308,N_8232);
xor U9334 (N_9334,N_7795,N_8417);
nand U9335 (N_9335,N_8607,N_7806);
or U9336 (N_9336,N_8562,N_7800);
xor U9337 (N_9337,N_8247,N_8205);
or U9338 (N_9338,N_7826,N_7592);
nand U9339 (N_9339,N_8374,N_8336);
nand U9340 (N_9340,N_7712,N_7572);
and U9341 (N_9341,N_8445,N_8575);
or U9342 (N_9342,N_7680,N_7859);
and U9343 (N_9343,N_8535,N_8538);
nor U9344 (N_9344,N_8069,N_8628);
xnor U9345 (N_9345,N_7880,N_7735);
or U9346 (N_9346,N_8656,N_7803);
or U9347 (N_9347,N_8370,N_8553);
xor U9348 (N_9348,N_8490,N_7903);
nand U9349 (N_9349,N_8366,N_8438);
nor U9350 (N_9350,N_7704,N_7746);
or U9351 (N_9351,N_7713,N_7822);
nand U9352 (N_9352,N_8118,N_8176);
nand U9353 (N_9353,N_7658,N_8270);
xnor U9354 (N_9354,N_8627,N_8674);
xnor U9355 (N_9355,N_8064,N_7736);
nor U9356 (N_9356,N_7608,N_7969);
or U9357 (N_9357,N_8742,N_8100);
nor U9358 (N_9358,N_8020,N_8471);
xor U9359 (N_9359,N_7952,N_7858);
and U9360 (N_9360,N_8074,N_8275);
nand U9361 (N_9361,N_7699,N_7645);
and U9362 (N_9362,N_7874,N_7771);
xnor U9363 (N_9363,N_8470,N_8040);
nand U9364 (N_9364,N_7809,N_7834);
and U9365 (N_9365,N_8533,N_8735);
xnor U9366 (N_9366,N_8089,N_7545);
nor U9367 (N_9367,N_7941,N_7743);
xnor U9368 (N_9368,N_7623,N_8326);
xor U9369 (N_9369,N_8213,N_8190);
nand U9370 (N_9370,N_8320,N_8616);
and U9371 (N_9371,N_8455,N_8380);
xnor U9372 (N_9372,N_7609,N_7954);
and U9373 (N_9373,N_8611,N_7831);
xnor U9374 (N_9374,N_8550,N_8381);
nor U9375 (N_9375,N_8313,N_8662);
xor U9376 (N_9376,N_7902,N_8014);
and U9377 (N_9377,N_8642,N_8254);
xnor U9378 (N_9378,N_8210,N_8232);
nand U9379 (N_9379,N_7907,N_7933);
nor U9380 (N_9380,N_8481,N_8037);
and U9381 (N_9381,N_8289,N_8726);
or U9382 (N_9382,N_8692,N_8169);
nand U9383 (N_9383,N_8021,N_7865);
and U9384 (N_9384,N_8281,N_7548);
or U9385 (N_9385,N_8574,N_8176);
xor U9386 (N_9386,N_7702,N_7649);
or U9387 (N_9387,N_8214,N_8582);
and U9388 (N_9388,N_8393,N_7758);
nor U9389 (N_9389,N_8342,N_7916);
xor U9390 (N_9390,N_8075,N_7718);
xnor U9391 (N_9391,N_7942,N_7779);
or U9392 (N_9392,N_8101,N_8486);
nor U9393 (N_9393,N_7604,N_8295);
and U9394 (N_9394,N_7598,N_7980);
and U9395 (N_9395,N_7673,N_7566);
nand U9396 (N_9396,N_7536,N_8008);
nand U9397 (N_9397,N_7897,N_8533);
and U9398 (N_9398,N_8227,N_8112);
or U9399 (N_9399,N_7919,N_8041);
xor U9400 (N_9400,N_8380,N_7836);
or U9401 (N_9401,N_7788,N_7568);
or U9402 (N_9402,N_7868,N_7793);
and U9403 (N_9403,N_7724,N_8586);
and U9404 (N_9404,N_8533,N_7878);
and U9405 (N_9405,N_8032,N_8405);
or U9406 (N_9406,N_7943,N_8149);
and U9407 (N_9407,N_8211,N_7966);
xnor U9408 (N_9408,N_7828,N_7855);
xor U9409 (N_9409,N_7637,N_8311);
or U9410 (N_9410,N_8176,N_8036);
or U9411 (N_9411,N_8554,N_7734);
nand U9412 (N_9412,N_7736,N_8426);
nand U9413 (N_9413,N_8623,N_8643);
nand U9414 (N_9414,N_7885,N_7676);
or U9415 (N_9415,N_8735,N_7859);
nand U9416 (N_9416,N_8143,N_8089);
nand U9417 (N_9417,N_8032,N_8647);
and U9418 (N_9418,N_7577,N_8721);
or U9419 (N_9419,N_8572,N_8041);
nand U9420 (N_9420,N_8559,N_8296);
and U9421 (N_9421,N_7625,N_8688);
or U9422 (N_9422,N_8106,N_7930);
or U9423 (N_9423,N_8225,N_8261);
nand U9424 (N_9424,N_7707,N_8295);
nor U9425 (N_9425,N_8109,N_7897);
xor U9426 (N_9426,N_8190,N_7604);
nor U9427 (N_9427,N_8581,N_7702);
and U9428 (N_9428,N_8503,N_8460);
nand U9429 (N_9429,N_8155,N_8127);
and U9430 (N_9430,N_7541,N_8574);
and U9431 (N_9431,N_7757,N_7978);
or U9432 (N_9432,N_7777,N_8429);
nand U9433 (N_9433,N_7796,N_8528);
xnor U9434 (N_9434,N_8629,N_7873);
nor U9435 (N_9435,N_8617,N_7565);
nand U9436 (N_9436,N_8392,N_8297);
or U9437 (N_9437,N_8676,N_7500);
nand U9438 (N_9438,N_8124,N_8519);
nor U9439 (N_9439,N_7620,N_8680);
and U9440 (N_9440,N_7734,N_8031);
nor U9441 (N_9441,N_8570,N_7877);
and U9442 (N_9442,N_8646,N_8102);
or U9443 (N_9443,N_7910,N_8251);
nor U9444 (N_9444,N_8467,N_8261);
nor U9445 (N_9445,N_7676,N_7843);
nor U9446 (N_9446,N_8023,N_8019);
nand U9447 (N_9447,N_8072,N_8062);
nor U9448 (N_9448,N_7564,N_7714);
xor U9449 (N_9449,N_8292,N_7875);
xor U9450 (N_9450,N_8267,N_8011);
or U9451 (N_9451,N_8537,N_7630);
or U9452 (N_9452,N_7923,N_8593);
or U9453 (N_9453,N_8110,N_8552);
xor U9454 (N_9454,N_8089,N_7662);
nand U9455 (N_9455,N_8244,N_7843);
xnor U9456 (N_9456,N_7885,N_7563);
or U9457 (N_9457,N_7886,N_7864);
nand U9458 (N_9458,N_7904,N_8308);
nor U9459 (N_9459,N_8571,N_8522);
nor U9460 (N_9460,N_8640,N_8657);
and U9461 (N_9461,N_8156,N_8407);
and U9462 (N_9462,N_7598,N_8034);
nand U9463 (N_9463,N_8627,N_8051);
and U9464 (N_9464,N_8703,N_8602);
or U9465 (N_9465,N_8689,N_8023);
nor U9466 (N_9466,N_7711,N_7520);
xor U9467 (N_9467,N_8205,N_7713);
nand U9468 (N_9468,N_8538,N_8327);
and U9469 (N_9469,N_7643,N_8413);
nand U9470 (N_9470,N_8494,N_8068);
nor U9471 (N_9471,N_8438,N_7955);
nor U9472 (N_9472,N_8495,N_8643);
nand U9473 (N_9473,N_7822,N_7897);
nor U9474 (N_9474,N_8058,N_8459);
nand U9475 (N_9475,N_8444,N_7989);
nand U9476 (N_9476,N_8213,N_8525);
nand U9477 (N_9477,N_8171,N_8629);
xor U9478 (N_9478,N_7937,N_7717);
nor U9479 (N_9479,N_7986,N_8591);
or U9480 (N_9480,N_7691,N_8360);
nor U9481 (N_9481,N_7831,N_7846);
xnor U9482 (N_9482,N_8126,N_8111);
and U9483 (N_9483,N_7671,N_8385);
nor U9484 (N_9484,N_7839,N_7714);
nor U9485 (N_9485,N_7556,N_8564);
and U9486 (N_9486,N_7830,N_8209);
and U9487 (N_9487,N_8458,N_8009);
and U9488 (N_9488,N_7501,N_7825);
nor U9489 (N_9489,N_7648,N_8146);
or U9490 (N_9490,N_8177,N_7814);
xnor U9491 (N_9491,N_8487,N_8659);
or U9492 (N_9492,N_7630,N_7883);
nand U9493 (N_9493,N_7861,N_7947);
nor U9494 (N_9494,N_7963,N_8679);
and U9495 (N_9495,N_8114,N_7800);
and U9496 (N_9496,N_8104,N_8156);
or U9497 (N_9497,N_8461,N_8041);
and U9498 (N_9498,N_8643,N_8449);
xor U9499 (N_9499,N_7709,N_7642);
and U9500 (N_9500,N_8655,N_7923);
nor U9501 (N_9501,N_7503,N_8696);
and U9502 (N_9502,N_8077,N_7978);
nand U9503 (N_9503,N_7789,N_8277);
nor U9504 (N_9504,N_8434,N_8641);
nor U9505 (N_9505,N_7878,N_8433);
or U9506 (N_9506,N_8402,N_7727);
nand U9507 (N_9507,N_8148,N_8057);
nand U9508 (N_9508,N_7569,N_8613);
nor U9509 (N_9509,N_8244,N_8216);
nand U9510 (N_9510,N_7639,N_7782);
or U9511 (N_9511,N_8107,N_8492);
nor U9512 (N_9512,N_7626,N_8482);
nand U9513 (N_9513,N_8053,N_8607);
and U9514 (N_9514,N_7889,N_7916);
and U9515 (N_9515,N_7844,N_8582);
or U9516 (N_9516,N_7521,N_8664);
and U9517 (N_9517,N_7651,N_8007);
xor U9518 (N_9518,N_8408,N_8667);
and U9519 (N_9519,N_8697,N_8549);
xor U9520 (N_9520,N_7581,N_7717);
nand U9521 (N_9521,N_8447,N_8043);
or U9522 (N_9522,N_7662,N_8679);
and U9523 (N_9523,N_8674,N_8649);
xnor U9524 (N_9524,N_8719,N_8445);
xor U9525 (N_9525,N_7926,N_7965);
and U9526 (N_9526,N_8189,N_8556);
or U9527 (N_9527,N_7815,N_8065);
nor U9528 (N_9528,N_8167,N_8096);
nand U9529 (N_9529,N_8730,N_7642);
nor U9530 (N_9530,N_7717,N_7966);
xnor U9531 (N_9531,N_7923,N_7655);
xor U9532 (N_9532,N_7606,N_7723);
nor U9533 (N_9533,N_8594,N_7509);
xor U9534 (N_9534,N_8426,N_7608);
nor U9535 (N_9535,N_8560,N_7642);
or U9536 (N_9536,N_7946,N_8315);
and U9537 (N_9537,N_8001,N_8368);
nor U9538 (N_9538,N_7654,N_8331);
nand U9539 (N_9539,N_8624,N_8276);
or U9540 (N_9540,N_8318,N_8529);
and U9541 (N_9541,N_8393,N_8283);
and U9542 (N_9542,N_7654,N_8164);
or U9543 (N_9543,N_8010,N_7777);
xor U9544 (N_9544,N_7566,N_7954);
xnor U9545 (N_9545,N_7806,N_8177);
or U9546 (N_9546,N_8127,N_8579);
and U9547 (N_9547,N_8449,N_8583);
and U9548 (N_9548,N_7538,N_8211);
xnor U9549 (N_9549,N_8695,N_8253);
xor U9550 (N_9550,N_7886,N_7973);
nand U9551 (N_9551,N_8027,N_8481);
xnor U9552 (N_9552,N_7808,N_7687);
nor U9553 (N_9553,N_7808,N_8487);
nand U9554 (N_9554,N_8321,N_7805);
nand U9555 (N_9555,N_7818,N_8418);
nor U9556 (N_9556,N_8625,N_7604);
xor U9557 (N_9557,N_8077,N_7797);
nand U9558 (N_9558,N_7764,N_7599);
or U9559 (N_9559,N_7659,N_7918);
nand U9560 (N_9560,N_7780,N_8445);
or U9561 (N_9561,N_7671,N_8356);
nor U9562 (N_9562,N_8203,N_7904);
xnor U9563 (N_9563,N_8599,N_7794);
nor U9564 (N_9564,N_7839,N_8127);
nor U9565 (N_9565,N_8563,N_8655);
nor U9566 (N_9566,N_8024,N_7638);
or U9567 (N_9567,N_7637,N_8465);
nor U9568 (N_9568,N_7711,N_8557);
or U9569 (N_9569,N_7820,N_8571);
and U9570 (N_9570,N_7670,N_7693);
and U9571 (N_9571,N_7997,N_8488);
and U9572 (N_9572,N_8508,N_8185);
and U9573 (N_9573,N_8283,N_8305);
nand U9574 (N_9574,N_7686,N_8062);
nand U9575 (N_9575,N_8696,N_8185);
or U9576 (N_9576,N_7739,N_7800);
nand U9577 (N_9577,N_8571,N_8419);
nand U9578 (N_9578,N_7895,N_8147);
or U9579 (N_9579,N_7859,N_8640);
and U9580 (N_9580,N_8568,N_7624);
and U9581 (N_9581,N_7503,N_8255);
and U9582 (N_9582,N_8503,N_7772);
xor U9583 (N_9583,N_7656,N_7863);
nor U9584 (N_9584,N_8699,N_8578);
nand U9585 (N_9585,N_7950,N_8279);
xor U9586 (N_9586,N_8735,N_7561);
xor U9587 (N_9587,N_8393,N_8107);
or U9588 (N_9588,N_8349,N_8517);
and U9589 (N_9589,N_7812,N_8648);
or U9590 (N_9590,N_7710,N_8321);
or U9591 (N_9591,N_8707,N_8518);
or U9592 (N_9592,N_7581,N_8532);
nand U9593 (N_9593,N_8085,N_7523);
nor U9594 (N_9594,N_8175,N_7628);
nor U9595 (N_9595,N_8715,N_8446);
nor U9596 (N_9596,N_8019,N_8270);
or U9597 (N_9597,N_8716,N_8631);
nand U9598 (N_9598,N_8182,N_7583);
xnor U9599 (N_9599,N_7724,N_7850);
xor U9600 (N_9600,N_8478,N_7606);
nor U9601 (N_9601,N_7792,N_7771);
xnor U9602 (N_9602,N_7747,N_7849);
or U9603 (N_9603,N_7642,N_7536);
nor U9604 (N_9604,N_7586,N_7736);
nand U9605 (N_9605,N_7842,N_8261);
and U9606 (N_9606,N_8534,N_7805);
nand U9607 (N_9607,N_8393,N_8367);
nand U9608 (N_9608,N_8727,N_8089);
and U9609 (N_9609,N_8367,N_8419);
nand U9610 (N_9610,N_8711,N_8505);
xnor U9611 (N_9611,N_7828,N_7883);
or U9612 (N_9612,N_8549,N_7621);
xor U9613 (N_9613,N_7846,N_8051);
and U9614 (N_9614,N_8357,N_8582);
and U9615 (N_9615,N_8078,N_8287);
or U9616 (N_9616,N_7686,N_8489);
nand U9617 (N_9617,N_7634,N_8126);
nand U9618 (N_9618,N_7609,N_8161);
xnor U9619 (N_9619,N_8094,N_7797);
or U9620 (N_9620,N_8570,N_8410);
nand U9621 (N_9621,N_8604,N_8208);
nand U9622 (N_9622,N_8049,N_8566);
or U9623 (N_9623,N_7597,N_8567);
xor U9624 (N_9624,N_7882,N_7926);
xor U9625 (N_9625,N_8033,N_8488);
or U9626 (N_9626,N_8404,N_8565);
and U9627 (N_9627,N_8299,N_7844);
nand U9628 (N_9628,N_7876,N_8143);
nor U9629 (N_9629,N_7926,N_7860);
nand U9630 (N_9630,N_8330,N_7567);
or U9631 (N_9631,N_8268,N_8194);
or U9632 (N_9632,N_8535,N_8667);
xor U9633 (N_9633,N_8335,N_7647);
xor U9634 (N_9634,N_7523,N_8136);
nand U9635 (N_9635,N_8668,N_8317);
and U9636 (N_9636,N_7697,N_8403);
nand U9637 (N_9637,N_8019,N_7624);
and U9638 (N_9638,N_8633,N_8695);
xor U9639 (N_9639,N_7768,N_7591);
and U9640 (N_9640,N_7893,N_8504);
nand U9641 (N_9641,N_8172,N_8127);
nand U9642 (N_9642,N_7931,N_8719);
xnor U9643 (N_9643,N_7938,N_7879);
xor U9644 (N_9644,N_8484,N_8225);
nor U9645 (N_9645,N_8068,N_8206);
or U9646 (N_9646,N_8321,N_8581);
and U9647 (N_9647,N_8435,N_7766);
nand U9648 (N_9648,N_7617,N_8413);
xor U9649 (N_9649,N_7524,N_7805);
xor U9650 (N_9650,N_8446,N_7512);
or U9651 (N_9651,N_7967,N_7987);
nor U9652 (N_9652,N_8009,N_8187);
and U9653 (N_9653,N_7952,N_8398);
nand U9654 (N_9654,N_7779,N_8594);
and U9655 (N_9655,N_7825,N_8746);
and U9656 (N_9656,N_7683,N_8606);
nand U9657 (N_9657,N_8161,N_7670);
nor U9658 (N_9658,N_7527,N_7676);
or U9659 (N_9659,N_7635,N_7934);
and U9660 (N_9660,N_8241,N_8258);
and U9661 (N_9661,N_7811,N_7779);
nand U9662 (N_9662,N_7845,N_8501);
xor U9663 (N_9663,N_8115,N_7667);
nand U9664 (N_9664,N_7795,N_7986);
nor U9665 (N_9665,N_8115,N_7669);
or U9666 (N_9666,N_8485,N_8500);
nand U9667 (N_9667,N_7810,N_7845);
nand U9668 (N_9668,N_7907,N_8159);
nand U9669 (N_9669,N_7601,N_8253);
nor U9670 (N_9670,N_8200,N_7973);
or U9671 (N_9671,N_7879,N_7683);
xnor U9672 (N_9672,N_8095,N_8651);
xnor U9673 (N_9673,N_7800,N_8352);
xnor U9674 (N_9674,N_8077,N_8329);
nor U9675 (N_9675,N_7689,N_7735);
xor U9676 (N_9676,N_8345,N_8154);
nor U9677 (N_9677,N_8607,N_8739);
nand U9678 (N_9678,N_7923,N_8553);
nor U9679 (N_9679,N_8521,N_8449);
nand U9680 (N_9680,N_7995,N_8035);
xor U9681 (N_9681,N_7762,N_7928);
or U9682 (N_9682,N_8707,N_7659);
nor U9683 (N_9683,N_7898,N_7823);
or U9684 (N_9684,N_7560,N_7801);
xnor U9685 (N_9685,N_8539,N_8512);
or U9686 (N_9686,N_7660,N_7693);
or U9687 (N_9687,N_7899,N_8422);
or U9688 (N_9688,N_8672,N_8642);
or U9689 (N_9689,N_8264,N_8523);
and U9690 (N_9690,N_7922,N_7615);
nor U9691 (N_9691,N_8394,N_7634);
or U9692 (N_9692,N_7595,N_8602);
and U9693 (N_9693,N_8056,N_7824);
nand U9694 (N_9694,N_8438,N_8251);
and U9695 (N_9695,N_7607,N_7715);
nor U9696 (N_9696,N_7926,N_8134);
nor U9697 (N_9697,N_7919,N_8198);
or U9698 (N_9698,N_8513,N_8510);
and U9699 (N_9699,N_8676,N_8094);
and U9700 (N_9700,N_8695,N_8278);
xor U9701 (N_9701,N_8515,N_7752);
or U9702 (N_9702,N_8141,N_7507);
or U9703 (N_9703,N_8015,N_7725);
nor U9704 (N_9704,N_8061,N_8256);
nor U9705 (N_9705,N_8518,N_7519);
and U9706 (N_9706,N_8296,N_8625);
nand U9707 (N_9707,N_7895,N_8144);
nor U9708 (N_9708,N_7646,N_8265);
and U9709 (N_9709,N_8313,N_7897);
nand U9710 (N_9710,N_7797,N_8162);
or U9711 (N_9711,N_8168,N_7842);
xor U9712 (N_9712,N_7586,N_8514);
and U9713 (N_9713,N_8220,N_8376);
nor U9714 (N_9714,N_8479,N_8043);
xor U9715 (N_9715,N_8155,N_7925);
nand U9716 (N_9716,N_7874,N_7831);
and U9717 (N_9717,N_8091,N_7834);
nand U9718 (N_9718,N_7829,N_8653);
or U9719 (N_9719,N_8740,N_8678);
nand U9720 (N_9720,N_7796,N_8207);
or U9721 (N_9721,N_8543,N_8134);
nand U9722 (N_9722,N_8091,N_7844);
and U9723 (N_9723,N_8260,N_7848);
nor U9724 (N_9724,N_8500,N_8300);
nand U9725 (N_9725,N_8403,N_8192);
and U9726 (N_9726,N_8736,N_8607);
xnor U9727 (N_9727,N_8398,N_8738);
or U9728 (N_9728,N_8178,N_8383);
xnor U9729 (N_9729,N_7615,N_8586);
nand U9730 (N_9730,N_8211,N_8006);
or U9731 (N_9731,N_8070,N_8469);
xnor U9732 (N_9732,N_8744,N_8683);
nand U9733 (N_9733,N_8066,N_8746);
nor U9734 (N_9734,N_8170,N_8528);
xor U9735 (N_9735,N_8431,N_8329);
and U9736 (N_9736,N_8642,N_8643);
nand U9737 (N_9737,N_7976,N_8109);
or U9738 (N_9738,N_7745,N_7707);
xnor U9739 (N_9739,N_8384,N_8558);
nor U9740 (N_9740,N_8664,N_8112);
or U9741 (N_9741,N_8654,N_7854);
nor U9742 (N_9742,N_7606,N_7994);
or U9743 (N_9743,N_8666,N_8561);
nor U9744 (N_9744,N_8384,N_8738);
nand U9745 (N_9745,N_8704,N_7618);
and U9746 (N_9746,N_8225,N_8577);
and U9747 (N_9747,N_8191,N_8569);
and U9748 (N_9748,N_8679,N_8301);
or U9749 (N_9749,N_7594,N_8547);
xnor U9750 (N_9750,N_8156,N_7891);
xor U9751 (N_9751,N_8459,N_8212);
nor U9752 (N_9752,N_7683,N_7749);
nand U9753 (N_9753,N_7820,N_8256);
nor U9754 (N_9754,N_8503,N_8179);
xor U9755 (N_9755,N_7642,N_8101);
nand U9756 (N_9756,N_8109,N_8296);
nand U9757 (N_9757,N_8530,N_8447);
xnor U9758 (N_9758,N_8107,N_8218);
nor U9759 (N_9759,N_8203,N_7558);
nor U9760 (N_9760,N_8234,N_7516);
or U9761 (N_9761,N_8745,N_7720);
nor U9762 (N_9762,N_7774,N_8341);
and U9763 (N_9763,N_8491,N_7938);
or U9764 (N_9764,N_8199,N_8304);
or U9765 (N_9765,N_8738,N_8355);
or U9766 (N_9766,N_8030,N_7943);
and U9767 (N_9767,N_7917,N_7931);
nand U9768 (N_9768,N_8372,N_8596);
nand U9769 (N_9769,N_8293,N_8747);
or U9770 (N_9770,N_7533,N_7864);
xnor U9771 (N_9771,N_7501,N_7888);
and U9772 (N_9772,N_8282,N_7721);
or U9773 (N_9773,N_8264,N_8514);
xnor U9774 (N_9774,N_8746,N_8486);
nor U9775 (N_9775,N_7722,N_8164);
and U9776 (N_9776,N_7822,N_8161);
and U9777 (N_9777,N_8742,N_7679);
and U9778 (N_9778,N_7650,N_8160);
or U9779 (N_9779,N_8026,N_8670);
nor U9780 (N_9780,N_7576,N_8164);
nor U9781 (N_9781,N_7610,N_8169);
nand U9782 (N_9782,N_7848,N_7869);
xnor U9783 (N_9783,N_8134,N_7665);
nand U9784 (N_9784,N_8660,N_8020);
nand U9785 (N_9785,N_8346,N_8459);
nor U9786 (N_9786,N_7577,N_8619);
nor U9787 (N_9787,N_8719,N_8081);
and U9788 (N_9788,N_7679,N_7545);
xnor U9789 (N_9789,N_7840,N_8162);
nor U9790 (N_9790,N_7711,N_8156);
or U9791 (N_9791,N_7508,N_7979);
or U9792 (N_9792,N_8632,N_8402);
nor U9793 (N_9793,N_8554,N_7905);
or U9794 (N_9794,N_8353,N_8038);
and U9795 (N_9795,N_7646,N_7583);
xnor U9796 (N_9796,N_7916,N_8719);
nand U9797 (N_9797,N_8291,N_8737);
nand U9798 (N_9798,N_8214,N_8514);
nand U9799 (N_9799,N_8634,N_8023);
or U9800 (N_9800,N_8013,N_8608);
and U9801 (N_9801,N_8172,N_8184);
and U9802 (N_9802,N_8394,N_8356);
xnor U9803 (N_9803,N_8086,N_8652);
xor U9804 (N_9804,N_8576,N_7824);
nor U9805 (N_9805,N_8133,N_7521);
and U9806 (N_9806,N_8672,N_8027);
or U9807 (N_9807,N_8355,N_7536);
or U9808 (N_9808,N_8527,N_8145);
xor U9809 (N_9809,N_8678,N_8743);
nand U9810 (N_9810,N_7886,N_8170);
nor U9811 (N_9811,N_7852,N_7627);
and U9812 (N_9812,N_7954,N_8496);
nand U9813 (N_9813,N_8363,N_7664);
and U9814 (N_9814,N_7962,N_7913);
xnor U9815 (N_9815,N_8492,N_8528);
nand U9816 (N_9816,N_7532,N_8639);
nand U9817 (N_9817,N_7714,N_7906);
or U9818 (N_9818,N_8252,N_8361);
xnor U9819 (N_9819,N_8568,N_8361);
nor U9820 (N_9820,N_7535,N_7524);
or U9821 (N_9821,N_8028,N_7539);
xor U9822 (N_9822,N_7982,N_8640);
or U9823 (N_9823,N_7548,N_7584);
or U9824 (N_9824,N_8708,N_8495);
and U9825 (N_9825,N_8217,N_7604);
nand U9826 (N_9826,N_8262,N_8222);
or U9827 (N_9827,N_7512,N_7633);
nor U9828 (N_9828,N_7824,N_7544);
or U9829 (N_9829,N_8745,N_7899);
and U9830 (N_9830,N_8580,N_8705);
and U9831 (N_9831,N_7558,N_7622);
or U9832 (N_9832,N_8264,N_8246);
nor U9833 (N_9833,N_8032,N_7744);
nor U9834 (N_9834,N_8659,N_8398);
and U9835 (N_9835,N_8005,N_7649);
nand U9836 (N_9836,N_7562,N_8371);
and U9837 (N_9837,N_7887,N_7706);
or U9838 (N_9838,N_7641,N_7957);
nand U9839 (N_9839,N_7929,N_8469);
nand U9840 (N_9840,N_8019,N_7521);
xor U9841 (N_9841,N_7890,N_8368);
and U9842 (N_9842,N_8212,N_8430);
or U9843 (N_9843,N_7799,N_7924);
nand U9844 (N_9844,N_7751,N_7979);
and U9845 (N_9845,N_8525,N_7922);
and U9846 (N_9846,N_7873,N_8743);
nor U9847 (N_9847,N_7759,N_8341);
nor U9848 (N_9848,N_7900,N_7552);
xor U9849 (N_9849,N_8184,N_7920);
and U9850 (N_9850,N_8427,N_8287);
nand U9851 (N_9851,N_8258,N_8201);
and U9852 (N_9852,N_7940,N_7511);
and U9853 (N_9853,N_8441,N_8095);
or U9854 (N_9854,N_7936,N_8626);
or U9855 (N_9855,N_8134,N_8360);
and U9856 (N_9856,N_7874,N_8260);
nand U9857 (N_9857,N_8669,N_8589);
nand U9858 (N_9858,N_8047,N_8449);
or U9859 (N_9859,N_8261,N_8096);
xnor U9860 (N_9860,N_7733,N_7877);
and U9861 (N_9861,N_7663,N_7774);
or U9862 (N_9862,N_8275,N_7939);
nor U9863 (N_9863,N_7771,N_7851);
and U9864 (N_9864,N_8670,N_7658);
xor U9865 (N_9865,N_8366,N_8290);
nand U9866 (N_9866,N_7554,N_8110);
xnor U9867 (N_9867,N_7714,N_8306);
nand U9868 (N_9868,N_7562,N_7669);
xor U9869 (N_9869,N_8277,N_8115);
nand U9870 (N_9870,N_8135,N_8362);
or U9871 (N_9871,N_7643,N_7669);
nor U9872 (N_9872,N_8123,N_7557);
nand U9873 (N_9873,N_7984,N_7743);
and U9874 (N_9874,N_7642,N_8715);
nand U9875 (N_9875,N_7672,N_7732);
and U9876 (N_9876,N_7550,N_7889);
nand U9877 (N_9877,N_7744,N_8333);
nand U9878 (N_9878,N_7999,N_7788);
nand U9879 (N_9879,N_8518,N_8650);
nand U9880 (N_9880,N_8287,N_7512);
nand U9881 (N_9881,N_7757,N_8371);
or U9882 (N_9882,N_8097,N_8517);
or U9883 (N_9883,N_8571,N_8150);
and U9884 (N_9884,N_8040,N_8287);
nor U9885 (N_9885,N_8285,N_8466);
xnor U9886 (N_9886,N_7926,N_8163);
or U9887 (N_9887,N_8716,N_8048);
and U9888 (N_9888,N_7627,N_8429);
and U9889 (N_9889,N_7501,N_7508);
and U9890 (N_9890,N_7838,N_7886);
nor U9891 (N_9891,N_7580,N_8428);
nand U9892 (N_9892,N_7757,N_8699);
nor U9893 (N_9893,N_8564,N_8716);
or U9894 (N_9894,N_8586,N_8448);
xnor U9895 (N_9895,N_8237,N_7897);
and U9896 (N_9896,N_8559,N_8053);
and U9897 (N_9897,N_8121,N_7637);
nor U9898 (N_9898,N_7987,N_7814);
xnor U9899 (N_9899,N_7817,N_7892);
xor U9900 (N_9900,N_7800,N_8561);
and U9901 (N_9901,N_8743,N_8441);
nand U9902 (N_9902,N_8200,N_8325);
or U9903 (N_9903,N_7709,N_8740);
nand U9904 (N_9904,N_8256,N_8706);
nor U9905 (N_9905,N_7703,N_8736);
or U9906 (N_9906,N_8686,N_8591);
or U9907 (N_9907,N_8328,N_8660);
nand U9908 (N_9908,N_7518,N_8312);
nor U9909 (N_9909,N_7811,N_7799);
xor U9910 (N_9910,N_7894,N_7737);
or U9911 (N_9911,N_8731,N_8536);
xor U9912 (N_9912,N_7830,N_7515);
nand U9913 (N_9913,N_8132,N_8149);
nor U9914 (N_9914,N_8328,N_7832);
and U9915 (N_9915,N_7805,N_8427);
nor U9916 (N_9916,N_8188,N_7882);
and U9917 (N_9917,N_7871,N_7952);
xor U9918 (N_9918,N_8175,N_8732);
nand U9919 (N_9919,N_7784,N_8201);
nand U9920 (N_9920,N_8011,N_8480);
and U9921 (N_9921,N_7971,N_8169);
or U9922 (N_9922,N_7797,N_8736);
nor U9923 (N_9923,N_7700,N_8323);
nor U9924 (N_9924,N_8454,N_8748);
xnor U9925 (N_9925,N_8139,N_7862);
xnor U9926 (N_9926,N_7512,N_7660);
or U9927 (N_9927,N_8317,N_8207);
nor U9928 (N_9928,N_7674,N_8713);
or U9929 (N_9929,N_8462,N_7857);
nor U9930 (N_9930,N_8668,N_7920);
xnor U9931 (N_9931,N_8679,N_8159);
or U9932 (N_9932,N_8212,N_8534);
and U9933 (N_9933,N_8297,N_7711);
nor U9934 (N_9934,N_8047,N_8342);
or U9935 (N_9935,N_7556,N_7926);
or U9936 (N_9936,N_8260,N_7893);
xnor U9937 (N_9937,N_8517,N_7633);
and U9938 (N_9938,N_8097,N_8303);
or U9939 (N_9939,N_7511,N_8742);
nor U9940 (N_9940,N_7670,N_8525);
and U9941 (N_9941,N_8281,N_7657);
xnor U9942 (N_9942,N_7965,N_8261);
and U9943 (N_9943,N_8639,N_7786);
nor U9944 (N_9944,N_8509,N_7844);
or U9945 (N_9945,N_8737,N_7713);
and U9946 (N_9946,N_7898,N_8275);
nor U9947 (N_9947,N_8258,N_7650);
nand U9948 (N_9948,N_8526,N_7673);
xnor U9949 (N_9949,N_7604,N_7834);
or U9950 (N_9950,N_8154,N_7878);
or U9951 (N_9951,N_8607,N_7581);
or U9952 (N_9952,N_7583,N_7769);
or U9953 (N_9953,N_8147,N_8444);
nor U9954 (N_9954,N_7956,N_8399);
or U9955 (N_9955,N_8130,N_7855);
or U9956 (N_9956,N_8171,N_8457);
and U9957 (N_9957,N_7534,N_8706);
or U9958 (N_9958,N_7570,N_8457);
or U9959 (N_9959,N_7928,N_8369);
and U9960 (N_9960,N_8640,N_8607);
xor U9961 (N_9961,N_8640,N_8723);
nor U9962 (N_9962,N_7648,N_8264);
nand U9963 (N_9963,N_7522,N_8535);
xnor U9964 (N_9964,N_8523,N_8696);
xnor U9965 (N_9965,N_8015,N_7906);
or U9966 (N_9966,N_7527,N_8539);
xor U9967 (N_9967,N_7657,N_7577);
and U9968 (N_9968,N_8359,N_8488);
nor U9969 (N_9969,N_8606,N_8072);
nor U9970 (N_9970,N_8035,N_7593);
xnor U9971 (N_9971,N_8539,N_8521);
and U9972 (N_9972,N_8145,N_8128);
or U9973 (N_9973,N_8052,N_7987);
nand U9974 (N_9974,N_7765,N_8301);
nor U9975 (N_9975,N_8692,N_7971);
xor U9976 (N_9976,N_7883,N_7879);
and U9977 (N_9977,N_7727,N_8117);
nand U9978 (N_9978,N_7974,N_7830);
and U9979 (N_9979,N_7974,N_8016);
and U9980 (N_9980,N_8165,N_7908);
and U9981 (N_9981,N_8626,N_8028);
or U9982 (N_9982,N_8354,N_8569);
nor U9983 (N_9983,N_7594,N_7554);
or U9984 (N_9984,N_7843,N_7984);
xor U9985 (N_9985,N_8360,N_7832);
and U9986 (N_9986,N_7825,N_7975);
nand U9987 (N_9987,N_8482,N_7650);
xor U9988 (N_9988,N_8271,N_8301);
xor U9989 (N_9989,N_8262,N_8018);
nor U9990 (N_9990,N_7541,N_8372);
xor U9991 (N_9991,N_8545,N_8511);
or U9992 (N_9992,N_8296,N_8123);
xor U9993 (N_9993,N_8015,N_8493);
or U9994 (N_9994,N_8194,N_8230);
nand U9995 (N_9995,N_7650,N_8113);
nand U9996 (N_9996,N_8654,N_7932);
nor U9997 (N_9997,N_7669,N_7647);
xor U9998 (N_9998,N_7574,N_8389);
xnor U9999 (N_9999,N_8259,N_8089);
xnor U10000 (N_10000,N_9619,N_9926);
nand U10001 (N_10001,N_9414,N_9431);
nand U10002 (N_10002,N_9039,N_9417);
nand U10003 (N_10003,N_9110,N_9690);
xnor U10004 (N_10004,N_8757,N_8952);
xnor U10005 (N_10005,N_9389,N_8922);
nand U10006 (N_10006,N_9382,N_9120);
and U10007 (N_10007,N_8800,N_9356);
nand U10008 (N_10008,N_9907,N_8762);
or U10009 (N_10009,N_9137,N_9374);
or U10010 (N_10010,N_9921,N_9524);
nand U10011 (N_10011,N_9986,N_8845);
nor U10012 (N_10012,N_8976,N_9892);
or U10013 (N_10013,N_9293,N_8989);
nand U10014 (N_10014,N_9254,N_8928);
and U10015 (N_10015,N_9673,N_9479);
xnor U10016 (N_10016,N_9401,N_9751);
or U10017 (N_10017,N_9993,N_9420);
nand U10018 (N_10018,N_9433,N_8823);
nor U10019 (N_10019,N_9896,N_9781);
nor U10020 (N_10020,N_9981,N_9552);
xor U10021 (N_10021,N_9027,N_9623);
xor U10022 (N_10022,N_9778,N_8916);
xnor U10023 (N_10023,N_9261,N_9017);
xnor U10024 (N_10024,N_9441,N_9483);
and U10025 (N_10025,N_8758,N_8780);
and U10026 (N_10026,N_9167,N_8893);
nor U10027 (N_10027,N_9286,N_8990);
xor U10028 (N_10028,N_9209,N_9422);
nand U10029 (N_10029,N_9753,N_9251);
xor U10030 (N_10030,N_9425,N_9544);
or U10031 (N_10031,N_8874,N_9192);
and U10032 (N_10032,N_8798,N_8931);
and U10033 (N_10033,N_9366,N_9657);
or U10034 (N_10034,N_9255,N_9691);
xor U10035 (N_10035,N_8847,N_9782);
xor U10036 (N_10036,N_9135,N_9074);
nor U10037 (N_10037,N_8796,N_9075);
xor U10038 (N_10038,N_9122,N_9170);
or U10039 (N_10039,N_9469,N_9296);
and U10040 (N_10040,N_9956,N_9330);
nor U10041 (N_10041,N_9735,N_8964);
nor U10042 (N_10042,N_9649,N_9791);
nor U10043 (N_10043,N_9920,N_9979);
nand U10044 (N_10044,N_9784,N_8871);
or U10045 (N_10045,N_9360,N_9612);
nor U10046 (N_10046,N_8837,N_9258);
or U10047 (N_10047,N_9653,N_9234);
and U10048 (N_10048,N_8977,N_9709);
and U10049 (N_10049,N_9622,N_9386);
nand U10050 (N_10050,N_9179,N_9598);
nand U10051 (N_10051,N_9243,N_9965);
nor U10052 (N_10052,N_9642,N_9221);
or U10053 (N_10053,N_9628,N_9652);
or U10054 (N_10054,N_8770,N_9011);
xnor U10055 (N_10055,N_9675,N_9134);
nor U10056 (N_10056,N_9766,N_8992);
nand U10057 (N_10057,N_9418,N_9439);
xor U10058 (N_10058,N_9563,N_9465);
nand U10059 (N_10059,N_9399,N_9725);
nand U10060 (N_10060,N_9335,N_9723);
nor U10061 (N_10061,N_9114,N_9082);
nand U10062 (N_10062,N_9253,N_9550);
nand U10063 (N_10063,N_9752,N_9555);
nand U10064 (N_10064,N_9842,N_9589);
and U10065 (N_10065,N_9952,N_9787);
xnor U10066 (N_10066,N_9034,N_9955);
nand U10067 (N_10067,N_9689,N_9950);
xor U10068 (N_10068,N_9924,N_8791);
or U10069 (N_10069,N_9284,N_9877);
or U10070 (N_10070,N_8973,N_8869);
xnor U10071 (N_10071,N_9174,N_9843);
nor U10072 (N_10072,N_9129,N_9520);
and U10073 (N_10073,N_9381,N_9162);
and U10074 (N_10074,N_9868,N_9083);
and U10075 (N_10075,N_9009,N_8759);
xor U10076 (N_10076,N_9757,N_8946);
nand U10077 (N_10077,N_9999,N_9805);
or U10078 (N_10078,N_9239,N_9367);
nor U10079 (N_10079,N_9428,N_8831);
or U10080 (N_10080,N_9499,N_8863);
xnor U10081 (N_10081,N_8889,N_9313);
nand U10082 (N_10082,N_9069,N_9117);
or U10083 (N_10083,N_9738,N_9963);
nand U10084 (N_10084,N_8828,N_9040);
or U10085 (N_10085,N_9046,N_9685);
and U10086 (N_10086,N_9756,N_9067);
and U10087 (N_10087,N_9404,N_9001);
xnor U10088 (N_10088,N_9664,N_9206);
nand U10089 (N_10089,N_8934,N_9827);
and U10090 (N_10090,N_9291,N_9373);
or U10091 (N_10091,N_9486,N_9852);
and U10092 (N_10092,N_9530,N_9475);
and U10093 (N_10093,N_9809,N_8811);
or U10094 (N_10094,N_8767,N_8755);
nand U10095 (N_10095,N_9858,N_9720);
or U10096 (N_10096,N_9108,N_9525);
and U10097 (N_10097,N_8962,N_9910);
and U10098 (N_10098,N_9825,N_8890);
and U10099 (N_10099,N_8904,N_9887);
nor U10100 (N_10100,N_9071,N_9925);
and U10101 (N_10101,N_9509,N_9247);
and U10102 (N_10102,N_8777,N_9201);
xor U10103 (N_10103,N_9904,N_9161);
or U10104 (N_10104,N_9383,N_9281);
nor U10105 (N_10105,N_9180,N_8887);
nand U10106 (N_10106,N_9014,N_9567);
or U10107 (N_10107,N_9307,N_9398);
or U10108 (N_10108,N_9283,N_9746);
nand U10109 (N_10109,N_9764,N_9372);
xnor U10110 (N_10110,N_9610,N_9343);
nand U10111 (N_10111,N_9015,N_9856);
or U10112 (N_10112,N_9616,N_9380);
nor U10113 (N_10113,N_8986,N_9779);
xnor U10114 (N_10114,N_9311,N_8998);
nand U10115 (N_10115,N_9005,N_9976);
or U10116 (N_10116,N_8877,N_9661);
and U10117 (N_10117,N_9866,N_9724);
nand U10118 (N_10118,N_9731,N_9080);
xor U10119 (N_10119,N_9964,N_8921);
and U10120 (N_10120,N_9237,N_9629);
xnor U10121 (N_10121,N_9996,N_9324);
xnor U10122 (N_10122,N_8833,N_9066);
nor U10123 (N_10123,N_9312,N_9156);
or U10124 (N_10124,N_9448,N_9309);
or U10125 (N_10125,N_9427,N_9743);
or U10126 (N_10126,N_9565,N_9620);
nand U10127 (N_10127,N_9785,N_9705);
or U10128 (N_10128,N_9190,N_9645);
nand U10129 (N_10129,N_8805,N_9157);
nand U10130 (N_10130,N_9534,N_8751);
or U10131 (N_10131,N_9477,N_9814);
and U10132 (N_10132,N_9348,N_9480);
or U10133 (N_10133,N_9061,N_8878);
xnor U10134 (N_10134,N_9365,N_9242);
nor U10135 (N_10135,N_9760,N_9495);
nor U10136 (N_10136,N_9513,N_8803);
xnor U10137 (N_10137,N_9194,N_9940);
nand U10138 (N_10138,N_9775,N_9604);
xnor U10139 (N_10139,N_9349,N_9767);
and U10140 (N_10140,N_8752,N_8854);
xor U10141 (N_10141,N_9630,N_9278);
nand U10142 (N_10142,N_9638,N_9023);
xor U10143 (N_10143,N_8974,N_8801);
or U10144 (N_10144,N_9870,N_9862);
xnor U10145 (N_10145,N_9079,N_9191);
and U10146 (N_10146,N_9199,N_9801);
nor U10147 (N_10147,N_9452,N_9517);
or U10148 (N_10148,N_9058,N_8781);
nor U10149 (N_10149,N_8985,N_8929);
nor U10150 (N_10150,N_9806,N_9531);
nor U10151 (N_10151,N_9086,N_9337);
nand U10152 (N_10152,N_9203,N_9466);
nand U10153 (N_10153,N_9406,N_9248);
nand U10154 (N_10154,N_8900,N_9139);
xor U10155 (N_10155,N_9244,N_9101);
xor U10156 (N_10156,N_9213,N_9793);
and U10157 (N_10157,N_9733,N_8840);
nor U10158 (N_10158,N_8813,N_9118);
nor U10159 (N_10159,N_9734,N_9432);
or U10160 (N_10160,N_9811,N_9917);
nand U10161 (N_10161,N_8794,N_9500);
or U10162 (N_10162,N_8814,N_9387);
nor U10163 (N_10163,N_9193,N_9091);
or U10164 (N_10164,N_9602,N_9217);
xnor U10165 (N_10165,N_8923,N_9676);
or U10166 (N_10166,N_9823,N_9100);
nor U10167 (N_10167,N_9197,N_9336);
xor U10168 (N_10168,N_9172,N_9489);
nand U10169 (N_10169,N_9304,N_9019);
nand U10170 (N_10170,N_9717,N_9831);
and U10171 (N_10171,N_8872,N_9429);
xnor U10172 (N_10172,N_9329,N_9613);
xor U10173 (N_10173,N_9561,N_9305);
xor U10174 (N_10174,N_9674,N_9759);
nor U10175 (N_10175,N_9872,N_9942);
or U10176 (N_10176,N_9798,N_9588);
and U10177 (N_10177,N_9245,N_9178);
and U10178 (N_10178,N_9656,N_8843);
nand U10179 (N_10179,N_9430,N_9570);
nor U10180 (N_10180,N_9096,N_8761);
xor U10181 (N_10181,N_9270,N_9906);
nand U10182 (N_10182,N_8786,N_9755);
and U10183 (N_10183,N_9155,N_9516);
xnor U10184 (N_10184,N_9817,N_9455);
xnor U10185 (N_10185,N_9147,N_9140);
nor U10186 (N_10186,N_8903,N_8797);
or U10187 (N_10187,N_9990,N_9663);
nor U10188 (N_10188,N_8884,N_9624);
or U10189 (N_10189,N_9944,N_9458);
and U10190 (N_10190,N_9092,N_9052);
and U10191 (N_10191,N_9405,N_9937);
nor U10192 (N_10192,N_9468,N_9218);
nand U10193 (N_10193,N_8880,N_9508);
nand U10194 (N_10194,N_9773,N_9594);
xor U10195 (N_10195,N_9539,N_9216);
xnor U10196 (N_10196,N_9712,N_9169);
or U10197 (N_10197,N_9163,N_8776);
xor U10198 (N_10198,N_8933,N_9476);
nand U10199 (N_10199,N_9851,N_9205);
nor U10200 (N_10200,N_8954,N_9158);
or U10201 (N_10201,N_9472,N_9953);
nand U10202 (N_10202,N_8766,N_9984);
nor U10203 (N_10203,N_8816,N_9655);
xor U10204 (N_10204,N_9395,N_9089);
or U10205 (N_10205,N_9423,N_9850);
nand U10206 (N_10206,N_9750,N_9224);
and U10207 (N_10207,N_9130,N_9124);
xnor U10208 (N_10208,N_9013,N_8821);
or U10209 (N_10209,N_8888,N_9277);
and U10210 (N_10210,N_9536,N_9359);
or U10211 (N_10211,N_9049,N_9447);
and U10212 (N_10212,N_9727,N_8939);
xor U10213 (N_10213,N_9350,N_9532);
or U10214 (N_10214,N_8760,N_9765);
or U10215 (N_10215,N_9370,N_9772);
and U10216 (N_10216,N_9646,N_9300);
nand U10217 (N_10217,N_8875,N_9543);
or U10218 (N_10218,N_9057,N_9686);
and U10219 (N_10219,N_9949,N_9869);
xnor U10220 (N_10220,N_8827,N_9780);
and U10221 (N_10221,N_9927,N_8835);
nand U10222 (N_10222,N_9113,N_9802);
or U10223 (N_10223,N_8945,N_8789);
or U10224 (N_10224,N_9796,N_9880);
and U10225 (N_10225,N_8784,N_9145);
and U10226 (N_10226,N_9094,N_9679);
nor U10227 (N_10227,N_9960,N_9871);
xnor U10228 (N_10228,N_9107,N_9585);
xor U10229 (N_10229,N_8993,N_9708);
nor U10230 (N_10230,N_9215,N_9435);
xor U10231 (N_10231,N_9368,N_9351);
nor U10232 (N_10232,N_8836,N_9220);
or U10233 (N_10233,N_9085,N_8915);
xnor U10234 (N_10234,N_8948,N_9650);
nor U10235 (N_10235,N_9473,N_9461);
nor U10236 (N_10236,N_9935,N_9551);
and U10237 (N_10237,N_9715,N_9160);
xor U10238 (N_10238,N_8925,N_9995);
or U10239 (N_10239,N_9403,N_8969);
xor U10240 (N_10240,N_9148,N_8818);
nand U10241 (N_10241,N_9202,N_9975);
nand U10242 (N_10242,N_9143,N_8865);
nand U10243 (N_10243,N_8942,N_8792);
or U10244 (N_10244,N_9671,N_9697);
or U10245 (N_10245,N_9314,N_9214);
nor U10246 (N_10246,N_9666,N_9542);
nand U10247 (N_10247,N_9838,N_9064);
or U10248 (N_10248,N_8941,N_9200);
and U10249 (N_10249,N_9334,N_9518);
nor U10250 (N_10250,N_9068,N_9834);
nor U10251 (N_10251,N_8795,N_8765);
or U10252 (N_10252,N_9886,N_9595);
nor U10253 (N_10253,N_8987,N_9047);
nand U10254 (N_10254,N_9928,N_9030);
nand U10255 (N_10255,N_9498,N_8943);
nor U10256 (N_10256,N_9867,N_8785);
nand U10257 (N_10257,N_8978,N_9164);
xor U10258 (N_10258,N_9295,N_8913);
xor U10259 (N_10259,N_8851,N_9770);
xor U10260 (N_10260,N_8950,N_9044);
xnor U10261 (N_10261,N_9865,N_9945);
nor U10262 (N_10262,N_9006,N_8901);
and U10263 (N_10263,N_9813,N_9012);
and U10264 (N_10264,N_9932,N_8824);
xnor U10265 (N_10265,N_9884,N_8826);
and U10266 (N_10266,N_9402,N_9881);
or U10267 (N_10267,N_9133,N_9824);
nor U10268 (N_10268,N_9810,N_9885);
nand U10269 (N_10269,N_8850,N_9592);
and U10270 (N_10270,N_9978,N_8858);
or U10271 (N_10271,N_9672,N_9583);
or U10272 (N_10272,N_9166,N_9821);
nor U10273 (N_10273,N_9832,N_9273);
nor U10274 (N_10274,N_8860,N_8932);
or U10275 (N_10275,N_9855,N_9128);
or U10276 (N_10276,N_9181,N_9090);
xor U10277 (N_10277,N_9299,N_9041);
nor U10278 (N_10278,N_9297,N_9424);
or U10279 (N_10279,N_9703,N_9228);
nor U10280 (N_10280,N_9152,N_9288);
xnor U10281 (N_10281,N_9694,N_9116);
and U10282 (N_10282,N_9988,N_8963);
or U10283 (N_10283,N_8778,N_9186);
or U10284 (N_10284,N_9319,N_9632);
and U10285 (N_10285,N_9864,N_9104);
nor U10286 (N_10286,N_9358,N_9246);
and U10287 (N_10287,N_9882,N_9891);
nor U10288 (N_10288,N_8807,N_9822);
xor U10289 (N_10289,N_8808,N_8855);
xnor U10290 (N_10290,N_9636,N_9758);
and U10291 (N_10291,N_9210,N_9501);
nand U10292 (N_10292,N_9700,N_9835);
nand U10293 (N_10293,N_9545,N_8873);
nand U10294 (N_10294,N_9303,N_9883);
and U10295 (N_10295,N_9577,N_8830);
or U10296 (N_10296,N_9590,N_9032);
xor U10297 (N_10297,N_9361,N_9994);
and U10298 (N_10298,N_9035,N_9861);
xnor U10299 (N_10299,N_8936,N_9002);
and U10300 (N_10300,N_8917,N_9553);
and U10301 (N_10301,N_9631,N_9911);
and U10302 (N_10302,N_9457,N_8809);
or U10303 (N_10303,N_9150,N_8820);
or U10304 (N_10304,N_9141,N_9878);
xor U10305 (N_10305,N_9637,N_9189);
and U10306 (N_10306,N_9493,N_9446);
or U10307 (N_10307,N_9322,N_9692);
or U10308 (N_10308,N_9571,N_9310);
or U10309 (N_10309,N_9898,N_9774);
and U10310 (N_10310,N_9776,N_9989);
nor U10311 (N_10311,N_9815,N_9879);
xor U10312 (N_10312,N_9260,N_9105);
xor U10313 (N_10313,N_9236,N_9177);
and U10314 (N_10314,N_8883,N_8935);
nor U10315 (N_10315,N_9505,N_9050);
nand U10316 (N_10316,N_8907,N_9957);
nor U10317 (N_10317,N_9808,N_9275);
and U10318 (N_10318,N_9506,N_9626);
or U10319 (N_10319,N_8815,N_9647);
xor U10320 (N_10320,N_9397,N_8898);
nor U10321 (N_10321,N_9923,N_8790);
and U10322 (N_10322,N_9434,N_9095);
xnor U10323 (N_10323,N_9639,N_9786);
nor U10324 (N_10324,N_9959,N_9151);
xnor U10325 (N_10325,N_9062,N_8853);
nor U10326 (N_10326,N_9377,N_9238);
and U10327 (N_10327,N_8832,N_9393);
nor U10328 (N_10328,N_9276,N_9392);
nor U10329 (N_10329,N_9769,N_8799);
and U10330 (N_10330,N_9048,N_9818);
xor U10331 (N_10331,N_9596,N_9568);
nor U10332 (N_10332,N_9026,N_9833);
nor U10333 (N_10333,N_9175,N_9326);
nand U10334 (N_10334,N_9948,N_9909);
and U10335 (N_10335,N_9608,N_8838);
nand U10336 (N_10336,N_8846,N_9693);
or U10337 (N_10337,N_9354,N_9056);
nand U10338 (N_10338,N_9346,N_9510);
or U10339 (N_10339,N_9249,N_9931);
and U10340 (N_10340,N_9918,N_9038);
nand U10341 (N_10341,N_8981,N_9970);
and U10342 (N_10342,N_9803,N_9732);
nand U10343 (N_10343,N_8841,N_9573);
xor U10344 (N_10344,N_8774,N_9938);
or U10345 (N_10345,N_9826,N_9274);
and U10346 (N_10346,N_9761,N_9841);
and U10347 (N_10347,N_9481,N_9371);
nor U10348 (N_10348,N_9073,N_9819);
or U10349 (N_10349,N_9388,N_8886);
and U10350 (N_10350,N_9951,N_9173);
nor U10351 (N_10351,N_9125,N_9138);
nand U10352 (N_10352,N_9688,N_8756);
nor U10353 (N_10353,N_9364,N_9271);
or U10354 (N_10354,N_8919,N_9208);
or U10355 (N_10355,N_9268,N_8970);
and U10356 (N_10356,N_9450,N_9933);
or U10357 (N_10357,N_9741,N_9974);
nor U10358 (N_10358,N_9264,N_9967);
or U10359 (N_10359,N_9947,N_9055);
or U10360 (N_10360,N_9492,N_9744);
xor U10361 (N_10361,N_9605,N_9033);
and U10362 (N_10362,N_9323,N_9837);
xor U10363 (N_10363,N_9470,N_8879);
and U10364 (N_10364,N_8772,N_9106);
or U10365 (N_10365,N_9207,N_8908);
and U10366 (N_10366,N_9449,N_9936);
or U10367 (N_10367,N_9941,N_8955);
or U10368 (N_10368,N_9719,N_9985);
or U10369 (N_10369,N_9681,N_8839);
and U10370 (N_10370,N_9292,N_9165);
xnor U10371 (N_10371,N_9451,N_9426);
or U10372 (N_10372,N_9250,N_9899);
and U10373 (N_10373,N_9227,N_9987);
or U10374 (N_10374,N_9266,N_9729);
nor U10375 (N_10375,N_9912,N_8842);
and U10376 (N_10376,N_9257,N_8979);
xnor U10377 (N_10377,N_9716,N_9853);
xor U10378 (N_10378,N_8856,N_9737);
and U10379 (N_10379,N_8859,N_9894);
and U10380 (N_10380,N_9929,N_9098);
and U10381 (N_10381,N_9718,N_9614);
xnor U10382 (N_10382,N_9900,N_9340);
or U10383 (N_10383,N_9229,N_9070);
xnor U10384 (N_10384,N_9528,N_9554);
xnor U10385 (N_10385,N_8997,N_9347);
nand U10386 (N_10386,N_9408,N_9302);
nor U10387 (N_10387,N_9280,N_9231);
nand U10388 (N_10388,N_9799,N_9682);
nor U10389 (N_10389,N_9627,N_8849);
nand U10390 (N_10390,N_9327,N_9232);
nand U10391 (N_10391,N_9204,N_9582);
nor U10392 (N_10392,N_9540,N_9512);
and U10393 (N_10393,N_9460,N_8937);
nand U10394 (N_10394,N_9437,N_9575);
nand U10395 (N_10395,N_9574,N_9847);
nor U10396 (N_10396,N_9601,N_9053);
xor U10397 (N_10397,N_9749,N_9306);
or U10398 (N_10398,N_8894,N_9004);
or U10399 (N_10399,N_9893,N_9962);
and U10400 (N_10400,N_8947,N_9076);
nor U10401 (N_10401,N_8967,N_8817);
nand U10402 (N_10402,N_8961,N_9634);
xnor U10403 (N_10403,N_9790,N_8899);
nor U10404 (N_10404,N_9262,N_9196);
and U10405 (N_10405,N_8980,N_9454);
xor U10406 (N_10406,N_9059,N_8864);
and U10407 (N_10407,N_9580,N_9287);
and U10408 (N_10408,N_9007,N_9581);
or U10409 (N_10409,N_9659,N_9897);
nand U10410 (N_10410,N_8882,N_9338);
nand U10411 (N_10411,N_9603,N_8787);
xnor U10412 (N_10412,N_8910,N_9812);
xor U10413 (N_10413,N_9903,N_9093);
xor U10414 (N_10414,N_9919,N_8892);
nand U10415 (N_10415,N_9529,N_8870);
nor U10416 (N_10416,N_9037,N_9294);
nor U10417 (N_10417,N_8881,N_9320);
nor U10418 (N_10418,N_9593,N_8912);
xnor U10419 (N_10419,N_9102,N_9579);
and U10420 (N_10420,N_9667,N_9747);
xor U10421 (N_10421,N_9054,N_9440);
nor U10422 (N_10422,N_9353,N_8991);
nor U10423 (N_10423,N_8906,N_8806);
xnor U10424 (N_10424,N_9618,N_9487);
and U10425 (N_10425,N_9783,N_9504);
or U10426 (N_10426,N_9088,N_8927);
and U10427 (N_10427,N_8788,N_9018);
nand U10428 (N_10428,N_9968,N_9860);
nor U10429 (N_10429,N_9131,N_9142);
xor U10430 (N_10430,N_9485,N_9547);
and U10431 (N_10431,N_9282,N_9185);
and U10432 (N_10432,N_8867,N_9713);
nor U10433 (N_10433,N_9409,N_8971);
or U10434 (N_10434,N_9654,N_9526);
nand U10435 (N_10435,N_9848,N_9474);
nor U10436 (N_10436,N_9111,N_9939);
nand U10437 (N_10437,N_9467,N_9849);
and U10438 (N_10438,N_9836,N_9235);
or U10439 (N_10439,N_9711,N_9168);
xnor U10440 (N_10440,N_9154,N_8822);
nand U10441 (N_10441,N_9464,N_9328);
or U10442 (N_10442,N_9020,N_9438);
nand U10443 (N_10443,N_9225,N_8966);
and U10444 (N_10444,N_9127,N_9357);
nand U10445 (N_10445,N_9680,N_8750);
nand U10446 (N_10446,N_8779,N_9376);
xnor U10447 (N_10447,N_9665,N_9797);
xnor U10448 (N_10448,N_9740,N_9222);
nor U10449 (N_10449,N_9490,N_9562);
nand U10450 (N_10450,N_9889,N_9149);
or U10451 (N_10451,N_9109,N_9739);
or U10452 (N_10452,N_8895,N_9043);
or U10453 (N_10453,N_9036,N_9198);
nor U10454 (N_10454,N_9569,N_9820);
xnor U10455 (N_10455,N_9507,N_9146);
or U10456 (N_10456,N_8930,N_9607);
xnor U10457 (N_10457,N_9123,N_9519);
nor U10458 (N_10458,N_9503,N_9648);
nand U10459 (N_10459,N_9259,N_8940);
xor U10460 (N_10460,N_9187,N_9321);
and U10461 (N_10461,N_9223,N_8911);
nor U10462 (N_10462,N_9859,N_9410);
or U10463 (N_10463,N_9285,N_9317);
and U10464 (N_10464,N_9643,N_9704);
nand U10465 (N_10465,N_9863,N_9669);
and U10466 (N_10466,N_9115,N_9339);
or U10467 (N_10467,N_8983,N_9839);
or U10468 (N_10468,N_9754,N_9789);
nand U10469 (N_10469,N_9816,N_9211);
nand U10470 (N_10470,N_9546,N_9771);
or U10471 (N_10471,N_8891,N_9230);
or U10472 (N_10472,N_9854,N_9060);
nor U10473 (N_10473,N_9980,N_9998);
nor U10474 (N_10474,N_9901,N_9184);
nor U10475 (N_10475,N_8896,N_9584);
xnor U10476 (N_10476,N_9930,N_9972);
xnor U10477 (N_10477,N_8852,N_9385);
or U10478 (N_10478,N_9934,N_9651);
nor U10479 (N_10479,N_9644,N_8769);
and U10480 (N_10480,N_9606,N_9830);
and U10481 (N_10481,N_8968,N_9394);
nand U10482 (N_10482,N_9463,N_9000);
or U10483 (N_10483,N_9991,N_9523);
nor U10484 (N_10484,N_9308,N_9706);
or U10485 (N_10485,N_8810,N_9600);
nor U10486 (N_10486,N_9252,N_9698);
xor U10487 (N_10487,N_9973,N_9511);
or U10488 (N_10488,N_8897,N_9456);
xor U10489 (N_10489,N_9908,N_9522);
nor U10490 (N_10490,N_9369,N_9971);
nand U10491 (N_10491,N_8982,N_9436);
xor U10492 (N_10492,N_9097,N_9029);
nor U10493 (N_10493,N_9421,N_9289);
nor U10494 (N_10494,N_8988,N_9412);
xnor U10495 (N_10495,N_9621,N_9265);
xor U10496 (N_10496,N_9514,N_9954);
nor U10497 (N_10497,N_9298,N_9625);
nand U10498 (N_10498,N_9640,N_8972);
nor U10499 (N_10499,N_9462,N_9591);
nor U10500 (N_10500,N_9515,N_9792);
xnor U10501 (N_10501,N_9958,N_9742);
nor U10502 (N_10502,N_9419,N_9662);
nor U10503 (N_10503,N_9888,N_9379);
or U10504 (N_10504,N_9290,N_8975);
or U10505 (N_10505,N_9396,N_8764);
xor U10506 (N_10506,N_9445,N_8868);
nor U10507 (N_10507,N_9969,N_9442);
nand U10508 (N_10508,N_9484,N_9804);
nor U10509 (N_10509,N_9391,N_9586);
nor U10510 (N_10510,N_9844,N_9548);
nor U10511 (N_10511,N_9176,N_9763);
nor U10512 (N_10512,N_9895,N_9025);
or U10513 (N_10513,N_8958,N_9016);
nor U10514 (N_10514,N_9087,N_9267);
nand U10515 (N_10515,N_9794,N_9699);
xnor U10516 (N_10516,N_8804,N_9660);
nand U10517 (N_10517,N_9045,N_8829);
and U10518 (N_10518,N_9576,N_9363);
or U10519 (N_10519,N_8848,N_9182);
and U10520 (N_10520,N_9777,N_8876);
xor U10521 (N_10521,N_9943,N_8938);
xor U10522 (N_10522,N_8812,N_9233);
and U10523 (N_10523,N_9762,N_9828);
nand U10524 (N_10524,N_9678,N_9722);
or U10525 (N_10525,N_8793,N_9617);
nand U10526 (N_10526,N_9344,N_8959);
nor U10527 (N_10527,N_8802,N_9263);
nand U10528 (N_10528,N_9683,N_9042);
or U10529 (N_10529,N_8834,N_9913);
and U10530 (N_10530,N_8951,N_9378);
or U10531 (N_10531,N_9800,N_9549);
nand U10532 (N_10532,N_9065,N_9922);
xnor U10533 (N_10533,N_9535,N_9564);
nor U10534 (N_10534,N_9875,N_9482);
xnor U10535 (N_10535,N_9099,N_9031);
nand U10536 (N_10536,N_9873,N_9977);
or U10537 (N_10537,N_9611,N_9840);
nor U10538 (N_10538,N_9084,N_9521);
nand U10539 (N_10539,N_9916,N_9641);
nand U10540 (N_10540,N_9992,N_9241);
nor U10541 (N_10541,N_9212,N_9721);
or U10542 (N_10542,N_9256,N_8953);
xor U10543 (N_10543,N_9345,N_9415);
nand U10544 (N_10544,N_9453,N_9876);
or U10545 (N_10545,N_8965,N_9730);
and U10546 (N_10546,N_8957,N_8999);
xnor U10547 (N_10547,N_9444,N_9795);
and U10548 (N_10548,N_9341,N_8924);
xor U10549 (N_10549,N_9494,N_9443);
or U10550 (N_10550,N_9566,N_9538);
nand U10551 (N_10551,N_9416,N_8861);
and U10552 (N_10552,N_9707,N_8956);
and U10553 (N_10553,N_9407,N_9541);
nand U10554 (N_10554,N_8984,N_9728);
and U10555 (N_10555,N_9587,N_8902);
xnor U10556 (N_10556,N_9171,N_8775);
nand U10557 (N_10557,N_8783,N_8949);
or U10558 (N_10558,N_9471,N_8753);
xor U10559 (N_10559,N_9668,N_9072);
nand U10560 (N_10560,N_9658,N_9609);
nor U10561 (N_10561,N_9279,N_8994);
nor U10562 (N_10562,N_8768,N_9745);
and U10563 (N_10563,N_9983,N_8819);
or U10564 (N_10564,N_9269,N_9961);
nand U10565 (N_10565,N_9112,N_9226);
nand U10566 (N_10566,N_9997,N_9845);
or U10567 (N_10567,N_9597,N_9829);
and U10568 (N_10568,N_9874,N_9558);
or U10569 (N_10569,N_9533,N_9670);
and U10570 (N_10570,N_9272,N_9021);
nand U10571 (N_10571,N_9768,N_8914);
xnor U10572 (N_10572,N_9890,N_9077);
or U10573 (N_10573,N_8754,N_9615);
xor U10574 (N_10574,N_9696,N_8825);
nand U10575 (N_10575,N_9063,N_9022);
xor U10576 (N_10576,N_9556,N_9684);
and U10577 (N_10577,N_9497,N_9677);
xor U10578 (N_10578,N_9578,N_9736);
or U10579 (N_10579,N_9219,N_9126);
or U10580 (N_10580,N_9301,N_9788);
or U10581 (N_10581,N_9807,N_9390);
and U10582 (N_10582,N_9478,N_9008);
or U10583 (N_10583,N_9411,N_9315);
or U10584 (N_10584,N_9183,N_9701);
xor U10585 (N_10585,N_8909,N_9496);
nor U10586 (N_10586,N_9857,N_9316);
nand U10587 (N_10587,N_9132,N_9560);
or U10588 (N_10588,N_9144,N_8857);
xor U10589 (N_10589,N_9332,N_9342);
and U10590 (N_10590,N_9413,N_8771);
or U10591 (N_10591,N_9384,N_9153);
xnor U10592 (N_10592,N_8926,N_8844);
xnor U10593 (N_10593,N_9051,N_9240);
xor U10594 (N_10594,N_8866,N_8944);
nand U10595 (N_10595,N_9748,N_9946);
or U10596 (N_10596,N_9188,N_9081);
or U10597 (N_10597,N_9362,N_9599);
nand U10598 (N_10598,N_9375,N_9331);
or U10599 (N_10599,N_9710,N_9010);
or U10600 (N_10600,N_8918,N_9352);
nand U10601 (N_10601,N_8862,N_9121);
nand U10602 (N_10602,N_9537,N_8782);
nor U10603 (N_10603,N_9502,N_9966);
nor U10604 (N_10604,N_9915,N_8996);
or U10605 (N_10605,N_9702,N_9982);
nand U10606 (N_10606,N_9559,N_9028);
nor U10607 (N_10607,N_9024,N_9695);
nand U10608 (N_10608,N_8773,N_9635);
nand U10609 (N_10609,N_9003,N_9527);
and U10610 (N_10610,N_9318,N_9355);
nand U10611 (N_10611,N_9687,N_8960);
and U10612 (N_10612,N_9195,N_8885);
nand U10613 (N_10613,N_9136,N_9557);
xor U10614 (N_10614,N_9103,N_9078);
and U10615 (N_10615,N_9633,N_9491);
xnor U10616 (N_10616,N_9846,N_9914);
xor U10617 (N_10617,N_9902,N_9400);
nand U10618 (N_10618,N_9905,N_9325);
or U10619 (N_10619,N_9459,N_9119);
and U10620 (N_10620,N_9159,N_9333);
and U10621 (N_10621,N_8905,N_9488);
nor U10622 (N_10622,N_9726,N_8763);
and U10623 (N_10623,N_8920,N_8995);
or U10624 (N_10624,N_9714,N_9572);
or U10625 (N_10625,N_9930,N_9209);
nor U10626 (N_10626,N_9461,N_9701);
xnor U10627 (N_10627,N_8982,N_9897);
nand U10628 (N_10628,N_9204,N_9285);
nor U10629 (N_10629,N_9383,N_9907);
nor U10630 (N_10630,N_9722,N_9217);
xnor U10631 (N_10631,N_9714,N_9371);
nand U10632 (N_10632,N_9252,N_9190);
nor U10633 (N_10633,N_9433,N_8917);
nor U10634 (N_10634,N_9330,N_9420);
nor U10635 (N_10635,N_9634,N_9136);
xnor U10636 (N_10636,N_8781,N_9388);
or U10637 (N_10637,N_9731,N_8988);
nand U10638 (N_10638,N_8804,N_9806);
nor U10639 (N_10639,N_9119,N_8997);
nor U10640 (N_10640,N_9397,N_9413);
xnor U10641 (N_10641,N_9044,N_9830);
or U10642 (N_10642,N_9366,N_9847);
nor U10643 (N_10643,N_9508,N_8828);
xnor U10644 (N_10644,N_9601,N_9883);
or U10645 (N_10645,N_9585,N_8855);
xnor U10646 (N_10646,N_9850,N_9210);
and U10647 (N_10647,N_9954,N_9910);
nand U10648 (N_10648,N_9879,N_9663);
and U10649 (N_10649,N_9405,N_9607);
xor U10650 (N_10650,N_8985,N_9133);
or U10651 (N_10651,N_9683,N_9465);
xor U10652 (N_10652,N_9491,N_9841);
or U10653 (N_10653,N_9538,N_8986);
nor U10654 (N_10654,N_9130,N_9625);
and U10655 (N_10655,N_8861,N_9049);
and U10656 (N_10656,N_9849,N_9249);
nand U10657 (N_10657,N_9063,N_9451);
nand U10658 (N_10658,N_8980,N_9676);
or U10659 (N_10659,N_9544,N_9495);
nand U10660 (N_10660,N_9767,N_8873);
nor U10661 (N_10661,N_9614,N_9713);
nand U10662 (N_10662,N_9808,N_9370);
or U10663 (N_10663,N_8794,N_9754);
and U10664 (N_10664,N_9992,N_9670);
xor U10665 (N_10665,N_9463,N_9422);
and U10666 (N_10666,N_9604,N_8809);
or U10667 (N_10667,N_9360,N_9862);
nand U10668 (N_10668,N_9815,N_9748);
xor U10669 (N_10669,N_9608,N_9652);
nand U10670 (N_10670,N_9876,N_8975);
nand U10671 (N_10671,N_8898,N_9755);
nor U10672 (N_10672,N_9002,N_9469);
nor U10673 (N_10673,N_9439,N_9909);
and U10674 (N_10674,N_9584,N_9321);
xnor U10675 (N_10675,N_9077,N_9893);
nand U10676 (N_10676,N_9704,N_9171);
and U10677 (N_10677,N_9626,N_9641);
and U10678 (N_10678,N_9657,N_9735);
nand U10679 (N_10679,N_9574,N_8894);
nor U10680 (N_10680,N_9451,N_9695);
nand U10681 (N_10681,N_8951,N_9478);
nor U10682 (N_10682,N_8867,N_9514);
or U10683 (N_10683,N_9849,N_8928);
and U10684 (N_10684,N_9667,N_8895);
and U10685 (N_10685,N_9152,N_9137);
nand U10686 (N_10686,N_9858,N_9548);
nor U10687 (N_10687,N_9346,N_8842);
nand U10688 (N_10688,N_9386,N_9389);
xnor U10689 (N_10689,N_9351,N_9027);
nand U10690 (N_10690,N_9047,N_9257);
xnor U10691 (N_10691,N_9899,N_9879);
nand U10692 (N_10692,N_9708,N_9055);
nand U10693 (N_10693,N_8873,N_9525);
nand U10694 (N_10694,N_9009,N_9648);
nor U10695 (N_10695,N_9932,N_9380);
and U10696 (N_10696,N_9347,N_9083);
xnor U10697 (N_10697,N_9899,N_8882);
or U10698 (N_10698,N_9783,N_9122);
or U10699 (N_10699,N_9980,N_8821);
xor U10700 (N_10700,N_8983,N_9687);
xor U10701 (N_10701,N_8769,N_9760);
and U10702 (N_10702,N_9573,N_8969);
and U10703 (N_10703,N_9569,N_9544);
or U10704 (N_10704,N_9681,N_9414);
nand U10705 (N_10705,N_9868,N_8900);
xor U10706 (N_10706,N_8766,N_8992);
nand U10707 (N_10707,N_9243,N_8773);
nor U10708 (N_10708,N_9325,N_9964);
or U10709 (N_10709,N_9405,N_9344);
nor U10710 (N_10710,N_9928,N_8912);
xnor U10711 (N_10711,N_9136,N_9834);
and U10712 (N_10712,N_9309,N_9206);
xor U10713 (N_10713,N_9146,N_9283);
xor U10714 (N_10714,N_9985,N_8818);
xor U10715 (N_10715,N_9307,N_9913);
and U10716 (N_10716,N_9516,N_9482);
nor U10717 (N_10717,N_9956,N_8951);
xnor U10718 (N_10718,N_9315,N_9776);
nand U10719 (N_10719,N_8792,N_8777);
or U10720 (N_10720,N_9921,N_9260);
nand U10721 (N_10721,N_9991,N_9865);
and U10722 (N_10722,N_9045,N_8995);
nor U10723 (N_10723,N_9955,N_9322);
nand U10724 (N_10724,N_8981,N_9779);
xnor U10725 (N_10725,N_9616,N_9098);
or U10726 (N_10726,N_9390,N_9906);
xor U10727 (N_10727,N_8880,N_8940);
and U10728 (N_10728,N_9617,N_9580);
or U10729 (N_10729,N_9238,N_9684);
nor U10730 (N_10730,N_9826,N_8815);
xor U10731 (N_10731,N_9066,N_9782);
or U10732 (N_10732,N_8841,N_9670);
or U10733 (N_10733,N_8873,N_8980);
and U10734 (N_10734,N_8791,N_9104);
and U10735 (N_10735,N_8835,N_9423);
xor U10736 (N_10736,N_8779,N_9790);
nand U10737 (N_10737,N_9037,N_9891);
and U10738 (N_10738,N_9696,N_8990);
and U10739 (N_10739,N_8907,N_9474);
and U10740 (N_10740,N_8954,N_9102);
or U10741 (N_10741,N_8825,N_9005);
nor U10742 (N_10742,N_9800,N_9574);
or U10743 (N_10743,N_9315,N_9829);
and U10744 (N_10744,N_8823,N_9402);
and U10745 (N_10745,N_8780,N_9132);
nor U10746 (N_10746,N_8867,N_9931);
and U10747 (N_10747,N_8983,N_9490);
and U10748 (N_10748,N_9328,N_9449);
or U10749 (N_10749,N_9872,N_9394);
and U10750 (N_10750,N_9649,N_9621);
and U10751 (N_10751,N_9396,N_8959);
or U10752 (N_10752,N_9030,N_9893);
nor U10753 (N_10753,N_9425,N_9655);
and U10754 (N_10754,N_9618,N_9723);
or U10755 (N_10755,N_9307,N_9915);
or U10756 (N_10756,N_8756,N_8804);
nand U10757 (N_10757,N_9030,N_8988);
and U10758 (N_10758,N_9914,N_9018);
xnor U10759 (N_10759,N_9099,N_9164);
nor U10760 (N_10760,N_8935,N_9490);
and U10761 (N_10761,N_9580,N_9928);
nand U10762 (N_10762,N_9777,N_9019);
and U10763 (N_10763,N_9754,N_8761);
xor U10764 (N_10764,N_9936,N_9943);
or U10765 (N_10765,N_8880,N_9217);
and U10766 (N_10766,N_9140,N_8815);
xnor U10767 (N_10767,N_8921,N_9281);
nor U10768 (N_10768,N_9675,N_9927);
nand U10769 (N_10769,N_8807,N_8863);
xor U10770 (N_10770,N_9348,N_9625);
nor U10771 (N_10771,N_9769,N_9158);
nand U10772 (N_10772,N_9256,N_8834);
nand U10773 (N_10773,N_9796,N_9172);
xnor U10774 (N_10774,N_9524,N_9640);
or U10775 (N_10775,N_9420,N_8974);
xnor U10776 (N_10776,N_9140,N_9950);
nand U10777 (N_10777,N_8886,N_9751);
xnor U10778 (N_10778,N_9809,N_9264);
xor U10779 (N_10779,N_9981,N_9100);
xnor U10780 (N_10780,N_9364,N_9749);
xor U10781 (N_10781,N_9881,N_9581);
and U10782 (N_10782,N_9047,N_9090);
and U10783 (N_10783,N_9186,N_9091);
xnor U10784 (N_10784,N_8896,N_9478);
nor U10785 (N_10785,N_9855,N_9558);
or U10786 (N_10786,N_8976,N_8974);
and U10787 (N_10787,N_8767,N_9896);
or U10788 (N_10788,N_9021,N_9170);
xor U10789 (N_10789,N_8945,N_9011);
nor U10790 (N_10790,N_9063,N_9398);
nor U10791 (N_10791,N_9388,N_8981);
and U10792 (N_10792,N_9595,N_8780);
nand U10793 (N_10793,N_9733,N_8853);
nor U10794 (N_10794,N_9133,N_9724);
and U10795 (N_10795,N_9230,N_9901);
and U10796 (N_10796,N_8997,N_9066);
or U10797 (N_10797,N_9070,N_9557);
xnor U10798 (N_10798,N_9918,N_9293);
or U10799 (N_10799,N_9704,N_9164);
or U10800 (N_10800,N_9600,N_9204);
nand U10801 (N_10801,N_9661,N_9493);
xor U10802 (N_10802,N_9947,N_9838);
nand U10803 (N_10803,N_8980,N_8847);
nor U10804 (N_10804,N_9045,N_9384);
xor U10805 (N_10805,N_9448,N_9275);
and U10806 (N_10806,N_9898,N_9391);
or U10807 (N_10807,N_9444,N_9912);
xor U10808 (N_10808,N_9287,N_9244);
xnor U10809 (N_10809,N_9201,N_9338);
and U10810 (N_10810,N_9114,N_9963);
xor U10811 (N_10811,N_8753,N_9178);
and U10812 (N_10812,N_9110,N_9116);
nand U10813 (N_10813,N_9239,N_8795);
or U10814 (N_10814,N_9517,N_9134);
nand U10815 (N_10815,N_9676,N_9323);
nor U10816 (N_10816,N_9237,N_9458);
nand U10817 (N_10817,N_9536,N_9512);
or U10818 (N_10818,N_9927,N_9504);
xor U10819 (N_10819,N_9281,N_9812);
xor U10820 (N_10820,N_9864,N_9531);
nand U10821 (N_10821,N_9978,N_9560);
nor U10822 (N_10822,N_9633,N_9110);
or U10823 (N_10823,N_9389,N_9035);
or U10824 (N_10824,N_9884,N_9119);
nor U10825 (N_10825,N_9074,N_9932);
and U10826 (N_10826,N_9935,N_9763);
xor U10827 (N_10827,N_9975,N_9144);
xor U10828 (N_10828,N_9322,N_8851);
xor U10829 (N_10829,N_9366,N_9895);
and U10830 (N_10830,N_9397,N_9163);
or U10831 (N_10831,N_8940,N_9965);
nor U10832 (N_10832,N_9563,N_9144);
and U10833 (N_10833,N_9898,N_8950);
and U10834 (N_10834,N_9362,N_9979);
nor U10835 (N_10835,N_9077,N_9577);
and U10836 (N_10836,N_9846,N_9027);
nor U10837 (N_10837,N_9907,N_9843);
and U10838 (N_10838,N_9556,N_8933);
nor U10839 (N_10839,N_9907,N_9786);
or U10840 (N_10840,N_8805,N_9727);
or U10841 (N_10841,N_9766,N_9367);
xnor U10842 (N_10842,N_9385,N_9068);
nor U10843 (N_10843,N_9806,N_9584);
or U10844 (N_10844,N_9043,N_9189);
and U10845 (N_10845,N_9518,N_8847);
nor U10846 (N_10846,N_9310,N_9395);
xnor U10847 (N_10847,N_9991,N_9438);
nand U10848 (N_10848,N_8873,N_9949);
nor U10849 (N_10849,N_8951,N_9231);
xnor U10850 (N_10850,N_9465,N_9913);
xnor U10851 (N_10851,N_9500,N_9401);
xor U10852 (N_10852,N_8882,N_8901);
nor U10853 (N_10853,N_9130,N_9956);
nand U10854 (N_10854,N_8813,N_8902);
or U10855 (N_10855,N_8855,N_8965);
nor U10856 (N_10856,N_9630,N_9353);
nand U10857 (N_10857,N_9738,N_9446);
or U10858 (N_10858,N_9633,N_9643);
and U10859 (N_10859,N_8783,N_9270);
nor U10860 (N_10860,N_9674,N_8775);
nor U10861 (N_10861,N_9426,N_9639);
or U10862 (N_10862,N_9274,N_9172);
and U10863 (N_10863,N_9204,N_9792);
nor U10864 (N_10864,N_9677,N_8828);
or U10865 (N_10865,N_9440,N_9728);
nand U10866 (N_10866,N_9819,N_9785);
or U10867 (N_10867,N_9205,N_9233);
nand U10868 (N_10868,N_9725,N_8782);
xnor U10869 (N_10869,N_9185,N_9298);
nor U10870 (N_10870,N_9875,N_9077);
xnor U10871 (N_10871,N_9551,N_9981);
nor U10872 (N_10872,N_9105,N_8864);
or U10873 (N_10873,N_8893,N_8776);
and U10874 (N_10874,N_9608,N_9726);
or U10875 (N_10875,N_9249,N_9256);
nor U10876 (N_10876,N_9822,N_9493);
nand U10877 (N_10877,N_9996,N_8823);
nor U10878 (N_10878,N_9271,N_9804);
and U10879 (N_10879,N_9658,N_9236);
nand U10880 (N_10880,N_9608,N_9851);
xnor U10881 (N_10881,N_9540,N_9931);
nand U10882 (N_10882,N_9312,N_9553);
or U10883 (N_10883,N_8880,N_8863);
nor U10884 (N_10884,N_9792,N_9968);
nor U10885 (N_10885,N_9921,N_9814);
nor U10886 (N_10886,N_9905,N_9365);
nand U10887 (N_10887,N_9081,N_8992);
or U10888 (N_10888,N_9725,N_9763);
nor U10889 (N_10889,N_9397,N_9677);
nor U10890 (N_10890,N_9929,N_8968);
and U10891 (N_10891,N_9279,N_8845);
and U10892 (N_10892,N_9914,N_9198);
nand U10893 (N_10893,N_9277,N_9430);
xnor U10894 (N_10894,N_9138,N_9855);
xor U10895 (N_10895,N_9600,N_9073);
and U10896 (N_10896,N_9610,N_9917);
or U10897 (N_10897,N_9907,N_8750);
or U10898 (N_10898,N_8764,N_9424);
nor U10899 (N_10899,N_9475,N_9666);
or U10900 (N_10900,N_9116,N_9069);
and U10901 (N_10901,N_9826,N_9857);
xor U10902 (N_10902,N_9458,N_8880);
or U10903 (N_10903,N_9112,N_9376);
and U10904 (N_10904,N_9291,N_8863);
xnor U10905 (N_10905,N_9293,N_9000);
xor U10906 (N_10906,N_9608,N_9538);
and U10907 (N_10907,N_9953,N_9043);
nand U10908 (N_10908,N_9689,N_8860);
and U10909 (N_10909,N_8913,N_9287);
nor U10910 (N_10910,N_8961,N_9575);
and U10911 (N_10911,N_9038,N_9022);
nand U10912 (N_10912,N_8797,N_9537);
and U10913 (N_10913,N_9706,N_8993);
or U10914 (N_10914,N_8887,N_9843);
or U10915 (N_10915,N_9612,N_9194);
or U10916 (N_10916,N_8975,N_9064);
and U10917 (N_10917,N_9007,N_9856);
or U10918 (N_10918,N_9949,N_9357);
or U10919 (N_10919,N_9659,N_9236);
nor U10920 (N_10920,N_9123,N_9742);
nor U10921 (N_10921,N_9753,N_9915);
nor U10922 (N_10922,N_9044,N_9401);
xor U10923 (N_10923,N_9391,N_9367);
or U10924 (N_10924,N_9080,N_9854);
nor U10925 (N_10925,N_9178,N_9175);
xnor U10926 (N_10926,N_9058,N_9050);
nor U10927 (N_10927,N_9977,N_9774);
and U10928 (N_10928,N_8876,N_9316);
nor U10929 (N_10929,N_8807,N_9009);
nor U10930 (N_10930,N_9418,N_9207);
and U10931 (N_10931,N_9804,N_9229);
and U10932 (N_10932,N_9698,N_9876);
xor U10933 (N_10933,N_9264,N_9042);
or U10934 (N_10934,N_9852,N_9916);
or U10935 (N_10935,N_8779,N_9620);
and U10936 (N_10936,N_9972,N_9218);
nor U10937 (N_10937,N_9013,N_9789);
or U10938 (N_10938,N_9499,N_9292);
nand U10939 (N_10939,N_9364,N_8881);
and U10940 (N_10940,N_9122,N_9800);
and U10941 (N_10941,N_9129,N_9488);
nor U10942 (N_10942,N_9267,N_8851);
or U10943 (N_10943,N_9152,N_9123);
and U10944 (N_10944,N_9057,N_9496);
xnor U10945 (N_10945,N_9140,N_9554);
or U10946 (N_10946,N_9932,N_9544);
and U10947 (N_10947,N_9449,N_9734);
nor U10948 (N_10948,N_8966,N_8964);
nor U10949 (N_10949,N_9108,N_8941);
and U10950 (N_10950,N_8851,N_9303);
nor U10951 (N_10951,N_9318,N_9952);
nor U10952 (N_10952,N_9625,N_9250);
xnor U10953 (N_10953,N_8897,N_8829);
and U10954 (N_10954,N_8887,N_8794);
and U10955 (N_10955,N_9373,N_9640);
xor U10956 (N_10956,N_9639,N_8920);
nand U10957 (N_10957,N_9812,N_8931);
xor U10958 (N_10958,N_8767,N_9912);
or U10959 (N_10959,N_8938,N_9362);
nor U10960 (N_10960,N_9689,N_9801);
or U10961 (N_10961,N_9752,N_9011);
nor U10962 (N_10962,N_9868,N_9218);
and U10963 (N_10963,N_9676,N_8905);
xor U10964 (N_10964,N_9486,N_9672);
nor U10965 (N_10965,N_8966,N_9026);
nor U10966 (N_10966,N_9872,N_9603);
or U10967 (N_10967,N_9756,N_9211);
and U10968 (N_10968,N_8855,N_9863);
nor U10969 (N_10969,N_9254,N_9031);
nor U10970 (N_10970,N_9438,N_9162);
or U10971 (N_10971,N_9558,N_9901);
and U10972 (N_10972,N_8881,N_9545);
or U10973 (N_10973,N_9985,N_9212);
xnor U10974 (N_10974,N_8755,N_9999);
nor U10975 (N_10975,N_9779,N_8877);
or U10976 (N_10976,N_9971,N_9935);
nor U10977 (N_10977,N_9616,N_9956);
xor U10978 (N_10978,N_9755,N_8905);
or U10979 (N_10979,N_9161,N_9415);
or U10980 (N_10980,N_9870,N_9276);
or U10981 (N_10981,N_9880,N_9812);
nor U10982 (N_10982,N_9747,N_9073);
nor U10983 (N_10983,N_9163,N_9729);
xor U10984 (N_10984,N_9079,N_9039);
nor U10985 (N_10985,N_9792,N_9794);
xnor U10986 (N_10986,N_9017,N_8773);
and U10987 (N_10987,N_9148,N_9153);
and U10988 (N_10988,N_9830,N_9287);
or U10989 (N_10989,N_9959,N_8945);
nand U10990 (N_10990,N_9015,N_8761);
nand U10991 (N_10991,N_9015,N_9370);
xor U10992 (N_10992,N_9625,N_9057);
nor U10993 (N_10993,N_8866,N_9394);
and U10994 (N_10994,N_9283,N_9239);
or U10995 (N_10995,N_9381,N_9670);
nor U10996 (N_10996,N_9952,N_9849);
or U10997 (N_10997,N_8935,N_9699);
nand U10998 (N_10998,N_9293,N_9171);
nor U10999 (N_10999,N_9045,N_9215);
nor U11000 (N_11000,N_9724,N_9823);
or U11001 (N_11001,N_8856,N_9742);
and U11002 (N_11002,N_8867,N_9261);
nand U11003 (N_11003,N_9501,N_9033);
and U11004 (N_11004,N_9205,N_8815);
xor U11005 (N_11005,N_9202,N_9164);
or U11006 (N_11006,N_9250,N_9999);
nor U11007 (N_11007,N_9345,N_9599);
or U11008 (N_11008,N_9103,N_9285);
nand U11009 (N_11009,N_9473,N_9367);
or U11010 (N_11010,N_8797,N_8837);
or U11011 (N_11011,N_8940,N_9566);
or U11012 (N_11012,N_9829,N_9612);
nand U11013 (N_11013,N_9354,N_9040);
nand U11014 (N_11014,N_9996,N_8937);
and U11015 (N_11015,N_9279,N_9216);
nand U11016 (N_11016,N_9627,N_8829);
and U11017 (N_11017,N_9636,N_9868);
nor U11018 (N_11018,N_9606,N_8865);
and U11019 (N_11019,N_9621,N_9485);
nand U11020 (N_11020,N_8860,N_9905);
and U11021 (N_11021,N_9997,N_9987);
xor U11022 (N_11022,N_9171,N_8895);
xor U11023 (N_11023,N_8979,N_9914);
and U11024 (N_11024,N_9625,N_8978);
nand U11025 (N_11025,N_8796,N_9535);
and U11026 (N_11026,N_9927,N_9013);
nor U11027 (N_11027,N_9224,N_9784);
and U11028 (N_11028,N_9118,N_9198);
nand U11029 (N_11029,N_9061,N_9471);
nand U11030 (N_11030,N_9083,N_9885);
nor U11031 (N_11031,N_9550,N_9276);
nor U11032 (N_11032,N_9740,N_9685);
nor U11033 (N_11033,N_9987,N_9540);
and U11034 (N_11034,N_9389,N_9327);
nand U11035 (N_11035,N_9658,N_9255);
nor U11036 (N_11036,N_9733,N_9524);
or U11037 (N_11037,N_9960,N_8807);
and U11038 (N_11038,N_9266,N_9113);
or U11039 (N_11039,N_9755,N_9332);
xnor U11040 (N_11040,N_9488,N_9573);
xnor U11041 (N_11041,N_9512,N_9478);
nand U11042 (N_11042,N_9209,N_9187);
or U11043 (N_11043,N_8794,N_9547);
nand U11044 (N_11044,N_9062,N_8935);
and U11045 (N_11045,N_9725,N_9070);
nor U11046 (N_11046,N_9139,N_9000);
nand U11047 (N_11047,N_8795,N_9134);
and U11048 (N_11048,N_9635,N_9274);
nor U11049 (N_11049,N_9685,N_9705);
xnor U11050 (N_11050,N_9165,N_8838);
nor U11051 (N_11051,N_9645,N_9635);
nand U11052 (N_11052,N_8773,N_8774);
xor U11053 (N_11053,N_9769,N_9248);
or U11054 (N_11054,N_9027,N_9971);
nand U11055 (N_11055,N_9935,N_9142);
nand U11056 (N_11056,N_9442,N_9832);
and U11057 (N_11057,N_9859,N_9910);
nor U11058 (N_11058,N_9412,N_9597);
and U11059 (N_11059,N_9062,N_9252);
xnor U11060 (N_11060,N_9977,N_9319);
or U11061 (N_11061,N_9985,N_9821);
nor U11062 (N_11062,N_9912,N_9407);
and U11063 (N_11063,N_9028,N_9025);
nor U11064 (N_11064,N_9415,N_8761);
nor U11065 (N_11065,N_9901,N_9008);
nand U11066 (N_11066,N_8817,N_8926);
nor U11067 (N_11067,N_9856,N_9751);
nor U11068 (N_11068,N_8759,N_8985);
or U11069 (N_11069,N_9580,N_9098);
nor U11070 (N_11070,N_8753,N_9841);
xnor U11071 (N_11071,N_9037,N_9831);
or U11072 (N_11072,N_9595,N_9760);
and U11073 (N_11073,N_9622,N_9398);
nand U11074 (N_11074,N_9660,N_9006);
nor U11075 (N_11075,N_9674,N_9682);
nand U11076 (N_11076,N_9889,N_8769);
and U11077 (N_11077,N_8886,N_9353);
nand U11078 (N_11078,N_8774,N_9809);
nor U11079 (N_11079,N_9422,N_9271);
nor U11080 (N_11080,N_9549,N_9521);
xor U11081 (N_11081,N_9912,N_8827);
or U11082 (N_11082,N_9721,N_9503);
nand U11083 (N_11083,N_9649,N_9062);
nor U11084 (N_11084,N_9029,N_9011);
or U11085 (N_11085,N_9255,N_9520);
nor U11086 (N_11086,N_8917,N_9793);
nand U11087 (N_11087,N_9110,N_8751);
nor U11088 (N_11088,N_8983,N_9717);
xnor U11089 (N_11089,N_8810,N_8880);
or U11090 (N_11090,N_8991,N_9461);
xnor U11091 (N_11091,N_9679,N_9897);
xnor U11092 (N_11092,N_8994,N_9268);
nor U11093 (N_11093,N_9697,N_9051);
and U11094 (N_11094,N_9466,N_9141);
or U11095 (N_11095,N_9008,N_9786);
nand U11096 (N_11096,N_8782,N_8836);
nand U11097 (N_11097,N_8862,N_8852);
nor U11098 (N_11098,N_9520,N_9541);
nor U11099 (N_11099,N_9542,N_9392);
xor U11100 (N_11100,N_9315,N_9288);
and U11101 (N_11101,N_9364,N_8987);
nor U11102 (N_11102,N_9613,N_8827);
nand U11103 (N_11103,N_9054,N_9304);
nand U11104 (N_11104,N_9564,N_9338);
or U11105 (N_11105,N_9084,N_9508);
nand U11106 (N_11106,N_8910,N_8957);
and U11107 (N_11107,N_8794,N_9556);
nand U11108 (N_11108,N_9600,N_9643);
nor U11109 (N_11109,N_9706,N_9201);
or U11110 (N_11110,N_8862,N_9313);
xor U11111 (N_11111,N_9740,N_8951);
nand U11112 (N_11112,N_9657,N_8898);
and U11113 (N_11113,N_9434,N_9541);
nor U11114 (N_11114,N_8881,N_8894);
or U11115 (N_11115,N_9794,N_9685);
nor U11116 (N_11116,N_8859,N_9506);
xor U11117 (N_11117,N_9741,N_9752);
nand U11118 (N_11118,N_9997,N_9921);
nor U11119 (N_11119,N_9103,N_9357);
or U11120 (N_11120,N_9211,N_9290);
nand U11121 (N_11121,N_8935,N_8969);
nand U11122 (N_11122,N_9062,N_8831);
or U11123 (N_11123,N_9982,N_9901);
or U11124 (N_11124,N_9045,N_9582);
nand U11125 (N_11125,N_9012,N_9191);
nor U11126 (N_11126,N_9262,N_9129);
or U11127 (N_11127,N_9174,N_9519);
and U11128 (N_11128,N_9123,N_9360);
xor U11129 (N_11129,N_9713,N_8910);
nor U11130 (N_11130,N_9624,N_9928);
and U11131 (N_11131,N_9356,N_9416);
xor U11132 (N_11132,N_9943,N_9960);
nand U11133 (N_11133,N_9861,N_9574);
and U11134 (N_11134,N_9661,N_8882);
nand U11135 (N_11135,N_9488,N_9826);
or U11136 (N_11136,N_9962,N_9306);
nor U11137 (N_11137,N_9418,N_9333);
xor U11138 (N_11138,N_9469,N_9914);
xor U11139 (N_11139,N_8964,N_9654);
nand U11140 (N_11140,N_9867,N_9568);
and U11141 (N_11141,N_9236,N_9977);
nor U11142 (N_11142,N_9532,N_9346);
nor U11143 (N_11143,N_9646,N_9143);
xnor U11144 (N_11144,N_9709,N_8948);
and U11145 (N_11145,N_9726,N_9165);
xnor U11146 (N_11146,N_9367,N_9316);
nor U11147 (N_11147,N_9471,N_9083);
nand U11148 (N_11148,N_8778,N_9653);
xnor U11149 (N_11149,N_9633,N_9570);
xnor U11150 (N_11150,N_9729,N_9686);
nor U11151 (N_11151,N_9838,N_9467);
and U11152 (N_11152,N_9803,N_8984);
nor U11153 (N_11153,N_9063,N_9459);
nand U11154 (N_11154,N_8803,N_9907);
nand U11155 (N_11155,N_9383,N_9926);
nor U11156 (N_11156,N_9143,N_8857);
and U11157 (N_11157,N_9803,N_9552);
nand U11158 (N_11158,N_9329,N_8898);
nor U11159 (N_11159,N_9377,N_9417);
or U11160 (N_11160,N_9969,N_9487);
nor U11161 (N_11161,N_9641,N_9455);
or U11162 (N_11162,N_9856,N_9655);
or U11163 (N_11163,N_9179,N_9209);
and U11164 (N_11164,N_9594,N_9632);
and U11165 (N_11165,N_9908,N_8852);
xnor U11166 (N_11166,N_8893,N_8864);
and U11167 (N_11167,N_9365,N_8979);
nor U11168 (N_11168,N_8899,N_9307);
and U11169 (N_11169,N_9906,N_9118);
and U11170 (N_11170,N_8809,N_8892);
nor U11171 (N_11171,N_8810,N_8780);
xor U11172 (N_11172,N_9972,N_9853);
nand U11173 (N_11173,N_9773,N_9990);
nand U11174 (N_11174,N_8968,N_9632);
nand U11175 (N_11175,N_8981,N_9221);
nor U11176 (N_11176,N_8904,N_9224);
or U11177 (N_11177,N_9466,N_9236);
nor U11178 (N_11178,N_9595,N_9829);
and U11179 (N_11179,N_9620,N_9563);
nand U11180 (N_11180,N_9455,N_9763);
or U11181 (N_11181,N_9309,N_9418);
nand U11182 (N_11182,N_9280,N_8872);
xnor U11183 (N_11183,N_8872,N_9525);
xor U11184 (N_11184,N_9522,N_9798);
nand U11185 (N_11185,N_8841,N_9488);
nand U11186 (N_11186,N_9865,N_9910);
or U11187 (N_11187,N_9418,N_9294);
nand U11188 (N_11188,N_9058,N_9801);
nand U11189 (N_11189,N_9426,N_9843);
or U11190 (N_11190,N_9381,N_8773);
or U11191 (N_11191,N_8798,N_9977);
nand U11192 (N_11192,N_9825,N_9351);
or U11193 (N_11193,N_9921,N_8928);
nor U11194 (N_11194,N_9017,N_9344);
and U11195 (N_11195,N_9108,N_9650);
xor U11196 (N_11196,N_9415,N_8985);
and U11197 (N_11197,N_9290,N_9957);
nor U11198 (N_11198,N_9622,N_9023);
nand U11199 (N_11199,N_9149,N_9405);
xnor U11200 (N_11200,N_9956,N_9904);
nand U11201 (N_11201,N_9809,N_8783);
nand U11202 (N_11202,N_8884,N_9551);
and U11203 (N_11203,N_9283,N_8859);
xnor U11204 (N_11204,N_9054,N_8933);
nand U11205 (N_11205,N_9591,N_9869);
xnor U11206 (N_11206,N_9099,N_9817);
nand U11207 (N_11207,N_9394,N_9496);
nor U11208 (N_11208,N_9368,N_9757);
xnor U11209 (N_11209,N_9961,N_8807);
nand U11210 (N_11210,N_9721,N_8766);
nand U11211 (N_11211,N_9653,N_9048);
or U11212 (N_11212,N_9436,N_9831);
nor U11213 (N_11213,N_9687,N_9156);
and U11214 (N_11214,N_9746,N_9255);
and U11215 (N_11215,N_9987,N_8922);
nand U11216 (N_11216,N_9155,N_9859);
and U11217 (N_11217,N_8937,N_9483);
and U11218 (N_11218,N_8946,N_8821);
nor U11219 (N_11219,N_9058,N_9033);
nor U11220 (N_11220,N_8827,N_9981);
and U11221 (N_11221,N_9281,N_9116);
nor U11222 (N_11222,N_9935,N_9639);
xnor U11223 (N_11223,N_9293,N_9581);
xnor U11224 (N_11224,N_9631,N_8804);
nor U11225 (N_11225,N_9066,N_9650);
nor U11226 (N_11226,N_9717,N_9550);
nor U11227 (N_11227,N_8842,N_9127);
nand U11228 (N_11228,N_9436,N_9452);
nand U11229 (N_11229,N_9898,N_8852);
nor U11230 (N_11230,N_9183,N_8954);
nand U11231 (N_11231,N_8963,N_9527);
nand U11232 (N_11232,N_8948,N_9393);
nand U11233 (N_11233,N_9697,N_9053);
nor U11234 (N_11234,N_8823,N_9612);
xor U11235 (N_11235,N_9093,N_9993);
nor U11236 (N_11236,N_9197,N_8868);
or U11237 (N_11237,N_8902,N_8814);
nor U11238 (N_11238,N_9484,N_9361);
nand U11239 (N_11239,N_9599,N_9429);
xnor U11240 (N_11240,N_9052,N_9961);
or U11241 (N_11241,N_9953,N_9954);
and U11242 (N_11242,N_9309,N_9334);
xnor U11243 (N_11243,N_9162,N_8896);
and U11244 (N_11244,N_8764,N_9578);
or U11245 (N_11245,N_8812,N_8919);
and U11246 (N_11246,N_9796,N_9879);
xor U11247 (N_11247,N_8767,N_8802);
nor U11248 (N_11248,N_9160,N_9915);
and U11249 (N_11249,N_8844,N_9182);
or U11250 (N_11250,N_10078,N_10902);
nor U11251 (N_11251,N_11167,N_10463);
nand U11252 (N_11252,N_10300,N_10788);
xor U11253 (N_11253,N_10830,N_10392);
and U11254 (N_11254,N_10688,N_11057);
or U11255 (N_11255,N_10455,N_11117);
nand U11256 (N_11256,N_10964,N_10292);
xor U11257 (N_11257,N_10501,N_10053);
xor U11258 (N_11258,N_10440,N_10293);
nor U11259 (N_11259,N_10593,N_10510);
xnor U11260 (N_11260,N_10175,N_10312);
nand U11261 (N_11261,N_10196,N_10228);
xnor U11262 (N_11262,N_11048,N_10184);
nor U11263 (N_11263,N_10426,N_10948);
nor U11264 (N_11264,N_10191,N_10225);
nand U11265 (N_11265,N_11190,N_10767);
nor U11266 (N_11266,N_10277,N_10558);
nand U11267 (N_11267,N_11075,N_11141);
and U11268 (N_11268,N_10047,N_10739);
nor U11269 (N_11269,N_10282,N_10405);
xnor U11270 (N_11270,N_10007,N_10816);
nor U11271 (N_11271,N_10470,N_10077);
and U11272 (N_11272,N_10853,N_10142);
or U11273 (N_11273,N_10466,N_11028);
nand U11274 (N_11274,N_10143,N_10779);
or U11275 (N_11275,N_10984,N_10321);
xor U11276 (N_11276,N_10546,N_10704);
and U11277 (N_11277,N_10591,N_10805);
nor U11278 (N_11278,N_10900,N_10492);
nand U11279 (N_11279,N_10766,N_10869);
nor U11280 (N_11280,N_10967,N_11245);
nand U11281 (N_11281,N_11180,N_10682);
nand U11282 (N_11282,N_10423,N_10696);
and U11283 (N_11283,N_11072,N_10118);
nand U11284 (N_11284,N_10317,N_10679);
or U11285 (N_11285,N_11225,N_10460);
nand U11286 (N_11286,N_10004,N_10429);
nor U11287 (N_11287,N_11202,N_10016);
xor U11288 (N_11288,N_10777,N_10486);
and U11289 (N_11289,N_11157,N_10488);
xnor U11290 (N_11290,N_10410,N_10462);
nand U11291 (N_11291,N_10549,N_10562);
nand U11292 (N_11292,N_10132,N_10314);
xnor U11293 (N_11293,N_10275,N_10122);
nand U11294 (N_11294,N_10947,N_10961);
nand U11295 (N_11295,N_10394,N_11034);
nor U11296 (N_11296,N_11161,N_10059);
nand U11297 (N_11297,N_10261,N_10815);
xnor U11298 (N_11298,N_10834,N_10190);
xnor U11299 (N_11299,N_11095,N_10038);
xor U11300 (N_11300,N_10083,N_11042);
and U11301 (N_11301,N_10071,N_10559);
nor U11302 (N_11302,N_11077,N_11114);
nand U11303 (N_11303,N_10491,N_10588);
nor U11304 (N_11304,N_11206,N_10454);
nor U11305 (N_11305,N_10754,N_10750);
and U11306 (N_11306,N_10039,N_11145);
xor U11307 (N_11307,N_10082,N_11195);
nand U11308 (N_11308,N_10407,N_10691);
or U11309 (N_11309,N_10844,N_10453);
xnor U11310 (N_11310,N_11239,N_10623);
and U11311 (N_11311,N_10298,N_11104);
nor U11312 (N_11312,N_10425,N_10345);
and U11313 (N_11313,N_11099,N_10305);
or U11314 (N_11314,N_11128,N_10302);
xnor U11315 (N_11315,N_10269,N_10189);
or U11316 (N_11316,N_10320,N_11199);
or U11317 (N_11317,N_10852,N_10450);
nor U11318 (N_11318,N_10433,N_10380);
nand U11319 (N_11319,N_10945,N_10791);
xnor U11320 (N_11320,N_10010,N_11210);
and U11321 (N_11321,N_10698,N_10829);
and U11322 (N_11322,N_11040,N_11170);
nand U11323 (N_11323,N_11232,N_10678);
or U11324 (N_11324,N_10362,N_10036);
nor U11325 (N_11325,N_10862,N_10249);
nor U11326 (N_11326,N_10182,N_10612);
nor U11327 (N_11327,N_11159,N_11220);
nor U11328 (N_11328,N_10119,N_10699);
nor U11329 (N_11329,N_10213,N_10656);
xnor U11330 (N_11330,N_10290,N_10280);
nor U11331 (N_11331,N_10103,N_10733);
and U11332 (N_11332,N_10875,N_10795);
nand U11333 (N_11333,N_10333,N_10975);
nor U11334 (N_11334,N_10776,N_11038);
and U11335 (N_11335,N_10346,N_10437);
xor U11336 (N_11336,N_11196,N_10056);
or U11337 (N_11337,N_10157,N_10540);
or U11338 (N_11338,N_10839,N_10605);
and U11339 (N_11339,N_11152,N_10657);
and U11340 (N_11340,N_10670,N_10564);
xor U11341 (N_11341,N_10896,N_10895);
nand U11342 (N_11342,N_10914,N_10404);
or U11343 (N_11343,N_10354,N_10397);
nor U11344 (N_11344,N_10114,N_10181);
nand U11345 (N_11345,N_10563,N_10057);
xnor U11346 (N_11346,N_10744,N_11050);
nand U11347 (N_11347,N_10028,N_10512);
nor U11348 (N_11348,N_11203,N_10718);
nand U11349 (N_11349,N_10993,N_10673);
nor U11350 (N_11350,N_10411,N_10216);
nand U11351 (N_11351,N_11115,N_11069);
nand U11352 (N_11352,N_10515,N_11148);
nand U11353 (N_11353,N_10538,N_10168);
nor U11354 (N_11354,N_10921,N_10624);
nand U11355 (N_11355,N_10652,N_10307);
or U11356 (N_11356,N_11108,N_11226);
or U11357 (N_11357,N_10838,N_10409);
nand U11358 (N_11358,N_10797,N_11123);
and U11359 (N_11359,N_10891,N_10676);
nor U11360 (N_11360,N_11020,N_10927);
xor U11361 (N_11361,N_11032,N_10813);
or U11362 (N_11362,N_10703,N_10257);
nand U11363 (N_11363,N_10369,N_10901);
xor U11364 (N_11364,N_11061,N_10390);
nor U11365 (N_11365,N_10044,N_10179);
nor U11366 (N_11366,N_10522,N_10729);
and U11367 (N_11367,N_10536,N_10490);
or U11368 (N_11368,N_10887,N_10582);
or U11369 (N_11369,N_10357,N_10185);
nor U11370 (N_11370,N_10669,N_10903);
or U11371 (N_11371,N_10343,N_10640);
and U11372 (N_11372,N_11213,N_11146);
and U11373 (N_11373,N_10498,N_10121);
nor U11374 (N_11374,N_11055,N_10263);
or U11375 (N_11375,N_10606,N_10929);
nand U11376 (N_11376,N_11150,N_10758);
or U11377 (N_11377,N_11184,N_10169);
nand U11378 (N_11378,N_11086,N_10291);
nand U11379 (N_11379,N_10924,N_10417);
xor U11380 (N_11380,N_10738,N_11139);
and U11381 (N_11381,N_10659,N_10211);
nor U11382 (N_11382,N_11087,N_10867);
and U11383 (N_11383,N_10660,N_10684);
nor U11384 (N_11384,N_10322,N_11124);
nor U11385 (N_11385,N_11079,N_11031);
nor U11386 (N_11386,N_10988,N_10804);
and U11387 (N_11387,N_10937,N_11004);
xor U11388 (N_11388,N_10388,N_11238);
nand U11389 (N_11389,N_10099,N_10458);
xor U11390 (N_11390,N_10446,N_10372);
and U11391 (N_11391,N_11097,N_10285);
nor U11392 (N_11392,N_10013,N_10907);
or U11393 (N_11393,N_10422,N_10974);
nor U11394 (N_11394,N_10205,N_10585);
nor U11395 (N_11395,N_10551,N_10812);
or U11396 (N_11396,N_10529,N_10613);
xor U11397 (N_11397,N_10557,N_10434);
and U11398 (N_11398,N_10970,N_10928);
xor U11399 (N_11399,N_11029,N_10267);
or U11400 (N_11400,N_11191,N_10416);
and U11401 (N_11401,N_11222,N_10756);
nor U11402 (N_11402,N_10101,N_11235);
nor U11403 (N_11403,N_10186,N_10352);
nand U11404 (N_11404,N_10857,N_10552);
xor U11405 (N_11405,N_10435,N_10811);
nor U11406 (N_11406,N_10637,N_10570);
and U11407 (N_11407,N_10835,N_11024);
nand U11408 (N_11408,N_10759,N_11130);
nand U11409 (N_11409,N_10148,N_10134);
xnor U11410 (N_11410,N_10006,N_10802);
nand U11411 (N_11411,N_10959,N_11112);
or U11412 (N_11412,N_10939,N_11081);
nor U11413 (N_11413,N_11151,N_10874);
nor U11414 (N_11414,N_11240,N_11092);
and U11415 (N_11415,N_10527,N_10609);
nand U11416 (N_11416,N_11053,N_10859);
and U11417 (N_11417,N_10803,N_10824);
and U11418 (N_11418,N_10663,N_10932);
and U11419 (N_11419,N_10725,N_11143);
xnor U11420 (N_11420,N_11074,N_10452);
xor U11421 (N_11421,N_11094,N_10368);
or U11422 (N_11422,N_10035,N_10722);
and U11423 (N_11423,N_10897,N_10913);
or U11424 (N_11424,N_10164,N_11192);
nand U11425 (N_11425,N_10560,N_10051);
nor U11426 (N_11426,N_10218,N_10861);
or U11427 (N_11427,N_10478,N_10431);
or U11428 (N_11428,N_10638,N_10001);
nor U11429 (N_11429,N_10230,N_10719);
and U11430 (N_11430,N_10209,N_10172);
xnor U11431 (N_11431,N_10781,N_11140);
nand U11432 (N_11432,N_10294,N_10573);
xor U11433 (N_11433,N_10479,N_10383);
nand U11434 (N_11434,N_10949,N_11037);
nor U11435 (N_11435,N_10705,N_10342);
and U11436 (N_11436,N_10286,N_10787);
or U11437 (N_11437,N_11118,N_10145);
xor U11438 (N_11438,N_10432,N_11105);
and U11439 (N_11439,N_11243,N_10589);
or U11440 (N_11440,N_10086,N_10014);
nand U11441 (N_11441,N_10850,N_10151);
xor U11442 (N_11442,N_10761,N_10012);
xnor U11443 (N_11443,N_10100,N_11223);
xor U11444 (N_11444,N_10938,N_10757);
or U11445 (N_11445,N_10910,N_10135);
and U11446 (N_11446,N_10102,N_10576);
nand U11447 (N_11447,N_10689,N_10849);
nor U11448 (N_11448,N_10614,N_10441);
xnor U11449 (N_11449,N_10306,N_10260);
and U11450 (N_11450,N_10973,N_10942);
xnor U11451 (N_11451,N_10129,N_10325);
or U11452 (N_11452,N_10675,N_10344);
or U11453 (N_11453,N_10634,N_10518);
nand U11454 (N_11454,N_10076,N_10149);
xor U11455 (N_11455,N_11162,N_11051);
nand U11456 (N_11456,N_11135,N_10885);
xnor U11457 (N_11457,N_10626,N_11197);
and U11458 (N_11458,N_10052,N_10532);
and U11459 (N_11459,N_10604,N_10063);
xnor U11460 (N_11460,N_10860,N_10141);
and U11461 (N_11461,N_11103,N_10116);
and U11462 (N_11462,N_10138,N_10365);
nand U11463 (N_11463,N_10265,N_10930);
xnor U11464 (N_11464,N_10769,N_11100);
nor U11465 (N_11465,N_10027,N_11006);
or U11466 (N_11466,N_10414,N_11198);
and U11467 (N_11467,N_10655,N_10156);
or U11468 (N_11468,N_10319,N_10093);
nor U11469 (N_11469,N_10413,N_10537);
xnor U11470 (N_11470,N_11026,N_10533);
nor U11471 (N_11471,N_10926,N_10996);
and U11472 (N_11472,N_10192,N_10109);
nor U11473 (N_11473,N_10734,N_11212);
nor U11474 (N_11474,N_10273,N_10361);
nand U11475 (N_11475,N_10207,N_11083);
xnor U11476 (N_11476,N_10798,N_11169);
xnor U11477 (N_11477,N_10545,N_10284);
nand U11478 (N_11478,N_10107,N_10508);
or U11479 (N_11479,N_11008,N_10117);
xor U11480 (N_11480,N_10889,N_10823);
nor U11481 (N_11481,N_10878,N_10456);
xnor U11482 (N_11482,N_10060,N_10041);
and U11483 (N_11483,N_10105,N_10598);
nor U11484 (N_11484,N_10616,N_10808);
xnor U11485 (N_11485,N_11209,N_10774);
nand U11486 (N_11486,N_10304,N_10943);
or U11487 (N_11487,N_10037,N_10775);
xnor U11488 (N_11488,N_11216,N_10992);
nand U11489 (N_11489,N_10106,N_10918);
or U11490 (N_11490,N_10144,N_10825);
xnor U11491 (N_11491,N_10956,N_10743);
nand U11492 (N_11492,N_10940,N_10893);
nor U11493 (N_11493,N_10922,N_11089);
and U11494 (N_11494,N_10509,N_10665);
xnor U11495 (N_11495,N_10370,N_10448);
nor U11496 (N_11496,N_10229,N_10375);
and U11497 (N_11497,N_10482,N_10055);
nand U11498 (N_11498,N_10746,N_10647);
and U11499 (N_11499,N_10318,N_10627);
or U11500 (N_11500,N_10310,N_10166);
or U11501 (N_11501,N_10247,N_10176);
and U11502 (N_11502,N_10313,N_10295);
nand U11503 (N_11503,N_10474,N_11088);
nand U11504 (N_11504,N_10752,N_10040);
and U11505 (N_11505,N_10385,N_10188);
and U11506 (N_11506,N_10994,N_10584);
nand U11507 (N_11507,N_10534,N_10341);
xnor U11508 (N_11508,N_10672,N_10223);
or U11509 (N_11509,N_10485,N_10111);
nand U11510 (N_11510,N_11023,N_10108);
nor U11511 (N_11511,N_10695,N_10617);
nor U11512 (N_11512,N_10873,N_10906);
nor U11513 (N_11513,N_10778,N_10991);
or U11514 (N_11514,N_10140,N_10421);
nor U11515 (N_11515,N_10240,N_10931);
nor U11516 (N_11516,N_10309,N_11147);
or U11517 (N_11517,N_10990,N_10256);
and U11518 (N_11518,N_10773,N_11237);
and U11519 (N_11519,N_10625,N_10245);
nand U11520 (N_11520,N_10858,N_10045);
xnor U11521 (N_11521,N_10832,N_10234);
nor U11522 (N_11522,N_10000,N_10236);
nor U11523 (N_11523,N_11013,N_10771);
nor U11524 (N_11524,N_10124,N_10387);
and U11525 (N_11525,N_10221,N_10566);
nand U11526 (N_11526,N_10976,N_10170);
or U11527 (N_11527,N_11085,N_10800);
nor U11528 (N_11528,N_10794,N_10917);
and U11529 (N_11529,N_10382,N_10713);
nand U11530 (N_11530,N_11018,N_10015);
xor U11531 (N_11531,N_10712,N_10158);
or U11532 (N_11532,N_10279,N_10630);
nand U11533 (N_11533,N_10098,N_10768);
xnor U11534 (N_11534,N_10898,N_10952);
nand U11535 (N_11535,N_10371,N_10396);
xnor U11536 (N_11536,N_10894,N_10685);
nand U11537 (N_11537,N_10619,N_10567);
xnor U11538 (N_11538,N_10031,N_10330);
xor U11539 (N_11539,N_10694,N_10868);
nor U11540 (N_11540,N_10554,N_10074);
nor U11541 (N_11541,N_10565,N_10180);
and U11542 (N_11542,N_10595,N_10528);
nor U11543 (N_11543,N_10841,N_10246);
and U11544 (N_11544,N_10139,N_10005);
nand U11545 (N_11545,N_11136,N_11166);
xnor U11546 (N_11546,N_10643,N_10373);
and U11547 (N_11547,N_10258,N_10415);
nand U11548 (N_11548,N_11021,N_10658);
nor U11549 (N_11549,N_10402,N_10755);
nor U11550 (N_11550,N_11035,N_10200);
or U11551 (N_11551,N_10535,N_11084);
nand U11552 (N_11552,N_10908,N_10977);
or U11553 (N_11553,N_10473,N_10715);
xnor U11554 (N_11554,N_10097,N_10241);
nor U11555 (N_11555,N_10586,N_10243);
and U11556 (N_11556,N_11082,N_10995);
or U11557 (N_11557,N_11054,N_10706);
or U11558 (N_11558,N_10748,N_10217);
xor U11559 (N_11559,N_11153,N_10731);
nand U11560 (N_11560,N_10963,N_10814);
or U11561 (N_11561,N_10709,N_10308);
and U11562 (N_11562,N_10519,N_10592);
xnor U11563 (N_11563,N_10187,N_10870);
nor U11564 (N_11564,N_10198,N_10541);
nor U11565 (N_11565,N_11000,N_11224);
xor U11566 (N_11566,N_10270,N_10631);
nor U11567 (N_11567,N_10299,N_11070);
or U11568 (N_11568,N_10328,N_10096);
nor U11569 (N_11569,N_10760,N_10222);
xor U11570 (N_11570,N_10274,N_11211);
nor U11571 (N_11571,N_10762,N_10475);
nand U11572 (N_11572,N_10951,N_10842);
and U11573 (N_11573,N_11076,N_11236);
nor U11574 (N_11574,N_10153,N_10581);
xnor U11575 (N_11575,N_10863,N_11012);
nand U11576 (N_11576,N_10851,N_10472);
nand U11577 (N_11577,N_10547,N_10866);
and U11578 (N_11578,N_10377,N_10502);
or U11579 (N_11579,N_10747,N_10026);
xor U11580 (N_11580,N_10311,N_10381);
or U11581 (N_11581,N_11144,N_10367);
or U11582 (N_11582,N_11046,N_10395);
xor U11583 (N_11583,N_10215,N_11110);
and U11584 (N_11584,N_11007,N_10772);
xor U11585 (N_11585,N_10253,N_10661);
nand U11586 (N_11586,N_10130,N_10120);
xor U11587 (N_11587,N_10208,N_10648);
nor U11588 (N_11588,N_10792,N_10666);
nand U11589 (N_11589,N_10935,N_10981);
or U11590 (N_11590,N_10030,N_10461);
xor U11591 (N_11591,N_10543,N_10248);
or U11592 (N_11592,N_10194,N_10969);
xnor U11593 (N_11593,N_10481,N_10524);
nand U11594 (N_11594,N_10810,N_10701);
and U11595 (N_11595,N_10050,N_10818);
nand U11596 (N_11596,N_11016,N_10262);
and U11597 (N_11597,N_10464,N_11163);
xor U11598 (N_11598,N_10183,N_11189);
nand U11599 (N_11599,N_10193,N_10687);
xor U11600 (N_11600,N_10468,N_10112);
or U11601 (N_11601,N_11119,N_10329);
nand U11602 (N_11602,N_10629,N_10058);
nand U11603 (N_11603,N_11096,N_10064);
or U11604 (N_11604,N_10572,N_10989);
nor U11605 (N_11605,N_11068,N_10436);
xor U11606 (N_11606,N_10674,N_10686);
and U11607 (N_11607,N_10548,N_11073);
xor U11608 (N_11608,N_11207,N_10590);
nor U11609 (N_11609,N_11080,N_10459);
nor U11610 (N_11610,N_11044,N_10556);
xnor U11611 (N_11611,N_10649,N_11227);
nor U11612 (N_11612,N_10427,N_11045);
or U11613 (N_11613,N_10062,N_11091);
nor U11614 (N_11614,N_10316,N_10578);
nand U11615 (N_11615,N_10732,N_10819);
xor U11616 (N_11616,N_10641,N_10020);
nand U11617 (N_11617,N_10065,N_10671);
nor U11618 (N_11618,N_10278,N_10982);
nand U11619 (N_11619,N_11134,N_11175);
xnor U11620 (N_11620,N_10968,N_10206);
or U11621 (N_11621,N_10363,N_10113);
or U11622 (N_11622,N_10358,N_10780);
and U11623 (N_11623,N_10327,N_10919);
or U11624 (N_11624,N_11058,N_10296);
nand U11625 (N_11625,N_10710,N_11234);
nor U11626 (N_11626,N_11160,N_10338);
and U11627 (N_11627,N_10827,N_10480);
xnor U11628 (N_11628,N_10882,N_10049);
or U11629 (N_11629,N_10272,N_10214);
and U11630 (N_11630,N_11177,N_10763);
nor U11631 (N_11631,N_10347,N_10334);
or U11632 (N_11632,N_11138,N_10561);
xor U11633 (N_11633,N_11186,N_10525);
or U11634 (N_11634,N_10493,N_10177);
nor U11635 (N_11635,N_10268,N_10024);
and U11636 (N_11636,N_10070,N_10043);
nor U11637 (N_11637,N_10946,N_10697);
and U11638 (N_11638,N_11248,N_11027);
nand U11639 (N_11639,N_10171,N_10276);
or U11640 (N_11640,N_10611,N_11228);
or U11641 (N_11641,N_10128,N_11231);
and U11642 (N_11642,N_10855,N_10846);
nand U11643 (N_11643,N_10707,N_11208);
nand U11644 (N_11644,N_10569,N_10966);
or U11645 (N_11645,N_10577,N_10349);
or U11646 (N_11646,N_10326,N_10224);
xnor U11647 (N_11647,N_10408,N_10596);
and U11648 (N_11648,N_11173,N_11002);
nor U11649 (N_11649,N_10465,N_10348);
xor U11650 (N_11650,N_11219,N_10847);
nand U11651 (N_11651,N_10283,N_10886);
nor U11652 (N_11652,N_10079,N_10513);
or U11653 (N_11653,N_10203,N_10287);
and U11654 (N_11654,N_10412,N_10133);
or U11655 (N_11655,N_10197,N_10084);
nand U11656 (N_11656,N_11102,N_10753);
xor U11657 (N_11657,N_10517,N_10483);
and U11658 (N_11658,N_10933,N_11181);
or U11659 (N_11659,N_10126,N_10848);
xor U11660 (N_11660,N_10965,N_10068);
nor U11661 (N_11661,N_10237,N_10449);
nor U11662 (N_11662,N_11172,N_10923);
nand U11663 (N_11663,N_11109,N_10487);
nand U11664 (N_11664,N_11062,N_11155);
nand U11665 (N_11665,N_10828,N_11065);
and U11666 (N_11666,N_10720,N_10254);
or U11667 (N_11667,N_11125,N_11176);
xnor U11668 (N_11668,N_10420,N_10856);
xor U11669 (N_11669,N_10378,N_10095);
nor U11670 (N_11670,N_11001,N_10837);
nand U11671 (N_11671,N_10199,N_10505);
nand U11672 (N_11672,N_10090,N_10066);
and U11673 (N_11673,N_10023,N_10708);
or U11674 (N_11674,N_10442,N_10801);
nor U11675 (N_11675,N_10822,N_10266);
or U11676 (N_11676,N_10212,N_10751);
nand U11677 (N_11677,N_10080,N_10046);
or U11678 (N_11678,N_10955,N_10231);
or U11679 (N_11679,N_11049,N_10997);
xnor U11680 (N_11680,N_10740,N_10008);
and U11681 (N_11681,N_10202,N_10620);
xor U11682 (N_11682,N_11093,N_11214);
or U11683 (N_11683,N_10443,N_11063);
or U11684 (N_11684,N_10444,N_10503);
nand U11685 (N_11685,N_10424,N_10909);
nand U11686 (N_11686,N_10419,N_10160);
nor U11687 (N_11687,N_10336,N_10364);
nor U11688 (N_11688,N_10072,N_11030);
nand U11689 (N_11689,N_11090,N_10048);
xnor U11690 (N_11690,N_10067,N_10809);
nor U11691 (N_11691,N_10782,N_10484);
nor U11692 (N_11692,N_10580,N_10622);
xor U11693 (N_11693,N_10635,N_10683);
xnor U11694 (N_11694,N_10600,N_11041);
xnor U11695 (N_11695,N_10137,N_10094);
nand U11696 (N_11696,N_10840,N_11164);
nand U11697 (N_11697,N_10081,N_10594);
or U11698 (N_11698,N_10636,N_10574);
or U11699 (N_11699,N_10520,N_10457);
and U11700 (N_11700,N_11064,N_10826);
nand U11701 (N_11701,N_11132,N_11188);
or U11702 (N_11702,N_10714,N_10088);
or U11703 (N_11703,N_10920,N_10152);
and U11704 (N_11704,N_10986,N_10022);
xor U11705 (N_11705,N_11171,N_11185);
nor U11706 (N_11706,N_10884,N_10796);
xor U11707 (N_11707,N_10978,N_10890);
and U11708 (N_11708,N_10340,N_11242);
or U11709 (N_11709,N_10351,N_11015);
or U11710 (N_11710,N_10603,N_10507);
or U11711 (N_11711,N_10724,N_10530);
xnor U11712 (N_11712,N_10165,N_10075);
nor U11713 (N_11713,N_10497,N_10876);
or U11714 (N_11714,N_10610,N_10980);
or U11715 (N_11715,N_10092,N_10727);
and U11716 (N_11716,N_10904,N_10360);
and U11717 (N_11717,N_10315,N_10721);
nor U11718 (N_11718,N_10618,N_11217);
and U11719 (N_11719,N_10833,N_10496);
xor U11720 (N_11720,N_10790,N_10147);
or U11721 (N_11721,N_10163,N_10854);
nand U11722 (N_11722,N_10971,N_11043);
nor U11723 (N_11723,N_11098,N_10944);
nand U11724 (N_11724,N_11221,N_10905);
xnor U11725 (N_11725,N_11121,N_10162);
or U11726 (N_11726,N_10195,N_11067);
nor U11727 (N_11727,N_10820,N_10469);
and U11728 (N_11728,N_10646,N_11003);
nor U11729 (N_11729,N_11230,N_10403);
xnor U11730 (N_11730,N_10003,N_10504);
xnor U11731 (N_11731,N_10500,N_11194);
or U11732 (N_11732,N_10201,N_10366);
and U11733 (N_11733,N_10332,N_10255);
nor U11734 (N_11734,N_10770,N_10252);
nand U11735 (N_11735,N_10353,N_10355);
xnor U11736 (N_11736,N_10735,N_11201);
xor U11737 (N_11737,N_10749,N_11133);
nand U11738 (N_11738,N_11200,N_10494);
nor U11739 (N_11739,N_11025,N_11014);
xnor U11740 (N_11740,N_10662,N_10999);
xnor U11741 (N_11741,N_10817,N_10438);
xor U11742 (N_11742,N_10745,N_11120);
nand U11743 (N_11743,N_11033,N_10785);
or U11744 (N_11744,N_11060,N_11205);
nor U11745 (N_11745,N_11182,N_11129);
nor U11746 (N_11746,N_10544,N_11066);
nand U11747 (N_11747,N_10428,N_11101);
nand U11748 (N_11748,N_10807,N_10110);
xnor U11749 (N_11749,N_10575,N_10021);
nor U11750 (N_11750,N_10467,N_10303);
nand U11751 (N_11751,N_10601,N_10693);
nor U11752 (N_11752,N_10987,N_10379);
and U11753 (N_11753,N_10471,N_11215);
nand U11754 (N_11754,N_10406,N_11183);
xnor U11755 (N_11755,N_10227,N_10737);
and U11756 (N_11756,N_10621,N_10324);
nor U11757 (N_11757,N_10281,N_10730);
and U11758 (N_11758,N_10793,N_10953);
and U11759 (N_11759,N_11005,N_10011);
nand U11760 (N_11760,N_10872,N_10061);
and U11761 (N_11761,N_10628,N_10957);
nor U11762 (N_11762,N_10167,N_10335);
nand U11763 (N_11763,N_10019,N_10633);
nor U11764 (N_11764,N_10526,N_10127);
nor U11765 (N_11765,N_10892,N_10711);
nand U11766 (N_11766,N_10159,N_10359);
or U11767 (N_11767,N_10998,N_11059);
nor U11768 (N_11768,N_10728,N_11122);
or U11769 (N_11769,N_11178,N_10376);
and U11770 (N_11770,N_10843,N_10089);
xnor U11771 (N_11771,N_11244,N_11011);
or U11772 (N_11772,N_10912,N_10690);
and U11773 (N_11773,N_11193,N_10960);
xor U11774 (N_11774,N_10650,N_10331);
or U11775 (N_11775,N_11126,N_10174);
xor U11776 (N_11776,N_10386,N_10391);
nand U11777 (N_11777,N_10521,N_11149);
xnor U11778 (N_11778,N_10915,N_11179);
and U11779 (N_11779,N_10883,N_10702);
xnor U11780 (N_11780,N_10136,N_10146);
nand U11781 (N_11781,N_10677,N_11052);
and U11782 (N_11782,N_11142,N_10664);
xor U11783 (N_11783,N_10009,N_10587);
nor U11784 (N_11784,N_10865,N_10418);
and U11785 (N_11785,N_10583,N_10911);
or U11786 (N_11786,N_11246,N_10161);
or U11787 (N_11787,N_10599,N_10821);
xor U11788 (N_11788,N_10210,N_10568);
or U11789 (N_11789,N_10680,N_10131);
nand U11790 (N_11790,N_10717,N_10123);
or U11791 (N_11791,N_10700,N_10881);
nand U11792 (N_11792,N_11137,N_10430);
nand U11793 (N_11793,N_11056,N_11019);
and U11794 (N_11794,N_10091,N_10389);
nor U11795 (N_11795,N_10539,N_11127);
or U11796 (N_11796,N_10297,N_10880);
nand U11797 (N_11797,N_10259,N_10954);
or U11798 (N_11798,N_10608,N_10799);
nand U11799 (N_11799,N_10374,N_10553);
nand U11800 (N_11800,N_10726,N_11022);
or U11801 (N_11801,N_10034,N_11218);
nor U11802 (N_11802,N_10506,N_10836);
xnor U11803 (N_11803,N_11168,N_10002);
xnor U11804 (N_11804,N_10271,N_10736);
or U11805 (N_11805,N_10653,N_10789);
nor U11806 (N_11806,N_10602,N_10936);
nor U11807 (N_11807,N_10399,N_10571);
xor U11808 (N_11808,N_10934,N_10716);
and U11809 (N_11809,N_10644,N_10783);
xnor U11810 (N_11810,N_10288,N_10555);
and U11811 (N_11811,N_10085,N_11158);
or U11812 (N_11812,N_10477,N_10925);
or U11813 (N_11813,N_10950,N_10916);
nand U11814 (N_11814,N_10579,N_11047);
nor U11815 (N_11815,N_11131,N_10400);
nand U11816 (N_11816,N_10054,N_10784);
and U11817 (N_11817,N_10972,N_11187);
and U11818 (N_11818,N_10029,N_10495);
nor U11819 (N_11819,N_11241,N_10523);
and U11820 (N_11820,N_10741,N_10806);
nand U11821 (N_11821,N_10615,N_10667);
xor U11822 (N_11822,N_10845,N_10250);
and U11823 (N_11823,N_10499,N_10042);
or U11824 (N_11824,N_11113,N_10226);
xor U11825 (N_11825,N_10632,N_10242);
nand U11826 (N_11826,N_11017,N_10447);
and U11827 (N_11827,N_10173,N_11116);
and U11828 (N_11828,N_10178,N_10398);
and U11829 (N_11829,N_11009,N_10516);
nor U11830 (N_11830,N_10888,N_10899);
xnor U11831 (N_11831,N_10742,N_10323);
nor U11832 (N_11832,N_10439,N_10025);
or U11833 (N_11833,N_11174,N_10069);
xnor U11834 (N_11834,N_10204,N_10764);
nor U11835 (N_11835,N_10104,N_10489);
or U11836 (N_11836,N_11204,N_10607);
or U11837 (N_11837,N_10356,N_10979);
nor U11838 (N_11838,N_10233,N_10681);
xor U11839 (N_11839,N_10831,N_10393);
and U11840 (N_11840,N_10651,N_10244);
nor U11841 (N_11841,N_10864,N_11071);
nor U11842 (N_11842,N_10339,N_10692);
or U11843 (N_11843,N_10264,N_11229);
xnor U11844 (N_11844,N_10219,N_10639);
nor U11845 (N_11845,N_10983,N_11156);
or U11846 (N_11846,N_10337,N_10962);
nand U11847 (N_11847,N_10511,N_10251);
nand U11848 (N_11848,N_10017,N_10289);
xnor U11849 (N_11849,N_10115,N_10018);
and U11850 (N_11850,N_10073,N_10597);
nor U11851 (N_11851,N_10445,N_10235);
and U11852 (N_11852,N_10786,N_10384);
xor U11853 (N_11853,N_10531,N_10668);
and U11854 (N_11854,N_10645,N_10401);
nor U11855 (N_11855,N_11233,N_10985);
nand U11856 (N_11856,N_10476,N_10542);
nand U11857 (N_11857,N_10958,N_10871);
nand U11858 (N_11858,N_10125,N_10877);
or U11859 (N_11859,N_10301,N_11107);
xor U11860 (N_11860,N_11247,N_10220);
xnor U11861 (N_11861,N_10723,N_11165);
nor U11862 (N_11862,N_11039,N_10032);
and U11863 (N_11863,N_11111,N_10642);
xor U11864 (N_11864,N_11010,N_11106);
nor U11865 (N_11865,N_10033,N_11036);
nor U11866 (N_11866,N_10238,N_11154);
nand U11867 (N_11867,N_10232,N_10150);
or U11868 (N_11868,N_10514,N_10239);
or U11869 (N_11869,N_10350,N_10451);
and U11870 (N_11870,N_10155,N_11249);
nand U11871 (N_11871,N_10765,N_10654);
xor U11872 (N_11872,N_10154,N_11078);
or U11873 (N_11873,N_10941,N_10550);
and U11874 (N_11874,N_10087,N_10879);
or U11875 (N_11875,N_10700,N_10131);
nand U11876 (N_11876,N_10311,N_11084);
nand U11877 (N_11877,N_10632,N_10286);
nor U11878 (N_11878,N_10577,N_10656);
and U11879 (N_11879,N_10066,N_10222);
xor U11880 (N_11880,N_10916,N_10297);
xor U11881 (N_11881,N_10280,N_10062);
nor U11882 (N_11882,N_10360,N_10442);
or U11883 (N_11883,N_11243,N_10112);
xnor U11884 (N_11884,N_10762,N_11227);
nor U11885 (N_11885,N_10615,N_11033);
or U11886 (N_11886,N_10647,N_10973);
or U11887 (N_11887,N_11115,N_10914);
xnor U11888 (N_11888,N_10482,N_10304);
and U11889 (N_11889,N_11202,N_10192);
xnor U11890 (N_11890,N_10331,N_10783);
or U11891 (N_11891,N_10811,N_10726);
or U11892 (N_11892,N_10205,N_10401);
xnor U11893 (N_11893,N_11240,N_10574);
nor U11894 (N_11894,N_10086,N_10369);
nor U11895 (N_11895,N_10334,N_11115);
and U11896 (N_11896,N_11145,N_10399);
nand U11897 (N_11897,N_10737,N_10516);
or U11898 (N_11898,N_10519,N_10126);
nand U11899 (N_11899,N_10802,N_11054);
nor U11900 (N_11900,N_11035,N_10040);
or U11901 (N_11901,N_10530,N_10844);
or U11902 (N_11902,N_10778,N_10700);
or U11903 (N_11903,N_10004,N_10884);
and U11904 (N_11904,N_11140,N_10807);
xnor U11905 (N_11905,N_10140,N_10119);
and U11906 (N_11906,N_11225,N_10626);
or U11907 (N_11907,N_10156,N_10768);
or U11908 (N_11908,N_10071,N_10408);
nand U11909 (N_11909,N_10201,N_10826);
or U11910 (N_11910,N_10596,N_10372);
and U11911 (N_11911,N_10541,N_11248);
and U11912 (N_11912,N_10193,N_10707);
xor U11913 (N_11913,N_10194,N_10648);
xnor U11914 (N_11914,N_10800,N_10920);
or U11915 (N_11915,N_10878,N_10306);
nor U11916 (N_11916,N_11060,N_11120);
or U11917 (N_11917,N_10496,N_11165);
or U11918 (N_11918,N_11034,N_10352);
nand U11919 (N_11919,N_10142,N_10839);
and U11920 (N_11920,N_10787,N_10324);
and U11921 (N_11921,N_10800,N_10542);
xor U11922 (N_11922,N_11167,N_10969);
or U11923 (N_11923,N_10395,N_11069);
and U11924 (N_11924,N_10698,N_10465);
xnor U11925 (N_11925,N_10759,N_10309);
and U11926 (N_11926,N_10785,N_10964);
nor U11927 (N_11927,N_10826,N_10620);
and U11928 (N_11928,N_10258,N_10224);
or U11929 (N_11929,N_10596,N_10103);
and U11930 (N_11930,N_10130,N_11108);
and U11931 (N_11931,N_11110,N_10846);
or U11932 (N_11932,N_11082,N_11114);
nor U11933 (N_11933,N_10294,N_10384);
nor U11934 (N_11934,N_10694,N_10355);
nor U11935 (N_11935,N_11134,N_11056);
or U11936 (N_11936,N_10278,N_10945);
nor U11937 (N_11937,N_10046,N_11041);
and U11938 (N_11938,N_10983,N_10149);
nand U11939 (N_11939,N_10142,N_10111);
xnor U11940 (N_11940,N_10617,N_10305);
xnor U11941 (N_11941,N_10587,N_11219);
nor U11942 (N_11942,N_10046,N_10332);
or U11943 (N_11943,N_10240,N_10483);
or U11944 (N_11944,N_10756,N_10694);
and U11945 (N_11945,N_10613,N_11010);
or U11946 (N_11946,N_11191,N_10082);
and U11947 (N_11947,N_10373,N_10204);
xnor U11948 (N_11948,N_10902,N_10650);
or U11949 (N_11949,N_10508,N_10789);
nand U11950 (N_11950,N_10017,N_10988);
xnor U11951 (N_11951,N_10395,N_11016);
or U11952 (N_11952,N_10106,N_10816);
nor U11953 (N_11953,N_10167,N_10285);
nand U11954 (N_11954,N_11072,N_11003);
nor U11955 (N_11955,N_10418,N_10741);
or U11956 (N_11956,N_11249,N_10070);
and U11957 (N_11957,N_11115,N_10466);
and U11958 (N_11958,N_10680,N_10876);
or U11959 (N_11959,N_10877,N_10298);
or U11960 (N_11960,N_10330,N_10014);
or U11961 (N_11961,N_11078,N_10283);
nand U11962 (N_11962,N_10430,N_11032);
xnor U11963 (N_11963,N_10713,N_10183);
or U11964 (N_11964,N_10371,N_10315);
and U11965 (N_11965,N_10332,N_10166);
or U11966 (N_11966,N_10322,N_10174);
or U11967 (N_11967,N_10239,N_10111);
or U11968 (N_11968,N_10143,N_10502);
xor U11969 (N_11969,N_11012,N_10460);
and U11970 (N_11970,N_10199,N_10846);
xor U11971 (N_11971,N_10993,N_10570);
or U11972 (N_11972,N_11249,N_10555);
nand U11973 (N_11973,N_10843,N_11233);
nand U11974 (N_11974,N_10129,N_10956);
nor U11975 (N_11975,N_10679,N_10571);
and U11976 (N_11976,N_10975,N_10923);
and U11977 (N_11977,N_10216,N_10653);
xnor U11978 (N_11978,N_11248,N_10874);
nor U11979 (N_11979,N_10503,N_10734);
nor U11980 (N_11980,N_10174,N_11231);
and U11981 (N_11981,N_10503,N_10477);
or U11982 (N_11982,N_11201,N_10288);
and U11983 (N_11983,N_10090,N_10481);
nor U11984 (N_11984,N_11226,N_11148);
or U11985 (N_11985,N_10353,N_10732);
and U11986 (N_11986,N_10296,N_10541);
nor U11987 (N_11987,N_10201,N_10327);
or U11988 (N_11988,N_11012,N_10699);
xor U11989 (N_11989,N_10674,N_10764);
or U11990 (N_11990,N_10601,N_10182);
or U11991 (N_11991,N_10417,N_11208);
nand U11992 (N_11992,N_11132,N_11161);
or U11993 (N_11993,N_10133,N_10011);
xor U11994 (N_11994,N_10195,N_10348);
and U11995 (N_11995,N_10027,N_10868);
or U11996 (N_11996,N_10868,N_10954);
nor U11997 (N_11997,N_10153,N_10508);
or U11998 (N_11998,N_10514,N_10535);
and U11999 (N_11999,N_10243,N_11005);
nor U12000 (N_12000,N_11181,N_10889);
nor U12001 (N_12001,N_11115,N_10884);
xor U12002 (N_12002,N_10451,N_10777);
nand U12003 (N_12003,N_11207,N_10344);
nand U12004 (N_12004,N_10653,N_10567);
or U12005 (N_12005,N_10297,N_11095);
nand U12006 (N_12006,N_11198,N_10894);
nor U12007 (N_12007,N_11165,N_10239);
nor U12008 (N_12008,N_10574,N_10854);
xnor U12009 (N_12009,N_10653,N_11153);
xor U12010 (N_12010,N_10537,N_10069);
nor U12011 (N_12011,N_10371,N_11206);
xnor U12012 (N_12012,N_10363,N_10355);
nand U12013 (N_12013,N_10343,N_10079);
and U12014 (N_12014,N_10259,N_10860);
and U12015 (N_12015,N_10346,N_11167);
and U12016 (N_12016,N_11178,N_10264);
and U12017 (N_12017,N_11058,N_10747);
nand U12018 (N_12018,N_10224,N_10320);
or U12019 (N_12019,N_10636,N_10807);
xor U12020 (N_12020,N_10091,N_10501);
nor U12021 (N_12021,N_10102,N_10404);
and U12022 (N_12022,N_10641,N_10819);
and U12023 (N_12023,N_10364,N_11147);
nor U12024 (N_12024,N_10656,N_10379);
nand U12025 (N_12025,N_11112,N_10589);
nand U12026 (N_12026,N_11228,N_10494);
and U12027 (N_12027,N_10593,N_10855);
xnor U12028 (N_12028,N_10249,N_10574);
and U12029 (N_12029,N_11032,N_11174);
xor U12030 (N_12030,N_10639,N_10709);
and U12031 (N_12031,N_10639,N_10233);
nor U12032 (N_12032,N_10896,N_10793);
xor U12033 (N_12033,N_10633,N_11135);
and U12034 (N_12034,N_10327,N_11014);
nand U12035 (N_12035,N_10159,N_10435);
and U12036 (N_12036,N_10889,N_10439);
and U12037 (N_12037,N_10033,N_10865);
or U12038 (N_12038,N_10497,N_11094);
nand U12039 (N_12039,N_10273,N_11140);
nand U12040 (N_12040,N_10624,N_10877);
and U12041 (N_12041,N_10054,N_10110);
nand U12042 (N_12042,N_10932,N_10194);
or U12043 (N_12043,N_10896,N_10126);
xnor U12044 (N_12044,N_10594,N_10916);
or U12045 (N_12045,N_11071,N_10629);
or U12046 (N_12046,N_11143,N_10569);
xnor U12047 (N_12047,N_10932,N_10789);
nand U12048 (N_12048,N_11202,N_10524);
nor U12049 (N_12049,N_11189,N_10060);
and U12050 (N_12050,N_10246,N_10783);
nor U12051 (N_12051,N_10418,N_10740);
xnor U12052 (N_12052,N_10270,N_10887);
nor U12053 (N_12053,N_10292,N_10145);
nand U12054 (N_12054,N_10921,N_10769);
or U12055 (N_12055,N_10798,N_11206);
and U12056 (N_12056,N_10847,N_10438);
and U12057 (N_12057,N_10144,N_10180);
xnor U12058 (N_12058,N_10638,N_11060);
or U12059 (N_12059,N_11070,N_10384);
nor U12060 (N_12060,N_11068,N_10505);
or U12061 (N_12061,N_10733,N_10210);
nor U12062 (N_12062,N_10466,N_10805);
nand U12063 (N_12063,N_10007,N_11103);
nand U12064 (N_12064,N_10018,N_10033);
nor U12065 (N_12065,N_10061,N_10588);
or U12066 (N_12066,N_10374,N_10728);
or U12067 (N_12067,N_10949,N_11189);
and U12068 (N_12068,N_10038,N_10810);
xor U12069 (N_12069,N_11028,N_10803);
or U12070 (N_12070,N_10523,N_10093);
and U12071 (N_12071,N_10789,N_10792);
nand U12072 (N_12072,N_11049,N_10537);
nor U12073 (N_12073,N_10065,N_10938);
or U12074 (N_12074,N_10095,N_10317);
nand U12075 (N_12075,N_10196,N_10045);
xor U12076 (N_12076,N_11131,N_10237);
or U12077 (N_12077,N_10199,N_10345);
xnor U12078 (N_12078,N_11171,N_10897);
and U12079 (N_12079,N_10172,N_10545);
or U12080 (N_12080,N_10739,N_10747);
and U12081 (N_12081,N_10614,N_10791);
nand U12082 (N_12082,N_11032,N_10950);
nand U12083 (N_12083,N_10385,N_10544);
and U12084 (N_12084,N_10521,N_10628);
or U12085 (N_12085,N_11181,N_10750);
xor U12086 (N_12086,N_10058,N_10540);
or U12087 (N_12087,N_10624,N_10161);
and U12088 (N_12088,N_11196,N_10289);
nand U12089 (N_12089,N_10550,N_10410);
or U12090 (N_12090,N_10198,N_10377);
xnor U12091 (N_12091,N_10693,N_10242);
xor U12092 (N_12092,N_11236,N_10976);
or U12093 (N_12093,N_10534,N_10559);
xor U12094 (N_12094,N_10944,N_10248);
and U12095 (N_12095,N_10296,N_10004);
or U12096 (N_12096,N_10141,N_10400);
and U12097 (N_12097,N_10667,N_10273);
nor U12098 (N_12098,N_10075,N_10998);
nand U12099 (N_12099,N_10518,N_10597);
nand U12100 (N_12100,N_10554,N_10733);
and U12101 (N_12101,N_10026,N_11226);
xor U12102 (N_12102,N_10079,N_10592);
nor U12103 (N_12103,N_10410,N_10231);
nand U12104 (N_12104,N_10012,N_10216);
or U12105 (N_12105,N_10072,N_10062);
nand U12106 (N_12106,N_10626,N_10094);
or U12107 (N_12107,N_10244,N_10904);
nor U12108 (N_12108,N_10273,N_10468);
nor U12109 (N_12109,N_10488,N_10479);
and U12110 (N_12110,N_10588,N_10338);
or U12111 (N_12111,N_10608,N_10446);
and U12112 (N_12112,N_11150,N_10851);
and U12113 (N_12113,N_10066,N_11128);
and U12114 (N_12114,N_10465,N_11151);
nand U12115 (N_12115,N_10596,N_11185);
nand U12116 (N_12116,N_10737,N_10721);
or U12117 (N_12117,N_10196,N_10305);
nand U12118 (N_12118,N_10992,N_10811);
nand U12119 (N_12119,N_10894,N_11234);
and U12120 (N_12120,N_10296,N_10323);
nand U12121 (N_12121,N_10523,N_10836);
or U12122 (N_12122,N_10049,N_10271);
nand U12123 (N_12123,N_10054,N_10463);
or U12124 (N_12124,N_10436,N_10879);
and U12125 (N_12125,N_10419,N_11104);
nor U12126 (N_12126,N_10343,N_10992);
or U12127 (N_12127,N_10130,N_10087);
nand U12128 (N_12128,N_10540,N_10599);
xnor U12129 (N_12129,N_10355,N_10584);
xnor U12130 (N_12130,N_10671,N_10148);
xnor U12131 (N_12131,N_10307,N_10234);
and U12132 (N_12132,N_10748,N_10867);
nor U12133 (N_12133,N_10345,N_10549);
and U12134 (N_12134,N_10559,N_10200);
nor U12135 (N_12135,N_10997,N_10460);
nand U12136 (N_12136,N_10300,N_11191);
or U12137 (N_12137,N_10183,N_10424);
or U12138 (N_12138,N_10095,N_10382);
xor U12139 (N_12139,N_10901,N_11225);
nand U12140 (N_12140,N_11018,N_10404);
nand U12141 (N_12141,N_11214,N_11219);
or U12142 (N_12142,N_10955,N_10265);
and U12143 (N_12143,N_10601,N_10927);
nand U12144 (N_12144,N_11004,N_10657);
nor U12145 (N_12145,N_11184,N_10568);
nor U12146 (N_12146,N_10961,N_11090);
xor U12147 (N_12147,N_10757,N_10035);
and U12148 (N_12148,N_10794,N_11220);
xor U12149 (N_12149,N_10226,N_10158);
nand U12150 (N_12150,N_10420,N_10303);
and U12151 (N_12151,N_10483,N_10352);
and U12152 (N_12152,N_10566,N_10911);
nand U12153 (N_12153,N_10745,N_11201);
or U12154 (N_12154,N_10374,N_10686);
xor U12155 (N_12155,N_10251,N_10909);
xnor U12156 (N_12156,N_10117,N_11041);
nand U12157 (N_12157,N_10500,N_10042);
and U12158 (N_12158,N_10860,N_10374);
or U12159 (N_12159,N_10232,N_10112);
nor U12160 (N_12160,N_10251,N_10721);
nor U12161 (N_12161,N_11199,N_10383);
nor U12162 (N_12162,N_11040,N_11094);
nand U12163 (N_12163,N_10944,N_10474);
or U12164 (N_12164,N_10957,N_10532);
nand U12165 (N_12165,N_10625,N_10804);
xor U12166 (N_12166,N_10230,N_11132);
xor U12167 (N_12167,N_10329,N_10169);
nor U12168 (N_12168,N_10114,N_10375);
xnor U12169 (N_12169,N_10745,N_10070);
xor U12170 (N_12170,N_11025,N_11058);
xnor U12171 (N_12171,N_10366,N_10069);
xnor U12172 (N_12172,N_10269,N_10273);
nand U12173 (N_12173,N_10885,N_10335);
nor U12174 (N_12174,N_10055,N_11033);
and U12175 (N_12175,N_10658,N_10850);
or U12176 (N_12176,N_11116,N_10717);
nor U12177 (N_12177,N_11139,N_10118);
and U12178 (N_12178,N_10659,N_10643);
and U12179 (N_12179,N_10259,N_10095);
or U12180 (N_12180,N_11028,N_10999);
or U12181 (N_12181,N_11088,N_10080);
and U12182 (N_12182,N_10396,N_10927);
or U12183 (N_12183,N_10418,N_10712);
nor U12184 (N_12184,N_10436,N_11167);
nand U12185 (N_12185,N_11170,N_10163);
xnor U12186 (N_12186,N_11004,N_10793);
or U12187 (N_12187,N_10772,N_10142);
xor U12188 (N_12188,N_10184,N_10335);
and U12189 (N_12189,N_11224,N_10916);
nand U12190 (N_12190,N_10210,N_10951);
xor U12191 (N_12191,N_11239,N_11140);
or U12192 (N_12192,N_10692,N_10554);
xor U12193 (N_12193,N_10051,N_10471);
xnor U12194 (N_12194,N_10377,N_11003);
and U12195 (N_12195,N_10610,N_10959);
nor U12196 (N_12196,N_10102,N_10912);
nand U12197 (N_12197,N_10725,N_10537);
xnor U12198 (N_12198,N_10651,N_10057);
xnor U12199 (N_12199,N_10269,N_10094);
xor U12200 (N_12200,N_11216,N_10341);
nand U12201 (N_12201,N_10466,N_10005);
or U12202 (N_12202,N_10005,N_10933);
xnor U12203 (N_12203,N_10543,N_10415);
or U12204 (N_12204,N_11119,N_11114);
xnor U12205 (N_12205,N_11189,N_10601);
and U12206 (N_12206,N_11119,N_10611);
xnor U12207 (N_12207,N_11209,N_10696);
and U12208 (N_12208,N_11229,N_10699);
and U12209 (N_12209,N_10410,N_11063);
nor U12210 (N_12210,N_10012,N_10372);
nand U12211 (N_12211,N_10220,N_10705);
or U12212 (N_12212,N_10922,N_10899);
xor U12213 (N_12213,N_10070,N_10873);
and U12214 (N_12214,N_10346,N_10858);
nand U12215 (N_12215,N_11070,N_10387);
or U12216 (N_12216,N_10811,N_10671);
or U12217 (N_12217,N_10937,N_10314);
xor U12218 (N_12218,N_10060,N_11219);
and U12219 (N_12219,N_10005,N_10017);
nand U12220 (N_12220,N_10730,N_10990);
nor U12221 (N_12221,N_10849,N_11086);
and U12222 (N_12222,N_10254,N_11023);
nand U12223 (N_12223,N_10637,N_11218);
or U12224 (N_12224,N_10496,N_10424);
nand U12225 (N_12225,N_10544,N_10732);
and U12226 (N_12226,N_10496,N_10590);
xnor U12227 (N_12227,N_10711,N_10976);
xor U12228 (N_12228,N_11043,N_10468);
nor U12229 (N_12229,N_11050,N_10680);
nor U12230 (N_12230,N_10873,N_10018);
or U12231 (N_12231,N_10593,N_10840);
nor U12232 (N_12232,N_11125,N_10940);
xor U12233 (N_12233,N_10218,N_10034);
xnor U12234 (N_12234,N_10410,N_10884);
or U12235 (N_12235,N_11004,N_10825);
or U12236 (N_12236,N_10719,N_11104);
and U12237 (N_12237,N_10896,N_10288);
and U12238 (N_12238,N_10589,N_10038);
or U12239 (N_12239,N_10199,N_11140);
nor U12240 (N_12240,N_10329,N_11086);
xnor U12241 (N_12241,N_10769,N_11044);
nor U12242 (N_12242,N_10570,N_10339);
or U12243 (N_12243,N_10002,N_11232);
xor U12244 (N_12244,N_10424,N_10599);
xnor U12245 (N_12245,N_11009,N_10245);
or U12246 (N_12246,N_10502,N_10519);
nand U12247 (N_12247,N_10606,N_10612);
nor U12248 (N_12248,N_10731,N_10683);
and U12249 (N_12249,N_11115,N_10856);
nand U12250 (N_12250,N_11241,N_10545);
or U12251 (N_12251,N_10545,N_10127);
nand U12252 (N_12252,N_11189,N_10427);
nand U12253 (N_12253,N_11248,N_10342);
xnor U12254 (N_12254,N_10911,N_10861);
or U12255 (N_12255,N_11019,N_10135);
nand U12256 (N_12256,N_10519,N_11030);
nor U12257 (N_12257,N_11072,N_10073);
nor U12258 (N_12258,N_11103,N_11159);
xor U12259 (N_12259,N_10465,N_10815);
xor U12260 (N_12260,N_10884,N_10769);
or U12261 (N_12261,N_10547,N_10777);
nor U12262 (N_12262,N_10811,N_10856);
and U12263 (N_12263,N_10423,N_10715);
xnor U12264 (N_12264,N_10688,N_10915);
or U12265 (N_12265,N_11132,N_10622);
nor U12266 (N_12266,N_11069,N_10827);
nor U12267 (N_12267,N_11204,N_10932);
or U12268 (N_12268,N_11228,N_10132);
xor U12269 (N_12269,N_10536,N_10621);
nand U12270 (N_12270,N_10797,N_10341);
nand U12271 (N_12271,N_10704,N_10527);
xor U12272 (N_12272,N_10522,N_10770);
nor U12273 (N_12273,N_10632,N_10333);
nor U12274 (N_12274,N_10476,N_10408);
xor U12275 (N_12275,N_10231,N_10743);
and U12276 (N_12276,N_10570,N_10289);
nor U12277 (N_12277,N_11081,N_10892);
nor U12278 (N_12278,N_10079,N_10358);
xor U12279 (N_12279,N_10825,N_11145);
and U12280 (N_12280,N_10478,N_11086);
and U12281 (N_12281,N_10674,N_11044);
nand U12282 (N_12282,N_11104,N_10771);
nand U12283 (N_12283,N_11032,N_11181);
nand U12284 (N_12284,N_10446,N_10917);
xnor U12285 (N_12285,N_10654,N_10730);
nor U12286 (N_12286,N_10710,N_10954);
or U12287 (N_12287,N_10890,N_10860);
or U12288 (N_12288,N_10137,N_11028);
xor U12289 (N_12289,N_10432,N_10778);
nor U12290 (N_12290,N_11089,N_10772);
nor U12291 (N_12291,N_10829,N_11214);
and U12292 (N_12292,N_11234,N_10954);
nor U12293 (N_12293,N_10865,N_10209);
nand U12294 (N_12294,N_10811,N_10812);
and U12295 (N_12295,N_10345,N_10736);
or U12296 (N_12296,N_10356,N_10971);
or U12297 (N_12297,N_10905,N_11117);
or U12298 (N_12298,N_10307,N_11143);
and U12299 (N_12299,N_10147,N_11172);
and U12300 (N_12300,N_11145,N_10445);
nand U12301 (N_12301,N_11174,N_10971);
nand U12302 (N_12302,N_10129,N_11174);
xnor U12303 (N_12303,N_10173,N_11189);
xor U12304 (N_12304,N_11092,N_10906);
or U12305 (N_12305,N_10288,N_10648);
nand U12306 (N_12306,N_10649,N_10555);
xor U12307 (N_12307,N_10171,N_10742);
nor U12308 (N_12308,N_10259,N_10572);
and U12309 (N_12309,N_10265,N_10481);
xnor U12310 (N_12310,N_10413,N_10611);
nor U12311 (N_12311,N_10358,N_11234);
xor U12312 (N_12312,N_10213,N_10843);
and U12313 (N_12313,N_10817,N_10233);
nor U12314 (N_12314,N_10746,N_10317);
and U12315 (N_12315,N_11074,N_10332);
nand U12316 (N_12316,N_10503,N_10781);
nand U12317 (N_12317,N_11200,N_10698);
nor U12318 (N_12318,N_10613,N_10132);
nand U12319 (N_12319,N_10318,N_10415);
nor U12320 (N_12320,N_11188,N_10335);
or U12321 (N_12321,N_10154,N_11013);
and U12322 (N_12322,N_11159,N_10349);
and U12323 (N_12323,N_10036,N_11038);
xor U12324 (N_12324,N_10178,N_10034);
nand U12325 (N_12325,N_10839,N_10162);
and U12326 (N_12326,N_10802,N_10664);
xnor U12327 (N_12327,N_10371,N_10482);
xnor U12328 (N_12328,N_10830,N_11064);
and U12329 (N_12329,N_10063,N_10632);
or U12330 (N_12330,N_10644,N_10607);
or U12331 (N_12331,N_11241,N_10453);
and U12332 (N_12332,N_10240,N_10561);
xor U12333 (N_12333,N_10762,N_10759);
or U12334 (N_12334,N_10206,N_10846);
nand U12335 (N_12335,N_10328,N_10941);
and U12336 (N_12336,N_11135,N_10006);
or U12337 (N_12337,N_10822,N_11138);
or U12338 (N_12338,N_10492,N_10415);
xor U12339 (N_12339,N_10428,N_10885);
or U12340 (N_12340,N_10355,N_10163);
and U12341 (N_12341,N_11197,N_10470);
or U12342 (N_12342,N_10067,N_10846);
nor U12343 (N_12343,N_10743,N_11231);
and U12344 (N_12344,N_10569,N_10394);
or U12345 (N_12345,N_11166,N_10280);
or U12346 (N_12346,N_11152,N_10431);
nor U12347 (N_12347,N_10357,N_10688);
or U12348 (N_12348,N_11022,N_11102);
nand U12349 (N_12349,N_10378,N_10479);
and U12350 (N_12350,N_10180,N_10190);
xnor U12351 (N_12351,N_10029,N_10182);
xor U12352 (N_12352,N_11190,N_10020);
nor U12353 (N_12353,N_11049,N_10384);
and U12354 (N_12354,N_10002,N_10314);
nor U12355 (N_12355,N_10442,N_10999);
nor U12356 (N_12356,N_11000,N_10442);
or U12357 (N_12357,N_11141,N_10849);
and U12358 (N_12358,N_10993,N_10789);
and U12359 (N_12359,N_11060,N_10828);
xnor U12360 (N_12360,N_10458,N_11156);
and U12361 (N_12361,N_10422,N_10199);
and U12362 (N_12362,N_10686,N_11161);
and U12363 (N_12363,N_10355,N_10216);
and U12364 (N_12364,N_10004,N_10767);
nor U12365 (N_12365,N_11200,N_10767);
or U12366 (N_12366,N_10491,N_11104);
nand U12367 (N_12367,N_10149,N_10639);
nor U12368 (N_12368,N_10490,N_11201);
xor U12369 (N_12369,N_10653,N_10695);
nand U12370 (N_12370,N_10633,N_10021);
xnor U12371 (N_12371,N_10370,N_10161);
or U12372 (N_12372,N_10104,N_11133);
xnor U12373 (N_12373,N_10361,N_10827);
nand U12374 (N_12374,N_10134,N_10489);
nor U12375 (N_12375,N_10971,N_10983);
or U12376 (N_12376,N_10621,N_11225);
nand U12377 (N_12377,N_10678,N_11077);
nor U12378 (N_12378,N_10510,N_11103);
xor U12379 (N_12379,N_10142,N_10181);
nand U12380 (N_12380,N_10673,N_10972);
or U12381 (N_12381,N_10729,N_11049);
and U12382 (N_12382,N_10383,N_10155);
and U12383 (N_12383,N_11063,N_10986);
nand U12384 (N_12384,N_10873,N_11001);
xor U12385 (N_12385,N_10610,N_10317);
nand U12386 (N_12386,N_10261,N_10126);
and U12387 (N_12387,N_10676,N_10321);
nor U12388 (N_12388,N_11100,N_10869);
xnor U12389 (N_12389,N_11058,N_10525);
and U12390 (N_12390,N_11060,N_10113);
xnor U12391 (N_12391,N_10960,N_11042);
nand U12392 (N_12392,N_10571,N_11151);
nand U12393 (N_12393,N_10944,N_10190);
and U12394 (N_12394,N_10959,N_10118);
and U12395 (N_12395,N_10398,N_11105);
nor U12396 (N_12396,N_10173,N_10072);
or U12397 (N_12397,N_11144,N_11062);
xnor U12398 (N_12398,N_10946,N_10965);
xnor U12399 (N_12399,N_10497,N_10400);
and U12400 (N_12400,N_10414,N_10436);
nor U12401 (N_12401,N_10180,N_11074);
nand U12402 (N_12402,N_10483,N_10953);
xnor U12403 (N_12403,N_11041,N_10570);
or U12404 (N_12404,N_11164,N_11243);
and U12405 (N_12405,N_10273,N_11091);
nand U12406 (N_12406,N_10069,N_10463);
xnor U12407 (N_12407,N_10306,N_10519);
and U12408 (N_12408,N_10213,N_10801);
and U12409 (N_12409,N_10842,N_10229);
or U12410 (N_12410,N_10029,N_10400);
or U12411 (N_12411,N_10645,N_11201);
nand U12412 (N_12412,N_11132,N_10424);
and U12413 (N_12413,N_10726,N_10490);
or U12414 (N_12414,N_10504,N_10879);
nor U12415 (N_12415,N_10465,N_10674);
xor U12416 (N_12416,N_10134,N_10784);
nand U12417 (N_12417,N_11063,N_10547);
nor U12418 (N_12418,N_10273,N_10980);
or U12419 (N_12419,N_11191,N_10509);
nor U12420 (N_12420,N_10593,N_11079);
and U12421 (N_12421,N_11195,N_10274);
nand U12422 (N_12422,N_10327,N_10813);
and U12423 (N_12423,N_10440,N_10418);
nor U12424 (N_12424,N_10353,N_11020);
nor U12425 (N_12425,N_11000,N_10297);
nor U12426 (N_12426,N_10470,N_10677);
xor U12427 (N_12427,N_10899,N_10548);
and U12428 (N_12428,N_10002,N_10715);
or U12429 (N_12429,N_10675,N_11017);
and U12430 (N_12430,N_11037,N_10115);
or U12431 (N_12431,N_10824,N_10621);
xnor U12432 (N_12432,N_10878,N_10137);
nor U12433 (N_12433,N_10848,N_10477);
or U12434 (N_12434,N_10457,N_10626);
nor U12435 (N_12435,N_10843,N_10098);
or U12436 (N_12436,N_10582,N_10393);
and U12437 (N_12437,N_10930,N_10412);
nand U12438 (N_12438,N_10725,N_10087);
xnor U12439 (N_12439,N_10987,N_11237);
nand U12440 (N_12440,N_10335,N_10491);
and U12441 (N_12441,N_10447,N_10767);
xor U12442 (N_12442,N_10255,N_10087);
nand U12443 (N_12443,N_10729,N_10678);
nor U12444 (N_12444,N_10533,N_10293);
nor U12445 (N_12445,N_10232,N_10159);
and U12446 (N_12446,N_10458,N_10317);
nor U12447 (N_12447,N_10204,N_11138);
xnor U12448 (N_12448,N_11072,N_11237);
nor U12449 (N_12449,N_10669,N_10183);
xnor U12450 (N_12450,N_10077,N_10497);
xor U12451 (N_12451,N_10345,N_10547);
xor U12452 (N_12452,N_10045,N_10756);
and U12453 (N_12453,N_10314,N_10867);
nand U12454 (N_12454,N_10291,N_11132);
or U12455 (N_12455,N_10048,N_10211);
and U12456 (N_12456,N_10304,N_10931);
and U12457 (N_12457,N_11184,N_10467);
nand U12458 (N_12458,N_11069,N_10210);
or U12459 (N_12459,N_10596,N_10154);
nor U12460 (N_12460,N_10690,N_11212);
and U12461 (N_12461,N_10903,N_10889);
nand U12462 (N_12462,N_10052,N_10036);
nand U12463 (N_12463,N_10382,N_11136);
xnor U12464 (N_12464,N_10758,N_10802);
nor U12465 (N_12465,N_10791,N_10446);
and U12466 (N_12466,N_10527,N_10327);
or U12467 (N_12467,N_11247,N_10093);
nand U12468 (N_12468,N_11154,N_10738);
nand U12469 (N_12469,N_10998,N_11145);
or U12470 (N_12470,N_10319,N_10982);
xnor U12471 (N_12471,N_11186,N_10345);
xnor U12472 (N_12472,N_10482,N_11131);
nor U12473 (N_12473,N_11031,N_10759);
and U12474 (N_12474,N_11183,N_10724);
and U12475 (N_12475,N_10314,N_10661);
and U12476 (N_12476,N_11217,N_11142);
and U12477 (N_12477,N_10757,N_10558);
nor U12478 (N_12478,N_10134,N_10023);
xor U12479 (N_12479,N_10884,N_10182);
nor U12480 (N_12480,N_10210,N_10630);
or U12481 (N_12481,N_10119,N_10292);
and U12482 (N_12482,N_10905,N_10664);
nand U12483 (N_12483,N_10173,N_11127);
or U12484 (N_12484,N_10203,N_10783);
and U12485 (N_12485,N_11024,N_10601);
nand U12486 (N_12486,N_10250,N_10268);
or U12487 (N_12487,N_10111,N_10062);
or U12488 (N_12488,N_10224,N_10026);
or U12489 (N_12489,N_10719,N_10191);
nand U12490 (N_12490,N_10642,N_11208);
xor U12491 (N_12491,N_10879,N_10874);
and U12492 (N_12492,N_10471,N_11044);
and U12493 (N_12493,N_10572,N_10788);
nand U12494 (N_12494,N_10655,N_11136);
or U12495 (N_12495,N_10775,N_10761);
xnor U12496 (N_12496,N_10423,N_10837);
or U12497 (N_12497,N_11074,N_10553);
nor U12498 (N_12498,N_11055,N_10576);
nand U12499 (N_12499,N_10140,N_11008);
nor U12500 (N_12500,N_12333,N_11358);
nand U12501 (N_12501,N_12390,N_11933);
and U12502 (N_12502,N_12007,N_11588);
and U12503 (N_12503,N_12376,N_12451);
nor U12504 (N_12504,N_11404,N_11342);
nand U12505 (N_12505,N_12171,N_11789);
nor U12506 (N_12506,N_11940,N_11313);
nand U12507 (N_12507,N_11997,N_11319);
nor U12508 (N_12508,N_12142,N_11350);
or U12509 (N_12509,N_11409,N_11993);
or U12510 (N_12510,N_12307,N_11939);
nor U12511 (N_12511,N_11912,N_12071);
xnor U12512 (N_12512,N_11649,N_12039);
nor U12513 (N_12513,N_12345,N_11639);
nand U12514 (N_12514,N_12306,N_11331);
nor U12515 (N_12515,N_11707,N_11802);
and U12516 (N_12516,N_12379,N_11426);
xor U12517 (N_12517,N_12153,N_12319);
and U12518 (N_12518,N_11434,N_11810);
nor U12519 (N_12519,N_12158,N_11349);
and U12520 (N_12520,N_11457,N_11296);
nand U12521 (N_12521,N_12320,N_11811);
nand U12522 (N_12522,N_11370,N_11935);
nand U12523 (N_12523,N_11446,N_12411);
or U12524 (N_12524,N_11376,N_12261);
nand U12525 (N_12525,N_11488,N_12363);
and U12526 (N_12526,N_12388,N_12354);
xor U12527 (N_12527,N_11579,N_11405);
nand U12528 (N_12528,N_11492,N_12485);
nand U12529 (N_12529,N_11936,N_11750);
nor U12530 (N_12530,N_12317,N_12035);
and U12531 (N_12531,N_11668,N_11968);
or U12532 (N_12532,N_11794,N_11969);
nor U12533 (N_12533,N_12003,N_12194);
and U12534 (N_12534,N_12160,N_12083);
nor U12535 (N_12535,N_12398,N_11980);
xor U12536 (N_12536,N_12298,N_12081);
nor U12537 (N_12537,N_11829,N_12286);
or U12538 (N_12538,N_11503,N_12095);
and U12539 (N_12539,N_11781,N_11410);
or U12540 (N_12540,N_12184,N_11419);
or U12541 (N_12541,N_11889,N_12339);
nand U12542 (N_12542,N_11506,N_12137);
or U12543 (N_12543,N_11608,N_11784);
or U12544 (N_12544,N_12330,N_11747);
xor U12545 (N_12545,N_11898,N_11334);
xor U12546 (N_12546,N_11398,N_11858);
nor U12547 (N_12547,N_11805,N_12212);
nand U12548 (N_12548,N_12167,N_12352);
nand U12549 (N_12549,N_11485,N_12334);
nor U12550 (N_12550,N_12116,N_11305);
xnor U12551 (N_12551,N_11850,N_11470);
nor U12552 (N_12552,N_12497,N_11388);
nand U12553 (N_12553,N_11763,N_12107);
xor U12554 (N_12554,N_11299,N_11537);
or U12555 (N_12555,N_11374,N_12271);
nand U12556 (N_12556,N_11830,N_11702);
xnor U12557 (N_12557,N_12449,N_11843);
nand U12558 (N_12558,N_11384,N_11880);
xor U12559 (N_12559,N_12047,N_11704);
or U12560 (N_12560,N_11658,N_12498);
nand U12561 (N_12561,N_12405,N_11516);
or U12562 (N_12562,N_12313,N_12227);
and U12563 (N_12563,N_11458,N_11844);
nor U12564 (N_12564,N_11859,N_12125);
xnor U12565 (N_12565,N_12268,N_11822);
and U12566 (N_12566,N_11631,N_12091);
and U12567 (N_12567,N_12481,N_11863);
nand U12568 (N_12568,N_11544,N_11486);
xnor U12569 (N_12569,N_12136,N_11460);
nor U12570 (N_12570,N_12359,N_11303);
xor U12571 (N_12571,N_12106,N_11766);
nor U12572 (N_12572,N_12471,N_12289);
xor U12573 (N_12573,N_12407,N_11720);
or U12574 (N_12574,N_11284,N_12311);
or U12575 (N_12575,N_12065,N_11380);
nand U12576 (N_12576,N_12474,N_11420);
nand U12577 (N_12577,N_11574,N_12084);
nand U12578 (N_12578,N_12037,N_12172);
nand U12579 (N_12579,N_11441,N_12001);
xor U12580 (N_12580,N_11394,N_11402);
xor U12581 (N_12581,N_11988,N_11686);
and U12582 (N_12582,N_12123,N_12438);
and U12583 (N_12583,N_12458,N_11857);
nor U12584 (N_12584,N_11254,N_11497);
or U12585 (N_12585,N_12143,N_12199);
xor U12586 (N_12586,N_12242,N_11634);
and U12587 (N_12587,N_12276,N_11317);
nand U12588 (N_12588,N_11575,N_11283);
xnor U12589 (N_12589,N_11530,N_11630);
nand U12590 (N_12590,N_12208,N_12312);
nand U12591 (N_12591,N_11941,N_12410);
nand U12592 (N_12592,N_11924,N_12214);
xnor U12593 (N_12593,N_11339,N_12254);
or U12594 (N_12594,N_11651,N_12145);
xor U12595 (N_12595,N_11392,N_12157);
nand U12596 (N_12596,N_11677,N_12032);
xor U12597 (N_12597,N_12338,N_11724);
nand U12598 (N_12598,N_11564,N_11834);
or U12599 (N_12599,N_12211,N_12428);
and U12600 (N_12600,N_11362,N_12206);
or U12601 (N_12601,N_11416,N_11333);
and U12602 (N_12602,N_12408,N_11694);
or U12603 (N_12603,N_11320,N_11555);
nor U12604 (N_12604,N_11761,N_12262);
nor U12605 (N_12605,N_12423,N_11562);
nor U12606 (N_12606,N_12302,N_11603);
nor U12607 (N_12607,N_11315,N_11351);
nor U12608 (N_12608,N_12465,N_11644);
xnor U12609 (N_12609,N_12100,N_12140);
nor U12610 (N_12610,N_11760,N_12183);
or U12611 (N_12611,N_12435,N_12228);
or U12612 (N_12612,N_11689,N_11353);
nand U12613 (N_12613,N_11893,N_12096);
xnor U12614 (N_12614,N_11583,N_11578);
nor U12615 (N_12615,N_12074,N_12285);
nand U12616 (N_12616,N_12490,N_11733);
nor U12617 (N_12617,N_11931,N_12443);
nand U12618 (N_12618,N_11674,N_12269);
or U12619 (N_12619,N_11451,N_11558);
nor U12620 (N_12620,N_11864,N_11919);
or U12621 (N_12621,N_11330,N_11846);
or U12622 (N_12622,N_12446,N_11874);
nand U12623 (N_12623,N_12279,N_11927);
nor U12624 (N_12624,N_12124,N_12392);
xor U12625 (N_12625,N_11517,N_11258);
and U12626 (N_12626,N_12274,N_11736);
and U12627 (N_12627,N_11838,N_11521);
nor U12628 (N_12628,N_12008,N_11982);
xnor U12629 (N_12629,N_12326,N_11401);
nand U12630 (N_12630,N_12168,N_11310);
xor U12631 (N_12631,N_11741,N_12174);
nand U12632 (N_12632,N_12480,N_11638);
and U12633 (N_12633,N_11918,N_11652);
or U12634 (N_12634,N_12150,N_11901);
and U12635 (N_12635,N_12267,N_12025);
nor U12636 (N_12636,N_11340,N_11383);
nand U12637 (N_12637,N_12432,N_12119);
xnor U12638 (N_12638,N_12078,N_12484);
and U12639 (N_12639,N_11526,N_12369);
xnor U12640 (N_12640,N_12063,N_11659);
nand U12641 (N_12641,N_12399,N_12133);
or U12642 (N_12642,N_12395,N_11915);
xnor U12643 (N_12643,N_11599,N_12004);
nand U12644 (N_12644,N_11951,N_12093);
nor U12645 (N_12645,N_11818,N_11567);
nand U12646 (N_12646,N_11954,N_11450);
nand U12647 (N_12647,N_11587,N_12053);
nand U12648 (N_12648,N_12135,N_12441);
nand U12649 (N_12649,N_11701,N_12290);
or U12650 (N_12650,N_12014,N_12353);
xor U12651 (N_12651,N_11633,N_11594);
and U12652 (N_12652,N_11336,N_12429);
nor U12653 (N_12653,N_12337,N_12452);
xnor U12654 (N_12654,N_12151,N_11788);
or U12655 (N_12655,N_12346,N_11713);
and U12656 (N_12656,N_11727,N_11831);
nor U12657 (N_12657,N_12023,N_12122);
xor U12658 (N_12658,N_11559,N_11718);
nor U12659 (N_12659,N_12495,N_11994);
nand U12660 (N_12660,N_11885,N_11253);
nor U12661 (N_12661,N_11892,N_12403);
nor U12662 (N_12662,N_12110,N_11545);
or U12663 (N_12663,N_11729,N_11297);
and U12664 (N_12664,N_11853,N_12420);
nor U12665 (N_12665,N_11617,N_12349);
nand U12666 (N_12666,N_12050,N_11602);
nor U12667 (N_12667,N_11697,N_11891);
xnor U12668 (N_12668,N_11953,N_11512);
nand U12669 (N_12669,N_11826,N_12204);
nand U12670 (N_12670,N_12041,N_12266);
xnor U12671 (N_12671,N_11740,N_12186);
or U12672 (N_12672,N_11318,N_12360);
xnor U12673 (N_12673,N_11683,N_11820);
nand U12674 (N_12674,N_11364,N_12460);
nor U12675 (N_12675,N_11779,N_11906);
xor U12676 (N_12676,N_11490,N_11515);
nor U12677 (N_12677,N_12464,N_12335);
xnor U12678 (N_12678,N_12163,N_11746);
and U12679 (N_12679,N_11828,N_11377);
nand U12680 (N_12680,N_11772,N_11817);
nor U12681 (N_12681,N_12139,N_12221);
xnor U12682 (N_12682,N_12182,N_11920);
nand U12683 (N_12683,N_11448,N_11700);
or U12684 (N_12684,N_11604,N_12389);
or U12685 (N_12685,N_11878,N_11730);
nand U12686 (N_12686,N_11796,N_11321);
nand U12687 (N_12687,N_11790,N_11580);
nand U12688 (N_12688,N_11967,N_11593);
nor U12689 (N_12689,N_11696,N_11698);
or U12690 (N_12690,N_11636,N_11705);
nand U12691 (N_12691,N_11501,N_12431);
nor U12692 (N_12692,N_12232,N_12016);
xor U12693 (N_12693,N_12404,N_11459);
xnor U12694 (N_12694,N_11447,N_11354);
or U12695 (N_12695,N_11807,N_11449);
xnor U12696 (N_12696,N_11412,N_11281);
nor U12697 (N_12697,N_12121,N_11871);
or U12698 (N_12698,N_12386,N_11987);
nand U12699 (N_12699,N_12223,N_11532);
or U12700 (N_12700,N_11431,N_12426);
or U12701 (N_12701,N_12219,N_12225);
xnor U12702 (N_12702,N_11533,N_11841);
xor U12703 (N_12703,N_11895,N_11302);
or U12704 (N_12704,N_12087,N_12365);
xnor U12705 (N_12705,N_11592,N_11679);
nand U12706 (N_12706,N_11365,N_11572);
xor U12707 (N_12707,N_11732,N_12134);
nor U12708 (N_12708,N_11263,N_11872);
or U12709 (N_12709,N_11801,N_12385);
nand U12710 (N_12710,N_12082,N_12409);
xnor U12711 (N_12711,N_11540,N_11637);
xnor U12712 (N_12712,N_11648,N_11922);
and U12713 (N_12713,N_11748,N_12327);
xor U12714 (N_12714,N_12419,N_11627);
and U12715 (N_12715,N_11287,N_12099);
and U12716 (N_12716,N_12246,N_11926);
and U12717 (N_12717,N_12475,N_11962);
and U12718 (N_12718,N_11643,N_11884);
nor U12719 (N_12719,N_11665,N_11780);
xor U12720 (N_12720,N_11433,N_11708);
nor U12721 (N_12721,N_11849,N_12056);
xnor U12722 (N_12722,N_12332,N_11681);
nor U12723 (N_12723,N_12299,N_11654);
nor U12724 (N_12724,N_12373,N_11466);
xnor U12725 (N_12725,N_12027,N_12038);
nand U12726 (N_12726,N_12367,N_11944);
and U12727 (N_12727,N_12115,N_12085);
and U12728 (N_12728,N_11456,N_12394);
nor U12729 (N_12729,N_12425,N_12259);
nand U12730 (N_12730,N_11723,N_11438);
nand U12731 (N_12731,N_11984,N_12051);
xnor U12732 (N_12732,N_11596,N_11851);
or U12733 (N_12733,N_12457,N_11355);
nand U12734 (N_12734,N_11605,N_12105);
nor U12735 (N_12735,N_11758,N_11989);
nor U12736 (N_12736,N_11856,N_11252);
nand U12737 (N_12737,N_11836,N_11972);
and U12738 (N_12738,N_12132,N_11271);
nand U12739 (N_12739,N_11749,N_11827);
xor U12740 (N_12740,N_11326,N_11908);
or U12741 (N_12741,N_11942,N_11514);
xnor U12742 (N_12742,N_11261,N_11928);
nor U12743 (N_12743,N_11511,N_12052);
xnor U12744 (N_12744,N_12434,N_12169);
or U12745 (N_12745,N_11929,N_11534);
xnor U12746 (N_12746,N_11671,N_11866);
and U12747 (N_12747,N_11563,N_11824);
nand U12748 (N_12748,N_11632,N_12479);
nor U12749 (N_12749,N_12287,N_11847);
xnor U12750 (N_12750,N_11304,N_12235);
or U12751 (N_12751,N_11484,N_11845);
and U12752 (N_12752,N_12483,N_12488);
and U12753 (N_12753,N_11372,N_11552);
nor U12754 (N_12754,N_12043,N_11755);
or U12755 (N_12755,N_12402,N_12278);
nand U12756 (N_12756,N_11257,N_11752);
or U12757 (N_12757,N_11472,N_11539);
and U12758 (N_12758,N_11549,N_12098);
xor U12759 (N_12759,N_12472,N_11565);
or U12760 (N_12760,N_12344,N_11369);
nor U12761 (N_12761,N_12155,N_12040);
and U12762 (N_12762,N_11877,N_12216);
and U12763 (N_12763,N_12297,N_11560);
or U12764 (N_12764,N_12120,N_11876);
xnor U12765 (N_12765,N_11273,N_12215);
xor U12766 (N_12766,N_11952,N_11546);
xor U12767 (N_12767,N_11797,N_11646);
nor U12768 (N_12768,N_12102,N_11306);
xor U12769 (N_12769,N_11421,N_11422);
and U12770 (N_12770,N_12048,N_11883);
and U12771 (N_12771,N_11992,N_12397);
and U12772 (N_12772,N_12197,N_11958);
and U12773 (N_12773,N_11622,N_11391);
and U12774 (N_12774,N_11991,N_11667);
nor U12775 (N_12775,N_11717,N_12138);
and U12776 (N_12776,N_11903,N_12476);
nor U12777 (N_12777,N_11480,N_12018);
nor U12778 (N_12778,N_11786,N_11468);
xnor U12779 (N_12779,N_11499,N_11453);
and U12780 (N_12780,N_11657,N_11452);
or U12781 (N_12781,N_12301,N_11629);
and U12782 (N_12782,N_11946,N_11739);
and U12783 (N_12783,N_12412,N_12079);
or U12784 (N_12784,N_12057,N_11323);
and U12785 (N_12785,N_11360,N_12076);
or U12786 (N_12786,N_11769,N_12196);
nand U12787 (N_12787,N_11692,N_11411);
nor U12788 (N_12788,N_12300,N_11782);
xor U12789 (N_12789,N_12034,N_12371);
nand U12790 (N_12790,N_11581,N_11478);
or U12791 (N_12791,N_12200,N_11494);
nor U12792 (N_12792,N_11616,N_12318);
and U12793 (N_12793,N_12439,N_12021);
or U12794 (N_12794,N_12413,N_12112);
nor U12795 (N_12795,N_11454,N_11791);
and U12796 (N_12796,N_11867,N_11439);
xor U12797 (N_12797,N_11428,N_11938);
xnor U12798 (N_12798,N_11571,N_12382);
nor U12799 (N_12799,N_11277,N_11329);
or U12800 (N_12800,N_11823,N_11710);
or U12801 (N_12801,N_12370,N_12396);
nor U12802 (N_12802,N_12226,N_11726);
nand U12803 (N_12803,N_11557,N_11798);
and U12804 (N_12804,N_12283,N_12209);
and U12805 (N_12805,N_11379,N_11314);
and U12806 (N_12806,N_11762,N_12170);
nor U12807 (N_12807,N_11868,N_11442);
xor U12808 (N_12808,N_12252,N_12070);
nand U12809 (N_12809,N_11647,N_11524);
and U12810 (N_12810,N_11819,N_11378);
xor U12811 (N_12811,N_11417,N_11645);
xnor U12812 (N_12812,N_11839,N_12064);
nor U12813 (N_12813,N_11731,N_11619);
nor U12814 (N_12814,N_11981,N_12230);
or U12815 (N_12815,N_11476,N_12418);
and U12816 (N_12816,N_11437,N_11860);
and U12817 (N_12817,N_12114,N_11553);
or U12818 (N_12818,N_11359,N_11338);
and U12819 (N_12819,N_11907,N_12291);
nor U12820 (N_12820,N_11301,N_11429);
and U12821 (N_12821,N_11275,N_11744);
nor U12822 (N_12822,N_12164,N_11900);
xor U12823 (N_12823,N_11424,N_11719);
nor U12824 (N_12824,N_12461,N_11745);
or U12825 (N_12825,N_12243,N_11289);
or U12826 (N_12826,N_11347,N_11662);
nor U12827 (N_12827,N_12055,N_11346);
and U12828 (N_12828,N_12308,N_12130);
nor U12829 (N_12829,N_11597,N_12336);
xor U12830 (N_12830,N_11923,N_11684);
xnor U12831 (N_12831,N_11861,N_12316);
and U12832 (N_12832,N_11474,N_11949);
and U12833 (N_12833,N_12203,N_12477);
nor U12834 (N_12834,N_11959,N_12128);
or U12835 (N_12835,N_11507,N_11787);
xnor U12836 (N_12836,N_12181,N_11806);
nor U12837 (N_12837,N_11777,N_11274);
or U12838 (N_12838,N_12455,N_11979);
xnor U12839 (N_12839,N_12068,N_11852);
or U12840 (N_12840,N_11664,N_11343);
xnor U12841 (N_12841,N_11937,N_11804);
or U12842 (N_12842,N_12383,N_11778);
and U12843 (N_12843,N_12077,N_11525);
xor U12844 (N_12844,N_11816,N_11276);
xor U12845 (N_12845,N_11496,N_12238);
xor U12846 (N_12846,N_12321,N_12207);
xor U12847 (N_12847,N_12378,N_11256);
nor U12848 (N_12848,N_11660,N_12011);
or U12849 (N_12849,N_12118,N_12478);
and U12850 (N_12850,N_11436,N_11479);
nand U12851 (N_12851,N_11482,N_11280);
xnor U12852 (N_12852,N_12453,N_11595);
or U12853 (N_12853,N_11842,N_11712);
and U12854 (N_12854,N_11635,N_12374);
xnor U12855 (N_12855,N_12280,N_11768);
xor U12856 (N_12856,N_12253,N_11875);
nor U12857 (N_12857,N_11309,N_12469);
nand U12858 (N_12858,N_12251,N_11332);
xor U12859 (N_12859,N_12424,N_11734);
nand U12860 (N_12860,N_12022,N_11785);
and U12861 (N_12861,N_11985,N_11978);
xor U12862 (N_12862,N_11570,N_11528);
nand U12863 (N_12863,N_11687,N_12444);
nor U12864 (N_12864,N_11945,N_12258);
and U12865 (N_12865,N_12141,N_11770);
nor U12866 (N_12866,N_12010,N_12342);
nand U12867 (N_12867,N_12176,N_11508);
nor U12868 (N_12868,N_11335,N_11523);
xnor U12869 (N_12869,N_12331,N_12146);
xnor U12870 (N_12870,N_11735,N_12159);
or U12871 (N_12871,N_11792,N_11676);
nor U12872 (N_12872,N_11835,N_12103);
and U12873 (N_12873,N_11754,N_12250);
nand U12874 (N_12874,N_12303,N_12218);
or U12875 (N_12875,N_12059,N_11345);
and U12876 (N_12876,N_12494,N_11609);
or U12877 (N_12877,N_12315,N_11624);
nand U12878 (N_12878,N_12012,N_11699);
nand U12879 (N_12879,N_11267,N_12355);
nand U12880 (N_12880,N_11475,N_11751);
and U12881 (N_12881,N_11688,N_11715);
nand U12882 (N_12882,N_12248,N_11585);
or U12883 (N_12883,N_12213,N_11990);
and U12884 (N_12884,N_12104,N_11491);
nand U12885 (N_12885,N_12234,N_12440);
xnor U12886 (N_12886,N_11373,N_11870);
nand U12887 (N_12887,N_11298,N_12245);
nor U12888 (N_12888,N_11661,N_12400);
or U12889 (N_12889,N_12005,N_12364);
nand U12890 (N_12890,N_11505,N_11809);
nor U12891 (N_12891,N_12073,N_12466);
xor U12892 (N_12892,N_12162,N_11904);
and U12893 (N_12893,N_12437,N_12387);
and U12894 (N_12894,N_11481,N_11278);
nand U12895 (N_12895,N_11998,N_11489);
xor U12896 (N_12896,N_12180,N_11666);
or U12897 (N_12897,N_12263,N_12422);
and U12898 (N_12898,N_12054,N_11932);
nand U12899 (N_12899,N_11408,N_12069);
xnor U12900 (N_12900,N_11894,N_11815);
or U12901 (N_12901,N_11757,N_11322);
and U12902 (N_12902,N_11327,N_11548);
nand U12903 (N_12903,N_11502,N_11921);
nor U12904 (N_12904,N_11890,N_12377);
or U12905 (N_12905,N_11612,N_12368);
nor U12906 (N_12906,N_11272,N_11620);
and U12907 (N_12907,N_12393,N_11328);
nand U12908 (N_12908,N_12058,N_11930);
or U12909 (N_12909,N_12433,N_11950);
nor U12910 (N_12910,N_11821,N_12066);
xor U12911 (N_12911,N_12357,N_12362);
nand U12912 (N_12912,N_11541,N_12482);
nor U12913 (N_12913,N_11282,N_12049);
xor U12914 (N_12914,N_11995,N_11837);
nand U12915 (N_12915,N_12080,N_11294);
nand U12916 (N_12916,N_12126,N_12414);
and U12917 (N_12917,N_12111,N_12361);
nand U12918 (N_12918,N_12177,N_11640);
xor U12919 (N_12919,N_12445,N_11312);
or U12920 (N_12920,N_12195,N_11799);
nand U12921 (N_12921,N_11293,N_11896);
or U12922 (N_12922,N_12129,N_12401);
nand U12923 (N_12923,N_12094,N_11576);
xor U12924 (N_12924,N_12487,N_12421);
nor U12925 (N_12925,N_12305,N_12217);
and U12926 (N_12926,N_11606,N_12173);
nand U12927 (N_12927,N_12036,N_12131);
or U12928 (N_12928,N_11825,N_11477);
nand U12929 (N_12929,N_12086,N_12323);
xor U12930 (N_12930,N_11387,N_12467);
nor U12931 (N_12931,N_12187,N_12447);
nor U12932 (N_12932,N_11414,N_11756);
and U12933 (N_12933,N_12281,N_12042);
or U12934 (N_12934,N_12454,N_12277);
and U12935 (N_12935,N_12324,N_11569);
nor U12936 (N_12936,N_12192,N_11464);
nand U12937 (N_12937,N_11610,N_12288);
nand U12938 (N_12938,N_12356,N_11415);
xnor U12939 (N_12939,N_12165,N_11543);
and U12940 (N_12940,N_12092,N_11531);
and U12941 (N_12941,N_11672,N_11965);
nor U12942 (N_12942,N_11406,N_11917);
and U12943 (N_12943,N_12044,N_11399);
nor U12944 (N_12944,N_11970,N_11996);
and U12945 (N_12945,N_11626,N_11607);
xnor U12946 (N_12946,N_11783,N_11693);
xnor U12947 (N_12947,N_11655,N_11400);
nand U12948 (N_12948,N_12375,N_12241);
nand U12949 (N_12949,N_11611,N_12006);
xnor U12950 (N_12950,N_12149,N_11483);
nor U12951 (N_12951,N_11773,N_11865);
and U12952 (N_12952,N_11325,N_11519);
or U12953 (N_12953,N_12075,N_11582);
or U12954 (N_12954,N_11879,N_12210);
nand U12955 (N_12955,N_11389,N_11255);
nand U12956 (N_12956,N_12470,N_12329);
and U12957 (N_12957,N_12109,N_11586);
nand U12958 (N_12958,N_11614,N_11737);
nor U12959 (N_12959,N_11547,N_12322);
xor U12960 (N_12960,N_12144,N_12060);
or U12961 (N_12961,N_11469,N_11909);
nand U12962 (N_12962,N_11250,N_12372);
xor U12963 (N_12963,N_11986,N_11800);
or U12964 (N_12964,N_12328,N_11337);
nand U12965 (N_12965,N_12416,N_12002);
or U12966 (N_12966,N_11598,N_11960);
or U12967 (N_12967,N_11957,N_11300);
or U12968 (N_12968,N_11445,N_11881);
xor U12969 (N_12969,N_11974,N_11682);
xor U12970 (N_12970,N_12030,N_12191);
xor U12971 (N_12971,N_12033,N_12061);
or U12972 (N_12972,N_11425,N_12152);
or U12973 (N_12973,N_11813,N_11396);
xnor U12974 (N_12974,N_12496,N_11561);
xnor U12975 (N_12975,N_12463,N_12000);
xor U12976 (N_12976,N_12296,N_11966);
nor U12977 (N_12977,N_11573,N_12282);
nor U12978 (N_12978,N_11887,N_12198);
nand U12979 (N_12979,N_11386,N_11440);
nand U12980 (N_12980,N_11691,N_11418);
or U12981 (N_12981,N_11971,N_11765);
and U12982 (N_12982,N_12240,N_11840);
nand U12983 (N_12983,N_11265,N_11706);
nor U12984 (N_12984,N_11324,N_11873);
nor U12985 (N_12985,N_11711,N_12249);
xor U12986 (N_12986,N_11613,N_12067);
xor U12987 (N_12987,N_11709,N_11520);
and U12988 (N_12988,N_12127,N_11366);
xor U12989 (N_12989,N_12450,N_11947);
nand U12990 (N_12990,N_11341,N_12247);
or U12991 (N_12991,N_11397,N_12117);
or U12992 (N_12992,N_11390,N_12202);
or U12993 (N_12993,N_11869,N_12045);
nor U12994 (N_12994,N_12350,N_12089);
nor U12995 (N_12995,N_12442,N_12156);
or U12996 (N_12996,N_12293,N_11291);
and U12997 (N_12997,N_11279,N_11721);
xor U12998 (N_12998,N_11642,N_11685);
and U12999 (N_12999,N_12265,N_11886);
or U13000 (N_13000,N_11356,N_11601);
nor U13001 (N_13001,N_11368,N_11382);
xnor U13002 (N_13002,N_11911,N_11621);
nor U13003 (N_13003,N_11882,N_12231);
nor U13004 (N_13004,N_11266,N_12189);
nor U13005 (N_13005,N_11509,N_11363);
nand U13006 (N_13006,N_11656,N_12244);
xnor U13007 (N_13007,N_11432,N_12270);
xor U13008 (N_13008,N_12220,N_12147);
or U13009 (N_13009,N_12491,N_12264);
xnor U13010 (N_13010,N_11500,N_12310);
and U13011 (N_13011,N_12351,N_11568);
xnor U13012 (N_13012,N_12314,N_12427);
nor U13013 (N_13013,N_11285,N_11529);
and U13014 (N_13014,N_11862,N_11535);
xnor U13015 (N_13015,N_11268,N_12459);
nand U13016 (N_13016,N_12304,N_11615);
nor U13017 (N_13017,N_11344,N_12154);
and U13018 (N_13018,N_12272,N_12233);
nand U13019 (N_13019,N_12161,N_12341);
and U13020 (N_13020,N_12489,N_11455);
and U13021 (N_13021,N_11977,N_11577);
nand U13022 (N_13022,N_11675,N_11943);
or U13023 (N_13023,N_12381,N_11375);
or U13024 (N_13024,N_11262,N_12229);
xor U13025 (N_13025,N_11975,N_11983);
and U13026 (N_13026,N_11286,N_12493);
nor U13027 (N_13027,N_11498,N_11403);
nor U13028 (N_13028,N_11307,N_11504);
xor U13029 (N_13029,N_11899,N_11738);
nand U13030 (N_13030,N_11650,N_11670);
or U13031 (N_13031,N_12256,N_11669);
xnor U13032 (N_13032,N_11916,N_11465);
or U13033 (N_13033,N_12222,N_12072);
xnor U13034 (N_13034,N_12294,N_12193);
xor U13035 (N_13035,N_11473,N_11308);
nor U13036 (N_13036,N_11803,N_11427);
nand U13037 (N_13037,N_11348,N_11510);
xor U13038 (N_13038,N_11352,N_11625);
nor U13039 (N_13039,N_12462,N_11753);
or U13040 (N_13040,N_12309,N_12101);
or U13041 (N_13041,N_11808,N_12430);
or U13042 (N_13042,N_11764,N_11269);
or U13043 (N_13043,N_11902,N_11848);
nand U13044 (N_13044,N_11260,N_12473);
and U13045 (N_13045,N_12468,N_12024);
nand U13046 (N_13046,N_11680,N_11367);
xor U13047 (N_13047,N_12179,N_11775);
xor U13048 (N_13048,N_11973,N_12236);
nand U13049 (N_13049,N_11742,N_11833);
xor U13050 (N_13050,N_12097,N_11393);
and U13051 (N_13051,N_11467,N_12325);
nor U13052 (N_13052,N_12448,N_11493);
nand U13053 (N_13053,N_11771,N_11759);
nor U13054 (N_13054,N_11423,N_11728);
xnor U13055 (N_13055,N_11897,N_11590);
nand U13056 (N_13056,N_12224,N_11538);
nor U13057 (N_13057,N_11443,N_11690);
nor U13058 (N_13058,N_11623,N_11407);
or U13059 (N_13059,N_11653,N_12273);
and U13060 (N_13060,N_11471,N_11513);
xor U13061 (N_13061,N_12380,N_12090);
or U13062 (N_13062,N_11495,N_12205);
xor U13063 (N_13063,N_11290,N_11381);
or U13064 (N_13064,N_12031,N_11311);
xor U13065 (N_13065,N_12201,N_11948);
nor U13066 (N_13066,N_11487,N_11295);
xor U13067 (N_13067,N_11812,N_11678);
xnor U13068 (N_13068,N_11855,N_11641);
or U13069 (N_13069,N_12358,N_11292);
nor U13070 (N_13070,N_12108,N_11554);
nand U13071 (N_13071,N_11955,N_11976);
nand U13072 (N_13072,N_11536,N_11551);
or U13073 (N_13073,N_11663,N_11910);
and U13074 (N_13074,N_11316,N_12486);
nand U13075 (N_13075,N_12029,N_12348);
nor U13076 (N_13076,N_11925,N_12347);
and U13077 (N_13077,N_11905,N_11430);
xor U13078 (N_13078,N_12088,N_11725);
and U13079 (N_13079,N_12384,N_11913);
or U13080 (N_13080,N_11793,N_12295);
xor U13081 (N_13081,N_12340,N_11385);
or U13082 (N_13082,N_12015,N_11357);
nor U13083 (N_13083,N_11703,N_11743);
and U13084 (N_13084,N_11964,N_12343);
and U13085 (N_13085,N_12013,N_11963);
nor U13086 (N_13086,N_12492,N_12026);
xnor U13087 (N_13087,N_12113,N_11444);
nor U13088 (N_13088,N_11264,N_12178);
xnor U13089 (N_13089,N_12260,N_12255);
nor U13090 (N_13090,N_11628,N_12239);
or U13091 (N_13091,N_11270,N_12366);
nand U13092 (N_13092,N_12436,N_11518);
nand U13093 (N_13093,N_12062,N_11888);
or U13094 (N_13094,N_11767,N_12284);
nor U13095 (N_13095,N_11251,N_11956);
nand U13096 (N_13096,N_11288,N_12406);
nor U13097 (N_13097,N_11600,N_11550);
xnor U13098 (N_13098,N_11361,N_12415);
nor U13099 (N_13099,N_11934,N_11591);
nand U13100 (N_13100,N_11832,N_11914);
and U13101 (N_13101,N_12188,N_11435);
nand U13102 (N_13102,N_11714,N_11814);
and U13103 (N_13103,N_12237,N_12185);
xor U13104 (N_13104,N_11259,N_11413);
xor U13105 (N_13105,N_11854,N_12009);
xnor U13106 (N_13106,N_11461,N_11776);
xor U13107 (N_13107,N_11542,N_12391);
xor U13108 (N_13108,N_11774,N_12020);
xnor U13109 (N_13109,N_12019,N_12275);
xnor U13110 (N_13110,N_11584,N_11522);
xnor U13111 (N_13111,N_12175,N_12148);
xnor U13112 (N_13112,N_11722,N_12017);
or U13113 (N_13113,N_11371,N_11618);
nand U13114 (N_13114,N_11695,N_11556);
or U13115 (N_13115,N_12190,N_11527);
nand U13116 (N_13116,N_12028,N_12292);
or U13117 (N_13117,N_12417,N_11589);
nor U13118 (N_13118,N_11961,N_11673);
and U13119 (N_13119,N_11462,N_12046);
or U13120 (N_13120,N_11463,N_11716);
xor U13121 (N_13121,N_12166,N_12257);
or U13122 (N_13122,N_11566,N_11999);
and U13123 (N_13123,N_11795,N_11395);
nand U13124 (N_13124,N_12456,N_12499);
or U13125 (N_13125,N_11510,N_11553);
nor U13126 (N_13126,N_11799,N_11280);
or U13127 (N_13127,N_11509,N_12226);
nand U13128 (N_13128,N_12230,N_11427);
nand U13129 (N_13129,N_12217,N_12442);
and U13130 (N_13130,N_11403,N_11623);
nand U13131 (N_13131,N_12450,N_11786);
or U13132 (N_13132,N_11268,N_12330);
xnor U13133 (N_13133,N_11798,N_11692);
nand U13134 (N_13134,N_11265,N_12231);
or U13135 (N_13135,N_11999,N_11293);
nand U13136 (N_13136,N_12357,N_11500);
xnor U13137 (N_13137,N_11693,N_12030);
xor U13138 (N_13138,N_11300,N_11913);
nor U13139 (N_13139,N_11746,N_12465);
nor U13140 (N_13140,N_11488,N_12331);
or U13141 (N_13141,N_11916,N_12200);
xor U13142 (N_13142,N_12415,N_12127);
xor U13143 (N_13143,N_11771,N_11301);
and U13144 (N_13144,N_11792,N_11317);
and U13145 (N_13145,N_12498,N_12235);
nor U13146 (N_13146,N_11377,N_12465);
xnor U13147 (N_13147,N_12311,N_11386);
nor U13148 (N_13148,N_12180,N_11746);
nand U13149 (N_13149,N_12316,N_11979);
or U13150 (N_13150,N_11900,N_12473);
nand U13151 (N_13151,N_11967,N_11789);
xor U13152 (N_13152,N_11317,N_11259);
or U13153 (N_13153,N_11505,N_11890);
nand U13154 (N_13154,N_11284,N_12458);
nor U13155 (N_13155,N_11867,N_12256);
or U13156 (N_13156,N_11829,N_12429);
xnor U13157 (N_13157,N_11726,N_12368);
and U13158 (N_13158,N_11811,N_11890);
xor U13159 (N_13159,N_11936,N_12165);
nor U13160 (N_13160,N_12040,N_11577);
nand U13161 (N_13161,N_11736,N_11322);
nand U13162 (N_13162,N_12120,N_12218);
nor U13163 (N_13163,N_11697,N_12406);
or U13164 (N_13164,N_11792,N_11966);
nand U13165 (N_13165,N_11539,N_12311);
and U13166 (N_13166,N_12074,N_11817);
or U13167 (N_13167,N_12495,N_11860);
and U13168 (N_13168,N_11786,N_11482);
or U13169 (N_13169,N_12485,N_12355);
nand U13170 (N_13170,N_11567,N_11506);
nand U13171 (N_13171,N_12270,N_11882);
nand U13172 (N_13172,N_11422,N_12309);
xor U13173 (N_13173,N_12303,N_12384);
and U13174 (N_13174,N_12437,N_12255);
xnor U13175 (N_13175,N_12409,N_12061);
nor U13176 (N_13176,N_12111,N_12057);
nor U13177 (N_13177,N_12262,N_11622);
nand U13178 (N_13178,N_11680,N_12270);
nor U13179 (N_13179,N_11736,N_11260);
and U13180 (N_13180,N_12037,N_12089);
nand U13181 (N_13181,N_11845,N_11477);
nor U13182 (N_13182,N_11610,N_11343);
nand U13183 (N_13183,N_11600,N_11903);
xnor U13184 (N_13184,N_12255,N_11278);
nor U13185 (N_13185,N_12224,N_12159);
or U13186 (N_13186,N_12146,N_11786);
nand U13187 (N_13187,N_12290,N_12106);
nand U13188 (N_13188,N_11825,N_11738);
or U13189 (N_13189,N_12137,N_12058);
xor U13190 (N_13190,N_12121,N_12438);
or U13191 (N_13191,N_11518,N_12213);
or U13192 (N_13192,N_11451,N_11867);
xor U13193 (N_13193,N_11390,N_11871);
or U13194 (N_13194,N_11434,N_12274);
and U13195 (N_13195,N_11512,N_11917);
nor U13196 (N_13196,N_11833,N_11474);
nor U13197 (N_13197,N_11563,N_12027);
xor U13198 (N_13198,N_11828,N_12182);
xor U13199 (N_13199,N_12218,N_11785);
xor U13200 (N_13200,N_11758,N_11984);
or U13201 (N_13201,N_12485,N_12401);
xor U13202 (N_13202,N_11544,N_12149);
or U13203 (N_13203,N_11985,N_11535);
xor U13204 (N_13204,N_11560,N_12143);
nand U13205 (N_13205,N_12085,N_12095);
nor U13206 (N_13206,N_11596,N_11976);
nand U13207 (N_13207,N_11834,N_12133);
nand U13208 (N_13208,N_12047,N_11478);
nand U13209 (N_13209,N_12089,N_12179);
xnor U13210 (N_13210,N_11826,N_12024);
nor U13211 (N_13211,N_12170,N_11806);
and U13212 (N_13212,N_12257,N_12365);
nand U13213 (N_13213,N_11989,N_11311);
nand U13214 (N_13214,N_12358,N_11258);
nand U13215 (N_13215,N_12191,N_12051);
or U13216 (N_13216,N_12149,N_11719);
nor U13217 (N_13217,N_11284,N_11657);
nand U13218 (N_13218,N_11659,N_11505);
nor U13219 (N_13219,N_12378,N_12020);
nand U13220 (N_13220,N_11783,N_11579);
or U13221 (N_13221,N_12429,N_11679);
or U13222 (N_13222,N_12350,N_11935);
nor U13223 (N_13223,N_12151,N_11823);
xnor U13224 (N_13224,N_12238,N_12173);
or U13225 (N_13225,N_12121,N_11610);
nor U13226 (N_13226,N_11974,N_12148);
nor U13227 (N_13227,N_11282,N_11299);
nand U13228 (N_13228,N_12297,N_12027);
xor U13229 (N_13229,N_12319,N_11280);
xnor U13230 (N_13230,N_11822,N_11580);
nand U13231 (N_13231,N_12005,N_11259);
or U13232 (N_13232,N_11286,N_11356);
or U13233 (N_13233,N_11584,N_12013);
nand U13234 (N_13234,N_11296,N_12245);
nor U13235 (N_13235,N_11435,N_12345);
nor U13236 (N_13236,N_11952,N_11461);
and U13237 (N_13237,N_12358,N_11695);
xnor U13238 (N_13238,N_11972,N_12056);
or U13239 (N_13239,N_12145,N_11668);
nand U13240 (N_13240,N_11812,N_12213);
nor U13241 (N_13241,N_12284,N_11994);
and U13242 (N_13242,N_11807,N_12412);
nor U13243 (N_13243,N_11496,N_11977);
or U13244 (N_13244,N_11587,N_11316);
nand U13245 (N_13245,N_11582,N_11934);
xor U13246 (N_13246,N_12215,N_12404);
xor U13247 (N_13247,N_11412,N_12163);
and U13248 (N_13248,N_12176,N_12128);
or U13249 (N_13249,N_11567,N_11480);
nor U13250 (N_13250,N_12323,N_12258);
nand U13251 (N_13251,N_11684,N_11937);
and U13252 (N_13252,N_12293,N_11366);
nor U13253 (N_13253,N_11468,N_12006);
or U13254 (N_13254,N_11354,N_11884);
or U13255 (N_13255,N_11876,N_11457);
and U13256 (N_13256,N_12016,N_11650);
and U13257 (N_13257,N_12151,N_12457);
nand U13258 (N_13258,N_11685,N_12203);
nor U13259 (N_13259,N_11353,N_11354);
xnor U13260 (N_13260,N_11258,N_11819);
nor U13261 (N_13261,N_11539,N_11694);
nand U13262 (N_13262,N_11279,N_11608);
or U13263 (N_13263,N_12090,N_11517);
nor U13264 (N_13264,N_11997,N_11984);
or U13265 (N_13265,N_12308,N_11342);
or U13266 (N_13266,N_12344,N_11561);
nor U13267 (N_13267,N_12387,N_11542);
or U13268 (N_13268,N_12215,N_12284);
and U13269 (N_13269,N_11515,N_12137);
nor U13270 (N_13270,N_11899,N_11772);
or U13271 (N_13271,N_11482,N_11683);
or U13272 (N_13272,N_11709,N_12033);
and U13273 (N_13273,N_11462,N_11536);
nor U13274 (N_13274,N_11894,N_12441);
or U13275 (N_13275,N_12466,N_12193);
and U13276 (N_13276,N_12359,N_11465);
nor U13277 (N_13277,N_11268,N_11675);
or U13278 (N_13278,N_12367,N_12005);
xor U13279 (N_13279,N_11777,N_12096);
nand U13280 (N_13280,N_11693,N_11838);
and U13281 (N_13281,N_11774,N_11615);
and U13282 (N_13282,N_11325,N_11290);
and U13283 (N_13283,N_11603,N_11951);
and U13284 (N_13284,N_11263,N_11687);
nand U13285 (N_13285,N_12377,N_11332);
or U13286 (N_13286,N_11885,N_11517);
nand U13287 (N_13287,N_11572,N_12362);
nand U13288 (N_13288,N_11436,N_12109);
xnor U13289 (N_13289,N_11446,N_12181);
xnor U13290 (N_13290,N_11611,N_12093);
nor U13291 (N_13291,N_12093,N_11468);
nor U13292 (N_13292,N_11540,N_11845);
and U13293 (N_13293,N_11871,N_12410);
and U13294 (N_13294,N_11406,N_11307);
and U13295 (N_13295,N_12456,N_12491);
nor U13296 (N_13296,N_11787,N_11743);
nand U13297 (N_13297,N_11407,N_11857);
or U13298 (N_13298,N_11693,N_12283);
or U13299 (N_13299,N_12004,N_11540);
xnor U13300 (N_13300,N_11861,N_11696);
nand U13301 (N_13301,N_11991,N_12495);
nand U13302 (N_13302,N_11633,N_11521);
nand U13303 (N_13303,N_11984,N_11746);
or U13304 (N_13304,N_11620,N_11825);
nand U13305 (N_13305,N_12236,N_11270);
xor U13306 (N_13306,N_11658,N_11631);
or U13307 (N_13307,N_11684,N_12170);
and U13308 (N_13308,N_12010,N_12070);
nor U13309 (N_13309,N_12329,N_12145);
nand U13310 (N_13310,N_12390,N_11767);
nor U13311 (N_13311,N_12160,N_11662);
nor U13312 (N_13312,N_11636,N_11434);
and U13313 (N_13313,N_11503,N_12398);
nor U13314 (N_13314,N_11325,N_12263);
xor U13315 (N_13315,N_11590,N_11428);
or U13316 (N_13316,N_11626,N_12018);
or U13317 (N_13317,N_11722,N_12076);
xnor U13318 (N_13318,N_12063,N_11738);
nand U13319 (N_13319,N_12336,N_11347);
nand U13320 (N_13320,N_11827,N_12228);
nand U13321 (N_13321,N_11287,N_11870);
nor U13322 (N_13322,N_11686,N_11596);
nand U13323 (N_13323,N_11797,N_11578);
nand U13324 (N_13324,N_11758,N_12081);
or U13325 (N_13325,N_11649,N_11795);
or U13326 (N_13326,N_11265,N_11931);
xor U13327 (N_13327,N_12358,N_11807);
nand U13328 (N_13328,N_11301,N_11633);
and U13329 (N_13329,N_11567,N_11908);
or U13330 (N_13330,N_12359,N_12347);
nand U13331 (N_13331,N_11922,N_11686);
and U13332 (N_13332,N_11971,N_11518);
xor U13333 (N_13333,N_11495,N_12473);
nor U13334 (N_13334,N_12068,N_11687);
or U13335 (N_13335,N_11275,N_11855);
nand U13336 (N_13336,N_11809,N_11890);
or U13337 (N_13337,N_12197,N_11415);
xor U13338 (N_13338,N_11265,N_12235);
xor U13339 (N_13339,N_11305,N_11256);
xor U13340 (N_13340,N_12146,N_11879);
xor U13341 (N_13341,N_11566,N_12445);
and U13342 (N_13342,N_11505,N_11896);
and U13343 (N_13343,N_11762,N_11465);
or U13344 (N_13344,N_11317,N_12299);
nand U13345 (N_13345,N_11301,N_11494);
nand U13346 (N_13346,N_12058,N_11585);
and U13347 (N_13347,N_12006,N_11445);
nand U13348 (N_13348,N_11302,N_12239);
xor U13349 (N_13349,N_12237,N_11302);
xnor U13350 (N_13350,N_11398,N_12065);
and U13351 (N_13351,N_11439,N_11487);
nor U13352 (N_13352,N_11281,N_12331);
and U13353 (N_13353,N_11551,N_11442);
and U13354 (N_13354,N_12451,N_11887);
nand U13355 (N_13355,N_12384,N_12116);
and U13356 (N_13356,N_11962,N_11399);
nand U13357 (N_13357,N_12148,N_12173);
or U13358 (N_13358,N_11615,N_12016);
xnor U13359 (N_13359,N_11786,N_12412);
xor U13360 (N_13360,N_12341,N_12024);
nand U13361 (N_13361,N_11925,N_11582);
or U13362 (N_13362,N_11901,N_12133);
and U13363 (N_13363,N_11902,N_11307);
xnor U13364 (N_13364,N_12012,N_11639);
and U13365 (N_13365,N_12382,N_11438);
nor U13366 (N_13366,N_11830,N_11304);
nand U13367 (N_13367,N_12283,N_11559);
nand U13368 (N_13368,N_12287,N_12121);
and U13369 (N_13369,N_12131,N_12066);
xor U13370 (N_13370,N_11567,N_12121);
and U13371 (N_13371,N_12288,N_11328);
nor U13372 (N_13372,N_12490,N_12042);
nor U13373 (N_13373,N_11927,N_11448);
nand U13374 (N_13374,N_11653,N_12093);
or U13375 (N_13375,N_12233,N_11683);
nor U13376 (N_13376,N_11575,N_12166);
and U13377 (N_13377,N_12269,N_11553);
nand U13378 (N_13378,N_11630,N_12270);
nor U13379 (N_13379,N_11292,N_12043);
xnor U13380 (N_13380,N_11817,N_11667);
or U13381 (N_13381,N_11432,N_11829);
xnor U13382 (N_13382,N_11470,N_11347);
nand U13383 (N_13383,N_11321,N_11718);
nand U13384 (N_13384,N_11948,N_11581);
nor U13385 (N_13385,N_12445,N_11314);
nand U13386 (N_13386,N_11271,N_11337);
nor U13387 (N_13387,N_11253,N_11995);
xor U13388 (N_13388,N_11660,N_11925);
xor U13389 (N_13389,N_12265,N_11930);
or U13390 (N_13390,N_12456,N_12024);
xnor U13391 (N_13391,N_11671,N_12482);
or U13392 (N_13392,N_11582,N_11878);
and U13393 (N_13393,N_11703,N_11837);
xor U13394 (N_13394,N_11768,N_12022);
and U13395 (N_13395,N_12447,N_11868);
nand U13396 (N_13396,N_11457,N_11473);
and U13397 (N_13397,N_12305,N_11910);
or U13398 (N_13398,N_12051,N_11367);
xor U13399 (N_13399,N_12140,N_11658);
or U13400 (N_13400,N_11910,N_12430);
or U13401 (N_13401,N_11625,N_11292);
or U13402 (N_13402,N_11570,N_11285);
nand U13403 (N_13403,N_12152,N_11891);
nand U13404 (N_13404,N_12131,N_12333);
and U13405 (N_13405,N_11252,N_12089);
xor U13406 (N_13406,N_12018,N_12189);
and U13407 (N_13407,N_11851,N_12467);
or U13408 (N_13408,N_12175,N_12117);
xor U13409 (N_13409,N_12385,N_12247);
nor U13410 (N_13410,N_11886,N_11817);
and U13411 (N_13411,N_11413,N_11377);
nor U13412 (N_13412,N_12362,N_12332);
and U13413 (N_13413,N_11255,N_12094);
or U13414 (N_13414,N_12201,N_12153);
and U13415 (N_13415,N_12317,N_11912);
xnor U13416 (N_13416,N_11963,N_12428);
nand U13417 (N_13417,N_11729,N_12424);
xor U13418 (N_13418,N_12207,N_11992);
xnor U13419 (N_13419,N_12142,N_12058);
xnor U13420 (N_13420,N_11701,N_11918);
nand U13421 (N_13421,N_11739,N_11431);
nor U13422 (N_13422,N_11647,N_11427);
nand U13423 (N_13423,N_11704,N_11919);
or U13424 (N_13424,N_11543,N_11289);
xor U13425 (N_13425,N_11605,N_11598);
and U13426 (N_13426,N_12230,N_11476);
nor U13427 (N_13427,N_11519,N_12401);
or U13428 (N_13428,N_11360,N_11625);
nor U13429 (N_13429,N_12273,N_11686);
xor U13430 (N_13430,N_12197,N_11999);
nand U13431 (N_13431,N_11548,N_12418);
nor U13432 (N_13432,N_11895,N_12261);
or U13433 (N_13433,N_12080,N_12146);
and U13434 (N_13434,N_12013,N_11848);
nor U13435 (N_13435,N_12125,N_11491);
and U13436 (N_13436,N_12241,N_11848);
and U13437 (N_13437,N_11332,N_11528);
nand U13438 (N_13438,N_11844,N_12302);
xnor U13439 (N_13439,N_11617,N_12065);
and U13440 (N_13440,N_12160,N_11509);
xnor U13441 (N_13441,N_12031,N_11921);
xor U13442 (N_13442,N_12075,N_12136);
nand U13443 (N_13443,N_12173,N_12473);
and U13444 (N_13444,N_11275,N_12115);
or U13445 (N_13445,N_12418,N_11919);
and U13446 (N_13446,N_11562,N_11967);
nand U13447 (N_13447,N_11699,N_11847);
nand U13448 (N_13448,N_12293,N_11315);
xnor U13449 (N_13449,N_11965,N_11298);
nor U13450 (N_13450,N_11618,N_11746);
and U13451 (N_13451,N_12105,N_11887);
or U13452 (N_13452,N_11459,N_12409);
nand U13453 (N_13453,N_11382,N_11912);
nand U13454 (N_13454,N_11727,N_12259);
nor U13455 (N_13455,N_11434,N_11723);
xnor U13456 (N_13456,N_11736,N_11378);
nand U13457 (N_13457,N_11290,N_11655);
and U13458 (N_13458,N_11641,N_11399);
xnor U13459 (N_13459,N_11724,N_12401);
nor U13460 (N_13460,N_11280,N_11736);
xnor U13461 (N_13461,N_12037,N_12055);
nand U13462 (N_13462,N_12487,N_12409);
and U13463 (N_13463,N_12456,N_11283);
nor U13464 (N_13464,N_12112,N_11295);
xor U13465 (N_13465,N_11811,N_11426);
or U13466 (N_13466,N_11768,N_11739);
nand U13467 (N_13467,N_12016,N_11634);
and U13468 (N_13468,N_11850,N_11836);
nor U13469 (N_13469,N_11308,N_11591);
nand U13470 (N_13470,N_11568,N_12303);
and U13471 (N_13471,N_11834,N_12194);
and U13472 (N_13472,N_11284,N_11473);
xor U13473 (N_13473,N_11540,N_12432);
and U13474 (N_13474,N_11528,N_11411);
xnor U13475 (N_13475,N_11943,N_12067);
or U13476 (N_13476,N_11643,N_12497);
or U13477 (N_13477,N_11959,N_12426);
or U13478 (N_13478,N_11568,N_12175);
and U13479 (N_13479,N_11342,N_11464);
and U13480 (N_13480,N_11356,N_11335);
and U13481 (N_13481,N_12248,N_12203);
nor U13482 (N_13482,N_11626,N_12284);
and U13483 (N_13483,N_12162,N_12193);
or U13484 (N_13484,N_12356,N_12004);
and U13485 (N_13485,N_12444,N_12112);
and U13486 (N_13486,N_11570,N_11376);
or U13487 (N_13487,N_11786,N_12096);
nand U13488 (N_13488,N_12490,N_11933);
xnor U13489 (N_13489,N_11583,N_11855);
nor U13490 (N_13490,N_12165,N_11468);
xor U13491 (N_13491,N_12139,N_11493);
nand U13492 (N_13492,N_12126,N_12252);
nor U13493 (N_13493,N_11963,N_11904);
xor U13494 (N_13494,N_11670,N_11343);
nor U13495 (N_13495,N_11463,N_11379);
or U13496 (N_13496,N_12193,N_11632);
xnor U13497 (N_13497,N_12155,N_11749);
nand U13498 (N_13498,N_12080,N_12179);
nor U13499 (N_13499,N_12463,N_11547);
nand U13500 (N_13500,N_12354,N_11553);
and U13501 (N_13501,N_11881,N_11266);
or U13502 (N_13502,N_12349,N_12240);
xnor U13503 (N_13503,N_11672,N_12466);
xor U13504 (N_13504,N_11787,N_12476);
xnor U13505 (N_13505,N_11302,N_11766);
xnor U13506 (N_13506,N_11950,N_11534);
xnor U13507 (N_13507,N_11897,N_11352);
xor U13508 (N_13508,N_12320,N_11606);
or U13509 (N_13509,N_11653,N_11454);
nand U13510 (N_13510,N_12139,N_11612);
and U13511 (N_13511,N_12406,N_11900);
nand U13512 (N_13512,N_12136,N_12214);
nor U13513 (N_13513,N_11968,N_11328);
nor U13514 (N_13514,N_12100,N_11598);
xor U13515 (N_13515,N_12013,N_12269);
nor U13516 (N_13516,N_12084,N_12074);
xnor U13517 (N_13517,N_11319,N_11613);
xnor U13518 (N_13518,N_12085,N_12070);
or U13519 (N_13519,N_11735,N_11918);
and U13520 (N_13520,N_11574,N_12485);
xor U13521 (N_13521,N_11374,N_11464);
xnor U13522 (N_13522,N_11253,N_12084);
or U13523 (N_13523,N_12361,N_11682);
or U13524 (N_13524,N_12268,N_12353);
and U13525 (N_13525,N_12479,N_11540);
and U13526 (N_13526,N_12217,N_11830);
nor U13527 (N_13527,N_12460,N_12432);
nor U13528 (N_13528,N_11546,N_11756);
nor U13529 (N_13529,N_12237,N_12423);
and U13530 (N_13530,N_11922,N_11940);
nor U13531 (N_13531,N_11922,N_11498);
or U13532 (N_13532,N_11470,N_12400);
nand U13533 (N_13533,N_11279,N_12099);
nor U13534 (N_13534,N_11390,N_11413);
xor U13535 (N_13535,N_12070,N_11693);
nand U13536 (N_13536,N_12329,N_12368);
nor U13537 (N_13537,N_12246,N_12196);
or U13538 (N_13538,N_12226,N_12367);
nand U13539 (N_13539,N_11623,N_11729);
and U13540 (N_13540,N_11951,N_11877);
and U13541 (N_13541,N_11262,N_11343);
or U13542 (N_13542,N_12488,N_11860);
nor U13543 (N_13543,N_12034,N_12460);
or U13544 (N_13544,N_11807,N_11487);
and U13545 (N_13545,N_12116,N_11354);
nand U13546 (N_13546,N_11442,N_11887);
nand U13547 (N_13547,N_11699,N_12097);
and U13548 (N_13548,N_11708,N_11874);
xnor U13549 (N_13549,N_11898,N_11329);
xnor U13550 (N_13550,N_11597,N_12210);
nand U13551 (N_13551,N_12146,N_12131);
nor U13552 (N_13552,N_12001,N_12189);
xnor U13553 (N_13553,N_11418,N_11400);
xor U13554 (N_13554,N_11606,N_12105);
nand U13555 (N_13555,N_11658,N_12130);
xnor U13556 (N_13556,N_11774,N_12325);
xor U13557 (N_13557,N_11587,N_11408);
nor U13558 (N_13558,N_12197,N_11639);
nor U13559 (N_13559,N_12022,N_11291);
nor U13560 (N_13560,N_11739,N_12238);
or U13561 (N_13561,N_11403,N_12050);
and U13562 (N_13562,N_11867,N_11790);
nand U13563 (N_13563,N_12052,N_11445);
and U13564 (N_13564,N_12479,N_11945);
nand U13565 (N_13565,N_12371,N_12122);
nor U13566 (N_13566,N_12306,N_12053);
xnor U13567 (N_13567,N_11839,N_11297);
nor U13568 (N_13568,N_12038,N_11418);
and U13569 (N_13569,N_11351,N_12067);
or U13570 (N_13570,N_11900,N_11539);
nand U13571 (N_13571,N_11697,N_12221);
nand U13572 (N_13572,N_11742,N_11871);
and U13573 (N_13573,N_12302,N_11551);
xnor U13574 (N_13574,N_11256,N_11649);
or U13575 (N_13575,N_12121,N_11994);
nand U13576 (N_13576,N_11602,N_11278);
nand U13577 (N_13577,N_12110,N_12273);
nor U13578 (N_13578,N_11570,N_12364);
and U13579 (N_13579,N_11421,N_11615);
or U13580 (N_13580,N_11346,N_11415);
xnor U13581 (N_13581,N_11769,N_12287);
nand U13582 (N_13582,N_11417,N_11506);
or U13583 (N_13583,N_11874,N_12433);
xor U13584 (N_13584,N_11308,N_12399);
or U13585 (N_13585,N_11534,N_11386);
and U13586 (N_13586,N_12024,N_11847);
xor U13587 (N_13587,N_11961,N_11474);
xor U13588 (N_13588,N_11270,N_12036);
or U13589 (N_13589,N_11965,N_11324);
xor U13590 (N_13590,N_11362,N_11803);
nor U13591 (N_13591,N_11397,N_11890);
or U13592 (N_13592,N_12409,N_12288);
xnor U13593 (N_13593,N_11460,N_12385);
and U13594 (N_13594,N_12275,N_12433);
or U13595 (N_13595,N_11746,N_11655);
nand U13596 (N_13596,N_11720,N_11266);
nor U13597 (N_13597,N_11737,N_11367);
nor U13598 (N_13598,N_11690,N_11644);
nor U13599 (N_13599,N_12224,N_11655);
and U13600 (N_13600,N_11925,N_11954);
nor U13601 (N_13601,N_12004,N_11668);
or U13602 (N_13602,N_11491,N_12154);
nor U13603 (N_13603,N_12293,N_12057);
or U13604 (N_13604,N_11260,N_11628);
nor U13605 (N_13605,N_12351,N_11468);
and U13606 (N_13606,N_12018,N_11994);
and U13607 (N_13607,N_11358,N_11823);
and U13608 (N_13608,N_12359,N_11348);
nor U13609 (N_13609,N_11919,N_12200);
nand U13610 (N_13610,N_11804,N_12180);
nand U13611 (N_13611,N_12162,N_11738);
and U13612 (N_13612,N_12196,N_12379);
nor U13613 (N_13613,N_12382,N_11616);
xor U13614 (N_13614,N_11799,N_11891);
or U13615 (N_13615,N_12289,N_12095);
nor U13616 (N_13616,N_11981,N_12223);
nand U13617 (N_13617,N_12068,N_11678);
nor U13618 (N_13618,N_11347,N_11864);
nand U13619 (N_13619,N_11407,N_12151);
xnor U13620 (N_13620,N_12453,N_11511);
xnor U13621 (N_13621,N_11899,N_12485);
xor U13622 (N_13622,N_12172,N_11401);
xnor U13623 (N_13623,N_11736,N_12325);
or U13624 (N_13624,N_11322,N_12206);
nand U13625 (N_13625,N_11314,N_11564);
or U13626 (N_13626,N_12250,N_11936);
and U13627 (N_13627,N_11811,N_11723);
and U13628 (N_13628,N_11983,N_12384);
nor U13629 (N_13629,N_12373,N_12132);
nand U13630 (N_13630,N_12331,N_12473);
nand U13631 (N_13631,N_11593,N_11649);
and U13632 (N_13632,N_11589,N_12353);
and U13633 (N_13633,N_11989,N_12117);
and U13634 (N_13634,N_12034,N_12025);
nand U13635 (N_13635,N_11728,N_12416);
nor U13636 (N_13636,N_12274,N_11517);
nor U13637 (N_13637,N_12347,N_12117);
xor U13638 (N_13638,N_11762,N_12156);
or U13639 (N_13639,N_12070,N_11726);
and U13640 (N_13640,N_11360,N_11861);
nor U13641 (N_13641,N_12194,N_11935);
nor U13642 (N_13642,N_12282,N_11831);
nand U13643 (N_13643,N_11528,N_12323);
nor U13644 (N_13644,N_12091,N_11252);
nor U13645 (N_13645,N_12209,N_11815);
xor U13646 (N_13646,N_12019,N_11812);
xor U13647 (N_13647,N_11305,N_11531);
and U13648 (N_13648,N_11864,N_11518);
or U13649 (N_13649,N_11740,N_12162);
xor U13650 (N_13650,N_11871,N_11639);
nor U13651 (N_13651,N_11311,N_11895);
and U13652 (N_13652,N_11321,N_12408);
xor U13653 (N_13653,N_12265,N_12232);
xor U13654 (N_13654,N_11736,N_11838);
nand U13655 (N_13655,N_11842,N_12462);
xor U13656 (N_13656,N_11580,N_12002);
xor U13657 (N_13657,N_12219,N_11709);
and U13658 (N_13658,N_11281,N_11661);
xor U13659 (N_13659,N_12366,N_12097);
nand U13660 (N_13660,N_11272,N_12034);
nor U13661 (N_13661,N_11957,N_12057);
nand U13662 (N_13662,N_12184,N_11559);
or U13663 (N_13663,N_11940,N_11733);
and U13664 (N_13664,N_12293,N_11402);
and U13665 (N_13665,N_11422,N_12151);
nand U13666 (N_13666,N_12292,N_11749);
nand U13667 (N_13667,N_11819,N_11506);
and U13668 (N_13668,N_11758,N_11764);
nor U13669 (N_13669,N_12327,N_11479);
xor U13670 (N_13670,N_11649,N_12433);
xnor U13671 (N_13671,N_12283,N_11938);
nor U13672 (N_13672,N_12492,N_12069);
or U13673 (N_13673,N_12296,N_11635);
or U13674 (N_13674,N_11919,N_11980);
or U13675 (N_13675,N_11487,N_12457);
nand U13676 (N_13676,N_11451,N_11963);
nor U13677 (N_13677,N_12272,N_12214);
xnor U13678 (N_13678,N_11778,N_11607);
nor U13679 (N_13679,N_11617,N_12482);
or U13680 (N_13680,N_11725,N_11403);
nand U13681 (N_13681,N_12276,N_11274);
nand U13682 (N_13682,N_11574,N_11929);
nand U13683 (N_13683,N_12286,N_11402);
xnor U13684 (N_13684,N_11392,N_11921);
nand U13685 (N_13685,N_11358,N_11674);
or U13686 (N_13686,N_12465,N_12008);
and U13687 (N_13687,N_12150,N_12169);
xnor U13688 (N_13688,N_12374,N_11250);
nand U13689 (N_13689,N_11955,N_11304);
nor U13690 (N_13690,N_12085,N_11557);
or U13691 (N_13691,N_11557,N_11765);
xnor U13692 (N_13692,N_12334,N_11439);
nand U13693 (N_13693,N_12295,N_11329);
nor U13694 (N_13694,N_11951,N_12382);
and U13695 (N_13695,N_12443,N_12107);
xnor U13696 (N_13696,N_11832,N_12449);
xor U13697 (N_13697,N_11803,N_11558);
nor U13698 (N_13698,N_11329,N_11841);
nor U13699 (N_13699,N_12379,N_11940);
nor U13700 (N_13700,N_11740,N_11971);
nor U13701 (N_13701,N_12306,N_12240);
nand U13702 (N_13702,N_12495,N_12369);
nand U13703 (N_13703,N_11859,N_12332);
nor U13704 (N_13704,N_11687,N_12102);
xnor U13705 (N_13705,N_11977,N_11460);
nand U13706 (N_13706,N_12189,N_11557);
nand U13707 (N_13707,N_12422,N_12448);
nor U13708 (N_13708,N_11550,N_12192);
and U13709 (N_13709,N_11572,N_12211);
or U13710 (N_13710,N_11374,N_11360);
and U13711 (N_13711,N_12083,N_11806);
nand U13712 (N_13712,N_12113,N_12119);
nand U13713 (N_13713,N_12390,N_11563);
xor U13714 (N_13714,N_12440,N_12384);
xor U13715 (N_13715,N_11641,N_11443);
xor U13716 (N_13716,N_11957,N_11749);
nor U13717 (N_13717,N_11586,N_11335);
nor U13718 (N_13718,N_11824,N_11999);
or U13719 (N_13719,N_12408,N_11441);
nor U13720 (N_13720,N_12027,N_12419);
xnor U13721 (N_13721,N_12352,N_12028);
and U13722 (N_13722,N_11757,N_11832);
xor U13723 (N_13723,N_12189,N_11989);
and U13724 (N_13724,N_11839,N_12415);
nand U13725 (N_13725,N_12446,N_11473);
nand U13726 (N_13726,N_11573,N_12260);
and U13727 (N_13727,N_11585,N_12481);
nor U13728 (N_13728,N_11595,N_12038);
nor U13729 (N_13729,N_12394,N_11947);
nor U13730 (N_13730,N_12076,N_11901);
nand U13731 (N_13731,N_11943,N_12331);
nand U13732 (N_13732,N_11947,N_12431);
xor U13733 (N_13733,N_11488,N_12497);
xnor U13734 (N_13734,N_11422,N_12347);
nand U13735 (N_13735,N_12336,N_11372);
and U13736 (N_13736,N_11949,N_11819);
and U13737 (N_13737,N_11677,N_12143);
nor U13738 (N_13738,N_11474,N_11946);
and U13739 (N_13739,N_11491,N_12445);
and U13740 (N_13740,N_12432,N_12148);
and U13741 (N_13741,N_11406,N_11780);
or U13742 (N_13742,N_12456,N_11660);
nor U13743 (N_13743,N_12154,N_12442);
xnor U13744 (N_13744,N_11920,N_11687);
nor U13745 (N_13745,N_11956,N_12369);
xnor U13746 (N_13746,N_11870,N_11400);
nor U13747 (N_13747,N_12198,N_11630);
or U13748 (N_13748,N_12237,N_11882);
xnor U13749 (N_13749,N_12458,N_11282);
nand U13750 (N_13750,N_13082,N_13208);
or U13751 (N_13751,N_12542,N_13196);
nor U13752 (N_13752,N_12688,N_13562);
or U13753 (N_13753,N_12922,N_12554);
nor U13754 (N_13754,N_12847,N_12608);
nor U13755 (N_13755,N_12728,N_12650);
or U13756 (N_13756,N_12888,N_12577);
nand U13757 (N_13757,N_13008,N_13539);
and U13758 (N_13758,N_13117,N_13192);
or U13759 (N_13759,N_13365,N_13722);
and U13760 (N_13760,N_12601,N_12759);
nor U13761 (N_13761,N_13526,N_12683);
nand U13762 (N_13762,N_13437,N_13364);
or U13763 (N_13763,N_12934,N_13337);
or U13764 (N_13764,N_12753,N_13018);
xor U13765 (N_13765,N_12588,N_12879);
xnor U13766 (N_13766,N_13669,N_13559);
and U13767 (N_13767,N_13657,N_13468);
xnor U13768 (N_13768,N_13300,N_12961);
nor U13769 (N_13769,N_13721,N_12782);
nor U13770 (N_13770,N_12779,N_12793);
xnor U13771 (N_13771,N_13376,N_13304);
or U13772 (N_13772,N_12526,N_13743);
xnor U13773 (N_13773,N_13504,N_13031);
nor U13774 (N_13774,N_13318,N_13396);
nand U13775 (N_13775,N_13435,N_12777);
nand U13776 (N_13776,N_13171,N_13591);
nand U13777 (N_13777,N_13628,N_13727);
nand U13778 (N_13778,N_12834,N_13507);
nand U13779 (N_13779,N_13642,N_12637);
nor U13780 (N_13780,N_12744,N_12614);
or U13781 (N_13781,N_13613,N_13546);
nand U13782 (N_13782,N_13204,N_12551);
or U13783 (N_13783,N_13086,N_13728);
nor U13784 (N_13784,N_12755,N_13427);
xor U13785 (N_13785,N_12991,N_12982);
or U13786 (N_13786,N_13747,N_13139);
nor U13787 (N_13787,N_12740,N_13395);
nor U13788 (N_13788,N_12868,N_13007);
nor U13789 (N_13789,N_12906,N_13338);
nand U13790 (N_13790,N_12886,N_13452);
nand U13791 (N_13791,N_13510,N_13239);
or U13792 (N_13792,N_12882,N_13401);
nor U13793 (N_13793,N_13462,N_12684);
nand U13794 (N_13794,N_13575,N_12701);
nand U13795 (N_13795,N_13113,N_13377);
and U13796 (N_13796,N_12833,N_13446);
and U13797 (N_13797,N_13548,N_13660);
and U13798 (N_13798,N_13379,N_13725);
xnor U13799 (N_13799,N_12792,N_13100);
nand U13800 (N_13800,N_12696,N_13381);
xnor U13801 (N_13801,N_13409,N_13420);
nand U13802 (N_13802,N_12939,N_12655);
or U13803 (N_13803,N_13339,N_13502);
and U13804 (N_13804,N_13220,N_13665);
and U13805 (N_13805,N_12843,N_13605);
nand U13806 (N_13806,N_13415,N_13658);
xor U13807 (N_13807,N_13612,N_12831);
nor U13808 (N_13808,N_13022,N_13463);
or U13809 (N_13809,N_12949,N_13101);
nor U13810 (N_13810,N_13630,N_12548);
and U13811 (N_13811,N_12691,N_13317);
nand U13812 (N_13812,N_13740,N_13623);
or U13813 (N_13813,N_13060,N_12837);
or U13814 (N_13814,N_12505,N_13719);
xnor U13815 (N_13815,N_12745,N_13584);
and U13816 (N_13816,N_12765,N_13104);
and U13817 (N_13817,N_12512,N_12803);
or U13818 (N_13818,N_12785,N_13049);
nand U13819 (N_13819,N_12662,N_12852);
nor U13820 (N_13820,N_13170,N_13729);
xor U13821 (N_13821,N_13640,N_13538);
nand U13822 (N_13822,N_12959,N_13635);
and U13823 (N_13823,N_13650,N_13044);
nor U13824 (N_13824,N_13443,N_13545);
xnor U13825 (N_13825,N_12929,N_12523);
nor U13826 (N_13826,N_12770,N_12794);
nor U13827 (N_13827,N_12648,N_13334);
nand U13828 (N_13828,N_12587,N_12907);
or U13829 (N_13829,N_13715,N_12724);
or U13830 (N_13830,N_12653,N_13255);
xnor U13831 (N_13831,N_12750,N_13058);
nor U13832 (N_13832,N_13013,N_12638);
nor U13833 (N_13833,N_13594,N_12507);
and U13834 (N_13834,N_12754,N_13470);
nor U13835 (N_13835,N_13258,N_13551);
xnor U13836 (N_13836,N_13614,N_13554);
nor U13837 (N_13837,N_12628,N_13251);
nand U13838 (N_13838,N_12621,N_13703);
nor U13839 (N_13839,N_12877,N_12585);
and U13840 (N_13840,N_13696,N_12965);
or U13841 (N_13841,N_13303,N_13151);
nand U13842 (N_13842,N_12594,N_13666);
nor U13843 (N_13843,N_13536,N_13676);
xnor U13844 (N_13844,N_12730,N_13212);
and U13845 (N_13845,N_12543,N_13424);
and U13846 (N_13846,N_13295,N_13585);
nor U13847 (N_13847,N_12589,N_13389);
and U13848 (N_13848,N_13601,N_12546);
nand U13849 (N_13849,N_13291,N_12593);
or U13850 (N_13850,N_13159,N_12578);
xnor U13851 (N_13851,N_12912,N_12511);
and U13852 (N_13852,N_12656,N_13603);
and U13853 (N_13853,N_13249,N_12856);
nor U13854 (N_13854,N_12702,N_12727);
and U13855 (N_13855,N_13678,N_12849);
and U13856 (N_13856,N_12689,N_12618);
and U13857 (N_13857,N_12780,N_13259);
xnor U13858 (N_13858,N_13579,N_13114);
or U13859 (N_13859,N_12705,N_12773);
nand U13860 (N_13860,N_13332,N_13039);
nor U13861 (N_13861,N_13272,N_13061);
nand U13862 (N_13862,N_12786,N_12956);
nand U13863 (N_13863,N_13157,N_12804);
nor U13864 (N_13864,N_12816,N_13439);
xor U13865 (N_13865,N_13260,N_13380);
nand U13866 (N_13866,N_12736,N_13501);
nor U13867 (N_13867,N_13353,N_13503);
and U13868 (N_13868,N_13116,N_13035);
nor U13869 (N_13869,N_13683,N_12903);
xor U13870 (N_13870,N_13425,N_13186);
nor U13871 (N_13871,N_12678,N_13610);
or U13872 (N_13872,N_13011,N_13213);
nand U13873 (N_13873,N_13019,N_12720);
nor U13874 (N_13874,N_13659,N_12969);
or U13875 (N_13875,N_12818,N_13229);
or U13876 (N_13876,N_13625,N_13277);
nor U13877 (N_13877,N_13471,N_13182);
nand U13878 (N_13878,N_13587,N_13433);
nor U13879 (N_13879,N_12930,N_12790);
nor U13880 (N_13880,N_12873,N_12642);
or U13881 (N_13881,N_13704,N_13549);
or U13882 (N_13882,N_13062,N_12682);
xor U13883 (N_13883,N_13412,N_13537);
nand U13884 (N_13884,N_13621,N_12996);
and U13885 (N_13885,N_12699,N_12590);
xnor U13886 (N_13886,N_13543,N_12742);
nor U13887 (N_13887,N_12845,N_12558);
nor U13888 (N_13888,N_13108,N_12559);
and U13889 (N_13889,N_13359,N_13455);
xnor U13890 (N_13890,N_13600,N_12685);
nand U13891 (N_13891,N_12784,N_13053);
nor U13892 (N_13892,N_13375,N_13201);
nor U13893 (N_13893,N_13476,N_13231);
nor U13894 (N_13894,N_13385,N_12998);
nand U13895 (N_13895,N_13024,N_13484);
nand U13896 (N_13896,N_12641,N_13202);
and U13897 (N_13897,N_12570,N_12992);
nand U13898 (N_13898,N_13467,N_12919);
xor U13899 (N_13899,N_13529,N_13520);
and U13900 (N_13900,N_12695,N_13081);
or U13901 (N_13901,N_13651,N_12566);
xor U13902 (N_13902,N_13234,N_13426);
or U13903 (N_13903,N_12899,N_12640);
and U13904 (N_13904,N_13112,N_12876);
and U13905 (N_13905,N_12550,N_12958);
nand U13906 (N_13906,N_12573,N_13006);
and U13907 (N_13907,N_13483,N_13228);
xnor U13908 (N_13908,N_13363,N_13709);
and U13909 (N_13909,N_13699,N_13497);
and U13910 (N_13910,N_13378,N_12801);
nand U13911 (N_13911,N_13616,N_13736);
xnor U13912 (N_13912,N_13327,N_12576);
and U13913 (N_13913,N_13662,N_12751);
nor U13914 (N_13914,N_12603,N_13005);
xor U13915 (N_13915,N_12997,N_13680);
nand U13916 (N_13916,N_13012,N_13315);
nor U13917 (N_13917,N_13142,N_12767);
nand U13918 (N_13918,N_12898,N_12883);
and U13919 (N_13919,N_13134,N_13017);
and U13920 (N_13920,N_13564,N_12710);
and U13921 (N_13921,N_13403,N_12606);
nor U13922 (N_13922,N_12987,N_12935);
nor U13923 (N_13923,N_13319,N_12737);
xnor U13924 (N_13924,N_13410,N_12781);
xnor U13925 (N_13925,N_13450,N_13451);
nor U13926 (N_13926,N_13029,N_12670);
and U13927 (N_13927,N_12824,N_12516);
and U13928 (N_13928,N_13098,N_13275);
and U13929 (N_13929,N_12936,N_13569);
nor U13930 (N_13930,N_13508,N_13485);
or U13931 (N_13931,N_13211,N_13674);
and U13932 (N_13932,N_13568,N_13595);
nand U13933 (N_13933,N_13348,N_13028);
or U13934 (N_13934,N_13178,N_12950);
nor U13935 (N_13935,N_12717,N_12651);
nand U13936 (N_13936,N_13193,N_12545);
or U13937 (N_13937,N_12968,N_12893);
or U13938 (N_13938,N_12675,N_13639);
and U13939 (N_13939,N_12908,N_13224);
xor U13940 (N_13940,N_12994,N_12537);
nand U13941 (N_13941,N_12680,N_13517);
nor U13942 (N_13942,N_12844,N_12605);
nor U13943 (N_13943,N_13237,N_12687);
nor U13944 (N_13944,N_13590,N_13391);
or U13945 (N_13945,N_13593,N_13701);
nor U13946 (N_13946,N_13219,N_13523);
xor U13947 (N_13947,N_13469,N_13631);
xor U13948 (N_13948,N_13074,N_12874);
nand U13949 (N_13949,N_13493,N_12851);
xor U13950 (N_13950,N_12889,N_13553);
nor U13951 (N_13951,N_13051,N_13447);
xor U13952 (N_13952,N_12774,N_13690);
or U13953 (N_13953,N_12762,N_12769);
and U13954 (N_13954,N_13405,N_12677);
xnor U13955 (N_13955,N_13698,N_13056);
nand U13956 (N_13956,N_13422,N_12798);
nor U13957 (N_13957,N_13694,N_13077);
and U13958 (N_13958,N_12993,N_12700);
xnor U13959 (N_13959,N_12574,N_13288);
nand U13960 (N_13960,N_13472,N_12890);
or U13961 (N_13961,N_12716,N_12839);
nand U13962 (N_13962,N_12787,N_13619);
or U13963 (N_13963,N_13495,N_13465);
xnor U13964 (N_13964,N_13294,N_13488);
nor U13965 (N_13965,N_13399,N_13563);
or U13966 (N_13966,N_12528,N_13132);
or U13967 (N_13967,N_13418,N_13388);
and U13968 (N_13968,N_13392,N_12826);
and U13969 (N_13969,N_13480,N_12832);
and U13970 (N_13970,N_12529,N_13482);
xor U13971 (N_13971,N_13583,N_13183);
nor U13972 (N_13972,N_12622,N_12825);
or U13973 (N_13973,N_12871,N_12829);
xor U13974 (N_13974,N_12714,N_12858);
and U13975 (N_13975,N_13199,N_13355);
nor U13976 (N_13976,N_13606,N_12966);
nor U13977 (N_13977,N_13148,N_13281);
nor U13978 (N_13978,N_12972,N_13205);
and U13979 (N_13979,N_13161,N_12807);
nor U13980 (N_13980,N_13276,N_13386);
nand U13981 (N_13981,N_12582,N_12715);
nor U13982 (N_13982,N_12501,N_13166);
or U13983 (N_13983,N_12812,N_12931);
nor U13984 (N_13984,N_12562,N_13298);
nor U13985 (N_13985,N_12796,N_12760);
nand U13986 (N_13986,N_12607,N_13033);
and U13987 (N_13987,N_12863,N_13009);
xnor U13988 (N_13988,N_12748,N_13442);
or U13989 (N_13989,N_12502,N_12722);
and U13990 (N_13990,N_13697,N_12821);
and U13991 (N_13991,N_13306,N_12942);
xnor U13992 (N_13992,N_12667,N_13528);
nor U13993 (N_13993,N_13322,N_13041);
nor U13994 (N_13994,N_13629,N_12560);
nor U13995 (N_13995,N_12517,N_12713);
nor U13996 (N_13996,N_13050,N_12575);
nand U13997 (N_13997,N_12527,N_13655);
or U13998 (N_13998,N_13215,N_12957);
nor U13999 (N_13999,N_13069,N_13498);
and U14000 (N_14000,N_12810,N_13030);
nor U14001 (N_14001,N_13607,N_13209);
nand U14002 (N_14002,N_13407,N_12703);
nor U14003 (N_14003,N_12897,N_12974);
nor U14004 (N_14004,N_13692,N_13416);
nor U14005 (N_14005,N_13287,N_13246);
nand U14006 (N_14006,N_12894,N_13441);
nand U14007 (N_14007,N_12733,N_12761);
or U14008 (N_14008,N_12827,N_13466);
xnor U14009 (N_14009,N_12654,N_13580);
nand U14010 (N_14010,N_12772,N_13571);
xor U14011 (N_14011,N_13748,N_12978);
nor U14012 (N_14012,N_13649,N_13084);
nor U14013 (N_14013,N_13194,N_12553);
or U14014 (N_14014,N_12565,N_13210);
and U14015 (N_14015,N_12521,N_12538);
nor U14016 (N_14016,N_13016,N_12623);
nand U14017 (N_14017,N_13064,N_13648);
xnor U14018 (N_14018,N_12625,N_12967);
and U14019 (N_14019,N_12896,N_13598);
nand U14020 (N_14020,N_12595,N_12884);
and U14021 (N_14021,N_12933,N_12869);
nor U14022 (N_14022,N_12955,N_13121);
xnor U14023 (N_14023,N_12531,N_13687);
nor U14024 (N_14024,N_13481,N_12980);
or U14025 (N_14025,N_13682,N_13373);
or U14026 (N_14026,N_13684,N_12694);
and U14027 (N_14027,N_13487,N_13341);
nor U14028 (N_14028,N_13043,N_12556);
xnor U14029 (N_14029,N_12747,N_13599);
nand U14030 (N_14030,N_13609,N_12658);
nand U14031 (N_14031,N_13506,N_13126);
nor U14032 (N_14032,N_13413,N_12630);
or U14033 (N_14033,N_12932,N_12711);
and U14034 (N_14034,N_13675,N_13459);
or U14035 (N_14035,N_12923,N_13511);
or U14036 (N_14036,N_13404,N_12510);
xnor U14037 (N_14037,N_13328,N_13262);
xor U14038 (N_14038,N_12811,N_12976);
and U14039 (N_14039,N_13478,N_13429);
nand U14040 (N_14040,N_12610,N_13066);
and U14041 (N_14041,N_13068,N_13269);
or U14042 (N_14042,N_13516,N_12563);
nand U14043 (N_14043,N_13394,N_13440);
and U14044 (N_14044,N_13744,N_12915);
and U14045 (N_14045,N_13641,N_13254);
nor U14046 (N_14046,N_13456,N_13225);
nor U14047 (N_14047,N_13707,N_13274);
nand U14048 (N_14048,N_13078,N_12739);
nand U14049 (N_14049,N_12666,N_13138);
xor U14050 (N_14050,N_13240,N_13241);
nor U14051 (N_14051,N_12515,N_12840);
or U14052 (N_14052,N_12660,N_13505);
xor U14053 (N_14053,N_13233,N_12676);
nor U14054 (N_14054,N_13522,N_12850);
nor U14055 (N_14055,N_13634,N_12539);
nand U14056 (N_14056,N_13279,N_12814);
and U14057 (N_14057,N_12731,N_13133);
nand U14058 (N_14058,N_12911,N_13573);
nor U14059 (N_14059,N_13103,N_13626);
or U14060 (N_14060,N_13344,N_13131);
nor U14061 (N_14061,N_13085,N_12661);
xnor U14062 (N_14062,N_13045,N_13489);
xnor U14063 (N_14063,N_13032,N_13280);
nor U14064 (N_14064,N_12709,N_13496);
or U14065 (N_14065,N_13163,N_12872);
nor U14066 (N_14066,N_13486,N_12624);
and U14067 (N_14067,N_12564,N_12602);
nand U14068 (N_14068,N_12615,N_13167);
nor U14069 (N_14069,N_12620,N_13118);
and U14070 (N_14070,N_12925,N_13737);
nor U14071 (N_14071,N_13530,N_13741);
and U14072 (N_14072,N_13685,N_13547);
nand U14073 (N_14073,N_12830,N_13397);
or U14074 (N_14074,N_13654,N_13611);
and U14075 (N_14075,N_13369,N_13408);
xnor U14076 (N_14076,N_13092,N_13661);
nand U14077 (N_14077,N_13638,N_13122);
and U14078 (N_14078,N_13187,N_13055);
or U14079 (N_14079,N_12860,N_13700);
xor U14080 (N_14080,N_13691,N_12776);
xnor U14081 (N_14081,N_12887,N_12920);
and U14082 (N_14082,N_12671,N_12892);
nor U14083 (N_14083,N_12500,N_13326);
and U14084 (N_14084,N_12504,N_13454);
and U14085 (N_14085,N_13127,N_13177);
and U14086 (N_14086,N_13176,N_13586);
xor U14087 (N_14087,N_13174,N_13689);
xnor U14088 (N_14088,N_12672,N_13109);
xor U14089 (N_14089,N_13330,N_13705);
nand U14090 (N_14090,N_13550,N_13312);
and U14091 (N_14091,N_13256,N_13561);
xor U14092 (N_14092,N_12509,N_13512);
nor U14093 (N_14093,N_13266,N_13110);
or U14094 (N_14094,N_12944,N_13336);
nor U14095 (N_14095,N_12584,N_13203);
or U14096 (N_14096,N_12766,N_13036);
xor U14097 (N_14097,N_13130,N_13500);
nor U14098 (N_14098,N_12609,N_13532);
or U14099 (N_14099,N_13738,N_12508);
and U14100 (N_14100,N_13710,N_13438);
nand U14101 (N_14101,N_12881,N_13627);
nand U14102 (N_14102,N_12657,N_13147);
nor U14103 (N_14103,N_13268,N_13604);
nand U14104 (N_14104,N_13168,N_12918);
or U14105 (N_14105,N_12617,N_13002);
nor U14106 (N_14106,N_13492,N_12698);
nand U14107 (N_14107,N_13038,N_13156);
and U14108 (N_14108,N_13316,N_12901);
nand U14109 (N_14109,N_13181,N_12557);
and U14110 (N_14110,N_12547,N_13023);
nand U14111 (N_14111,N_13042,N_12866);
xor U14112 (N_14112,N_13475,N_12693);
nor U14113 (N_14113,N_13226,N_12729);
or U14114 (N_14114,N_12647,N_13278);
and U14115 (N_14115,N_13608,N_13264);
or U14116 (N_14116,N_13681,N_12819);
xnor U14117 (N_14117,N_13457,N_13524);
nor U14118 (N_14118,N_13308,N_13449);
nand U14119 (N_14119,N_13667,N_13668);
nor U14120 (N_14120,N_13393,N_12988);
nor U14121 (N_14121,N_13025,N_12914);
or U14122 (N_14122,N_13672,N_12581);
nor U14123 (N_14123,N_13048,N_13301);
nand U14124 (N_14124,N_13188,N_13592);
and U14125 (N_14125,N_13102,N_13444);
and U14126 (N_14126,N_13216,N_13430);
nand U14127 (N_14127,N_13144,N_13253);
nand U14128 (N_14128,N_12846,N_13617);
nor U14129 (N_14129,N_12917,N_13180);
nand U14130 (N_14130,N_12743,N_13097);
xor U14131 (N_14131,N_12928,N_12686);
and U14132 (N_14132,N_12791,N_12536);
xor U14133 (N_14133,N_13146,N_12544);
and U14134 (N_14134,N_12970,N_12864);
and U14135 (N_14135,N_12916,N_13745);
and U14136 (N_14136,N_12948,N_12947);
nand U14137 (N_14137,N_13285,N_12971);
and U14138 (N_14138,N_12867,N_13702);
and U14139 (N_14139,N_12530,N_13556);
xnor U14140 (N_14140,N_13054,N_13671);
xor U14141 (N_14141,N_13140,N_12652);
nor U14142 (N_14142,N_12808,N_12945);
nand U14143 (N_14143,N_13749,N_12885);
and U14144 (N_14144,N_13540,N_13414);
nand U14145 (N_14145,N_13206,N_12937);
nand U14146 (N_14146,N_12636,N_12532);
or U14147 (N_14147,N_13434,N_13350);
nor U14148 (N_14148,N_12712,N_13010);
or U14149 (N_14149,N_13313,N_12809);
nor U14150 (N_14150,N_13622,N_13080);
xnor U14151 (N_14151,N_13340,N_13624);
xnor U14152 (N_14152,N_13431,N_12778);
nor U14153 (N_14153,N_13015,N_13534);
nor U14154 (N_14154,N_13347,N_13693);
and U14155 (N_14155,N_12855,N_12749);
and U14156 (N_14156,N_13521,N_12708);
and U14157 (N_14157,N_13565,N_13198);
or U14158 (N_14158,N_13479,N_12758);
or U14159 (N_14159,N_13165,N_13282);
and U14160 (N_14160,N_13004,N_13128);
and U14161 (N_14161,N_12659,N_12631);
nand U14162 (N_14162,N_12878,N_12668);
nor U14163 (N_14163,N_13515,N_12597);
xnor U14164 (N_14164,N_12592,N_13644);
or U14165 (N_14165,N_13227,N_13111);
nor U14166 (N_14166,N_12768,N_12552);
xor U14167 (N_14167,N_12951,N_12895);
xor U14168 (N_14168,N_13552,N_12665);
xnor U14169 (N_14169,N_13154,N_13230);
nand U14170 (N_14170,N_13739,N_13073);
nand U14171 (N_14171,N_13735,N_13297);
nand U14172 (N_14172,N_13162,N_13267);
nand U14173 (N_14173,N_13115,N_13250);
or U14174 (N_14174,N_12946,N_13021);
nand U14175 (N_14175,N_13284,N_12938);
or U14176 (N_14176,N_12817,N_12572);
or U14177 (N_14177,N_12891,N_13576);
or U14178 (N_14178,N_13656,N_13270);
and U14179 (N_14179,N_12561,N_13652);
nor U14180 (N_14180,N_12862,N_12836);
and U14181 (N_14181,N_13419,N_12627);
or U14182 (N_14182,N_13160,N_13372);
xnor U14183 (N_14183,N_13531,N_13519);
and U14184 (N_14184,N_12706,N_12822);
nor U14185 (N_14185,N_13717,N_12802);
xor U14186 (N_14186,N_13223,N_13514);
nor U14187 (N_14187,N_13075,N_13293);
nand U14188 (N_14188,N_12764,N_13083);
nand U14189 (N_14189,N_12952,N_13302);
and U14190 (N_14190,N_12789,N_13597);
and U14191 (N_14191,N_12823,N_13314);
nand U14192 (N_14192,N_12861,N_13362);
nor U14193 (N_14193,N_13620,N_13191);
or U14194 (N_14194,N_13345,N_13323);
nor U14195 (N_14195,N_12646,N_13020);
and U14196 (N_14196,N_13653,N_13141);
xnor U14197 (N_14197,N_13245,N_13686);
and U14198 (N_14198,N_13273,N_12815);
xor U14199 (N_14199,N_13136,N_13361);
nor U14200 (N_14200,N_13286,N_12841);
nor U14201 (N_14201,N_13324,N_13236);
xor U14202 (N_14202,N_13292,N_12799);
nor U14203 (N_14203,N_13718,N_13417);
nand U14204 (N_14204,N_13172,N_12735);
xnor U14205 (N_14205,N_12756,N_12611);
xor U14206 (N_14206,N_12813,N_13664);
or U14207 (N_14207,N_13555,N_12853);
nand U14208 (N_14208,N_13351,N_12697);
nor U14209 (N_14209,N_13093,N_13195);
xor U14210 (N_14210,N_12525,N_13207);
nand U14211 (N_14211,N_13222,N_13059);
and U14212 (N_14212,N_13733,N_12674);
nand U14213 (N_14213,N_12738,N_12979);
and U14214 (N_14214,N_13560,N_13290);
and U14215 (N_14215,N_12986,N_13706);
xnor U14216 (N_14216,N_13164,N_12503);
or U14217 (N_14217,N_13357,N_13732);
xor U14218 (N_14218,N_12604,N_13087);
and U14219 (N_14219,N_13535,N_12519);
xnor U14220 (N_14220,N_13106,N_13309);
and U14221 (N_14221,N_13052,N_13574);
nor U14222 (N_14222,N_13089,N_12612);
or U14223 (N_14223,N_12909,N_13076);
nor U14224 (N_14224,N_12619,N_13398);
or U14225 (N_14225,N_12984,N_12848);
and U14226 (N_14226,N_12783,N_12788);
nand U14227 (N_14227,N_13003,N_12643);
nor U14228 (N_14228,N_12513,N_13299);
or U14229 (N_14229,N_13063,N_13037);
nor U14230 (N_14230,N_12870,N_13411);
and U14231 (N_14231,N_13349,N_13129);
nor U14232 (N_14232,N_13421,N_12690);
and U14233 (N_14233,N_12805,N_12859);
xnor U14234 (N_14234,N_13238,N_13637);
and U14235 (N_14235,N_13001,N_12953);
xor U14236 (N_14236,N_13402,N_13310);
xnor U14237 (N_14237,N_12910,N_12632);
or U14238 (N_14238,N_12943,N_13368);
nor U14239 (N_14239,N_13383,N_13445);
nand U14240 (N_14240,N_13150,N_13366);
and U14241 (N_14241,N_13325,N_12596);
nand U14242 (N_14242,N_12989,N_12854);
or U14243 (N_14243,N_13184,N_13090);
or U14244 (N_14244,N_12977,N_13000);
and U14245 (N_14245,N_13577,N_13169);
nand U14246 (N_14246,N_13726,N_12567);
and U14247 (N_14247,N_12880,N_13602);
nor U14248 (N_14248,N_13329,N_13572);
xnor U14249 (N_14249,N_12990,N_13582);
and U14250 (N_14250,N_13567,N_13645);
nor U14251 (N_14251,N_13096,N_13248);
nand U14252 (N_14252,N_13541,N_12865);
xor U14253 (N_14253,N_13730,N_13716);
and U14254 (N_14254,N_13646,N_13153);
xor U14255 (N_14255,N_12940,N_13513);
or U14256 (N_14256,N_13305,N_12540);
nor U14257 (N_14257,N_12549,N_13509);
and U14258 (N_14258,N_12571,N_12900);
nor U14259 (N_14259,N_13647,N_13119);
nor U14260 (N_14260,N_12555,N_12579);
xnor U14261 (N_14261,N_12681,N_13588);
xnor U14262 (N_14262,N_13723,N_12635);
nor U14263 (N_14263,N_13244,N_12522);
nand U14264 (N_14264,N_13367,N_13217);
nand U14265 (N_14265,N_13643,N_13218);
nor U14266 (N_14266,N_12902,N_12857);
xor U14267 (N_14267,N_13200,N_13542);
xor U14268 (N_14268,N_13499,N_12664);
or U14269 (N_14269,N_12960,N_13734);
and U14270 (N_14270,N_13065,N_13027);
xor U14271 (N_14271,N_13670,N_13677);
xnor U14272 (N_14272,N_13034,N_13448);
or U14273 (N_14273,N_13589,N_12973);
nor U14274 (N_14274,N_13107,N_12999);
nor U14275 (N_14275,N_12704,N_13387);
xor U14276 (N_14276,N_13307,N_12626);
or U14277 (N_14277,N_13342,N_13221);
nand U14278 (N_14278,N_13143,N_13358);
and U14279 (N_14279,N_12975,N_13474);
and U14280 (N_14280,N_13453,N_13370);
nor U14281 (N_14281,N_12820,N_13354);
nand U14282 (N_14282,N_13428,N_13046);
and U14283 (N_14283,N_12725,N_12962);
nor U14284 (N_14284,N_13578,N_13158);
nand U14285 (N_14285,N_13558,N_13123);
nor U14286 (N_14286,N_12629,N_13711);
and U14287 (N_14287,N_12669,N_13633);
nor U14288 (N_14288,N_13175,N_12600);
xor U14289 (N_14289,N_12963,N_13040);
or U14290 (N_14290,N_12741,N_13321);
nor U14291 (N_14291,N_12533,N_13533);
nand U14292 (N_14292,N_12828,N_13712);
nand U14293 (N_14293,N_13557,N_13688);
and U14294 (N_14294,N_13283,N_13149);
xor U14295 (N_14295,N_13527,N_12541);
xor U14296 (N_14296,N_13371,N_12757);
xor U14297 (N_14297,N_13179,N_13615);
nor U14298 (N_14298,N_12634,N_13464);
and U14299 (N_14299,N_12726,N_13261);
nor U14300 (N_14300,N_13570,N_13461);
xnor U14301 (N_14301,N_12663,N_12927);
and U14302 (N_14302,N_13406,N_12795);
or U14303 (N_14303,N_12718,N_12520);
and U14304 (N_14304,N_13423,N_13458);
or U14305 (N_14305,N_13343,N_13400);
nor U14306 (N_14306,N_13360,N_12734);
or U14307 (N_14307,N_12613,N_13243);
xnor U14308 (N_14308,N_12645,N_13724);
xnor U14309 (N_14309,N_13331,N_13636);
and U14310 (N_14310,N_13746,N_12995);
xnor U14311 (N_14311,N_13374,N_12721);
nor U14312 (N_14312,N_13477,N_13026);
nor U14313 (N_14313,N_13296,N_13197);
and U14314 (N_14314,N_12586,N_12763);
and U14315 (N_14315,N_13190,N_13072);
xor U14316 (N_14316,N_13094,N_13095);
or U14317 (N_14317,N_13581,N_12842);
or U14318 (N_14318,N_13432,N_13695);
nor U14319 (N_14319,N_13352,N_12800);
xor U14320 (N_14320,N_12644,N_13679);
xor U14321 (N_14321,N_13596,N_12921);
or U14322 (N_14322,N_12524,N_13252);
xnor U14323 (N_14323,N_13105,N_13632);
xnor U14324 (N_14324,N_12580,N_13333);
nor U14325 (N_14325,N_13014,N_12633);
or U14326 (N_14326,N_13460,N_12913);
xnor U14327 (N_14327,N_12506,N_13120);
nand U14328 (N_14328,N_13491,N_12616);
xnor U14329 (N_14329,N_13289,N_13566);
or U14330 (N_14330,N_12924,N_12964);
or U14331 (N_14331,N_12835,N_12983);
and U14332 (N_14332,N_13091,N_13271);
or U14333 (N_14333,N_12583,N_12639);
xor U14334 (N_14334,N_13346,N_13124);
nand U14335 (N_14335,N_13708,N_13382);
nor U14336 (N_14336,N_12692,N_13214);
and U14337 (N_14337,N_13257,N_12838);
xnor U14338 (N_14338,N_13071,N_12797);
nor U14339 (N_14339,N_13320,N_13079);
xnor U14340 (N_14340,N_12904,N_13125);
or U14341 (N_14341,N_12875,N_13335);
nor U14342 (N_14342,N_13185,N_12568);
nand U14343 (N_14343,N_12707,N_13525);
nand U14344 (N_14344,N_13618,N_13518);
and U14345 (N_14345,N_13070,N_13742);
and U14346 (N_14346,N_13173,N_13384);
or U14347 (N_14347,N_12534,N_12535);
and U14348 (N_14348,N_13494,N_13242);
and U14349 (N_14349,N_13673,N_12926);
nor U14350 (N_14350,N_13311,N_12752);
nand U14351 (N_14351,N_12649,N_13247);
and U14352 (N_14352,N_12746,N_12591);
xor U14353 (N_14353,N_12518,N_12905);
and U14354 (N_14354,N_12598,N_13137);
nand U14355 (N_14355,N_13436,N_12775);
and U14356 (N_14356,N_13731,N_13235);
nor U14357 (N_14357,N_12806,N_13490);
xnor U14358 (N_14358,N_12679,N_12673);
nor U14359 (N_14359,N_13544,N_13714);
or U14360 (N_14360,N_13720,N_12771);
nand U14361 (N_14361,N_13713,N_13145);
nand U14362 (N_14362,N_13663,N_13099);
nand U14363 (N_14363,N_13135,N_13356);
or U14364 (N_14364,N_12569,N_12723);
nand U14365 (N_14365,N_12981,N_12985);
and U14366 (N_14366,N_12514,N_12719);
or U14367 (N_14367,N_12954,N_13189);
or U14368 (N_14368,N_13390,N_12732);
nor U14369 (N_14369,N_13152,N_13155);
nor U14370 (N_14370,N_13473,N_12941);
nand U14371 (N_14371,N_13057,N_13088);
nand U14372 (N_14372,N_13263,N_13067);
xnor U14373 (N_14373,N_12599,N_13232);
or U14374 (N_14374,N_13265,N_13047);
or U14375 (N_14375,N_13641,N_13024);
nor U14376 (N_14376,N_13359,N_12650);
xnor U14377 (N_14377,N_13734,N_13361);
or U14378 (N_14378,N_13244,N_13266);
and U14379 (N_14379,N_13684,N_13670);
nor U14380 (N_14380,N_12797,N_13733);
nand U14381 (N_14381,N_13577,N_13226);
and U14382 (N_14382,N_13454,N_12576);
and U14383 (N_14383,N_13324,N_13173);
xnor U14384 (N_14384,N_13267,N_12576);
xor U14385 (N_14385,N_12733,N_12559);
nand U14386 (N_14386,N_12946,N_12707);
or U14387 (N_14387,N_13354,N_13701);
or U14388 (N_14388,N_13444,N_13424);
nand U14389 (N_14389,N_13115,N_12853);
nand U14390 (N_14390,N_13421,N_13186);
xnor U14391 (N_14391,N_12899,N_12658);
nand U14392 (N_14392,N_12882,N_13004);
xnor U14393 (N_14393,N_12761,N_13026);
and U14394 (N_14394,N_12900,N_12511);
and U14395 (N_14395,N_12675,N_13102);
xnor U14396 (N_14396,N_13276,N_13425);
and U14397 (N_14397,N_13282,N_12620);
or U14398 (N_14398,N_13606,N_13313);
nor U14399 (N_14399,N_13613,N_13740);
or U14400 (N_14400,N_12700,N_13541);
nand U14401 (N_14401,N_13703,N_12686);
or U14402 (N_14402,N_13579,N_12880);
or U14403 (N_14403,N_13381,N_12757);
xnor U14404 (N_14404,N_13046,N_13112);
nand U14405 (N_14405,N_13420,N_13033);
or U14406 (N_14406,N_13040,N_13007);
and U14407 (N_14407,N_12843,N_12743);
or U14408 (N_14408,N_13729,N_13291);
nand U14409 (N_14409,N_13104,N_13503);
nand U14410 (N_14410,N_12856,N_13561);
and U14411 (N_14411,N_12755,N_12917);
nand U14412 (N_14412,N_12712,N_12559);
xnor U14413 (N_14413,N_13677,N_13610);
nor U14414 (N_14414,N_13420,N_13264);
nor U14415 (N_14415,N_13396,N_13724);
nor U14416 (N_14416,N_12982,N_13461);
and U14417 (N_14417,N_12522,N_12942);
nand U14418 (N_14418,N_13439,N_12601);
and U14419 (N_14419,N_13185,N_13486);
nor U14420 (N_14420,N_12535,N_13146);
nor U14421 (N_14421,N_13660,N_13607);
and U14422 (N_14422,N_13021,N_13081);
nor U14423 (N_14423,N_13125,N_12711);
nor U14424 (N_14424,N_13170,N_13513);
xnor U14425 (N_14425,N_12527,N_13406);
xnor U14426 (N_14426,N_13172,N_12543);
and U14427 (N_14427,N_13198,N_12844);
xor U14428 (N_14428,N_13509,N_13002);
nor U14429 (N_14429,N_12545,N_13284);
or U14430 (N_14430,N_13398,N_13359);
xor U14431 (N_14431,N_12909,N_13381);
and U14432 (N_14432,N_13025,N_13553);
or U14433 (N_14433,N_12673,N_13687);
nand U14434 (N_14434,N_13571,N_12522);
and U14435 (N_14435,N_13738,N_13666);
nand U14436 (N_14436,N_13050,N_13562);
nor U14437 (N_14437,N_13742,N_12632);
xnor U14438 (N_14438,N_13748,N_13057);
nor U14439 (N_14439,N_13727,N_12687);
xor U14440 (N_14440,N_13470,N_13483);
nor U14441 (N_14441,N_12733,N_13176);
nand U14442 (N_14442,N_13684,N_12795);
nand U14443 (N_14443,N_13404,N_13403);
and U14444 (N_14444,N_13277,N_13500);
xnor U14445 (N_14445,N_13253,N_12507);
or U14446 (N_14446,N_12967,N_13327);
or U14447 (N_14447,N_13466,N_12848);
and U14448 (N_14448,N_13431,N_12519);
xor U14449 (N_14449,N_13358,N_13573);
xnor U14450 (N_14450,N_13694,N_12544);
nor U14451 (N_14451,N_13433,N_12649);
nand U14452 (N_14452,N_12520,N_13301);
and U14453 (N_14453,N_13069,N_13273);
nor U14454 (N_14454,N_13264,N_13266);
or U14455 (N_14455,N_13637,N_13646);
nor U14456 (N_14456,N_13073,N_13219);
nand U14457 (N_14457,N_13593,N_13324);
nand U14458 (N_14458,N_13219,N_12918);
nor U14459 (N_14459,N_13238,N_13450);
nand U14460 (N_14460,N_12899,N_12712);
nor U14461 (N_14461,N_13198,N_12597);
and U14462 (N_14462,N_12893,N_12895);
xor U14463 (N_14463,N_13550,N_12863);
xnor U14464 (N_14464,N_12610,N_12884);
nand U14465 (N_14465,N_12843,N_12715);
and U14466 (N_14466,N_12567,N_12997);
nand U14467 (N_14467,N_12509,N_12515);
xnor U14468 (N_14468,N_12695,N_12567);
xnor U14469 (N_14469,N_13606,N_12755);
nand U14470 (N_14470,N_13024,N_13363);
nand U14471 (N_14471,N_12986,N_12752);
nor U14472 (N_14472,N_13444,N_13649);
nor U14473 (N_14473,N_12991,N_12725);
xor U14474 (N_14474,N_13068,N_12862);
and U14475 (N_14475,N_12572,N_12598);
nand U14476 (N_14476,N_13744,N_12845);
or U14477 (N_14477,N_12859,N_12633);
xnor U14478 (N_14478,N_13235,N_12573);
xor U14479 (N_14479,N_12883,N_12524);
or U14480 (N_14480,N_13664,N_12671);
and U14481 (N_14481,N_13399,N_12741);
and U14482 (N_14482,N_13615,N_13094);
xnor U14483 (N_14483,N_12548,N_13275);
or U14484 (N_14484,N_12950,N_13056);
nand U14485 (N_14485,N_13685,N_12709);
nor U14486 (N_14486,N_12832,N_13318);
nand U14487 (N_14487,N_12750,N_12602);
xnor U14488 (N_14488,N_12672,N_12847);
nor U14489 (N_14489,N_12571,N_12517);
or U14490 (N_14490,N_13711,N_13328);
nor U14491 (N_14491,N_13166,N_12847);
xor U14492 (N_14492,N_12564,N_12660);
and U14493 (N_14493,N_12800,N_13448);
nor U14494 (N_14494,N_12759,N_13310);
or U14495 (N_14495,N_13483,N_12661);
nor U14496 (N_14496,N_13151,N_12572);
or U14497 (N_14497,N_13386,N_12742);
nand U14498 (N_14498,N_12918,N_13630);
and U14499 (N_14499,N_13652,N_13137);
nand U14500 (N_14500,N_13191,N_13185);
xnor U14501 (N_14501,N_13405,N_13416);
or U14502 (N_14502,N_13161,N_12611);
nand U14503 (N_14503,N_12869,N_13443);
nand U14504 (N_14504,N_12566,N_13539);
nand U14505 (N_14505,N_13174,N_12698);
xor U14506 (N_14506,N_13257,N_13403);
or U14507 (N_14507,N_13713,N_13665);
or U14508 (N_14508,N_13354,N_13516);
nand U14509 (N_14509,N_13471,N_13240);
or U14510 (N_14510,N_12835,N_12963);
nand U14511 (N_14511,N_12735,N_13135);
xnor U14512 (N_14512,N_12899,N_13510);
nand U14513 (N_14513,N_12713,N_12879);
nand U14514 (N_14514,N_12712,N_13693);
and U14515 (N_14515,N_13470,N_13322);
or U14516 (N_14516,N_13676,N_13592);
xnor U14517 (N_14517,N_12880,N_12868);
or U14518 (N_14518,N_13482,N_12952);
or U14519 (N_14519,N_13323,N_12745);
nor U14520 (N_14520,N_13269,N_13333);
nor U14521 (N_14521,N_13361,N_13079);
xor U14522 (N_14522,N_13469,N_12602);
and U14523 (N_14523,N_12606,N_12782);
or U14524 (N_14524,N_13723,N_13594);
nor U14525 (N_14525,N_12971,N_13378);
and U14526 (N_14526,N_13526,N_12584);
or U14527 (N_14527,N_13487,N_13519);
or U14528 (N_14528,N_13366,N_12628);
nand U14529 (N_14529,N_13284,N_12917);
xnor U14530 (N_14530,N_12840,N_13485);
nand U14531 (N_14531,N_13572,N_13246);
nand U14532 (N_14532,N_12811,N_13595);
xor U14533 (N_14533,N_13504,N_12633);
and U14534 (N_14534,N_12696,N_12886);
xnor U14535 (N_14535,N_13522,N_12694);
nand U14536 (N_14536,N_13304,N_13000);
or U14537 (N_14537,N_13195,N_13504);
nor U14538 (N_14538,N_13580,N_13708);
or U14539 (N_14539,N_13263,N_12614);
nor U14540 (N_14540,N_13300,N_13016);
and U14541 (N_14541,N_13349,N_12829);
nor U14542 (N_14542,N_13239,N_13390);
nand U14543 (N_14543,N_12805,N_12927);
xor U14544 (N_14544,N_13295,N_12845);
or U14545 (N_14545,N_12829,N_13026);
or U14546 (N_14546,N_12800,N_13325);
or U14547 (N_14547,N_12752,N_12888);
and U14548 (N_14548,N_12515,N_13440);
nand U14549 (N_14549,N_13670,N_12926);
nand U14550 (N_14550,N_13242,N_13194);
xor U14551 (N_14551,N_13108,N_12592);
or U14552 (N_14552,N_13510,N_13700);
nand U14553 (N_14553,N_13748,N_12731);
nor U14554 (N_14554,N_13098,N_13253);
and U14555 (N_14555,N_13535,N_12566);
nor U14556 (N_14556,N_13407,N_12763);
nand U14557 (N_14557,N_12922,N_13631);
and U14558 (N_14558,N_13554,N_12502);
or U14559 (N_14559,N_12794,N_13724);
or U14560 (N_14560,N_13065,N_12674);
xor U14561 (N_14561,N_13437,N_13283);
and U14562 (N_14562,N_13423,N_12887);
nor U14563 (N_14563,N_13189,N_13370);
or U14564 (N_14564,N_12901,N_12580);
xor U14565 (N_14565,N_13251,N_12513);
or U14566 (N_14566,N_12611,N_13489);
and U14567 (N_14567,N_13589,N_13286);
and U14568 (N_14568,N_13713,N_12766);
and U14569 (N_14569,N_12920,N_13079);
nand U14570 (N_14570,N_12856,N_13215);
and U14571 (N_14571,N_13430,N_13656);
nand U14572 (N_14572,N_13693,N_12927);
xor U14573 (N_14573,N_13093,N_13662);
and U14574 (N_14574,N_12841,N_13434);
or U14575 (N_14575,N_13522,N_13262);
and U14576 (N_14576,N_12977,N_13349);
xor U14577 (N_14577,N_12752,N_13660);
xnor U14578 (N_14578,N_12622,N_12678);
nor U14579 (N_14579,N_12695,N_13111);
nor U14580 (N_14580,N_13544,N_13624);
nand U14581 (N_14581,N_12832,N_12910);
nor U14582 (N_14582,N_13295,N_13298);
xor U14583 (N_14583,N_13260,N_12778);
xnor U14584 (N_14584,N_13727,N_12539);
xor U14585 (N_14585,N_13495,N_13654);
nor U14586 (N_14586,N_13499,N_13217);
xor U14587 (N_14587,N_13009,N_12645);
xnor U14588 (N_14588,N_13178,N_13427);
or U14589 (N_14589,N_13015,N_13395);
or U14590 (N_14590,N_12688,N_12912);
nor U14591 (N_14591,N_13026,N_13340);
nor U14592 (N_14592,N_13597,N_13517);
nor U14593 (N_14593,N_12978,N_13393);
nor U14594 (N_14594,N_13238,N_13499);
nand U14595 (N_14595,N_13573,N_13123);
nor U14596 (N_14596,N_12851,N_13573);
xor U14597 (N_14597,N_13636,N_13042);
xor U14598 (N_14598,N_13080,N_12566);
and U14599 (N_14599,N_13517,N_13036);
nand U14600 (N_14600,N_13144,N_13039);
nand U14601 (N_14601,N_12918,N_13391);
nor U14602 (N_14602,N_12879,N_12645);
and U14603 (N_14603,N_13671,N_12517);
or U14604 (N_14604,N_13526,N_12622);
and U14605 (N_14605,N_13367,N_13390);
nand U14606 (N_14606,N_13498,N_13446);
xor U14607 (N_14607,N_12764,N_13320);
or U14608 (N_14608,N_13282,N_12968);
xor U14609 (N_14609,N_13215,N_13197);
or U14610 (N_14610,N_13148,N_13287);
xnor U14611 (N_14611,N_12575,N_12735);
and U14612 (N_14612,N_13054,N_12505);
nand U14613 (N_14613,N_13715,N_13177);
xnor U14614 (N_14614,N_13321,N_13239);
nand U14615 (N_14615,N_12873,N_13719);
and U14616 (N_14616,N_13005,N_13445);
xnor U14617 (N_14617,N_12514,N_12981);
nor U14618 (N_14618,N_13608,N_12956);
xnor U14619 (N_14619,N_13681,N_13087);
xnor U14620 (N_14620,N_13599,N_13035);
and U14621 (N_14621,N_12504,N_13112);
and U14622 (N_14622,N_13591,N_13165);
or U14623 (N_14623,N_13340,N_12911);
nor U14624 (N_14624,N_13653,N_13450);
nand U14625 (N_14625,N_13237,N_13252);
and U14626 (N_14626,N_13366,N_13655);
xor U14627 (N_14627,N_12995,N_12747);
and U14628 (N_14628,N_13621,N_12919);
nand U14629 (N_14629,N_12983,N_12794);
nor U14630 (N_14630,N_12817,N_12578);
or U14631 (N_14631,N_13063,N_13162);
or U14632 (N_14632,N_12844,N_13401);
nor U14633 (N_14633,N_12713,N_12946);
or U14634 (N_14634,N_13144,N_13238);
nand U14635 (N_14635,N_12934,N_13213);
or U14636 (N_14636,N_12798,N_13680);
nand U14637 (N_14637,N_13312,N_13371);
xnor U14638 (N_14638,N_13284,N_12749);
xnor U14639 (N_14639,N_12531,N_12828);
nand U14640 (N_14640,N_13552,N_12627);
or U14641 (N_14641,N_13264,N_12861);
or U14642 (N_14642,N_13532,N_13410);
nor U14643 (N_14643,N_13450,N_13580);
or U14644 (N_14644,N_12559,N_13159);
nand U14645 (N_14645,N_13720,N_13345);
and U14646 (N_14646,N_13145,N_13033);
xor U14647 (N_14647,N_13200,N_13308);
or U14648 (N_14648,N_13371,N_13703);
nor U14649 (N_14649,N_12922,N_12866);
or U14650 (N_14650,N_13695,N_13022);
and U14651 (N_14651,N_13020,N_13473);
and U14652 (N_14652,N_13446,N_12554);
xnor U14653 (N_14653,N_13006,N_13294);
and U14654 (N_14654,N_12925,N_12779);
and U14655 (N_14655,N_13341,N_13404);
xnor U14656 (N_14656,N_13219,N_13512);
and U14657 (N_14657,N_12875,N_13656);
xnor U14658 (N_14658,N_12945,N_12700);
or U14659 (N_14659,N_13100,N_12810);
and U14660 (N_14660,N_13706,N_13414);
nand U14661 (N_14661,N_13717,N_13195);
nor U14662 (N_14662,N_13264,N_13319);
xnor U14663 (N_14663,N_13309,N_13305);
xor U14664 (N_14664,N_13141,N_13736);
and U14665 (N_14665,N_13354,N_13381);
and U14666 (N_14666,N_12893,N_12689);
nand U14667 (N_14667,N_12754,N_13376);
nor U14668 (N_14668,N_13111,N_13365);
nor U14669 (N_14669,N_12712,N_12806);
and U14670 (N_14670,N_13178,N_12727);
nand U14671 (N_14671,N_12647,N_13299);
nor U14672 (N_14672,N_13050,N_12695);
and U14673 (N_14673,N_13630,N_12625);
nand U14674 (N_14674,N_12966,N_13643);
and U14675 (N_14675,N_13198,N_13428);
nand U14676 (N_14676,N_13111,N_13462);
xor U14677 (N_14677,N_13242,N_13360);
or U14678 (N_14678,N_13113,N_13513);
and U14679 (N_14679,N_13452,N_13185);
and U14680 (N_14680,N_13156,N_13507);
or U14681 (N_14681,N_12946,N_13492);
nor U14682 (N_14682,N_13362,N_13197);
and U14683 (N_14683,N_12746,N_13232);
nor U14684 (N_14684,N_12705,N_13663);
xor U14685 (N_14685,N_13081,N_13001);
or U14686 (N_14686,N_12717,N_13435);
and U14687 (N_14687,N_12812,N_13220);
nor U14688 (N_14688,N_12911,N_13294);
xor U14689 (N_14689,N_13076,N_12620);
xor U14690 (N_14690,N_13024,N_13714);
nor U14691 (N_14691,N_12660,N_13508);
xnor U14692 (N_14692,N_12790,N_13591);
or U14693 (N_14693,N_12782,N_13408);
nand U14694 (N_14694,N_13269,N_12505);
nor U14695 (N_14695,N_13088,N_13638);
nor U14696 (N_14696,N_12778,N_13280);
and U14697 (N_14697,N_13642,N_13610);
xnor U14698 (N_14698,N_13065,N_12798);
nor U14699 (N_14699,N_13191,N_12561);
or U14700 (N_14700,N_13232,N_12630);
nor U14701 (N_14701,N_12771,N_12638);
nand U14702 (N_14702,N_13483,N_12642);
xor U14703 (N_14703,N_12712,N_13587);
xnor U14704 (N_14704,N_13556,N_13585);
nor U14705 (N_14705,N_13439,N_13267);
nand U14706 (N_14706,N_12536,N_13177);
nand U14707 (N_14707,N_13648,N_13426);
or U14708 (N_14708,N_13207,N_13273);
or U14709 (N_14709,N_13159,N_12936);
nor U14710 (N_14710,N_12631,N_13681);
nor U14711 (N_14711,N_12533,N_12929);
nor U14712 (N_14712,N_12976,N_12846);
nand U14713 (N_14713,N_12815,N_13272);
and U14714 (N_14714,N_12757,N_12976);
xnor U14715 (N_14715,N_12706,N_12971);
or U14716 (N_14716,N_13543,N_12514);
xor U14717 (N_14717,N_13142,N_13135);
nor U14718 (N_14718,N_13314,N_13196);
or U14719 (N_14719,N_13016,N_13154);
or U14720 (N_14720,N_13311,N_13151);
nor U14721 (N_14721,N_13552,N_13639);
xor U14722 (N_14722,N_13154,N_12752);
xor U14723 (N_14723,N_13379,N_13319);
nor U14724 (N_14724,N_13351,N_12882);
or U14725 (N_14725,N_12811,N_12634);
nor U14726 (N_14726,N_12527,N_13618);
nand U14727 (N_14727,N_12759,N_13549);
nand U14728 (N_14728,N_13643,N_13672);
and U14729 (N_14729,N_12923,N_12990);
nor U14730 (N_14730,N_13356,N_13564);
nand U14731 (N_14731,N_13178,N_13028);
nand U14732 (N_14732,N_12744,N_13462);
xnor U14733 (N_14733,N_12798,N_13458);
nand U14734 (N_14734,N_12714,N_13061);
or U14735 (N_14735,N_12828,N_12523);
nor U14736 (N_14736,N_13525,N_13567);
and U14737 (N_14737,N_12957,N_12509);
nand U14738 (N_14738,N_12564,N_13434);
or U14739 (N_14739,N_12744,N_13470);
nand U14740 (N_14740,N_13673,N_13620);
or U14741 (N_14741,N_13728,N_12775);
or U14742 (N_14742,N_12664,N_13271);
nor U14743 (N_14743,N_12781,N_13626);
nand U14744 (N_14744,N_12884,N_13613);
nor U14745 (N_14745,N_13541,N_12795);
xor U14746 (N_14746,N_12571,N_13575);
xnor U14747 (N_14747,N_13605,N_12560);
nor U14748 (N_14748,N_13268,N_12631);
and U14749 (N_14749,N_12763,N_13258);
xor U14750 (N_14750,N_13195,N_13246);
xnor U14751 (N_14751,N_12706,N_13333);
nor U14752 (N_14752,N_13298,N_13210);
nand U14753 (N_14753,N_13135,N_13107);
and U14754 (N_14754,N_12612,N_13546);
or U14755 (N_14755,N_12689,N_12913);
or U14756 (N_14756,N_13465,N_13709);
xor U14757 (N_14757,N_13596,N_13081);
or U14758 (N_14758,N_13747,N_12961);
or U14759 (N_14759,N_12871,N_13308);
nand U14760 (N_14760,N_13633,N_13727);
and U14761 (N_14761,N_13320,N_13323);
or U14762 (N_14762,N_13334,N_13581);
nor U14763 (N_14763,N_12595,N_13485);
and U14764 (N_14764,N_13176,N_13394);
xnor U14765 (N_14765,N_13341,N_13603);
or U14766 (N_14766,N_12853,N_13427);
and U14767 (N_14767,N_13204,N_13003);
and U14768 (N_14768,N_13708,N_12511);
nand U14769 (N_14769,N_13003,N_13361);
xnor U14770 (N_14770,N_13402,N_12944);
or U14771 (N_14771,N_12713,N_13154);
nand U14772 (N_14772,N_13133,N_12593);
nand U14773 (N_14773,N_12644,N_12932);
nor U14774 (N_14774,N_12512,N_13379);
nand U14775 (N_14775,N_12669,N_13423);
or U14776 (N_14776,N_12889,N_13233);
or U14777 (N_14777,N_12811,N_13487);
nor U14778 (N_14778,N_12525,N_13663);
nand U14779 (N_14779,N_13575,N_13531);
or U14780 (N_14780,N_13588,N_13494);
nand U14781 (N_14781,N_13467,N_12908);
or U14782 (N_14782,N_13203,N_13564);
nor U14783 (N_14783,N_13177,N_12907);
or U14784 (N_14784,N_13333,N_13559);
nand U14785 (N_14785,N_13721,N_13131);
and U14786 (N_14786,N_12800,N_12737);
nor U14787 (N_14787,N_13349,N_13402);
or U14788 (N_14788,N_12802,N_13511);
and U14789 (N_14789,N_13022,N_13020);
nor U14790 (N_14790,N_12882,N_13666);
or U14791 (N_14791,N_13236,N_12713);
and U14792 (N_14792,N_13330,N_13114);
xor U14793 (N_14793,N_13386,N_13687);
and U14794 (N_14794,N_13348,N_12763);
and U14795 (N_14795,N_13161,N_13434);
and U14796 (N_14796,N_13061,N_13710);
nand U14797 (N_14797,N_12900,N_12728);
xnor U14798 (N_14798,N_12683,N_13261);
nand U14799 (N_14799,N_13605,N_13731);
or U14800 (N_14800,N_12705,N_13519);
or U14801 (N_14801,N_13144,N_13134);
xor U14802 (N_14802,N_13643,N_12588);
xor U14803 (N_14803,N_13582,N_12568);
or U14804 (N_14804,N_13206,N_12592);
and U14805 (N_14805,N_13598,N_13238);
nand U14806 (N_14806,N_13197,N_13665);
nor U14807 (N_14807,N_13682,N_13482);
xnor U14808 (N_14808,N_13605,N_12851);
nor U14809 (N_14809,N_12933,N_12934);
xnor U14810 (N_14810,N_12889,N_12552);
xnor U14811 (N_14811,N_12569,N_13200);
or U14812 (N_14812,N_12698,N_13453);
nor U14813 (N_14813,N_13419,N_12725);
nand U14814 (N_14814,N_12747,N_12513);
nand U14815 (N_14815,N_13026,N_13475);
nand U14816 (N_14816,N_12910,N_13089);
nor U14817 (N_14817,N_13284,N_13485);
nor U14818 (N_14818,N_12615,N_12756);
nor U14819 (N_14819,N_12994,N_13332);
nand U14820 (N_14820,N_13273,N_12627);
and U14821 (N_14821,N_13585,N_12844);
nor U14822 (N_14822,N_13204,N_13084);
nand U14823 (N_14823,N_13171,N_12929);
nor U14824 (N_14824,N_13178,N_13014);
nand U14825 (N_14825,N_13578,N_12542);
nor U14826 (N_14826,N_13186,N_13295);
nand U14827 (N_14827,N_13538,N_13070);
nand U14828 (N_14828,N_13747,N_13262);
and U14829 (N_14829,N_13654,N_13133);
and U14830 (N_14830,N_13658,N_12834);
and U14831 (N_14831,N_13263,N_12896);
nand U14832 (N_14832,N_13633,N_13189);
xor U14833 (N_14833,N_13682,N_12678);
nand U14834 (N_14834,N_12506,N_13053);
nand U14835 (N_14835,N_12694,N_13351);
and U14836 (N_14836,N_12846,N_13115);
and U14837 (N_14837,N_13648,N_12515);
and U14838 (N_14838,N_13442,N_13323);
xnor U14839 (N_14839,N_12538,N_13711);
nor U14840 (N_14840,N_12541,N_12784);
nand U14841 (N_14841,N_13100,N_13639);
nor U14842 (N_14842,N_13611,N_13597);
nand U14843 (N_14843,N_13709,N_12677);
and U14844 (N_14844,N_13382,N_12826);
nor U14845 (N_14845,N_13163,N_12668);
and U14846 (N_14846,N_13215,N_13547);
and U14847 (N_14847,N_13304,N_13677);
nand U14848 (N_14848,N_12560,N_13118);
nand U14849 (N_14849,N_13543,N_13498);
or U14850 (N_14850,N_12692,N_12932);
and U14851 (N_14851,N_13060,N_13734);
nor U14852 (N_14852,N_12813,N_13481);
xor U14853 (N_14853,N_13087,N_13537);
xor U14854 (N_14854,N_13109,N_13695);
xor U14855 (N_14855,N_12904,N_12654);
nor U14856 (N_14856,N_13143,N_13386);
and U14857 (N_14857,N_12923,N_12889);
and U14858 (N_14858,N_12873,N_12976);
xnor U14859 (N_14859,N_12937,N_12655);
xnor U14860 (N_14860,N_13446,N_13668);
nor U14861 (N_14861,N_13151,N_12627);
or U14862 (N_14862,N_13519,N_13140);
nor U14863 (N_14863,N_12692,N_13417);
nand U14864 (N_14864,N_12757,N_12863);
nand U14865 (N_14865,N_13130,N_12857);
nor U14866 (N_14866,N_13182,N_13697);
xnor U14867 (N_14867,N_12641,N_12799);
nor U14868 (N_14868,N_12881,N_13211);
and U14869 (N_14869,N_13360,N_13387);
and U14870 (N_14870,N_12931,N_13208);
or U14871 (N_14871,N_13577,N_12536);
nand U14872 (N_14872,N_12762,N_13007);
nor U14873 (N_14873,N_13156,N_13395);
or U14874 (N_14874,N_12999,N_13017);
and U14875 (N_14875,N_13486,N_13080);
and U14876 (N_14876,N_12940,N_13111);
nor U14877 (N_14877,N_13120,N_13451);
and U14878 (N_14878,N_13486,N_13600);
nand U14879 (N_14879,N_12726,N_13454);
nand U14880 (N_14880,N_13298,N_13558);
xnor U14881 (N_14881,N_12519,N_13208);
or U14882 (N_14882,N_12730,N_13065);
nor U14883 (N_14883,N_12709,N_13099);
nor U14884 (N_14884,N_12988,N_13356);
and U14885 (N_14885,N_13249,N_13564);
nand U14886 (N_14886,N_13276,N_13731);
nor U14887 (N_14887,N_13176,N_13308);
nor U14888 (N_14888,N_13198,N_12614);
or U14889 (N_14889,N_12704,N_13615);
or U14890 (N_14890,N_12606,N_13588);
nand U14891 (N_14891,N_12978,N_13014);
and U14892 (N_14892,N_13564,N_13682);
xnor U14893 (N_14893,N_13412,N_13073);
or U14894 (N_14894,N_13442,N_13139);
nand U14895 (N_14895,N_13341,N_13079);
and U14896 (N_14896,N_12675,N_13425);
and U14897 (N_14897,N_13375,N_13051);
nand U14898 (N_14898,N_13009,N_13557);
nor U14899 (N_14899,N_12552,N_13434);
and U14900 (N_14900,N_13056,N_13345);
or U14901 (N_14901,N_13710,N_13464);
xor U14902 (N_14902,N_13671,N_13126);
nand U14903 (N_14903,N_13153,N_12902);
nor U14904 (N_14904,N_12966,N_13023);
nor U14905 (N_14905,N_13349,N_13729);
and U14906 (N_14906,N_13742,N_12709);
nor U14907 (N_14907,N_13499,N_12601);
nor U14908 (N_14908,N_12729,N_13563);
or U14909 (N_14909,N_12910,N_12710);
or U14910 (N_14910,N_13644,N_13140);
nand U14911 (N_14911,N_12948,N_12614);
and U14912 (N_14912,N_13709,N_12879);
or U14913 (N_14913,N_13254,N_13023);
nand U14914 (N_14914,N_13440,N_13508);
xor U14915 (N_14915,N_12651,N_12513);
nand U14916 (N_14916,N_13161,N_13688);
nand U14917 (N_14917,N_12627,N_12816);
nor U14918 (N_14918,N_13679,N_13429);
nor U14919 (N_14919,N_13694,N_13090);
xnor U14920 (N_14920,N_12790,N_12967);
and U14921 (N_14921,N_13636,N_13088);
or U14922 (N_14922,N_13737,N_13261);
nand U14923 (N_14923,N_12869,N_12813);
xor U14924 (N_14924,N_13366,N_13269);
and U14925 (N_14925,N_13360,N_13652);
nor U14926 (N_14926,N_13313,N_12666);
xnor U14927 (N_14927,N_13697,N_13041);
xnor U14928 (N_14928,N_13057,N_12904);
xnor U14929 (N_14929,N_13559,N_13744);
nand U14930 (N_14930,N_13598,N_12534);
or U14931 (N_14931,N_13718,N_13156);
and U14932 (N_14932,N_13201,N_13650);
xnor U14933 (N_14933,N_13254,N_12649);
xor U14934 (N_14934,N_13559,N_13022);
or U14935 (N_14935,N_13156,N_12806);
nand U14936 (N_14936,N_13142,N_13192);
nor U14937 (N_14937,N_13228,N_12810);
nand U14938 (N_14938,N_13350,N_13383);
and U14939 (N_14939,N_12823,N_12841);
or U14940 (N_14940,N_12685,N_12921);
xor U14941 (N_14941,N_13685,N_13347);
nand U14942 (N_14942,N_13032,N_13651);
and U14943 (N_14943,N_12822,N_12721);
xnor U14944 (N_14944,N_13353,N_13425);
and U14945 (N_14945,N_13563,N_13593);
xor U14946 (N_14946,N_12994,N_13385);
nor U14947 (N_14947,N_12920,N_13502);
nand U14948 (N_14948,N_13457,N_12630);
xor U14949 (N_14949,N_13400,N_13732);
or U14950 (N_14950,N_13326,N_13325);
or U14951 (N_14951,N_12877,N_13380);
or U14952 (N_14952,N_12853,N_12687);
or U14953 (N_14953,N_13148,N_13455);
nand U14954 (N_14954,N_13742,N_13329);
and U14955 (N_14955,N_12772,N_13133);
nor U14956 (N_14956,N_13316,N_13020);
or U14957 (N_14957,N_13075,N_12568);
xnor U14958 (N_14958,N_12784,N_13369);
nor U14959 (N_14959,N_13184,N_13200);
and U14960 (N_14960,N_13511,N_12970);
and U14961 (N_14961,N_13676,N_12716);
nor U14962 (N_14962,N_12719,N_13618);
nor U14963 (N_14963,N_13587,N_12691);
or U14964 (N_14964,N_13471,N_12797);
or U14965 (N_14965,N_13124,N_13035);
nand U14966 (N_14966,N_12868,N_13521);
and U14967 (N_14967,N_12713,N_12607);
nor U14968 (N_14968,N_13680,N_13229);
and U14969 (N_14969,N_13494,N_12595);
and U14970 (N_14970,N_12754,N_13630);
nand U14971 (N_14971,N_12680,N_13454);
nand U14972 (N_14972,N_12625,N_13687);
nor U14973 (N_14973,N_13349,N_12554);
nand U14974 (N_14974,N_13395,N_12714);
nand U14975 (N_14975,N_12779,N_13156);
and U14976 (N_14976,N_13465,N_12701);
nor U14977 (N_14977,N_13741,N_12985);
nand U14978 (N_14978,N_13539,N_12635);
or U14979 (N_14979,N_13276,N_13531);
and U14980 (N_14980,N_12664,N_13367);
nor U14981 (N_14981,N_13325,N_13484);
nor U14982 (N_14982,N_12863,N_13002);
xor U14983 (N_14983,N_13618,N_13134);
nand U14984 (N_14984,N_13208,N_13468);
xor U14985 (N_14985,N_13541,N_12512);
nor U14986 (N_14986,N_12778,N_13121);
nor U14987 (N_14987,N_13262,N_12611);
xnor U14988 (N_14988,N_12672,N_13164);
nand U14989 (N_14989,N_12776,N_13008);
and U14990 (N_14990,N_12875,N_13006);
or U14991 (N_14991,N_13355,N_13237);
or U14992 (N_14992,N_12714,N_13398);
and U14993 (N_14993,N_13240,N_13593);
xor U14994 (N_14994,N_12531,N_12963);
or U14995 (N_14995,N_13214,N_12658);
xnor U14996 (N_14996,N_12700,N_13435);
nor U14997 (N_14997,N_12678,N_13215);
and U14998 (N_14998,N_12765,N_13197);
nor U14999 (N_14999,N_13507,N_12661);
nor U15000 (N_15000,N_14441,N_14569);
and U15001 (N_15001,N_14493,N_14464);
xor U15002 (N_15002,N_14728,N_14394);
nor U15003 (N_15003,N_13759,N_14781);
xnor U15004 (N_15004,N_14962,N_13947);
xor U15005 (N_15005,N_14011,N_14621);
nand U15006 (N_15006,N_13770,N_14788);
or U15007 (N_15007,N_14852,N_14793);
nor U15008 (N_15008,N_14666,N_14660);
and U15009 (N_15009,N_13940,N_14300);
and U15010 (N_15010,N_13804,N_14632);
xnor U15011 (N_15011,N_14599,N_14035);
and U15012 (N_15012,N_14884,N_14880);
nor U15013 (N_15013,N_13831,N_14401);
or U15014 (N_15014,N_14506,N_14164);
and U15015 (N_15015,N_14996,N_14715);
and U15016 (N_15016,N_14610,N_14624);
xor U15017 (N_15017,N_14501,N_14130);
nand U15018 (N_15018,N_14020,N_14830);
and U15019 (N_15019,N_14120,N_14053);
xor U15020 (N_15020,N_14057,N_14301);
nor U15021 (N_15021,N_14922,N_14832);
nand U15022 (N_15022,N_13873,N_14315);
xnor U15023 (N_15023,N_14959,N_13994);
xnor U15024 (N_15024,N_14477,N_14458);
nand U15025 (N_15025,N_14491,N_14432);
and U15026 (N_15026,N_14245,N_14606);
xor U15027 (N_15027,N_14290,N_14356);
nand U15028 (N_15028,N_13837,N_13761);
xnor U15029 (N_15029,N_14986,N_14088);
or U15030 (N_15030,N_14327,N_14400);
and U15031 (N_15031,N_14982,N_14620);
and U15032 (N_15032,N_13984,N_14083);
nand U15033 (N_15033,N_13787,N_14670);
or U15034 (N_15034,N_14039,N_14686);
nor U15035 (N_15035,N_14304,N_13754);
xor U15036 (N_15036,N_13893,N_13896);
and U15037 (N_15037,N_14641,N_14581);
nand U15038 (N_15038,N_13806,N_14177);
xor U15039 (N_15039,N_13865,N_14133);
xor U15040 (N_15040,N_14752,N_14135);
nand U15041 (N_15041,N_14407,N_14071);
xnor U15042 (N_15042,N_14764,N_14845);
and U15043 (N_15043,N_13906,N_14368);
or U15044 (N_15044,N_14612,N_14643);
or U15045 (N_15045,N_14224,N_13939);
nor U15046 (N_15046,N_14983,N_14722);
or U15047 (N_15047,N_14635,N_14556);
and U15048 (N_15048,N_14820,N_14408);
or U15049 (N_15049,N_14848,N_14834);
nand U15050 (N_15050,N_14495,N_14257);
and U15051 (N_15051,N_14345,N_13913);
xnor U15052 (N_15052,N_13857,N_14409);
nor U15053 (N_15053,N_13853,N_14534);
or U15054 (N_15054,N_13842,N_14840);
xor U15055 (N_15055,N_13963,N_13983);
or U15056 (N_15056,N_14141,N_14402);
nor U15057 (N_15057,N_13791,N_14759);
nand U15058 (N_15058,N_14067,N_14069);
xor U15059 (N_15059,N_14523,N_14530);
or U15060 (N_15060,N_14614,N_14563);
and U15061 (N_15061,N_14335,N_14961);
nor U15062 (N_15062,N_13960,N_14077);
nand U15063 (N_15063,N_14924,N_13845);
nor U15064 (N_15064,N_13860,N_14931);
nand U15065 (N_15065,N_14898,N_14994);
nor U15066 (N_15066,N_13779,N_14419);
nand U15067 (N_15067,N_14700,N_14453);
xor U15068 (N_15068,N_13861,N_14242);
nor U15069 (N_15069,N_14307,N_14566);
nand U15070 (N_15070,N_14559,N_14062);
or U15071 (N_15071,N_14956,N_13924);
nor U15072 (N_15072,N_14582,N_14321);
or U15073 (N_15073,N_14010,N_14138);
and U15074 (N_15074,N_14425,N_14452);
xnor U15075 (N_15075,N_14763,N_14435);
nor U15076 (N_15076,N_14705,N_14951);
or U15077 (N_15077,N_13829,N_14762);
and U15078 (N_15078,N_14656,N_14333);
and U15079 (N_15079,N_14704,N_14339);
xnor U15080 (N_15080,N_14689,N_13941);
nand U15081 (N_15081,N_14917,N_14776);
and U15082 (N_15082,N_14462,N_14919);
xnor U15083 (N_15083,N_14168,N_14483);
and U15084 (N_15084,N_14795,N_14151);
nand U15085 (N_15085,N_13858,N_13789);
or U15086 (N_15086,N_14433,N_14388);
xnor U15087 (N_15087,N_14169,N_14851);
and U15088 (N_15088,N_14343,N_14977);
or U15089 (N_15089,N_14743,N_14264);
or U15090 (N_15090,N_14791,N_14017);
and U15091 (N_15091,N_14831,N_13768);
or U15092 (N_15092,N_14420,N_14351);
nand U15093 (N_15093,N_14357,N_13929);
and U15094 (N_15094,N_14173,N_14219);
xor U15095 (N_15095,N_14756,N_14591);
nand U15096 (N_15096,N_14080,N_14730);
xor U15097 (N_15097,N_14528,N_13894);
or U15098 (N_15098,N_14204,N_14803);
or U15099 (N_15099,N_14214,N_14933);
nor U15100 (N_15100,N_14480,N_13822);
or U15101 (N_15101,N_14560,N_14627);
nand U15102 (N_15102,N_14004,N_14934);
or U15103 (N_15103,N_14985,N_14331);
nor U15104 (N_15104,N_13867,N_13952);
nor U15105 (N_15105,N_14529,N_14045);
and U15106 (N_15106,N_13883,N_13820);
or U15107 (N_15107,N_14023,N_13840);
nor U15108 (N_15108,N_14340,N_14174);
or U15109 (N_15109,N_14690,N_13856);
and U15110 (N_15110,N_14395,N_14222);
xnor U15111 (N_15111,N_13943,N_14892);
and U15112 (N_15112,N_14123,N_14719);
and U15113 (N_15113,N_13846,N_14829);
nor U15114 (N_15114,N_14548,N_13854);
nand U15115 (N_15115,N_14244,N_14811);
or U15116 (N_15116,N_14552,N_14481);
or U15117 (N_15117,N_14276,N_14887);
or U15118 (N_15118,N_14555,N_13922);
nand U15119 (N_15119,N_14541,N_14472);
and U15120 (N_15120,N_14052,N_14850);
or U15121 (N_15121,N_14981,N_14201);
and U15122 (N_15122,N_14826,N_13851);
nor U15123 (N_15123,N_14187,N_13895);
nor U15124 (N_15124,N_14888,N_14303);
nor U15125 (N_15125,N_14094,N_13830);
xnor U15126 (N_15126,N_14103,N_14058);
and U15127 (N_15127,N_14841,N_14564);
xnor U15128 (N_15128,N_14590,N_13821);
nand U15129 (N_15129,N_14682,N_14142);
nand U15130 (N_15130,N_13987,N_14007);
and U15131 (N_15131,N_14256,N_14298);
or U15132 (N_15132,N_14267,N_14740);
nand U15133 (N_15133,N_14212,N_14218);
xor U15134 (N_15134,N_14270,N_14097);
xnor U15135 (N_15135,N_13931,N_14248);
and U15136 (N_15136,N_14561,N_14325);
and U15137 (N_15137,N_13801,N_14733);
xor U15138 (N_15138,N_14623,N_14678);
nor U15139 (N_15139,N_13962,N_14991);
nor U15140 (N_15140,N_14289,N_14794);
or U15141 (N_15141,N_14939,N_14968);
or U15142 (N_15142,N_14283,N_14596);
and U15143 (N_15143,N_13833,N_14954);
xor U15144 (N_15144,N_14551,N_14602);
and U15145 (N_15145,N_14717,N_14751);
or U15146 (N_15146,N_14935,N_14595);
and U15147 (N_15147,N_14861,N_13781);
xor U15148 (N_15148,N_14215,N_14777);
nand U15149 (N_15149,N_14577,N_14466);
and U15150 (N_15150,N_14771,N_14953);
nor U15151 (N_15151,N_14238,N_14901);
nor U15152 (N_15152,N_13797,N_13888);
nor U15153 (N_15153,N_14874,N_14391);
nor U15154 (N_15154,N_14658,N_13911);
nor U15155 (N_15155,N_14191,N_14636);
nor U15156 (N_15156,N_14910,N_14765);
nor U15157 (N_15157,N_14909,N_13945);
xor U15158 (N_15158,N_14687,N_13998);
nand U15159 (N_15159,N_14363,N_14118);
xor U15160 (N_15160,N_14279,N_14378);
nor U15161 (N_15161,N_13881,N_14948);
nand U15162 (N_15162,N_14511,N_13986);
xnor U15163 (N_15163,N_14475,N_14463);
xor U15164 (N_15164,N_14639,N_14676);
and U15165 (N_15165,N_14825,N_14865);
or U15166 (N_15166,N_14457,N_14504);
nand U15167 (N_15167,N_14448,N_14027);
xnor U15168 (N_15168,N_13902,N_14306);
and U15169 (N_15169,N_14232,N_14586);
xor U15170 (N_15170,N_14359,N_14099);
nor U15171 (N_15171,N_14593,N_14072);
nand U15172 (N_15172,N_13850,N_14611);
xor U15173 (N_15173,N_14040,N_14721);
xor U15174 (N_15174,N_14854,N_13967);
and U15175 (N_15175,N_14437,N_14942);
xnor U15176 (N_15176,N_14720,N_14474);
or U15177 (N_15177,N_13874,N_14422);
and U15178 (N_15178,N_14317,N_13961);
or U15179 (N_15179,N_14927,N_14813);
xor U15180 (N_15180,N_14877,N_14410);
nor U15181 (N_15181,N_14881,N_14055);
nand U15182 (N_15182,N_14833,N_13977);
xor U15183 (N_15183,N_14239,N_14698);
nor U15184 (N_15184,N_14426,N_14160);
nand U15185 (N_15185,N_14443,N_14312);
xnor U15186 (N_15186,N_14945,N_14478);
and U15187 (N_15187,N_13969,N_14638);
or U15188 (N_15188,N_14159,N_14546);
or U15189 (N_15189,N_14873,N_14059);
xor U15190 (N_15190,N_14181,N_14547);
and U15191 (N_15191,N_13944,N_14882);
nor U15192 (N_15192,N_14872,N_14185);
or U15193 (N_15193,N_14914,N_14467);
or U15194 (N_15194,N_13885,N_14015);
or U15195 (N_15195,N_14140,N_14487);
xnor U15196 (N_15196,N_14253,N_14685);
xnor U15197 (N_15197,N_14585,N_14318);
or U15198 (N_15198,N_14309,N_14930);
or U15199 (N_15199,N_14411,N_14938);
nor U15200 (N_15200,N_13920,N_14489);
nand U15201 (N_15201,N_14579,N_14696);
xor U15202 (N_15202,N_14347,N_14255);
nand U15203 (N_15203,N_14320,N_13886);
xor U15204 (N_15204,N_14943,N_14600);
nor U15205 (N_15205,N_14044,N_14194);
and U15206 (N_15206,N_14659,N_14093);
and U15207 (N_15207,N_14384,N_13777);
nand U15208 (N_15208,N_14758,N_14047);
and U15209 (N_15209,N_14139,N_14060);
or U15210 (N_15210,N_14005,N_14221);
xnor U15211 (N_15211,N_14937,N_13774);
nor U15212 (N_15212,N_14427,N_13869);
or U15213 (N_15213,N_13772,N_14625);
or U15214 (N_15214,N_14000,N_14476);
or U15215 (N_15215,N_13852,N_14512);
and U15216 (N_15216,N_14054,N_14184);
and U15217 (N_15217,N_14471,N_14513);
nor U15218 (N_15218,N_14669,N_13786);
xnor U15219 (N_15219,N_13766,N_14167);
xor U15220 (N_15220,N_13762,N_14397);
or U15221 (N_15221,N_13782,N_14598);
or U15222 (N_15222,N_14175,N_14308);
xnor U15223 (N_15223,N_14389,N_13892);
nor U15224 (N_15224,N_14946,N_14087);
nand U15225 (N_15225,N_14226,N_14386);
and U15226 (N_15226,N_14490,N_14692);
xor U15227 (N_15227,N_14860,N_14430);
xnor U15228 (N_15228,N_13758,N_13810);
and U15229 (N_15229,N_14744,N_14774);
xnor U15230 (N_15230,N_14371,N_14905);
nand U15231 (N_15231,N_14580,N_13949);
or U15232 (N_15232,N_14767,N_13799);
xor U15233 (N_15233,N_14147,N_14583);
and U15234 (N_15234,N_13910,N_14172);
nor U15235 (N_15235,N_14111,N_14890);
nand U15236 (N_15236,N_14739,N_13903);
nor U15237 (N_15237,N_14979,N_14429);
and U15238 (N_15238,N_14835,N_14274);
or U15239 (N_15239,N_14233,N_14112);
nor U15240 (N_15240,N_14036,N_14646);
and U15241 (N_15241,N_14921,N_14916);
nand U15242 (N_15242,N_13790,N_13993);
and U15243 (N_15243,N_14864,N_14906);
or U15244 (N_15244,N_13841,N_14545);
and U15245 (N_15245,N_14502,N_14373);
xor U15246 (N_15246,N_13935,N_14500);
and U15247 (N_15247,N_14984,N_14869);
or U15248 (N_15248,N_14423,N_14271);
nand U15249 (N_15249,N_14246,N_14786);
or U15250 (N_15250,N_14361,N_14497);
nand U15251 (N_15251,N_13832,N_14154);
xnor U15252 (N_15252,N_14724,N_13926);
xor U15253 (N_15253,N_14405,N_14428);
and U15254 (N_15254,N_13909,N_14499);
nor U15255 (N_15255,N_13828,N_14421);
nand U15256 (N_15256,N_14323,N_13763);
nand U15257 (N_15257,N_14104,N_14209);
and U15258 (N_15258,N_14971,N_13827);
nor U15259 (N_15259,N_13976,N_14470);
or U15260 (N_15260,N_13991,N_14285);
nand U15261 (N_15261,N_14542,N_14671);
xor U15262 (N_15262,N_14714,N_14216);
and U15263 (N_15263,N_14261,N_14498);
xnor U15264 (N_15264,N_14012,N_14859);
nand U15265 (N_15265,N_14137,N_14263);
nor U15266 (N_15266,N_13925,N_14353);
nand U15267 (N_15267,N_14090,N_14597);
or U15268 (N_15268,N_14667,N_14073);
or U15269 (N_15269,N_14182,N_14757);
nand U15270 (N_15270,N_14379,N_14157);
xor U15271 (N_15271,N_14124,N_14867);
and U15272 (N_15272,N_14192,N_13788);
nor U15273 (N_15273,N_14230,N_14125);
nand U15274 (N_15274,N_14254,N_14642);
xor U15275 (N_15275,N_14640,N_14179);
nand U15276 (N_15276,N_14079,N_13884);
or U15277 (N_15277,N_14695,N_14899);
nand U15278 (N_15278,N_14568,N_14608);
nand U15279 (N_15279,N_14106,N_14521);
or U15280 (N_15280,N_13819,N_14358);
nor U15281 (N_15281,N_14710,N_14749);
nand U15282 (N_15282,N_14115,N_14114);
nor U15283 (N_15283,N_14348,N_14615);
and U15284 (N_15284,N_14101,N_14863);
nand U15285 (N_15285,N_14839,N_14126);
nor U15286 (N_15286,N_14197,N_14494);
nor U15287 (N_15287,N_14925,N_14664);
and U15288 (N_15288,N_14171,N_14442);
xnor U15289 (N_15289,N_14107,N_14134);
nand U15290 (N_15290,N_14769,N_14156);
xor U15291 (N_15291,N_14703,N_14964);
xnor U15292 (N_15292,N_14484,N_14170);
nand U15293 (N_15293,N_14006,N_14155);
and U15294 (N_15294,N_14034,N_14188);
or U15295 (N_15295,N_13900,N_14683);
nor U15296 (N_15296,N_14431,N_14247);
or U15297 (N_15297,N_13959,N_13890);
nand U15298 (N_15298,N_14085,N_14203);
xnor U15299 (N_15299,N_14165,N_13907);
and U15300 (N_15300,N_14234,N_14081);
nor U15301 (N_15301,N_14775,N_14902);
or U15302 (N_15302,N_14305,N_14990);
nand U15303 (N_15303,N_14396,N_13934);
or U15304 (N_15304,N_14824,N_13870);
and U15305 (N_15305,N_14413,N_13859);
nor U15306 (N_15306,N_14381,N_14009);
nor U15307 (N_15307,N_14893,N_13995);
xnor U15308 (N_15308,N_14316,N_14460);
nor U15309 (N_15309,N_13921,N_13773);
nand U15310 (N_15310,N_13955,N_14755);
nand U15311 (N_15311,N_13985,N_14849);
or U15312 (N_15312,N_13807,N_13775);
and U15313 (N_15313,N_14868,N_14385);
or U15314 (N_15314,N_14987,N_14070);
xor U15315 (N_15315,N_14592,N_14449);
nor U15316 (N_15316,N_14024,N_14236);
and U15317 (N_15317,N_14878,N_14821);
nand U15318 (N_15318,N_14999,N_14018);
nand U15319 (N_15319,N_13942,N_13877);
and U15320 (N_15320,N_14819,N_14797);
and U15321 (N_15321,N_14282,N_14311);
xnor U15322 (N_15322,N_14208,N_14180);
and U15323 (N_15323,N_14326,N_14108);
or U15324 (N_15324,N_14619,N_14908);
or U15325 (N_15325,N_13818,N_14609);
xor U15326 (N_15326,N_14697,N_14796);
nand U15327 (N_15327,N_14176,N_14536);
nand U15328 (N_15328,N_13912,N_13805);
nand U15329 (N_15329,N_14158,N_14785);
xor U15330 (N_15330,N_14288,N_14383);
or U15331 (N_15331,N_14622,N_14613);
nor U15332 (N_15332,N_14787,N_14166);
nand U15333 (N_15333,N_14603,N_14198);
nand U15334 (N_15334,N_14508,N_14119);
and U15335 (N_15335,N_13794,N_14258);
nand U15336 (N_15336,N_14399,N_14095);
xnor U15337 (N_15337,N_14444,N_14663);
and U15338 (N_15338,N_14616,N_14189);
or U15339 (N_15339,N_14629,N_14190);
and U15340 (N_15340,N_13776,N_13798);
nand U15341 (N_15341,N_14195,N_14780);
nor U15342 (N_15342,N_14778,N_14746);
xnor U15343 (N_15343,N_13808,N_14145);
and U15344 (N_15344,N_14424,N_14926);
xnor U15345 (N_15345,N_14149,N_14417);
nor U15346 (N_15346,N_14369,N_14436);
or U15347 (N_15347,N_14136,N_14346);
xor U15348 (N_15348,N_14028,N_14048);
xnor U15349 (N_15349,N_14645,N_13956);
and U15350 (N_15350,N_14681,N_14066);
and U15351 (N_15351,N_13815,N_13802);
nand U15352 (N_15352,N_14567,N_14292);
or U15353 (N_15353,N_14207,N_14266);
xor U15354 (N_15354,N_14390,N_14310);
and U15355 (N_15355,N_14651,N_14816);
nor U15356 (N_15356,N_14100,N_13793);
and U15357 (N_15357,N_13918,N_14550);
nor U15358 (N_15358,N_14299,N_14969);
xor U15359 (N_15359,N_14706,N_13965);
xor U15360 (N_15360,N_14798,N_14679);
xor U15361 (N_15361,N_14434,N_13999);
xor U15362 (N_15362,N_14492,N_14161);
and U15363 (N_15363,N_14008,N_14105);
xor U15364 (N_15364,N_14382,N_14735);
xnor U15365 (N_15365,N_14923,N_13936);
or U15366 (N_15366,N_14132,N_14021);
nor U15367 (N_15367,N_14295,N_14957);
nor U15368 (N_15368,N_14549,N_14110);
nand U15369 (N_15369,N_13765,N_13996);
nor U15370 (N_15370,N_14912,N_13997);
and U15371 (N_15371,N_14857,N_14505);
or U15372 (N_15372,N_14847,N_14885);
nand U15373 (N_15373,N_14228,N_14684);
and U15374 (N_15374,N_14488,N_13780);
nor U15375 (N_15375,N_14708,N_14302);
nand U15376 (N_15376,N_14268,N_14374);
nand U15377 (N_15377,N_14732,N_14631);
or U15378 (N_15378,N_14742,N_14862);
nand U15379 (N_15379,N_13839,N_14940);
or U15380 (N_15380,N_14799,N_14178);
xnor U15381 (N_15381,N_14661,N_14644);
nor U15382 (N_15382,N_14360,N_14540);
and U15383 (N_15383,N_14972,N_14790);
xnor U15384 (N_15384,N_14313,N_14146);
or U15385 (N_15385,N_13966,N_13825);
xor U15386 (N_15386,N_13803,N_14673);
or U15387 (N_15387,N_14225,N_14186);
xnor U15388 (N_15388,N_13914,N_14768);
xor U15389 (N_15389,N_14291,N_14789);
nand U15390 (N_15390,N_14287,N_13928);
xnor U15391 (N_15391,N_14503,N_14955);
and U15392 (N_15392,N_14524,N_13875);
or U15393 (N_15393,N_14517,N_13923);
or U15394 (N_15394,N_14677,N_14162);
nor U15395 (N_15395,N_13968,N_14766);
xnor U15396 (N_15396,N_13769,N_14808);
or U15397 (N_15397,N_14252,N_14876);
xnor U15398 (N_15398,N_13950,N_14456);
and U15399 (N_15399,N_14725,N_14152);
nor U15400 (N_15400,N_14702,N_14947);
nor U15401 (N_15401,N_14366,N_14836);
nor U15402 (N_15402,N_14974,N_14997);
and U15403 (N_15403,N_14293,N_14589);
and U15404 (N_15404,N_14866,N_14455);
xor U15405 (N_15405,N_14750,N_14607);
nand U15406 (N_15406,N_14944,N_13980);
nand U15407 (N_15407,N_14200,N_14376);
or U15408 (N_15408,N_14447,N_14998);
or U15409 (N_15409,N_14950,N_14647);
xor U15410 (N_15410,N_13753,N_13862);
nand U15411 (N_15411,N_14822,N_14729);
or U15412 (N_15412,N_14805,N_14754);
and U15413 (N_15413,N_14707,N_14102);
and U15414 (N_15414,N_14127,N_14241);
nor U15415 (N_15415,N_14674,N_14482);
xnor U15416 (N_15416,N_14507,N_14029);
nor U15417 (N_15417,N_13948,N_14913);
nor U15418 (N_15418,N_14486,N_13756);
nand U15419 (N_15419,N_14978,N_14096);
nand U15420 (N_15420,N_14260,N_13871);
and U15421 (N_15421,N_13953,N_13835);
nor U15422 (N_15422,N_13916,N_14713);
or U15423 (N_15423,N_14928,N_14469);
xnor U15424 (N_15424,N_13783,N_14199);
nor U15425 (N_15425,N_14064,N_14630);
and U15426 (N_15426,N_14403,N_14653);
and U15427 (N_15427,N_14761,N_14963);
or U15428 (N_15428,N_14856,N_13836);
nor U15429 (N_15429,N_14870,N_14043);
nor U15430 (N_15430,N_14618,N_14479);
and U15431 (N_15431,N_14051,N_13823);
nand U15432 (N_15432,N_14535,N_14539);
nand U15433 (N_15433,N_14806,N_14050);
or U15434 (N_15434,N_14445,N_14038);
nor U15435 (N_15435,N_14022,N_14668);
xnor U15436 (N_15436,N_14284,N_13848);
nor U15437 (N_15437,N_14019,N_14911);
xnor U15438 (N_15438,N_13989,N_14056);
xnor U15439 (N_15439,N_14416,N_14131);
or U15440 (N_15440,N_14897,N_13933);
nand U15441 (N_15441,N_14414,N_13978);
xor U15442 (N_15442,N_14016,N_13905);
xor U15443 (N_15443,N_14652,N_14573);
or U15444 (N_15444,N_14213,N_13868);
xor U15445 (N_15445,N_13880,N_14734);
nand U15446 (N_15446,N_14074,N_13879);
xnor U15447 (N_15447,N_14709,N_13838);
xnor U15448 (N_15448,N_14634,N_14543);
nor U15449 (N_15449,N_14042,N_14770);
and U15450 (N_15450,N_14889,N_14605);
or U15451 (N_15451,N_14193,N_14509);
or U15452 (N_15452,N_13767,N_14362);
xor U15453 (N_15453,N_14375,N_14594);
nor U15454 (N_15454,N_14341,N_14628);
or U15455 (N_15455,N_14574,N_14844);
or U15456 (N_15456,N_14275,N_14183);
or U15457 (N_15457,N_14783,N_14030);
and U15458 (N_15458,N_13752,N_14525);
or U15459 (N_15459,N_14014,N_14370);
xor U15460 (N_15460,N_14518,N_14588);
nand U15461 (N_15461,N_14748,N_14468);
nor U15462 (N_15462,N_14894,N_13817);
and U15463 (N_15463,N_14680,N_14392);
nand U15464 (N_15464,N_14063,N_14344);
nand U15465 (N_15465,N_14450,N_14827);
and U15466 (N_15466,N_14076,N_13855);
nor U15467 (N_15467,N_14026,N_13951);
nor U15468 (N_15468,N_14807,N_14886);
nand U15469 (N_15469,N_14727,N_14975);
and U15470 (N_15470,N_14049,N_13979);
or U15471 (N_15471,N_13970,N_13904);
or U15472 (N_15472,N_14699,N_13843);
or U15473 (N_15473,N_14037,N_14741);
nor U15474 (N_15474,N_14075,N_14163);
nand U15475 (N_15475,N_14952,N_14654);
xnor U15476 (N_15476,N_14065,N_14516);
nand U15477 (N_15477,N_14086,N_14879);
xor U15478 (N_15478,N_13866,N_13785);
nor U15479 (N_15479,N_14451,N_14404);
or U15480 (N_15480,N_14334,N_14281);
and U15481 (N_15481,N_14993,N_13826);
or U15482 (N_15482,N_14143,N_14601);
or U15483 (N_15483,N_14041,N_14153);
xnor U15484 (N_15484,N_14328,N_13990);
nand U15485 (N_15485,N_14286,N_14496);
xnor U15486 (N_15486,N_14558,N_14461);
nand U15487 (N_15487,N_14688,N_14249);
and U15488 (N_15488,N_14753,N_13864);
nand U15489 (N_15489,N_14025,N_14932);
or U15490 (N_15490,N_14329,N_14812);
and U15491 (N_15491,N_14838,N_14235);
xnor U15492 (N_15492,N_14691,N_14823);
nor U15493 (N_15493,N_13938,N_13812);
nor U15494 (N_15494,N_13760,N_14989);
nor U15495 (N_15495,N_14297,N_14965);
xor U15496 (N_15496,N_14737,N_14280);
and U15497 (N_15497,N_14314,N_14002);
xor U15498 (N_15498,N_14515,N_14760);
nand U15499 (N_15499,N_14220,N_14526);
or U15500 (N_15500,N_14915,N_14078);
or U15501 (N_15501,N_13813,N_14745);
nor U15502 (N_15502,N_14693,N_14532);
or U15503 (N_15503,N_13988,N_14694);
or U15504 (N_15504,N_14372,N_13891);
xnor U15505 (N_15505,N_14089,N_14001);
nand U15506 (N_15506,N_14520,N_14240);
xor U15507 (N_15507,N_14415,N_14092);
xor U15508 (N_15508,N_14259,N_13981);
nand U15509 (N_15509,N_14439,N_13778);
nand U15510 (N_15510,N_14800,N_14810);
nand U15511 (N_15511,N_14229,N_14904);
nand U15512 (N_15512,N_14227,N_14617);
or U15513 (N_15513,N_13897,N_14109);
nand U15514 (N_15514,N_14784,N_14575);
nor U15515 (N_15515,N_14726,N_14958);
and U15516 (N_15516,N_14061,N_14815);
nor U15517 (N_15517,N_14336,N_14296);
nor U15518 (N_15518,N_14973,N_14804);
xor U15519 (N_15519,N_14113,N_14332);
nand U15520 (N_15520,N_14398,N_13849);
xnor U15521 (N_15521,N_14324,N_14527);
nor U15522 (N_15522,N_14570,N_14920);
xnor U15523 (N_15523,N_13755,N_14723);
xnor U15524 (N_15524,N_14802,N_14747);
nor U15525 (N_15525,N_14858,N_13751);
or U15526 (N_15526,N_14243,N_14855);
xnor U15527 (N_15527,N_14736,N_13795);
or U15528 (N_15528,N_13816,N_13847);
nand U15529 (N_15529,N_14205,N_13937);
nor U15530 (N_15530,N_13800,N_14003);
and U15531 (N_15531,N_14533,N_14231);
nor U15532 (N_15532,N_14514,N_14262);
or U15533 (N_15533,N_14949,N_14553);
or U15534 (N_15534,N_13946,N_14365);
nand U15535 (N_15535,N_14626,N_13844);
and U15536 (N_15536,N_14738,N_14406);
or U15537 (N_15537,N_14967,N_14895);
nand U15538 (N_15538,N_14554,N_14251);
or U15539 (N_15539,N_14322,N_14217);
or U15540 (N_15540,N_14731,N_13882);
and U15541 (N_15541,N_14519,N_14557);
nand U15542 (N_15542,N_14537,N_14121);
and U15543 (N_15543,N_14903,N_14465);
xnor U15544 (N_15544,N_13973,N_14082);
nand U15545 (N_15545,N_14718,N_14128);
and U15546 (N_15546,N_14773,N_13834);
xnor U15547 (N_15547,N_13917,N_14980);
xor U15548 (N_15548,N_13915,N_14223);
xnor U15549 (N_15549,N_14510,N_14779);
and U15550 (N_15550,N_13982,N_14250);
and U15551 (N_15551,N_14604,N_14387);
nor U15552 (N_15552,N_14571,N_13971);
xor U15553 (N_15553,N_14918,N_14672);
nor U15554 (N_15554,N_14995,N_14068);
or U15555 (N_15555,N_14896,N_14377);
nor U15556 (N_15556,N_14976,N_14446);
nor U15557 (N_15557,N_14196,N_14817);
and U15558 (N_15558,N_14459,N_14665);
xor U15559 (N_15559,N_13972,N_14853);
xnor U15560 (N_15560,N_14891,N_13919);
xnor U15561 (N_15561,N_14144,N_14988);
xnor U15562 (N_15562,N_14900,N_14772);
nor U15563 (N_15563,N_13964,N_14210);
nand U15564 (N_15564,N_13899,N_14587);
nand U15565 (N_15565,N_14237,N_14828);
nor U15566 (N_15566,N_13792,N_14936);
and U15567 (N_15567,N_13764,N_14960);
nand U15568 (N_15568,N_14875,N_13927);
nand U15569 (N_15569,N_14150,N_14837);
and U15570 (N_15570,N_13750,N_14538);
xor U15571 (N_15571,N_14883,N_14655);
xnor U15572 (N_15572,N_14801,N_14084);
xor U15573 (N_15573,N_13796,N_14633);
and U15574 (N_15574,N_14122,N_14117);
nand U15575 (N_15575,N_13809,N_14531);
and U15576 (N_15576,N_14485,N_13771);
nand U15577 (N_15577,N_14907,N_14992);
nand U15578 (N_15578,N_14572,N_14576);
or U15579 (N_15579,N_13954,N_14330);
or U15580 (N_15580,N_13863,N_14843);
xor U15581 (N_15581,N_14970,N_14650);
nand U15582 (N_15582,N_13876,N_13901);
nand U15583 (N_15583,N_14454,N_14319);
nor U15584 (N_15584,N_14350,N_14701);
or U15585 (N_15585,N_14032,N_14929);
or U15586 (N_15586,N_14657,N_14211);
nand U15587 (N_15587,N_14675,N_14584);
nand U15588 (N_15588,N_14814,N_13930);
and U15589 (N_15589,N_13757,N_14438);
or U15590 (N_15590,N_13784,N_14565);
nor U15591 (N_15591,N_14941,N_13992);
nor U15592 (N_15592,N_14294,N_14716);
and U15593 (N_15593,N_14033,N_14364);
or U15594 (N_15594,N_14562,N_14418);
nand U15595 (N_15595,N_14782,N_13872);
nand U15596 (N_15596,N_14354,N_14342);
nand U15597 (N_15597,N_14273,N_13898);
xor U15598 (N_15598,N_14046,N_14966);
nor U15599 (N_15599,N_13887,N_14269);
and U15600 (N_15600,N_13811,N_14272);
nor U15601 (N_15601,N_14367,N_13975);
and U15602 (N_15602,N_14649,N_14031);
or U15603 (N_15603,N_14809,N_14206);
xnor U15604 (N_15604,N_14648,N_14412);
nor U15605 (N_15605,N_14355,N_14637);
nand U15606 (N_15606,N_14338,N_13814);
or U15607 (N_15607,N_14380,N_14544);
nand U15608 (N_15608,N_14277,N_14842);
or U15609 (N_15609,N_13957,N_13908);
xor U15610 (N_15610,N_14116,N_14278);
nor U15611 (N_15611,N_14792,N_14148);
nand U15612 (N_15612,N_14013,N_14578);
nor U15613 (N_15613,N_13932,N_14712);
or U15614 (N_15614,N_14711,N_14337);
nand U15615 (N_15615,N_14871,N_14393);
nor U15616 (N_15616,N_14846,N_14202);
and U15617 (N_15617,N_14440,N_14522);
nand U15618 (N_15618,N_14818,N_13824);
xor U15619 (N_15619,N_13958,N_14662);
xor U15620 (N_15620,N_14473,N_14098);
nand U15621 (N_15621,N_13878,N_14091);
or U15622 (N_15622,N_13889,N_13974);
or U15623 (N_15623,N_14265,N_14352);
and U15624 (N_15624,N_14349,N_14129);
nand U15625 (N_15625,N_14754,N_14614);
nor U15626 (N_15626,N_14551,N_13987);
or U15627 (N_15627,N_14725,N_13949);
nand U15628 (N_15628,N_14456,N_14415);
xor U15629 (N_15629,N_14072,N_14838);
or U15630 (N_15630,N_14461,N_14418);
or U15631 (N_15631,N_14375,N_13953);
and U15632 (N_15632,N_14201,N_14872);
nor U15633 (N_15633,N_14233,N_14934);
xor U15634 (N_15634,N_14740,N_14633);
nand U15635 (N_15635,N_13999,N_13879);
nor U15636 (N_15636,N_14597,N_14309);
and U15637 (N_15637,N_14384,N_14750);
xor U15638 (N_15638,N_14297,N_14617);
nand U15639 (N_15639,N_14988,N_14327);
nor U15640 (N_15640,N_14412,N_14706);
nor U15641 (N_15641,N_14503,N_14590);
xor U15642 (N_15642,N_14619,N_14630);
and U15643 (N_15643,N_13776,N_14096);
or U15644 (N_15644,N_14814,N_14656);
xor U15645 (N_15645,N_14383,N_14502);
xnor U15646 (N_15646,N_14190,N_14073);
nand U15647 (N_15647,N_13925,N_14855);
and U15648 (N_15648,N_13916,N_14225);
or U15649 (N_15649,N_14328,N_13769);
nor U15650 (N_15650,N_14229,N_14735);
or U15651 (N_15651,N_14623,N_13838);
and U15652 (N_15652,N_14279,N_14440);
and U15653 (N_15653,N_14075,N_14231);
and U15654 (N_15654,N_14878,N_13765);
xnor U15655 (N_15655,N_13898,N_14381);
and U15656 (N_15656,N_14653,N_14637);
nand U15657 (N_15657,N_14968,N_14777);
and U15658 (N_15658,N_14440,N_14232);
and U15659 (N_15659,N_14523,N_14053);
or U15660 (N_15660,N_14465,N_14899);
and U15661 (N_15661,N_14229,N_14305);
xnor U15662 (N_15662,N_14525,N_14635);
nand U15663 (N_15663,N_13974,N_13849);
xnor U15664 (N_15664,N_13777,N_13938);
or U15665 (N_15665,N_14324,N_14311);
nor U15666 (N_15666,N_14150,N_14798);
xor U15667 (N_15667,N_14106,N_14880);
or U15668 (N_15668,N_14006,N_13792);
and U15669 (N_15669,N_14001,N_14724);
and U15670 (N_15670,N_13796,N_14654);
nand U15671 (N_15671,N_14404,N_14641);
nor U15672 (N_15672,N_13783,N_14974);
nor U15673 (N_15673,N_13992,N_14297);
nand U15674 (N_15674,N_14743,N_14359);
and U15675 (N_15675,N_14560,N_14224);
and U15676 (N_15676,N_13970,N_14667);
and U15677 (N_15677,N_14215,N_14755);
and U15678 (N_15678,N_14740,N_14194);
nor U15679 (N_15679,N_13880,N_14321);
xnor U15680 (N_15680,N_14402,N_14577);
or U15681 (N_15681,N_14436,N_14695);
nand U15682 (N_15682,N_14889,N_14092);
xnor U15683 (N_15683,N_14846,N_14891);
nor U15684 (N_15684,N_14055,N_13916);
nand U15685 (N_15685,N_14219,N_14394);
nor U15686 (N_15686,N_14893,N_14565);
nand U15687 (N_15687,N_14851,N_13821);
and U15688 (N_15688,N_14798,N_14517);
or U15689 (N_15689,N_14964,N_14652);
nor U15690 (N_15690,N_14601,N_14852);
nor U15691 (N_15691,N_14626,N_14258);
xnor U15692 (N_15692,N_14951,N_14111);
nand U15693 (N_15693,N_14008,N_14412);
nor U15694 (N_15694,N_13928,N_14930);
nand U15695 (N_15695,N_14022,N_14106);
nand U15696 (N_15696,N_14873,N_14741);
nor U15697 (N_15697,N_14590,N_14946);
nor U15698 (N_15698,N_13889,N_14145);
nand U15699 (N_15699,N_14163,N_14695);
and U15700 (N_15700,N_14079,N_14920);
or U15701 (N_15701,N_14776,N_14574);
or U15702 (N_15702,N_14830,N_14384);
and U15703 (N_15703,N_14412,N_14792);
xnor U15704 (N_15704,N_14211,N_14301);
nor U15705 (N_15705,N_14868,N_13957);
or U15706 (N_15706,N_14177,N_14108);
or U15707 (N_15707,N_14549,N_14514);
nand U15708 (N_15708,N_14823,N_14379);
nor U15709 (N_15709,N_14008,N_14812);
xnor U15710 (N_15710,N_14459,N_14119);
nor U15711 (N_15711,N_14265,N_14221);
or U15712 (N_15712,N_14752,N_14545);
or U15713 (N_15713,N_14588,N_14894);
nor U15714 (N_15714,N_13772,N_14124);
nor U15715 (N_15715,N_14486,N_14922);
xnor U15716 (N_15716,N_14669,N_14738);
and U15717 (N_15717,N_14342,N_13768);
nand U15718 (N_15718,N_14219,N_14087);
or U15719 (N_15719,N_14816,N_14795);
nand U15720 (N_15720,N_14574,N_14806);
nor U15721 (N_15721,N_14014,N_14353);
nand U15722 (N_15722,N_14633,N_14778);
and U15723 (N_15723,N_14245,N_14266);
or U15724 (N_15724,N_14387,N_13970);
nand U15725 (N_15725,N_13791,N_13776);
and U15726 (N_15726,N_13838,N_14216);
xnor U15727 (N_15727,N_14834,N_14761);
and U15728 (N_15728,N_14462,N_14746);
nand U15729 (N_15729,N_14615,N_14382);
and U15730 (N_15730,N_14533,N_14121);
nor U15731 (N_15731,N_14226,N_14230);
and U15732 (N_15732,N_14666,N_14451);
nand U15733 (N_15733,N_14822,N_14545);
and U15734 (N_15734,N_14687,N_13899);
and U15735 (N_15735,N_14647,N_14396);
xnor U15736 (N_15736,N_13852,N_14046);
nand U15737 (N_15737,N_14002,N_14114);
nand U15738 (N_15738,N_14212,N_14147);
or U15739 (N_15739,N_14624,N_13926);
or U15740 (N_15740,N_14612,N_14718);
nand U15741 (N_15741,N_13814,N_14584);
and U15742 (N_15742,N_14210,N_13889);
nor U15743 (N_15743,N_14104,N_14276);
xnor U15744 (N_15744,N_14510,N_14731);
nand U15745 (N_15745,N_14988,N_14697);
xor U15746 (N_15746,N_14658,N_14140);
xor U15747 (N_15747,N_14234,N_14897);
and U15748 (N_15748,N_14349,N_14669);
and U15749 (N_15749,N_14302,N_14352);
or U15750 (N_15750,N_14569,N_14502);
or U15751 (N_15751,N_14397,N_13828);
or U15752 (N_15752,N_14022,N_14706);
xnor U15753 (N_15753,N_14887,N_14180);
nand U15754 (N_15754,N_14426,N_14788);
or U15755 (N_15755,N_14289,N_14968);
and U15756 (N_15756,N_14557,N_14124);
or U15757 (N_15757,N_14019,N_14547);
nand U15758 (N_15758,N_14927,N_14512);
and U15759 (N_15759,N_14115,N_14127);
xnor U15760 (N_15760,N_13903,N_13818);
or U15761 (N_15761,N_14019,N_14606);
and U15762 (N_15762,N_14599,N_14460);
xor U15763 (N_15763,N_14933,N_14919);
nand U15764 (N_15764,N_13973,N_14767);
and U15765 (N_15765,N_14872,N_13758);
and U15766 (N_15766,N_14849,N_14612);
or U15767 (N_15767,N_14371,N_14638);
and U15768 (N_15768,N_14364,N_14587);
nor U15769 (N_15769,N_14371,N_14425);
nor U15770 (N_15770,N_14405,N_13862);
nor U15771 (N_15771,N_13969,N_14794);
nor U15772 (N_15772,N_13994,N_14633);
or U15773 (N_15773,N_13803,N_14759);
nor U15774 (N_15774,N_13762,N_13780);
or U15775 (N_15775,N_14350,N_14208);
nand U15776 (N_15776,N_14196,N_14131);
nand U15777 (N_15777,N_14094,N_14452);
xnor U15778 (N_15778,N_14387,N_14877);
and U15779 (N_15779,N_14618,N_14519);
and U15780 (N_15780,N_14145,N_14901);
or U15781 (N_15781,N_13773,N_14407);
or U15782 (N_15782,N_13987,N_14587);
nor U15783 (N_15783,N_14959,N_13852);
xnor U15784 (N_15784,N_13869,N_13804);
nand U15785 (N_15785,N_13936,N_14228);
and U15786 (N_15786,N_14547,N_14683);
or U15787 (N_15787,N_14174,N_14838);
or U15788 (N_15788,N_13873,N_14828);
nand U15789 (N_15789,N_14728,N_14532);
xnor U15790 (N_15790,N_14295,N_14394);
xor U15791 (N_15791,N_14189,N_14885);
nand U15792 (N_15792,N_14789,N_14086);
nand U15793 (N_15793,N_13858,N_14310);
or U15794 (N_15794,N_14057,N_14720);
nand U15795 (N_15795,N_14989,N_14721);
nand U15796 (N_15796,N_14592,N_13943);
and U15797 (N_15797,N_14924,N_14181);
and U15798 (N_15798,N_13962,N_14826);
nor U15799 (N_15799,N_13753,N_14587);
nor U15800 (N_15800,N_14738,N_14944);
nor U15801 (N_15801,N_14996,N_14156);
nand U15802 (N_15802,N_14267,N_13836);
xnor U15803 (N_15803,N_13850,N_14618);
or U15804 (N_15804,N_14099,N_14536);
nor U15805 (N_15805,N_13830,N_14557);
nand U15806 (N_15806,N_14430,N_14399);
and U15807 (N_15807,N_14812,N_14612);
and U15808 (N_15808,N_14673,N_14360);
and U15809 (N_15809,N_14849,N_13787);
nor U15810 (N_15810,N_13839,N_14594);
and U15811 (N_15811,N_14027,N_14552);
and U15812 (N_15812,N_14440,N_14717);
and U15813 (N_15813,N_13892,N_14046);
nand U15814 (N_15814,N_14078,N_14953);
or U15815 (N_15815,N_14157,N_14951);
nor U15816 (N_15816,N_14420,N_14589);
nand U15817 (N_15817,N_13768,N_14487);
nand U15818 (N_15818,N_14018,N_14144);
xnor U15819 (N_15819,N_14708,N_14710);
and U15820 (N_15820,N_14906,N_13800);
nor U15821 (N_15821,N_14743,N_14648);
nand U15822 (N_15822,N_14549,N_13780);
nand U15823 (N_15823,N_14844,N_14596);
nand U15824 (N_15824,N_14706,N_13842);
or U15825 (N_15825,N_13910,N_14782);
nand U15826 (N_15826,N_14223,N_14314);
and U15827 (N_15827,N_14725,N_14833);
nand U15828 (N_15828,N_14152,N_14679);
and U15829 (N_15829,N_14756,N_14724);
and U15830 (N_15830,N_14364,N_14188);
and U15831 (N_15831,N_14550,N_13826);
nand U15832 (N_15832,N_14870,N_14346);
nor U15833 (N_15833,N_14350,N_14964);
and U15834 (N_15834,N_13854,N_14597);
and U15835 (N_15835,N_14883,N_14075);
or U15836 (N_15836,N_14940,N_14417);
and U15837 (N_15837,N_13794,N_14030);
nand U15838 (N_15838,N_14503,N_14674);
and U15839 (N_15839,N_14179,N_14722);
or U15840 (N_15840,N_14912,N_14390);
or U15841 (N_15841,N_14339,N_14927);
nor U15842 (N_15842,N_14204,N_14652);
or U15843 (N_15843,N_14548,N_14819);
and U15844 (N_15844,N_14242,N_14536);
or U15845 (N_15845,N_14055,N_14378);
xnor U15846 (N_15846,N_14782,N_14324);
nor U15847 (N_15847,N_14559,N_13940);
xor U15848 (N_15848,N_13781,N_14507);
or U15849 (N_15849,N_14359,N_14691);
or U15850 (N_15850,N_14632,N_13896);
nor U15851 (N_15851,N_14271,N_14657);
or U15852 (N_15852,N_14461,N_14976);
nand U15853 (N_15853,N_14806,N_13980);
nor U15854 (N_15854,N_13782,N_13809);
and U15855 (N_15855,N_14433,N_14499);
nor U15856 (N_15856,N_14021,N_13849);
nand U15857 (N_15857,N_14762,N_14016);
xor U15858 (N_15858,N_14944,N_14428);
nand U15859 (N_15859,N_13997,N_14364);
nand U15860 (N_15860,N_13917,N_14694);
nand U15861 (N_15861,N_13811,N_14785);
nor U15862 (N_15862,N_14066,N_13900);
nor U15863 (N_15863,N_14868,N_13849);
nor U15864 (N_15864,N_14378,N_14074);
or U15865 (N_15865,N_14132,N_14820);
nor U15866 (N_15866,N_13881,N_14943);
nand U15867 (N_15867,N_14739,N_14560);
or U15868 (N_15868,N_13940,N_14700);
xnor U15869 (N_15869,N_14537,N_13792);
nand U15870 (N_15870,N_14682,N_14618);
or U15871 (N_15871,N_13840,N_14917);
nand U15872 (N_15872,N_13868,N_14932);
and U15873 (N_15873,N_14528,N_14933);
and U15874 (N_15874,N_14020,N_14055);
nor U15875 (N_15875,N_14399,N_13914);
or U15876 (N_15876,N_14459,N_13926);
or U15877 (N_15877,N_14272,N_14764);
and U15878 (N_15878,N_14906,N_14244);
or U15879 (N_15879,N_13822,N_14094);
nand U15880 (N_15880,N_14298,N_14386);
nand U15881 (N_15881,N_14215,N_14739);
nor U15882 (N_15882,N_14124,N_14852);
nand U15883 (N_15883,N_13801,N_13785);
xor U15884 (N_15884,N_14069,N_14784);
nand U15885 (N_15885,N_14089,N_14103);
nor U15886 (N_15886,N_14160,N_13841);
xnor U15887 (N_15887,N_14219,N_14919);
or U15888 (N_15888,N_13993,N_14208);
xor U15889 (N_15889,N_14842,N_14496);
nor U15890 (N_15890,N_14547,N_14014);
or U15891 (N_15891,N_14549,N_14860);
or U15892 (N_15892,N_14930,N_13785);
nor U15893 (N_15893,N_13861,N_14339);
xnor U15894 (N_15894,N_14658,N_14032);
and U15895 (N_15895,N_13974,N_14293);
and U15896 (N_15896,N_14665,N_14111);
and U15897 (N_15897,N_14253,N_14114);
and U15898 (N_15898,N_14550,N_13957);
or U15899 (N_15899,N_14154,N_14338);
xnor U15900 (N_15900,N_14779,N_14047);
nor U15901 (N_15901,N_14588,N_14768);
or U15902 (N_15902,N_14417,N_13858);
xnor U15903 (N_15903,N_13940,N_14984);
or U15904 (N_15904,N_14584,N_14040);
nand U15905 (N_15905,N_13756,N_14585);
and U15906 (N_15906,N_14775,N_14208);
and U15907 (N_15907,N_13863,N_13949);
xor U15908 (N_15908,N_14025,N_14718);
or U15909 (N_15909,N_14361,N_13880);
nand U15910 (N_15910,N_14923,N_14900);
nor U15911 (N_15911,N_14489,N_14171);
xnor U15912 (N_15912,N_14929,N_14302);
xor U15913 (N_15913,N_14548,N_14081);
nor U15914 (N_15914,N_14535,N_14449);
xor U15915 (N_15915,N_14739,N_14869);
and U15916 (N_15916,N_14881,N_14346);
xnor U15917 (N_15917,N_13921,N_14897);
or U15918 (N_15918,N_14003,N_14897);
nand U15919 (N_15919,N_14394,N_14584);
nand U15920 (N_15920,N_14847,N_13895);
nor U15921 (N_15921,N_14246,N_14018);
and U15922 (N_15922,N_14547,N_14498);
nor U15923 (N_15923,N_14810,N_14189);
and U15924 (N_15924,N_14777,N_13871);
or U15925 (N_15925,N_13911,N_13766);
and U15926 (N_15926,N_14772,N_14871);
xnor U15927 (N_15927,N_14462,N_13889);
or U15928 (N_15928,N_13940,N_14238);
or U15929 (N_15929,N_13842,N_14204);
xor U15930 (N_15930,N_14860,N_13840);
nor U15931 (N_15931,N_14948,N_14078);
and U15932 (N_15932,N_14211,N_14542);
nor U15933 (N_15933,N_14529,N_14803);
nand U15934 (N_15934,N_14478,N_13850);
nor U15935 (N_15935,N_14378,N_14659);
xnor U15936 (N_15936,N_14130,N_14507);
or U15937 (N_15937,N_14238,N_14027);
nor U15938 (N_15938,N_13762,N_14788);
nand U15939 (N_15939,N_13778,N_14102);
xnor U15940 (N_15940,N_14956,N_14250);
xor U15941 (N_15941,N_14671,N_14401);
nand U15942 (N_15942,N_14592,N_13887);
nand U15943 (N_15943,N_14067,N_14836);
or U15944 (N_15944,N_13967,N_14299);
nand U15945 (N_15945,N_13996,N_14919);
nand U15946 (N_15946,N_14084,N_14636);
and U15947 (N_15947,N_13774,N_14675);
nor U15948 (N_15948,N_14907,N_14561);
and U15949 (N_15949,N_14068,N_14679);
nor U15950 (N_15950,N_14435,N_14695);
nand U15951 (N_15951,N_14419,N_14367);
nand U15952 (N_15952,N_14137,N_14179);
or U15953 (N_15953,N_14236,N_14368);
nand U15954 (N_15954,N_14605,N_14514);
and U15955 (N_15955,N_14065,N_14130);
and U15956 (N_15956,N_13921,N_14915);
and U15957 (N_15957,N_14169,N_14997);
xnor U15958 (N_15958,N_14390,N_14794);
xor U15959 (N_15959,N_14032,N_14624);
xnor U15960 (N_15960,N_14283,N_13860);
and U15961 (N_15961,N_14143,N_14045);
xnor U15962 (N_15962,N_14177,N_13943);
nor U15963 (N_15963,N_13977,N_14989);
nand U15964 (N_15964,N_14077,N_14457);
nor U15965 (N_15965,N_14894,N_14746);
xnor U15966 (N_15966,N_14072,N_14999);
or U15967 (N_15967,N_13805,N_14659);
nor U15968 (N_15968,N_14301,N_13964);
nor U15969 (N_15969,N_13894,N_14356);
xnor U15970 (N_15970,N_14612,N_13787);
or U15971 (N_15971,N_14981,N_13928);
or U15972 (N_15972,N_13847,N_13786);
nor U15973 (N_15973,N_14256,N_14079);
xor U15974 (N_15974,N_14919,N_14346);
and U15975 (N_15975,N_14002,N_13901);
xnor U15976 (N_15976,N_14120,N_14863);
or U15977 (N_15977,N_14931,N_14319);
and U15978 (N_15978,N_14567,N_14817);
nor U15979 (N_15979,N_14826,N_14772);
or U15980 (N_15980,N_13791,N_14407);
or U15981 (N_15981,N_13947,N_13982);
xor U15982 (N_15982,N_14430,N_13814);
or U15983 (N_15983,N_14165,N_14170);
or U15984 (N_15984,N_13902,N_13880);
nand U15985 (N_15985,N_13766,N_13894);
and U15986 (N_15986,N_14141,N_14565);
xnor U15987 (N_15987,N_13986,N_14527);
and U15988 (N_15988,N_14700,N_14431);
nor U15989 (N_15989,N_14244,N_13996);
or U15990 (N_15990,N_14709,N_14500);
nor U15991 (N_15991,N_14694,N_14939);
nand U15992 (N_15992,N_14876,N_14123);
or U15993 (N_15993,N_14094,N_14555);
or U15994 (N_15994,N_14463,N_14184);
nand U15995 (N_15995,N_13845,N_14917);
and U15996 (N_15996,N_13964,N_14215);
nand U15997 (N_15997,N_14304,N_14235);
or U15998 (N_15998,N_14804,N_14884);
and U15999 (N_15999,N_14581,N_14750);
and U16000 (N_16000,N_14170,N_13769);
nand U16001 (N_16001,N_14174,N_14636);
nor U16002 (N_16002,N_14329,N_14392);
and U16003 (N_16003,N_14156,N_13804);
or U16004 (N_16004,N_13920,N_14038);
or U16005 (N_16005,N_14719,N_14619);
nor U16006 (N_16006,N_14402,N_14241);
nor U16007 (N_16007,N_14833,N_14826);
nor U16008 (N_16008,N_13938,N_13886);
xnor U16009 (N_16009,N_14687,N_14528);
or U16010 (N_16010,N_14069,N_14715);
and U16011 (N_16011,N_13880,N_13879);
nor U16012 (N_16012,N_14019,N_14685);
xor U16013 (N_16013,N_14204,N_14969);
nor U16014 (N_16014,N_14998,N_14042);
and U16015 (N_16015,N_14611,N_14979);
nor U16016 (N_16016,N_14297,N_14103);
and U16017 (N_16017,N_13830,N_14277);
and U16018 (N_16018,N_14426,N_14172);
and U16019 (N_16019,N_14093,N_14914);
nor U16020 (N_16020,N_14339,N_14673);
and U16021 (N_16021,N_14473,N_14486);
nor U16022 (N_16022,N_14603,N_14568);
xor U16023 (N_16023,N_14828,N_14219);
nand U16024 (N_16024,N_14205,N_14537);
and U16025 (N_16025,N_14871,N_13954);
and U16026 (N_16026,N_13841,N_14650);
and U16027 (N_16027,N_13781,N_14455);
and U16028 (N_16028,N_14299,N_14690);
nand U16029 (N_16029,N_14345,N_13866);
nor U16030 (N_16030,N_14055,N_14534);
xor U16031 (N_16031,N_14718,N_14091);
nor U16032 (N_16032,N_13951,N_14433);
nor U16033 (N_16033,N_14930,N_14031);
nor U16034 (N_16034,N_14585,N_14522);
nor U16035 (N_16035,N_14059,N_13990);
and U16036 (N_16036,N_14262,N_14165);
xnor U16037 (N_16037,N_14427,N_14729);
nand U16038 (N_16038,N_14249,N_14997);
and U16039 (N_16039,N_14922,N_14527);
and U16040 (N_16040,N_14230,N_14727);
xnor U16041 (N_16041,N_14007,N_14433);
or U16042 (N_16042,N_14592,N_14271);
nand U16043 (N_16043,N_13970,N_13780);
and U16044 (N_16044,N_14091,N_14316);
and U16045 (N_16045,N_13990,N_14359);
and U16046 (N_16046,N_13943,N_14748);
nor U16047 (N_16047,N_13944,N_13785);
or U16048 (N_16048,N_14755,N_14244);
or U16049 (N_16049,N_14112,N_14942);
nor U16050 (N_16050,N_14238,N_14630);
and U16051 (N_16051,N_14337,N_14930);
nand U16052 (N_16052,N_14100,N_13837);
or U16053 (N_16053,N_14443,N_14018);
nand U16054 (N_16054,N_14694,N_14593);
or U16055 (N_16055,N_14827,N_14497);
or U16056 (N_16056,N_13838,N_14893);
nand U16057 (N_16057,N_13967,N_14054);
or U16058 (N_16058,N_14338,N_14326);
or U16059 (N_16059,N_14048,N_14692);
or U16060 (N_16060,N_14329,N_14612);
nand U16061 (N_16061,N_13910,N_13824);
xnor U16062 (N_16062,N_13841,N_14272);
and U16063 (N_16063,N_14466,N_13992);
nand U16064 (N_16064,N_13769,N_14023);
and U16065 (N_16065,N_14988,N_14505);
and U16066 (N_16066,N_14693,N_14454);
and U16067 (N_16067,N_14062,N_14349);
and U16068 (N_16068,N_13858,N_14730);
and U16069 (N_16069,N_14966,N_14100);
and U16070 (N_16070,N_13968,N_13959);
nand U16071 (N_16071,N_14558,N_14377);
and U16072 (N_16072,N_14105,N_14863);
or U16073 (N_16073,N_14321,N_13838);
and U16074 (N_16074,N_14509,N_14899);
xnor U16075 (N_16075,N_14276,N_14418);
and U16076 (N_16076,N_14139,N_14592);
nand U16077 (N_16077,N_14510,N_14801);
and U16078 (N_16078,N_14644,N_14217);
and U16079 (N_16079,N_14234,N_14374);
xnor U16080 (N_16080,N_13949,N_14047);
xnor U16081 (N_16081,N_14318,N_14627);
xor U16082 (N_16082,N_14351,N_14546);
xor U16083 (N_16083,N_14937,N_14682);
nor U16084 (N_16084,N_14547,N_14449);
nor U16085 (N_16085,N_14088,N_14961);
nor U16086 (N_16086,N_14415,N_14801);
nand U16087 (N_16087,N_14273,N_14799);
nor U16088 (N_16088,N_14885,N_13865);
nand U16089 (N_16089,N_14990,N_14862);
and U16090 (N_16090,N_14091,N_13847);
nand U16091 (N_16091,N_14384,N_14886);
and U16092 (N_16092,N_14479,N_14281);
xnor U16093 (N_16093,N_13883,N_13948);
and U16094 (N_16094,N_14551,N_14939);
nand U16095 (N_16095,N_13875,N_14339);
and U16096 (N_16096,N_13775,N_14182);
xnor U16097 (N_16097,N_13876,N_14074);
nand U16098 (N_16098,N_13776,N_14361);
xnor U16099 (N_16099,N_14256,N_13847);
and U16100 (N_16100,N_14335,N_14380);
nor U16101 (N_16101,N_14821,N_14592);
nand U16102 (N_16102,N_14777,N_14752);
nor U16103 (N_16103,N_14044,N_13964);
and U16104 (N_16104,N_13895,N_13911);
nor U16105 (N_16105,N_14643,N_14835);
nand U16106 (N_16106,N_13866,N_14541);
nor U16107 (N_16107,N_14103,N_14806);
nand U16108 (N_16108,N_14366,N_13852);
nand U16109 (N_16109,N_14385,N_14751);
and U16110 (N_16110,N_13914,N_14572);
xnor U16111 (N_16111,N_13755,N_14349);
nor U16112 (N_16112,N_14452,N_13909);
xnor U16113 (N_16113,N_14487,N_14041);
nor U16114 (N_16114,N_14561,N_14247);
nor U16115 (N_16115,N_14607,N_14071);
or U16116 (N_16116,N_13885,N_14316);
and U16117 (N_16117,N_14152,N_13885);
and U16118 (N_16118,N_14928,N_13809);
nand U16119 (N_16119,N_14228,N_14475);
nand U16120 (N_16120,N_14265,N_14372);
nand U16121 (N_16121,N_14527,N_14997);
xnor U16122 (N_16122,N_14696,N_13794);
xor U16123 (N_16123,N_14805,N_13807);
nand U16124 (N_16124,N_14024,N_14536);
xor U16125 (N_16125,N_14054,N_14639);
nor U16126 (N_16126,N_14452,N_14253);
and U16127 (N_16127,N_14736,N_14819);
or U16128 (N_16128,N_14048,N_14064);
or U16129 (N_16129,N_13902,N_14693);
and U16130 (N_16130,N_14245,N_14382);
xnor U16131 (N_16131,N_14634,N_13775);
xnor U16132 (N_16132,N_14884,N_14561);
nand U16133 (N_16133,N_14712,N_14647);
and U16134 (N_16134,N_14775,N_14083);
nand U16135 (N_16135,N_14813,N_14448);
nand U16136 (N_16136,N_14202,N_14753);
xor U16137 (N_16137,N_13938,N_14223);
or U16138 (N_16138,N_13857,N_14214);
nor U16139 (N_16139,N_13967,N_14690);
nand U16140 (N_16140,N_14575,N_14750);
xor U16141 (N_16141,N_13767,N_14470);
nor U16142 (N_16142,N_14193,N_14692);
and U16143 (N_16143,N_14323,N_13775);
or U16144 (N_16144,N_14160,N_14397);
xnor U16145 (N_16145,N_14786,N_14889);
xnor U16146 (N_16146,N_14360,N_14650);
or U16147 (N_16147,N_13892,N_13829);
nor U16148 (N_16148,N_14433,N_14205);
xor U16149 (N_16149,N_14039,N_14545);
nor U16150 (N_16150,N_14607,N_14568);
or U16151 (N_16151,N_13942,N_14148);
or U16152 (N_16152,N_13929,N_13793);
and U16153 (N_16153,N_14374,N_14175);
nor U16154 (N_16154,N_14066,N_13960);
and U16155 (N_16155,N_14244,N_14700);
or U16156 (N_16156,N_13756,N_14736);
nand U16157 (N_16157,N_14143,N_14653);
xor U16158 (N_16158,N_14833,N_13855);
nand U16159 (N_16159,N_14875,N_14595);
or U16160 (N_16160,N_13995,N_13773);
nor U16161 (N_16161,N_14105,N_14244);
or U16162 (N_16162,N_14571,N_14140);
and U16163 (N_16163,N_14557,N_14695);
xor U16164 (N_16164,N_13851,N_14880);
nand U16165 (N_16165,N_13820,N_14535);
xor U16166 (N_16166,N_14085,N_13928);
or U16167 (N_16167,N_14426,N_14650);
and U16168 (N_16168,N_14765,N_14792);
or U16169 (N_16169,N_14090,N_14899);
or U16170 (N_16170,N_13886,N_14137);
nor U16171 (N_16171,N_14170,N_13872);
nor U16172 (N_16172,N_13950,N_14105);
or U16173 (N_16173,N_14942,N_14623);
nor U16174 (N_16174,N_14329,N_14595);
and U16175 (N_16175,N_14820,N_13898);
xor U16176 (N_16176,N_14804,N_14708);
nor U16177 (N_16177,N_14087,N_14533);
and U16178 (N_16178,N_14362,N_13841);
nand U16179 (N_16179,N_14674,N_14877);
and U16180 (N_16180,N_14472,N_13824);
and U16181 (N_16181,N_14662,N_14709);
nor U16182 (N_16182,N_14573,N_14642);
or U16183 (N_16183,N_14834,N_13987);
xnor U16184 (N_16184,N_14349,N_14184);
nor U16185 (N_16185,N_14286,N_14187);
nand U16186 (N_16186,N_13924,N_14976);
nand U16187 (N_16187,N_14389,N_14970);
xnor U16188 (N_16188,N_14865,N_14349);
nor U16189 (N_16189,N_14037,N_13811);
and U16190 (N_16190,N_14638,N_14453);
nand U16191 (N_16191,N_14342,N_14918);
xnor U16192 (N_16192,N_14612,N_14121);
xnor U16193 (N_16193,N_14016,N_14165);
nand U16194 (N_16194,N_14432,N_13896);
or U16195 (N_16195,N_14237,N_14163);
xor U16196 (N_16196,N_13770,N_14680);
or U16197 (N_16197,N_14594,N_14366);
or U16198 (N_16198,N_13869,N_14338);
nor U16199 (N_16199,N_14715,N_14766);
nor U16200 (N_16200,N_14899,N_14361);
xnor U16201 (N_16201,N_14868,N_14998);
or U16202 (N_16202,N_14467,N_14090);
xor U16203 (N_16203,N_13793,N_14073);
nand U16204 (N_16204,N_13854,N_14938);
and U16205 (N_16205,N_14001,N_14657);
or U16206 (N_16206,N_14643,N_14004);
or U16207 (N_16207,N_14136,N_14776);
or U16208 (N_16208,N_14082,N_14339);
nand U16209 (N_16209,N_14777,N_14334);
nor U16210 (N_16210,N_14322,N_14627);
nor U16211 (N_16211,N_14326,N_14646);
nand U16212 (N_16212,N_14961,N_14425);
or U16213 (N_16213,N_13874,N_14731);
nor U16214 (N_16214,N_14830,N_14808);
xor U16215 (N_16215,N_14323,N_14585);
or U16216 (N_16216,N_14234,N_13820);
or U16217 (N_16217,N_14811,N_14792);
or U16218 (N_16218,N_14676,N_13899);
xnor U16219 (N_16219,N_14430,N_14601);
nand U16220 (N_16220,N_14004,N_14140);
nor U16221 (N_16221,N_14341,N_14814);
or U16222 (N_16222,N_14306,N_14267);
and U16223 (N_16223,N_14189,N_14530);
nor U16224 (N_16224,N_13824,N_14942);
xnor U16225 (N_16225,N_14139,N_14622);
nand U16226 (N_16226,N_14004,N_14283);
nor U16227 (N_16227,N_14305,N_14058);
nor U16228 (N_16228,N_14593,N_13809);
and U16229 (N_16229,N_13807,N_14395);
or U16230 (N_16230,N_13864,N_14789);
xnor U16231 (N_16231,N_14996,N_13818);
or U16232 (N_16232,N_13758,N_14524);
and U16233 (N_16233,N_14003,N_14498);
xor U16234 (N_16234,N_14166,N_14508);
xnor U16235 (N_16235,N_13895,N_14194);
or U16236 (N_16236,N_13928,N_13897);
nand U16237 (N_16237,N_13944,N_14201);
and U16238 (N_16238,N_14750,N_14703);
and U16239 (N_16239,N_14005,N_14804);
nor U16240 (N_16240,N_14873,N_14822);
xnor U16241 (N_16241,N_14897,N_14102);
xor U16242 (N_16242,N_14400,N_14418);
nor U16243 (N_16243,N_13750,N_13996);
and U16244 (N_16244,N_14416,N_14792);
and U16245 (N_16245,N_14730,N_13879);
nor U16246 (N_16246,N_13809,N_14731);
xnor U16247 (N_16247,N_13823,N_14841);
nor U16248 (N_16248,N_14349,N_14532);
or U16249 (N_16249,N_14496,N_14832);
nor U16250 (N_16250,N_15852,N_16195);
nand U16251 (N_16251,N_15323,N_16008);
nor U16252 (N_16252,N_15639,N_15511);
nand U16253 (N_16253,N_15370,N_15487);
or U16254 (N_16254,N_15339,N_16226);
and U16255 (N_16255,N_15754,N_16200);
nor U16256 (N_16256,N_15427,N_15608);
xnor U16257 (N_16257,N_16207,N_16243);
nand U16258 (N_16258,N_15766,N_16208);
or U16259 (N_16259,N_15879,N_15127);
xnor U16260 (N_16260,N_16031,N_16040);
and U16261 (N_16261,N_15501,N_15731);
nand U16262 (N_16262,N_15738,N_15818);
and U16263 (N_16263,N_15165,N_15168);
xor U16264 (N_16264,N_16189,N_15552);
nor U16265 (N_16265,N_15000,N_15118);
nor U16266 (N_16266,N_15987,N_15609);
and U16267 (N_16267,N_15260,N_15214);
or U16268 (N_16268,N_16073,N_15983);
nand U16269 (N_16269,N_15962,N_15304);
nand U16270 (N_16270,N_15992,N_15549);
xnor U16271 (N_16271,N_15030,N_15712);
or U16272 (N_16272,N_15177,N_16131);
nor U16273 (N_16273,N_15756,N_15869);
nor U16274 (N_16274,N_16017,N_15572);
xnor U16275 (N_16275,N_15972,N_15775);
xor U16276 (N_16276,N_15056,N_15574);
nor U16277 (N_16277,N_16196,N_15587);
xor U16278 (N_16278,N_15167,N_16053);
xnor U16279 (N_16279,N_15788,N_16234);
or U16280 (N_16280,N_15259,N_15548);
nor U16281 (N_16281,N_16174,N_15790);
and U16282 (N_16282,N_15443,N_15313);
nor U16283 (N_16283,N_15789,N_15029);
nand U16284 (N_16284,N_15543,N_15134);
nor U16285 (N_16285,N_15054,N_15402);
and U16286 (N_16286,N_15171,N_15507);
xnor U16287 (N_16287,N_16068,N_15346);
and U16288 (N_16288,N_16125,N_16016);
xnor U16289 (N_16289,N_15556,N_15349);
nor U16290 (N_16290,N_15568,N_15036);
or U16291 (N_16291,N_16223,N_15090);
xor U16292 (N_16292,N_15931,N_15272);
and U16293 (N_16293,N_15045,N_15954);
or U16294 (N_16294,N_15482,N_16020);
and U16295 (N_16295,N_16218,N_15286);
xnor U16296 (N_16296,N_16116,N_16041);
xnor U16297 (N_16297,N_15673,N_15493);
and U16298 (N_16298,N_15761,N_15941);
nor U16299 (N_16299,N_16128,N_16092);
or U16300 (N_16300,N_15374,N_15436);
and U16301 (N_16301,N_15964,N_15336);
nor U16302 (N_16302,N_16090,N_15829);
and U16303 (N_16303,N_15031,N_15465);
and U16304 (N_16304,N_15799,N_15094);
or U16305 (N_16305,N_16069,N_15541);
xor U16306 (N_16306,N_16089,N_15918);
and U16307 (N_16307,N_16175,N_15515);
nor U16308 (N_16308,N_15656,N_15407);
nand U16309 (N_16309,N_15864,N_16214);
xor U16310 (N_16310,N_15269,N_16224);
xor U16311 (N_16311,N_15180,N_15975);
or U16312 (N_16312,N_16097,N_15748);
xor U16313 (N_16313,N_15395,N_15804);
xnor U16314 (N_16314,N_15133,N_15181);
nand U16315 (N_16315,N_16233,N_15371);
nor U16316 (N_16316,N_15331,N_15688);
nand U16317 (N_16317,N_16099,N_15989);
and U16318 (N_16318,N_15854,N_15569);
xnor U16319 (N_16319,N_15320,N_15711);
or U16320 (N_16320,N_15533,N_15236);
nand U16321 (N_16321,N_16101,N_16036);
xor U16322 (N_16322,N_15650,N_15274);
nor U16323 (N_16323,N_15704,N_16048);
xor U16324 (N_16324,N_16084,N_16145);
and U16325 (N_16325,N_15623,N_15980);
or U16326 (N_16326,N_15522,N_15098);
and U16327 (N_16327,N_15640,N_15702);
nor U16328 (N_16328,N_15179,N_15473);
nor U16329 (N_16329,N_15889,N_15225);
xnor U16330 (N_16330,N_16023,N_15886);
nand U16331 (N_16331,N_15648,N_15922);
nand U16332 (N_16332,N_15409,N_15201);
nor U16333 (N_16333,N_15288,N_15300);
nand U16334 (N_16334,N_15950,N_15900);
or U16335 (N_16335,N_15567,N_16194);
nand U16336 (N_16336,N_15981,N_16035);
xor U16337 (N_16337,N_16204,N_15278);
nor U16338 (N_16338,N_15596,N_15723);
xor U16339 (N_16339,N_15223,N_15246);
nor U16340 (N_16340,N_15666,N_15840);
nand U16341 (N_16341,N_15555,N_15542);
nand U16342 (N_16342,N_15477,N_15318);
nand U16343 (N_16343,N_15537,N_16057);
or U16344 (N_16344,N_15327,N_16037);
nor U16345 (N_16345,N_15678,N_16185);
and U16346 (N_16346,N_16049,N_15810);
and U16347 (N_16347,N_16183,N_15872);
xor U16348 (N_16348,N_16162,N_15285);
or U16349 (N_16349,N_15464,N_15590);
nand U16350 (N_16350,N_15050,N_16002);
and U16351 (N_16351,N_15920,N_15446);
or U16352 (N_16352,N_15600,N_15633);
or U16353 (N_16353,N_16029,N_15364);
nand U16354 (N_16354,N_15204,N_16216);
or U16355 (N_16355,N_15203,N_16199);
or U16356 (N_16356,N_15803,N_16159);
xor U16357 (N_16357,N_16170,N_16058);
and U16358 (N_16358,N_15459,N_15116);
or U16359 (N_16359,N_15513,N_15562);
nor U16360 (N_16360,N_16028,N_15794);
or U16361 (N_16361,N_15945,N_15669);
nand U16362 (N_16362,N_15827,N_15379);
xnor U16363 (N_16363,N_15044,N_16177);
nor U16364 (N_16364,N_16138,N_15915);
nand U16365 (N_16365,N_16184,N_15063);
xor U16366 (N_16366,N_16045,N_15998);
or U16367 (N_16367,N_15077,N_16222);
nor U16368 (N_16368,N_15113,N_15164);
nor U16369 (N_16369,N_15111,N_15720);
and U16370 (N_16370,N_15721,N_15797);
and U16371 (N_16371,N_15586,N_15088);
nor U16372 (N_16372,N_15885,N_15658);
xnor U16373 (N_16373,N_15891,N_15451);
xnor U16374 (N_16374,N_15976,N_16152);
nor U16375 (N_16375,N_15396,N_15420);
xor U16376 (N_16376,N_15001,N_15588);
xor U16377 (N_16377,N_15610,N_15399);
xnor U16378 (N_16378,N_15003,N_16211);
or U16379 (N_16379,N_15632,N_16239);
nor U16380 (N_16380,N_15469,N_15069);
or U16381 (N_16381,N_15281,N_15226);
nand U16382 (N_16382,N_15536,N_16228);
nor U16383 (N_16383,N_15314,N_16160);
or U16384 (N_16384,N_15247,N_15488);
or U16385 (N_16385,N_15051,N_15853);
or U16386 (N_16386,N_15103,N_15192);
xor U16387 (N_16387,N_15876,N_15937);
xnor U16388 (N_16388,N_15004,N_15530);
xnor U16389 (N_16389,N_15771,N_16122);
and U16390 (N_16390,N_15892,N_15636);
and U16391 (N_16391,N_15630,N_15557);
xor U16392 (N_16392,N_16236,N_15652);
and U16393 (N_16393,N_15757,N_15257);
or U16394 (N_16394,N_15674,N_16178);
nor U16395 (N_16395,N_15565,N_15765);
xor U16396 (N_16396,N_15714,N_16051);
and U16397 (N_16397,N_15126,N_15628);
nor U16398 (N_16398,N_16004,N_15499);
and U16399 (N_16399,N_16019,N_15816);
nor U16400 (N_16400,N_15150,N_15241);
nor U16401 (N_16401,N_16190,N_16182);
nor U16402 (N_16402,N_15532,N_15747);
nor U16403 (N_16403,N_15500,N_15856);
nor U16404 (N_16404,N_15277,N_15725);
nand U16405 (N_16405,N_15412,N_15579);
nor U16406 (N_16406,N_15660,N_15935);
nor U16407 (N_16407,N_15040,N_15137);
and U16408 (N_16408,N_15121,N_16072);
and U16409 (N_16409,N_15907,N_16168);
nor U16410 (N_16410,N_15439,N_16030);
nand U16411 (N_16411,N_15325,N_16098);
and U16412 (N_16412,N_15831,N_15763);
or U16413 (N_16413,N_15946,N_15786);
nor U16414 (N_16414,N_16056,N_15566);
or U16415 (N_16415,N_15060,N_16240);
and U16416 (N_16416,N_15926,N_15701);
and U16417 (N_16417,N_15117,N_16033);
nor U16418 (N_16418,N_15115,N_16007);
or U16419 (N_16419,N_15011,N_15461);
and U16420 (N_16420,N_15048,N_15329);
and U16421 (N_16421,N_15531,N_15071);
nor U16422 (N_16422,N_15708,N_16210);
and U16423 (N_16423,N_15087,N_15235);
nand U16424 (N_16424,N_15049,N_15143);
or U16425 (N_16425,N_15070,N_15967);
nor U16426 (N_16426,N_15523,N_15248);
nor U16427 (N_16427,N_15114,N_15847);
nand U16428 (N_16428,N_16237,N_15401);
nor U16429 (N_16429,N_15099,N_15929);
and U16430 (N_16430,N_16034,N_15333);
nor U16431 (N_16431,N_16150,N_15729);
nor U16432 (N_16432,N_15159,N_15514);
or U16433 (N_16433,N_16107,N_15474);
nand U16434 (N_16434,N_16203,N_15538);
xnor U16435 (N_16435,N_16187,N_15382);
xor U16436 (N_16436,N_15993,N_15219);
or U16437 (N_16437,N_15437,N_15153);
or U16438 (N_16438,N_15102,N_16061);
nand U16439 (N_16439,N_15611,N_15254);
or U16440 (N_16440,N_15850,N_15503);
xnor U16441 (N_16441,N_15010,N_15619);
xnor U16442 (N_16442,N_15166,N_15138);
and U16443 (N_16443,N_15713,N_15863);
nand U16444 (N_16444,N_15082,N_15564);
or U16445 (N_16445,N_16085,N_16246);
nor U16446 (N_16446,N_15559,N_16094);
and U16447 (N_16447,N_15791,N_15642);
xnor U16448 (N_16448,N_15904,N_15517);
nor U16449 (N_16449,N_15061,N_16047);
and U16450 (N_16450,N_15074,N_16143);
xnor U16451 (N_16451,N_15584,N_15434);
nand U16452 (N_16452,N_15463,N_15172);
nor U16453 (N_16453,N_15047,N_15505);
nand U16454 (N_16454,N_15957,N_15080);
nor U16455 (N_16455,N_15234,N_15097);
nand U16456 (N_16456,N_15306,N_15635);
or U16457 (N_16457,N_15681,N_16024);
xnor U16458 (N_16458,N_15059,N_15846);
and U16459 (N_16459,N_15250,N_15661);
nand U16460 (N_16460,N_15842,N_15388);
and U16461 (N_16461,N_16163,N_15366);
or U16462 (N_16462,N_15970,N_15356);
xor U16463 (N_16463,N_15602,N_15156);
or U16464 (N_16464,N_15836,N_16102);
nand U16465 (N_16465,N_16014,N_15141);
or U16466 (N_16466,N_15629,N_16071);
nor U16467 (N_16467,N_15762,N_16018);
nand U16468 (N_16468,N_15359,N_15140);
or U16469 (N_16469,N_15744,N_15966);
nand U16470 (N_16470,N_15693,N_15732);
nor U16471 (N_16471,N_15147,N_15749);
xor U16472 (N_16472,N_15547,N_15719);
nor U16473 (N_16473,N_15825,N_16201);
or U16474 (N_16474,N_15131,N_16188);
nor U16475 (N_16475,N_15389,N_15175);
nand U16476 (N_16476,N_15750,N_15550);
or U16477 (N_16477,N_15107,N_15258);
nor U16478 (N_16478,N_15968,N_16142);
nor U16479 (N_16479,N_15026,N_15317);
or U16480 (N_16480,N_15545,N_15780);
and U16481 (N_16481,N_15662,N_15092);
and U16482 (N_16482,N_15358,N_15654);
or U16483 (N_16483,N_15185,N_15734);
or U16484 (N_16484,N_15252,N_15837);
nand U16485 (N_16485,N_15284,N_16130);
and U16486 (N_16486,N_15301,N_15826);
or U16487 (N_16487,N_15264,N_15350);
or U16488 (N_16488,N_15450,N_16217);
xnor U16489 (N_16489,N_16249,N_15458);
nand U16490 (N_16490,N_15471,N_15724);
nand U16491 (N_16491,N_15527,N_16082);
or U16492 (N_16492,N_15974,N_15709);
or U16493 (N_16493,N_15476,N_16126);
nor U16494 (N_16494,N_15617,N_15381);
nor U16495 (N_16495,N_15183,N_15824);
or U16496 (N_16496,N_15400,N_15062);
or U16497 (N_16497,N_15079,N_15940);
or U16498 (N_16498,N_15170,N_16077);
and U16499 (N_16499,N_15188,N_15135);
xnor U16500 (N_16500,N_15934,N_15085);
nor U16501 (N_16501,N_15859,N_15037);
nor U16502 (N_16502,N_16022,N_15109);
xor U16503 (N_16503,N_15735,N_15534);
xor U16504 (N_16504,N_16050,N_15018);
xor U16505 (N_16505,N_15406,N_15665);
xor U16506 (N_16506,N_15122,N_15835);
nand U16507 (N_16507,N_15008,N_15174);
nor U16508 (N_16508,N_15032,N_16156);
xnor U16509 (N_16509,N_15783,N_15643);
and U16510 (N_16510,N_15132,N_15575);
or U16511 (N_16511,N_15647,N_15490);
nand U16512 (N_16512,N_15393,N_15279);
and U16513 (N_16513,N_15418,N_15367);
nor U16514 (N_16514,N_16167,N_15948);
and U16515 (N_16515,N_15667,N_15986);
and U16516 (N_16516,N_15035,N_15956);
nand U16517 (N_16517,N_15741,N_15322);
and U16518 (N_16518,N_15270,N_15220);
nand U16519 (N_16519,N_15951,N_16103);
nor U16520 (N_16520,N_15144,N_15043);
nand U16521 (N_16521,N_15430,N_15064);
nor U16522 (N_16522,N_15193,N_15139);
nand U16523 (N_16523,N_15873,N_15597);
nand U16524 (N_16524,N_15808,N_15798);
or U16525 (N_16525,N_15508,N_16039);
nand U16526 (N_16526,N_15066,N_15200);
xnor U16527 (N_16527,N_16165,N_16006);
xnor U16528 (N_16528,N_15449,N_15930);
and U16529 (N_16529,N_16078,N_16245);
or U16530 (N_16530,N_15577,N_15233);
nand U16531 (N_16531,N_15089,N_15425);
xor U16532 (N_16532,N_15052,N_16060);
xnor U16533 (N_16533,N_15222,N_15736);
and U16534 (N_16534,N_15484,N_15676);
xor U16535 (N_16535,N_16021,N_15700);
and U16536 (N_16536,N_16225,N_16070);
xor U16537 (N_16537,N_16075,N_15007);
nand U16538 (N_16538,N_15718,N_15483);
or U16539 (N_16539,N_15638,N_15108);
xnor U16540 (N_16540,N_16105,N_15255);
and U16541 (N_16541,N_16112,N_15291);
xor U16542 (N_16542,N_15782,N_15737);
and U16543 (N_16543,N_15142,N_15973);
or U16544 (N_16544,N_15888,N_15942);
nor U16545 (N_16545,N_15625,N_15013);
and U16546 (N_16546,N_15195,N_16065);
or U16547 (N_16547,N_15563,N_15106);
xnor U16548 (N_16548,N_15104,N_15302);
and U16549 (N_16549,N_15595,N_15354);
xor U16550 (N_16550,N_15145,N_15697);
xor U16551 (N_16551,N_15698,N_15182);
nor U16552 (N_16552,N_15385,N_15240);
nor U16553 (N_16553,N_15423,N_16123);
or U16554 (N_16554,N_15232,N_15519);
nand U16555 (N_16555,N_15843,N_15478);
nand U16556 (N_16556,N_15154,N_15751);
or U16557 (N_16557,N_15161,N_15310);
nand U16558 (N_16558,N_15813,N_15841);
and U16559 (N_16559,N_15578,N_16100);
nor U16560 (N_16560,N_16003,N_15119);
xor U16561 (N_16561,N_16074,N_15100);
nor U16562 (N_16562,N_16108,N_15020);
and U16563 (N_16563,N_15862,N_15733);
and U16564 (N_16564,N_15178,N_16119);
and U16565 (N_16565,N_15861,N_15546);
nand U16566 (N_16566,N_15641,N_15448);
and U16567 (N_16567,N_16135,N_15256);
xnor U16568 (N_16568,N_15271,N_15454);
xor U16569 (N_16569,N_16169,N_16172);
nand U16570 (N_16570,N_15727,N_16011);
and U16571 (N_16571,N_15305,N_15447);
and U16572 (N_16572,N_15238,N_15939);
nand U16573 (N_16573,N_15710,N_15249);
nand U16574 (N_16574,N_15938,N_15149);
nand U16575 (N_16575,N_15591,N_16215);
nand U16576 (N_16576,N_15282,N_15944);
nor U16577 (N_16577,N_15072,N_15884);
xor U16578 (N_16578,N_15491,N_15955);
xnor U16579 (N_16579,N_15985,N_15839);
and U16580 (N_16580,N_15042,N_15294);
xnor U16581 (N_16581,N_16059,N_15245);
or U16582 (N_16582,N_15814,N_15883);
or U16583 (N_16583,N_16171,N_15960);
or U16584 (N_16584,N_15787,N_15509);
xnor U16585 (N_16585,N_15624,N_16202);
xor U16586 (N_16586,N_15332,N_15677);
nor U16587 (N_16587,N_15205,N_15781);
nand U16588 (N_16588,N_16127,N_16147);
and U16589 (N_16589,N_15592,N_15832);
nor U16590 (N_16590,N_15497,N_15849);
nand U16591 (N_16591,N_15309,N_16118);
xnor U16592 (N_16592,N_16044,N_15176);
nand U16593 (N_16593,N_16241,N_15479);
nand U16594 (N_16594,N_15978,N_15820);
xor U16595 (N_16595,N_15275,N_15173);
and U16596 (N_16596,N_15570,N_15742);
xnor U16597 (N_16597,N_15913,N_15769);
nand U16598 (N_16598,N_15760,N_15927);
and U16599 (N_16599,N_15758,N_15021);
nor U16600 (N_16600,N_15615,N_16153);
nor U16601 (N_16601,N_15961,N_15199);
xnor U16602 (N_16602,N_15081,N_15984);
nand U16603 (N_16603,N_15158,N_16139);
nand U16604 (N_16604,N_16104,N_16166);
and U16605 (N_16605,N_15583,N_15576);
nor U16606 (N_16606,N_16193,N_15373);
xor U16607 (N_16607,N_16027,N_15540);
and U16608 (N_16608,N_15002,N_15912);
xnor U16609 (N_16609,N_15812,N_15330);
nor U16610 (N_16610,N_15206,N_15009);
xnor U16611 (N_16611,N_15699,N_16081);
nor U16612 (N_16612,N_15337,N_15809);
or U16613 (N_16613,N_15157,N_15387);
xor U16614 (N_16614,N_15792,N_15441);
and U16615 (N_16615,N_15715,N_15838);
xor U16616 (N_16616,N_15746,N_15867);
nand U16617 (N_16617,N_16197,N_15865);
nor U16618 (N_16618,N_15426,N_15753);
nand U16619 (N_16619,N_16164,N_15796);
xnor U16620 (N_16620,N_15593,N_15785);
and U16621 (N_16621,N_15560,N_16005);
nand U16622 (N_16622,N_16198,N_15405);
and U16623 (N_16623,N_15457,N_15598);
xnor U16624 (N_16624,N_15404,N_15162);
or U16625 (N_16625,N_15403,N_15807);
nor U16626 (N_16626,N_15263,N_15991);
nand U16627 (N_16627,N_15777,N_16013);
or U16628 (N_16628,N_15994,N_15024);
and U16629 (N_16629,N_15506,N_16080);
nor U16630 (N_16630,N_15351,N_15287);
and U16631 (N_16631,N_15027,N_15445);
and U16632 (N_16632,N_15218,N_15198);
nor U16633 (N_16633,N_15504,N_15801);
nand U16634 (N_16634,N_15229,N_15589);
and U16635 (N_16635,N_15759,N_15726);
nor U16636 (N_16636,N_15995,N_15695);
or U16637 (N_16637,N_15811,N_16012);
xor U16638 (N_16638,N_15874,N_16086);
and U16639 (N_16639,N_15455,N_16096);
nor U16640 (N_16640,N_15187,N_15415);
nor U16641 (N_16641,N_15594,N_15462);
or U16642 (N_16642,N_15899,N_16212);
and U16643 (N_16643,N_15717,N_15902);
nand U16644 (N_16644,N_15386,N_16132);
and U16645 (N_16645,N_15068,N_15129);
xnor U16646 (N_16646,N_15347,N_15034);
nand U16647 (N_16647,N_15599,N_16064);
nand U16648 (N_16648,N_15516,N_15215);
nor U16649 (N_16649,N_15355,N_15703);
nand U16650 (N_16650,N_16010,N_15905);
xor U16651 (N_16651,N_15202,N_15209);
nor U16652 (N_16652,N_15039,N_16244);
xnor U16653 (N_16653,N_15148,N_15988);
or U16654 (N_16654,N_15408,N_15016);
or U16655 (N_16655,N_16000,N_15303);
and U16656 (N_16656,N_16158,N_15384);
nand U16657 (N_16657,N_15308,N_15324);
and U16658 (N_16658,N_15554,N_15773);
xnor U16659 (N_16659,N_15932,N_16181);
and U16660 (N_16660,N_15774,N_15919);
nor U16661 (N_16661,N_15028,N_15844);
or U16662 (N_16662,N_15571,N_15101);
and U16663 (N_16663,N_15645,N_16242);
and U16664 (N_16664,N_15878,N_15690);
or U16665 (N_16665,N_15631,N_15413);
or U16666 (N_16666,N_15372,N_15296);
or U16667 (N_16667,N_15805,N_15467);
or U16668 (N_16668,N_15685,N_15495);
and U16669 (N_16669,N_15340,N_15914);
xor U16670 (N_16670,N_15058,N_16247);
nand U16671 (N_16671,N_15391,N_15558);
or U16672 (N_16672,N_15521,N_15151);
or U16673 (N_16673,N_15283,N_16087);
nor U16674 (N_16674,N_15684,N_15696);
nand U16675 (N_16675,N_15764,N_15925);
nor U16676 (N_16676,N_16043,N_15217);
nor U16677 (N_16677,N_15075,N_15855);
nand U16678 (N_16678,N_16144,N_15411);
or U16679 (N_16679,N_15261,N_15438);
or U16680 (N_16680,N_15452,N_15924);
or U16681 (N_16681,N_15834,N_16157);
or U16682 (N_16682,N_15416,N_15307);
nand U16683 (N_16683,N_15128,N_15784);
xor U16684 (N_16684,N_15680,N_15917);
or U16685 (N_16685,N_16124,N_15996);
nand U16686 (N_16686,N_15928,N_15237);
or U16687 (N_16687,N_16230,N_15655);
xor U16688 (N_16688,N_15520,N_15417);
xor U16689 (N_16689,N_15823,N_15605);
xor U16690 (N_16690,N_15230,N_15694);
nor U16691 (N_16691,N_15155,N_15357);
xnor U16692 (N_16692,N_15496,N_15014);
and U16693 (N_16693,N_15163,N_15953);
and U16694 (N_16694,N_15422,N_15553);
or U16695 (N_16695,N_15038,N_15730);
nand U16696 (N_16696,N_15707,N_15908);
and U16697 (N_16697,N_16079,N_15344);
and U16698 (N_16698,N_15890,N_15963);
and U16699 (N_16699,N_15815,N_15679);
or U16700 (N_16700,N_15860,N_15472);
and U16701 (N_16701,N_15015,N_15319);
xnor U16702 (N_16702,N_15898,N_15244);
or U16703 (N_16703,N_15909,N_15273);
xor U16704 (N_16704,N_15489,N_15073);
nor U16705 (N_16705,N_15671,N_15321);
nand U16706 (N_16706,N_16180,N_15041);
nand U16707 (N_16707,N_15239,N_15216);
and U16708 (N_16708,N_15341,N_15526);
or U16709 (N_16709,N_15194,N_15189);
or U16710 (N_16710,N_15947,N_15949);
nor U16711 (N_16711,N_15880,N_15691);
nor U16712 (N_16712,N_16062,N_16088);
and U16713 (N_16713,N_15745,N_15378);
xnor U16714 (N_16714,N_15644,N_15512);
or U16715 (N_16715,N_15453,N_15670);
or U16716 (N_16716,N_15312,N_16229);
and U16717 (N_16717,N_16042,N_16161);
nor U16718 (N_16718,N_16248,N_15466);
nor U16719 (N_16719,N_16232,N_16121);
or U16720 (N_16720,N_15475,N_15936);
xnor U16721 (N_16721,N_16151,N_15124);
nand U16722 (N_16722,N_15335,N_15375);
nor U16723 (N_16723,N_15136,N_15772);
nor U16724 (N_16724,N_15268,N_15510);
nor U16725 (N_16725,N_16148,N_15017);
nand U16726 (N_16726,N_15524,N_15293);
xor U16727 (N_16727,N_15440,N_15767);
nand U16728 (N_16728,N_15295,N_15982);
or U16729 (N_16729,N_15326,N_15768);
nor U16730 (N_16730,N_15429,N_15752);
xor U16731 (N_16731,N_15906,N_15299);
nor U16732 (N_16732,N_16149,N_15755);
xnor U16733 (N_16733,N_15999,N_15424);
xnor U16734 (N_16734,N_15006,N_15857);
nor U16735 (N_16735,N_15663,N_15152);
xor U16736 (N_16736,N_15672,N_15086);
nand U16737 (N_16737,N_15848,N_15916);
or U16738 (N_16738,N_15057,N_15398);
nand U16739 (N_16739,N_15581,N_15377);
or U16740 (N_16740,N_16206,N_15779);
nor U16741 (N_16741,N_15146,N_16106);
or U16742 (N_16742,N_15706,N_15620);
or U16743 (N_16743,N_15601,N_15776);
or U16744 (N_16744,N_15561,N_15535);
nand U16745 (N_16745,N_15675,N_15743);
nand U16746 (N_16746,N_15191,N_15169);
nand U16747 (N_16747,N_15486,N_15646);
nand U16748 (N_16748,N_15213,N_15683);
nor U16749 (N_16749,N_15830,N_15903);
or U16750 (N_16750,N_15800,N_15093);
or U16751 (N_16751,N_16113,N_15055);
and U16752 (N_16752,N_15125,N_15612);
and U16753 (N_16753,N_15431,N_15289);
nor U16754 (N_16754,N_15046,N_15078);
nor U16755 (N_16755,N_15227,N_15091);
nor U16756 (N_16756,N_15444,N_15297);
nand U16757 (N_16757,N_15971,N_15502);
nor U16758 (N_16758,N_15637,N_15253);
nand U16759 (N_16759,N_15362,N_15428);
and U16760 (N_16760,N_15692,N_15210);
xor U16761 (N_16761,N_16238,N_15130);
or U16762 (N_16762,N_15770,N_15910);
and U16763 (N_16763,N_15539,N_16066);
nand U16764 (N_16764,N_15582,N_15952);
nand U16765 (N_16765,N_16205,N_15893);
or U16766 (N_16766,N_15875,N_15023);
nand U16767 (N_16767,N_15316,N_15292);
xnor U16768 (N_16768,N_16137,N_15614);
nor U16769 (N_16769,N_16055,N_15033);
and U16770 (N_16770,N_15969,N_15328);
nand U16771 (N_16771,N_15435,N_15460);
and U16772 (N_16772,N_15368,N_15481);
nor U16773 (N_16773,N_15977,N_15649);
or U16774 (N_16774,N_15267,N_15342);
or U16775 (N_16775,N_16091,N_16140);
nand U16776 (N_16776,N_15470,N_15518);
xor U16777 (N_16777,N_16146,N_15627);
nor U16778 (N_16778,N_15828,N_15979);
nand U16779 (N_16779,N_16117,N_15485);
nor U16780 (N_16780,N_16063,N_15687);
nand U16781 (N_16781,N_15456,N_15468);
nand U16782 (N_16782,N_15338,N_16038);
nand U16783 (N_16783,N_16001,N_16154);
or U16784 (N_16784,N_15432,N_15160);
nor U16785 (N_16785,N_15871,N_15740);
and U16786 (N_16786,N_15616,N_15958);
nand U16787 (N_16787,N_15224,N_15123);
xor U16788 (N_16788,N_15603,N_15266);
and U16789 (N_16789,N_15498,N_15795);
or U16790 (N_16790,N_15585,N_15228);
xor U16791 (N_16791,N_16186,N_16025);
xnor U16792 (N_16792,N_15618,N_15851);
nor U16793 (N_16793,N_15728,N_16179);
xnor U16794 (N_16794,N_15207,N_16114);
nor U16795 (N_16795,N_15397,N_16095);
nand U16796 (N_16796,N_15894,N_15383);
nand U16797 (N_16797,N_15419,N_15414);
xor U16798 (N_16798,N_15739,N_15005);
or U16799 (N_16799,N_15525,N_16231);
and U16800 (N_16800,N_16192,N_16054);
and U16801 (N_16801,N_16083,N_15421);
and U16802 (N_16802,N_15613,N_15881);
nor U16803 (N_16803,N_15353,N_15221);
nor U16804 (N_16804,N_15716,N_15604);
and U16805 (N_16805,N_16026,N_15345);
and U16806 (N_16806,N_16015,N_15433);
nand U16807 (N_16807,N_16093,N_15821);
xor U16808 (N_16808,N_16115,N_16141);
nor U16809 (N_16809,N_15231,N_15012);
nor U16810 (N_16810,N_15529,N_16227);
or U16811 (N_16811,N_15651,N_15943);
or U16812 (N_16812,N_16176,N_15208);
or U16813 (N_16813,N_15363,N_15190);
or U16814 (N_16814,N_15211,N_15664);
nand U16815 (N_16815,N_15494,N_15921);
nand U16816 (N_16816,N_15870,N_15095);
and U16817 (N_16817,N_15186,N_15280);
nor U16818 (N_16818,N_15622,N_15394);
and U16819 (N_16819,N_15315,N_15096);
nor U16820 (N_16820,N_15778,N_16076);
nor U16821 (N_16821,N_15657,N_15895);
and U16822 (N_16822,N_15022,N_15933);
nand U16823 (N_16823,N_15897,N_15290);
xnor U16824 (N_16824,N_16209,N_15689);
or U16825 (N_16825,N_15390,N_15360);
nor U16826 (N_16826,N_15065,N_15242);
nor U16827 (N_16827,N_15997,N_15668);
and U16828 (N_16828,N_15365,N_15480);
and U16829 (N_16829,N_16111,N_15858);
and U16830 (N_16830,N_15705,N_16173);
nor U16831 (N_16831,N_16109,N_15334);
nand U16832 (N_16832,N_15959,N_15802);
and U16833 (N_16833,N_15817,N_15243);
nor U16834 (N_16834,N_15822,N_15806);
xnor U16835 (N_16835,N_16009,N_16136);
and U16836 (N_16836,N_15544,N_16120);
and U16837 (N_16837,N_15053,N_15311);
or U16838 (N_16838,N_15686,N_15634);
and U16839 (N_16839,N_15376,N_15076);
xor U16840 (N_16840,N_15251,N_15580);
and U16841 (N_16841,N_15887,N_15025);
nand U16842 (N_16842,N_15262,N_16191);
nand U16843 (N_16843,N_15392,N_16155);
nand U16844 (N_16844,N_15682,N_15492);
xnor U16845 (N_16845,N_15105,N_15265);
nand U16846 (N_16846,N_15621,N_15833);
and U16847 (N_16847,N_15793,N_15369);
or U16848 (N_16848,N_15877,N_15276);
xor U16849 (N_16849,N_15067,N_15868);
and U16850 (N_16850,N_15606,N_15083);
nor U16851 (N_16851,N_15626,N_16110);
nand U16852 (N_16852,N_16032,N_15722);
xnor U16853 (N_16853,N_15348,N_15019);
xor U16854 (N_16854,N_15551,N_15659);
nand U16855 (N_16855,N_16052,N_15528);
nor U16856 (N_16856,N_15896,N_15442);
or U16857 (N_16857,N_15380,N_15361);
nor U16858 (N_16858,N_16129,N_16221);
nor U16859 (N_16859,N_15410,N_15352);
nor U16860 (N_16860,N_15120,N_15343);
nor U16861 (N_16861,N_15196,N_15110);
nor U16862 (N_16862,N_15845,N_15990);
xnor U16863 (N_16863,N_15212,N_16220);
nor U16864 (N_16864,N_15901,N_15965);
xor U16865 (N_16865,N_16133,N_15607);
and U16866 (N_16866,N_15084,N_16067);
or U16867 (N_16867,N_15112,N_16219);
nand U16868 (N_16868,N_15923,N_15882);
nor U16869 (N_16869,N_15819,N_16235);
xor U16870 (N_16870,N_15866,N_15653);
nand U16871 (N_16871,N_15298,N_16213);
xor U16872 (N_16872,N_16046,N_15573);
nand U16873 (N_16873,N_15184,N_16134);
and U16874 (N_16874,N_15911,N_15197);
nor U16875 (N_16875,N_16043,N_15201);
nor U16876 (N_16876,N_16225,N_15159);
nand U16877 (N_16877,N_15260,N_16061);
and U16878 (N_16878,N_15032,N_15737);
nor U16879 (N_16879,N_15949,N_16224);
nand U16880 (N_16880,N_15543,N_16121);
and U16881 (N_16881,N_15513,N_15587);
nor U16882 (N_16882,N_16184,N_15548);
xor U16883 (N_16883,N_15337,N_15126);
nand U16884 (N_16884,N_15161,N_15317);
xor U16885 (N_16885,N_16068,N_15497);
xor U16886 (N_16886,N_15660,N_15543);
xor U16887 (N_16887,N_15162,N_15431);
nor U16888 (N_16888,N_15202,N_16188);
nand U16889 (N_16889,N_16169,N_16242);
or U16890 (N_16890,N_15174,N_15819);
nand U16891 (N_16891,N_16099,N_15879);
nand U16892 (N_16892,N_15068,N_15065);
nand U16893 (N_16893,N_15415,N_16085);
nor U16894 (N_16894,N_16070,N_15808);
nand U16895 (N_16895,N_15830,N_16145);
nand U16896 (N_16896,N_15368,N_15156);
nand U16897 (N_16897,N_15958,N_15340);
nor U16898 (N_16898,N_16156,N_15052);
or U16899 (N_16899,N_15680,N_15775);
or U16900 (N_16900,N_15497,N_15158);
or U16901 (N_16901,N_15697,N_16082);
or U16902 (N_16902,N_15433,N_15471);
and U16903 (N_16903,N_15323,N_15348);
nand U16904 (N_16904,N_15235,N_16020);
and U16905 (N_16905,N_15127,N_16085);
nand U16906 (N_16906,N_15751,N_15456);
xor U16907 (N_16907,N_15075,N_15641);
and U16908 (N_16908,N_15860,N_15077);
nand U16909 (N_16909,N_15600,N_15610);
nand U16910 (N_16910,N_15539,N_15343);
or U16911 (N_16911,N_16038,N_15452);
nand U16912 (N_16912,N_15185,N_15368);
or U16913 (N_16913,N_15787,N_15550);
and U16914 (N_16914,N_15272,N_15518);
or U16915 (N_16915,N_16218,N_15543);
and U16916 (N_16916,N_15249,N_15387);
nor U16917 (N_16917,N_15035,N_16015);
and U16918 (N_16918,N_15679,N_15787);
nor U16919 (N_16919,N_15850,N_15453);
nand U16920 (N_16920,N_16012,N_16080);
and U16921 (N_16921,N_15944,N_15203);
xor U16922 (N_16922,N_15437,N_15581);
nand U16923 (N_16923,N_16109,N_15348);
and U16924 (N_16924,N_15670,N_15522);
and U16925 (N_16925,N_15442,N_16128);
nand U16926 (N_16926,N_15389,N_16053);
or U16927 (N_16927,N_16114,N_16043);
xor U16928 (N_16928,N_15967,N_16234);
nor U16929 (N_16929,N_15045,N_15305);
and U16930 (N_16930,N_15998,N_15453);
nor U16931 (N_16931,N_15077,N_15467);
xor U16932 (N_16932,N_15651,N_15556);
and U16933 (N_16933,N_16049,N_15676);
xor U16934 (N_16934,N_15822,N_15812);
or U16935 (N_16935,N_15052,N_15453);
xor U16936 (N_16936,N_15793,N_16078);
nor U16937 (N_16937,N_15901,N_15894);
and U16938 (N_16938,N_16088,N_15021);
or U16939 (N_16939,N_15005,N_15881);
xor U16940 (N_16940,N_16190,N_15495);
or U16941 (N_16941,N_16229,N_15167);
nor U16942 (N_16942,N_15297,N_15731);
and U16943 (N_16943,N_15557,N_15588);
and U16944 (N_16944,N_16149,N_15762);
and U16945 (N_16945,N_15714,N_15559);
xor U16946 (N_16946,N_15903,N_15416);
and U16947 (N_16947,N_15930,N_16173);
or U16948 (N_16948,N_15204,N_15088);
or U16949 (N_16949,N_16145,N_15804);
nand U16950 (N_16950,N_16153,N_15534);
xor U16951 (N_16951,N_15817,N_15810);
nor U16952 (N_16952,N_15328,N_16140);
xnor U16953 (N_16953,N_15009,N_15230);
nand U16954 (N_16954,N_15405,N_15741);
or U16955 (N_16955,N_15598,N_15340);
nand U16956 (N_16956,N_15450,N_15676);
nand U16957 (N_16957,N_15526,N_15087);
or U16958 (N_16958,N_15997,N_15827);
and U16959 (N_16959,N_15032,N_16248);
and U16960 (N_16960,N_16002,N_15286);
nor U16961 (N_16961,N_15258,N_16053);
and U16962 (N_16962,N_15156,N_15214);
and U16963 (N_16963,N_16080,N_15245);
and U16964 (N_16964,N_15001,N_15780);
nor U16965 (N_16965,N_16191,N_15830);
nand U16966 (N_16966,N_15004,N_15493);
nor U16967 (N_16967,N_15497,N_15322);
nand U16968 (N_16968,N_15581,N_16244);
nand U16969 (N_16969,N_15225,N_16222);
nand U16970 (N_16970,N_15328,N_16218);
xor U16971 (N_16971,N_15335,N_15708);
nor U16972 (N_16972,N_15618,N_15839);
nor U16973 (N_16973,N_15838,N_15360);
xnor U16974 (N_16974,N_15196,N_15214);
and U16975 (N_16975,N_15246,N_15171);
xnor U16976 (N_16976,N_15713,N_15622);
nand U16977 (N_16977,N_15895,N_15883);
nand U16978 (N_16978,N_15158,N_15814);
nor U16979 (N_16979,N_15323,N_15013);
and U16980 (N_16980,N_15809,N_15254);
or U16981 (N_16981,N_15558,N_15282);
nand U16982 (N_16982,N_15639,N_16074);
xnor U16983 (N_16983,N_15336,N_15102);
and U16984 (N_16984,N_16115,N_15278);
xor U16985 (N_16985,N_16046,N_15002);
and U16986 (N_16986,N_15963,N_15171);
and U16987 (N_16987,N_15002,N_15700);
nand U16988 (N_16988,N_15758,N_16153);
and U16989 (N_16989,N_15640,N_16208);
and U16990 (N_16990,N_15013,N_15252);
nor U16991 (N_16991,N_15396,N_15419);
xor U16992 (N_16992,N_15446,N_16181);
nor U16993 (N_16993,N_15431,N_15484);
and U16994 (N_16994,N_16136,N_15940);
or U16995 (N_16995,N_15502,N_15799);
nand U16996 (N_16996,N_16241,N_15510);
xnor U16997 (N_16997,N_15428,N_16135);
nand U16998 (N_16998,N_15919,N_15908);
xnor U16999 (N_16999,N_16160,N_16228);
or U17000 (N_17000,N_16033,N_15148);
xnor U17001 (N_17001,N_15339,N_15189);
or U17002 (N_17002,N_15275,N_15267);
nor U17003 (N_17003,N_15686,N_15333);
xor U17004 (N_17004,N_15131,N_15205);
or U17005 (N_17005,N_16080,N_15098);
xor U17006 (N_17006,N_15067,N_15186);
nand U17007 (N_17007,N_16025,N_15381);
or U17008 (N_17008,N_15325,N_15126);
nand U17009 (N_17009,N_15756,N_15779);
or U17010 (N_17010,N_15122,N_15018);
and U17011 (N_17011,N_15954,N_15133);
nand U17012 (N_17012,N_15150,N_15220);
and U17013 (N_17013,N_15196,N_15207);
or U17014 (N_17014,N_15142,N_15069);
or U17015 (N_17015,N_15453,N_16102);
and U17016 (N_17016,N_15654,N_15439);
and U17017 (N_17017,N_15812,N_15375);
and U17018 (N_17018,N_15046,N_15155);
xor U17019 (N_17019,N_16224,N_15592);
nor U17020 (N_17020,N_15918,N_15699);
nand U17021 (N_17021,N_15679,N_16143);
or U17022 (N_17022,N_16196,N_16022);
and U17023 (N_17023,N_15626,N_15485);
xnor U17024 (N_17024,N_16247,N_15621);
and U17025 (N_17025,N_15780,N_15796);
xor U17026 (N_17026,N_15658,N_16105);
and U17027 (N_17027,N_15066,N_15636);
and U17028 (N_17028,N_15868,N_15191);
and U17029 (N_17029,N_15371,N_15306);
and U17030 (N_17030,N_15425,N_15840);
xnor U17031 (N_17031,N_15966,N_15143);
or U17032 (N_17032,N_15355,N_15136);
nor U17033 (N_17033,N_15780,N_15581);
xor U17034 (N_17034,N_15848,N_16132);
nand U17035 (N_17035,N_15354,N_15849);
and U17036 (N_17036,N_15498,N_15742);
nand U17037 (N_17037,N_15356,N_15344);
nor U17038 (N_17038,N_16130,N_15148);
nor U17039 (N_17039,N_16107,N_16100);
nand U17040 (N_17040,N_15767,N_15755);
nand U17041 (N_17041,N_15870,N_15219);
and U17042 (N_17042,N_16060,N_15708);
xnor U17043 (N_17043,N_15079,N_15424);
xnor U17044 (N_17044,N_15740,N_15054);
xnor U17045 (N_17045,N_15942,N_16113);
nand U17046 (N_17046,N_15109,N_15997);
and U17047 (N_17047,N_15133,N_15610);
nor U17048 (N_17048,N_15921,N_15172);
nor U17049 (N_17049,N_15360,N_15658);
xnor U17050 (N_17050,N_16184,N_15750);
xor U17051 (N_17051,N_15692,N_15287);
nand U17052 (N_17052,N_16123,N_15098);
or U17053 (N_17053,N_15175,N_15991);
nor U17054 (N_17054,N_15758,N_16151);
xor U17055 (N_17055,N_15730,N_15958);
nand U17056 (N_17056,N_15794,N_15566);
nor U17057 (N_17057,N_15623,N_15557);
nand U17058 (N_17058,N_15035,N_16106);
and U17059 (N_17059,N_15191,N_15859);
nor U17060 (N_17060,N_15879,N_15322);
or U17061 (N_17061,N_15695,N_16078);
xnor U17062 (N_17062,N_16249,N_15697);
nand U17063 (N_17063,N_15768,N_15221);
and U17064 (N_17064,N_15606,N_15835);
and U17065 (N_17065,N_15364,N_15116);
or U17066 (N_17066,N_15359,N_15912);
nor U17067 (N_17067,N_15935,N_16182);
nand U17068 (N_17068,N_15472,N_15367);
xor U17069 (N_17069,N_15330,N_16140);
or U17070 (N_17070,N_16226,N_15538);
xnor U17071 (N_17071,N_15011,N_15880);
nand U17072 (N_17072,N_15762,N_15606);
nor U17073 (N_17073,N_15061,N_15850);
or U17074 (N_17074,N_15587,N_15580);
and U17075 (N_17075,N_15660,N_15930);
and U17076 (N_17076,N_15674,N_15384);
or U17077 (N_17077,N_15398,N_15009);
nand U17078 (N_17078,N_15691,N_15710);
nor U17079 (N_17079,N_15869,N_15201);
nor U17080 (N_17080,N_15116,N_15612);
nor U17081 (N_17081,N_15911,N_16113);
or U17082 (N_17082,N_15490,N_15481);
nor U17083 (N_17083,N_16202,N_16164);
or U17084 (N_17084,N_15864,N_16229);
and U17085 (N_17085,N_15562,N_15286);
xnor U17086 (N_17086,N_15433,N_15604);
or U17087 (N_17087,N_16212,N_15457);
and U17088 (N_17088,N_15072,N_16138);
nor U17089 (N_17089,N_15617,N_15902);
xnor U17090 (N_17090,N_15734,N_15872);
nand U17091 (N_17091,N_15551,N_16195);
and U17092 (N_17092,N_15750,N_15397);
or U17093 (N_17093,N_15363,N_15823);
and U17094 (N_17094,N_15270,N_16135);
nor U17095 (N_17095,N_15377,N_15606);
nor U17096 (N_17096,N_15310,N_16167);
nand U17097 (N_17097,N_15310,N_16092);
xor U17098 (N_17098,N_15780,N_15494);
or U17099 (N_17099,N_15593,N_15757);
and U17100 (N_17100,N_15251,N_16029);
nand U17101 (N_17101,N_15469,N_15037);
xnor U17102 (N_17102,N_15635,N_15070);
and U17103 (N_17103,N_15443,N_15283);
nor U17104 (N_17104,N_16091,N_15189);
nand U17105 (N_17105,N_15649,N_15093);
nand U17106 (N_17106,N_15341,N_15156);
nor U17107 (N_17107,N_15084,N_15220);
nand U17108 (N_17108,N_15721,N_15075);
nand U17109 (N_17109,N_15443,N_16218);
and U17110 (N_17110,N_15612,N_15338);
or U17111 (N_17111,N_15999,N_15847);
nand U17112 (N_17112,N_16202,N_15161);
nand U17113 (N_17113,N_15357,N_16160);
xor U17114 (N_17114,N_15688,N_15161);
or U17115 (N_17115,N_15439,N_15729);
nor U17116 (N_17116,N_16230,N_16203);
or U17117 (N_17117,N_16039,N_16166);
and U17118 (N_17118,N_15702,N_16213);
nand U17119 (N_17119,N_15730,N_15755);
xor U17120 (N_17120,N_16241,N_15757);
nand U17121 (N_17121,N_15686,N_15642);
and U17122 (N_17122,N_16015,N_15512);
nand U17123 (N_17123,N_15611,N_15980);
nor U17124 (N_17124,N_15270,N_15332);
and U17125 (N_17125,N_15863,N_15435);
or U17126 (N_17126,N_15798,N_15319);
xor U17127 (N_17127,N_15258,N_15494);
nor U17128 (N_17128,N_15372,N_15234);
nor U17129 (N_17129,N_15531,N_15664);
nor U17130 (N_17130,N_16188,N_15066);
xor U17131 (N_17131,N_15446,N_15402);
or U17132 (N_17132,N_15914,N_15873);
nor U17133 (N_17133,N_15356,N_15217);
nand U17134 (N_17134,N_16144,N_15094);
xor U17135 (N_17135,N_15290,N_15860);
nand U17136 (N_17136,N_16064,N_15252);
nand U17137 (N_17137,N_15909,N_15224);
nor U17138 (N_17138,N_15461,N_15241);
and U17139 (N_17139,N_15582,N_15352);
xor U17140 (N_17140,N_15126,N_15355);
nor U17141 (N_17141,N_16028,N_16185);
xor U17142 (N_17142,N_15113,N_15803);
nand U17143 (N_17143,N_15481,N_15802);
or U17144 (N_17144,N_15675,N_15288);
nor U17145 (N_17145,N_15384,N_15557);
xnor U17146 (N_17146,N_16210,N_15986);
xor U17147 (N_17147,N_15230,N_15006);
nor U17148 (N_17148,N_15419,N_16020);
xor U17149 (N_17149,N_16198,N_15908);
and U17150 (N_17150,N_15866,N_15428);
and U17151 (N_17151,N_15764,N_16108);
or U17152 (N_17152,N_15215,N_15430);
and U17153 (N_17153,N_15501,N_16207);
and U17154 (N_17154,N_15303,N_16089);
xor U17155 (N_17155,N_15604,N_15019);
and U17156 (N_17156,N_16092,N_15717);
nor U17157 (N_17157,N_16138,N_15207);
or U17158 (N_17158,N_15701,N_15847);
nor U17159 (N_17159,N_16065,N_15788);
xor U17160 (N_17160,N_15149,N_15998);
nor U17161 (N_17161,N_15431,N_15595);
and U17162 (N_17162,N_15380,N_15850);
or U17163 (N_17163,N_16226,N_16055);
or U17164 (N_17164,N_15092,N_15038);
xor U17165 (N_17165,N_15151,N_15654);
xor U17166 (N_17166,N_15478,N_15553);
and U17167 (N_17167,N_15971,N_15145);
nor U17168 (N_17168,N_16035,N_15461);
nor U17169 (N_17169,N_15221,N_15756);
xnor U17170 (N_17170,N_15025,N_16157);
nor U17171 (N_17171,N_16186,N_15322);
nand U17172 (N_17172,N_15491,N_15541);
and U17173 (N_17173,N_15776,N_16107);
nor U17174 (N_17174,N_15307,N_16118);
nor U17175 (N_17175,N_15010,N_15322);
and U17176 (N_17176,N_15754,N_16053);
or U17177 (N_17177,N_15407,N_15609);
or U17178 (N_17178,N_16109,N_15618);
xor U17179 (N_17179,N_15869,N_15101);
and U17180 (N_17180,N_15839,N_15276);
nor U17181 (N_17181,N_15085,N_15299);
and U17182 (N_17182,N_15695,N_16028);
nor U17183 (N_17183,N_16180,N_15048);
nand U17184 (N_17184,N_15627,N_16159);
nand U17185 (N_17185,N_15994,N_15161);
and U17186 (N_17186,N_15931,N_16236);
nand U17187 (N_17187,N_15128,N_16187);
and U17188 (N_17188,N_16090,N_15511);
nand U17189 (N_17189,N_15925,N_15053);
or U17190 (N_17190,N_15969,N_15136);
or U17191 (N_17191,N_15950,N_16110);
and U17192 (N_17192,N_16243,N_15968);
xor U17193 (N_17193,N_15795,N_15941);
xor U17194 (N_17194,N_15241,N_15454);
xor U17195 (N_17195,N_15158,N_15867);
nand U17196 (N_17196,N_15001,N_15759);
xnor U17197 (N_17197,N_15588,N_15562);
or U17198 (N_17198,N_15457,N_15939);
and U17199 (N_17199,N_16209,N_15987);
nor U17200 (N_17200,N_15732,N_15225);
nand U17201 (N_17201,N_15526,N_15522);
and U17202 (N_17202,N_15872,N_15935);
nand U17203 (N_17203,N_15681,N_15983);
xor U17204 (N_17204,N_15378,N_15123);
or U17205 (N_17205,N_15392,N_15219);
nor U17206 (N_17206,N_15938,N_15852);
xnor U17207 (N_17207,N_16232,N_15704);
or U17208 (N_17208,N_15069,N_16243);
or U17209 (N_17209,N_15731,N_15580);
nand U17210 (N_17210,N_15038,N_15823);
and U17211 (N_17211,N_16118,N_16024);
nor U17212 (N_17212,N_15195,N_15342);
nor U17213 (N_17213,N_15739,N_15451);
and U17214 (N_17214,N_15605,N_15588);
nand U17215 (N_17215,N_15724,N_15942);
or U17216 (N_17216,N_15286,N_15814);
or U17217 (N_17217,N_15739,N_16034);
or U17218 (N_17218,N_15381,N_15161);
xnor U17219 (N_17219,N_15100,N_15949);
nor U17220 (N_17220,N_16014,N_16161);
nand U17221 (N_17221,N_15946,N_15811);
xor U17222 (N_17222,N_15037,N_16101);
nand U17223 (N_17223,N_15572,N_15901);
nor U17224 (N_17224,N_16125,N_15248);
nor U17225 (N_17225,N_15457,N_16015);
xnor U17226 (N_17226,N_15982,N_15707);
nor U17227 (N_17227,N_15577,N_15897);
nand U17228 (N_17228,N_15294,N_15838);
or U17229 (N_17229,N_15090,N_15926);
and U17230 (N_17230,N_15164,N_15515);
nor U17231 (N_17231,N_16185,N_15967);
xnor U17232 (N_17232,N_15172,N_15918);
nor U17233 (N_17233,N_16209,N_15127);
and U17234 (N_17234,N_15288,N_15958);
nor U17235 (N_17235,N_16034,N_15187);
and U17236 (N_17236,N_15025,N_15483);
xor U17237 (N_17237,N_15993,N_15263);
nor U17238 (N_17238,N_15955,N_16165);
nand U17239 (N_17239,N_15662,N_15005);
or U17240 (N_17240,N_16034,N_15502);
or U17241 (N_17241,N_15552,N_15415);
and U17242 (N_17242,N_16029,N_15720);
nor U17243 (N_17243,N_15964,N_15263);
or U17244 (N_17244,N_15932,N_15271);
xnor U17245 (N_17245,N_16230,N_15233);
and U17246 (N_17246,N_15600,N_15778);
nor U17247 (N_17247,N_15198,N_16198);
nor U17248 (N_17248,N_15979,N_15844);
nor U17249 (N_17249,N_15551,N_15529);
or U17250 (N_17250,N_16116,N_15058);
or U17251 (N_17251,N_15606,N_15757);
xor U17252 (N_17252,N_15618,N_15800);
and U17253 (N_17253,N_15352,N_15888);
nor U17254 (N_17254,N_15404,N_15515);
or U17255 (N_17255,N_15245,N_15028);
nor U17256 (N_17256,N_15242,N_15154);
nand U17257 (N_17257,N_15392,N_15686);
or U17258 (N_17258,N_15730,N_15514);
and U17259 (N_17259,N_15855,N_15613);
nor U17260 (N_17260,N_15502,N_15444);
and U17261 (N_17261,N_16022,N_15972);
nor U17262 (N_17262,N_15709,N_16112);
xor U17263 (N_17263,N_15522,N_15060);
nand U17264 (N_17264,N_15213,N_15510);
and U17265 (N_17265,N_15004,N_15606);
nand U17266 (N_17266,N_15058,N_15094);
xnor U17267 (N_17267,N_15740,N_16032);
xnor U17268 (N_17268,N_15242,N_16053);
xnor U17269 (N_17269,N_15818,N_16134);
nand U17270 (N_17270,N_15274,N_15878);
and U17271 (N_17271,N_15704,N_15710);
nor U17272 (N_17272,N_15838,N_15809);
nand U17273 (N_17273,N_15667,N_15560);
or U17274 (N_17274,N_16224,N_15473);
and U17275 (N_17275,N_15796,N_15425);
nor U17276 (N_17276,N_15125,N_15016);
nor U17277 (N_17277,N_15321,N_15406);
or U17278 (N_17278,N_15059,N_16153);
nor U17279 (N_17279,N_16056,N_16127);
nor U17280 (N_17280,N_15423,N_15828);
nor U17281 (N_17281,N_15831,N_15854);
xor U17282 (N_17282,N_15518,N_16051);
nor U17283 (N_17283,N_15895,N_15772);
nor U17284 (N_17284,N_15915,N_15149);
or U17285 (N_17285,N_15917,N_15781);
or U17286 (N_17286,N_16191,N_16023);
nor U17287 (N_17287,N_15110,N_16131);
xnor U17288 (N_17288,N_15968,N_15554);
nand U17289 (N_17289,N_15921,N_16177);
and U17290 (N_17290,N_16199,N_15338);
nand U17291 (N_17291,N_15228,N_15970);
xnor U17292 (N_17292,N_16135,N_15726);
nor U17293 (N_17293,N_15829,N_15174);
and U17294 (N_17294,N_15208,N_16217);
xnor U17295 (N_17295,N_15256,N_16175);
nand U17296 (N_17296,N_15152,N_15131);
or U17297 (N_17297,N_15326,N_15025);
nand U17298 (N_17298,N_15519,N_16111);
nor U17299 (N_17299,N_15403,N_15718);
nor U17300 (N_17300,N_15009,N_15902);
xnor U17301 (N_17301,N_16137,N_15680);
nand U17302 (N_17302,N_16033,N_15524);
or U17303 (N_17303,N_15046,N_16150);
xor U17304 (N_17304,N_15977,N_15560);
nand U17305 (N_17305,N_15454,N_15742);
nand U17306 (N_17306,N_16214,N_15338);
xor U17307 (N_17307,N_16169,N_16083);
and U17308 (N_17308,N_15422,N_15094);
or U17309 (N_17309,N_15770,N_15174);
xnor U17310 (N_17310,N_15380,N_15782);
nor U17311 (N_17311,N_15823,N_15669);
and U17312 (N_17312,N_15213,N_15426);
nand U17313 (N_17313,N_15020,N_15848);
xnor U17314 (N_17314,N_16190,N_15147);
nand U17315 (N_17315,N_15068,N_15460);
nand U17316 (N_17316,N_15025,N_15963);
or U17317 (N_17317,N_16111,N_15510);
nor U17318 (N_17318,N_15611,N_15512);
xnor U17319 (N_17319,N_15661,N_16236);
nor U17320 (N_17320,N_16165,N_16215);
or U17321 (N_17321,N_15212,N_15493);
and U17322 (N_17322,N_16106,N_15282);
nor U17323 (N_17323,N_16241,N_15061);
xor U17324 (N_17324,N_15995,N_15783);
nand U17325 (N_17325,N_16161,N_15718);
and U17326 (N_17326,N_15401,N_15893);
nand U17327 (N_17327,N_15534,N_16115);
and U17328 (N_17328,N_15322,N_15128);
or U17329 (N_17329,N_15247,N_16015);
or U17330 (N_17330,N_15528,N_15622);
xor U17331 (N_17331,N_15529,N_15897);
and U17332 (N_17332,N_15040,N_16177);
and U17333 (N_17333,N_16105,N_15999);
xor U17334 (N_17334,N_15013,N_15343);
nor U17335 (N_17335,N_15302,N_15132);
xnor U17336 (N_17336,N_15246,N_15474);
nand U17337 (N_17337,N_15728,N_15703);
or U17338 (N_17338,N_15697,N_15426);
nor U17339 (N_17339,N_15167,N_16106);
nand U17340 (N_17340,N_15216,N_15384);
or U17341 (N_17341,N_15633,N_15061);
xor U17342 (N_17342,N_16029,N_15932);
nand U17343 (N_17343,N_15908,N_15849);
or U17344 (N_17344,N_15717,N_15224);
xnor U17345 (N_17345,N_16188,N_15763);
and U17346 (N_17346,N_15289,N_15019);
or U17347 (N_17347,N_16211,N_15789);
and U17348 (N_17348,N_15887,N_15169);
and U17349 (N_17349,N_15151,N_15987);
nor U17350 (N_17350,N_15372,N_15594);
nor U17351 (N_17351,N_15367,N_15280);
and U17352 (N_17352,N_16113,N_16010);
or U17353 (N_17353,N_15223,N_15153);
and U17354 (N_17354,N_15352,N_15258);
and U17355 (N_17355,N_16033,N_15526);
or U17356 (N_17356,N_15013,N_15530);
nand U17357 (N_17357,N_15225,N_16064);
nand U17358 (N_17358,N_15850,N_15457);
and U17359 (N_17359,N_15955,N_15404);
nor U17360 (N_17360,N_15877,N_15670);
or U17361 (N_17361,N_15260,N_15351);
and U17362 (N_17362,N_15325,N_15213);
nor U17363 (N_17363,N_15328,N_15402);
nand U17364 (N_17364,N_15250,N_15546);
or U17365 (N_17365,N_15551,N_15983);
or U17366 (N_17366,N_16115,N_15356);
nand U17367 (N_17367,N_15933,N_16109);
nand U17368 (N_17368,N_15644,N_15558);
and U17369 (N_17369,N_15578,N_16129);
and U17370 (N_17370,N_15938,N_15185);
nor U17371 (N_17371,N_15739,N_15467);
xor U17372 (N_17372,N_15780,N_15645);
nand U17373 (N_17373,N_15972,N_15654);
and U17374 (N_17374,N_15175,N_15960);
xor U17375 (N_17375,N_16149,N_15659);
nand U17376 (N_17376,N_15774,N_15838);
or U17377 (N_17377,N_16069,N_15732);
xor U17378 (N_17378,N_15060,N_15380);
nand U17379 (N_17379,N_15035,N_15141);
or U17380 (N_17380,N_15277,N_15654);
and U17381 (N_17381,N_15020,N_16246);
xnor U17382 (N_17382,N_16075,N_15739);
nor U17383 (N_17383,N_15774,N_16152);
or U17384 (N_17384,N_15769,N_15133);
and U17385 (N_17385,N_15355,N_15437);
xor U17386 (N_17386,N_16074,N_15111);
nor U17387 (N_17387,N_15203,N_15416);
nor U17388 (N_17388,N_15187,N_15705);
nand U17389 (N_17389,N_15659,N_16190);
nor U17390 (N_17390,N_15825,N_16119);
or U17391 (N_17391,N_15595,N_15578);
xnor U17392 (N_17392,N_15066,N_15575);
nor U17393 (N_17393,N_15692,N_15967);
xor U17394 (N_17394,N_16244,N_15328);
or U17395 (N_17395,N_16070,N_15735);
and U17396 (N_17396,N_16152,N_15605);
nand U17397 (N_17397,N_15100,N_15964);
or U17398 (N_17398,N_15569,N_16130);
nand U17399 (N_17399,N_15432,N_15502);
nor U17400 (N_17400,N_15565,N_15170);
xnor U17401 (N_17401,N_15163,N_15909);
and U17402 (N_17402,N_16107,N_15306);
xor U17403 (N_17403,N_15893,N_15546);
nand U17404 (N_17404,N_15440,N_15495);
nand U17405 (N_17405,N_15737,N_15017);
or U17406 (N_17406,N_15705,N_15429);
and U17407 (N_17407,N_15034,N_15878);
and U17408 (N_17408,N_16153,N_15494);
or U17409 (N_17409,N_15865,N_15132);
xnor U17410 (N_17410,N_15817,N_15219);
nor U17411 (N_17411,N_15345,N_15047);
and U17412 (N_17412,N_15631,N_16101);
xnor U17413 (N_17413,N_15056,N_16109);
xnor U17414 (N_17414,N_15864,N_16065);
or U17415 (N_17415,N_15517,N_15453);
nand U17416 (N_17416,N_15636,N_15428);
nand U17417 (N_17417,N_15713,N_15107);
nor U17418 (N_17418,N_15731,N_15446);
xnor U17419 (N_17419,N_15558,N_16134);
xnor U17420 (N_17420,N_15005,N_15205);
xor U17421 (N_17421,N_15163,N_15148);
nor U17422 (N_17422,N_15149,N_15744);
nand U17423 (N_17423,N_16058,N_15830);
xnor U17424 (N_17424,N_15832,N_15409);
nand U17425 (N_17425,N_15864,N_15830);
nor U17426 (N_17426,N_15883,N_16180);
nand U17427 (N_17427,N_15671,N_15361);
xnor U17428 (N_17428,N_15001,N_15091);
xnor U17429 (N_17429,N_15943,N_15491);
and U17430 (N_17430,N_15078,N_15468);
nand U17431 (N_17431,N_16226,N_15914);
xnor U17432 (N_17432,N_15714,N_15754);
nand U17433 (N_17433,N_15045,N_15955);
or U17434 (N_17434,N_15025,N_15301);
nor U17435 (N_17435,N_15048,N_15113);
and U17436 (N_17436,N_15081,N_15428);
or U17437 (N_17437,N_16131,N_15024);
xnor U17438 (N_17438,N_15908,N_15571);
xnor U17439 (N_17439,N_15391,N_15201);
nor U17440 (N_17440,N_15129,N_15517);
xor U17441 (N_17441,N_15324,N_15416);
nor U17442 (N_17442,N_15496,N_15339);
nor U17443 (N_17443,N_16167,N_16112);
xnor U17444 (N_17444,N_15740,N_16036);
and U17445 (N_17445,N_15429,N_15311);
xor U17446 (N_17446,N_16078,N_15002);
nand U17447 (N_17447,N_16214,N_15606);
or U17448 (N_17448,N_16093,N_16221);
nor U17449 (N_17449,N_15067,N_15674);
nor U17450 (N_17450,N_15314,N_15066);
nor U17451 (N_17451,N_15712,N_15827);
nand U17452 (N_17452,N_15691,N_15070);
nand U17453 (N_17453,N_15361,N_15342);
nor U17454 (N_17454,N_15709,N_16081);
and U17455 (N_17455,N_15201,N_15069);
nand U17456 (N_17456,N_15739,N_15460);
and U17457 (N_17457,N_15906,N_15670);
or U17458 (N_17458,N_15054,N_16113);
nand U17459 (N_17459,N_15595,N_15269);
nor U17460 (N_17460,N_15111,N_15385);
nor U17461 (N_17461,N_16063,N_15636);
nand U17462 (N_17462,N_15391,N_15788);
nand U17463 (N_17463,N_15671,N_15839);
and U17464 (N_17464,N_16177,N_15362);
or U17465 (N_17465,N_15316,N_15198);
or U17466 (N_17466,N_15509,N_15123);
and U17467 (N_17467,N_15754,N_15646);
nand U17468 (N_17468,N_15107,N_15901);
and U17469 (N_17469,N_15903,N_15559);
nand U17470 (N_17470,N_16135,N_15371);
and U17471 (N_17471,N_15222,N_16003);
nor U17472 (N_17472,N_15009,N_15959);
xor U17473 (N_17473,N_15101,N_15587);
nand U17474 (N_17474,N_15874,N_15053);
nor U17475 (N_17475,N_16128,N_15115);
and U17476 (N_17476,N_15398,N_15479);
and U17477 (N_17477,N_15681,N_16059);
or U17478 (N_17478,N_15030,N_15726);
or U17479 (N_17479,N_15082,N_15931);
or U17480 (N_17480,N_15378,N_16221);
nand U17481 (N_17481,N_15697,N_16201);
and U17482 (N_17482,N_16052,N_15514);
nand U17483 (N_17483,N_15829,N_15124);
xnor U17484 (N_17484,N_15728,N_15602);
xor U17485 (N_17485,N_16056,N_15981);
and U17486 (N_17486,N_15797,N_16123);
xnor U17487 (N_17487,N_15663,N_15680);
xnor U17488 (N_17488,N_15583,N_15569);
or U17489 (N_17489,N_16248,N_15446);
nor U17490 (N_17490,N_16165,N_15252);
nand U17491 (N_17491,N_16113,N_16048);
and U17492 (N_17492,N_15084,N_15146);
and U17493 (N_17493,N_15691,N_16106);
or U17494 (N_17494,N_15065,N_15161);
and U17495 (N_17495,N_15583,N_15002);
or U17496 (N_17496,N_15746,N_15460);
nand U17497 (N_17497,N_15979,N_15234);
nor U17498 (N_17498,N_15541,N_16028);
and U17499 (N_17499,N_15230,N_16221);
or U17500 (N_17500,N_17258,N_17349);
or U17501 (N_17501,N_17365,N_16801);
and U17502 (N_17502,N_17462,N_16846);
nand U17503 (N_17503,N_17484,N_17239);
and U17504 (N_17504,N_16566,N_17392);
xnor U17505 (N_17505,N_17219,N_17480);
or U17506 (N_17506,N_16989,N_16759);
and U17507 (N_17507,N_17034,N_17256);
or U17508 (N_17508,N_16441,N_16769);
nor U17509 (N_17509,N_16406,N_16474);
nand U17510 (N_17510,N_16900,N_16520);
nand U17511 (N_17511,N_16516,N_16512);
and U17512 (N_17512,N_16903,N_17037);
nand U17513 (N_17513,N_17470,N_16673);
and U17514 (N_17514,N_17402,N_16352);
xor U17515 (N_17515,N_17001,N_17445);
and U17516 (N_17516,N_16944,N_17129);
nand U17517 (N_17517,N_16264,N_17060);
and U17518 (N_17518,N_16605,N_16467);
and U17519 (N_17519,N_17061,N_16997);
nand U17520 (N_17520,N_17430,N_17389);
nand U17521 (N_17521,N_16761,N_17393);
xor U17522 (N_17522,N_16282,N_16356);
or U17523 (N_17523,N_17083,N_16712);
nor U17524 (N_17524,N_16935,N_16483);
and U17525 (N_17525,N_16401,N_16511);
or U17526 (N_17526,N_17319,N_17420);
and U17527 (N_17527,N_16702,N_16598);
and U17528 (N_17528,N_16305,N_17082);
xnor U17529 (N_17529,N_17433,N_16921);
and U17530 (N_17530,N_16789,N_16945);
nor U17531 (N_17531,N_16841,N_16699);
nand U17532 (N_17532,N_16535,N_17472);
or U17533 (N_17533,N_16973,N_16528);
and U17534 (N_17534,N_16351,N_16650);
or U17535 (N_17535,N_17443,N_16951);
and U17536 (N_17536,N_16328,N_16400);
xor U17537 (N_17537,N_16440,N_17442);
nor U17538 (N_17538,N_16668,N_17459);
or U17539 (N_17539,N_17031,N_17407);
nor U17540 (N_17540,N_17355,N_16344);
and U17541 (N_17541,N_17321,N_17063);
nand U17542 (N_17542,N_17250,N_16901);
or U17543 (N_17543,N_16738,N_17202);
nor U17544 (N_17544,N_17141,N_16552);
or U17545 (N_17545,N_16860,N_16882);
nor U17546 (N_17546,N_17255,N_16251);
nor U17547 (N_17547,N_16695,N_17253);
and U17548 (N_17548,N_16827,N_16472);
xor U17549 (N_17549,N_16655,N_17376);
or U17550 (N_17550,N_16959,N_17434);
nand U17551 (N_17551,N_16659,N_17327);
nand U17552 (N_17552,N_17014,N_16775);
nand U17553 (N_17553,N_17095,N_17452);
or U17554 (N_17554,N_17068,N_16438);
nor U17555 (N_17555,N_16476,N_16275);
nor U17556 (N_17556,N_16749,N_16785);
xnor U17557 (N_17557,N_17481,N_17312);
and U17558 (N_17558,N_17271,N_16933);
and U17559 (N_17559,N_16631,N_17415);
nand U17560 (N_17560,N_16696,N_16479);
nand U17561 (N_17561,N_17294,N_17002);
and U17562 (N_17562,N_16286,N_17311);
nand U17563 (N_17563,N_17020,N_16326);
xor U17564 (N_17564,N_16355,N_16602);
xnor U17565 (N_17565,N_17118,N_16619);
nor U17566 (N_17566,N_16623,N_17336);
and U17567 (N_17567,N_16526,N_17309);
and U17568 (N_17568,N_17286,N_17266);
nor U17569 (N_17569,N_17328,N_17069);
nor U17570 (N_17570,N_16701,N_16430);
xnor U17571 (N_17571,N_16469,N_16728);
or U17572 (N_17572,N_16360,N_16622);
nand U17573 (N_17573,N_17025,N_16947);
xnor U17574 (N_17574,N_16980,N_17013);
xor U17575 (N_17575,N_17230,N_17302);
or U17576 (N_17576,N_16966,N_17399);
and U17577 (N_17577,N_16490,N_16575);
xor U17578 (N_17578,N_17164,N_16839);
xor U17579 (N_17579,N_17058,N_16875);
and U17580 (N_17580,N_16791,N_17485);
nor U17581 (N_17581,N_16744,N_17425);
or U17582 (N_17582,N_16859,N_17085);
and U17583 (N_17583,N_16589,N_16250);
xnor U17584 (N_17584,N_16455,N_16502);
xor U17585 (N_17585,N_16804,N_17026);
xor U17586 (N_17586,N_17391,N_16273);
and U17587 (N_17587,N_16606,N_17173);
xor U17588 (N_17588,N_17306,N_16307);
or U17589 (N_17589,N_17201,N_17176);
xor U17590 (N_17590,N_16818,N_16869);
xor U17591 (N_17591,N_16703,N_16942);
or U17592 (N_17592,N_17215,N_17358);
xor U17593 (N_17593,N_16564,N_16928);
and U17594 (N_17594,N_16965,N_17172);
or U17595 (N_17595,N_17424,N_16465);
nor U17596 (N_17596,N_16770,N_16887);
nand U17597 (N_17597,N_16613,N_17222);
xnor U17598 (N_17598,N_16266,N_16379);
nand U17599 (N_17599,N_16601,N_16932);
nand U17600 (N_17600,N_16724,N_17496);
nand U17601 (N_17601,N_16862,N_16337);
xnor U17602 (N_17602,N_16847,N_16995);
xor U17603 (N_17603,N_17439,N_17388);
xor U17604 (N_17604,N_17130,N_16988);
and U17605 (N_17605,N_16544,N_17205);
nor U17606 (N_17606,N_16506,N_17438);
and U17607 (N_17607,N_16260,N_17211);
nand U17608 (N_17608,N_16676,N_16413);
nand U17609 (N_17609,N_16281,N_17143);
nand U17610 (N_17610,N_16393,N_17251);
and U17611 (N_17611,N_17482,N_16905);
or U17612 (N_17612,N_17366,N_16717);
or U17613 (N_17613,N_16332,N_17423);
xor U17614 (N_17614,N_16309,N_16704);
xnor U17615 (N_17615,N_16718,N_16715);
or U17616 (N_17616,N_17383,N_17346);
nand U17617 (N_17617,N_16664,N_17120);
nor U17618 (N_17618,N_16462,N_16559);
nand U17619 (N_17619,N_16481,N_16808);
nand U17620 (N_17620,N_17209,N_16291);
nor U17621 (N_17621,N_16262,N_16886);
or U17622 (N_17622,N_16579,N_17107);
nor U17623 (N_17623,N_16641,N_17494);
nor U17624 (N_17624,N_16920,N_16913);
nand U17625 (N_17625,N_16384,N_17006);
and U17626 (N_17626,N_16364,N_16873);
xor U17627 (N_17627,N_16371,N_16614);
xnor U17628 (N_17628,N_16957,N_16568);
nand U17629 (N_17629,N_17027,N_16625);
or U17630 (N_17630,N_16346,N_17186);
or U17631 (N_17631,N_16572,N_16555);
nand U17632 (N_17632,N_17320,N_16357);
nor U17633 (N_17633,N_16505,N_16359);
or U17634 (N_17634,N_17090,N_16633);
nand U17635 (N_17635,N_16743,N_17374);
or U17636 (N_17636,N_16970,N_17204);
xor U17637 (N_17637,N_16493,N_16587);
and U17638 (N_17638,N_16689,N_17275);
nor U17639 (N_17639,N_16537,N_16259);
nand U17640 (N_17640,N_16842,N_16972);
or U17641 (N_17641,N_17300,N_17023);
nor U17642 (N_17642,N_16377,N_16964);
xor U17643 (N_17643,N_16720,N_17183);
xor U17644 (N_17644,N_16542,N_16786);
and U17645 (N_17645,N_17017,N_16848);
xnor U17646 (N_17646,N_16381,N_17162);
nor U17647 (N_17647,N_17228,N_17322);
nor U17648 (N_17648,N_16644,N_16652);
nand U17649 (N_17649,N_16853,N_16949);
nand U17650 (N_17650,N_16603,N_17166);
xor U17651 (N_17651,N_17193,N_17436);
xnor U17652 (N_17652,N_17435,N_17267);
nor U17653 (N_17653,N_17140,N_17054);
or U17654 (N_17654,N_16557,N_17105);
xnor U17655 (N_17655,N_16727,N_16297);
nor U17656 (N_17656,N_16278,N_16663);
and U17657 (N_17657,N_17015,N_16308);
xnor U17658 (N_17658,N_17032,N_16313);
and U17659 (N_17659,N_17421,N_17282);
nor U17660 (N_17660,N_16856,N_16496);
or U17661 (N_17661,N_17345,N_17313);
or U17662 (N_17662,N_16803,N_16434);
and U17663 (N_17663,N_16926,N_16287);
or U17664 (N_17664,N_16939,N_17078);
xnor U17665 (N_17665,N_16794,N_16924);
nand U17666 (N_17666,N_16560,N_17064);
or U17667 (N_17667,N_17053,N_17160);
nor U17668 (N_17668,N_16312,N_16647);
xor U17669 (N_17669,N_16651,N_17021);
nor U17670 (N_17670,N_16283,N_17299);
nor U17671 (N_17671,N_17126,N_17127);
xor U17672 (N_17672,N_17348,N_16363);
nand U17673 (N_17673,N_16253,N_16817);
or U17674 (N_17674,N_17367,N_16883);
or U17675 (N_17675,N_17122,N_16333);
nor U17676 (N_17676,N_16661,N_16914);
and U17677 (N_17677,N_17397,N_17454);
and U17678 (N_17678,N_16551,N_17416);
and U17679 (N_17679,N_17229,N_16675);
nor U17680 (N_17680,N_17281,N_17161);
and U17681 (N_17681,N_17136,N_17088);
nand U17682 (N_17682,N_16783,N_17288);
nor U17683 (N_17683,N_17177,N_16398);
and U17684 (N_17684,N_17012,N_16854);
or U17685 (N_17685,N_17226,N_16806);
nor U17686 (N_17686,N_16936,N_16709);
nor U17687 (N_17687,N_16721,N_17360);
xor U17688 (N_17688,N_16310,N_17331);
and U17689 (N_17689,N_16289,N_17351);
nand U17690 (N_17690,N_16279,N_17035);
or U17691 (N_17691,N_16658,N_17379);
nor U17692 (N_17692,N_16338,N_17075);
nor U17693 (N_17693,N_17451,N_16762);
or U17694 (N_17694,N_16742,N_17181);
nand U17695 (N_17695,N_16684,N_16265);
and U17696 (N_17696,N_17106,N_17314);
or U17697 (N_17697,N_16495,N_16778);
or U17698 (N_17698,N_16958,N_17487);
nor U17699 (N_17699,N_16261,N_17466);
or U17700 (N_17700,N_16909,N_16284);
nand U17701 (N_17701,N_16732,N_17332);
xnor U17702 (N_17702,N_16577,N_17269);
nor U17703 (N_17703,N_16953,N_16318);
and U17704 (N_17704,N_16439,N_16811);
and U17705 (N_17705,N_16437,N_16594);
and U17706 (N_17706,N_17398,N_17432);
nor U17707 (N_17707,N_16876,N_17469);
xor U17708 (N_17708,N_16776,N_16864);
and U17709 (N_17709,N_17038,N_17401);
and U17710 (N_17710,N_16304,N_16447);
or U17711 (N_17711,N_16532,N_17386);
nor U17712 (N_17712,N_16740,N_16303);
and U17713 (N_17713,N_17489,N_16501);
and U17714 (N_17714,N_16697,N_16630);
nand U17715 (N_17715,N_16531,N_17493);
nand U17716 (N_17716,N_16375,N_16489);
nand U17717 (N_17717,N_17184,N_16435);
xor U17718 (N_17718,N_16380,N_17121);
nand U17719 (N_17719,N_17235,N_17133);
xor U17720 (N_17720,N_16763,N_16402);
xor U17721 (N_17721,N_16576,N_16518);
nor U17722 (N_17722,N_16581,N_16367);
or U17723 (N_17723,N_17352,N_16960);
and U17724 (N_17724,N_16979,N_16460);
and U17725 (N_17725,N_16617,N_17403);
and U17726 (N_17726,N_16996,N_16394);
xnor U17727 (N_17727,N_16342,N_16331);
xnor U17728 (N_17728,N_17124,N_16475);
nor U17729 (N_17729,N_16399,N_16832);
and U17730 (N_17730,N_17047,N_16632);
xnor U17731 (N_17731,N_17317,N_16492);
or U17732 (N_17732,N_16971,N_17243);
nand U17733 (N_17733,N_17040,N_16396);
and U17734 (N_17734,N_16376,N_16523);
nor U17735 (N_17735,N_16730,N_17216);
nand U17736 (N_17736,N_16975,N_16741);
or U17737 (N_17737,N_16277,N_16865);
or U17738 (N_17738,N_16923,N_16897);
and U17739 (N_17739,N_17033,N_16896);
nand U17740 (N_17740,N_16565,N_16588);
nor U17741 (N_17741,N_17467,N_16403);
nand U17742 (N_17742,N_17149,N_16772);
nand U17743 (N_17743,N_17298,N_17057);
xor U17744 (N_17744,N_16777,N_16610);
or U17745 (N_17745,N_17241,N_17237);
and U17746 (N_17746,N_16295,N_17394);
or U17747 (N_17747,N_17465,N_17463);
nand U17748 (N_17748,N_17297,N_16828);
xnor U17749 (N_17749,N_17108,N_17076);
nand U17750 (N_17750,N_16522,N_16509);
and U17751 (N_17751,N_16692,N_16986);
or U17752 (N_17752,N_16654,N_16754);
xor U17753 (N_17753,N_16497,N_16358);
and U17754 (N_17754,N_16733,N_17029);
nand U17755 (N_17755,N_17159,N_16993);
nor U17756 (N_17756,N_16934,N_17052);
or U17757 (N_17757,N_16851,N_17024);
nor U17758 (N_17758,N_16863,N_16368);
nand U17759 (N_17759,N_17059,N_16391);
xnor U17760 (N_17760,N_16317,N_16288);
nor U17761 (N_17761,N_17390,N_17084);
and U17762 (N_17762,N_17418,N_16274);
and U17763 (N_17763,N_17370,N_17200);
nand U17764 (N_17764,N_16653,N_17431);
nand U17765 (N_17765,N_17158,N_16477);
nor U17766 (N_17766,N_17110,N_17016);
nand U17767 (N_17767,N_17169,N_16764);
nor U17768 (N_17768,N_16524,N_17384);
or U17769 (N_17769,N_16722,N_17203);
nor U17770 (N_17770,N_17338,N_16758);
or U17771 (N_17771,N_17499,N_17174);
nand U17772 (N_17772,N_16634,N_17307);
xnor U17773 (N_17773,N_16950,N_16411);
xor U17774 (N_17774,N_17214,N_16713);
xor U17775 (N_17775,N_16417,N_16629);
and U17776 (N_17776,N_16280,N_16795);
xnor U17777 (N_17777,N_16812,N_16790);
xnor U17778 (N_17778,N_17363,N_16272);
and U17779 (N_17779,N_17139,N_17460);
xnor U17780 (N_17780,N_16824,N_17100);
or U17781 (N_17781,N_17233,N_17097);
nand U17782 (N_17782,N_17457,N_16955);
xor U17783 (N_17783,N_17483,N_17019);
xor U17784 (N_17784,N_17030,N_16624);
nand U17785 (N_17785,N_17491,N_17427);
nor U17786 (N_17786,N_16731,N_17206);
or U17787 (N_17787,N_17111,N_16574);
and U17788 (N_17788,N_16880,N_16292);
nor U17789 (N_17789,N_17180,N_16395);
nor U17790 (N_17790,N_16729,N_17217);
nor U17791 (N_17791,N_16919,N_16327);
and U17792 (N_17792,N_16604,N_16814);
nor U17793 (N_17793,N_16451,N_16482);
xnor U17794 (N_17794,N_17213,N_16685);
and U17795 (N_17795,N_16878,N_16719);
nor U17796 (N_17796,N_16940,N_16334);
and U17797 (N_17797,N_16750,N_17109);
or U17798 (N_17798,N_17380,N_16500);
nand U17799 (N_17799,N_16657,N_16449);
or U17800 (N_17800,N_17179,N_16616);
nand U17801 (N_17801,N_16445,N_16627);
nand U17802 (N_17802,N_16825,N_17244);
nand U17803 (N_17803,N_16872,N_16840);
nand U17804 (N_17804,N_16311,N_16938);
and U17805 (N_17805,N_17155,N_17151);
or U17806 (N_17806,N_16388,N_16299);
nand U17807 (N_17807,N_16888,N_17357);
or U17808 (N_17808,N_16885,N_16499);
xor U17809 (N_17809,N_16454,N_17458);
or U17810 (N_17810,N_17410,N_16548);
nor U17811 (N_17811,N_17197,N_17000);
nor U17812 (N_17812,N_16507,N_16609);
nor U17813 (N_17813,N_17198,N_16267);
nor U17814 (N_17814,N_16366,N_16365);
nor U17815 (N_17815,N_16683,N_16466);
nand U17816 (N_17816,N_16612,N_17188);
and U17817 (N_17817,N_17498,N_17448);
or U17818 (N_17818,N_16582,N_16670);
and U17819 (N_17819,N_17042,N_16912);
nor U17820 (N_17820,N_16766,N_17028);
nor U17821 (N_17821,N_16826,N_16443);
or U17822 (N_17822,N_17131,N_17242);
or U17823 (N_17823,N_16679,N_16792);
and U17824 (N_17824,N_16714,N_17134);
or U17825 (N_17825,N_16855,N_16788);
xnor U17826 (N_17826,N_16301,N_16322);
nor U17827 (N_17827,N_17453,N_17150);
xnor U17828 (N_17828,N_17412,N_16590);
and U17829 (N_17829,N_17007,N_17074);
or U17830 (N_17830,N_16407,N_16674);
and U17831 (N_17831,N_16640,N_17417);
and U17832 (N_17832,N_17208,N_17265);
nand U17833 (N_17833,N_17289,N_16665);
and U17834 (N_17834,N_16941,N_16831);
and U17835 (N_17835,N_16908,N_16597);
xor U17836 (N_17836,N_16796,N_17167);
xor U17837 (N_17837,N_17456,N_17284);
and U17838 (N_17838,N_17210,N_16271);
or U17839 (N_17839,N_16906,N_16892);
and U17840 (N_17840,N_17187,N_17277);
nor U17841 (N_17841,N_17165,N_16992);
nor U17842 (N_17842,N_17369,N_16488);
xor U17843 (N_17843,N_16436,N_17375);
nor U17844 (N_17844,N_16444,N_17046);
or U17845 (N_17845,N_17192,N_17147);
nor U17846 (N_17846,N_17062,N_17333);
or U17847 (N_17847,N_16821,N_17245);
nand U17848 (N_17848,N_16561,N_16829);
nand U17849 (N_17849,N_17372,N_16263);
nand U17850 (N_17850,N_17236,N_16768);
or U17851 (N_17851,N_17171,N_16752);
nand U17852 (N_17852,N_16751,N_16527);
and U17853 (N_17853,N_16793,N_17497);
nand U17854 (N_17854,N_16536,N_16756);
or U17855 (N_17855,N_16898,N_16484);
or U17856 (N_17856,N_16723,N_16525);
or U17857 (N_17857,N_17293,N_16450);
nand U17858 (N_17858,N_17194,N_16943);
xor U17859 (N_17859,N_17094,N_16296);
nor U17860 (N_17860,N_16463,N_16866);
xor U17861 (N_17861,N_16563,N_17305);
or U17862 (N_17862,N_16420,N_16845);
or U17863 (N_17863,N_17157,N_16690);
nor U17864 (N_17864,N_16370,N_17295);
xnor U17865 (N_17865,N_16990,N_17036);
nand U17866 (N_17866,N_16642,N_17422);
and U17867 (N_17867,N_16553,N_17447);
nor U17868 (N_17868,N_16343,N_16387);
and U17869 (N_17869,N_16468,N_16349);
nor U17870 (N_17870,N_17310,N_17290);
nor U17871 (N_17871,N_17444,N_17099);
nor U17872 (N_17872,N_16546,N_16646);
or U17873 (N_17873,N_16890,N_16779);
nand U17874 (N_17874,N_16968,N_16969);
nand U17875 (N_17875,N_16857,N_16416);
nand U17876 (N_17876,N_17406,N_16998);
nand U17877 (N_17877,N_17359,N_16494);
nor U17878 (N_17878,N_17249,N_16877);
xnor U17879 (N_17879,N_17079,N_17071);
nor U17880 (N_17880,N_17170,N_16929);
nand U17881 (N_17881,N_16256,N_17404);
and U17882 (N_17882,N_17223,N_16294);
and U17883 (N_17883,N_17315,N_16432);
xor U17884 (N_17884,N_16583,N_17257);
xor U17885 (N_17885,N_16615,N_16600);
xnor U17886 (N_17886,N_16409,N_17009);
or U17887 (N_17887,N_17381,N_16671);
and U17888 (N_17888,N_17091,N_16879);
nand U17889 (N_17889,N_16907,N_16765);
xnor U17890 (N_17890,N_17081,N_17207);
and U17891 (N_17891,N_16910,N_17154);
nand U17892 (N_17892,N_16948,N_16805);
or U17893 (N_17893,N_16822,N_17276);
nor U17894 (N_17894,N_17220,N_17148);
or U17895 (N_17895,N_16554,N_16798);
nor U17896 (N_17896,N_17405,N_17478);
and U17897 (N_17897,N_17440,N_16480);
xor U17898 (N_17898,N_17087,N_16385);
xnor U17899 (N_17899,N_16858,N_16666);
nand U17900 (N_17900,N_16611,N_16823);
nand U17901 (N_17901,N_16956,N_17373);
and U17902 (N_17902,N_17318,N_16620);
and U17903 (N_17903,N_16835,N_16471);
and U17904 (N_17904,N_16425,N_16636);
and U17905 (N_17905,N_16347,N_16362);
or U17906 (N_17906,N_16556,N_16735);
or U17907 (N_17907,N_17382,N_17343);
or U17908 (N_17908,N_17005,N_16787);
or U17909 (N_17909,N_17261,N_17128);
nor U17910 (N_17910,N_16503,N_16491);
nand U17911 (N_17911,N_17051,N_16498);
nor U17912 (N_17912,N_16739,N_17231);
and U17913 (N_17913,N_17304,N_16392);
and U17914 (N_17914,N_17329,N_16874);
nand U17915 (N_17915,N_17114,N_17341);
and U17916 (N_17916,N_17125,N_16335);
and U17917 (N_17917,N_17175,N_16421);
nor U17918 (N_17918,N_16915,N_16660);
xnor U17919 (N_17919,N_17010,N_16911);
nand U17920 (N_17920,N_16963,N_17342);
xor U17921 (N_17921,N_16771,N_17003);
nor U17922 (N_17922,N_17093,N_16747);
nand U17923 (N_17923,N_16974,N_16538);
xor U17924 (N_17924,N_16345,N_17490);
xnor U17925 (N_17925,N_16290,N_16889);
nand U17926 (N_17926,N_16596,N_17495);
and U17927 (N_17927,N_16987,N_16374);
and U17928 (N_17928,N_17378,N_16734);
nand U17929 (N_17929,N_17263,N_16639);
xor U17930 (N_17930,N_17279,N_17153);
xnor U17931 (N_17931,N_17104,N_17476);
nor U17932 (N_17932,N_17011,N_16737);
nor U17933 (N_17933,N_16255,N_16849);
xnor U17934 (N_17934,N_17224,N_16530);
or U17935 (N_17935,N_16962,N_16424);
xor U17936 (N_17936,N_17191,N_16431);
nand U17937 (N_17937,N_16706,N_16780);
nand U17938 (N_17938,N_17098,N_17185);
or U17939 (N_17939,N_16784,N_16843);
nand U17940 (N_17940,N_17248,N_16781);
nand U17941 (N_17941,N_17117,N_16810);
nor U17942 (N_17942,N_16270,N_16807);
or U17943 (N_17943,N_16545,N_16994);
nand U17944 (N_17944,N_16700,N_17419);
and U17945 (N_17945,N_17004,N_17112);
and U17946 (N_17946,N_16461,N_16984);
or U17947 (N_17947,N_16871,N_16599);
xnor U17948 (N_17948,N_16918,N_16300);
and U17949 (N_17949,N_16446,N_17137);
or U17950 (N_17950,N_16946,N_16837);
and U17951 (N_17951,N_16412,N_16894);
nand U17952 (N_17952,N_16645,N_16677);
or U17953 (N_17953,N_16844,N_16961);
nor U17954 (N_17954,N_16580,N_16442);
and U17955 (N_17955,N_16931,N_17273);
xnor U17956 (N_17956,N_16422,N_17232);
nand U17957 (N_17957,N_16904,N_16694);
or U17958 (N_17958,N_17070,N_17272);
and U17959 (N_17959,N_16578,N_16504);
and U17960 (N_17960,N_17471,N_16452);
nor U17961 (N_17961,N_17450,N_16513);
nor U17962 (N_17962,N_16453,N_16314);
nor U17963 (N_17963,N_17252,N_17486);
xnor U17964 (N_17964,N_17377,N_17168);
nand U17965 (N_17965,N_16638,N_16382);
or U17966 (N_17966,N_16927,N_17285);
and U17967 (N_17967,N_17195,N_16608);
nand U17968 (N_17968,N_16725,N_16868);
nand U17969 (N_17969,N_17326,N_16426);
nand U17970 (N_17970,N_16833,N_17218);
nand U17971 (N_17971,N_16571,N_16348);
xnor U17972 (N_17972,N_16514,N_16967);
nor U17973 (N_17973,N_16649,N_16405);
xor U17974 (N_17974,N_17283,N_17247);
or U17975 (N_17975,N_16298,N_16850);
nor U17976 (N_17976,N_16473,N_17429);
or U17977 (N_17977,N_16410,N_16954);
and U17978 (N_17978,N_16350,N_16628);
nand U17979 (N_17979,N_16378,N_16643);
or U17980 (N_17980,N_17400,N_16325);
nand U17981 (N_17981,N_16820,N_16541);
or U17982 (N_17982,N_16558,N_17437);
nor U17983 (N_17983,N_16285,N_17492);
nor U17984 (N_17984,N_16427,N_16711);
or U17985 (N_17985,N_17190,N_16891);
nand U17986 (N_17986,N_16316,N_16459);
or U17987 (N_17987,N_17103,N_16293);
and U17988 (N_17988,N_16448,N_16419);
and U17989 (N_17989,N_16517,N_16428);
xor U17990 (N_17990,N_17262,N_17474);
xnor U17991 (N_17991,N_16534,N_17396);
and U17992 (N_17992,N_17385,N_16258);
nand U17993 (N_17993,N_17182,N_16329);
and U17994 (N_17994,N_16917,N_16925);
or U17995 (N_17995,N_17361,N_17387);
or U17996 (N_17996,N_17479,N_16302);
nor U17997 (N_17997,N_16930,N_17050);
xor U17998 (N_17998,N_17145,N_16802);
nor U17999 (N_17999,N_17268,N_16315);
and U18000 (N_18000,N_17146,N_17337);
and U18001 (N_18001,N_16753,N_16852);
xor U18002 (N_18002,N_16457,N_17344);
and U18003 (N_18003,N_16767,N_17196);
and U18004 (N_18004,N_16681,N_17354);
xnor U18005 (N_18005,N_17408,N_16306);
or U18006 (N_18006,N_16339,N_16543);
nand U18007 (N_18007,N_16341,N_17323);
xor U18008 (N_18008,N_16487,N_16815);
nor U18009 (N_18009,N_16937,N_17189);
nor U18010 (N_18010,N_16521,N_16757);
or U18011 (N_18011,N_17072,N_16895);
nor U18012 (N_18012,N_17475,N_16745);
xnor U18013 (N_18013,N_16710,N_16688);
nor U18014 (N_18014,N_17234,N_17259);
or U18015 (N_18015,N_16404,N_17362);
or U18016 (N_18016,N_17449,N_17411);
xnor U18017 (N_18017,N_16867,N_16705);
nand U18018 (N_18018,N_16648,N_16321);
or U18019 (N_18019,N_16797,N_17364);
nand U18020 (N_18020,N_17080,N_17246);
and U18021 (N_18021,N_16607,N_17339);
xnor U18022 (N_18022,N_16952,N_17488);
nand U18023 (N_18023,N_17056,N_17055);
nor U18024 (N_18024,N_17101,N_17067);
nand U18025 (N_18025,N_16870,N_16257);
nor U18026 (N_18026,N_16626,N_16716);
xnor U18027 (N_18027,N_16830,N_16397);
nor U18028 (N_18028,N_16893,N_16976);
nand U18029 (N_18029,N_16336,N_17163);
xnor U18030 (N_18030,N_17240,N_16458);
nor U18031 (N_18031,N_16773,N_17347);
nor U18032 (N_18032,N_16585,N_16669);
or U18033 (N_18033,N_16637,N_16423);
or U18034 (N_18034,N_16977,N_17119);
or U18035 (N_18035,N_17303,N_17092);
or U18036 (N_18036,N_17086,N_16414);
and U18037 (N_18037,N_16621,N_17044);
or U18038 (N_18038,N_16922,N_16760);
nand U18039 (N_18039,N_16884,N_16429);
xnor U18040 (N_18040,N_17371,N_16678);
nand U18041 (N_18041,N_16748,N_16508);
and U18042 (N_18042,N_16361,N_16510);
nor U18043 (N_18043,N_17225,N_16902);
or U18044 (N_18044,N_17264,N_17018);
nor U18045 (N_18045,N_16515,N_16635);
xnor U18046 (N_18046,N_17041,N_17464);
xor U18047 (N_18047,N_16320,N_17446);
nor U18048 (N_18048,N_17287,N_17102);
and U18049 (N_18049,N_16464,N_17008);
nand U18050 (N_18050,N_16667,N_16680);
nand U18051 (N_18051,N_16570,N_17043);
nor U18052 (N_18052,N_17132,N_17049);
nor U18053 (N_18053,N_17113,N_16708);
or U18054 (N_18054,N_16586,N_16591);
xnor U18055 (N_18055,N_16595,N_16816);
xnor U18056 (N_18056,N_16687,N_17308);
and U18057 (N_18057,N_16573,N_16593);
nor U18058 (N_18058,N_17270,N_17089);
nand U18059 (N_18059,N_17325,N_17212);
and U18060 (N_18060,N_16836,N_16478);
nand U18061 (N_18061,N_17156,N_16899);
nand U18062 (N_18062,N_16549,N_17334);
and U18063 (N_18063,N_16369,N_17221);
and U18064 (N_18064,N_16529,N_16383);
or U18065 (N_18065,N_17274,N_16656);
and U18066 (N_18066,N_16319,N_16562);
nor U18067 (N_18067,N_16470,N_16340);
nor U18068 (N_18068,N_16691,N_16372);
xnor U18069 (N_18069,N_16418,N_17368);
and U18070 (N_18070,N_16539,N_17340);
nand U18071 (N_18071,N_16799,N_17178);
or U18072 (N_18072,N_16415,N_16800);
or U18073 (N_18073,N_16486,N_17350);
and U18074 (N_18074,N_16276,N_17426);
nand U18075 (N_18075,N_16693,N_16456);
or U18076 (N_18076,N_16540,N_17335);
or U18077 (N_18077,N_16861,N_16682);
or U18078 (N_18078,N_17142,N_16707);
nor U18079 (N_18079,N_16755,N_16323);
nor U18080 (N_18080,N_16991,N_17353);
and U18081 (N_18081,N_16547,N_16252);
nor U18082 (N_18082,N_17039,N_16834);
nor U18083 (N_18083,N_17292,N_16354);
xor U18084 (N_18084,N_17441,N_16698);
or U18085 (N_18085,N_16269,N_17301);
or U18086 (N_18086,N_17227,N_16519);
and U18087 (N_18087,N_17073,N_17414);
nor U18088 (N_18088,N_16736,N_16386);
or U18089 (N_18089,N_16838,N_16782);
nor U18090 (N_18090,N_16672,N_17066);
and U18091 (N_18091,N_17123,N_17280);
or U18092 (N_18092,N_16881,N_16983);
xor U18093 (N_18093,N_16268,N_17395);
nand U18094 (N_18094,N_16533,N_16254);
and U18095 (N_18095,N_17428,N_16584);
and U18096 (N_18096,N_16999,N_17144);
xor U18097 (N_18097,N_16618,N_16389);
and U18098 (N_18098,N_16686,N_17477);
or U18099 (N_18099,N_17455,N_17135);
nand U18100 (N_18100,N_16550,N_16982);
or U18101 (N_18101,N_16485,N_17116);
nor U18102 (N_18102,N_16324,N_17096);
and U18103 (N_18103,N_16433,N_16746);
nand U18104 (N_18104,N_17077,N_17296);
or U18105 (N_18105,N_16978,N_16390);
or U18106 (N_18106,N_17291,N_17115);
or U18107 (N_18107,N_16819,N_17022);
xor U18108 (N_18108,N_16373,N_17473);
nor U18109 (N_18109,N_17199,N_16567);
and U18110 (N_18110,N_16916,N_16774);
nor U18111 (N_18111,N_17152,N_16353);
xnor U18112 (N_18112,N_17238,N_16569);
nor U18113 (N_18113,N_17468,N_16813);
xnor U18114 (N_18114,N_17260,N_17324);
or U18115 (N_18115,N_16592,N_17254);
or U18116 (N_18116,N_16662,N_17409);
nor U18117 (N_18117,N_17316,N_17461);
nor U18118 (N_18118,N_16726,N_16330);
xnor U18119 (N_18119,N_16985,N_17330);
and U18120 (N_18120,N_17356,N_16981);
nor U18121 (N_18121,N_17138,N_16809);
xnor U18122 (N_18122,N_17045,N_17413);
xnor U18123 (N_18123,N_17278,N_17048);
and U18124 (N_18124,N_17065,N_16408);
nor U18125 (N_18125,N_16554,N_16300);
and U18126 (N_18126,N_17001,N_16553);
nor U18127 (N_18127,N_16525,N_17072);
nor U18128 (N_18128,N_16610,N_16824);
nor U18129 (N_18129,N_16736,N_16963);
nand U18130 (N_18130,N_17426,N_17307);
nand U18131 (N_18131,N_17197,N_17313);
and U18132 (N_18132,N_17241,N_16689);
nor U18133 (N_18133,N_16887,N_17276);
or U18134 (N_18134,N_16619,N_16583);
nor U18135 (N_18135,N_17017,N_17443);
nor U18136 (N_18136,N_17417,N_16569);
and U18137 (N_18137,N_16715,N_16654);
nand U18138 (N_18138,N_16653,N_17371);
xor U18139 (N_18139,N_16715,N_16348);
xnor U18140 (N_18140,N_17223,N_17114);
or U18141 (N_18141,N_17299,N_17417);
and U18142 (N_18142,N_16866,N_17054);
or U18143 (N_18143,N_16396,N_17114);
xor U18144 (N_18144,N_16451,N_16347);
nand U18145 (N_18145,N_17327,N_16354);
and U18146 (N_18146,N_17145,N_17133);
or U18147 (N_18147,N_17419,N_16395);
or U18148 (N_18148,N_16507,N_16877);
xor U18149 (N_18149,N_16454,N_16391);
xnor U18150 (N_18150,N_17431,N_17492);
nand U18151 (N_18151,N_16330,N_16306);
xnor U18152 (N_18152,N_16254,N_16753);
nand U18153 (N_18153,N_16565,N_17199);
nor U18154 (N_18154,N_16773,N_17273);
and U18155 (N_18155,N_16436,N_17320);
xor U18156 (N_18156,N_16875,N_17235);
and U18157 (N_18157,N_16780,N_17218);
xnor U18158 (N_18158,N_16767,N_17162);
nor U18159 (N_18159,N_17113,N_16865);
nor U18160 (N_18160,N_17084,N_16865);
nand U18161 (N_18161,N_16995,N_17357);
or U18162 (N_18162,N_16836,N_17128);
nor U18163 (N_18163,N_16431,N_16338);
nand U18164 (N_18164,N_17086,N_16483);
or U18165 (N_18165,N_16714,N_17299);
nor U18166 (N_18166,N_17388,N_16531);
nor U18167 (N_18167,N_16717,N_16332);
nand U18168 (N_18168,N_16263,N_17294);
and U18169 (N_18169,N_17334,N_16398);
nor U18170 (N_18170,N_16361,N_17098);
and U18171 (N_18171,N_16586,N_16583);
nor U18172 (N_18172,N_16461,N_17302);
xnor U18173 (N_18173,N_17306,N_17172);
or U18174 (N_18174,N_16625,N_16705);
nand U18175 (N_18175,N_16339,N_17293);
nor U18176 (N_18176,N_16783,N_16272);
and U18177 (N_18177,N_17290,N_16694);
and U18178 (N_18178,N_16583,N_17490);
nor U18179 (N_18179,N_17219,N_17234);
nand U18180 (N_18180,N_17444,N_17403);
xor U18181 (N_18181,N_17456,N_16514);
nor U18182 (N_18182,N_17012,N_16458);
or U18183 (N_18183,N_17210,N_16535);
nor U18184 (N_18184,N_16461,N_16436);
or U18185 (N_18185,N_16993,N_16912);
nor U18186 (N_18186,N_17222,N_16884);
xor U18187 (N_18187,N_17144,N_16948);
or U18188 (N_18188,N_17377,N_17436);
nand U18189 (N_18189,N_16734,N_17453);
nor U18190 (N_18190,N_17159,N_17427);
nor U18191 (N_18191,N_16589,N_17310);
nor U18192 (N_18192,N_16471,N_17156);
nor U18193 (N_18193,N_16824,N_16700);
nand U18194 (N_18194,N_16268,N_16488);
or U18195 (N_18195,N_16654,N_17046);
nor U18196 (N_18196,N_16283,N_17091);
nor U18197 (N_18197,N_16868,N_16408);
and U18198 (N_18198,N_16348,N_16801);
xnor U18199 (N_18199,N_16380,N_17155);
or U18200 (N_18200,N_16735,N_16483);
nand U18201 (N_18201,N_16991,N_16785);
and U18202 (N_18202,N_17051,N_16749);
nor U18203 (N_18203,N_16936,N_17145);
and U18204 (N_18204,N_16994,N_16378);
and U18205 (N_18205,N_16423,N_17170);
nand U18206 (N_18206,N_17170,N_16443);
xor U18207 (N_18207,N_17179,N_16833);
nor U18208 (N_18208,N_16384,N_17203);
or U18209 (N_18209,N_17281,N_16343);
and U18210 (N_18210,N_16506,N_17297);
xnor U18211 (N_18211,N_17014,N_17008);
nor U18212 (N_18212,N_16950,N_17363);
or U18213 (N_18213,N_16431,N_17426);
xor U18214 (N_18214,N_17120,N_17447);
xnor U18215 (N_18215,N_17428,N_16409);
nor U18216 (N_18216,N_17453,N_16639);
nand U18217 (N_18217,N_17269,N_17101);
and U18218 (N_18218,N_16772,N_16400);
xor U18219 (N_18219,N_16565,N_17131);
or U18220 (N_18220,N_16344,N_17344);
and U18221 (N_18221,N_17003,N_16779);
or U18222 (N_18222,N_16607,N_17319);
xnor U18223 (N_18223,N_16275,N_16879);
xor U18224 (N_18224,N_16895,N_16290);
xor U18225 (N_18225,N_16902,N_16601);
and U18226 (N_18226,N_16961,N_16525);
and U18227 (N_18227,N_17257,N_17076);
and U18228 (N_18228,N_17240,N_16894);
nand U18229 (N_18229,N_16455,N_16774);
or U18230 (N_18230,N_16817,N_16998);
xor U18231 (N_18231,N_16521,N_17395);
and U18232 (N_18232,N_16968,N_17299);
or U18233 (N_18233,N_17385,N_16811);
nor U18234 (N_18234,N_17339,N_17114);
xor U18235 (N_18235,N_17125,N_17361);
nand U18236 (N_18236,N_16987,N_16764);
nand U18237 (N_18237,N_17386,N_16986);
and U18238 (N_18238,N_16491,N_16259);
nor U18239 (N_18239,N_17114,N_17408);
nor U18240 (N_18240,N_17129,N_16685);
and U18241 (N_18241,N_17332,N_16932);
and U18242 (N_18242,N_16281,N_17243);
and U18243 (N_18243,N_17475,N_16608);
or U18244 (N_18244,N_16622,N_16692);
nand U18245 (N_18245,N_16308,N_17213);
and U18246 (N_18246,N_17499,N_17113);
or U18247 (N_18247,N_16474,N_16570);
nand U18248 (N_18248,N_16275,N_17129);
nor U18249 (N_18249,N_16997,N_16891);
nand U18250 (N_18250,N_17104,N_16357);
and U18251 (N_18251,N_17477,N_16464);
nor U18252 (N_18252,N_16907,N_16596);
and U18253 (N_18253,N_16800,N_17119);
or U18254 (N_18254,N_17140,N_16819);
and U18255 (N_18255,N_16517,N_17064);
xor U18256 (N_18256,N_17315,N_16871);
nand U18257 (N_18257,N_16250,N_16363);
or U18258 (N_18258,N_16906,N_17388);
nor U18259 (N_18259,N_16658,N_17117);
and U18260 (N_18260,N_17497,N_17016);
nor U18261 (N_18261,N_17435,N_17231);
and U18262 (N_18262,N_16361,N_16732);
or U18263 (N_18263,N_17253,N_17082);
or U18264 (N_18264,N_16846,N_17080);
xnor U18265 (N_18265,N_16663,N_16581);
xor U18266 (N_18266,N_17091,N_16369);
nand U18267 (N_18267,N_16988,N_16461);
nor U18268 (N_18268,N_16344,N_17257);
or U18269 (N_18269,N_16544,N_16877);
and U18270 (N_18270,N_17027,N_17285);
nand U18271 (N_18271,N_16879,N_16414);
nor U18272 (N_18272,N_16478,N_16501);
and U18273 (N_18273,N_16587,N_17226);
xor U18274 (N_18274,N_16809,N_16851);
xor U18275 (N_18275,N_16330,N_16951);
xor U18276 (N_18276,N_17247,N_16442);
and U18277 (N_18277,N_16549,N_16825);
xor U18278 (N_18278,N_17181,N_16848);
nor U18279 (N_18279,N_17222,N_16902);
nand U18280 (N_18280,N_17279,N_16913);
and U18281 (N_18281,N_16460,N_16757);
and U18282 (N_18282,N_16657,N_17288);
nor U18283 (N_18283,N_17242,N_16562);
or U18284 (N_18284,N_16354,N_17093);
and U18285 (N_18285,N_16499,N_17113);
and U18286 (N_18286,N_16298,N_16908);
nand U18287 (N_18287,N_17029,N_17118);
xor U18288 (N_18288,N_16341,N_16967);
nand U18289 (N_18289,N_16323,N_16920);
or U18290 (N_18290,N_16825,N_16384);
nor U18291 (N_18291,N_16419,N_16589);
and U18292 (N_18292,N_16914,N_16299);
and U18293 (N_18293,N_17265,N_17215);
or U18294 (N_18294,N_16480,N_16486);
xor U18295 (N_18295,N_16956,N_17291);
nand U18296 (N_18296,N_16466,N_16839);
xor U18297 (N_18297,N_17471,N_17402);
and U18298 (N_18298,N_16758,N_16709);
nor U18299 (N_18299,N_16679,N_17364);
or U18300 (N_18300,N_16986,N_16898);
or U18301 (N_18301,N_16272,N_16871);
and U18302 (N_18302,N_17246,N_17264);
nor U18303 (N_18303,N_17368,N_16952);
nor U18304 (N_18304,N_16403,N_17199);
and U18305 (N_18305,N_17210,N_16257);
nand U18306 (N_18306,N_17320,N_17013);
xnor U18307 (N_18307,N_16539,N_16657);
xor U18308 (N_18308,N_16979,N_16902);
or U18309 (N_18309,N_16649,N_17189);
nor U18310 (N_18310,N_17004,N_17293);
nor U18311 (N_18311,N_16376,N_17147);
and U18312 (N_18312,N_16310,N_16361);
and U18313 (N_18313,N_17406,N_16611);
or U18314 (N_18314,N_17302,N_16913);
nand U18315 (N_18315,N_16506,N_16277);
and U18316 (N_18316,N_16426,N_16318);
nand U18317 (N_18317,N_17315,N_16324);
and U18318 (N_18318,N_17495,N_16493);
xor U18319 (N_18319,N_17027,N_17171);
nand U18320 (N_18320,N_17339,N_16802);
and U18321 (N_18321,N_17431,N_17280);
xor U18322 (N_18322,N_16469,N_17035);
nand U18323 (N_18323,N_16890,N_16595);
and U18324 (N_18324,N_16671,N_17343);
nor U18325 (N_18325,N_16932,N_16929);
nand U18326 (N_18326,N_17075,N_17113);
or U18327 (N_18327,N_17156,N_17059);
xnor U18328 (N_18328,N_17045,N_16698);
nand U18329 (N_18329,N_17480,N_16990);
and U18330 (N_18330,N_16327,N_17113);
and U18331 (N_18331,N_17484,N_16493);
nand U18332 (N_18332,N_16601,N_16453);
and U18333 (N_18333,N_16640,N_16671);
xnor U18334 (N_18334,N_17429,N_16615);
nand U18335 (N_18335,N_16339,N_17371);
and U18336 (N_18336,N_16569,N_16835);
and U18337 (N_18337,N_16462,N_16353);
nand U18338 (N_18338,N_17010,N_17043);
xor U18339 (N_18339,N_16496,N_16549);
nor U18340 (N_18340,N_16406,N_16933);
nand U18341 (N_18341,N_17142,N_16324);
xnor U18342 (N_18342,N_17146,N_16748);
nor U18343 (N_18343,N_16329,N_17226);
or U18344 (N_18344,N_17479,N_16424);
nor U18345 (N_18345,N_16466,N_16450);
xor U18346 (N_18346,N_16372,N_16252);
or U18347 (N_18347,N_17309,N_16287);
nand U18348 (N_18348,N_16830,N_16497);
or U18349 (N_18349,N_16918,N_16356);
or U18350 (N_18350,N_16767,N_16753);
and U18351 (N_18351,N_17237,N_17060);
nand U18352 (N_18352,N_16319,N_16484);
or U18353 (N_18353,N_17048,N_16279);
nand U18354 (N_18354,N_17441,N_16675);
or U18355 (N_18355,N_16669,N_16475);
xnor U18356 (N_18356,N_17278,N_17362);
xor U18357 (N_18357,N_16922,N_17419);
xor U18358 (N_18358,N_16325,N_17119);
and U18359 (N_18359,N_17476,N_16296);
and U18360 (N_18360,N_17337,N_17029);
and U18361 (N_18361,N_17259,N_17366);
and U18362 (N_18362,N_16368,N_16906);
or U18363 (N_18363,N_16719,N_17079);
nor U18364 (N_18364,N_16332,N_16437);
nand U18365 (N_18365,N_17384,N_17073);
and U18366 (N_18366,N_16923,N_16778);
and U18367 (N_18367,N_16355,N_17397);
xor U18368 (N_18368,N_16832,N_17226);
nand U18369 (N_18369,N_16547,N_16954);
and U18370 (N_18370,N_16546,N_17265);
xnor U18371 (N_18371,N_17035,N_17318);
xnor U18372 (N_18372,N_16392,N_17099);
nor U18373 (N_18373,N_17033,N_17094);
or U18374 (N_18374,N_16778,N_16678);
and U18375 (N_18375,N_16689,N_17477);
nand U18376 (N_18376,N_17409,N_16676);
and U18377 (N_18377,N_16657,N_17370);
nand U18378 (N_18378,N_17114,N_17374);
and U18379 (N_18379,N_16643,N_17086);
or U18380 (N_18380,N_17376,N_16322);
and U18381 (N_18381,N_16946,N_16662);
and U18382 (N_18382,N_17163,N_17194);
and U18383 (N_18383,N_16835,N_16610);
nor U18384 (N_18384,N_16268,N_16775);
and U18385 (N_18385,N_17037,N_17332);
or U18386 (N_18386,N_16674,N_17461);
and U18387 (N_18387,N_17373,N_16427);
nand U18388 (N_18388,N_17403,N_16909);
xor U18389 (N_18389,N_17481,N_16956);
nor U18390 (N_18390,N_16890,N_16387);
and U18391 (N_18391,N_16252,N_17046);
xor U18392 (N_18392,N_17184,N_16296);
xor U18393 (N_18393,N_16590,N_17284);
xnor U18394 (N_18394,N_17272,N_16390);
xnor U18395 (N_18395,N_16487,N_17471);
xor U18396 (N_18396,N_16643,N_17323);
or U18397 (N_18397,N_17406,N_16677);
and U18398 (N_18398,N_17378,N_17028);
nand U18399 (N_18399,N_17166,N_17207);
or U18400 (N_18400,N_17202,N_16753);
nor U18401 (N_18401,N_16848,N_17484);
or U18402 (N_18402,N_17354,N_16851);
or U18403 (N_18403,N_17251,N_16724);
or U18404 (N_18404,N_16463,N_16345);
nand U18405 (N_18405,N_17280,N_16546);
nor U18406 (N_18406,N_16304,N_16302);
and U18407 (N_18407,N_17049,N_16583);
nor U18408 (N_18408,N_16704,N_17211);
nor U18409 (N_18409,N_16836,N_16411);
and U18410 (N_18410,N_16582,N_16722);
nor U18411 (N_18411,N_16369,N_16625);
nor U18412 (N_18412,N_16571,N_16271);
or U18413 (N_18413,N_17284,N_16557);
or U18414 (N_18414,N_16951,N_16455);
nand U18415 (N_18415,N_16894,N_17096);
and U18416 (N_18416,N_16731,N_17142);
and U18417 (N_18417,N_16622,N_16441);
and U18418 (N_18418,N_16283,N_16575);
or U18419 (N_18419,N_16492,N_16788);
nand U18420 (N_18420,N_16707,N_17298);
xor U18421 (N_18421,N_16670,N_16547);
and U18422 (N_18422,N_16935,N_16622);
nand U18423 (N_18423,N_16950,N_16476);
or U18424 (N_18424,N_17424,N_17013);
nand U18425 (N_18425,N_16719,N_16813);
and U18426 (N_18426,N_16941,N_16485);
xnor U18427 (N_18427,N_17309,N_16767);
or U18428 (N_18428,N_16983,N_16404);
or U18429 (N_18429,N_17341,N_17489);
nand U18430 (N_18430,N_16916,N_16917);
or U18431 (N_18431,N_16297,N_17307);
and U18432 (N_18432,N_16886,N_17409);
or U18433 (N_18433,N_17261,N_16390);
and U18434 (N_18434,N_16723,N_16395);
nor U18435 (N_18435,N_16335,N_17457);
nor U18436 (N_18436,N_17446,N_17380);
xnor U18437 (N_18437,N_17476,N_17007);
xnor U18438 (N_18438,N_16862,N_16449);
and U18439 (N_18439,N_16722,N_17479);
nand U18440 (N_18440,N_17244,N_16689);
xnor U18441 (N_18441,N_17025,N_16406);
nor U18442 (N_18442,N_16911,N_16871);
nor U18443 (N_18443,N_17084,N_17356);
nor U18444 (N_18444,N_16776,N_16922);
xor U18445 (N_18445,N_16783,N_17204);
nand U18446 (N_18446,N_16524,N_16471);
nand U18447 (N_18447,N_17094,N_16599);
nor U18448 (N_18448,N_17406,N_16446);
and U18449 (N_18449,N_17077,N_16508);
nor U18450 (N_18450,N_17051,N_17394);
and U18451 (N_18451,N_16374,N_17264);
nand U18452 (N_18452,N_16457,N_16393);
xnor U18453 (N_18453,N_16551,N_16887);
nor U18454 (N_18454,N_16276,N_16289);
xor U18455 (N_18455,N_16840,N_16612);
and U18456 (N_18456,N_16606,N_17247);
xor U18457 (N_18457,N_16434,N_17464);
nand U18458 (N_18458,N_16657,N_16771);
and U18459 (N_18459,N_16612,N_16352);
nor U18460 (N_18460,N_17288,N_17423);
nand U18461 (N_18461,N_16850,N_16667);
nand U18462 (N_18462,N_17102,N_17146);
and U18463 (N_18463,N_16753,N_17482);
nor U18464 (N_18464,N_17079,N_16930);
nand U18465 (N_18465,N_17017,N_16969);
and U18466 (N_18466,N_17321,N_16563);
nor U18467 (N_18467,N_17057,N_16986);
or U18468 (N_18468,N_17079,N_16402);
or U18469 (N_18469,N_16936,N_16787);
and U18470 (N_18470,N_17493,N_16504);
nand U18471 (N_18471,N_16859,N_16403);
xor U18472 (N_18472,N_17291,N_17256);
and U18473 (N_18473,N_17238,N_16365);
nor U18474 (N_18474,N_16371,N_17438);
xor U18475 (N_18475,N_17267,N_17164);
and U18476 (N_18476,N_16696,N_16909);
nand U18477 (N_18477,N_16374,N_17395);
nor U18478 (N_18478,N_16404,N_16913);
and U18479 (N_18479,N_16476,N_16363);
or U18480 (N_18480,N_17163,N_17228);
xor U18481 (N_18481,N_16492,N_16649);
nand U18482 (N_18482,N_17101,N_17195);
or U18483 (N_18483,N_16293,N_16353);
xnor U18484 (N_18484,N_16565,N_16406);
and U18485 (N_18485,N_17328,N_16538);
or U18486 (N_18486,N_16984,N_16412);
and U18487 (N_18487,N_16684,N_17417);
or U18488 (N_18488,N_16278,N_16470);
and U18489 (N_18489,N_16714,N_17263);
or U18490 (N_18490,N_17069,N_16653);
nand U18491 (N_18491,N_16854,N_17420);
nand U18492 (N_18492,N_16973,N_16708);
xor U18493 (N_18493,N_16480,N_17133);
nor U18494 (N_18494,N_16498,N_17483);
and U18495 (N_18495,N_16767,N_16875);
and U18496 (N_18496,N_16662,N_16338);
nor U18497 (N_18497,N_16920,N_17255);
or U18498 (N_18498,N_16359,N_16633);
nand U18499 (N_18499,N_16977,N_17045);
nor U18500 (N_18500,N_17177,N_16590);
or U18501 (N_18501,N_16384,N_17402);
or U18502 (N_18502,N_17279,N_16781);
nand U18503 (N_18503,N_17256,N_17466);
and U18504 (N_18504,N_16611,N_16956);
xor U18505 (N_18505,N_17072,N_16292);
nand U18506 (N_18506,N_16948,N_16270);
nor U18507 (N_18507,N_16258,N_17337);
nand U18508 (N_18508,N_16872,N_16426);
xor U18509 (N_18509,N_16383,N_16502);
and U18510 (N_18510,N_16462,N_16937);
xnor U18511 (N_18511,N_16574,N_16984);
xnor U18512 (N_18512,N_16740,N_16586);
nor U18513 (N_18513,N_17482,N_17005);
or U18514 (N_18514,N_16472,N_17354);
xnor U18515 (N_18515,N_16518,N_17392);
nor U18516 (N_18516,N_16678,N_17067);
nor U18517 (N_18517,N_16944,N_17260);
and U18518 (N_18518,N_16886,N_16694);
xnor U18519 (N_18519,N_17042,N_17390);
nand U18520 (N_18520,N_16726,N_16282);
nand U18521 (N_18521,N_17477,N_16678);
and U18522 (N_18522,N_17321,N_16936);
nand U18523 (N_18523,N_16774,N_16508);
nand U18524 (N_18524,N_17387,N_17439);
and U18525 (N_18525,N_17138,N_16796);
nor U18526 (N_18526,N_16367,N_17412);
nand U18527 (N_18527,N_16964,N_16490);
and U18528 (N_18528,N_16902,N_16597);
nor U18529 (N_18529,N_16620,N_17458);
xor U18530 (N_18530,N_16953,N_17030);
or U18531 (N_18531,N_16930,N_16860);
and U18532 (N_18532,N_17375,N_16422);
and U18533 (N_18533,N_17126,N_17202);
nand U18534 (N_18534,N_16773,N_16446);
and U18535 (N_18535,N_16266,N_17290);
nor U18536 (N_18536,N_17050,N_17183);
nand U18537 (N_18537,N_16916,N_16754);
xor U18538 (N_18538,N_17316,N_16933);
nor U18539 (N_18539,N_17318,N_16804);
xnor U18540 (N_18540,N_16491,N_16614);
or U18541 (N_18541,N_16351,N_16832);
nand U18542 (N_18542,N_16562,N_16881);
xnor U18543 (N_18543,N_16364,N_16696);
nor U18544 (N_18544,N_17257,N_16659);
or U18545 (N_18545,N_17330,N_17026);
or U18546 (N_18546,N_17407,N_16622);
nand U18547 (N_18547,N_16661,N_16327);
and U18548 (N_18548,N_16859,N_17247);
and U18549 (N_18549,N_17309,N_16316);
nand U18550 (N_18550,N_16314,N_16796);
nand U18551 (N_18551,N_17195,N_16419);
or U18552 (N_18552,N_16973,N_16530);
nor U18553 (N_18553,N_17333,N_16856);
nor U18554 (N_18554,N_16289,N_16954);
nor U18555 (N_18555,N_17090,N_16279);
and U18556 (N_18556,N_16858,N_16690);
and U18557 (N_18557,N_16715,N_16406);
nand U18558 (N_18558,N_17465,N_16789);
and U18559 (N_18559,N_17270,N_16265);
and U18560 (N_18560,N_16503,N_17208);
nand U18561 (N_18561,N_16396,N_16852);
nor U18562 (N_18562,N_16790,N_16940);
nand U18563 (N_18563,N_16321,N_17348);
xor U18564 (N_18564,N_17438,N_16678);
nand U18565 (N_18565,N_16575,N_16728);
xnor U18566 (N_18566,N_16489,N_16548);
xnor U18567 (N_18567,N_16257,N_16682);
nor U18568 (N_18568,N_16447,N_17343);
or U18569 (N_18569,N_16501,N_17093);
nand U18570 (N_18570,N_17445,N_16920);
xnor U18571 (N_18571,N_16250,N_17056);
and U18572 (N_18572,N_16478,N_17054);
xor U18573 (N_18573,N_17407,N_17172);
nor U18574 (N_18574,N_16838,N_16936);
and U18575 (N_18575,N_17399,N_16301);
or U18576 (N_18576,N_16753,N_16651);
nor U18577 (N_18577,N_16551,N_17135);
or U18578 (N_18578,N_16360,N_16895);
or U18579 (N_18579,N_17369,N_16606);
xnor U18580 (N_18580,N_16618,N_17475);
or U18581 (N_18581,N_16716,N_16539);
xor U18582 (N_18582,N_17343,N_17001);
and U18583 (N_18583,N_17035,N_16575);
nor U18584 (N_18584,N_17473,N_16998);
xor U18585 (N_18585,N_16902,N_16293);
xor U18586 (N_18586,N_17069,N_16609);
nor U18587 (N_18587,N_17233,N_17457);
nand U18588 (N_18588,N_17297,N_17400);
nand U18589 (N_18589,N_17484,N_16789);
nand U18590 (N_18590,N_16910,N_16789);
and U18591 (N_18591,N_16250,N_16259);
or U18592 (N_18592,N_16297,N_16328);
xor U18593 (N_18593,N_16856,N_16393);
and U18594 (N_18594,N_17222,N_17318);
xnor U18595 (N_18595,N_16454,N_16475);
xor U18596 (N_18596,N_16689,N_17223);
nand U18597 (N_18597,N_16676,N_16899);
and U18598 (N_18598,N_17090,N_16767);
nor U18599 (N_18599,N_16736,N_16794);
xor U18600 (N_18600,N_16703,N_17036);
xor U18601 (N_18601,N_16447,N_16603);
nand U18602 (N_18602,N_17242,N_16626);
nor U18603 (N_18603,N_16662,N_17059);
nand U18604 (N_18604,N_17386,N_17382);
or U18605 (N_18605,N_16371,N_16984);
and U18606 (N_18606,N_16480,N_16736);
and U18607 (N_18607,N_16790,N_16431);
nand U18608 (N_18608,N_16396,N_17025);
and U18609 (N_18609,N_17414,N_17498);
xor U18610 (N_18610,N_17063,N_17040);
xnor U18611 (N_18611,N_16759,N_16953);
or U18612 (N_18612,N_17066,N_16987);
or U18613 (N_18613,N_16719,N_17399);
or U18614 (N_18614,N_16413,N_16788);
or U18615 (N_18615,N_16769,N_16837);
nand U18616 (N_18616,N_16332,N_17105);
nor U18617 (N_18617,N_16638,N_16643);
nor U18618 (N_18618,N_17343,N_16336);
nor U18619 (N_18619,N_17380,N_16586);
nand U18620 (N_18620,N_16688,N_17412);
xor U18621 (N_18621,N_17002,N_16965);
or U18622 (N_18622,N_16372,N_16352);
and U18623 (N_18623,N_16623,N_16790);
xnor U18624 (N_18624,N_17357,N_17347);
nor U18625 (N_18625,N_16307,N_17243);
xor U18626 (N_18626,N_16382,N_16473);
nand U18627 (N_18627,N_16808,N_17155);
or U18628 (N_18628,N_17397,N_16795);
and U18629 (N_18629,N_17311,N_16589);
nand U18630 (N_18630,N_16622,N_17058);
and U18631 (N_18631,N_16289,N_16676);
nand U18632 (N_18632,N_16632,N_17307);
and U18633 (N_18633,N_17365,N_16947);
or U18634 (N_18634,N_17011,N_16890);
or U18635 (N_18635,N_17091,N_16414);
xor U18636 (N_18636,N_16940,N_16727);
nand U18637 (N_18637,N_17455,N_16660);
nor U18638 (N_18638,N_16623,N_16548);
nand U18639 (N_18639,N_17326,N_17472);
or U18640 (N_18640,N_16346,N_17261);
nand U18641 (N_18641,N_17281,N_16277);
xor U18642 (N_18642,N_17382,N_16727);
or U18643 (N_18643,N_16838,N_17246);
xnor U18644 (N_18644,N_16517,N_17102);
nor U18645 (N_18645,N_17295,N_16627);
or U18646 (N_18646,N_17368,N_16393);
xor U18647 (N_18647,N_16371,N_16763);
nor U18648 (N_18648,N_16906,N_16470);
or U18649 (N_18649,N_17293,N_16726);
nand U18650 (N_18650,N_17217,N_16726);
nor U18651 (N_18651,N_16793,N_16456);
nor U18652 (N_18652,N_17255,N_17288);
and U18653 (N_18653,N_17316,N_17019);
nor U18654 (N_18654,N_16716,N_16560);
or U18655 (N_18655,N_16760,N_16642);
xnor U18656 (N_18656,N_16808,N_16817);
nor U18657 (N_18657,N_16378,N_17109);
nor U18658 (N_18658,N_16739,N_16575);
xnor U18659 (N_18659,N_17060,N_16617);
nand U18660 (N_18660,N_16326,N_16928);
xor U18661 (N_18661,N_16826,N_16444);
or U18662 (N_18662,N_16278,N_16563);
nor U18663 (N_18663,N_16919,N_17096);
xnor U18664 (N_18664,N_16938,N_17153);
xnor U18665 (N_18665,N_16524,N_16344);
or U18666 (N_18666,N_16898,N_16630);
and U18667 (N_18667,N_17065,N_16683);
xnor U18668 (N_18668,N_16281,N_17023);
xnor U18669 (N_18669,N_16710,N_17368);
nor U18670 (N_18670,N_16551,N_16684);
xor U18671 (N_18671,N_16969,N_16848);
nand U18672 (N_18672,N_16542,N_16528);
nor U18673 (N_18673,N_16940,N_16651);
nor U18674 (N_18674,N_16404,N_16621);
nand U18675 (N_18675,N_17064,N_16705);
nand U18676 (N_18676,N_17456,N_16777);
or U18677 (N_18677,N_17421,N_17021);
xnor U18678 (N_18678,N_16843,N_16955);
xnor U18679 (N_18679,N_17124,N_16519);
and U18680 (N_18680,N_16910,N_17167);
nor U18681 (N_18681,N_16927,N_17213);
xnor U18682 (N_18682,N_16250,N_16916);
and U18683 (N_18683,N_16340,N_17243);
and U18684 (N_18684,N_16597,N_16620);
nand U18685 (N_18685,N_16529,N_17039);
or U18686 (N_18686,N_17443,N_16758);
or U18687 (N_18687,N_16487,N_16261);
nand U18688 (N_18688,N_17467,N_16823);
and U18689 (N_18689,N_16291,N_16407);
xnor U18690 (N_18690,N_17482,N_17490);
and U18691 (N_18691,N_17265,N_17176);
nor U18692 (N_18692,N_17113,N_17190);
or U18693 (N_18693,N_17010,N_16996);
nand U18694 (N_18694,N_17414,N_16506);
nor U18695 (N_18695,N_17205,N_16670);
or U18696 (N_18696,N_16809,N_17083);
nor U18697 (N_18697,N_17468,N_16459);
xnor U18698 (N_18698,N_16594,N_16551);
and U18699 (N_18699,N_16907,N_16913);
nor U18700 (N_18700,N_17342,N_16588);
xor U18701 (N_18701,N_16883,N_16857);
xnor U18702 (N_18702,N_16620,N_17012);
nand U18703 (N_18703,N_16261,N_16633);
and U18704 (N_18704,N_16514,N_17188);
nand U18705 (N_18705,N_16609,N_17317);
or U18706 (N_18706,N_16821,N_16919);
and U18707 (N_18707,N_16322,N_16522);
or U18708 (N_18708,N_16296,N_16755);
nor U18709 (N_18709,N_16984,N_17416);
or U18710 (N_18710,N_16358,N_16279);
and U18711 (N_18711,N_16546,N_16757);
nand U18712 (N_18712,N_17057,N_17338);
and U18713 (N_18713,N_16527,N_16581);
nand U18714 (N_18714,N_16966,N_17117);
and U18715 (N_18715,N_17488,N_16671);
nor U18716 (N_18716,N_16889,N_16759);
nor U18717 (N_18717,N_16664,N_16409);
and U18718 (N_18718,N_17185,N_16503);
and U18719 (N_18719,N_16662,N_16945);
xnor U18720 (N_18720,N_17497,N_16304);
and U18721 (N_18721,N_16317,N_17044);
or U18722 (N_18722,N_16981,N_17389);
xor U18723 (N_18723,N_17396,N_17484);
and U18724 (N_18724,N_17262,N_17030);
or U18725 (N_18725,N_16504,N_17397);
nor U18726 (N_18726,N_17143,N_17218);
xnor U18727 (N_18727,N_17266,N_16607);
nor U18728 (N_18728,N_17244,N_17454);
nor U18729 (N_18729,N_16966,N_17400);
or U18730 (N_18730,N_16571,N_16646);
xor U18731 (N_18731,N_16506,N_17074);
or U18732 (N_18732,N_16615,N_16326);
xor U18733 (N_18733,N_17218,N_16744);
nor U18734 (N_18734,N_17425,N_16910);
or U18735 (N_18735,N_16657,N_17357);
or U18736 (N_18736,N_17392,N_16702);
nor U18737 (N_18737,N_16441,N_16415);
nand U18738 (N_18738,N_16641,N_16286);
xnor U18739 (N_18739,N_16965,N_16306);
nor U18740 (N_18740,N_17381,N_16355);
nor U18741 (N_18741,N_17281,N_16584);
or U18742 (N_18742,N_16603,N_16387);
or U18743 (N_18743,N_17440,N_16524);
and U18744 (N_18744,N_16945,N_16475);
or U18745 (N_18745,N_16858,N_16555);
or U18746 (N_18746,N_17409,N_16816);
nor U18747 (N_18747,N_17438,N_16814);
xor U18748 (N_18748,N_16717,N_17300);
nor U18749 (N_18749,N_16993,N_17178);
nor U18750 (N_18750,N_17644,N_17765);
nand U18751 (N_18751,N_17934,N_18369);
or U18752 (N_18752,N_18548,N_18327);
nand U18753 (N_18753,N_18378,N_18269);
or U18754 (N_18754,N_18550,N_17935);
or U18755 (N_18755,N_17691,N_17685);
nand U18756 (N_18756,N_17673,N_18163);
nor U18757 (N_18757,N_18415,N_17723);
nand U18758 (N_18758,N_17928,N_18153);
nor U18759 (N_18759,N_18296,N_17834);
xor U18760 (N_18760,N_18497,N_17949);
nand U18761 (N_18761,N_17604,N_18399);
nand U18762 (N_18762,N_17745,N_18741);
nor U18763 (N_18763,N_17826,N_17915);
xor U18764 (N_18764,N_18610,N_17579);
xor U18765 (N_18765,N_17594,N_18037);
or U18766 (N_18766,N_17965,N_17818);
xor U18767 (N_18767,N_18594,N_18410);
and U18768 (N_18768,N_17791,N_18141);
and U18769 (N_18769,N_18329,N_18182);
and U18770 (N_18770,N_17546,N_18565);
xnor U18771 (N_18771,N_18374,N_18189);
nand U18772 (N_18772,N_18590,N_18098);
nand U18773 (N_18773,N_18036,N_18744);
nor U18774 (N_18774,N_18718,N_18161);
xnor U18775 (N_18775,N_18241,N_18411);
xor U18776 (N_18776,N_17982,N_18691);
and U18777 (N_18777,N_17681,N_18686);
nand U18778 (N_18778,N_18668,N_18462);
and U18779 (N_18779,N_18186,N_18035);
or U18780 (N_18780,N_17764,N_18057);
or U18781 (N_18781,N_18704,N_17952);
nand U18782 (N_18782,N_18480,N_17812);
xnor U18783 (N_18783,N_18513,N_18087);
nand U18784 (N_18784,N_18324,N_17777);
nand U18785 (N_18785,N_17648,N_18725);
xor U18786 (N_18786,N_17809,N_18575);
nand U18787 (N_18787,N_18446,N_18094);
xnor U18788 (N_18788,N_18661,N_17666);
and U18789 (N_18789,N_18109,N_18184);
or U18790 (N_18790,N_18009,N_17823);
or U18791 (N_18791,N_18309,N_17600);
xor U18792 (N_18792,N_18564,N_17801);
xnor U18793 (N_18793,N_17899,N_18418);
nor U18794 (N_18794,N_18165,N_17758);
or U18795 (N_18795,N_18567,N_18681);
and U18796 (N_18796,N_18099,N_17802);
nor U18797 (N_18797,N_17531,N_18749);
and U18798 (N_18798,N_17654,N_18102);
or U18799 (N_18799,N_17612,N_18217);
or U18800 (N_18800,N_17845,N_17969);
xor U18801 (N_18801,N_17553,N_17533);
nor U18802 (N_18802,N_18291,N_18322);
nor U18803 (N_18803,N_18563,N_17943);
and U18804 (N_18804,N_17995,N_18007);
and U18805 (N_18805,N_17857,N_17595);
nor U18806 (N_18806,N_17505,N_18675);
and U18807 (N_18807,N_18438,N_18655);
xor U18808 (N_18808,N_17716,N_18043);
nand U18809 (N_18809,N_18233,N_18597);
xor U18810 (N_18810,N_17848,N_17903);
nor U18811 (N_18811,N_18601,N_18008);
or U18812 (N_18812,N_18228,N_17994);
or U18813 (N_18813,N_18142,N_18650);
nand U18814 (N_18814,N_18721,N_18637);
nand U18815 (N_18815,N_18658,N_17709);
nor U18816 (N_18816,N_18237,N_17862);
nand U18817 (N_18817,N_18295,N_18254);
or U18818 (N_18818,N_18458,N_17762);
nand U18819 (N_18819,N_18204,N_18040);
or U18820 (N_18820,N_18588,N_18058);
nor U18821 (N_18821,N_18128,N_17635);
nand U18822 (N_18822,N_17798,N_18012);
nor U18823 (N_18823,N_18112,N_17643);
nor U18824 (N_18824,N_17755,N_17910);
or U18825 (N_18825,N_17953,N_17835);
xnor U18826 (N_18826,N_18486,N_17732);
nor U18827 (N_18827,N_18049,N_18320);
and U18828 (N_18828,N_18314,N_17997);
nand U18829 (N_18829,N_18738,N_18346);
and U18830 (N_18830,N_18245,N_18337);
and U18831 (N_18831,N_18286,N_18046);
or U18832 (N_18832,N_18589,N_18420);
and U18833 (N_18833,N_17895,N_17627);
nand U18834 (N_18834,N_18617,N_17854);
and U18835 (N_18835,N_18274,N_18465);
xnor U18836 (N_18836,N_18082,N_17678);
nor U18837 (N_18837,N_17660,N_18727);
nand U18838 (N_18838,N_17573,N_18443);
xnor U18839 (N_18839,N_18440,N_17789);
nor U18840 (N_18840,N_17571,N_18249);
or U18841 (N_18841,N_17617,N_18527);
nor U18842 (N_18842,N_18229,N_18384);
and U18843 (N_18843,N_18074,N_17879);
nor U18844 (N_18844,N_17704,N_18195);
or U18845 (N_18845,N_18679,N_18626);
and U18846 (N_18846,N_17568,N_17547);
and U18847 (N_18847,N_17615,N_18522);
nand U18848 (N_18848,N_17872,N_18580);
and U18849 (N_18849,N_18545,N_18717);
xor U18850 (N_18850,N_18654,N_18516);
nor U18851 (N_18851,N_17596,N_17698);
nand U18852 (N_18852,N_17833,N_17729);
xor U18853 (N_18853,N_17944,N_18022);
nor U18854 (N_18854,N_18616,N_17774);
nor U18855 (N_18855,N_17780,N_18431);
nor U18856 (N_18856,N_18192,N_17775);
and U18857 (N_18857,N_18119,N_17610);
nor U18858 (N_18858,N_17913,N_17770);
and U18859 (N_18859,N_18200,N_17530);
and U18860 (N_18860,N_18129,N_18305);
or U18861 (N_18861,N_17737,N_18501);
and U18862 (N_18862,N_18653,N_17511);
nand U18863 (N_18863,N_18735,N_17683);
and U18864 (N_18864,N_17890,N_18151);
nand U18865 (N_18865,N_18212,N_17750);
or U18866 (N_18866,N_18439,N_18147);
xor U18867 (N_18867,N_17649,N_18317);
and U18868 (N_18868,N_18338,N_18648);
and U18869 (N_18869,N_17911,N_17696);
xnor U18870 (N_18870,N_18521,N_18412);
nor U18871 (N_18871,N_18600,N_18507);
nand U18872 (N_18872,N_18070,N_18408);
or U18873 (N_18873,N_17695,N_18061);
or U18874 (N_18874,N_18619,N_17708);
nand U18875 (N_18875,N_18013,N_17877);
xnor U18876 (N_18876,N_18724,N_18442);
nor U18877 (N_18877,N_17688,N_18244);
xor U18878 (N_18878,N_18183,N_17807);
or U18879 (N_18879,N_17527,N_17856);
nand U18880 (N_18880,N_18341,N_17622);
nor U18881 (N_18881,N_18086,N_17677);
nand U18882 (N_18882,N_18194,N_17738);
nand U18883 (N_18883,N_17880,N_18703);
xnor U18884 (N_18884,N_17513,N_18559);
or U18885 (N_18885,N_18288,N_18586);
and U18886 (N_18886,N_18067,N_18253);
or U18887 (N_18887,N_17817,N_18282);
or U18888 (N_18888,N_18148,N_17693);
nor U18889 (N_18889,N_17984,N_18172);
or U18890 (N_18890,N_17979,N_18323);
xnor U18891 (N_18891,N_17878,N_18390);
xor U18892 (N_18892,N_18268,N_17523);
nand U18893 (N_18893,N_18598,N_18330);
and U18894 (N_18894,N_17931,N_18199);
xnor U18895 (N_18895,N_17597,N_18391);
nor U18896 (N_18896,N_17728,N_17510);
and U18897 (N_18897,N_18020,N_17633);
or U18898 (N_18898,N_18325,N_17968);
and U18899 (N_18899,N_17605,N_18731);
nor U18900 (N_18900,N_17850,N_18169);
nor U18901 (N_18901,N_18145,N_17672);
xnor U18902 (N_18902,N_18072,N_18419);
nand U18903 (N_18903,N_17796,N_18352);
and U18904 (N_18904,N_18572,N_17577);
xnor U18905 (N_18905,N_18478,N_18092);
or U18906 (N_18906,N_18059,N_18311);
and U18907 (N_18907,N_18555,N_17908);
nor U18908 (N_18908,N_18488,N_17947);
xor U18909 (N_18909,N_18298,N_18685);
nor U18910 (N_18910,N_17822,N_17957);
nand U18911 (N_18911,N_17570,N_17967);
xnor U18912 (N_18912,N_18080,N_17682);
nand U18913 (N_18913,N_18001,N_18400);
or U18914 (N_18914,N_18381,N_17790);
xnor U18915 (N_18915,N_18706,N_18726);
xor U18916 (N_18916,N_18417,N_18505);
xnor U18917 (N_18917,N_18160,N_18236);
and U18918 (N_18918,N_18582,N_18697);
nand U18919 (N_18919,N_18719,N_18243);
or U18920 (N_18920,N_18068,N_18468);
nor U18921 (N_18921,N_18225,N_17532);
xor U18922 (N_18922,N_18720,N_17506);
and U18923 (N_18923,N_18302,N_17501);
or U18924 (N_18924,N_17656,N_18124);
or U18925 (N_18925,N_18174,N_18081);
xnor U18926 (N_18926,N_17588,N_18461);
nand U18927 (N_18927,N_17827,N_17962);
and U18928 (N_18928,N_17689,N_18078);
nor U18929 (N_18929,N_18613,N_18167);
nor U18930 (N_18930,N_18076,N_18742);
or U18931 (N_18931,N_18517,N_17528);
xnor U18932 (N_18932,N_18052,N_18694);
xnor U18933 (N_18933,N_17863,N_17629);
or U18934 (N_18934,N_17799,N_18427);
nor U18935 (N_18935,N_18005,N_18349);
or U18936 (N_18936,N_18010,N_18606);
xor U18937 (N_18937,N_18248,N_17983);
or U18938 (N_18938,N_17989,N_18596);
or U18939 (N_18939,N_17876,N_17832);
and U18940 (N_18940,N_17902,N_18357);
nand U18941 (N_18941,N_17509,N_17507);
and U18942 (N_18942,N_18413,N_18259);
nor U18943 (N_18943,N_18403,N_17756);
nand U18944 (N_18944,N_17580,N_18041);
nand U18945 (N_18945,N_17724,N_18529);
xor U18946 (N_18946,N_18592,N_18624);
nor U18947 (N_18947,N_17893,N_17946);
nand U18948 (N_18948,N_18437,N_17592);
nand U18949 (N_18949,N_18304,N_17978);
xnor U18950 (N_18950,N_18159,N_18347);
nor U18951 (N_18951,N_17831,N_18371);
nor U18952 (N_18952,N_18034,N_18045);
xnor U18953 (N_18953,N_18083,N_18331);
or U18954 (N_18954,N_17922,N_18515);
nand U18955 (N_18955,N_18230,N_17529);
xor U18956 (N_18956,N_17519,N_18105);
or U18957 (N_18957,N_17961,N_17917);
nand U18958 (N_18958,N_18278,N_18472);
xnor U18959 (N_18959,N_18353,N_17587);
nor U18960 (N_18960,N_17853,N_17987);
nor U18961 (N_18961,N_17992,N_18451);
xnor U18962 (N_18962,N_18239,N_17690);
nor U18963 (N_18963,N_17508,N_18541);
and U18964 (N_18964,N_18232,N_17930);
nand U18965 (N_18965,N_18047,N_18688);
xor U18966 (N_18966,N_17646,N_17981);
nor U18967 (N_18967,N_18342,N_17674);
nand U18968 (N_18968,N_18700,N_18503);
nand U18969 (N_18969,N_18250,N_18348);
xnor U18970 (N_18970,N_17858,N_18262);
nand U18971 (N_18971,N_17891,N_18463);
or U18972 (N_18972,N_18170,N_18379);
nor U18973 (N_18973,N_17933,N_18428);
and U18974 (N_18974,N_18133,N_17904);
nand U18975 (N_18975,N_18635,N_17781);
or U18976 (N_18976,N_17515,N_18711);
xor U18977 (N_18977,N_17558,N_18456);
nor U18978 (N_18978,N_17616,N_18623);
nand U18979 (N_18979,N_18090,N_18602);
or U18980 (N_18980,N_17581,N_18270);
nand U18981 (N_18981,N_17972,N_17684);
nand U18982 (N_18982,N_17563,N_18445);
and U18983 (N_18983,N_17898,N_17793);
and U18984 (N_18984,N_17794,N_18748);
xnor U18985 (N_18985,N_18543,N_17769);
nor U18986 (N_18986,N_17540,N_18044);
or U18987 (N_18987,N_18407,N_18432);
and U18988 (N_18988,N_18321,N_18690);
xnor U18989 (N_18989,N_18401,N_17544);
and U18990 (N_18990,N_18475,N_18332);
and U18991 (N_18991,N_17759,N_18476);
nand U18992 (N_18992,N_18227,N_17667);
xnor U18993 (N_18993,N_17557,N_17866);
or U18994 (N_18994,N_18743,N_18271);
and U18995 (N_18995,N_18028,N_18131);
xor U18996 (N_18996,N_17868,N_18179);
or U18997 (N_18997,N_18389,N_17865);
and U18998 (N_18998,N_17749,N_18190);
nand U18999 (N_18999,N_17779,N_18123);
nand U19000 (N_19000,N_18143,N_17657);
xnor U19001 (N_19001,N_17645,N_18662);
nand U19002 (N_19002,N_17717,N_18669);
or U19003 (N_19003,N_18649,N_18627);
or U19004 (N_19004,N_18651,N_18642);
and U19005 (N_19005,N_17734,N_18027);
or U19006 (N_19006,N_18433,N_17813);
or U19007 (N_19007,N_17929,N_17719);
nor U19008 (N_19008,N_18361,N_17601);
or U19009 (N_19009,N_17885,N_17718);
and U19010 (N_19010,N_17614,N_17819);
nor U19011 (N_19011,N_18453,N_18292);
or U19012 (N_19012,N_17840,N_18496);
and U19013 (N_19013,N_18483,N_18523);
and U19014 (N_19014,N_17503,N_17516);
and U19015 (N_19015,N_18603,N_17680);
and U19016 (N_19016,N_18150,N_17650);
xor U19017 (N_19017,N_18025,N_17603);
or U19018 (N_19018,N_18493,N_18033);
xor U19019 (N_19019,N_18444,N_17748);
xor U19020 (N_19020,N_18712,N_18604);
nor U19021 (N_19021,N_18158,N_17782);
nor U19022 (N_19022,N_18376,N_18615);
nand U19023 (N_19023,N_17959,N_17873);
or U19024 (N_19024,N_18581,N_17720);
and U19025 (N_19025,N_18645,N_18577);
or U19026 (N_19026,N_18100,N_17535);
xnor U19027 (N_19027,N_18614,N_18152);
or U19028 (N_19028,N_17816,N_18089);
and U19029 (N_19029,N_18104,N_17804);
and U19030 (N_19030,N_18071,N_18457);
and U19031 (N_19031,N_17730,N_18514);
and U19032 (N_19032,N_18287,N_17653);
nor U19033 (N_19033,N_17549,N_18739);
nand U19034 (N_19034,N_17569,N_18121);
nand U19035 (N_19035,N_18538,N_17555);
or U19036 (N_19036,N_18238,N_18211);
nor U19037 (N_19037,N_17806,N_18696);
or U19038 (N_19038,N_17733,N_17619);
nand U19039 (N_19039,N_18519,N_17537);
nand U19040 (N_19040,N_18546,N_18388);
nand U19041 (N_19041,N_18032,N_17810);
nand U19042 (N_19042,N_18737,N_18224);
nand U19043 (N_19043,N_18272,N_18019);
nor U19044 (N_19044,N_18713,N_18672);
nor U19045 (N_19045,N_18307,N_18447);
xnor U19046 (N_19046,N_17640,N_18290);
or U19047 (N_19047,N_18063,N_17921);
xnor U19048 (N_19048,N_17602,N_17520);
or U19049 (N_19049,N_18740,N_18464);
or U19050 (N_19050,N_17955,N_18530);
or U19051 (N_19051,N_18017,N_18149);
nand U19052 (N_19052,N_17889,N_18671);
or U19053 (N_19053,N_18116,N_17638);
xor U19054 (N_19054,N_18065,N_17963);
nand U19055 (N_19055,N_17714,N_17901);
nor U19056 (N_19056,N_17954,N_17974);
xor U19057 (N_19057,N_18485,N_17783);
nand U19058 (N_19058,N_18518,N_18511);
xor U19059 (N_19059,N_17937,N_17578);
nor U19060 (N_19060,N_18042,N_17741);
or U19061 (N_19061,N_17788,N_18351);
or U19062 (N_19062,N_18197,N_18144);
or U19063 (N_19063,N_17652,N_17727);
nor U19064 (N_19064,N_18266,N_17642);
nor U19065 (N_19065,N_18684,N_18356);
or U19066 (N_19066,N_17631,N_18409);
nand U19067 (N_19067,N_17907,N_18069);
xnor U19068 (N_19068,N_18556,N_18535);
or U19069 (N_19069,N_18628,N_18364);
nand U19070 (N_19070,N_18695,N_18216);
nand U19071 (N_19071,N_18360,N_18449);
nor U19072 (N_19072,N_17940,N_17665);
and U19073 (N_19073,N_18492,N_18608);
nor U19074 (N_19074,N_18732,N_18736);
nor U19075 (N_19075,N_17998,N_18607);
nand U19076 (N_19076,N_17960,N_18632);
or U19077 (N_19077,N_18441,N_18095);
and U19078 (N_19078,N_17882,N_18355);
xor U19079 (N_19079,N_18051,N_17566);
xor U19080 (N_19080,N_17773,N_18162);
nor U19081 (N_19081,N_18377,N_18508);
or U19082 (N_19082,N_17636,N_17609);
or U19083 (N_19083,N_17512,N_18459);
and U19084 (N_19084,N_17875,N_18715);
or U19085 (N_19085,N_18297,N_17837);
or U19086 (N_19086,N_17990,N_18576);
and U19087 (N_19087,N_18281,N_18023);
nand U19088 (N_19088,N_18294,N_17739);
nand U19089 (N_19089,N_18710,N_17658);
nor U19090 (N_19090,N_18219,N_18692);
nand U19091 (N_19091,N_18643,N_17870);
nor U19092 (N_19092,N_18506,N_18641);
and U19093 (N_19093,N_18114,N_17800);
and U19094 (N_19094,N_18549,N_17589);
nand U19095 (N_19095,N_18479,N_17668);
and U19096 (N_19096,N_18584,N_18489);
xor U19097 (N_19097,N_17561,N_18373);
and U19098 (N_19098,N_18689,N_18639);
and U19099 (N_19099,N_17628,N_17771);
xor U19100 (N_19100,N_17585,N_17951);
nand U19101 (N_19101,N_18264,N_17766);
nor U19102 (N_19102,N_17575,N_18175);
or U19103 (N_19103,N_18263,N_18132);
xnor U19104 (N_19104,N_17752,N_18191);
xnor U19105 (N_19105,N_17829,N_18289);
and U19106 (N_19106,N_18004,N_18499);
or U19107 (N_19107,N_18510,N_17787);
nand U19108 (N_19108,N_18716,N_17836);
or U19109 (N_19109,N_18405,N_17841);
or U19110 (N_19110,N_17613,N_18509);
xnor U19111 (N_19111,N_17792,N_18599);
or U19112 (N_19112,N_17582,N_18339);
or U19113 (N_19113,N_17500,N_18385);
nand U19114 (N_19114,N_18531,N_18595);
xnor U19115 (N_19115,N_18504,N_18319);
and U19116 (N_19116,N_18280,N_17590);
and U19117 (N_19117,N_17687,N_18612);
nor U19118 (N_19118,N_18201,N_18676);
nand U19119 (N_19119,N_18055,N_17864);
and U19120 (N_19120,N_18106,N_18484);
nand U19121 (N_19121,N_18406,N_18512);
xor U19122 (N_19122,N_17844,N_18647);
and U19123 (N_19123,N_18487,N_18425);
and U19124 (N_19124,N_18630,N_17715);
nor U19125 (N_19125,N_18118,N_18629);
nor U19126 (N_19126,N_17938,N_18421);
and U19127 (N_19127,N_17639,N_18404);
nor U19128 (N_19128,N_17504,N_18178);
nand U19129 (N_19129,N_17705,N_18392);
nor U19130 (N_19130,N_17991,N_18285);
nand U19131 (N_19131,N_18202,N_18326);
nor U19132 (N_19132,N_17669,N_18312);
xnor U19133 (N_19133,N_17784,N_18173);
and U19134 (N_19134,N_18242,N_17583);
xor U19135 (N_19135,N_17620,N_18283);
xor U19136 (N_19136,N_17526,N_18103);
and U19137 (N_19137,N_18176,N_17932);
or U19138 (N_19138,N_18481,N_18164);
xnor U19139 (N_19139,N_17598,N_18091);
nor U19140 (N_19140,N_18466,N_18016);
or U19141 (N_19141,N_17985,N_17754);
or U19142 (N_19142,N_18247,N_18634);
or U19143 (N_19143,N_18702,N_17624);
nor U19144 (N_19144,N_17626,N_18031);
nor U19145 (N_19145,N_17536,N_18663);
nor U19146 (N_19146,N_18609,N_17725);
xnor U19147 (N_19147,N_18308,N_18030);
and U19148 (N_19148,N_17753,N_18062);
nand U19149 (N_19149,N_18115,N_17942);
or U19150 (N_19150,N_18315,N_18048);
nand U19151 (N_19151,N_17637,N_17726);
nor U19152 (N_19152,N_18520,N_17892);
nand U19153 (N_19153,N_17824,N_17926);
nor U19154 (N_19154,N_17702,N_18450);
nor U19155 (N_19155,N_17980,N_17538);
nor U19156 (N_19156,N_17552,N_18747);
and U19157 (N_19157,N_18122,N_17534);
nand U19158 (N_19158,N_17852,N_18370);
nand U19159 (N_19159,N_17973,N_18677);
nand U19160 (N_19160,N_17867,N_18723);
nand U19161 (N_19161,N_18430,N_17785);
xor U19162 (N_19162,N_17971,N_17647);
or U19163 (N_19163,N_17861,N_17805);
or U19164 (N_19164,N_18220,N_18185);
or U19165 (N_19165,N_17927,N_18208);
xor U19166 (N_19166,N_18591,N_18002);
and U19167 (N_19167,N_17662,N_17735);
or U19168 (N_19168,N_17760,N_17918);
nor U19169 (N_19169,N_18198,N_17710);
nand U19170 (N_19170,N_18344,N_18255);
xor U19171 (N_19171,N_18235,N_18557);
xnor U19172 (N_19172,N_18097,N_17591);
nor U19173 (N_19173,N_17999,N_18386);
and U19174 (N_19174,N_18154,N_17939);
nor U19175 (N_19175,N_17977,N_18746);
or U19176 (N_19176,N_18073,N_18640);
nor U19177 (N_19177,N_17699,N_18011);
and U19178 (N_19178,N_17542,N_18310);
nand U19179 (N_19179,N_17675,N_18644);
or U19180 (N_19180,N_18275,N_17686);
or U19181 (N_19181,N_18587,N_18365);
xor U19182 (N_19182,N_18015,N_18279);
or U19183 (N_19183,N_18166,N_18687);
nand U19184 (N_19184,N_18318,N_18273);
nor U19185 (N_19185,N_17948,N_18181);
xnor U19186 (N_19186,N_17886,N_17966);
nor U19187 (N_19187,N_18056,N_18205);
nand U19188 (N_19188,N_18424,N_17517);
xnor U19189 (N_19189,N_18656,N_17945);
and U19190 (N_19190,N_18490,N_18053);
nand U19191 (N_19191,N_18659,N_18638);
and U19192 (N_19192,N_18678,N_18135);
nor U19193 (N_19193,N_18673,N_18108);
nand U19194 (N_19194,N_17659,N_17846);
nor U19195 (N_19195,N_18079,N_17545);
or U19196 (N_19196,N_17814,N_18500);
nor U19197 (N_19197,N_17843,N_17996);
or U19198 (N_19198,N_17751,N_18745);
xnor U19199 (N_19199,N_18633,N_17900);
xor U19200 (N_19200,N_18222,N_18372);
and U19201 (N_19201,N_18335,N_18064);
nor U19202 (N_19202,N_18708,N_17713);
nor U19203 (N_19203,N_17518,N_18120);
and U19204 (N_19204,N_17664,N_18260);
nand U19205 (N_19205,N_17554,N_18050);
xnor U19206 (N_19206,N_18395,N_17707);
or U19207 (N_19207,N_18382,N_18699);
nor U19208 (N_19208,N_18491,N_17884);
nor U19209 (N_19209,N_18667,N_17923);
or U19210 (N_19210,N_17721,N_18452);
xor U19211 (N_19211,N_18605,N_18526);
nand U19212 (N_19212,N_18525,N_18474);
or U19213 (N_19213,N_18110,N_18375);
nand U19214 (N_19214,N_18171,N_18705);
xor U19215 (N_19215,N_18561,N_18547);
xnor U19216 (N_19216,N_17941,N_18593);
xor U19217 (N_19217,N_18434,N_18729);
or U19218 (N_19218,N_17871,N_18502);
and U19219 (N_19219,N_18252,N_18136);
nand U19220 (N_19220,N_17916,N_18117);
or U19221 (N_19221,N_18733,N_18139);
xnor U19222 (N_19222,N_17711,N_17576);
nand U19223 (N_19223,N_18196,N_18209);
xnor U19224 (N_19224,N_17851,N_17679);
xnor U19225 (N_19225,N_18084,N_18670);
nor U19226 (N_19226,N_17869,N_17820);
and U19227 (N_19227,N_18231,N_18714);
or U19228 (N_19228,N_18240,N_18101);
or U19229 (N_19229,N_18498,N_17768);
and U19230 (N_19230,N_17838,N_18652);
or U19231 (N_19231,N_18306,N_18534);
xor U19232 (N_19232,N_18680,N_17584);
or U19233 (N_19233,N_18018,N_18157);
xnor U19234 (N_19234,N_18460,N_18660);
or U19235 (N_19235,N_18218,N_17740);
and U19236 (N_19236,N_18397,N_18223);
and U19237 (N_19237,N_17747,N_17525);
nand U19238 (N_19238,N_17502,N_18207);
xnor U19239 (N_19239,N_18316,N_18631);
nand U19240 (N_19240,N_17608,N_18300);
nand U19241 (N_19241,N_17888,N_18210);
nor U19242 (N_19242,N_17821,N_17572);
xor U19243 (N_19243,N_18569,N_18585);
and U19244 (N_19244,N_18414,N_18187);
nand U19245 (N_19245,N_18455,N_18665);
nor U19246 (N_19246,N_17611,N_17847);
and U19247 (N_19247,N_18477,N_18093);
and U19248 (N_19248,N_17958,N_17883);
or U19249 (N_19249,N_17860,N_18276);
or U19250 (N_19250,N_18571,N_17559);
xor U19251 (N_19251,N_18127,N_18618);
xnor U19252 (N_19252,N_18396,N_18734);
nor U19253 (N_19253,N_18709,N_17564);
xnor U19254 (N_19254,N_18088,N_18293);
and U19255 (N_19255,N_18066,N_17988);
nor U19256 (N_19256,N_17606,N_17543);
nand U19257 (N_19257,N_17618,N_18552);
xnor U19258 (N_19258,N_18203,N_17541);
or U19259 (N_19259,N_18636,N_18664);
nand U19260 (N_19260,N_18038,N_17855);
nand U19261 (N_19261,N_18698,N_17731);
and U19262 (N_19262,N_17706,N_18544);
xnor U19263 (N_19263,N_18054,N_17919);
and U19264 (N_19264,N_17651,N_18226);
xnor U19265 (N_19265,N_17976,N_17522);
xor U19266 (N_19266,N_17663,N_18573);
nand U19267 (N_19267,N_18553,N_18267);
nor U19268 (N_19268,N_18125,N_17670);
or U19269 (N_19269,N_18363,N_18560);
or U19270 (N_19270,N_18558,N_17767);
nand U19271 (N_19271,N_18621,N_18256);
xor U19272 (N_19272,N_18536,N_18693);
and U19273 (N_19273,N_18435,N_17905);
nand U19274 (N_19274,N_17986,N_18137);
nor U19275 (N_19275,N_18354,N_17887);
and U19276 (N_19276,N_18328,N_18029);
xor U19277 (N_19277,N_18146,N_18138);
nand U19278 (N_19278,N_17521,N_18473);
nand U19279 (N_19279,N_18570,N_18215);
nor U19280 (N_19280,N_17742,N_17925);
and U19281 (N_19281,N_18026,N_18206);
nand U19282 (N_19282,N_18537,N_18021);
xor U19283 (N_19283,N_17842,N_18368);
xor U19284 (N_19284,N_18542,N_18578);
xor U19285 (N_19285,N_17632,N_18429);
xor U19286 (N_19286,N_18394,N_18682);
nor U19287 (N_19287,N_18221,N_18334);
xnor U19288 (N_19288,N_18214,N_18625);
and U19289 (N_19289,N_18284,N_17763);
and U19290 (N_19290,N_18111,N_18257);
xnor U19291 (N_19291,N_17593,N_18494);
xor U19292 (N_19292,N_17703,N_18728);
nor U19293 (N_19293,N_18188,N_17736);
and U19294 (N_19294,N_17599,N_18155);
nand U19295 (N_19295,N_18701,N_17797);
or U19296 (N_19296,N_18393,N_17808);
xnor U19297 (N_19297,N_18060,N_18467);
and U19298 (N_19298,N_17803,N_18422);
nand U19299 (N_19299,N_18367,N_17897);
and U19300 (N_19300,N_18333,N_18471);
and U19301 (N_19301,N_18448,N_18539);
or U19302 (N_19302,N_17993,N_17815);
and U19303 (N_19303,N_17744,N_17676);
xor U19304 (N_19304,N_18343,N_17811);
nor U19305 (N_19305,N_18707,N_18730);
xnor U19306 (N_19306,N_17964,N_18134);
nand U19307 (N_19307,N_17722,N_18107);
nor U19308 (N_19308,N_18562,N_18383);
xor U19309 (N_19309,N_17700,N_17641);
or U19310 (N_19310,N_18579,N_17562);
xnor U19311 (N_19311,N_17912,N_18213);
xor U19312 (N_19312,N_17630,N_18657);
nand U19313 (N_19313,N_18168,N_18622);
or U19314 (N_19314,N_18611,N_18126);
and U19315 (N_19315,N_18039,N_18426);
xnor U19316 (N_19316,N_18416,N_17621);
or U19317 (N_19317,N_17881,N_18566);
nand U19318 (N_19318,N_18554,N_18436);
xnor U19319 (N_19319,N_18077,N_17694);
nand U19320 (N_19320,N_17975,N_18620);
nand U19321 (N_19321,N_17556,N_18362);
nand U19322 (N_19322,N_18299,N_18140);
nand U19323 (N_19323,N_17551,N_18246);
xnor U19324 (N_19324,N_18524,N_17936);
nor U19325 (N_19325,N_17712,N_17586);
and U19326 (N_19326,N_17692,N_18340);
nor U19327 (N_19327,N_17548,N_18303);
nand U19328 (N_19328,N_18193,N_17743);
and U19329 (N_19329,N_18096,N_17786);
nand U19330 (N_19330,N_17514,N_18234);
xor U19331 (N_19331,N_17896,N_18533);
or U19332 (N_19332,N_18683,N_18532);
nor U19333 (N_19333,N_17746,N_18345);
xor U19334 (N_19334,N_18006,N_18551);
nand U19335 (N_19335,N_17655,N_18265);
xor U19336 (N_19336,N_18469,N_18350);
nand U19337 (N_19337,N_18313,N_18540);
and U19338 (N_19338,N_18387,N_17634);
nand U19339 (N_19339,N_18366,N_18180);
or U19340 (N_19340,N_17567,N_17574);
nand U19341 (N_19341,N_17839,N_17956);
and U19342 (N_19342,N_17565,N_17607);
nor U19343 (N_19343,N_17924,N_18075);
and U19344 (N_19344,N_18258,N_18574);
nor U19345 (N_19345,N_17701,N_18423);
xnor U19346 (N_19346,N_18113,N_18130);
or U19347 (N_19347,N_18085,N_17623);
or U19348 (N_19348,N_17920,N_17970);
nor U19349 (N_19349,N_17950,N_17906);
or U19350 (N_19350,N_17849,N_18277);
nor U19351 (N_19351,N_17761,N_18402);
or U19352 (N_19352,N_18261,N_18177);
nor U19353 (N_19353,N_17909,N_17894);
xnor U19354 (N_19354,N_17550,N_18482);
xnor U19355 (N_19355,N_17539,N_18000);
and U19356 (N_19356,N_18666,N_18583);
nand U19357 (N_19357,N_18454,N_18301);
and U19358 (N_19358,N_18398,N_18336);
or U19359 (N_19359,N_17874,N_17795);
xor U19360 (N_19360,N_18024,N_17778);
and U19361 (N_19361,N_18003,N_17828);
nor U19362 (N_19362,N_17825,N_17776);
xor U19363 (N_19363,N_18470,N_18014);
or U19364 (N_19364,N_18358,N_17625);
or U19365 (N_19365,N_17661,N_18646);
xor U19366 (N_19366,N_17914,N_18156);
nand U19367 (N_19367,N_18528,N_18495);
and U19368 (N_19368,N_17830,N_17524);
xnor U19369 (N_19369,N_18722,N_18359);
or U19370 (N_19370,N_18380,N_17757);
or U19371 (N_19371,N_18568,N_17772);
and U19372 (N_19372,N_17560,N_17859);
nand U19373 (N_19373,N_17697,N_18251);
nand U19374 (N_19374,N_18674,N_17671);
nand U19375 (N_19375,N_17555,N_17790);
and U19376 (N_19376,N_18257,N_18457);
nand U19377 (N_19377,N_17988,N_18094);
xnor U19378 (N_19378,N_17840,N_17632);
nand U19379 (N_19379,N_17960,N_18224);
xor U19380 (N_19380,N_17570,N_17632);
nand U19381 (N_19381,N_18661,N_17657);
nand U19382 (N_19382,N_17713,N_18044);
or U19383 (N_19383,N_18159,N_18623);
nand U19384 (N_19384,N_18618,N_17597);
or U19385 (N_19385,N_18056,N_17842);
nand U19386 (N_19386,N_18359,N_17500);
and U19387 (N_19387,N_18430,N_17835);
xor U19388 (N_19388,N_18482,N_17795);
xnor U19389 (N_19389,N_17544,N_18159);
nand U19390 (N_19390,N_17649,N_17887);
xor U19391 (N_19391,N_18489,N_18223);
nand U19392 (N_19392,N_18502,N_18563);
or U19393 (N_19393,N_17522,N_17781);
and U19394 (N_19394,N_18274,N_18036);
nor U19395 (N_19395,N_17665,N_17912);
or U19396 (N_19396,N_18060,N_17877);
or U19397 (N_19397,N_17613,N_17904);
or U19398 (N_19398,N_17908,N_18351);
and U19399 (N_19399,N_17838,N_18023);
and U19400 (N_19400,N_18539,N_18247);
nand U19401 (N_19401,N_18236,N_17790);
and U19402 (N_19402,N_18092,N_18505);
and U19403 (N_19403,N_18097,N_17517);
xor U19404 (N_19404,N_18206,N_17585);
xnor U19405 (N_19405,N_18257,N_17715);
and U19406 (N_19406,N_18594,N_17915);
or U19407 (N_19407,N_17665,N_18002);
and U19408 (N_19408,N_17551,N_18719);
xor U19409 (N_19409,N_17846,N_18393);
and U19410 (N_19410,N_18018,N_17741);
xor U19411 (N_19411,N_17548,N_18059);
and U19412 (N_19412,N_18079,N_18037);
nand U19413 (N_19413,N_17853,N_17776);
nand U19414 (N_19414,N_18669,N_17908);
xor U19415 (N_19415,N_18624,N_17621);
and U19416 (N_19416,N_18586,N_18038);
nor U19417 (N_19417,N_18562,N_17685);
or U19418 (N_19418,N_18250,N_18098);
nor U19419 (N_19419,N_18070,N_17992);
nand U19420 (N_19420,N_18709,N_18273);
xor U19421 (N_19421,N_17740,N_17933);
or U19422 (N_19422,N_17659,N_17647);
nand U19423 (N_19423,N_18165,N_17994);
xor U19424 (N_19424,N_18643,N_18354);
and U19425 (N_19425,N_17840,N_18418);
or U19426 (N_19426,N_18182,N_17623);
and U19427 (N_19427,N_17782,N_18016);
or U19428 (N_19428,N_18124,N_17872);
nand U19429 (N_19429,N_17698,N_17711);
or U19430 (N_19430,N_18190,N_18497);
nor U19431 (N_19431,N_18048,N_17823);
and U19432 (N_19432,N_17943,N_17579);
or U19433 (N_19433,N_17852,N_18644);
and U19434 (N_19434,N_17727,N_17986);
xor U19435 (N_19435,N_18564,N_18639);
nand U19436 (N_19436,N_18019,N_18028);
xor U19437 (N_19437,N_17842,N_18428);
nand U19438 (N_19438,N_17854,N_17816);
nor U19439 (N_19439,N_18250,N_18339);
nor U19440 (N_19440,N_18424,N_18255);
nand U19441 (N_19441,N_18146,N_18402);
or U19442 (N_19442,N_18285,N_18415);
nor U19443 (N_19443,N_18548,N_18423);
nand U19444 (N_19444,N_18057,N_18161);
nor U19445 (N_19445,N_17998,N_18399);
or U19446 (N_19446,N_17509,N_18210);
or U19447 (N_19447,N_18513,N_17835);
and U19448 (N_19448,N_18135,N_18193);
nor U19449 (N_19449,N_17981,N_18360);
nand U19450 (N_19450,N_18283,N_17900);
xor U19451 (N_19451,N_18262,N_17741);
or U19452 (N_19452,N_17727,N_18184);
and U19453 (N_19453,N_18230,N_18726);
xor U19454 (N_19454,N_18545,N_17701);
and U19455 (N_19455,N_18287,N_18564);
xnor U19456 (N_19456,N_17789,N_17799);
nand U19457 (N_19457,N_18710,N_18061);
nor U19458 (N_19458,N_18633,N_18508);
xnor U19459 (N_19459,N_18366,N_17683);
and U19460 (N_19460,N_18524,N_18084);
nand U19461 (N_19461,N_17859,N_17834);
nor U19462 (N_19462,N_18282,N_18329);
and U19463 (N_19463,N_17908,N_18088);
or U19464 (N_19464,N_17575,N_18418);
or U19465 (N_19465,N_18669,N_18522);
nand U19466 (N_19466,N_18177,N_18187);
xor U19467 (N_19467,N_18729,N_17791);
or U19468 (N_19468,N_17849,N_18429);
or U19469 (N_19469,N_18486,N_17824);
nand U19470 (N_19470,N_17737,N_17924);
and U19471 (N_19471,N_17885,N_18342);
nor U19472 (N_19472,N_17640,N_17723);
nand U19473 (N_19473,N_18422,N_18290);
nand U19474 (N_19474,N_17832,N_18543);
xor U19475 (N_19475,N_18389,N_17506);
or U19476 (N_19476,N_18504,N_18172);
and U19477 (N_19477,N_18034,N_18638);
xnor U19478 (N_19478,N_18403,N_18746);
nand U19479 (N_19479,N_18154,N_17958);
nor U19480 (N_19480,N_18321,N_17650);
xnor U19481 (N_19481,N_17544,N_18261);
or U19482 (N_19482,N_17707,N_17917);
xnor U19483 (N_19483,N_17660,N_18728);
nand U19484 (N_19484,N_18261,N_18023);
or U19485 (N_19485,N_18032,N_18730);
nand U19486 (N_19486,N_18696,N_18437);
nand U19487 (N_19487,N_18081,N_18305);
or U19488 (N_19488,N_17665,N_18378);
or U19489 (N_19489,N_18304,N_18366);
nor U19490 (N_19490,N_17650,N_17733);
nand U19491 (N_19491,N_18613,N_17658);
xnor U19492 (N_19492,N_17571,N_17781);
nor U19493 (N_19493,N_17859,N_17755);
nand U19494 (N_19494,N_17610,N_18046);
nand U19495 (N_19495,N_17660,N_18392);
xnor U19496 (N_19496,N_18498,N_18268);
or U19497 (N_19497,N_18698,N_18357);
nor U19498 (N_19498,N_18106,N_17631);
xor U19499 (N_19499,N_17852,N_17878);
nand U19500 (N_19500,N_18389,N_17627);
and U19501 (N_19501,N_18489,N_18695);
or U19502 (N_19502,N_18395,N_18573);
nand U19503 (N_19503,N_18391,N_17568);
nand U19504 (N_19504,N_18160,N_18091);
or U19505 (N_19505,N_17644,N_18063);
nand U19506 (N_19506,N_18243,N_17752);
nor U19507 (N_19507,N_18092,N_18648);
nor U19508 (N_19508,N_17603,N_18447);
nor U19509 (N_19509,N_17534,N_18162);
or U19510 (N_19510,N_17761,N_18613);
nor U19511 (N_19511,N_17861,N_18004);
nand U19512 (N_19512,N_18462,N_18433);
or U19513 (N_19513,N_17780,N_17891);
nor U19514 (N_19514,N_18602,N_18411);
or U19515 (N_19515,N_18033,N_18231);
and U19516 (N_19516,N_18280,N_18500);
or U19517 (N_19517,N_18072,N_18354);
xnor U19518 (N_19518,N_18519,N_18369);
xnor U19519 (N_19519,N_17846,N_18730);
nor U19520 (N_19520,N_17682,N_17811);
nand U19521 (N_19521,N_17820,N_18371);
or U19522 (N_19522,N_18563,N_17726);
and U19523 (N_19523,N_17532,N_17706);
nor U19524 (N_19524,N_18728,N_17849);
or U19525 (N_19525,N_17505,N_18159);
nor U19526 (N_19526,N_18604,N_18334);
xor U19527 (N_19527,N_18332,N_18244);
xor U19528 (N_19528,N_18599,N_18038);
or U19529 (N_19529,N_17906,N_18291);
xnor U19530 (N_19530,N_17876,N_18436);
nand U19531 (N_19531,N_18058,N_18576);
xnor U19532 (N_19532,N_18701,N_18499);
xor U19533 (N_19533,N_18505,N_18158);
nor U19534 (N_19534,N_18249,N_18353);
nor U19535 (N_19535,N_17696,N_17561);
nand U19536 (N_19536,N_18589,N_17830);
xor U19537 (N_19537,N_17629,N_17645);
nand U19538 (N_19538,N_18697,N_17740);
and U19539 (N_19539,N_17895,N_17552);
xor U19540 (N_19540,N_18510,N_17859);
nor U19541 (N_19541,N_17837,N_18486);
nand U19542 (N_19542,N_17799,N_18062);
nand U19543 (N_19543,N_18453,N_17786);
and U19544 (N_19544,N_18373,N_17733);
or U19545 (N_19545,N_17727,N_18167);
or U19546 (N_19546,N_17703,N_17560);
or U19547 (N_19547,N_18474,N_18048);
nand U19548 (N_19548,N_17854,N_17732);
and U19549 (N_19549,N_17762,N_17949);
nor U19550 (N_19550,N_17628,N_18568);
nand U19551 (N_19551,N_18643,N_18177);
or U19552 (N_19552,N_18634,N_18050);
and U19553 (N_19553,N_18468,N_18264);
xnor U19554 (N_19554,N_17681,N_18612);
nand U19555 (N_19555,N_18262,N_18696);
or U19556 (N_19556,N_17819,N_17873);
nor U19557 (N_19557,N_18695,N_17806);
or U19558 (N_19558,N_18278,N_18080);
nor U19559 (N_19559,N_17942,N_17995);
xor U19560 (N_19560,N_18535,N_18146);
nor U19561 (N_19561,N_18085,N_18747);
or U19562 (N_19562,N_17775,N_18240);
nand U19563 (N_19563,N_18586,N_18718);
or U19564 (N_19564,N_17608,N_18382);
xnor U19565 (N_19565,N_18722,N_18337);
nand U19566 (N_19566,N_17608,N_18483);
nor U19567 (N_19567,N_17875,N_17705);
nand U19568 (N_19568,N_17695,N_18504);
nor U19569 (N_19569,N_17916,N_18125);
or U19570 (N_19570,N_17512,N_17837);
nand U19571 (N_19571,N_17649,N_18378);
and U19572 (N_19572,N_18176,N_18486);
or U19573 (N_19573,N_17864,N_18394);
xor U19574 (N_19574,N_17687,N_18506);
nor U19575 (N_19575,N_18711,N_18705);
nand U19576 (N_19576,N_17753,N_18116);
nor U19577 (N_19577,N_18305,N_17705);
and U19578 (N_19578,N_17581,N_18666);
nor U19579 (N_19579,N_17794,N_18328);
and U19580 (N_19580,N_18359,N_18619);
and U19581 (N_19581,N_17947,N_18382);
xor U19582 (N_19582,N_18635,N_18623);
or U19583 (N_19583,N_18288,N_18734);
nor U19584 (N_19584,N_18729,N_17775);
xor U19585 (N_19585,N_17536,N_18331);
nor U19586 (N_19586,N_17691,N_17573);
xor U19587 (N_19587,N_17716,N_17936);
nor U19588 (N_19588,N_18663,N_18045);
nor U19589 (N_19589,N_18454,N_18191);
xor U19590 (N_19590,N_17551,N_17789);
xnor U19591 (N_19591,N_18415,N_17973);
and U19592 (N_19592,N_17904,N_17505);
and U19593 (N_19593,N_18631,N_17780);
or U19594 (N_19594,N_18669,N_18206);
and U19595 (N_19595,N_18070,N_17759);
nand U19596 (N_19596,N_18360,N_18588);
xnor U19597 (N_19597,N_18692,N_17643);
nand U19598 (N_19598,N_18549,N_18284);
nand U19599 (N_19599,N_18156,N_18517);
and U19600 (N_19600,N_17933,N_17705);
xor U19601 (N_19601,N_18720,N_18478);
or U19602 (N_19602,N_18688,N_18081);
nand U19603 (N_19603,N_18143,N_18512);
nor U19604 (N_19604,N_18571,N_18093);
xnor U19605 (N_19605,N_18733,N_18337);
and U19606 (N_19606,N_18273,N_17701);
xnor U19607 (N_19607,N_18652,N_17790);
xor U19608 (N_19608,N_17533,N_18285);
and U19609 (N_19609,N_18684,N_18105);
nand U19610 (N_19610,N_18218,N_18162);
and U19611 (N_19611,N_18224,N_17567);
xnor U19612 (N_19612,N_18603,N_17959);
xnor U19613 (N_19613,N_17512,N_17720);
xnor U19614 (N_19614,N_18097,N_17790);
and U19615 (N_19615,N_18619,N_18732);
and U19616 (N_19616,N_18230,N_18484);
and U19617 (N_19617,N_18266,N_18676);
nand U19618 (N_19618,N_17520,N_18370);
nand U19619 (N_19619,N_18622,N_18713);
or U19620 (N_19620,N_17598,N_17515);
nand U19621 (N_19621,N_18263,N_17889);
nor U19622 (N_19622,N_18563,N_18493);
xnor U19623 (N_19623,N_18349,N_17642);
nor U19624 (N_19624,N_18076,N_18743);
nor U19625 (N_19625,N_18369,N_18508);
xnor U19626 (N_19626,N_18214,N_17836);
xor U19627 (N_19627,N_17770,N_18621);
and U19628 (N_19628,N_18185,N_18439);
xor U19629 (N_19629,N_17599,N_18614);
or U19630 (N_19630,N_18242,N_18674);
and U19631 (N_19631,N_18616,N_18283);
nand U19632 (N_19632,N_17906,N_17516);
and U19633 (N_19633,N_18463,N_18325);
nand U19634 (N_19634,N_17869,N_18607);
nand U19635 (N_19635,N_18379,N_17808);
xnor U19636 (N_19636,N_17874,N_17761);
and U19637 (N_19637,N_18704,N_18475);
and U19638 (N_19638,N_18387,N_17908);
nand U19639 (N_19639,N_17852,N_18241);
xnor U19640 (N_19640,N_17847,N_17842);
xor U19641 (N_19641,N_18637,N_18062);
and U19642 (N_19642,N_17742,N_18124);
nand U19643 (N_19643,N_17592,N_17775);
nor U19644 (N_19644,N_17726,N_17980);
or U19645 (N_19645,N_18410,N_18557);
and U19646 (N_19646,N_18046,N_18034);
xnor U19647 (N_19647,N_18630,N_18692);
xnor U19648 (N_19648,N_17732,N_18011);
and U19649 (N_19649,N_18714,N_18253);
nor U19650 (N_19650,N_17522,N_18109);
nor U19651 (N_19651,N_18457,N_17622);
xor U19652 (N_19652,N_17800,N_17775);
nand U19653 (N_19653,N_18662,N_17921);
and U19654 (N_19654,N_18188,N_17586);
and U19655 (N_19655,N_18608,N_18624);
xnor U19656 (N_19656,N_17652,N_17960);
nor U19657 (N_19657,N_18430,N_18610);
or U19658 (N_19658,N_17933,N_17610);
nand U19659 (N_19659,N_17964,N_18720);
xnor U19660 (N_19660,N_18671,N_17923);
nand U19661 (N_19661,N_17793,N_17646);
or U19662 (N_19662,N_17620,N_18146);
nor U19663 (N_19663,N_17971,N_17608);
nand U19664 (N_19664,N_17903,N_18749);
xor U19665 (N_19665,N_18448,N_18611);
and U19666 (N_19666,N_18089,N_17792);
xor U19667 (N_19667,N_17942,N_18541);
and U19668 (N_19668,N_18034,N_18649);
xor U19669 (N_19669,N_17570,N_18184);
and U19670 (N_19670,N_18015,N_18720);
xor U19671 (N_19671,N_18383,N_18590);
or U19672 (N_19672,N_17647,N_18706);
or U19673 (N_19673,N_18178,N_18285);
and U19674 (N_19674,N_18410,N_18283);
and U19675 (N_19675,N_17979,N_18727);
and U19676 (N_19676,N_18129,N_17547);
nor U19677 (N_19677,N_17585,N_17533);
nand U19678 (N_19678,N_18363,N_18640);
and U19679 (N_19679,N_18064,N_17776);
nor U19680 (N_19680,N_17823,N_17710);
and U19681 (N_19681,N_18096,N_18016);
and U19682 (N_19682,N_17828,N_18619);
or U19683 (N_19683,N_18005,N_17836);
or U19684 (N_19684,N_17818,N_17532);
xor U19685 (N_19685,N_18101,N_18344);
nor U19686 (N_19686,N_17930,N_17663);
or U19687 (N_19687,N_17716,N_17695);
or U19688 (N_19688,N_18042,N_17514);
or U19689 (N_19689,N_18712,N_18003);
nand U19690 (N_19690,N_17699,N_17870);
xor U19691 (N_19691,N_17795,N_17546);
and U19692 (N_19692,N_18186,N_18231);
nor U19693 (N_19693,N_18208,N_17871);
xor U19694 (N_19694,N_17890,N_18586);
and U19695 (N_19695,N_17957,N_18371);
and U19696 (N_19696,N_18184,N_18535);
nand U19697 (N_19697,N_18368,N_17980);
xnor U19698 (N_19698,N_18597,N_18639);
or U19699 (N_19699,N_18334,N_18315);
and U19700 (N_19700,N_18709,N_17935);
nand U19701 (N_19701,N_18383,N_17734);
or U19702 (N_19702,N_17749,N_17913);
nor U19703 (N_19703,N_17537,N_18716);
xor U19704 (N_19704,N_18144,N_17530);
or U19705 (N_19705,N_17583,N_18719);
nand U19706 (N_19706,N_18396,N_17502);
xnor U19707 (N_19707,N_18479,N_17969);
and U19708 (N_19708,N_17813,N_18679);
xor U19709 (N_19709,N_18162,N_18149);
xor U19710 (N_19710,N_18065,N_17758);
xor U19711 (N_19711,N_18271,N_17617);
nand U19712 (N_19712,N_18301,N_17913);
and U19713 (N_19713,N_18495,N_17726);
xnor U19714 (N_19714,N_17553,N_18702);
nor U19715 (N_19715,N_17879,N_18042);
and U19716 (N_19716,N_17875,N_17864);
nor U19717 (N_19717,N_17862,N_17588);
and U19718 (N_19718,N_18453,N_18575);
xnor U19719 (N_19719,N_17853,N_18716);
and U19720 (N_19720,N_18228,N_18473);
xor U19721 (N_19721,N_18681,N_17812);
and U19722 (N_19722,N_18725,N_18547);
or U19723 (N_19723,N_17556,N_18201);
nand U19724 (N_19724,N_18607,N_18088);
nor U19725 (N_19725,N_17899,N_17750);
and U19726 (N_19726,N_18484,N_18493);
xor U19727 (N_19727,N_18734,N_18592);
xor U19728 (N_19728,N_17757,N_18033);
or U19729 (N_19729,N_17679,N_17696);
nor U19730 (N_19730,N_17738,N_17692);
or U19731 (N_19731,N_18371,N_17801);
nor U19732 (N_19732,N_17795,N_17777);
nor U19733 (N_19733,N_17749,N_17523);
xor U19734 (N_19734,N_17721,N_18226);
and U19735 (N_19735,N_18571,N_17508);
nand U19736 (N_19736,N_18005,N_18387);
nand U19737 (N_19737,N_17520,N_18641);
nand U19738 (N_19738,N_18362,N_18400);
xor U19739 (N_19739,N_17848,N_17773);
nand U19740 (N_19740,N_18293,N_18030);
nor U19741 (N_19741,N_18100,N_18305);
or U19742 (N_19742,N_17655,N_18695);
xor U19743 (N_19743,N_18143,N_17724);
or U19744 (N_19744,N_18531,N_17661);
nand U19745 (N_19745,N_17987,N_18114);
xor U19746 (N_19746,N_17566,N_18538);
and U19747 (N_19747,N_18284,N_18658);
or U19748 (N_19748,N_18656,N_18186);
nand U19749 (N_19749,N_17586,N_17896);
and U19750 (N_19750,N_18150,N_18179);
xnor U19751 (N_19751,N_17644,N_17793);
nand U19752 (N_19752,N_17790,N_18057);
nor U19753 (N_19753,N_17703,N_17821);
nor U19754 (N_19754,N_18523,N_18490);
nor U19755 (N_19755,N_18432,N_17790);
or U19756 (N_19756,N_18267,N_18406);
and U19757 (N_19757,N_17563,N_18488);
and U19758 (N_19758,N_18487,N_18237);
nand U19759 (N_19759,N_18520,N_18518);
xor U19760 (N_19760,N_17892,N_17704);
nand U19761 (N_19761,N_18281,N_18667);
nor U19762 (N_19762,N_17585,N_17801);
and U19763 (N_19763,N_18240,N_18575);
nand U19764 (N_19764,N_17651,N_17728);
or U19765 (N_19765,N_18513,N_18709);
or U19766 (N_19766,N_18032,N_17787);
and U19767 (N_19767,N_18000,N_18275);
or U19768 (N_19768,N_18696,N_17957);
nor U19769 (N_19769,N_17779,N_18513);
nor U19770 (N_19770,N_18407,N_17998);
and U19771 (N_19771,N_17819,N_18616);
nor U19772 (N_19772,N_17861,N_17939);
xor U19773 (N_19773,N_18653,N_18039);
nor U19774 (N_19774,N_18713,N_17564);
xor U19775 (N_19775,N_18354,N_17808);
nor U19776 (N_19776,N_18444,N_17937);
xnor U19777 (N_19777,N_18254,N_18429);
nor U19778 (N_19778,N_18198,N_18031);
and U19779 (N_19779,N_17929,N_18242);
nor U19780 (N_19780,N_17839,N_18080);
nor U19781 (N_19781,N_18633,N_17688);
or U19782 (N_19782,N_18134,N_18606);
and U19783 (N_19783,N_18287,N_18708);
or U19784 (N_19784,N_18089,N_17694);
xnor U19785 (N_19785,N_18500,N_17697);
and U19786 (N_19786,N_17796,N_18001);
nand U19787 (N_19787,N_18011,N_18033);
xor U19788 (N_19788,N_17783,N_17830);
xor U19789 (N_19789,N_18703,N_18710);
xnor U19790 (N_19790,N_17649,N_18456);
and U19791 (N_19791,N_18440,N_17514);
xnor U19792 (N_19792,N_18618,N_17951);
and U19793 (N_19793,N_18499,N_18669);
nand U19794 (N_19794,N_17740,N_17605);
and U19795 (N_19795,N_17833,N_18065);
and U19796 (N_19796,N_17500,N_17675);
nor U19797 (N_19797,N_18631,N_18200);
xor U19798 (N_19798,N_18574,N_17566);
and U19799 (N_19799,N_17724,N_17904);
nand U19800 (N_19800,N_18467,N_18003);
and U19801 (N_19801,N_18554,N_17945);
xnor U19802 (N_19802,N_17765,N_17817);
or U19803 (N_19803,N_17566,N_18651);
and U19804 (N_19804,N_18227,N_17521);
nor U19805 (N_19805,N_18403,N_17831);
nand U19806 (N_19806,N_18411,N_18471);
and U19807 (N_19807,N_17913,N_18733);
nor U19808 (N_19808,N_18228,N_17755);
nand U19809 (N_19809,N_18066,N_17609);
nand U19810 (N_19810,N_18406,N_17878);
nand U19811 (N_19811,N_17947,N_17827);
nor U19812 (N_19812,N_18043,N_17938);
and U19813 (N_19813,N_18065,N_18022);
nor U19814 (N_19814,N_18698,N_17648);
nor U19815 (N_19815,N_18274,N_18451);
nand U19816 (N_19816,N_18346,N_17638);
nor U19817 (N_19817,N_18101,N_18366);
nand U19818 (N_19818,N_17718,N_18066);
xnor U19819 (N_19819,N_18375,N_18344);
and U19820 (N_19820,N_18562,N_17972);
nand U19821 (N_19821,N_17802,N_17743);
and U19822 (N_19822,N_18100,N_17557);
xnor U19823 (N_19823,N_17788,N_17604);
xor U19824 (N_19824,N_18350,N_17879);
nand U19825 (N_19825,N_17902,N_18196);
nor U19826 (N_19826,N_17948,N_17968);
or U19827 (N_19827,N_18553,N_18435);
and U19828 (N_19828,N_17710,N_18682);
or U19829 (N_19829,N_17601,N_18266);
nand U19830 (N_19830,N_18334,N_17639);
and U19831 (N_19831,N_17773,N_18450);
xnor U19832 (N_19832,N_17640,N_18711);
xor U19833 (N_19833,N_18163,N_17771);
nor U19834 (N_19834,N_18477,N_18415);
xor U19835 (N_19835,N_18295,N_18440);
or U19836 (N_19836,N_17910,N_18426);
nor U19837 (N_19837,N_18514,N_18272);
nor U19838 (N_19838,N_18170,N_18342);
or U19839 (N_19839,N_18447,N_18644);
xnor U19840 (N_19840,N_18269,N_17507);
xnor U19841 (N_19841,N_18155,N_18472);
nor U19842 (N_19842,N_18337,N_17816);
xor U19843 (N_19843,N_18423,N_18409);
xnor U19844 (N_19844,N_18633,N_18614);
nand U19845 (N_19845,N_17920,N_18214);
xnor U19846 (N_19846,N_18734,N_17531);
nand U19847 (N_19847,N_18522,N_17558);
nor U19848 (N_19848,N_17776,N_18547);
xor U19849 (N_19849,N_18476,N_18744);
nor U19850 (N_19850,N_17876,N_17884);
nor U19851 (N_19851,N_18309,N_18277);
nor U19852 (N_19852,N_17790,N_18709);
and U19853 (N_19853,N_18616,N_17829);
nand U19854 (N_19854,N_18640,N_18685);
and U19855 (N_19855,N_17963,N_17897);
xnor U19856 (N_19856,N_18301,N_17839);
xnor U19857 (N_19857,N_17963,N_18003);
xor U19858 (N_19858,N_17766,N_17753);
nor U19859 (N_19859,N_17596,N_18461);
xnor U19860 (N_19860,N_17966,N_18182);
nand U19861 (N_19861,N_18152,N_17691);
or U19862 (N_19862,N_18594,N_18105);
nand U19863 (N_19863,N_18224,N_18360);
or U19864 (N_19864,N_17865,N_18701);
xnor U19865 (N_19865,N_17710,N_18013);
and U19866 (N_19866,N_18721,N_18128);
xor U19867 (N_19867,N_18345,N_17996);
nor U19868 (N_19868,N_18488,N_17658);
xnor U19869 (N_19869,N_18747,N_18702);
nor U19870 (N_19870,N_17594,N_18385);
or U19871 (N_19871,N_18545,N_18365);
and U19872 (N_19872,N_18152,N_17749);
nor U19873 (N_19873,N_17846,N_17571);
or U19874 (N_19874,N_18532,N_17901);
or U19875 (N_19875,N_17712,N_17564);
nor U19876 (N_19876,N_18292,N_17794);
nor U19877 (N_19877,N_18361,N_17857);
xor U19878 (N_19878,N_18093,N_18055);
and U19879 (N_19879,N_17557,N_17569);
or U19880 (N_19880,N_18469,N_18062);
and U19881 (N_19881,N_17957,N_18621);
nor U19882 (N_19882,N_18134,N_17966);
or U19883 (N_19883,N_18348,N_18666);
nor U19884 (N_19884,N_17657,N_18734);
nand U19885 (N_19885,N_18081,N_18247);
nand U19886 (N_19886,N_17686,N_17810);
nor U19887 (N_19887,N_18332,N_18219);
xor U19888 (N_19888,N_17564,N_18120);
nand U19889 (N_19889,N_18522,N_17901);
nand U19890 (N_19890,N_18487,N_17693);
or U19891 (N_19891,N_18427,N_17683);
and U19892 (N_19892,N_18375,N_18028);
or U19893 (N_19893,N_17627,N_18338);
nor U19894 (N_19894,N_18602,N_17805);
and U19895 (N_19895,N_17635,N_18026);
xnor U19896 (N_19896,N_18603,N_18052);
or U19897 (N_19897,N_17525,N_18621);
xnor U19898 (N_19898,N_18639,N_18661);
nor U19899 (N_19899,N_18329,N_17627);
and U19900 (N_19900,N_18680,N_18225);
nor U19901 (N_19901,N_18514,N_17924);
xor U19902 (N_19902,N_17802,N_17871);
nor U19903 (N_19903,N_18109,N_18081);
xnor U19904 (N_19904,N_17665,N_17877);
xnor U19905 (N_19905,N_17820,N_18738);
or U19906 (N_19906,N_17816,N_17967);
xor U19907 (N_19907,N_18581,N_18453);
nor U19908 (N_19908,N_18468,N_17733);
nand U19909 (N_19909,N_17916,N_18572);
xnor U19910 (N_19910,N_18378,N_18430);
and U19911 (N_19911,N_17521,N_17707);
xor U19912 (N_19912,N_17748,N_18091);
or U19913 (N_19913,N_18257,N_18382);
xor U19914 (N_19914,N_17738,N_17590);
nand U19915 (N_19915,N_18543,N_18087);
xor U19916 (N_19916,N_18122,N_18289);
xor U19917 (N_19917,N_18113,N_17937);
and U19918 (N_19918,N_18491,N_17751);
nor U19919 (N_19919,N_17706,N_18280);
or U19920 (N_19920,N_17565,N_18643);
nor U19921 (N_19921,N_18449,N_17965);
nand U19922 (N_19922,N_18735,N_18689);
nand U19923 (N_19923,N_18169,N_18589);
and U19924 (N_19924,N_18647,N_18666);
nand U19925 (N_19925,N_18330,N_18635);
nand U19926 (N_19926,N_18501,N_18627);
and U19927 (N_19927,N_17911,N_18261);
nor U19928 (N_19928,N_17542,N_18060);
xnor U19929 (N_19929,N_17865,N_17722);
nor U19930 (N_19930,N_17848,N_18280);
and U19931 (N_19931,N_18348,N_18190);
and U19932 (N_19932,N_18582,N_18333);
nand U19933 (N_19933,N_18339,N_17988);
nor U19934 (N_19934,N_18062,N_18548);
and U19935 (N_19935,N_18480,N_17721);
or U19936 (N_19936,N_17668,N_18580);
nor U19937 (N_19937,N_18100,N_17615);
nand U19938 (N_19938,N_18446,N_18530);
nor U19939 (N_19939,N_17753,N_17611);
and U19940 (N_19940,N_18359,N_18430);
xor U19941 (N_19941,N_17795,N_18449);
or U19942 (N_19942,N_18651,N_17986);
nand U19943 (N_19943,N_18674,N_17666);
and U19944 (N_19944,N_18511,N_17766);
or U19945 (N_19945,N_18718,N_17523);
nand U19946 (N_19946,N_17922,N_18199);
nand U19947 (N_19947,N_18640,N_18300);
xor U19948 (N_19948,N_17916,N_17984);
nand U19949 (N_19949,N_17955,N_18520);
nand U19950 (N_19950,N_17655,N_18669);
and U19951 (N_19951,N_17740,N_18108);
or U19952 (N_19952,N_18360,N_18580);
nand U19953 (N_19953,N_17640,N_17500);
nor U19954 (N_19954,N_17631,N_18602);
nand U19955 (N_19955,N_18275,N_18587);
nor U19956 (N_19956,N_18017,N_18485);
nor U19957 (N_19957,N_18314,N_17582);
and U19958 (N_19958,N_17771,N_18550);
xnor U19959 (N_19959,N_17785,N_18180);
xor U19960 (N_19960,N_17630,N_18349);
nand U19961 (N_19961,N_17620,N_17860);
xnor U19962 (N_19962,N_17999,N_18574);
or U19963 (N_19963,N_18314,N_17708);
and U19964 (N_19964,N_17612,N_18632);
nand U19965 (N_19965,N_18492,N_17743);
nor U19966 (N_19966,N_17713,N_17608);
xor U19967 (N_19967,N_17933,N_18109);
and U19968 (N_19968,N_17765,N_17707);
xnor U19969 (N_19969,N_18089,N_17930);
nor U19970 (N_19970,N_17945,N_18423);
and U19971 (N_19971,N_17956,N_17693);
nand U19972 (N_19972,N_18649,N_17563);
nand U19973 (N_19973,N_18586,N_17640);
nor U19974 (N_19974,N_17523,N_17577);
nand U19975 (N_19975,N_18132,N_18390);
nor U19976 (N_19976,N_17612,N_18683);
xor U19977 (N_19977,N_17568,N_18698);
nor U19978 (N_19978,N_18485,N_17977);
nor U19979 (N_19979,N_18121,N_18047);
nand U19980 (N_19980,N_18558,N_17588);
or U19981 (N_19981,N_18028,N_18198);
nor U19982 (N_19982,N_17781,N_18121);
nor U19983 (N_19983,N_17593,N_17548);
xnor U19984 (N_19984,N_17653,N_18021);
xor U19985 (N_19985,N_18002,N_17997);
xor U19986 (N_19986,N_18419,N_17596);
nor U19987 (N_19987,N_17564,N_17540);
nand U19988 (N_19988,N_17547,N_18665);
xnor U19989 (N_19989,N_17591,N_18223);
xnor U19990 (N_19990,N_18194,N_18688);
or U19991 (N_19991,N_18628,N_18483);
nand U19992 (N_19992,N_18021,N_18039);
or U19993 (N_19993,N_18336,N_17547);
nor U19994 (N_19994,N_17798,N_18437);
xnor U19995 (N_19995,N_18732,N_17600);
nand U19996 (N_19996,N_17659,N_18475);
or U19997 (N_19997,N_18302,N_18398);
nand U19998 (N_19998,N_17643,N_18427);
or U19999 (N_19999,N_18653,N_18014);
nor U20000 (N_20000,N_19736,N_19152);
nor U20001 (N_20001,N_19934,N_19318);
xor U20002 (N_20002,N_19267,N_19630);
nor U20003 (N_20003,N_19916,N_18919);
and U20004 (N_20004,N_19082,N_19748);
nor U20005 (N_20005,N_19779,N_19487);
nand U20006 (N_20006,N_19590,N_19425);
and U20007 (N_20007,N_19313,N_19551);
and U20008 (N_20008,N_19079,N_19801);
or U20009 (N_20009,N_19175,N_19050);
or U20010 (N_20010,N_19228,N_19909);
nand U20011 (N_20011,N_19334,N_19545);
nor U20012 (N_20012,N_19264,N_19508);
or U20013 (N_20013,N_19843,N_18797);
or U20014 (N_20014,N_19100,N_19147);
xnor U20015 (N_20015,N_19058,N_19210);
xor U20016 (N_20016,N_18843,N_19981);
nor U20017 (N_20017,N_19149,N_19066);
nand U20018 (N_20018,N_19835,N_19054);
and U20019 (N_20019,N_19823,N_19641);
xnor U20020 (N_20020,N_19656,N_18760);
or U20021 (N_20021,N_19467,N_18801);
xor U20022 (N_20022,N_19134,N_18834);
nand U20023 (N_20023,N_18967,N_19599);
nor U20024 (N_20024,N_19416,N_19192);
xor U20025 (N_20025,N_19906,N_19400);
xor U20026 (N_20026,N_18921,N_19824);
and U20027 (N_20027,N_19026,N_18966);
and U20028 (N_20028,N_19056,N_19456);
nand U20029 (N_20029,N_19997,N_18751);
nor U20030 (N_20030,N_19486,N_19349);
nand U20031 (N_20031,N_19095,N_19345);
or U20032 (N_20032,N_19238,N_19196);
nand U20033 (N_20033,N_19504,N_19584);
and U20034 (N_20034,N_18856,N_18934);
nand U20035 (N_20035,N_19772,N_19266);
nand U20036 (N_20036,N_19585,N_19690);
nand U20037 (N_20037,N_19493,N_19161);
and U20038 (N_20038,N_18877,N_18960);
nor U20039 (N_20039,N_19018,N_19621);
and U20040 (N_20040,N_19683,N_18917);
and U20041 (N_20041,N_18952,N_19742);
and U20042 (N_20042,N_19223,N_19326);
or U20043 (N_20043,N_19681,N_19327);
and U20044 (N_20044,N_19567,N_19650);
nor U20045 (N_20045,N_19502,N_18852);
xor U20046 (N_20046,N_19988,N_19432);
and U20047 (N_20047,N_19468,N_18903);
nor U20048 (N_20048,N_19787,N_18773);
and U20049 (N_20049,N_18823,N_19068);
nand U20050 (N_20050,N_19834,N_19112);
xor U20051 (N_20051,N_19254,N_19342);
and U20052 (N_20052,N_19568,N_18872);
nor U20053 (N_20053,N_19735,N_19029);
and U20054 (N_20054,N_19629,N_19007);
and U20055 (N_20055,N_19881,N_18962);
xnor U20056 (N_20056,N_19122,N_19308);
and U20057 (N_20057,N_19938,N_19440);
nor U20058 (N_20058,N_19057,N_19414);
nand U20059 (N_20059,N_19965,N_18763);
or U20060 (N_20060,N_19503,N_19732);
and U20061 (N_20061,N_18826,N_18774);
nor U20062 (N_20062,N_19789,N_19359);
nor U20063 (N_20063,N_19800,N_19478);
and U20064 (N_20064,N_19500,N_19218);
nand U20065 (N_20065,N_19514,N_19365);
nor U20066 (N_20066,N_19399,N_19880);
nor U20067 (N_20067,N_18887,N_19524);
nor U20068 (N_20068,N_19321,N_18997);
nand U20069 (N_20069,N_19290,N_19310);
xnor U20070 (N_20070,N_19461,N_19233);
xor U20071 (N_20071,N_19710,N_19804);
or U20072 (N_20072,N_19067,N_19372);
nand U20073 (N_20073,N_19806,N_19472);
nand U20074 (N_20074,N_19278,N_18758);
and U20075 (N_20075,N_18946,N_19113);
xor U20076 (N_20076,N_19548,N_19603);
xor U20077 (N_20077,N_19311,N_19395);
or U20078 (N_20078,N_19393,N_19918);
nor U20079 (N_20079,N_19251,N_19170);
and U20080 (N_20080,N_19247,N_18968);
nor U20081 (N_20081,N_18977,N_19505);
and U20082 (N_20082,N_19145,N_19755);
nand U20083 (N_20083,N_19573,N_19538);
and U20084 (N_20084,N_19968,N_19168);
nand U20085 (N_20085,N_19529,N_19929);
and U20086 (N_20086,N_18959,N_19914);
nor U20087 (N_20087,N_19867,N_19660);
and U20088 (N_20088,N_19604,N_19151);
nor U20089 (N_20089,N_18926,N_18750);
nand U20090 (N_20090,N_19385,N_18787);
and U20091 (N_20091,N_19544,N_19963);
nand U20092 (N_20092,N_19436,N_19108);
or U20093 (N_20093,N_19687,N_18838);
and U20094 (N_20094,N_19647,N_18886);
nor U20095 (N_20095,N_19291,N_19438);
and U20096 (N_20096,N_19088,N_19155);
nor U20097 (N_20097,N_19143,N_19745);
nor U20098 (N_20098,N_18756,N_19002);
or U20099 (N_20099,N_19759,N_18777);
xnor U20100 (N_20100,N_19454,N_19105);
nor U20101 (N_20101,N_19315,N_19542);
or U20102 (N_20102,N_19442,N_19336);
and U20103 (N_20103,N_19212,N_19350);
and U20104 (N_20104,N_19171,N_19827);
xor U20105 (N_20105,N_18931,N_19086);
xor U20106 (N_20106,N_19751,N_19571);
nand U20107 (N_20107,N_18900,N_19130);
or U20108 (N_20108,N_18815,N_19921);
or U20109 (N_20109,N_19976,N_19047);
or U20110 (N_20110,N_19966,N_19646);
nor U20111 (N_20111,N_19951,N_19878);
xnor U20112 (N_20112,N_19701,N_19672);
or U20113 (N_20113,N_19841,N_19733);
nor U20114 (N_20114,N_19126,N_19942);
nor U20115 (N_20115,N_18892,N_19236);
nand U20116 (N_20116,N_19366,N_19183);
nor U20117 (N_20117,N_18809,N_19932);
nand U20118 (N_20118,N_19260,N_19812);
nor U20119 (N_20119,N_19474,N_18840);
and U20120 (N_20120,N_18942,N_19839);
or U20121 (N_20121,N_19940,N_19977);
or U20122 (N_20122,N_19324,N_19106);
xor U20123 (N_20123,N_19415,N_19084);
or U20124 (N_20124,N_18998,N_19908);
xor U20125 (N_20125,N_19949,N_19999);
and U20126 (N_20126,N_18939,N_19319);
nor U20127 (N_20127,N_19314,N_19718);
and U20128 (N_20128,N_18907,N_19844);
nand U20129 (N_20129,N_19437,N_19148);
nand U20130 (N_20130,N_19727,N_19618);
and U20131 (N_20131,N_18824,N_18905);
nor U20132 (N_20132,N_19899,N_18794);
nor U20133 (N_20133,N_19541,N_19825);
xor U20134 (N_20134,N_18920,N_19182);
nor U20135 (N_20135,N_18890,N_19819);
nor U20136 (N_20136,N_19009,N_19035);
and U20137 (N_20137,N_19226,N_19782);
nand U20138 (N_20138,N_19281,N_19097);
nor U20139 (N_20139,N_19531,N_19747);
xnor U20140 (N_20140,N_18795,N_18891);
xnor U20141 (N_20141,N_19396,N_19587);
nor U20142 (N_20142,N_18902,N_19110);
nand U20143 (N_20143,N_19583,N_19131);
and U20144 (N_20144,N_19527,N_19022);
xor U20145 (N_20145,N_19103,N_19329);
or U20146 (N_20146,N_18893,N_19610);
xor U20147 (N_20147,N_19511,N_19144);
or U20148 (N_20148,N_19282,N_19377);
nor U20149 (N_20149,N_19870,N_19596);
nand U20150 (N_20150,N_19879,N_19159);
nor U20151 (N_20151,N_19215,N_18965);
and U20152 (N_20152,N_19957,N_19332);
or U20153 (N_20153,N_19992,N_19443);
nor U20154 (N_20154,N_19459,N_19591);
nor U20155 (N_20155,N_18901,N_19141);
nand U20156 (N_20156,N_19609,N_18844);
or U20157 (N_20157,N_19635,N_19617);
xor U20158 (N_20158,N_19348,N_19677);
nor U20159 (N_20159,N_19803,N_18833);
nand U20160 (N_20160,N_19030,N_19632);
and U20161 (N_20161,N_19275,N_19244);
nor U20162 (N_20162,N_19911,N_19252);
nor U20163 (N_20163,N_19640,N_19770);
or U20164 (N_20164,N_19555,N_19575);
and U20165 (N_20165,N_19337,N_18812);
nand U20166 (N_20166,N_19937,N_19785);
nor U20167 (N_20167,N_19749,N_19081);
and U20168 (N_20168,N_19605,N_19369);
nand U20169 (N_20169,N_19322,N_18954);
xnor U20170 (N_20170,N_19547,N_19513);
nand U20171 (N_20171,N_18767,N_19187);
nand U20172 (N_20172,N_19767,N_19743);
nor U20173 (N_20173,N_19179,N_19200);
and U20174 (N_20174,N_18867,N_19361);
nand U20175 (N_20175,N_19760,N_19905);
nor U20176 (N_20176,N_18781,N_19840);
nor U20177 (N_20177,N_18980,N_19012);
and U20178 (N_20178,N_19913,N_19875);
nand U20179 (N_20179,N_19962,N_19015);
xnor U20180 (N_20180,N_19490,N_19896);
nor U20181 (N_20181,N_19540,N_18854);
nand U20182 (N_20182,N_19277,N_19895);
xor U20183 (N_20183,N_19910,N_19116);
and U20184 (N_20184,N_18836,N_18964);
xor U20185 (N_20185,N_19598,N_18849);
and U20186 (N_20186,N_19792,N_19011);
and U20187 (N_20187,N_19089,N_18841);
and U20188 (N_20188,N_19008,N_18923);
xor U20189 (N_20189,N_19552,N_18799);
nor U20190 (N_20190,N_18858,N_19943);
or U20191 (N_20191,N_18853,N_19091);
or U20192 (N_20192,N_19661,N_19768);
nor U20193 (N_20193,N_19405,N_19495);
xor U20194 (N_20194,N_19070,N_19613);
or U20195 (N_20195,N_19697,N_18880);
and U20196 (N_20196,N_18904,N_19863);
nor U20197 (N_20197,N_19764,N_19814);
or U20198 (N_20198,N_19292,N_19219);
xnor U20199 (N_20199,N_19519,N_19273);
or U20200 (N_20200,N_19707,N_19802);
nor U20201 (N_20201,N_19649,N_19658);
xor U20202 (N_20202,N_19102,N_19889);
nand U20203 (N_20203,N_19499,N_19984);
nor U20204 (N_20204,N_18814,N_18888);
nor U20205 (N_20205,N_19430,N_19845);
nand U20206 (N_20206,N_18789,N_18911);
nand U20207 (N_20207,N_18828,N_19577);
nand U20208 (N_20208,N_18863,N_19027);
xor U20209 (N_20209,N_19589,N_18754);
nor U20210 (N_20210,N_19510,N_18783);
and U20211 (N_20211,N_19738,N_18974);
nand U20212 (N_20212,N_19719,N_19852);
or U20213 (N_20213,N_19832,N_19360);
nand U20214 (N_20214,N_18989,N_19331);
and U20215 (N_20215,N_18889,N_19995);
nand U20216 (N_20216,N_19586,N_19076);
nor U20217 (N_20217,N_19692,N_19229);
xor U20218 (N_20218,N_19522,N_19203);
nor U20219 (N_20219,N_19996,N_19856);
nand U20220 (N_20220,N_19428,N_19869);
nor U20221 (N_20221,N_19028,N_18915);
and U20222 (N_20222,N_19706,N_19362);
xor U20223 (N_20223,N_18969,N_19368);
nor U20224 (N_20224,N_19391,N_19959);
nor U20225 (N_20225,N_19257,N_19847);
xnor U20226 (N_20226,N_19158,N_19668);
nand U20227 (N_20227,N_19305,N_19739);
and U20228 (N_20228,N_19607,N_18805);
or U20229 (N_20229,N_18793,N_18818);
and U20230 (N_20230,N_19558,N_19915);
nor U20231 (N_20231,N_18827,N_18957);
and U20232 (N_20232,N_19872,N_19475);
nor U20233 (N_20233,N_19858,N_19588);
nor U20234 (N_20234,N_19859,N_18775);
xor U20235 (N_20235,N_19338,N_18786);
or U20236 (N_20236,N_19031,N_19927);
nand U20237 (N_20237,N_19973,N_19439);
xor U20238 (N_20238,N_19003,N_19922);
nand U20239 (N_20239,N_19411,N_19245);
xor U20240 (N_20240,N_19017,N_18855);
and U20241 (N_20241,N_19563,N_19163);
nor U20242 (N_20242,N_18932,N_19398);
and U20243 (N_20243,N_19280,N_19628);
or U20244 (N_20244,N_18940,N_19506);
nand U20245 (N_20245,N_19901,N_19044);
nand U20246 (N_20246,N_19713,N_19601);
xnor U20247 (N_20247,N_18829,N_19788);
or U20248 (N_20248,N_19941,N_19039);
or U20249 (N_20249,N_19670,N_19284);
nor U20250 (N_20250,N_18837,N_19036);
xor U20251 (N_20251,N_18983,N_19045);
and U20252 (N_20252,N_19128,N_19265);
nand U20253 (N_20253,N_19501,N_18779);
xnor U20254 (N_20254,N_18993,N_18961);
nand U20255 (N_20255,N_19268,N_19815);
xnor U20256 (N_20256,N_19295,N_19253);
or U20257 (N_20257,N_19700,N_18943);
xor U20258 (N_20258,N_19000,N_19831);
nand U20259 (N_20259,N_19286,N_19665);
and U20260 (N_20260,N_19484,N_19694);
xor U20261 (N_20261,N_18796,N_18807);
and U20262 (N_20262,N_19711,N_19794);
nor U20263 (N_20263,N_18896,N_19557);
nand U20264 (N_20264,N_19258,N_19928);
nor U20265 (N_20265,N_19691,N_19861);
or U20266 (N_20266,N_19673,N_19293);
nand U20267 (N_20267,N_19450,N_19185);
or U20268 (N_20268,N_19065,N_19761);
or U20269 (N_20269,N_19418,N_18876);
or U20270 (N_20270,N_19408,N_19139);
and U20271 (N_20271,N_19688,N_19205);
xnor U20272 (N_20272,N_19453,N_19777);
xnor U20273 (N_20273,N_18808,N_19682);
nor U20274 (N_20274,N_19190,N_19230);
or U20275 (N_20275,N_19897,N_19480);
nand U20276 (N_20276,N_19793,N_19926);
nand U20277 (N_20277,N_19309,N_19114);
nand U20278 (N_20278,N_19645,N_19902);
nor U20279 (N_20279,N_19256,N_19828);
and U20280 (N_20280,N_19776,N_19964);
and U20281 (N_20281,N_19850,N_19750);
xnor U20282 (N_20282,N_19619,N_19730);
or U20283 (N_20283,N_18990,N_19887);
or U20284 (N_20284,N_19556,N_19952);
and U20285 (N_20285,N_19240,N_18925);
nor U20286 (N_20286,N_19644,N_18871);
xnor U20287 (N_20287,N_18816,N_19498);
xor U20288 (N_20288,N_19217,N_19463);
and U20289 (N_20289,N_19680,N_19207);
nor U20290 (N_20290,N_19572,N_19669);
xnor U20291 (N_20291,N_19894,N_19614);
and U20292 (N_20292,N_19521,N_19954);
or U20293 (N_20293,N_19945,N_19312);
and U20294 (N_20294,N_19580,N_19891);
or U20295 (N_20295,N_19675,N_19339);
nor U20296 (N_20296,N_18963,N_18924);
nand U20297 (N_20297,N_19156,N_19559);
or U20298 (N_20298,N_19986,N_19409);
nor U20299 (N_20299,N_19213,N_18879);
xor U20300 (N_20300,N_19160,N_19197);
or U20301 (N_20301,N_19307,N_19154);
xor U20302 (N_20302,N_19272,N_18970);
nand U20303 (N_20303,N_19837,N_19982);
nor U20304 (N_20304,N_19709,N_19092);
nor U20305 (N_20305,N_19569,N_19133);
xnor U20306 (N_20306,N_19374,N_19127);
and U20307 (N_20307,N_19447,N_19402);
and U20308 (N_20308,N_19714,N_19662);
nand U20309 (N_20309,N_19367,N_19109);
xnor U20310 (N_20310,N_19765,N_19758);
and U20311 (N_20311,N_18755,N_19032);
nor U20312 (N_20312,N_18938,N_18782);
xnor U20313 (N_20313,N_19882,N_19564);
or U20314 (N_20314,N_19497,N_18912);
nor U20315 (N_20315,N_19830,N_19351);
nand U20316 (N_20316,N_19390,N_19021);
nor U20317 (N_20317,N_19167,N_18778);
or U20318 (N_20318,N_19346,N_19255);
or U20319 (N_20319,N_19449,N_19451);
xor U20320 (N_20320,N_19539,N_18865);
nor U20321 (N_20321,N_19052,N_19080);
nor U20322 (N_20322,N_19378,N_19703);
and U20323 (N_20323,N_19686,N_18895);
or U20324 (N_20324,N_19594,N_18869);
xor U20325 (N_20325,N_19972,N_18922);
nand U20326 (N_20326,N_19693,N_19485);
or U20327 (N_20327,N_19446,N_18761);
and U20328 (N_20328,N_19237,N_19098);
nor U20329 (N_20329,N_19898,N_19199);
nand U20330 (N_20330,N_19403,N_19471);
xor U20331 (N_20331,N_18948,N_18979);
nor U20332 (N_20332,N_19093,N_19698);
xor U20333 (N_20333,N_19441,N_19034);
nor U20334 (N_20334,N_19689,N_19597);
or U20335 (N_20335,N_19358,N_19448);
nand U20336 (N_20336,N_19626,N_19162);
or U20337 (N_20337,N_19038,N_19379);
xnor U20338 (N_20338,N_19294,N_19797);
nand U20339 (N_20339,N_19987,N_19923);
xnor U20340 (N_20340,N_19234,N_19546);
or U20341 (N_20341,N_19534,N_19807);
nor U20342 (N_20342,N_18800,N_18884);
and U20343 (N_20343,N_19434,N_19469);
xnor U20344 (N_20344,N_19671,N_19757);
nor U20345 (N_20345,N_19364,N_19401);
nand U20346 (N_20346,N_19413,N_19612);
or U20347 (N_20347,N_19222,N_19970);
nand U20348 (N_20348,N_19094,N_19061);
xor U20349 (N_20349,N_19020,N_19176);
and U20350 (N_20350,N_19925,N_19317);
or U20351 (N_20351,N_19579,N_19829);
xor U20352 (N_20352,N_19298,N_19460);
xnor U20353 (N_20353,N_19933,N_18882);
xor U20354 (N_20354,N_19239,N_19198);
nand U20355 (N_20355,N_19010,N_19221);
xor U20356 (N_20356,N_19989,N_19301);
nand U20357 (N_20357,N_19994,N_18804);
and U20358 (N_20358,N_19716,N_19853);
and U20359 (N_20359,N_18784,N_19423);
and U20360 (N_20360,N_18770,N_19874);
nand U20361 (N_20361,N_19971,N_19132);
and U20362 (N_20362,N_19947,N_19518);
nand U20363 (N_20363,N_19530,N_19985);
nand U20364 (N_20364,N_19404,N_19983);
xnor U20365 (N_20365,N_18762,N_19115);
xnor U20366 (N_20366,N_19388,N_19948);
nor U20367 (N_20367,N_19784,N_19473);
nor U20368 (N_20368,N_19023,N_19944);
xor U20369 (N_20369,N_19269,N_19356);
or U20370 (N_20370,N_18936,N_19549);
and U20371 (N_20371,N_19136,N_18883);
nor U20372 (N_20372,N_18791,N_18862);
nor U20373 (N_20373,N_19796,N_19525);
or U20374 (N_20374,N_19259,N_18986);
and U20375 (N_20375,N_19912,N_19939);
or U20376 (N_20376,N_19462,N_18916);
and U20377 (N_20377,N_19826,N_19570);
nand U20378 (N_20378,N_19842,N_19328);
or U20379 (N_20379,N_19778,N_19191);
and U20380 (N_20380,N_19188,N_19846);
or U20381 (N_20381,N_18830,N_19775);
nand U20382 (N_20382,N_19025,N_19389);
nor U20383 (N_20383,N_19616,N_19195);
and U20384 (N_20384,N_19135,N_19330);
or U20385 (N_20385,N_19746,N_19553);
xor U20386 (N_20386,N_18820,N_19592);
xnor U20387 (N_20387,N_19381,N_19004);
nand U20388 (N_20388,N_19373,N_19235);
nand U20389 (N_20389,N_19465,N_19189);
nand U20390 (N_20390,N_19561,N_18988);
or U20391 (N_20391,N_19865,N_18947);
and U20392 (N_20392,N_19422,N_19520);
and U20393 (N_20393,N_19125,N_19476);
nand U20394 (N_20394,N_19166,N_18764);
nor U20395 (N_20395,N_18785,N_18835);
xor U20396 (N_20396,N_18825,N_19666);
xnor U20397 (N_20397,N_19809,N_19333);
nand U20398 (N_20398,N_18866,N_18832);
nand U20399 (N_20399,N_19752,N_19455);
and U20400 (N_20400,N_19704,N_19615);
and U20401 (N_20401,N_19276,N_19107);
nor U20402 (N_20402,N_19412,N_19435);
xor U20403 (N_20403,N_19833,N_18978);
xnor U20404 (N_20404,N_19608,N_18753);
and U20405 (N_20405,N_19157,N_18909);
xor U20406 (N_20406,N_19663,N_19496);
nand U20407 (N_20407,N_19383,N_19876);
nor U20408 (N_20408,N_19888,N_19457);
nor U20409 (N_20409,N_18992,N_19118);
nor U20410 (N_20410,N_19678,N_19602);
nand U20411 (N_20411,N_18982,N_18910);
nor U20412 (N_20412,N_19515,N_18999);
nand U20413 (N_20413,N_18996,N_19069);
or U20414 (N_20414,N_18848,N_19077);
or U20415 (N_20415,N_19458,N_19124);
nor U20416 (N_20416,N_18802,N_19655);
nand U20417 (N_20417,N_19781,N_19643);
nand U20418 (N_20418,N_19483,N_18870);
nand U20419 (N_20419,N_19274,N_19873);
xor U20420 (N_20420,N_19180,N_19444);
nor U20421 (N_20421,N_19920,N_19370);
xor U20422 (N_20422,N_19811,N_18851);
nand U20423 (N_20423,N_19153,N_19808);
and U20424 (N_20424,N_18845,N_18765);
xnor U20425 (N_20425,N_19737,N_18958);
nor U20426 (N_20426,N_19406,N_19231);
xor U20427 (N_20427,N_19325,N_19734);
nor U20428 (N_20428,N_18822,N_18766);
and U20429 (N_20429,N_19805,N_18987);
and U20430 (N_20430,N_19717,N_19990);
or U20431 (N_20431,N_19820,N_19090);
xnor U20432 (N_20432,N_19582,N_19172);
xor U20433 (N_20433,N_18780,N_19958);
nor U20434 (N_20434,N_18899,N_19304);
and U20435 (N_20435,N_18981,N_19699);
nand U20436 (N_20436,N_18850,N_19795);
or U20437 (N_20437,N_19287,N_19357);
nor U20438 (N_20438,N_19063,N_19464);
and U20439 (N_20439,N_19821,N_19554);
nor U20440 (N_20440,N_19303,N_19574);
and U20441 (N_20441,N_19715,N_19936);
nor U20442 (N_20442,N_19001,N_19517);
xnor U20443 (N_20443,N_19537,N_19043);
nor U20444 (N_20444,N_18821,N_19410);
or U20445 (N_20445,N_18984,N_19224);
and U20446 (N_20446,N_19283,N_19382);
or U20447 (N_20447,N_19363,N_19101);
or U20448 (N_20448,N_19684,N_19279);
and U20449 (N_20449,N_19648,N_19250);
or U20450 (N_20450,N_19013,N_19731);
nand U20451 (N_20451,N_19627,N_19774);
nor U20452 (N_20452,N_19523,N_18881);
or U20453 (N_20453,N_19762,N_19705);
or U20454 (N_20454,N_19866,N_19214);
and U20455 (N_20455,N_19978,N_19893);
nand U20456 (N_20456,N_19445,N_19376);
nand U20457 (N_20457,N_19073,N_18995);
or U20458 (N_20458,N_19193,N_18897);
and U20459 (N_20459,N_19169,N_18776);
nor U20460 (N_20460,N_19791,N_19974);
or U20461 (N_20461,N_19270,N_19320);
nand U20462 (N_20462,N_18906,N_19917);
xnor U20463 (N_20463,N_19786,N_19754);
nand U20464 (N_20464,N_19652,N_18792);
nand U20465 (N_20465,N_19062,N_18771);
and U20466 (N_20466,N_18941,N_18810);
xnor U20467 (N_20467,N_19960,N_19838);
xor U20468 (N_20468,N_19186,N_19593);
and U20469 (N_20469,N_18788,N_18951);
xor U20470 (N_20470,N_18864,N_18975);
nor U20471 (N_20471,N_19634,N_18976);
nand U20472 (N_20472,N_19046,N_19862);
nand U20473 (N_20473,N_19516,N_19729);
nand U20474 (N_20474,N_19299,N_19885);
nand U20475 (N_20475,N_19907,N_19536);
nor U20476 (N_20476,N_19216,N_19813);
nand U20477 (N_20477,N_19340,N_19854);
nor U20478 (N_20478,N_19857,N_19685);
nand U20479 (N_20479,N_19877,N_19816);
or U20480 (N_20480,N_19639,N_18868);
or U20481 (N_20481,N_19726,N_19433);
nand U20482 (N_20482,N_19006,N_19930);
or U20483 (N_20483,N_18898,N_19969);
nand U20484 (N_20484,N_18955,N_19654);
nor U20485 (N_20485,N_19347,N_19071);
and U20486 (N_20486,N_19741,N_19723);
or U20487 (N_20487,N_18878,N_19622);
nand U20488 (N_20488,N_19740,N_19818);
and U20489 (N_20489,N_19600,N_18973);
nand U20490 (N_20490,N_18806,N_19297);
and U20491 (N_20491,N_19883,N_19146);
nand U20492 (N_20492,N_19387,N_19051);
nand U20493 (N_20493,N_19241,N_19904);
nand U20494 (N_20494,N_19955,N_19783);
nand U20495 (N_20495,N_19227,N_19288);
nand U20496 (N_20496,N_19263,N_19085);
xor U20497 (N_20497,N_19798,N_19397);
or U20498 (N_20498,N_19019,N_19353);
nand U20499 (N_20499,N_19033,N_19211);
and U20500 (N_20500,N_19016,N_19676);
xnor U20501 (N_20501,N_19679,N_19481);
nor U20502 (N_20502,N_19728,N_19494);
nor U20503 (N_20503,N_19780,N_19037);
nand U20504 (N_20504,N_19562,N_19104);
or U20505 (N_20505,N_19202,N_19392);
xnor U20506 (N_20506,N_19137,N_19142);
xor U20507 (N_20507,N_18908,N_19753);
or U20508 (N_20508,N_19452,N_19919);
or U20509 (N_20509,N_19871,N_18953);
and U20510 (N_20510,N_19611,N_19625);
xnor U20511 (N_20511,N_19111,N_19053);
nand U20512 (N_20512,N_19296,N_19246);
nor U20513 (N_20513,N_19075,N_19005);
or U20514 (N_20514,N_19533,N_19072);
and U20515 (N_20515,N_18927,N_19578);
and U20516 (N_20516,N_19249,N_19316);
nor U20517 (N_20517,N_19024,N_19855);
xor U20518 (N_20518,N_18861,N_18873);
and U20519 (N_20519,N_19177,N_19201);
nand U20520 (N_20520,N_19078,N_19232);
nand U20521 (N_20521,N_19535,N_19766);
nand U20522 (N_20522,N_19771,N_19119);
and U20523 (N_20523,N_19424,N_19956);
nand U20524 (N_20524,N_18914,N_19674);
xor U20525 (N_20525,N_18768,N_19890);
nand U20526 (N_20526,N_19431,N_19492);
xor U20527 (N_20527,N_19064,N_18935);
xor U20528 (N_20528,N_19712,N_19744);
and U20529 (N_20529,N_19248,N_19344);
or U20530 (N_20530,N_19642,N_18937);
and U20531 (N_20531,N_19375,N_19394);
nor U20532 (N_20532,N_19595,N_19993);
xor U20533 (N_20533,N_19961,N_18757);
nand U20534 (N_20534,N_18885,N_19306);
nor U20535 (N_20535,N_18933,N_19799);
nand U20536 (N_20536,N_19543,N_19208);
or U20537 (N_20537,N_19657,N_19836);
nand U20538 (N_20538,N_19708,N_19631);
xnor U20539 (N_20539,N_19623,N_19722);
and U20540 (N_20540,N_19242,N_19150);
or U20541 (N_20541,N_19323,N_19868);
nor U20542 (N_20542,N_19491,N_19289);
xnor U20543 (N_20543,N_19123,N_19164);
nand U20544 (N_20544,N_18894,N_19998);
nand U20545 (N_20545,N_19121,N_19756);
nand U20546 (N_20546,N_19178,N_19822);
nand U20547 (N_20547,N_19042,N_19924);
and U20548 (N_20548,N_19060,N_18913);
nor U20549 (N_20549,N_19509,N_19174);
or U20550 (N_20550,N_19206,N_19946);
nand U20551 (N_20551,N_19532,N_18819);
nor U20552 (N_20552,N_19470,N_19341);
nand U20553 (N_20553,N_19427,N_18971);
and U20554 (N_20554,N_19243,N_19931);
or U20555 (N_20555,N_19566,N_19851);
nor U20556 (N_20556,N_19041,N_19421);
and U20557 (N_20557,N_19773,N_19407);
nand U20558 (N_20558,N_19083,N_18972);
or U20559 (N_20559,N_19014,N_18991);
and U20560 (N_20560,N_18842,N_19271);
or U20561 (N_20561,N_18859,N_19049);
or U20562 (N_20562,N_18769,N_18860);
nand U20563 (N_20563,N_18847,N_19636);
nand U20564 (N_20564,N_19419,N_19953);
nor U20565 (N_20565,N_18945,N_19040);
and U20566 (N_20566,N_19129,N_19724);
xnor U20567 (N_20567,N_18929,N_19638);
and U20568 (N_20568,N_19386,N_18817);
and U20569 (N_20569,N_19725,N_19117);
xnor U20570 (N_20570,N_19225,N_19967);
nand U20571 (N_20571,N_19565,N_19417);
or U20572 (N_20572,N_18875,N_18839);
or U20573 (N_20573,N_19849,N_19702);
nand U20574 (N_20574,N_19120,N_18944);
nor U20575 (N_20575,N_18798,N_19181);
xnor U20576 (N_20576,N_19664,N_19526);
nand U20577 (N_20577,N_19384,N_18994);
xnor U20578 (N_20578,N_19576,N_19209);
or U20579 (N_20579,N_19560,N_19489);
or U20580 (N_20580,N_18918,N_18752);
xor U20581 (N_20581,N_19720,N_19352);
and U20582 (N_20582,N_18790,N_19900);
xor U20583 (N_20583,N_19935,N_19769);
xnor U20584 (N_20584,N_18772,N_19512);
or U20585 (N_20585,N_18803,N_19903);
nor U20586 (N_20586,N_19659,N_19354);
nand U20587 (N_20587,N_19864,N_19975);
nor U20588 (N_20588,N_19055,N_19721);
nand U20589 (N_20589,N_19138,N_19184);
or U20590 (N_20590,N_19048,N_19335);
or U20591 (N_20591,N_19482,N_18949);
and U20592 (N_20592,N_19488,N_19096);
and U20593 (N_20593,N_19884,N_19528);
xor U20594 (N_20594,N_19763,N_19507);
nand U20595 (N_20595,N_19420,N_19204);
and U20596 (N_20596,N_19991,N_19173);
nor U20597 (N_20597,N_18930,N_19620);
or U20598 (N_20598,N_19371,N_19074);
nand U20599 (N_20599,N_19633,N_19087);
nand U20600 (N_20600,N_19140,N_19980);
xnor U20601 (N_20601,N_19886,N_19637);
nor U20602 (N_20602,N_19696,N_19343);
xor U20603 (N_20603,N_18813,N_19285);
xor U20604 (N_20604,N_19099,N_18928);
and U20605 (N_20605,N_19653,N_18956);
and U20606 (N_20606,N_19477,N_18874);
xor U20607 (N_20607,N_19860,N_19606);
xnor U20608 (N_20608,N_19194,N_19667);
nand U20609 (N_20609,N_18831,N_18950);
and U20610 (N_20610,N_19892,N_19950);
nand U20611 (N_20611,N_19380,N_18857);
xnor U20612 (N_20612,N_19262,N_19624);
and U20613 (N_20613,N_19848,N_18759);
or U20614 (N_20614,N_19979,N_19810);
or U20615 (N_20615,N_18846,N_19355);
nand U20616 (N_20616,N_19302,N_19790);
or U20617 (N_20617,N_19651,N_19479);
or U20618 (N_20618,N_19550,N_18811);
and U20619 (N_20619,N_19426,N_19817);
nand U20620 (N_20620,N_19429,N_19300);
nor U20621 (N_20621,N_19220,N_19059);
or U20622 (N_20622,N_19695,N_19165);
and U20623 (N_20623,N_18985,N_19466);
or U20624 (N_20624,N_19581,N_19261);
nand U20625 (N_20625,N_19328,N_19903);
nor U20626 (N_20626,N_19906,N_19818);
xor U20627 (N_20627,N_19743,N_19138);
nand U20628 (N_20628,N_19631,N_19323);
nand U20629 (N_20629,N_19198,N_19234);
nand U20630 (N_20630,N_19494,N_19921);
xnor U20631 (N_20631,N_19204,N_18760);
xnor U20632 (N_20632,N_19918,N_18948);
nor U20633 (N_20633,N_19127,N_19243);
xor U20634 (N_20634,N_19454,N_19737);
and U20635 (N_20635,N_19641,N_19355);
nand U20636 (N_20636,N_18981,N_18925);
xnor U20637 (N_20637,N_19515,N_19706);
nor U20638 (N_20638,N_19248,N_19996);
nor U20639 (N_20639,N_19412,N_19141);
or U20640 (N_20640,N_19611,N_19420);
nor U20641 (N_20641,N_19958,N_19063);
xnor U20642 (N_20642,N_19996,N_19230);
or U20643 (N_20643,N_19407,N_19836);
xnor U20644 (N_20644,N_19867,N_19435);
nor U20645 (N_20645,N_19049,N_19142);
nor U20646 (N_20646,N_19986,N_19228);
nor U20647 (N_20647,N_19438,N_19105);
xor U20648 (N_20648,N_19895,N_19547);
xor U20649 (N_20649,N_19843,N_18894);
nor U20650 (N_20650,N_18983,N_19211);
xnor U20651 (N_20651,N_19813,N_19887);
xnor U20652 (N_20652,N_19045,N_19515);
nand U20653 (N_20653,N_19841,N_19987);
xor U20654 (N_20654,N_19871,N_19803);
nand U20655 (N_20655,N_18886,N_18961);
and U20656 (N_20656,N_18967,N_19449);
nor U20657 (N_20657,N_19383,N_19457);
nor U20658 (N_20658,N_19231,N_19653);
nor U20659 (N_20659,N_19194,N_19129);
nand U20660 (N_20660,N_19676,N_19566);
and U20661 (N_20661,N_19379,N_19334);
or U20662 (N_20662,N_19214,N_19130);
xor U20663 (N_20663,N_19444,N_19842);
xnor U20664 (N_20664,N_19495,N_19838);
nand U20665 (N_20665,N_19740,N_18815);
nand U20666 (N_20666,N_18853,N_19526);
or U20667 (N_20667,N_18904,N_19695);
xnor U20668 (N_20668,N_19041,N_18856);
xor U20669 (N_20669,N_19294,N_18849);
nand U20670 (N_20670,N_19159,N_19677);
and U20671 (N_20671,N_19902,N_19738);
nand U20672 (N_20672,N_19995,N_19751);
nor U20673 (N_20673,N_19047,N_19371);
nand U20674 (N_20674,N_18874,N_19204);
or U20675 (N_20675,N_19263,N_19172);
nor U20676 (N_20676,N_18921,N_19865);
or U20677 (N_20677,N_19349,N_19126);
xor U20678 (N_20678,N_19406,N_19713);
xor U20679 (N_20679,N_19820,N_19645);
nand U20680 (N_20680,N_19259,N_19847);
or U20681 (N_20681,N_18787,N_19757);
or U20682 (N_20682,N_19955,N_19349);
nand U20683 (N_20683,N_18754,N_19617);
xor U20684 (N_20684,N_19402,N_19064);
or U20685 (N_20685,N_19744,N_19819);
nand U20686 (N_20686,N_18833,N_19758);
nand U20687 (N_20687,N_18858,N_19093);
and U20688 (N_20688,N_19358,N_19932);
xor U20689 (N_20689,N_19073,N_19809);
nand U20690 (N_20690,N_19744,N_19284);
nor U20691 (N_20691,N_19372,N_18874);
nand U20692 (N_20692,N_19295,N_19026);
and U20693 (N_20693,N_18945,N_18899);
and U20694 (N_20694,N_19530,N_18759);
xnor U20695 (N_20695,N_19667,N_19401);
and U20696 (N_20696,N_19199,N_18934);
or U20697 (N_20697,N_19727,N_19222);
or U20698 (N_20698,N_19941,N_19785);
and U20699 (N_20699,N_18970,N_19652);
and U20700 (N_20700,N_19447,N_19454);
xnor U20701 (N_20701,N_19276,N_19393);
nand U20702 (N_20702,N_19135,N_19684);
nor U20703 (N_20703,N_19740,N_19195);
and U20704 (N_20704,N_19458,N_18849);
nor U20705 (N_20705,N_19874,N_19689);
and U20706 (N_20706,N_19583,N_19772);
xnor U20707 (N_20707,N_19756,N_18829);
nor U20708 (N_20708,N_19828,N_18842);
or U20709 (N_20709,N_19791,N_19340);
or U20710 (N_20710,N_19451,N_19883);
and U20711 (N_20711,N_18896,N_18999);
and U20712 (N_20712,N_19058,N_18782);
and U20713 (N_20713,N_19013,N_19021);
and U20714 (N_20714,N_19551,N_19814);
xnor U20715 (N_20715,N_19014,N_18894);
nand U20716 (N_20716,N_19149,N_19312);
or U20717 (N_20717,N_19152,N_18939);
and U20718 (N_20718,N_19724,N_18793);
nor U20719 (N_20719,N_18816,N_19277);
xnor U20720 (N_20720,N_19397,N_19071);
xor U20721 (N_20721,N_19608,N_18936);
or U20722 (N_20722,N_19459,N_19672);
nand U20723 (N_20723,N_19629,N_18877);
nand U20724 (N_20724,N_19468,N_19466);
nor U20725 (N_20725,N_19343,N_19136);
or U20726 (N_20726,N_19173,N_19771);
nor U20727 (N_20727,N_19322,N_19103);
or U20728 (N_20728,N_19589,N_19531);
nor U20729 (N_20729,N_19288,N_19780);
nor U20730 (N_20730,N_19202,N_18853);
and U20731 (N_20731,N_19632,N_19252);
and U20732 (N_20732,N_19165,N_19029);
nor U20733 (N_20733,N_19409,N_19896);
and U20734 (N_20734,N_18846,N_18792);
and U20735 (N_20735,N_18849,N_19188);
and U20736 (N_20736,N_18753,N_19677);
and U20737 (N_20737,N_19827,N_19291);
and U20738 (N_20738,N_19077,N_19045);
nand U20739 (N_20739,N_19381,N_19159);
xnor U20740 (N_20740,N_19382,N_18958);
and U20741 (N_20741,N_18828,N_19262);
or U20742 (N_20742,N_19289,N_19870);
nand U20743 (N_20743,N_19900,N_19166);
and U20744 (N_20744,N_19496,N_18918);
and U20745 (N_20745,N_19726,N_18788);
xor U20746 (N_20746,N_19585,N_19841);
nand U20747 (N_20747,N_19969,N_19609);
nand U20748 (N_20748,N_19294,N_19819);
or U20749 (N_20749,N_19211,N_19950);
or U20750 (N_20750,N_19996,N_19020);
nor U20751 (N_20751,N_18958,N_19666);
and U20752 (N_20752,N_19834,N_19685);
or U20753 (N_20753,N_19151,N_18906);
nor U20754 (N_20754,N_19896,N_18813);
nor U20755 (N_20755,N_19195,N_19461);
nand U20756 (N_20756,N_19009,N_18792);
nand U20757 (N_20757,N_19404,N_19916);
nor U20758 (N_20758,N_19592,N_19084);
or U20759 (N_20759,N_18809,N_19490);
or U20760 (N_20760,N_19180,N_19308);
nand U20761 (N_20761,N_19624,N_19852);
and U20762 (N_20762,N_19232,N_19611);
and U20763 (N_20763,N_19109,N_19383);
xnor U20764 (N_20764,N_19422,N_18831);
nand U20765 (N_20765,N_19000,N_19357);
xnor U20766 (N_20766,N_19141,N_19902);
or U20767 (N_20767,N_19616,N_19610);
or U20768 (N_20768,N_19725,N_19508);
and U20769 (N_20769,N_19996,N_19210);
or U20770 (N_20770,N_19287,N_19657);
or U20771 (N_20771,N_19322,N_19049);
or U20772 (N_20772,N_18867,N_19282);
xnor U20773 (N_20773,N_19851,N_19989);
xor U20774 (N_20774,N_19812,N_19993);
xnor U20775 (N_20775,N_19903,N_19605);
or U20776 (N_20776,N_19087,N_19842);
nand U20777 (N_20777,N_18762,N_19089);
xor U20778 (N_20778,N_19100,N_19569);
and U20779 (N_20779,N_19202,N_19927);
xor U20780 (N_20780,N_19895,N_19675);
or U20781 (N_20781,N_19089,N_19360);
and U20782 (N_20782,N_19441,N_18922);
nand U20783 (N_20783,N_19901,N_19262);
nand U20784 (N_20784,N_19085,N_19722);
nor U20785 (N_20785,N_18846,N_18789);
nor U20786 (N_20786,N_19984,N_19874);
and U20787 (N_20787,N_19041,N_19553);
and U20788 (N_20788,N_19215,N_18803);
nor U20789 (N_20789,N_18947,N_19488);
nor U20790 (N_20790,N_19772,N_19552);
nor U20791 (N_20791,N_19155,N_18777);
and U20792 (N_20792,N_19737,N_19762);
and U20793 (N_20793,N_19948,N_19846);
nor U20794 (N_20794,N_19624,N_19503);
nor U20795 (N_20795,N_19207,N_19745);
nor U20796 (N_20796,N_19064,N_19777);
or U20797 (N_20797,N_19715,N_19132);
nand U20798 (N_20798,N_19386,N_19982);
xnor U20799 (N_20799,N_19733,N_19695);
xor U20800 (N_20800,N_19614,N_19493);
xor U20801 (N_20801,N_19627,N_19525);
nor U20802 (N_20802,N_18807,N_19927);
nand U20803 (N_20803,N_19162,N_19502);
nor U20804 (N_20804,N_19147,N_18955);
or U20805 (N_20805,N_19383,N_19522);
xor U20806 (N_20806,N_19361,N_19023);
and U20807 (N_20807,N_18994,N_18853);
nand U20808 (N_20808,N_19156,N_18951);
nand U20809 (N_20809,N_19448,N_19144);
and U20810 (N_20810,N_19600,N_19453);
nor U20811 (N_20811,N_18766,N_19108);
or U20812 (N_20812,N_19112,N_19034);
nand U20813 (N_20813,N_19553,N_19779);
or U20814 (N_20814,N_19902,N_18766);
xor U20815 (N_20815,N_19302,N_19788);
nand U20816 (N_20816,N_18835,N_19545);
xnor U20817 (N_20817,N_19919,N_18843);
or U20818 (N_20818,N_19647,N_19343);
or U20819 (N_20819,N_19022,N_19257);
xor U20820 (N_20820,N_18753,N_19352);
nor U20821 (N_20821,N_19510,N_19927);
or U20822 (N_20822,N_19988,N_19909);
xor U20823 (N_20823,N_19893,N_19428);
nor U20824 (N_20824,N_19013,N_19100);
and U20825 (N_20825,N_19426,N_19868);
or U20826 (N_20826,N_19271,N_19192);
xor U20827 (N_20827,N_19518,N_19165);
or U20828 (N_20828,N_19880,N_19728);
nand U20829 (N_20829,N_19534,N_19458);
and U20830 (N_20830,N_18842,N_19170);
xnor U20831 (N_20831,N_18794,N_19773);
xnor U20832 (N_20832,N_19934,N_19955);
nand U20833 (N_20833,N_19392,N_19130);
or U20834 (N_20834,N_19701,N_19356);
nand U20835 (N_20835,N_19724,N_19299);
xnor U20836 (N_20836,N_18894,N_19284);
nor U20837 (N_20837,N_19563,N_19321);
xor U20838 (N_20838,N_19759,N_19449);
nor U20839 (N_20839,N_19846,N_18757);
or U20840 (N_20840,N_19324,N_19846);
or U20841 (N_20841,N_18795,N_19902);
xnor U20842 (N_20842,N_19899,N_19148);
and U20843 (N_20843,N_19484,N_19738);
nand U20844 (N_20844,N_19859,N_19345);
nor U20845 (N_20845,N_18887,N_19676);
or U20846 (N_20846,N_19133,N_19522);
xor U20847 (N_20847,N_18877,N_19432);
or U20848 (N_20848,N_19128,N_19137);
and U20849 (N_20849,N_19797,N_19655);
xor U20850 (N_20850,N_19375,N_19086);
nand U20851 (N_20851,N_18895,N_19349);
nor U20852 (N_20852,N_19461,N_19645);
nor U20853 (N_20853,N_19471,N_18891);
nor U20854 (N_20854,N_19392,N_19759);
nor U20855 (N_20855,N_19003,N_19034);
and U20856 (N_20856,N_19615,N_19409);
nand U20857 (N_20857,N_18768,N_19785);
nand U20858 (N_20858,N_18833,N_19150);
nand U20859 (N_20859,N_19731,N_19946);
nor U20860 (N_20860,N_19354,N_19431);
nand U20861 (N_20861,N_19795,N_19124);
nand U20862 (N_20862,N_19420,N_19168);
and U20863 (N_20863,N_19294,N_19699);
nor U20864 (N_20864,N_19954,N_19001);
and U20865 (N_20865,N_19338,N_19884);
and U20866 (N_20866,N_19131,N_19055);
nor U20867 (N_20867,N_18986,N_18789);
xnor U20868 (N_20868,N_19778,N_19805);
nor U20869 (N_20869,N_19967,N_19507);
nor U20870 (N_20870,N_18946,N_19094);
and U20871 (N_20871,N_19596,N_19960);
xor U20872 (N_20872,N_19256,N_19422);
and U20873 (N_20873,N_18955,N_19113);
or U20874 (N_20874,N_19092,N_18903);
and U20875 (N_20875,N_19194,N_19622);
or U20876 (N_20876,N_19588,N_18791);
or U20877 (N_20877,N_19511,N_19870);
or U20878 (N_20878,N_19044,N_19808);
nand U20879 (N_20879,N_19622,N_18917);
nor U20880 (N_20880,N_19944,N_19677);
xnor U20881 (N_20881,N_19091,N_19979);
and U20882 (N_20882,N_19916,N_19353);
or U20883 (N_20883,N_19129,N_19479);
or U20884 (N_20884,N_19502,N_19051);
nand U20885 (N_20885,N_18939,N_19993);
and U20886 (N_20886,N_19181,N_19408);
nor U20887 (N_20887,N_19216,N_18917);
and U20888 (N_20888,N_18982,N_19383);
nor U20889 (N_20889,N_19235,N_19360);
and U20890 (N_20890,N_19581,N_19241);
nor U20891 (N_20891,N_19164,N_18915);
nor U20892 (N_20892,N_18761,N_18824);
xnor U20893 (N_20893,N_19220,N_19399);
xnor U20894 (N_20894,N_18854,N_18840);
and U20895 (N_20895,N_19194,N_19539);
nand U20896 (N_20896,N_18824,N_18994);
or U20897 (N_20897,N_19586,N_19514);
or U20898 (N_20898,N_19082,N_18873);
nor U20899 (N_20899,N_19663,N_18864);
and U20900 (N_20900,N_18879,N_18825);
nor U20901 (N_20901,N_19362,N_19640);
or U20902 (N_20902,N_19694,N_19991);
nor U20903 (N_20903,N_19640,N_19254);
and U20904 (N_20904,N_19115,N_19095);
nor U20905 (N_20905,N_19220,N_19288);
or U20906 (N_20906,N_19011,N_18769);
nand U20907 (N_20907,N_19489,N_19535);
xnor U20908 (N_20908,N_18984,N_18991);
and U20909 (N_20909,N_19697,N_19056);
nor U20910 (N_20910,N_19903,N_19165);
nor U20911 (N_20911,N_19129,N_19873);
xor U20912 (N_20912,N_19149,N_19593);
xnor U20913 (N_20913,N_19486,N_19809);
nor U20914 (N_20914,N_19159,N_19358);
and U20915 (N_20915,N_19837,N_19035);
and U20916 (N_20916,N_19689,N_19450);
or U20917 (N_20917,N_18990,N_18848);
nand U20918 (N_20918,N_19254,N_19885);
xor U20919 (N_20919,N_19329,N_19858);
or U20920 (N_20920,N_18902,N_19835);
nor U20921 (N_20921,N_19534,N_19446);
xor U20922 (N_20922,N_19738,N_18964);
nor U20923 (N_20923,N_19971,N_19033);
xor U20924 (N_20924,N_19819,N_19238);
nor U20925 (N_20925,N_19115,N_19961);
and U20926 (N_20926,N_19193,N_19306);
or U20927 (N_20927,N_19236,N_18809);
nor U20928 (N_20928,N_19603,N_19943);
nor U20929 (N_20929,N_18917,N_19433);
xor U20930 (N_20930,N_19414,N_19423);
nor U20931 (N_20931,N_19958,N_18902);
nor U20932 (N_20932,N_19488,N_19440);
nand U20933 (N_20933,N_19074,N_19599);
xnor U20934 (N_20934,N_19064,N_18960);
nand U20935 (N_20935,N_19164,N_19947);
or U20936 (N_20936,N_19036,N_19372);
or U20937 (N_20937,N_19596,N_19874);
or U20938 (N_20938,N_18860,N_19399);
or U20939 (N_20939,N_19220,N_19099);
xnor U20940 (N_20940,N_19560,N_19417);
or U20941 (N_20941,N_18971,N_19015);
nand U20942 (N_20942,N_19420,N_18970);
nand U20943 (N_20943,N_18953,N_19458);
xnor U20944 (N_20944,N_19507,N_19625);
nand U20945 (N_20945,N_19991,N_19195);
nor U20946 (N_20946,N_19218,N_19185);
nor U20947 (N_20947,N_19313,N_19849);
and U20948 (N_20948,N_19672,N_19074);
xor U20949 (N_20949,N_19097,N_19647);
nor U20950 (N_20950,N_19868,N_19460);
and U20951 (N_20951,N_18851,N_19747);
nor U20952 (N_20952,N_19321,N_19340);
and U20953 (N_20953,N_19072,N_19911);
nor U20954 (N_20954,N_19537,N_19067);
xnor U20955 (N_20955,N_18769,N_19798);
and U20956 (N_20956,N_19692,N_19816);
nand U20957 (N_20957,N_19854,N_18880);
xor U20958 (N_20958,N_18833,N_19081);
or U20959 (N_20959,N_19100,N_19161);
and U20960 (N_20960,N_19499,N_19172);
or U20961 (N_20961,N_19446,N_19094);
and U20962 (N_20962,N_19821,N_19952);
nor U20963 (N_20963,N_19581,N_19082);
and U20964 (N_20964,N_19841,N_19017);
or U20965 (N_20965,N_19298,N_19138);
nor U20966 (N_20966,N_19453,N_19331);
and U20967 (N_20967,N_18767,N_19556);
nor U20968 (N_20968,N_19242,N_18900);
nor U20969 (N_20969,N_19491,N_18974);
and U20970 (N_20970,N_19362,N_19991);
nand U20971 (N_20971,N_19738,N_19048);
and U20972 (N_20972,N_18783,N_18913);
xnor U20973 (N_20973,N_19035,N_19005);
or U20974 (N_20974,N_19735,N_19574);
xor U20975 (N_20975,N_19382,N_19341);
xnor U20976 (N_20976,N_19701,N_19615);
nor U20977 (N_20977,N_19709,N_19044);
and U20978 (N_20978,N_19097,N_19026);
and U20979 (N_20979,N_19366,N_19867);
xor U20980 (N_20980,N_19860,N_18828);
nand U20981 (N_20981,N_19907,N_18973);
and U20982 (N_20982,N_19042,N_19320);
xnor U20983 (N_20983,N_19862,N_19446);
xnor U20984 (N_20984,N_19778,N_18789);
nand U20985 (N_20985,N_19819,N_18798);
nand U20986 (N_20986,N_19504,N_18916);
or U20987 (N_20987,N_19715,N_19280);
xor U20988 (N_20988,N_19044,N_18782);
or U20989 (N_20989,N_19116,N_19695);
or U20990 (N_20990,N_18931,N_19129);
nor U20991 (N_20991,N_18889,N_19944);
or U20992 (N_20992,N_18867,N_18758);
and U20993 (N_20993,N_19458,N_18876);
and U20994 (N_20994,N_18938,N_18914);
and U20995 (N_20995,N_19984,N_19426);
nor U20996 (N_20996,N_18769,N_18771);
nand U20997 (N_20997,N_19507,N_19519);
and U20998 (N_20998,N_18832,N_19456);
nand U20999 (N_20999,N_19022,N_19262);
nor U21000 (N_21000,N_19322,N_19935);
nor U21001 (N_21001,N_19219,N_18839);
nor U21002 (N_21002,N_19342,N_19242);
and U21003 (N_21003,N_18913,N_18948);
or U21004 (N_21004,N_19883,N_19372);
and U21005 (N_21005,N_19607,N_19187);
nor U21006 (N_21006,N_19114,N_19421);
or U21007 (N_21007,N_18924,N_19771);
xnor U21008 (N_21008,N_19753,N_19731);
and U21009 (N_21009,N_19453,N_18875);
and U21010 (N_21010,N_19424,N_19793);
nor U21011 (N_21011,N_19216,N_19058);
or U21012 (N_21012,N_19639,N_19380);
nor U21013 (N_21013,N_19602,N_19141);
nor U21014 (N_21014,N_19847,N_19537);
and U21015 (N_21015,N_19847,N_18965);
or U21016 (N_21016,N_19106,N_19520);
or U21017 (N_21017,N_19600,N_19227);
or U21018 (N_21018,N_19038,N_19971);
nor U21019 (N_21019,N_19826,N_19418);
xor U21020 (N_21020,N_19398,N_19265);
and U21021 (N_21021,N_19529,N_19662);
and U21022 (N_21022,N_19798,N_19844);
xnor U21023 (N_21023,N_19228,N_18776);
and U21024 (N_21024,N_19255,N_18768);
nor U21025 (N_21025,N_19176,N_19334);
nor U21026 (N_21026,N_19013,N_19687);
xor U21027 (N_21027,N_18948,N_19809);
or U21028 (N_21028,N_19621,N_19694);
and U21029 (N_21029,N_18958,N_18970);
or U21030 (N_21030,N_19602,N_19728);
or U21031 (N_21031,N_19508,N_19831);
or U21032 (N_21032,N_19398,N_19031);
and U21033 (N_21033,N_19120,N_19159);
nor U21034 (N_21034,N_19823,N_19260);
nand U21035 (N_21035,N_19846,N_18811);
xor U21036 (N_21036,N_19292,N_19636);
and U21037 (N_21037,N_19212,N_19169);
nand U21038 (N_21038,N_19522,N_19385);
nor U21039 (N_21039,N_19533,N_19385);
nor U21040 (N_21040,N_19409,N_19329);
nand U21041 (N_21041,N_19279,N_19443);
xor U21042 (N_21042,N_18946,N_19023);
nand U21043 (N_21043,N_19285,N_19974);
xnor U21044 (N_21044,N_18815,N_19665);
nor U21045 (N_21045,N_18931,N_19376);
and U21046 (N_21046,N_18775,N_19147);
and U21047 (N_21047,N_19456,N_19117);
nor U21048 (N_21048,N_19801,N_19327);
nand U21049 (N_21049,N_19322,N_19923);
and U21050 (N_21050,N_19937,N_19066);
and U21051 (N_21051,N_19567,N_19510);
nor U21052 (N_21052,N_19002,N_19185);
and U21053 (N_21053,N_19110,N_18838);
and U21054 (N_21054,N_19399,N_19367);
xor U21055 (N_21055,N_19268,N_18959);
nor U21056 (N_21056,N_19473,N_18964);
nor U21057 (N_21057,N_19422,N_19872);
and U21058 (N_21058,N_19250,N_19952);
or U21059 (N_21059,N_18793,N_19524);
nand U21060 (N_21060,N_19925,N_19239);
nand U21061 (N_21061,N_19271,N_19714);
or U21062 (N_21062,N_19519,N_19101);
and U21063 (N_21063,N_19677,N_19010);
xnor U21064 (N_21064,N_18899,N_19524);
xor U21065 (N_21065,N_18751,N_19285);
nand U21066 (N_21066,N_18816,N_18998);
or U21067 (N_21067,N_19574,N_19156);
and U21068 (N_21068,N_19850,N_19110);
nand U21069 (N_21069,N_19684,N_19751);
xnor U21070 (N_21070,N_18914,N_19586);
or U21071 (N_21071,N_19157,N_19656);
xor U21072 (N_21072,N_19468,N_19662);
nor U21073 (N_21073,N_19552,N_19176);
or U21074 (N_21074,N_19565,N_18952);
or U21075 (N_21075,N_19189,N_18896);
or U21076 (N_21076,N_19401,N_18876);
or U21077 (N_21077,N_19078,N_19158);
or U21078 (N_21078,N_19549,N_18935);
nand U21079 (N_21079,N_19577,N_18983);
and U21080 (N_21080,N_19525,N_18994);
or U21081 (N_21081,N_19980,N_19917);
nor U21082 (N_21082,N_19363,N_19674);
or U21083 (N_21083,N_18866,N_19178);
and U21084 (N_21084,N_19568,N_19338);
nor U21085 (N_21085,N_19364,N_19285);
nand U21086 (N_21086,N_19613,N_19114);
and U21087 (N_21087,N_19938,N_18974);
or U21088 (N_21088,N_19477,N_18918);
xnor U21089 (N_21089,N_19233,N_19632);
xor U21090 (N_21090,N_19072,N_19942);
xnor U21091 (N_21091,N_18839,N_19983);
nand U21092 (N_21092,N_19190,N_19267);
xnor U21093 (N_21093,N_19264,N_19207);
nand U21094 (N_21094,N_19481,N_19443);
nand U21095 (N_21095,N_19276,N_19980);
nor U21096 (N_21096,N_18765,N_18981);
nor U21097 (N_21097,N_19355,N_19025);
xnor U21098 (N_21098,N_18902,N_18954);
nand U21099 (N_21099,N_19714,N_18797);
and U21100 (N_21100,N_19800,N_18973);
and U21101 (N_21101,N_19228,N_19017);
nor U21102 (N_21102,N_19692,N_18972);
and U21103 (N_21103,N_19660,N_18829);
xnor U21104 (N_21104,N_18955,N_18893);
nor U21105 (N_21105,N_19670,N_19162);
and U21106 (N_21106,N_19578,N_19397);
or U21107 (N_21107,N_19884,N_19574);
xnor U21108 (N_21108,N_19204,N_19956);
xnor U21109 (N_21109,N_18803,N_19047);
and U21110 (N_21110,N_19757,N_19994);
xnor U21111 (N_21111,N_18971,N_19222);
or U21112 (N_21112,N_19013,N_19918);
nand U21113 (N_21113,N_19383,N_18762);
or U21114 (N_21114,N_19017,N_19667);
nor U21115 (N_21115,N_18986,N_18833);
nor U21116 (N_21116,N_19453,N_19764);
xnor U21117 (N_21117,N_19713,N_19888);
or U21118 (N_21118,N_18788,N_19163);
or U21119 (N_21119,N_19266,N_19793);
and U21120 (N_21120,N_19810,N_19716);
nor U21121 (N_21121,N_19925,N_19384);
or U21122 (N_21122,N_18957,N_19927);
nor U21123 (N_21123,N_19090,N_19608);
nand U21124 (N_21124,N_19810,N_19772);
nor U21125 (N_21125,N_19257,N_19374);
or U21126 (N_21126,N_19817,N_19464);
nor U21127 (N_21127,N_19015,N_18955);
nand U21128 (N_21128,N_19625,N_19571);
nand U21129 (N_21129,N_19570,N_19134);
nor U21130 (N_21130,N_19246,N_19349);
nand U21131 (N_21131,N_19076,N_18783);
or U21132 (N_21132,N_19766,N_19051);
xnor U21133 (N_21133,N_19693,N_18877);
nor U21134 (N_21134,N_19981,N_18962);
xor U21135 (N_21135,N_19463,N_19359);
or U21136 (N_21136,N_18795,N_19276);
nor U21137 (N_21137,N_19946,N_18888);
and U21138 (N_21138,N_19785,N_19442);
and U21139 (N_21139,N_19072,N_19227);
nand U21140 (N_21140,N_19607,N_19721);
nand U21141 (N_21141,N_19661,N_19963);
nor U21142 (N_21142,N_18932,N_19799);
or U21143 (N_21143,N_19888,N_19123);
xnor U21144 (N_21144,N_19263,N_19938);
and U21145 (N_21145,N_19725,N_18863);
nand U21146 (N_21146,N_19312,N_19942);
nor U21147 (N_21147,N_19710,N_19312);
and U21148 (N_21148,N_19414,N_19129);
nor U21149 (N_21149,N_19922,N_19352);
or U21150 (N_21150,N_19577,N_18774);
and U21151 (N_21151,N_19062,N_19494);
or U21152 (N_21152,N_19659,N_19151);
nor U21153 (N_21153,N_19092,N_18988);
nand U21154 (N_21154,N_19560,N_19492);
and U21155 (N_21155,N_19223,N_19405);
or U21156 (N_21156,N_19472,N_18840);
and U21157 (N_21157,N_19937,N_19143);
nand U21158 (N_21158,N_19706,N_19886);
and U21159 (N_21159,N_19877,N_19326);
and U21160 (N_21160,N_18939,N_19257);
nand U21161 (N_21161,N_19991,N_19568);
or U21162 (N_21162,N_19731,N_18972);
or U21163 (N_21163,N_19002,N_19877);
nand U21164 (N_21164,N_19033,N_19624);
nand U21165 (N_21165,N_18881,N_19345);
and U21166 (N_21166,N_19542,N_19333);
or U21167 (N_21167,N_19612,N_19273);
xor U21168 (N_21168,N_18974,N_19269);
or U21169 (N_21169,N_19626,N_19114);
or U21170 (N_21170,N_19538,N_19257);
and U21171 (N_21171,N_19806,N_19558);
nand U21172 (N_21172,N_19790,N_18989);
nor U21173 (N_21173,N_18952,N_19653);
xor U21174 (N_21174,N_18975,N_18845);
nand U21175 (N_21175,N_18876,N_19528);
and U21176 (N_21176,N_19172,N_18893);
and U21177 (N_21177,N_18766,N_19355);
nor U21178 (N_21178,N_19788,N_19495);
xnor U21179 (N_21179,N_18885,N_19272);
xor U21180 (N_21180,N_18847,N_19965);
and U21181 (N_21181,N_19784,N_19761);
or U21182 (N_21182,N_19047,N_19652);
and U21183 (N_21183,N_18954,N_19269);
nor U21184 (N_21184,N_19297,N_18814);
nor U21185 (N_21185,N_19179,N_19988);
or U21186 (N_21186,N_19582,N_19166);
nor U21187 (N_21187,N_19702,N_18973);
or U21188 (N_21188,N_19129,N_19989);
nor U21189 (N_21189,N_19984,N_19297);
nor U21190 (N_21190,N_18944,N_19340);
nand U21191 (N_21191,N_18959,N_19810);
or U21192 (N_21192,N_18913,N_19708);
nand U21193 (N_21193,N_19548,N_19061);
nand U21194 (N_21194,N_19881,N_19760);
and U21195 (N_21195,N_19341,N_19207);
xor U21196 (N_21196,N_19828,N_18997);
xnor U21197 (N_21197,N_19740,N_19561);
nand U21198 (N_21198,N_19813,N_19186);
xnor U21199 (N_21199,N_19854,N_19364);
or U21200 (N_21200,N_19434,N_19749);
nor U21201 (N_21201,N_18959,N_18770);
nand U21202 (N_21202,N_19735,N_18858);
xor U21203 (N_21203,N_18957,N_19836);
xor U21204 (N_21204,N_19603,N_19985);
or U21205 (N_21205,N_18781,N_19461);
nor U21206 (N_21206,N_19489,N_19435);
xor U21207 (N_21207,N_18786,N_19697);
xnor U21208 (N_21208,N_19694,N_19765);
or U21209 (N_21209,N_19917,N_19966);
nand U21210 (N_21210,N_19858,N_19601);
and U21211 (N_21211,N_19109,N_18906);
xnor U21212 (N_21212,N_19436,N_18772);
xor U21213 (N_21213,N_19567,N_19869);
nand U21214 (N_21214,N_19275,N_19159);
or U21215 (N_21215,N_19908,N_19082);
or U21216 (N_21216,N_19770,N_19447);
nor U21217 (N_21217,N_18988,N_19397);
nor U21218 (N_21218,N_18903,N_18750);
and U21219 (N_21219,N_18780,N_19771);
nand U21220 (N_21220,N_19899,N_18989);
xor U21221 (N_21221,N_19662,N_19696);
and U21222 (N_21222,N_19795,N_19257);
and U21223 (N_21223,N_19308,N_19280);
xnor U21224 (N_21224,N_19511,N_19084);
xor U21225 (N_21225,N_19845,N_19653);
or U21226 (N_21226,N_19334,N_18886);
or U21227 (N_21227,N_19481,N_19039);
nand U21228 (N_21228,N_19812,N_19378);
or U21229 (N_21229,N_18904,N_18798);
nand U21230 (N_21230,N_19235,N_19717);
nand U21231 (N_21231,N_18976,N_19359);
xor U21232 (N_21232,N_19594,N_18933);
xnor U21233 (N_21233,N_18765,N_19811);
or U21234 (N_21234,N_19747,N_19697);
nand U21235 (N_21235,N_19122,N_19377);
and U21236 (N_21236,N_18763,N_18885);
and U21237 (N_21237,N_19777,N_19602);
or U21238 (N_21238,N_19062,N_19694);
or U21239 (N_21239,N_18992,N_19763);
nor U21240 (N_21240,N_19990,N_18877);
or U21241 (N_21241,N_19064,N_19528);
nor U21242 (N_21242,N_19253,N_19852);
nor U21243 (N_21243,N_19947,N_19047);
nor U21244 (N_21244,N_19452,N_19362);
or U21245 (N_21245,N_19180,N_19111);
xor U21246 (N_21246,N_18833,N_19639);
xor U21247 (N_21247,N_19472,N_19840);
and U21248 (N_21248,N_18829,N_19581);
or U21249 (N_21249,N_18960,N_19315);
or U21250 (N_21250,N_21037,N_20457);
xnor U21251 (N_21251,N_20190,N_20366);
xnor U21252 (N_21252,N_20494,N_20128);
nand U21253 (N_21253,N_20837,N_20788);
or U21254 (N_21254,N_20519,N_20689);
or U21255 (N_21255,N_20380,N_21112);
nand U21256 (N_21256,N_20351,N_20402);
or U21257 (N_21257,N_20182,N_20969);
nand U21258 (N_21258,N_20866,N_20423);
nor U21259 (N_21259,N_20898,N_20473);
xnor U21260 (N_21260,N_20259,N_20195);
nor U21261 (N_21261,N_21132,N_20826);
and U21262 (N_21262,N_20000,N_20130);
or U21263 (N_21263,N_20513,N_20174);
nand U21264 (N_21264,N_21053,N_20159);
nand U21265 (N_21265,N_21044,N_20908);
and U21266 (N_21266,N_20528,N_20296);
nand U21267 (N_21267,N_20574,N_21061);
nand U21268 (N_21268,N_20461,N_21203);
or U21269 (N_21269,N_20620,N_21114);
xnor U21270 (N_21270,N_20045,N_20421);
or U21271 (N_21271,N_20120,N_20643);
nand U21272 (N_21272,N_20726,N_20716);
xor U21273 (N_21273,N_20083,N_20743);
xnor U21274 (N_21274,N_20966,N_20485);
nor U21275 (N_21275,N_20290,N_20853);
nand U21276 (N_21276,N_20993,N_21165);
xor U21277 (N_21277,N_20074,N_21167);
xnor U21278 (N_21278,N_20187,N_20142);
nor U21279 (N_21279,N_20915,N_21038);
nand U21280 (N_21280,N_20859,N_20081);
nor U21281 (N_21281,N_21057,N_20718);
and U21282 (N_21282,N_21238,N_20458);
nand U21283 (N_21283,N_20084,N_20923);
xnor U21284 (N_21284,N_20410,N_20735);
and U21285 (N_21285,N_20241,N_20870);
nand U21286 (N_21286,N_20659,N_20450);
nor U21287 (N_21287,N_21122,N_20036);
xnor U21288 (N_21288,N_20286,N_20227);
or U21289 (N_21289,N_20373,N_20326);
and U21290 (N_21290,N_20878,N_20525);
nor U21291 (N_21291,N_20035,N_20323);
nand U21292 (N_21292,N_20037,N_20847);
nand U21293 (N_21293,N_20792,N_21213);
xnor U21294 (N_21294,N_20972,N_20971);
nor U21295 (N_21295,N_20362,N_20379);
or U21296 (N_21296,N_20235,N_20670);
and U21297 (N_21297,N_20526,N_20765);
nand U21298 (N_21298,N_20695,N_20717);
or U21299 (N_21299,N_20684,N_21022);
nand U21300 (N_21300,N_21102,N_20575);
xor U21301 (N_21301,N_20066,N_21175);
nor U21302 (N_21302,N_20921,N_20938);
and U21303 (N_21303,N_20600,N_20427);
nor U21304 (N_21304,N_21050,N_20376);
nand U21305 (N_21305,N_20129,N_20904);
nor U21306 (N_21306,N_20989,N_20625);
and U21307 (N_21307,N_20677,N_20946);
xnor U21308 (N_21308,N_20137,N_20231);
and U21309 (N_21309,N_20442,N_21212);
xnor U21310 (N_21310,N_21239,N_20459);
and U21311 (N_21311,N_20869,N_21120);
and U21312 (N_21312,N_20002,N_20539);
nor U21313 (N_21313,N_20426,N_20723);
nor U21314 (N_21314,N_20367,N_20704);
nor U21315 (N_21315,N_20750,N_20642);
xnor U21316 (N_21316,N_21101,N_21187);
or U21317 (N_21317,N_20477,N_21123);
or U21318 (N_21318,N_20221,N_20185);
nand U21319 (N_21319,N_20798,N_20087);
and U21320 (N_21320,N_20167,N_20504);
xnor U21321 (N_21321,N_21182,N_20668);
nor U21322 (N_21322,N_20154,N_20073);
nand U21323 (N_21323,N_20919,N_20958);
nor U21324 (N_21324,N_20484,N_20731);
nand U21325 (N_21325,N_20926,N_20149);
nor U21326 (N_21326,N_20498,N_20455);
nor U21327 (N_21327,N_20722,N_20542);
nor U21328 (N_21328,N_20777,N_20452);
and U21329 (N_21329,N_20469,N_20424);
and U21330 (N_21330,N_20573,N_20780);
and U21331 (N_21331,N_20356,N_20360);
nor U21332 (N_21332,N_20611,N_20481);
or U21333 (N_21333,N_20829,N_20814);
nand U21334 (N_21334,N_21124,N_20057);
nand U21335 (N_21335,N_20827,N_20291);
nor U21336 (N_21336,N_20548,N_21012);
nor U21337 (N_21337,N_20489,N_20093);
nand U21338 (N_21338,N_21130,N_20747);
or U21339 (N_21339,N_20559,N_20601);
nand U21340 (N_21340,N_20646,N_20236);
and U21341 (N_21341,N_20618,N_20856);
xnor U21342 (N_21342,N_20739,N_20635);
nor U21343 (N_21343,N_20666,N_20407);
xor U21344 (N_21344,N_21091,N_20245);
and U21345 (N_21345,N_20994,N_20786);
nand U21346 (N_21346,N_20067,N_20558);
nor U21347 (N_21347,N_20209,N_20400);
xor U21348 (N_21348,N_20738,N_20740);
and U21349 (N_21349,N_21249,N_21228);
xor U21350 (N_21350,N_20163,N_20077);
and U21351 (N_21351,N_20508,N_20181);
xor U21352 (N_21352,N_20604,N_21148);
nand U21353 (N_21353,N_20085,N_20011);
and U21354 (N_21354,N_20721,N_21077);
nand U21355 (N_21355,N_20454,N_20346);
xor U21356 (N_21356,N_20627,N_21045);
and U21357 (N_21357,N_20664,N_20315);
or U21358 (N_21358,N_21002,N_20340);
and U21359 (N_21359,N_21161,N_21026);
xnor U21360 (N_21360,N_20456,N_20783);
nand U21361 (N_21361,N_20748,N_20629);
or U21362 (N_21362,N_20842,N_20590);
or U21363 (N_21363,N_20439,N_20701);
nand U21364 (N_21364,N_20110,N_20321);
nor U21365 (N_21365,N_21219,N_20314);
nand U21366 (N_21366,N_20692,N_20411);
nand U21367 (N_21367,N_20431,N_21007);
nand U21368 (N_21368,N_20238,N_20127);
xor U21369 (N_21369,N_20854,N_20417);
nor U21370 (N_21370,N_20720,N_21116);
or U21371 (N_21371,N_20425,N_20233);
and U21372 (N_21372,N_20913,N_20225);
nor U21373 (N_21373,N_21232,N_20358);
nand U21374 (N_21374,N_20339,N_20957);
and U21375 (N_21375,N_20515,N_21189);
nand U21376 (N_21376,N_20416,N_20215);
nor U21377 (N_21377,N_20433,N_20117);
nor U21378 (N_21378,N_21208,N_20509);
nand U21379 (N_21379,N_20025,N_21195);
and U21380 (N_21380,N_20125,N_21226);
or U21381 (N_21381,N_20071,N_20403);
nand U21382 (N_21382,N_21149,N_20636);
nor U21383 (N_21383,N_21031,N_21090);
nor U21384 (N_21384,N_20895,N_21020);
xor U21385 (N_21385,N_20864,N_21089);
nand U21386 (N_21386,N_20708,N_21158);
and U21387 (N_21387,N_21009,N_20429);
nor U21388 (N_21388,N_20696,N_21121);
or U21389 (N_21389,N_20602,N_20927);
or U21390 (N_21390,N_20404,N_21244);
or U21391 (N_21391,N_20732,N_20343);
or U21392 (N_21392,N_20947,N_20292);
nand U21393 (N_21393,N_20724,N_20341);
nor U21394 (N_21394,N_20186,N_20283);
xnor U21395 (N_21395,N_20211,N_20806);
and U21396 (N_21396,N_20309,N_20121);
nor U21397 (N_21397,N_21140,N_20164);
and U21398 (N_21398,N_20800,N_20293);
xor U21399 (N_21399,N_20942,N_20333);
or U21400 (N_21400,N_20703,N_21128);
nor U21401 (N_21401,N_20658,N_20986);
xor U21402 (N_21402,N_20147,N_21183);
or U21403 (N_21403,N_20448,N_20753);
nor U21404 (N_21404,N_20375,N_21198);
nor U21405 (N_21405,N_20387,N_20543);
or U21406 (N_21406,N_20445,N_20911);
or U21407 (N_21407,N_21115,N_20887);
xor U21408 (N_21408,N_20799,N_20131);
nor U21409 (N_21409,N_21117,N_20384);
nand U21410 (N_21410,N_21056,N_21001);
nor U21411 (N_21411,N_20550,N_21069);
or U21412 (N_21412,N_20116,N_20967);
and U21413 (N_21413,N_20157,N_21233);
xnor U21414 (N_21414,N_20428,N_20082);
nand U21415 (N_21415,N_21176,N_20063);
nand U21416 (N_21416,N_20446,N_20886);
or U21417 (N_21417,N_20940,N_20289);
nor U21418 (N_21418,N_21242,N_20569);
and U21419 (N_21419,N_20549,N_20165);
nand U21420 (N_21420,N_21047,N_20823);
xor U21421 (N_21421,N_20160,N_21042);
and U21422 (N_21422,N_20383,N_20839);
xnor U21423 (N_21423,N_20582,N_21019);
and U21424 (N_21424,N_20830,N_21025);
or U21425 (N_21425,N_20746,N_20390);
xnor U21426 (N_21426,N_20336,N_20766);
or U21427 (N_21427,N_20026,N_20273);
nor U21428 (N_21428,N_20307,N_20843);
nand U21429 (N_21429,N_20928,N_20662);
nand U21430 (N_21430,N_20172,N_20930);
xor U21431 (N_21431,N_20464,N_20626);
or U21432 (N_21432,N_20101,N_20902);
or U21433 (N_21433,N_20813,N_20909);
or U21434 (N_21434,N_20188,N_20420);
nor U21435 (N_21435,N_20937,N_20062);
and U21436 (N_21436,N_21154,N_20785);
nand U21437 (N_21437,N_20476,N_20821);
and U21438 (N_21438,N_20568,N_20492);
and U21439 (N_21439,N_20031,N_20903);
and U21440 (N_21440,N_20530,N_20020);
nand U21441 (N_21441,N_20941,N_20929);
or U21442 (N_21442,N_20516,N_20808);
xor U21443 (N_21443,N_20891,N_20672);
and U21444 (N_21444,N_20949,N_20311);
or U21445 (N_21445,N_20070,N_21191);
or U21446 (N_21446,N_21241,N_20086);
and U21447 (N_21447,N_20179,N_20220);
and U21448 (N_21448,N_21085,N_20441);
nand U21449 (N_21449,N_20222,N_21146);
xnor U21450 (N_21450,N_21129,N_20041);
nand U21451 (N_21451,N_20271,N_20505);
xnor U21452 (N_21452,N_20016,N_20624);
and U21453 (N_21453,N_20998,N_20547);
nand U21454 (N_21454,N_20284,N_20706);
nor U21455 (N_21455,N_20983,N_20579);
nand U21456 (N_21456,N_21086,N_20522);
nand U21457 (N_21457,N_20488,N_20261);
nor U21458 (N_21458,N_20155,N_20034);
xnor U21459 (N_21459,N_20007,N_20763);
and U21460 (N_21460,N_21168,N_20453);
nor U21461 (N_21461,N_20963,N_20742);
or U21462 (N_21462,N_20201,N_20419);
or U21463 (N_21463,N_20355,N_20955);
nor U21464 (N_21464,N_20363,N_20310);
xor U21465 (N_21465,N_20764,N_20653);
xnor U21466 (N_21466,N_21109,N_20345);
and U21467 (N_21467,N_20719,N_20254);
and U21468 (N_21468,N_20369,N_20888);
nand U21469 (N_21469,N_21014,N_20496);
nor U21470 (N_21470,N_21245,N_20462);
and U21471 (N_21471,N_20124,N_20274);
nor U21472 (N_21472,N_20216,N_20418);
nor U21473 (N_21473,N_21078,N_20534);
nor U21474 (N_21474,N_20444,N_20329);
or U21475 (N_21475,N_20920,N_20977);
xor U21476 (N_21476,N_20171,N_20503);
xor U21477 (N_21477,N_21214,N_20019);
or U21478 (N_21478,N_21147,N_21184);
nor U21479 (N_21479,N_21083,N_20050);
xor U21480 (N_21480,N_20180,N_21032);
and U21481 (N_21481,N_21151,N_21193);
nor U21482 (N_21482,N_20874,N_21105);
nor U21483 (N_21483,N_20838,N_21243);
nand U21484 (N_21484,N_20108,N_21013);
nor U21485 (N_21485,N_20266,N_20388);
nor U21486 (N_21486,N_20332,N_20776);
and U21487 (N_21487,N_21076,N_20578);
nand U21488 (N_21488,N_20751,N_20612);
or U21489 (N_21489,N_21048,N_20631);
or U21490 (N_21490,N_21204,N_20816);
nand U21491 (N_21491,N_20399,N_20507);
nand U21492 (N_21492,N_20916,N_20372);
or U21493 (N_21493,N_20665,N_20104);
xor U21494 (N_21494,N_20102,N_21153);
nor U21495 (N_21495,N_20594,N_20762);
nor U21496 (N_21496,N_20111,N_20487);
xnor U21497 (N_21497,N_20145,N_20634);
nor U21498 (N_21498,N_20858,N_20285);
xor U21499 (N_21499,N_20848,N_20828);
nor U21500 (N_21500,N_20393,N_20583);
and U21501 (N_21501,N_20774,N_21100);
nand U21502 (N_21502,N_20368,N_20178);
xor U21503 (N_21503,N_21231,N_20552);
nor U21504 (N_21504,N_20493,N_20268);
nor U21505 (N_21505,N_20595,N_20027);
nand U21506 (N_21506,N_20771,N_20514);
and U21507 (N_21507,N_20939,N_20688);
nor U21508 (N_21508,N_20619,N_20834);
or U21509 (N_21509,N_21136,N_21246);
nor U21510 (N_21510,N_20652,N_20694);
xnor U21511 (N_21511,N_21040,N_20194);
and U21512 (N_21512,N_20365,N_21202);
xor U21513 (N_21513,N_20354,N_21084);
nand U21514 (N_21514,N_20175,N_20756);
xnor U21515 (N_21515,N_21209,N_20080);
and U21516 (N_21516,N_20661,N_20510);
and U21517 (N_21517,N_21028,N_20820);
xor U21518 (N_21518,N_20076,N_20091);
and U21519 (N_21519,N_21099,N_20791);
nor U21520 (N_21520,N_20324,N_20557);
nor U21521 (N_21521,N_20890,N_20749);
nor U21522 (N_21522,N_20541,N_20924);
or U21523 (N_21523,N_20981,N_21177);
nor U21524 (N_21524,N_20072,N_21156);
or U21525 (N_21525,N_20055,N_20945);
xnor U21526 (N_21526,N_20674,N_21055);
xnor U21527 (N_21527,N_20278,N_20079);
xnor U21528 (N_21528,N_20951,N_20320);
and U21529 (N_21529,N_20303,N_20391);
nor U21530 (N_21530,N_20538,N_20934);
and U21531 (N_21531,N_21131,N_20412);
nand U21532 (N_21532,N_20685,N_20432);
and U21533 (N_21533,N_21006,N_20506);
nand U21534 (N_21534,N_20103,N_21186);
or U21535 (N_21535,N_20030,N_20841);
nor U21536 (N_21536,N_20678,N_20608);
nand U21537 (N_21537,N_20206,N_21034);
nor U21538 (N_21538,N_20435,N_20537);
xnor U21539 (N_21539,N_21024,N_20733);
xor U21540 (N_21540,N_20305,N_20012);
nor U21541 (N_21541,N_20871,N_20961);
xnor U21542 (N_21542,N_20168,N_20812);
nor U21543 (N_21543,N_20302,N_20217);
xor U21544 (N_21544,N_20191,N_20205);
nand U21545 (N_21545,N_20710,N_20013);
xnor U21546 (N_21546,N_20047,N_21110);
nand U21547 (N_21547,N_20563,N_20553);
and U21548 (N_21548,N_20023,N_21138);
or U21549 (N_21549,N_20396,N_20294);
xnor U21550 (N_21550,N_21072,N_20156);
nor U21551 (N_21551,N_20571,N_20647);
xnor U21552 (N_21552,N_20831,N_20861);
or U21553 (N_21553,N_20727,N_20654);
nor U21554 (N_21554,N_20879,N_20529);
nand U21555 (N_21555,N_20728,N_20546);
xnor U21556 (N_21556,N_21096,N_21097);
xnor U21557 (N_21557,N_20249,N_20803);
and U21558 (N_21558,N_20232,N_20682);
nor U21559 (N_21559,N_20767,N_20099);
nand U21560 (N_21560,N_20374,N_20385);
xor U21561 (N_21561,N_20158,N_20234);
or U21562 (N_21562,N_20198,N_20204);
xnor U21563 (N_21563,N_20781,N_20622);
nand U21564 (N_21564,N_21133,N_20141);
and U21565 (N_21565,N_20637,N_21200);
nor U21566 (N_21566,N_20985,N_20250);
nor U21567 (N_21567,N_20230,N_20299);
nand U21568 (N_21568,N_20975,N_20973);
nor U21569 (N_21569,N_20844,N_20581);
nor U21570 (N_21570,N_20730,N_20357);
nor U21571 (N_21571,N_20894,N_21143);
xnor U21572 (N_21572,N_20440,N_20381);
xor U21573 (N_21573,N_20202,N_20857);
or U21574 (N_21574,N_21169,N_20944);
or U21575 (N_21575,N_20655,N_20014);
xor U21576 (N_21576,N_20338,N_20851);
nor U21577 (N_21577,N_20593,N_20962);
nand U21578 (N_21578,N_21141,N_20483);
xor U21579 (N_21579,N_20935,N_20304);
nor U21580 (N_21580,N_20527,N_20901);
and U21581 (N_21581,N_20475,N_20449);
and U21582 (N_21582,N_20832,N_20010);
nand U21583 (N_21583,N_20193,N_20922);
or U21584 (N_21584,N_20460,N_20161);
xnor U21585 (N_21585,N_20032,N_20334);
and U21586 (N_21586,N_20673,N_20835);
nand U21587 (N_21587,N_20247,N_20545);
and U21588 (N_21588,N_20196,N_20219);
and U21589 (N_21589,N_20097,N_20337);
nand U21590 (N_21590,N_21188,N_20882);
and U21591 (N_21591,N_20576,N_20897);
or U21592 (N_21592,N_20257,N_20580);
or U21593 (N_21593,N_20645,N_21218);
xor U21594 (N_21594,N_20151,N_20018);
and U21595 (N_21595,N_20166,N_21205);
nand U21596 (N_21596,N_20094,N_20996);
nor U21597 (N_21597,N_20224,N_20997);
nor U21598 (N_21598,N_20822,N_21179);
and U21599 (N_21599,N_20702,N_20797);
nand U21600 (N_21600,N_20173,N_20144);
xor U21601 (N_21601,N_20825,N_20621);
xnor U21602 (N_21602,N_20386,N_20005);
and U21603 (N_21603,N_20714,N_20239);
or U21604 (N_21604,N_20042,N_20004);
nor U21605 (N_21605,N_20199,N_20352);
xnor U21606 (N_21606,N_21051,N_20775);
xor U21607 (N_21607,N_21126,N_20572);
nor U21608 (N_21608,N_21065,N_20984);
nand U21609 (N_21609,N_20115,N_20306);
and U21610 (N_21610,N_20451,N_20098);
nor U21611 (N_21611,N_20592,N_21067);
or U21612 (N_21612,N_20555,N_20422);
or U21613 (N_21613,N_20377,N_20933);
and U21614 (N_21614,N_21155,N_20787);
nand U21615 (N_21615,N_20148,N_20521);
and U21616 (N_21616,N_20881,N_20610);
nor U21617 (N_21617,N_20015,N_20263);
nor U21618 (N_21618,N_20139,N_21210);
xnor U21619 (N_21619,N_21075,N_20632);
nand U21620 (N_21620,N_20846,N_20650);
xnor U21621 (N_21621,N_20965,N_20855);
and U21622 (N_21622,N_20092,N_20395);
nor U21623 (N_21623,N_21058,N_21027);
or U21624 (N_21624,N_20840,N_20804);
nor U21625 (N_21625,N_21018,N_20599);
or U21626 (N_21626,N_20331,N_20480);
and U21627 (N_21627,N_20954,N_20090);
nand U21628 (N_21628,N_20176,N_20075);
nand U21629 (N_21629,N_20860,N_20133);
xnor U21630 (N_21630,N_20316,N_20512);
and U21631 (N_21631,N_21137,N_20565);
or U21632 (N_21632,N_20782,N_20370);
or U21633 (N_21633,N_21021,N_20544);
and U21634 (N_21634,N_20065,N_21224);
and U21635 (N_21635,N_21171,N_20039);
and U21636 (N_21636,N_20438,N_20761);
or U21637 (N_21637,N_21192,N_20226);
and U21638 (N_21638,N_20868,N_20189);
nand U21639 (N_21639,N_20577,N_21030);
or U21640 (N_21640,N_20607,N_21119);
and U21641 (N_21641,N_21197,N_21150);
nor U21642 (N_21642,N_20912,N_20415);
xnor U21643 (N_21643,N_20006,N_20288);
and U21644 (N_21644,N_20656,N_20712);
and U21645 (N_21645,N_20676,N_21247);
or U21646 (N_21646,N_20524,N_21163);
nor U21647 (N_21647,N_20240,N_20298);
nor U21648 (N_21648,N_20135,N_20531);
or U21649 (N_21649,N_20889,N_21071);
nor U21650 (N_21650,N_20499,N_20212);
or U21651 (N_21651,N_20471,N_20342);
nand U21652 (N_21652,N_20143,N_20414);
nand U21653 (N_21653,N_20089,N_20591);
nand U21654 (N_21654,N_20648,N_20200);
xnor U21655 (N_21655,N_20279,N_20349);
nor U21656 (N_21656,N_20533,N_20687);
and U21657 (N_21657,N_20262,N_21070);
nor U21658 (N_21658,N_20693,N_21139);
nor U21659 (N_21659,N_20043,N_21217);
or U21660 (N_21660,N_20203,N_20392);
and U21661 (N_21661,N_20389,N_20849);
nand U21662 (N_21662,N_21073,N_20876);
xnor U21663 (N_21663,N_20606,N_21222);
and U21664 (N_21664,N_20008,N_20614);
or U21665 (N_21665,N_20361,N_20406);
xor U21666 (N_21666,N_20691,N_20109);
or U21667 (N_21667,N_20639,N_20896);
or U21668 (N_21668,N_20952,N_20197);
nand U21669 (N_21669,N_20709,N_21201);
xnor U21670 (N_21670,N_20999,N_20138);
and U21671 (N_21671,N_20443,N_21196);
nor U21672 (N_21672,N_20122,N_20312);
nand U21673 (N_21673,N_21081,N_20192);
or U21674 (N_21674,N_21068,N_20589);
and U21675 (N_21675,N_20409,N_20229);
nor U21676 (N_21676,N_20585,N_20146);
xnor U21677 (N_21677,N_20795,N_20644);
nor U21678 (N_21678,N_20651,N_20466);
nor U21679 (N_21679,N_21094,N_20478);
and U21680 (N_21680,N_21010,N_20815);
nor U21681 (N_21681,N_20501,N_21064);
xor U21682 (N_21682,N_20755,N_20244);
xnor U21683 (N_21683,N_20603,N_20246);
or U21684 (N_21684,N_20772,N_20056);
xor U21685 (N_21685,N_20001,N_20140);
or U21686 (N_21686,N_20183,N_21049);
nand U21687 (N_21687,N_20784,N_21060);
nor U21688 (N_21688,N_20623,N_20132);
nor U21689 (N_21689,N_21066,N_20276);
nand U21690 (N_21690,N_20567,N_20520);
nor U21691 (N_21691,N_21108,N_20096);
and U21692 (N_21692,N_21079,N_20350);
xor U21693 (N_21693,N_20605,N_21107);
or U21694 (N_21694,N_20914,N_20995);
or U21695 (N_21695,N_20883,N_20667);
and U21696 (N_21696,N_20300,N_20807);
and U21697 (N_21697,N_20327,N_20686);
xnor U21698 (N_21698,N_20532,N_20769);
xor U21699 (N_21699,N_20382,N_20184);
or U21700 (N_21700,N_20207,N_21220);
and U21701 (N_21701,N_20932,N_21229);
or U21702 (N_21702,N_20170,N_20873);
nor U21703 (N_21703,N_21093,N_20152);
xor U21704 (N_21704,N_21215,N_20982);
and U21705 (N_21705,N_20757,N_20518);
or U21706 (N_21706,N_20744,N_21017);
and U21707 (N_21707,N_20264,N_20068);
and U21708 (N_21708,N_20628,N_21180);
and U21709 (N_21709,N_21103,N_20551);
nand U21710 (N_21710,N_20267,N_20463);
nand U21711 (N_21711,N_20009,N_20126);
nor U21712 (N_21712,N_20884,N_20925);
or U21713 (N_21713,N_20313,N_20907);
nand U21714 (N_21714,N_20752,N_20401);
or U21715 (N_21715,N_21240,N_20208);
nand U21716 (N_21716,N_20741,N_20214);
xor U21717 (N_21717,N_21127,N_20308);
and U21718 (N_21718,N_20564,N_20474);
or U21719 (N_21719,N_21043,N_20675);
xor U21720 (N_21720,N_20046,N_20818);
xnor U21721 (N_21721,N_20758,N_21207);
and U21722 (N_21722,N_20408,N_20586);
nand U21723 (N_21723,N_20554,N_21036);
and U21724 (N_21724,N_20990,N_20638);
nand U21725 (N_21725,N_21113,N_20397);
xor U21726 (N_21726,N_20495,N_20280);
xnor U21727 (N_21727,N_20671,N_21145);
xor U21728 (N_21728,N_20681,N_20470);
nand U21729 (N_21729,N_20003,N_20123);
nor U21730 (N_21730,N_20255,N_20561);
nand U21731 (N_21731,N_20248,N_20237);
nand U21732 (N_21732,N_20778,N_20824);
or U21733 (N_21733,N_20811,N_20169);
nand U21734 (N_21734,N_21199,N_21023);
nand U21735 (N_21735,N_21074,N_21111);
or U21736 (N_21736,N_20613,N_21011);
or U21737 (N_21737,N_21172,N_20317);
nand U21738 (N_21738,N_21135,N_20892);
xor U21739 (N_21739,N_20479,N_20213);
nor U21740 (N_21740,N_20021,N_21004);
or U21741 (N_21741,N_21087,N_20497);
nand U21742 (N_21742,N_20865,N_21095);
or U21743 (N_21743,N_20413,N_20700);
nand U21744 (N_21744,N_20364,N_20760);
nand U21745 (N_21745,N_20281,N_21157);
xor U21746 (N_21746,N_20029,N_20258);
nor U21747 (N_21747,N_20863,N_21106);
nand U21748 (N_21748,N_21054,N_21118);
or U21749 (N_21749,N_20051,N_20095);
xnor U21750 (N_21750,N_20150,N_21166);
or U21751 (N_21751,N_20991,N_20679);
xor U21752 (N_21752,N_20344,N_20669);
and U21753 (N_21753,N_20069,N_20980);
nand U21754 (N_21754,N_20773,N_20598);
xnor U21755 (N_21755,N_21206,N_20918);
xor U21756 (N_21756,N_20588,N_21134);
nor U21757 (N_21757,N_20100,N_20950);
nand U21758 (N_21758,N_21173,N_20905);
nand U21759 (N_21759,N_21174,N_20270);
nor U21760 (N_21760,N_20136,N_21234);
or U21761 (N_21761,N_20953,N_20272);
nor U21762 (N_21762,N_20319,N_20347);
nand U21763 (N_21763,N_20680,N_20789);
and U21764 (N_21764,N_20570,N_20486);
nor U21765 (N_21765,N_20058,N_20833);
xor U21766 (N_21766,N_21178,N_20615);
nand U21767 (N_21767,N_20482,N_20113);
nand U21768 (N_21768,N_20875,N_20500);
or U21769 (N_21769,N_20322,N_20112);
xnor U21770 (N_21770,N_20943,N_20660);
and U21771 (N_21771,N_21000,N_20880);
xor U21772 (N_21772,N_21194,N_20437);
nor U21773 (N_21773,N_20088,N_20282);
nor U21774 (N_21774,N_20048,N_21170);
xor U21775 (N_21775,N_20044,N_21227);
nor U21776 (N_21776,N_20134,N_20275);
nor U21777 (N_21777,N_20251,N_20318);
nand U21778 (N_21778,N_20713,N_20022);
xnor U21779 (N_21779,N_20810,N_20745);
nor U21780 (N_21780,N_20640,N_20434);
nand U21781 (N_21781,N_20737,N_21211);
nor U21782 (N_21782,N_20430,N_20328);
nand U21783 (N_21783,N_20794,N_20223);
or U21784 (N_21784,N_21104,N_20867);
or U21785 (N_21785,N_21033,N_20301);
nor U21786 (N_21786,N_21144,N_20040);
or U21787 (N_21787,N_20394,N_20436);
xor U21788 (N_21788,N_20053,N_20033);
xnor U21789 (N_21789,N_20979,N_20597);
or U21790 (N_21790,N_20699,N_20260);
xor U21791 (N_21791,N_21159,N_20348);
or U21792 (N_21792,N_20243,N_21052);
nor U21793 (N_21793,N_20024,N_21005);
nor U21794 (N_21794,N_20729,N_20900);
and U21795 (N_21795,N_21088,N_21185);
nor U21796 (N_21796,N_20295,N_20378);
or U21797 (N_21797,N_20060,N_21162);
nor U21798 (N_21798,N_20405,N_20490);
nor U21799 (N_21799,N_20725,N_20609);
nor U21800 (N_21800,N_20802,N_20162);
nand U21801 (N_21801,N_21237,N_21016);
nand U21802 (N_21802,N_20218,N_20596);
nand U21803 (N_21803,N_20910,N_21062);
nand U21804 (N_21804,N_20988,N_21003);
xor U21805 (N_21805,N_21092,N_20917);
nand U21806 (N_21806,N_20540,N_20335);
nand U21807 (N_21807,N_20893,N_20956);
and U21808 (N_21808,N_20153,N_20970);
or U21809 (N_21809,N_20119,N_20277);
and U21810 (N_21810,N_20584,N_20059);
nand U21811 (N_21811,N_20960,N_21039);
nor U21812 (N_21812,N_20398,N_20936);
xor U21813 (N_21813,N_21152,N_21235);
and U21814 (N_21814,N_20465,N_21181);
xnor U21815 (N_21815,N_20562,N_20359);
nand U21816 (N_21816,N_20017,N_21223);
and U21817 (N_21817,N_20736,N_20177);
nand U21818 (N_21818,N_20697,N_20964);
or U21819 (N_21819,N_20523,N_20535);
nand U21820 (N_21820,N_20845,N_21164);
and U21821 (N_21821,N_20472,N_20228);
xor U21822 (N_21822,N_20630,N_21142);
and U21823 (N_21823,N_20560,N_20974);
nor U21824 (N_21824,N_20054,N_21190);
nor U21825 (N_21825,N_20491,N_21080);
or U21826 (N_21826,N_21035,N_20633);
or U21827 (N_21827,N_20850,N_20616);
xnor U21828 (N_21828,N_20566,N_20105);
nor U21829 (N_21829,N_20049,N_20253);
nor U21830 (N_21830,N_20325,N_21082);
nand U21831 (N_21831,N_20817,N_21221);
xnor U21832 (N_21832,N_20793,N_20759);
or U21833 (N_21833,N_20698,N_20061);
and U21834 (N_21834,N_20801,N_21059);
nand U21835 (N_21835,N_21015,N_20906);
nand U21836 (N_21836,N_20118,N_21225);
or U21837 (N_21837,N_20467,N_20705);
nand U21838 (N_21838,N_20617,N_20269);
nand U21839 (N_21839,N_20511,N_21041);
and U21840 (N_21840,N_20252,N_20978);
or U21841 (N_21841,N_20556,N_20028);
or U21842 (N_21842,N_20297,N_21160);
and U21843 (N_21843,N_21046,N_21236);
or U21844 (N_21844,N_20353,N_20447);
nand U21845 (N_21845,N_20715,N_20587);
nand U21846 (N_21846,N_20852,N_20256);
and U21847 (N_21847,N_20872,N_20330);
nor U21848 (N_21848,N_20779,N_20649);
and U21849 (N_21849,N_20819,N_20770);
or U21850 (N_21850,N_20711,N_20517);
xnor U21851 (N_21851,N_20078,N_21029);
or U21852 (N_21852,N_20987,N_20690);
nor U21853 (N_21853,N_20210,N_20641);
nor U21854 (N_21854,N_20948,N_20968);
xnor U21855 (N_21855,N_20862,N_20754);
nand U21856 (N_21856,N_21098,N_20790);
nor U21857 (N_21857,N_20992,N_20106);
and U21858 (N_21858,N_20707,N_20287);
or U21859 (N_21859,N_20734,N_20796);
xor U21860 (N_21860,N_20683,N_21230);
xor U21861 (N_21861,N_20663,N_20959);
xnor U21862 (N_21862,N_20836,N_20877);
nor U21863 (N_21863,N_20976,N_20899);
nor U21864 (N_21864,N_20885,N_21248);
or U21865 (N_21865,N_21125,N_21063);
nor U21866 (N_21866,N_20265,N_20536);
nand U21867 (N_21867,N_20768,N_20107);
and U21868 (N_21868,N_20064,N_21008);
or U21869 (N_21869,N_20114,N_20052);
or U21870 (N_21870,N_20805,N_20371);
and U21871 (N_21871,N_20502,N_20038);
xor U21872 (N_21872,N_20931,N_20809);
or U21873 (N_21873,N_21216,N_20657);
or U21874 (N_21874,N_20242,N_20468);
or U21875 (N_21875,N_20170,N_20113);
nand U21876 (N_21876,N_20034,N_20193);
nand U21877 (N_21877,N_20994,N_20388);
nor U21878 (N_21878,N_20907,N_20549);
or U21879 (N_21879,N_20191,N_20612);
nand U21880 (N_21880,N_20484,N_20620);
and U21881 (N_21881,N_20843,N_20338);
nor U21882 (N_21882,N_20654,N_20786);
xnor U21883 (N_21883,N_20079,N_21159);
xnor U21884 (N_21884,N_20081,N_20082);
and U21885 (N_21885,N_20613,N_21127);
xor U21886 (N_21886,N_20695,N_21040);
or U21887 (N_21887,N_20189,N_20732);
nor U21888 (N_21888,N_20787,N_20126);
nor U21889 (N_21889,N_20667,N_20203);
xnor U21890 (N_21890,N_20428,N_20583);
nor U21891 (N_21891,N_21090,N_20012);
or U21892 (N_21892,N_21087,N_20579);
nor U21893 (N_21893,N_21126,N_20589);
nor U21894 (N_21894,N_20753,N_20756);
nor U21895 (N_21895,N_20924,N_20574);
nand U21896 (N_21896,N_21036,N_20500);
and U21897 (N_21897,N_20718,N_20882);
nor U21898 (N_21898,N_20191,N_20436);
nor U21899 (N_21899,N_20201,N_20720);
or U21900 (N_21900,N_21118,N_20483);
nand U21901 (N_21901,N_21131,N_20764);
nor U21902 (N_21902,N_20475,N_20421);
xor U21903 (N_21903,N_21182,N_20290);
nor U21904 (N_21904,N_20786,N_20494);
or U21905 (N_21905,N_20103,N_21224);
nor U21906 (N_21906,N_20896,N_21150);
nor U21907 (N_21907,N_20181,N_20150);
nand U21908 (N_21908,N_20728,N_21203);
xor U21909 (N_21909,N_20204,N_20946);
and U21910 (N_21910,N_20045,N_21241);
and U21911 (N_21911,N_20044,N_21058);
xnor U21912 (N_21912,N_20608,N_20721);
nor U21913 (N_21913,N_21014,N_21168);
xnor U21914 (N_21914,N_20440,N_20783);
or U21915 (N_21915,N_20311,N_21073);
xnor U21916 (N_21916,N_20623,N_20530);
or U21917 (N_21917,N_20621,N_20509);
and U21918 (N_21918,N_20389,N_20994);
and U21919 (N_21919,N_21103,N_20628);
or U21920 (N_21920,N_20242,N_20552);
or U21921 (N_21921,N_20175,N_20635);
or U21922 (N_21922,N_20085,N_21024);
nor U21923 (N_21923,N_20184,N_20802);
and U21924 (N_21924,N_20996,N_20629);
and U21925 (N_21925,N_20373,N_20003);
or U21926 (N_21926,N_20809,N_20894);
and U21927 (N_21927,N_20857,N_20377);
nand U21928 (N_21928,N_20054,N_20008);
xnor U21929 (N_21929,N_20741,N_20394);
and U21930 (N_21930,N_21086,N_20373);
and U21931 (N_21931,N_20738,N_20311);
nand U21932 (N_21932,N_21200,N_21238);
or U21933 (N_21933,N_20101,N_20702);
or U21934 (N_21934,N_21245,N_21141);
xnor U21935 (N_21935,N_20785,N_20464);
or U21936 (N_21936,N_20743,N_20112);
and U21937 (N_21937,N_20369,N_20052);
nand U21938 (N_21938,N_20974,N_20562);
nand U21939 (N_21939,N_20362,N_20043);
nor U21940 (N_21940,N_20414,N_20811);
xnor U21941 (N_21941,N_20345,N_20862);
and U21942 (N_21942,N_21210,N_20315);
nand U21943 (N_21943,N_20162,N_20955);
nand U21944 (N_21944,N_20489,N_20088);
nand U21945 (N_21945,N_20939,N_21153);
xor U21946 (N_21946,N_20166,N_20590);
xnor U21947 (N_21947,N_21022,N_20515);
and U21948 (N_21948,N_20008,N_21183);
or U21949 (N_21949,N_20615,N_20764);
nor U21950 (N_21950,N_20887,N_21041);
nand U21951 (N_21951,N_21201,N_20356);
or U21952 (N_21952,N_20212,N_20824);
and U21953 (N_21953,N_20035,N_20674);
and U21954 (N_21954,N_20864,N_20987);
nor U21955 (N_21955,N_20323,N_21154);
and U21956 (N_21956,N_20682,N_20629);
nor U21957 (N_21957,N_20191,N_20744);
or U21958 (N_21958,N_21012,N_20749);
xnor U21959 (N_21959,N_20132,N_20604);
and U21960 (N_21960,N_20881,N_20792);
or U21961 (N_21961,N_20436,N_20928);
xor U21962 (N_21962,N_20093,N_20544);
nor U21963 (N_21963,N_20494,N_20773);
xor U21964 (N_21964,N_20524,N_20087);
nand U21965 (N_21965,N_20600,N_20987);
or U21966 (N_21966,N_20730,N_21191);
nand U21967 (N_21967,N_20833,N_20808);
or U21968 (N_21968,N_20585,N_20426);
xor U21969 (N_21969,N_20197,N_20105);
or U21970 (N_21970,N_20535,N_20266);
or U21971 (N_21971,N_20908,N_20369);
and U21972 (N_21972,N_20279,N_20070);
xor U21973 (N_21973,N_20933,N_20517);
or U21974 (N_21974,N_20236,N_20486);
and U21975 (N_21975,N_20431,N_21164);
and U21976 (N_21976,N_20477,N_20799);
nor U21977 (N_21977,N_20047,N_21054);
or U21978 (N_21978,N_21023,N_20378);
nand U21979 (N_21979,N_20625,N_20630);
nor U21980 (N_21980,N_20896,N_20563);
nor U21981 (N_21981,N_20619,N_20964);
or U21982 (N_21982,N_20808,N_20847);
nor U21983 (N_21983,N_20266,N_21093);
and U21984 (N_21984,N_20488,N_20620);
xor U21985 (N_21985,N_21058,N_21020);
and U21986 (N_21986,N_20452,N_20587);
nor U21987 (N_21987,N_20830,N_20411);
or U21988 (N_21988,N_20954,N_20049);
nand U21989 (N_21989,N_20204,N_20332);
nor U21990 (N_21990,N_20452,N_20931);
xnor U21991 (N_21991,N_20395,N_20060);
or U21992 (N_21992,N_20164,N_20313);
or U21993 (N_21993,N_21130,N_20706);
and U21994 (N_21994,N_21192,N_20070);
and U21995 (N_21995,N_20774,N_20533);
xor U21996 (N_21996,N_20903,N_20050);
nor U21997 (N_21997,N_20991,N_20651);
or U21998 (N_21998,N_20548,N_20280);
or U21999 (N_21999,N_20662,N_21203);
nand U22000 (N_22000,N_20323,N_21025);
nand U22001 (N_22001,N_21159,N_21084);
or U22002 (N_22002,N_20143,N_20865);
or U22003 (N_22003,N_21092,N_20345);
nand U22004 (N_22004,N_20612,N_20225);
xor U22005 (N_22005,N_20290,N_20384);
nand U22006 (N_22006,N_21046,N_20436);
or U22007 (N_22007,N_20897,N_20003);
and U22008 (N_22008,N_21161,N_20833);
and U22009 (N_22009,N_21207,N_20800);
nor U22010 (N_22010,N_20646,N_20258);
nand U22011 (N_22011,N_20669,N_20946);
or U22012 (N_22012,N_20396,N_20425);
nor U22013 (N_22013,N_21216,N_20002);
nor U22014 (N_22014,N_21043,N_20170);
nor U22015 (N_22015,N_20011,N_20368);
nand U22016 (N_22016,N_20897,N_20034);
and U22017 (N_22017,N_20117,N_20038);
nor U22018 (N_22018,N_20127,N_20299);
and U22019 (N_22019,N_20481,N_20927);
xnor U22020 (N_22020,N_21022,N_20760);
or U22021 (N_22021,N_20212,N_20006);
nand U22022 (N_22022,N_20251,N_21230);
nor U22023 (N_22023,N_20362,N_20805);
nor U22024 (N_22024,N_20420,N_20010);
nand U22025 (N_22025,N_20443,N_21094);
and U22026 (N_22026,N_20286,N_20244);
or U22027 (N_22027,N_20900,N_20393);
nor U22028 (N_22028,N_20849,N_20556);
and U22029 (N_22029,N_20759,N_20156);
and U22030 (N_22030,N_21149,N_20933);
and U22031 (N_22031,N_20156,N_20471);
nor U22032 (N_22032,N_20426,N_21081);
and U22033 (N_22033,N_20817,N_20866);
nor U22034 (N_22034,N_20773,N_20101);
nor U22035 (N_22035,N_20116,N_20275);
or U22036 (N_22036,N_20366,N_20167);
or U22037 (N_22037,N_20130,N_20863);
or U22038 (N_22038,N_20595,N_20129);
or U22039 (N_22039,N_20116,N_20292);
or U22040 (N_22040,N_20508,N_20452);
xnor U22041 (N_22041,N_20108,N_21207);
nand U22042 (N_22042,N_20826,N_20870);
nand U22043 (N_22043,N_20294,N_20054);
nand U22044 (N_22044,N_20091,N_20749);
and U22045 (N_22045,N_20643,N_20142);
nor U22046 (N_22046,N_20981,N_20873);
xnor U22047 (N_22047,N_20004,N_20508);
nor U22048 (N_22048,N_20441,N_21022);
or U22049 (N_22049,N_21238,N_20010);
and U22050 (N_22050,N_20968,N_21184);
xor U22051 (N_22051,N_20010,N_20118);
or U22052 (N_22052,N_20593,N_20681);
xnor U22053 (N_22053,N_21175,N_20290);
or U22054 (N_22054,N_20046,N_21043);
xnor U22055 (N_22055,N_20613,N_21145);
and U22056 (N_22056,N_21060,N_20828);
or U22057 (N_22057,N_20889,N_20159);
nand U22058 (N_22058,N_20655,N_20708);
nand U22059 (N_22059,N_21142,N_20176);
xor U22060 (N_22060,N_20088,N_21180);
or U22061 (N_22061,N_21126,N_20214);
nor U22062 (N_22062,N_20078,N_20483);
nor U22063 (N_22063,N_21008,N_20040);
xnor U22064 (N_22064,N_21236,N_20517);
or U22065 (N_22065,N_21158,N_20511);
and U22066 (N_22066,N_20196,N_20234);
nor U22067 (N_22067,N_20411,N_20581);
xnor U22068 (N_22068,N_20689,N_20768);
and U22069 (N_22069,N_20567,N_20145);
or U22070 (N_22070,N_20476,N_21142);
or U22071 (N_22071,N_20578,N_21193);
xor U22072 (N_22072,N_20270,N_20853);
nor U22073 (N_22073,N_20909,N_20693);
or U22074 (N_22074,N_21061,N_20380);
nor U22075 (N_22075,N_20142,N_20825);
or U22076 (N_22076,N_20673,N_20414);
or U22077 (N_22077,N_20178,N_20527);
nand U22078 (N_22078,N_20170,N_20127);
nand U22079 (N_22079,N_20207,N_20500);
or U22080 (N_22080,N_20455,N_20117);
and U22081 (N_22081,N_20625,N_20110);
xnor U22082 (N_22082,N_20423,N_20189);
nand U22083 (N_22083,N_20181,N_20488);
nand U22084 (N_22084,N_20258,N_20070);
or U22085 (N_22085,N_20459,N_20308);
or U22086 (N_22086,N_20324,N_21222);
nand U22087 (N_22087,N_21008,N_20820);
xor U22088 (N_22088,N_20534,N_20094);
or U22089 (N_22089,N_20535,N_20584);
xor U22090 (N_22090,N_20318,N_20765);
nor U22091 (N_22091,N_20737,N_20375);
nor U22092 (N_22092,N_20831,N_20092);
or U22093 (N_22093,N_21202,N_20538);
and U22094 (N_22094,N_20203,N_20985);
and U22095 (N_22095,N_20254,N_20579);
or U22096 (N_22096,N_20992,N_20434);
or U22097 (N_22097,N_21212,N_20203);
xnor U22098 (N_22098,N_21079,N_20975);
and U22099 (N_22099,N_20893,N_20583);
xor U22100 (N_22100,N_21181,N_20484);
xor U22101 (N_22101,N_20662,N_20503);
xnor U22102 (N_22102,N_21013,N_20419);
nor U22103 (N_22103,N_20087,N_20511);
and U22104 (N_22104,N_20606,N_20231);
or U22105 (N_22105,N_20840,N_20412);
xnor U22106 (N_22106,N_20546,N_20539);
nor U22107 (N_22107,N_20319,N_20086);
and U22108 (N_22108,N_20454,N_20149);
nand U22109 (N_22109,N_20880,N_20505);
nand U22110 (N_22110,N_20986,N_20305);
xnor U22111 (N_22111,N_20477,N_21230);
or U22112 (N_22112,N_20960,N_21102);
nor U22113 (N_22113,N_21055,N_21043);
nor U22114 (N_22114,N_20302,N_20660);
nand U22115 (N_22115,N_20349,N_21119);
nor U22116 (N_22116,N_21231,N_20621);
xnor U22117 (N_22117,N_20961,N_20280);
nor U22118 (N_22118,N_20713,N_20691);
nand U22119 (N_22119,N_20388,N_20356);
nand U22120 (N_22120,N_20884,N_21212);
and U22121 (N_22121,N_21036,N_20168);
nand U22122 (N_22122,N_20730,N_20559);
xnor U22123 (N_22123,N_20898,N_21006);
nor U22124 (N_22124,N_20941,N_20103);
nand U22125 (N_22125,N_21097,N_20614);
nor U22126 (N_22126,N_20452,N_21208);
nor U22127 (N_22127,N_20173,N_20268);
xnor U22128 (N_22128,N_21023,N_21106);
xnor U22129 (N_22129,N_20185,N_21039);
xnor U22130 (N_22130,N_21128,N_20995);
xor U22131 (N_22131,N_20189,N_21070);
or U22132 (N_22132,N_20083,N_20882);
xnor U22133 (N_22133,N_20330,N_20770);
xnor U22134 (N_22134,N_20468,N_20829);
nor U22135 (N_22135,N_20014,N_20571);
xnor U22136 (N_22136,N_20072,N_20544);
xnor U22137 (N_22137,N_20480,N_20824);
and U22138 (N_22138,N_20362,N_20831);
nor U22139 (N_22139,N_20627,N_20547);
and U22140 (N_22140,N_20945,N_20514);
xor U22141 (N_22141,N_20184,N_21178);
nand U22142 (N_22142,N_20201,N_20139);
and U22143 (N_22143,N_20078,N_20081);
and U22144 (N_22144,N_20198,N_20062);
and U22145 (N_22145,N_21204,N_21110);
nand U22146 (N_22146,N_20134,N_20801);
or U22147 (N_22147,N_20721,N_20210);
nand U22148 (N_22148,N_20397,N_20204);
or U22149 (N_22149,N_21185,N_20850);
nand U22150 (N_22150,N_20899,N_20113);
xor U22151 (N_22151,N_20706,N_20936);
and U22152 (N_22152,N_20263,N_20708);
and U22153 (N_22153,N_20512,N_21178);
and U22154 (N_22154,N_20904,N_20847);
and U22155 (N_22155,N_20326,N_20522);
nand U22156 (N_22156,N_21178,N_20549);
nor U22157 (N_22157,N_21229,N_20263);
or U22158 (N_22158,N_20066,N_21062);
xnor U22159 (N_22159,N_20067,N_20331);
xor U22160 (N_22160,N_21231,N_20932);
xor U22161 (N_22161,N_21023,N_20072);
and U22162 (N_22162,N_21194,N_20220);
xor U22163 (N_22163,N_20865,N_20234);
nor U22164 (N_22164,N_21020,N_20733);
or U22165 (N_22165,N_20066,N_21110);
xor U22166 (N_22166,N_21145,N_20137);
and U22167 (N_22167,N_20498,N_20973);
nor U22168 (N_22168,N_20991,N_20054);
xnor U22169 (N_22169,N_20641,N_20476);
xor U22170 (N_22170,N_20540,N_20967);
nand U22171 (N_22171,N_20128,N_21214);
or U22172 (N_22172,N_20869,N_20322);
or U22173 (N_22173,N_20732,N_20701);
and U22174 (N_22174,N_20180,N_20098);
and U22175 (N_22175,N_20171,N_21158);
and U22176 (N_22176,N_20080,N_20252);
nand U22177 (N_22177,N_20691,N_20637);
xnor U22178 (N_22178,N_20797,N_20506);
or U22179 (N_22179,N_21043,N_20002);
and U22180 (N_22180,N_20240,N_20917);
nor U22181 (N_22181,N_20528,N_21208);
nor U22182 (N_22182,N_20517,N_20341);
xnor U22183 (N_22183,N_20367,N_20412);
nand U22184 (N_22184,N_20577,N_20078);
nand U22185 (N_22185,N_20994,N_21157);
xnor U22186 (N_22186,N_21044,N_20004);
xor U22187 (N_22187,N_20252,N_20515);
and U22188 (N_22188,N_20581,N_20585);
nand U22189 (N_22189,N_20581,N_21196);
and U22190 (N_22190,N_20584,N_20743);
nand U22191 (N_22191,N_20518,N_20022);
nand U22192 (N_22192,N_20014,N_20920);
xnor U22193 (N_22193,N_20189,N_20878);
and U22194 (N_22194,N_20322,N_20141);
or U22195 (N_22195,N_20993,N_20134);
nor U22196 (N_22196,N_21177,N_20078);
xnor U22197 (N_22197,N_20131,N_20812);
xnor U22198 (N_22198,N_20672,N_20132);
or U22199 (N_22199,N_20310,N_20758);
xnor U22200 (N_22200,N_20883,N_21026);
and U22201 (N_22201,N_20438,N_20671);
and U22202 (N_22202,N_20178,N_20017);
and U22203 (N_22203,N_21111,N_21006);
xnor U22204 (N_22204,N_20616,N_20497);
xnor U22205 (N_22205,N_21107,N_20458);
and U22206 (N_22206,N_20352,N_20561);
nand U22207 (N_22207,N_20620,N_20509);
nand U22208 (N_22208,N_20297,N_20160);
nor U22209 (N_22209,N_20570,N_21110);
xor U22210 (N_22210,N_21183,N_20094);
nor U22211 (N_22211,N_20791,N_20719);
xnor U22212 (N_22212,N_20648,N_20987);
or U22213 (N_22213,N_21068,N_21188);
and U22214 (N_22214,N_20027,N_21067);
or U22215 (N_22215,N_21023,N_21236);
or U22216 (N_22216,N_20675,N_20671);
and U22217 (N_22217,N_20546,N_20435);
and U22218 (N_22218,N_20171,N_20966);
and U22219 (N_22219,N_20436,N_20258);
and U22220 (N_22220,N_20038,N_20614);
nand U22221 (N_22221,N_20798,N_20205);
nand U22222 (N_22222,N_21021,N_20815);
nand U22223 (N_22223,N_21081,N_20664);
xor U22224 (N_22224,N_20307,N_20373);
or U22225 (N_22225,N_20569,N_20389);
nor U22226 (N_22226,N_20231,N_21152);
or U22227 (N_22227,N_20929,N_20461);
xor U22228 (N_22228,N_21194,N_20943);
xnor U22229 (N_22229,N_21117,N_21238);
xnor U22230 (N_22230,N_20678,N_20762);
or U22231 (N_22231,N_20781,N_20181);
nor U22232 (N_22232,N_20912,N_20114);
and U22233 (N_22233,N_20656,N_20572);
nand U22234 (N_22234,N_20528,N_21083);
or U22235 (N_22235,N_20190,N_20895);
xor U22236 (N_22236,N_20147,N_20708);
and U22237 (N_22237,N_20512,N_21157);
xor U22238 (N_22238,N_21090,N_20951);
nand U22239 (N_22239,N_20580,N_20145);
or U22240 (N_22240,N_20016,N_21163);
or U22241 (N_22241,N_20218,N_20489);
nor U22242 (N_22242,N_20427,N_21050);
xnor U22243 (N_22243,N_20428,N_20788);
xor U22244 (N_22244,N_21125,N_20775);
nor U22245 (N_22245,N_20659,N_20013);
nor U22246 (N_22246,N_20264,N_20712);
nand U22247 (N_22247,N_20614,N_21236);
xor U22248 (N_22248,N_20974,N_20292);
xnor U22249 (N_22249,N_20435,N_20290);
or U22250 (N_22250,N_20407,N_20903);
or U22251 (N_22251,N_20326,N_20371);
nor U22252 (N_22252,N_20964,N_21185);
xor U22253 (N_22253,N_21135,N_20754);
xor U22254 (N_22254,N_20042,N_20706);
xor U22255 (N_22255,N_21141,N_20992);
nor U22256 (N_22256,N_20116,N_20591);
nand U22257 (N_22257,N_20643,N_20404);
or U22258 (N_22258,N_20424,N_20002);
xor U22259 (N_22259,N_20895,N_21052);
nand U22260 (N_22260,N_20052,N_20664);
xor U22261 (N_22261,N_20413,N_20538);
xor U22262 (N_22262,N_20168,N_20868);
nand U22263 (N_22263,N_20419,N_20199);
and U22264 (N_22264,N_20448,N_20757);
nor U22265 (N_22265,N_20535,N_20030);
or U22266 (N_22266,N_20963,N_21029);
or U22267 (N_22267,N_20163,N_20615);
and U22268 (N_22268,N_20705,N_21220);
or U22269 (N_22269,N_20184,N_20141);
or U22270 (N_22270,N_20896,N_20274);
or U22271 (N_22271,N_20823,N_20564);
nor U22272 (N_22272,N_20461,N_20137);
or U22273 (N_22273,N_20420,N_20918);
nor U22274 (N_22274,N_21169,N_20044);
and U22275 (N_22275,N_20875,N_20249);
nand U22276 (N_22276,N_20594,N_20931);
and U22277 (N_22277,N_20482,N_20693);
and U22278 (N_22278,N_21058,N_21131);
and U22279 (N_22279,N_20578,N_20642);
xor U22280 (N_22280,N_20780,N_20813);
nor U22281 (N_22281,N_20655,N_20394);
or U22282 (N_22282,N_20491,N_20589);
and U22283 (N_22283,N_20228,N_20716);
or U22284 (N_22284,N_20413,N_20189);
nand U22285 (N_22285,N_20855,N_20003);
or U22286 (N_22286,N_20460,N_20097);
nand U22287 (N_22287,N_21165,N_20898);
and U22288 (N_22288,N_20067,N_20894);
xnor U22289 (N_22289,N_20610,N_20974);
or U22290 (N_22290,N_20935,N_20290);
nand U22291 (N_22291,N_20163,N_20429);
nor U22292 (N_22292,N_20385,N_20665);
and U22293 (N_22293,N_20587,N_20641);
or U22294 (N_22294,N_20854,N_20478);
or U22295 (N_22295,N_20722,N_20713);
or U22296 (N_22296,N_21213,N_21223);
and U22297 (N_22297,N_20791,N_21029);
nand U22298 (N_22298,N_21061,N_20137);
nor U22299 (N_22299,N_20370,N_21215);
or U22300 (N_22300,N_20147,N_20617);
nor U22301 (N_22301,N_21126,N_20797);
xor U22302 (N_22302,N_20685,N_20917);
and U22303 (N_22303,N_20154,N_21180);
xnor U22304 (N_22304,N_20935,N_20403);
or U22305 (N_22305,N_21099,N_20674);
or U22306 (N_22306,N_20494,N_20308);
and U22307 (N_22307,N_20986,N_20091);
xnor U22308 (N_22308,N_20556,N_20975);
and U22309 (N_22309,N_20084,N_20946);
or U22310 (N_22310,N_20227,N_20540);
or U22311 (N_22311,N_20691,N_20678);
or U22312 (N_22312,N_20120,N_21124);
nand U22313 (N_22313,N_20551,N_20146);
nor U22314 (N_22314,N_20140,N_20828);
or U22315 (N_22315,N_20270,N_20088);
nand U22316 (N_22316,N_20965,N_21049);
or U22317 (N_22317,N_21232,N_20846);
or U22318 (N_22318,N_20217,N_20956);
or U22319 (N_22319,N_20112,N_21227);
nand U22320 (N_22320,N_21127,N_20489);
or U22321 (N_22321,N_20595,N_20540);
nand U22322 (N_22322,N_20465,N_20195);
or U22323 (N_22323,N_20054,N_20325);
nand U22324 (N_22324,N_20812,N_20251);
or U22325 (N_22325,N_20487,N_20032);
and U22326 (N_22326,N_20134,N_20863);
nor U22327 (N_22327,N_20687,N_20266);
nor U22328 (N_22328,N_20751,N_20194);
and U22329 (N_22329,N_20074,N_21247);
xnor U22330 (N_22330,N_21205,N_20674);
nand U22331 (N_22331,N_20298,N_21202);
xnor U22332 (N_22332,N_20785,N_21071);
xor U22333 (N_22333,N_20529,N_20375);
or U22334 (N_22334,N_20166,N_20079);
xnor U22335 (N_22335,N_20451,N_20138);
xor U22336 (N_22336,N_20253,N_20899);
nand U22337 (N_22337,N_20432,N_20561);
or U22338 (N_22338,N_20718,N_20119);
or U22339 (N_22339,N_20092,N_20253);
xnor U22340 (N_22340,N_20273,N_20638);
and U22341 (N_22341,N_20873,N_20349);
nand U22342 (N_22342,N_20173,N_20765);
and U22343 (N_22343,N_20034,N_20900);
nor U22344 (N_22344,N_20533,N_20892);
nand U22345 (N_22345,N_20911,N_21053);
xor U22346 (N_22346,N_20011,N_21055);
and U22347 (N_22347,N_20484,N_20290);
nand U22348 (N_22348,N_20549,N_20916);
and U22349 (N_22349,N_21116,N_21170);
nor U22350 (N_22350,N_20177,N_20935);
nand U22351 (N_22351,N_20889,N_20586);
xor U22352 (N_22352,N_20063,N_21044);
and U22353 (N_22353,N_20587,N_20322);
nand U22354 (N_22354,N_20755,N_20471);
or U22355 (N_22355,N_20730,N_21228);
and U22356 (N_22356,N_21135,N_20570);
or U22357 (N_22357,N_20310,N_20551);
xor U22358 (N_22358,N_20366,N_20487);
nand U22359 (N_22359,N_21067,N_21000);
nor U22360 (N_22360,N_20521,N_20540);
nor U22361 (N_22361,N_20932,N_20944);
and U22362 (N_22362,N_20849,N_20280);
or U22363 (N_22363,N_20573,N_21167);
xnor U22364 (N_22364,N_20780,N_20142);
nand U22365 (N_22365,N_21009,N_20281);
xnor U22366 (N_22366,N_21199,N_20621);
nand U22367 (N_22367,N_21086,N_20284);
xnor U22368 (N_22368,N_20557,N_20693);
xor U22369 (N_22369,N_20597,N_21191);
or U22370 (N_22370,N_21046,N_20109);
xor U22371 (N_22371,N_20672,N_20326);
nand U22372 (N_22372,N_20913,N_20515);
xor U22373 (N_22373,N_20170,N_20630);
xor U22374 (N_22374,N_20575,N_20155);
nor U22375 (N_22375,N_20390,N_20191);
nand U22376 (N_22376,N_20131,N_21053);
xor U22377 (N_22377,N_20964,N_20807);
and U22378 (N_22378,N_21150,N_20760);
nand U22379 (N_22379,N_21147,N_20967);
xnor U22380 (N_22380,N_20182,N_20795);
nor U22381 (N_22381,N_21139,N_20208);
and U22382 (N_22382,N_20747,N_20324);
or U22383 (N_22383,N_20688,N_20003);
and U22384 (N_22384,N_21009,N_20130);
or U22385 (N_22385,N_21237,N_20798);
nand U22386 (N_22386,N_20923,N_21000);
nor U22387 (N_22387,N_20243,N_20847);
or U22388 (N_22388,N_20290,N_20191);
or U22389 (N_22389,N_20707,N_20321);
and U22390 (N_22390,N_20177,N_20943);
nand U22391 (N_22391,N_20738,N_20986);
or U22392 (N_22392,N_20161,N_20400);
nor U22393 (N_22393,N_20074,N_21095);
nand U22394 (N_22394,N_21197,N_20460);
nand U22395 (N_22395,N_20489,N_21189);
xor U22396 (N_22396,N_20187,N_20844);
and U22397 (N_22397,N_20169,N_20390);
and U22398 (N_22398,N_20852,N_20760);
and U22399 (N_22399,N_20422,N_20539);
nand U22400 (N_22400,N_21123,N_21114);
xor U22401 (N_22401,N_20453,N_20185);
nor U22402 (N_22402,N_20258,N_20849);
xor U22403 (N_22403,N_21168,N_20953);
xnor U22404 (N_22404,N_20405,N_20253);
xnor U22405 (N_22405,N_20447,N_20076);
or U22406 (N_22406,N_20834,N_20640);
or U22407 (N_22407,N_20702,N_20774);
and U22408 (N_22408,N_20016,N_20293);
nand U22409 (N_22409,N_20046,N_21131);
nand U22410 (N_22410,N_20672,N_20620);
or U22411 (N_22411,N_20492,N_20490);
or U22412 (N_22412,N_20785,N_21086);
or U22413 (N_22413,N_20148,N_20036);
nor U22414 (N_22414,N_20325,N_20367);
nand U22415 (N_22415,N_20523,N_20237);
nor U22416 (N_22416,N_21177,N_20928);
nand U22417 (N_22417,N_20576,N_20062);
and U22418 (N_22418,N_21158,N_20777);
and U22419 (N_22419,N_20110,N_20449);
and U22420 (N_22420,N_21196,N_20945);
xor U22421 (N_22421,N_21019,N_20091);
nor U22422 (N_22422,N_20880,N_20688);
nand U22423 (N_22423,N_20595,N_21112);
or U22424 (N_22424,N_20933,N_20316);
xor U22425 (N_22425,N_20328,N_20281);
and U22426 (N_22426,N_21135,N_20505);
xor U22427 (N_22427,N_20167,N_20524);
or U22428 (N_22428,N_21077,N_20629);
or U22429 (N_22429,N_21150,N_20953);
and U22430 (N_22430,N_20351,N_21009);
nand U22431 (N_22431,N_20551,N_21115);
nor U22432 (N_22432,N_20441,N_20949);
or U22433 (N_22433,N_20670,N_20373);
nor U22434 (N_22434,N_20091,N_20295);
and U22435 (N_22435,N_20284,N_20954);
nor U22436 (N_22436,N_20423,N_20438);
and U22437 (N_22437,N_20460,N_20074);
nor U22438 (N_22438,N_20866,N_20595);
nor U22439 (N_22439,N_20116,N_20125);
or U22440 (N_22440,N_20117,N_20274);
xnor U22441 (N_22441,N_20419,N_20629);
or U22442 (N_22442,N_20135,N_20262);
xor U22443 (N_22443,N_20297,N_21238);
nand U22444 (N_22444,N_20332,N_20369);
nor U22445 (N_22445,N_20518,N_21197);
or U22446 (N_22446,N_20583,N_20124);
and U22447 (N_22447,N_21067,N_20237);
nand U22448 (N_22448,N_20769,N_20287);
nor U22449 (N_22449,N_20098,N_20968);
nand U22450 (N_22450,N_21194,N_20269);
nor U22451 (N_22451,N_20759,N_20444);
or U22452 (N_22452,N_20068,N_20120);
xor U22453 (N_22453,N_20915,N_20141);
and U22454 (N_22454,N_21169,N_20150);
xor U22455 (N_22455,N_20428,N_20353);
nor U22456 (N_22456,N_20563,N_20175);
nor U22457 (N_22457,N_20092,N_20991);
or U22458 (N_22458,N_21016,N_20706);
and U22459 (N_22459,N_21048,N_20051);
or U22460 (N_22460,N_21158,N_20218);
xor U22461 (N_22461,N_20739,N_20914);
xor U22462 (N_22462,N_21107,N_20669);
nand U22463 (N_22463,N_21123,N_21040);
nor U22464 (N_22464,N_20049,N_20347);
xor U22465 (N_22465,N_21042,N_20131);
and U22466 (N_22466,N_20104,N_21018);
nand U22467 (N_22467,N_20027,N_20183);
nor U22468 (N_22468,N_20091,N_20366);
and U22469 (N_22469,N_20974,N_20469);
and U22470 (N_22470,N_21141,N_21182);
xnor U22471 (N_22471,N_20161,N_20747);
and U22472 (N_22472,N_20368,N_20332);
xor U22473 (N_22473,N_21244,N_20225);
nor U22474 (N_22474,N_20698,N_20635);
nor U22475 (N_22475,N_20966,N_20336);
nand U22476 (N_22476,N_20206,N_20792);
xor U22477 (N_22477,N_20032,N_20062);
xnor U22478 (N_22478,N_20402,N_20577);
or U22479 (N_22479,N_20778,N_20423);
xor U22480 (N_22480,N_20921,N_21176);
xnor U22481 (N_22481,N_21068,N_20474);
or U22482 (N_22482,N_21033,N_21088);
xor U22483 (N_22483,N_20133,N_21004);
nand U22484 (N_22484,N_20014,N_21231);
or U22485 (N_22485,N_20203,N_20702);
nor U22486 (N_22486,N_20476,N_20607);
and U22487 (N_22487,N_20116,N_20433);
and U22488 (N_22488,N_21207,N_21006);
or U22489 (N_22489,N_20198,N_21081);
and U22490 (N_22490,N_20168,N_20094);
nor U22491 (N_22491,N_20160,N_20124);
xnor U22492 (N_22492,N_20823,N_20813);
xor U22493 (N_22493,N_21230,N_20438);
and U22494 (N_22494,N_20670,N_21158);
or U22495 (N_22495,N_20594,N_20567);
or U22496 (N_22496,N_20055,N_20283);
xor U22497 (N_22497,N_21140,N_20942);
nand U22498 (N_22498,N_20900,N_20101);
xor U22499 (N_22499,N_20715,N_21177);
nor U22500 (N_22500,N_22405,N_21281);
nor U22501 (N_22501,N_21641,N_22193);
nor U22502 (N_22502,N_21259,N_22179);
nor U22503 (N_22503,N_22186,N_21990);
nor U22504 (N_22504,N_22477,N_21595);
and U22505 (N_22505,N_21956,N_22252);
or U22506 (N_22506,N_21932,N_21526);
or U22507 (N_22507,N_21862,N_22402);
and U22508 (N_22508,N_22297,N_22492);
nor U22509 (N_22509,N_22011,N_22033);
xnor U22510 (N_22510,N_22429,N_22127);
or U22511 (N_22511,N_21663,N_21537);
or U22512 (N_22512,N_21940,N_22034);
or U22513 (N_22513,N_21412,N_21458);
nor U22514 (N_22514,N_21606,N_22028);
xnor U22515 (N_22515,N_22201,N_22263);
xor U22516 (N_22516,N_21823,N_22370);
or U22517 (N_22517,N_22436,N_22215);
or U22518 (N_22518,N_21450,N_22187);
and U22519 (N_22519,N_21425,N_21931);
xnor U22520 (N_22520,N_21430,N_21715);
xor U22521 (N_22521,N_22262,N_21445);
nand U22522 (N_22522,N_21778,N_21390);
or U22523 (N_22523,N_22257,N_21810);
xnor U22524 (N_22524,N_21948,N_21547);
nor U22525 (N_22525,N_21542,N_22237);
or U22526 (N_22526,N_21367,N_22414);
xor U22527 (N_22527,N_22242,N_22108);
xnor U22528 (N_22528,N_21876,N_21311);
nand U22529 (N_22529,N_21973,N_22393);
nor U22530 (N_22530,N_22132,N_21900);
or U22531 (N_22531,N_22185,N_21636);
xnor U22532 (N_22532,N_21275,N_22059);
or U22533 (N_22533,N_21438,N_21489);
or U22534 (N_22534,N_22497,N_21747);
nor U22535 (N_22535,N_21803,N_22403);
or U22536 (N_22536,N_22341,N_21677);
nand U22537 (N_22537,N_22366,N_22231);
nor U22538 (N_22538,N_22360,N_22418);
xor U22539 (N_22539,N_21396,N_21896);
xor U22540 (N_22540,N_21370,N_21361);
or U22541 (N_22541,N_21734,N_21714);
or U22542 (N_22542,N_22220,N_21303);
and U22543 (N_22543,N_22427,N_22382);
nor U22544 (N_22544,N_21617,N_22443);
and U22545 (N_22545,N_21284,N_22009);
xor U22546 (N_22546,N_21704,N_22157);
or U22547 (N_22547,N_21764,N_21433);
xor U22548 (N_22548,N_22441,N_21996);
nor U22549 (N_22549,N_22480,N_21944);
nor U22550 (N_22550,N_22364,N_21987);
or U22551 (N_22551,N_22378,N_22347);
nand U22552 (N_22552,N_22162,N_21437);
nor U22553 (N_22553,N_21988,N_21552);
and U22554 (N_22554,N_22498,N_22333);
or U22555 (N_22555,N_21880,N_22239);
xnor U22556 (N_22556,N_22408,N_21611);
xor U22557 (N_22557,N_21925,N_22250);
nor U22558 (N_22558,N_21665,N_22145);
and U22559 (N_22559,N_22043,N_22222);
xnor U22560 (N_22560,N_21680,N_22007);
or U22561 (N_22561,N_22103,N_22339);
xnor U22562 (N_22562,N_21411,N_21378);
and U22563 (N_22563,N_21258,N_21863);
or U22564 (N_22564,N_22189,N_21524);
nor U22565 (N_22565,N_21495,N_21858);
or U22566 (N_22566,N_21364,N_21564);
and U22567 (N_22567,N_21352,N_21793);
nand U22568 (N_22568,N_21723,N_21777);
nand U22569 (N_22569,N_22207,N_21942);
or U22570 (N_22570,N_21720,N_21969);
nand U22571 (N_22571,N_21737,N_21291);
nor U22572 (N_22572,N_21400,N_22042);
nor U22573 (N_22573,N_21502,N_22381);
or U22574 (N_22574,N_22357,N_21625);
xor U22575 (N_22575,N_22340,N_22013);
or U22576 (N_22576,N_21512,N_21365);
xnor U22577 (N_22577,N_21368,N_22183);
or U22578 (N_22578,N_21414,N_22149);
xnor U22579 (N_22579,N_21434,N_21510);
and U22580 (N_22580,N_22123,N_21846);
and U22581 (N_22581,N_22284,N_21519);
nand U22582 (N_22582,N_21724,N_22107);
and U22583 (N_22583,N_21757,N_21590);
nand U22584 (N_22584,N_21687,N_21253);
nand U22585 (N_22585,N_21428,N_21279);
nor U22586 (N_22586,N_22051,N_21933);
or U22587 (N_22587,N_21451,N_21923);
and U22588 (N_22588,N_22165,N_22040);
or U22589 (N_22589,N_22072,N_21692);
nand U22590 (N_22590,N_22411,N_22261);
nor U22591 (N_22591,N_21683,N_21917);
nand U22592 (N_22592,N_22368,N_21538);
nand U22593 (N_22593,N_22392,N_21706);
or U22594 (N_22594,N_21268,N_21946);
xnor U22595 (N_22595,N_22096,N_21276);
nor U22596 (N_22596,N_21310,N_22062);
nor U22597 (N_22597,N_21593,N_21600);
nor U22598 (N_22598,N_22109,N_22211);
xnor U22599 (N_22599,N_22318,N_21264);
nand U22600 (N_22600,N_22117,N_21882);
and U22601 (N_22601,N_22060,N_21662);
nor U22602 (N_22602,N_21958,N_21832);
or U22603 (N_22603,N_22337,N_22037);
and U22604 (N_22604,N_22012,N_21496);
or U22605 (N_22605,N_22039,N_22045);
and U22606 (N_22606,N_21758,N_21295);
or U22607 (N_22607,N_21885,N_21316);
xor U22608 (N_22608,N_22345,N_22273);
and U22609 (N_22609,N_21745,N_21561);
or U22610 (N_22610,N_21820,N_21350);
nor U22611 (N_22611,N_21760,N_22272);
nor U22612 (N_22612,N_22195,N_21460);
or U22613 (N_22613,N_22151,N_22468);
and U22614 (N_22614,N_21783,N_21825);
nand U22615 (N_22615,N_21672,N_21500);
nor U22616 (N_22616,N_21884,N_22387);
and U22617 (N_22617,N_21700,N_21667);
nor U22618 (N_22618,N_21659,N_21725);
nor U22619 (N_22619,N_21528,N_22097);
nor U22620 (N_22620,N_22088,N_21297);
nand U22621 (N_22621,N_21817,N_21573);
and U22622 (N_22622,N_21399,N_21380);
nor U22623 (N_22623,N_22140,N_22199);
and U22624 (N_22624,N_21815,N_22305);
nand U22625 (N_22625,N_22134,N_21601);
or U22626 (N_22626,N_21550,N_21572);
and U22627 (N_22627,N_22331,N_22432);
xnor U22628 (N_22628,N_21916,N_21325);
and U22629 (N_22629,N_22457,N_21827);
xnor U22630 (N_22630,N_22322,N_22154);
nand U22631 (N_22631,N_22113,N_21269);
and U22632 (N_22632,N_21807,N_21415);
xnor U22633 (N_22633,N_21675,N_21753);
xor U22634 (N_22634,N_21980,N_22421);
nand U22635 (N_22635,N_22281,N_22143);
xor U22636 (N_22636,N_22166,N_21616);
nor U22637 (N_22637,N_21462,N_21837);
or U22638 (N_22638,N_22463,N_22479);
or U22639 (N_22639,N_22248,N_22052);
nor U22640 (N_22640,N_21525,N_21466);
nor U22641 (N_22641,N_21849,N_21997);
nand U22642 (N_22642,N_22150,N_21355);
xnor U22643 (N_22643,N_21455,N_21543);
or U22644 (N_22644,N_21892,N_21494);
xor U22645 (N_22645,N_21392,N_21620);
or U22646 (N_22646,N_21304,N_21469);
nand U22647 (N_22647,N_21257,N_21541);
and U22648 (N_22648,N_22079,N_21794);
or U22649 (N_22649,N_21811,N_21331);
and U22650 (N_22650,N_21727,N_21599);
nand U22651 (N_22651,N_22080,N_21417);
and U22652 (N_22652,N_21787,N_21853);
xor U22653 (N_22653,N_22044,N_22424);
and U22654 (N_22654,N_21865,N_21797);
xor U22655 (N_22655,N_22235,N_21515);
or U22656 (N_22656,N_21372,N_22452);
nand U22657 (N_22657,N_21308,N_21947);
or U22658 (N_22658,N_21490,N_22131);
nand U22659 (N_22659,N_21324,N_22233);
or U22660 (N_22660,N_22081,N_22024);
nor U22661 (N_22661,N_21650,N_21909);
nor U22662 (N_22662,N_22067,N_21965);
and U22663 (N_22663,N_21901,N_22412);
or U22664 (N_22664,N_22425,N_21781);
and U22665 (N_22665,N_22354,N_22456);
nor U22666 (N_22666,N_21618,N_21471);
nor U22667 (N_22667,N_21637,N_22216);
or U22668 (N_22668,N_21749,N_22229);
nand U22669 (N_22669,N_21635,N_21251);
or U22670 (N_22670,N_22346,N_22178);
and U22671 (N_22671,N_21740,N_21371);
xnor U22672 (N_22672,N_21449,N_21523);
or U22673 (N_22673,N_21767,N_22208);
or U22674 (N_22674,N_21333,N_22482);
and U22675 (N_22675,N_21513,N_21682);
and U22676 (N_22676,N_22214,N_22086);
and U22677 (N_22677,N_22404,N_22061);
xnor U22678 (N_22678,N_22218,N_22232);
or U22679 (N_22679,N_22221,N_22258);
and U22680 (N_22680,N_22098,N_22176);
and U22681 (N_22681,N_22309,N_21613);
or U22682 (N_22682,N_22133,N_22047);
xor U22683 (N_22683,N_21703,N_21594);
nor U22684 (N_22684,N_22116,N_21904);
xor U22685 (N_22685,N_21729,N_22310);
or U22686 (N_22686,N_21999,N_22415);
and U22687 (N_22687,N_21349,N_21713);
or U22688 (N_22688,N_21407,N_21605);
and U22689 (N_22689,N_22275,N_22200);
or U22690 (N_22690,N_21406,N_21939);
and U22691 (N_22691,N_22192,N_21383);
or U22692 (N_22692,N_21328,N_22295);
nor U22693 (N_22693,N_21698,N_21435);
and U22694 (N_22694,N_21560,N_22064);
nand U22695 (N_22695,N_22264,N_22374);
nor U22696 (N_22696,N_21679,N_22385);
or U22697 (N_22697,N_22153,N_22148);
or U22698 (N_22698,N_21954,N_22303);
nand U22699 (N_22699,N_21338,N_22138);
and U22700 (N_22700,N_21621,N_22465);
xor U22701 (N_22701,N_21584,N_21648);
nor U22702 (N_22702,N_22173,N_21574);
or U22703 (N_22703,N_21267,N_21696);
nand U22704 (N_22704,N_21597,N_21989);
or U22705 (N_22705,N_21423,N_21824);
and U22706 (N_22706,N_21646,N_21929);
xnor U22707 (N_22707,N_22306,N_21468);
and U22708 (N_22708,N_22266,N_22450);
nor U22709 (N_22709,N_22371,N_21986);
xor U22710 (N_22710,N_21395,N_22319);
and U22711 (N_22711,N_21711,N_22289);
or U22712 (N_22712,N_22156,N_22074);
or U22713 (N_22713,N_22353,N_21688);
nor U22714 (N_22714,N_21889,N_22175);
nand U22715 (N_22715,N_21819,N_22105);
xor U22716 (N_22716,N_21624,N_21848);
and U22717 (N_22717,N_21805,N_22065);
nor U22718 (N_22718,N_21610,N_21263);
xor U22719 (N_22719,N_22190,N_21754);
or U22720 (N_22720,N_21277,N_22085);
xnor U22721 (N_22721,N_21287,N_22152);
and U22722 (N_22722,N_22486,N_21792);
and U22723 (N_22723,N_21983,N_22400);
or U22724 (N_22724,N_21649,N_22472);
or U22725 (N_22725,N_21254,N_21964);
nand U22726 (N_22726,N_21664,N_21271);
and U22727 (N_22727,N_21479,N_21746);
xor U22728 (N_22728,N_21615,N_21282);
nor U22729 (N_22729,N_21461,N_21346);
nor U22730 (N_22730,N_22329,N_22022);
and U22731 (N_22731,N_22006,N_22290);
and U22732 (N_22732,N_22351,N_21791);
nor U22733 (N_22733,N_21498,N_21930);
nor U22734 (N_22734,N_21431,N_21376);
xor U22735 (N_22735,N_21373,N_21936);
and U22736 (N_22736,N_22398,N_21867);
nor U22737 (N_22737,N_21501,N_22338);
xor U22738 (N_22738,N_21532,N_22202);
nor U22739 (N_22739,N_21554,N_21356);
xnor U22740 (N_22740,N_21798,N_21306);
or U22741 (N_22741,N_21717,N_22372);
xor U22742 (N_22742,N_21567,N_22269);
and U22743 (N_22743,N_21926,N_21632);
nand U22744 (N_22744,N_22070,N_22182);
and U22745 (N_22745,N_22448,N_21847);
nand U22746 (N_22746,N_22119,N_22212);
and U22747 (N_22747,N_21266,N_21353);
nor U22748 (N_22748,N_22082,N_22391);
or U22749 (N_22749,N_21937,N_21375);
nor U22750 (N_22750,N_22055,N_22496);
nand U22751 (N_22751,N_21393,N_21529);
and U22752 (N_22752,N_21897,N_22460);
xor U22753 (N_22753,N_21307,N_21492);
and U22754 (N_22754,N_21465,N_21286);
nand U22755 (N_22755,N_21972,N_21483);
nor U22756 (N_22756,N_21726,N_21583);
or U22757 (N_22757,N_21866,N_22174);
xnor U22758 (N_22758,N_21878,N_21546);
xnor U22759 (N_22759,N_21861,N_21920);
xor U22760 (N_22760,N_22327,N_21273);
xor U22761 (N_22761,N_21906,N_22026);
nand U22762 (N_22762,N_21558,N_22219);
or U22763 (N_22763,N_21709,N_21622);
xnor U22764 (N_22764,N_22321,N_21446);
xnor U22765 (N_22765,N_22375,N_21432);
nor U22766 (N_22766,N_21718,N_21540);
xnor U22767 (N_22767,N_22313,N_21786);
and U22768 (N_22768,N_21755,N_21397);
and U22769 (N_22769,N_22168,N_21531);
nor U22770 (N_22770,N_21436,N_21410);
and U22771 (N_22771,N_22246,N_21485);
nor U22772 (N_22772,N_22406,N_21871);
nand U22773 (N_22773,N_21785,N_22125);
nor U22774 (N_22774,N_21256,N_21943);
nand U22775 (N_22775,N_21893,N_22335);
or U22776 (N_22776,N_21442,N_22268);
and U22777 (N_22777,N_22316,N_21914);
or U22778 (N_22778,N_21589,N_22462);
or U22779 (N_22779,N_21503,N_21752);
or U22780 (N_22780,N_21318,N_22466);
xor U22781 (N_22781,N_21634,N_21568);
or U22782 (N_22782,N_21592,N_22395);
xnor U22783 (N_22783,N_21915,N_21447);
or U22784 (N_22784,N_22299,N_21934);
nor U22785 (N_22785,N_21860,N_21768);
xor U22786 (N_22786,N_22287,N_22386);
and U22787 (N_22787,N_21950,N_21913);
or U22788 (N_22788,N_21669,N_22094);
or U22789 (N_22789,N_21668,N_21470);
or U22790 (N_22790,N_21475,N_21522);
or U22791 (N_22791,N_21300,N_22455);
xnor U22792 (N_22792,N_21384,N_21982);
and U22793 (N_22793,N_21883,N_22092);
xor U22794 (N_22794,N_22430,N_21654);
and U22795 (N_22795,N_21774,N_22197);
and U22796 (N_22796,N_22128,N_21326);
and U22797 (N_22797,N_22367,N_21480);
and U22798 (N_22798,N_22280,N_22315);
or U22799 (N_22799,N_21626,N_22349);
or U22800 (N_22800,N_21949,N_21551);
or U22801 (N_22801,N_21639,N_21454);
nand U22802 (N_22802,N_22376,N_21619);
and U22803 (N_22803,N_21802,N_22461);
xor U22804 (N_22804,N_21759,N_21686);
xor U22805 (N_22805,N_21517,N_21653);
nor U22806 (N_22806,N_21813,N_22388);
or U22807 (N_22807,N_22475,N_22018);
xor U22808 (N_22808,N_21486,N_21674);
xnor U22809 (N_22809,N_21971,N_21309);
xnor U22810 (N_22810,N_21875,N_21302);
nand U22811 (N_22811,N_22027,N_22431);
and U22812 (N_22812,N_21332,N_21655);
or U22813 (N_22813,N_21801,N_22343);
or U22814 (N_22814,N_22194,N_21440);
xnor U22815 (N_22815,N_21358,N_22203);
and U22816 (N_22816,N_21544,N_22288);
or U22817 (N_22817,N_21716,N_21869);
xor U22818 (N_22818,N_22253,N_22478);
xnor U22819 (N_22819,N_21429,N_21313);
xnor U22820 (N_22820,N_21784,N_21985);
nand U22821 (N_22821,N_22120,N_21800);
nor U22822 (N_22822,N_21576,N_21736);
nor U22823 (N_22823,N_21348,N_21995);
nand U22824 (N_22824,N_21323,N_21545);
xnor U22825 (N_22825,N_22177,N_22390);
nor U22826 (N_22826,N_22251,N_21967);
xor U22827 (N_22827,N_21587,N_22118);
and U22828 (N_22828,N_21658,N_21836);
or U22829 (N_22829,N_22314,N_22433);
or U22830 (N_22830,N_21270,N_22014);
nor U22831 (N_22831,N_22110,N_21488);
and U22832 (N_22832,N_21623,N_21961);
nor U22833 (N_22833,N_22076,N_22330);
or U22834 (N_22834,N_22171,N_22419);
xor U22835 (N_22835,N_22083,N_21602);
or U22836 (N_22836,N_22102,N_21322);
and U22837 (N_22837,N_22442,N_21705);
or U22838 (N_22838,N_21775,N_21571);
xor U22839 (N_22839,N_21533,N_22025);
nor U22840 (N_22840,N_21416,N_22311);
nor U22841 (N_22841,N_21344,N_21330);
nor U22842 (N_22842,N_21661,N_22244);
nand U22843 (N_22843,N_21633,N_22423);
nand U22844 (N_22844,N_21992,N_22236);
and U22845 (N_22845,N_21441,N_21877);
nor U22846 (N_22846,N_22147,N_21733);
nand U22847 (N_22847,N_21666,N_21402);
nand U22848 (N_22848,N_21835,N_21738);
nor U22849 (N_22849,N_22111,N_21298);
xnor U22850 (N_22850,N_22300,N_21782);
nor U22851 (N_22851,N_21638,N_21343);
nor U22852 (N_22852,N_22439,N_21293);
and U22853 (N_22853,N_22015,N_22036);
or U22854 (N_22854,N_21690,N_22093);
and U22855 (N_22855,N_21556,N_21631);
and U22856 (N_22856,N_21722,N_22464);
or U22857 (N_22857,N_21899,N_22249);
nand U22858 (N_22858,N_22240,N_21296);
nor U22859 (N_22859,N_22359,N_21651);
xnor U22860 (N_22860,N_21289,N_22075);
xnor U22861 (N_22861,N_22066,N_22021);
or U22862 (N_22862,N_21314,N_21385);
nor U22863 (N_22863,N_22467,N_21527);
xnor U22864 (N_22864,N_22091,N_22095);
nor U22865 (N_22865,N_21347,N_21831);
nand U22866 (N_22866,N_22001,N_21317);
xor U22867 (N_22867,N_22379,N_21676);
nor U22868 (N_22868,N_22328,N_22228);
nor U22869 (N_22869,N_21911,N_22426);
xnor U22870 (N_22870,N_21499,N_21761);
and U22871 (N_22871,N_22407,N_21748);
or U22872 (N_22872,N_21991,N_21928);
xnor U22873 (N_22873,N_22458,N_21739);
xnor U22874 (N_22874,N_21643,N_22104);
xnor U22875 (N_22875,N_21844,N_21872);
nand U22876 (N_22876,N_21588,N_22493);
or U22877 (N_22877,N_21389,N_22344);
nor U22878 (N_22878,N_21978,N_21750);
and U22879 (N_22879,N_21957,N_22198);
xnor U22880 (N_22880,N_21630,N_21320);
or U22881 (N_22881,N_22348,N_21464);
xor U22882 (N_22882,N_22369,N_22271);
nor U22883 (N_22883,N_21530,N_22326);
and U22884 (N_22884,N_22445,N_21840);
or U22885 (N_22885,N_21873,N_21685);
nor U22886 (N_22886,N_21548,N_22172);
nor U22887 (N_22887,N_21250,N_21608);
nand U22888 (N_22888,N_21382,N_21809);
or U22889 (N_22889,N_21895,N_22129);
xnor U22890 (N_22890,N_21660,N_21569);
or U22891 (N_22891,N_21506,N_21476);
and U22892 (N_22892,N_21874,N_21453);
nand U22893 (N_22893,N_21391,N_22361);
nor U22894 (N_22894,N_22396,N_22164);
nor U22895 (N_22895,N_21463,N_22063);
nand U22896 (N_22896,N_22279,N_21959);
or U22897 (N_22897,N_22491,N_22003);
xor U22898 (N_22898,N_22334,N_22301);
nor U22899 (N_22899,N_21830,N_21744);
nor U22900 (N_22900,N_21580,N_21657);
nor U22901 (N_22901,N_21881,N_22020);
and U22902 (N_22902,N_22383,N_22255);
or U22903 (N_22903,N_21772,N_22444);
and U22904 (N_22904,N_21780,N_21652);
nor U22905 (N_22905,N_22473,N_22077);
nor U22906 (N_22906,N_21769,N_22023);
nor U22907 (N_22907,N_22205,N_22170);
and U22908 (N_22908,N_21857,N_21357);
or U22909 (N_22909,N_21927,N_21694);
nor U22910 (N_22910,N_22476,N_21681);
nor U22911 (N_22911,N_22122,N_21707);
nor U22912 (N_22912,N_21452,N_21508);
xor U22913 (N_22913,N_22484,N_21354);
xor U22914 (N_22914,N_22293,N_21398);
and U22915 (N_22915,N_22260,N_22399);
or U22916 (N_22916,N_21843,N_22294);
nor U22917 (N_22917,N_21799,N_21838);
xor U22918 (N_22918,N_22270,N_22495);
nor U22919 (N_22919,N_21386,N_21482);
or U22920 (N_22920,N_22420,N_21612);
nor U22921 (N_22921,N_21366,N_21689);
nor U22922 (N_22922,N_21301,N_22282);
nor U22923 (N_22923,N_21312,N_21788);
xor U22924 (N_22924,N_21285,N_21966);
nand U22925 (N_22925,N_22435,N_21553);
nor U22926 (N_22926,N_22474,N_22217);
xnor U22927 (N_22927,N_21363,N_21401);
and U22928 (N_22928,N_21582,N_22454);
nor U22929 (N_22929,N_21918,N_21628);
or U22930 (N_22930,N_21265,N_22336);
and U22931 (N_22931,N_21579,N_22410);
xnor U22932 (N_22932,N_21607,N_21336);
nand U22933 (N_22933,N_22286,N_22161);
xor U22934 (N_22934,N_22155,N_21274);
nand U22935 (N_22935,N_22146,N_21294);
nand U22936 (N_22936,N_21962,N_22068);
and U22937 (N_22937,N_21993,N_21477);
xnor U22938 (N_22938,N_22278,N_22238);
or U22939 (N_22939,N_21751,N_22397);
and U22940 (N_22940,N_22078,N_21891);
nand U22941 (N_22941,N_21902,N_22087);
nor U22942 (N_22942,N_21864,N_21319);
and U22943 (N_22943,N_21362,N_22144);
nand U22944 (N_22944,N_22409,N_22413);
xor U22945 (N_22945,N_21459,N_22488);
nand U22946 (N_22946,N_21535,N_22469);
xor U22947 (N_22947,N_21816,N_21487);
nor U22948 (N_22948,N_21856,N_22356);
or U22949 (N_22949,N_22283,N_21381);
nand U22950 (N_22950,N_21968,N_22160);
or U22951 (N_22951,N_21334,N_21497);
and U22952 (N_22952,N_21945,N_21955);
nor U22953 (N_22953,N_21821,N_21854);
nor U22954 (N_22954,N_21329,N_21719);
nor U22955 (N_22955,N_21647,N_22099);
nor U22956 (N_22956,N_21762,N_22114);
nand U22957 (N_22957,N_22401,N_21521);
or U22958 (N_22958,N_22048,N_21640);
xor U22959 (N_22959,N_22447,N_21342);
nand U22960 (N_22960,N_22243,N_22241);
or U22961 (N_22961,N_21841,N_21387);
xor U22962 (N_22962,N_21779,N_21735);
or U22963 (N_22963,N_21413,N_21491);
nand U22964 (N_22964,N_22159,N_21842);
xnor U22965 (N_22965,N_21963,N_22490);
nor U22966 (N_22966,N_21952,N_22245);
or U22967 (N_22967,N_22101,N_22030);
or U22968 (N_22968,N_22142,N_22362);
and U22969 (N_22969,N_22324,N_22206);
nand U22970 (N_22970,N_22004,N_22308);
or U22971 (N_22971,N_21514,N_21870);
nor U22972 (N_22972,N_21283,N_22332);
and U22973 (N_22973,N_22247,N_22029);
or U22974 (N_22974,N_21335,N_21272);
nand U22975 (N_22975,N_21818,N_21555);
and U22976 (N_22976,N_22471,N_21426);
xor U22977 (N_22977,N_22363,N_21260);
xnor U22978 (N_22978,N_21981,N_21409);
or U22979 (N_22979,N_22481,N_22451);
nand U22980 (N_22980,N_22276,N_21562);
nand U22981 (N_22981,N_22470,N_21627);
and U22982 (N_22982,N_22041,N_21278);
nor U22983 (N_22983,N_22453,N_21656);
or U22984 (N_22984,N_21351,N_22489);
nor U22985 (N_22985,N_21379,N_22188);
and U22986 (N_22986,N_22038,N_22384);
or U22987 (N_22987,N_22184,N_21305);
nor U22988 (N_22988,N_21670,N_22428);
nand U22989 (N_22989,N_22223,N_21290);
nor U22990 (N_22990,N_22084,N_21255);
and U22991 (N_22991,N_21953,N_21741);
nand U22992 (N_22992,N_22049,N_21776);
xor U22993 (N_22993,N_22487,N_22158);
nand U22994 (N_22994,N_22254,N_21742);
or U22995 (N_22995,N_22073,N_22163);
or U22996 (N_22996,N_21691,N_22196);
nand U22997 (N_22997,N_21505,N_22434);
xnor U22998 (N_22998,N_21790,N_21422);
or U22999 (N_22999,N_21478,N_21565);
nor U23000 (N_23000,N_21806,N_21976);
nand U23001 (N_23001,N_22181,N_21766);
nor U23002 (N_23002,N_22121,N_21845);
nor U23003 (N_23003,N_21879,N_22046);
nor U23004 (N_23004,N_21907,N_21975);
or U23005 (N_23005,N_21340,N_21796);
nor U23006 (N_23006,N_21979,N_22230);
and U23007 (N_23007,N_21578,N_21905);
nand U23008 (N_23008,N_21456,N_21596);
xnor U23009 (N_23009,N_22112,N_22019);
or U23010 (N_23010,N_21511,N_21509);
and U23011 (N_23011,N_21549,N_21974);
nor U23012 (N_23012,N_22483,N_22224);
nand U23013 (N_23013,N_21684,N_21886);
nand U23014 (N_23014,N_21828,N_21374);
and U23015 (N_23015,N_21804,N_21702);
nor U23016 (N_23016,N_21369,N_22210);
xor U23017 (N_23017,N_21795,N_22274);
and U23018 (N_23018,N_22494,N_22016);
nand U23019 (N_23019,N_21888,N_22139);
or U23020 (N_23020,N_21394,N_22106);
xor U23021 (N_23021,N_21337,N_21339);
nor U23022 (N_23022,N_22304,N_21868);
or U23023 (N_23023,N_21262,N_21935);
nand U23024 (N_23024,N_21252,N_21504);
or U23025 (N_23025,N_21756,N_22002);
xor U23026 (N_23026,N_21712,N_22449);
nand U23027 (N_23027,N_21941,N_21481);
xor U23028 (N_23028,N_22031,N_22365);
or U23029 (N_23029,N_21708,N_21288);
xor U23030 (N_23030,N_21765,N_22302);
nor U23031 (N_23031,N_21292,N_21721);
and U23032 (N_23032,N_22325,N_21591);
nand U23033 (N_23033,N_22054,N_21559);
or U23034 (N_23034,N_22234,N_21894);
nor U23035 (N_23035,N_21424,N_22035);
or U23036 (N_23036,N_21699,N_22296);
or U23037 (N_23037,N_22446,N_22267);
nand U23038 (N_23038,N_21516,N_21829);
nand U23039 (N_23039,N_22180,N_21518);
nor U23040 (N_23040,N_21910,N_21912);
nor U23041 (N_23041,N_22017,N_21730);
xnor U23042 (N_23042,N_21570,N_21408);
xor U23043 (N_23043,N_22000,N_21405);
and U23044 (N_23044,N_22417,N_21457);
and U23045 (N_23045,N_22265,N_22130);
nor U23046 (N_23046,N_22292,N_22256);
nand U23047 (N_23047,N_21321,N_21448);
or U23048 (N_23048,N_21280,N_22032);
and U23049 (N_23049,N_21697,N_21644);
nor U23050 (N_23050,N_22167,N_21903);
nand U23051 (N_23051,N_22285,N_21855);
or U23052 (N_23052,N_21577,N_22100);
and U23053 (N_23053,N_22352,N_21603);
or U23054 (N_23054,N_22136,N_21604);
nand U23055 (N_23055,N_21539,N_21507);
nand U23056 (N_23056,N_21970,N_21557);
and U23057 (N_23057,N_21671,N_22373);
xnor U23058 (N_23058,N_22057,N_22358);
or U23059 (N_23059,N_22213,N_21418);
or U23060 (N_23060,N_21743,N_22307);
xnor U23061 (N_23061,N_22440,N_21673);
and U23062 (N_23062,N_21420,N_21388);
xnor U23063 (N_23063,N_21642,N_21851);
xnor U23064 (N_23064,N_21359,N_22422);
nand U23065 (N_23065,N_22169,N_22227);
xor U23066 (N_23066,N_21701,N_21444);
xnor U23067 (N_23067,N_21922,N_21822);
nor U23068 (N_23068,N_21467,N_21581);
nor U23069 (N_23069,N_21345,N_22204);
nor U23070 (N_23070,N_22010,N_22438);
or U23071 (N_23071,N_21585,N_22209);
xnor U23072 (N_23072,N_21403,N_21484);
or U23073 (N_23073,N_21771,N_22355);
or U23074 (N_23074,N_22090,N_21812);
xor U23075 (N_23075,N_21474,N_22226);
and U23076 (N_23076,N_22416,N_22225);
and U23077 (N_23077,N_22053,N_22124);
or U23078 (N_23078,N_22137,N_21645);
and U23079 (N_23079,N_22089,N_22069);
nand U23080 (N_23080,N_21833,N_21360);
or U23081 (N_23081,N_22317,N_22071);
nor U23082 (N_23082,N_21919,N_21789);
and U23083 (N_23083,N_22056,N_22312);
nor U23084 (N_23084,N_22259,N_21908);
xnor U23085 (N_23085,N_21563,N_22126);
xnor U23086 (N_23086,N_21984,N_21404);
nand U23087 (N_23087,N_21536,N_21341);
nand U23088 (N_23088,N_22005,N_21834);
or U23089 (N_23089,N_21520,N_21598);
and U23090 (N_23090,N_22291,N_22050);
nor U23091 (N_23091,N_21808,N_22135);
and U23092 (N_23092,N_22115,N_21299);
xor U23093 (N_23093,N_21473,N_21763);
nor U23094 (N_23094,N_22191,N_21693);
xor U23095 (N_23095,N_21586,N_22141);
or U23096 (N_23096,N_22459,N_22380);
nand U23097 (N_23097,N_21826,N_21998);
nand U23098 (N_23098,N_21315,N_21732);
or U23099 (N_23099,N_22485,N_21977);
and U23100 (N_23100,N_21731,N_21710);
and U23101 (N_23101,N_21773,N_21609);
nor U23102 (N_23102,N_21421,N_21427);
and U23103 (N_23103,N_21575,N_21770);
and U23104 (N_23104,N_21839,N_21859);
nand U23105 (N_23105,N_21924,N_21960);
nor U23106 (N_23106,N_22499,N_22058);
and U23107 (N_23107,N_21261,N_22008);
or U23108 (N_23108,N_21327,N_22277);
nand U23109 (N_23109,N_21566,N_21695);
xor U23110 (N_23110,N_21443,N_21852);
nor U23111 (N_23111,N_22389,N_21493);
or U23112 (N_23112,N_21728,N_22437);
xnor U23113 (N_23113,N_22342,N_21938);
nand U23114 (N_23114,N_21814,N_21890);
nor U23115 (N_23115,N_21921,N_21850);
or U23116 (N_23116,N_21898,N_21887);
and U23117 (N_23117,N_22377,N_22323);
nor U23118 (N_23118,N_21472,N_22394);
nor U23119 (N_23119,N_21439,N_21614);
nor U23120 (N_23120,N_22350,N_21534);
and U23121 (N_23121,N_21994,N_22298);
and U23122 (N_23122,N_21678,N_21377);
nand U23123 (N_23123,N_22320,N_21629);
or U23124 (N_23124,N_21419,N_21951);
nor U23125 (N_23125,N_21510,N_22329);
and U23126 (N_23126,N_21337,N_21733);
and U23127 (N_23127,N_21976,N_21340);
xor U23128 (N_23128,N_21480,N_21496);
or U23129 (N_23129,N_21955,N_21780);
nand U23130 (N_23130,N_21291,N_21478);
or U23131 (N_23131,N_21250,N_21541);
xor U23132 (N_23132,N_22365,N_22429);
xnor U23133 (N_23133,N_21310,N_22262);
nor U23134 (N_23134,N_21844,N_21966);
and U23135 (N_23135,N_22280,N_21772);
and U23136 (N_23136,N_22296,N_22435);
xnor U23137 (N_23137,N_21531,N_21771);
nand U23138 (N_23138,N_21794,N_22209);
or U23139 (N_23139,N_21560,N_21522);
xor U23140 (N_23140,N_21567,N_21876);
and U23141 (N_23141,N_22368,N_22417);
nand U23142 (N_23142,N_21325,N_22381);
or U23143 (N_23143,N_21624,N_22111);
and U23144 (N_23144,N_21371,N_21274);
xnor U23145 (N_23145,N_21731,N_21836);
or U23146 (N_23146,N_21908,N_21674);
xor U23147 (N_23147,N_22358,N_21311);
xnor U23148 (N_23148,N_21679,N_22285);
or U23149 (N_23149,N_21413,N_21969);
nor U23150 (N_23150,N_21942,N_21957);
nor U23151 (N_23151,N_21520,N_21870);
xor U23152 (N_23152,N_21295,N_22453);
and U23153 (N_23153,N_21720,N_21799);
nor U23154 (N_23154,N_21955,N_21983);
and U23155 (N_23155,N_22340,N_22275);
xnor U23156 (N_23156,N_22020,N_22165);
nand U23157 (N_23157,N_22321,N_21984);
xnor U23158 (N_23158,N_21822,N_21563);
nand U23159 (N_23159,N_22389,N_21551);
nor U23160 (N_23160,N_21522,N_21929);
nand U23161 (N_23161,N_21540,N_22258);
xor U23162 (N_23162,N_21679,N_21954);
nand U23163 (N_23163,N_21339,N_22347);
nand U23164 (N_23164,N_21880,N_22176);
nor U23165 (N_23165,N_21904,N_22209);
xnor U23166 (N_23166,N_22404,N_21412);
nor U23167 (N_23167,N_22366,N_22010);
nor U23168 (N_23168,N_21743,N_21989);
xnor U23169 (N_23169,N_21892,N_21419);
nand U23170 (N_23170,N_22336,N_21736);
or U23171 (N_23171,N_21511,N_21768);
nand U23172 (N_23172,N_21622,N_21289);
nor U23173 (N_23173,N_21360,N_22057);
xor U23174 (N_23174,N_22496,N_21413);
nand U23175 (N_23175,N_22439,N_22024);
xor U23176 (N_23176,N_21723,N_22051);
or U23177 (N_23177,N_21663,N_21656);
nand U23178 (N_23178,N_21882,N_22072);
and U23179 (N_23179,N_21365,N_22471);
and U23180 (N_23180,N_22122,N_21344);
nand U23181 (N_23181,N_22141,N_22230);
nor U23182 (N_23182,N_21957,N_21662);
and U23183 (N_23183,N_21313,N_21549);
or U23184 (N_23184,N_22282,N_21274);
and U23185 (N_23185,N_21481,N_22051);
xnor U23186 (N_23186,N_21964,N_21461);
or U23187 (N_23187,N_21948,N_21400);
and U23188 (N_23188,N_21785,N_22134);
xor U23189 (N_23189,N_22046,N_21387);
nand U23190 (N_23190,N_22406,N_22454);
and U23191 (N_23191,N_21869,N_21641);
or U23192 (N_23192,N_21935,N_21385);
or U23193 (N_23193,N_21369,N_21555);
nand U23194 (N_23194,N_22288,N_21296);
nor U23195 (N_23195,N_21803,N_22209);
xor U23196 (N_23196,N_21716,N_22104);
nand U23197 (N_23197,N_21672,N_22162);
nor U23198 (N_23198,N_21349,N_22477);
nand U23199 (N_23199,N_22124,N_22349);
or U23200 (N_23200,N_22044,N_21289);
nand U23201 (N_23201,N_22282,N_21359);
nand U23202 (N_23202,N_22360,N_21408);
xor U23203 (N_23203,N_21773,N_22219);
and U23204 (N_23204,N_21948,N_22206);
and U23205 (N_23205,N_21679,N_22175);
xor U23206 (N_23206,N_21535,N_22272);
or U23207 (N_23207,N_21262,N_21347);
and U23208 (N_23208,N_22428,N_21325);
or U23209 (N_23209,N_22435,N_21762);
nand U23210 (N_23210,N_21640,N_22497);
and U23211 (N_23211,N_21380,N_21968);
nor U23212 (N_23212,N_21663,N_22197);
nand U23213 (N_23213,N_21870,N_21632);
xor U23214 (N_23214,N_21591,N_22086);
nor U23215 (N_23215,N_22350,N_21454);
or U23216 (N_23216,N_21380,N_21556);
or U23217 (N_23217,N_21907,N_21697);
and U23218 (N_23218,N_22059,N_21737);
xnor U23219 (N_23219,N_22470,N_21464);
nand U23220 (N_23220,N_22112,N_22362);
nand U23221 (N_23221,N_22088,N_21625);
nor U23222 (N_23222,N_22291,N_22148);
nor U23223 (N_23223,N_22367,N_21970);
nor U23224 (N_23224,N_22264,N_22063);
or U23225 (N_23225,N_21274,N_22096);
or U23226 (N_23226,N_21428,N_21264);
nor U23227 (N_23227,N_22058,N_21467);
or U23228 (N_23228,N_21401,N_22375);
xnor U23229 (N_23229,N_21950,N_21584);
xor U23230 (N_23230,N_21470,N_22349);
nor U23231 (N_23231,N_22357,N_21669);
xnor U23232 (N_23232,N_21546,N_21660);
nor U23233 (N_23233,N_22018,N_22053);
nand U23234 (N_23234,N_21781,N_21422);
nand U23235 (N_23235,N_22450,N_21865);
nand U23236 (N_23236,N_22209,N_21707);
xor U23237 (N_23237,N_22222,N_22433);
nor U23238 (N_23238,N_21332,N_21562);
nor U23239 (N_23239,N_22322,N_21961);
nand U23240 (N_23240,N_22203,N_21960);
nand U23241 (N_23241,N_22383,N_21706);
nand U23242 (N_23242,N_22491,N_22064);
nand U23243 (N_23243,N_21378,N_21752);
nand U23244 (N_23244,N_21274,N_22303);
and U23245 (N_23245,N_22095,N_22289);
and U23246 (N_23246,N_21870,N_22374);
xor U23247 (N_23247,N_21721,N_22064);
xnor U23248 (N_23248,N_21837,N_22352);
or U23249 (N_23249,N_22064,N_21958);
nand U23250 (N_23250,N_22147,N_21690);
xor U23251 (N_23251,N_22085,N_22408);
nand U23252 (N_23252,N_22151,N_21839);
nor U23253 (N_23253,N_22184,N_21448);
or U23254 (N_23254,N_21346,N_21567);
and U23255 (N_23255,N_21938,N_21458);
xor U23256 (N_23256,N_22461,N_21766);
nand U23257 (N_23257,N_21539,N_21616);
xnor U23258 (N_23258,N_21677,N_22025);
and U23259 (N_23259,N_21280,N_22064);
or U23260 (N_23260,N_21662,N_22054);
and U23261 (N_23261,N_22059,N_22238);
nor U23262 (N_23262,N_21715,N_21988);
nor U23263 (N_23263,N_21737,N_21855);
nor U23264 (N_23264,N_21796,N_21883);
and U23265 (N_23265,N_22233,N_21552);
xnor U23266 (N_23266,N_22472,N_22105);
xor U23267 (N_23267,N_21584,N_21374);
and U23268 (N_23268,N_22102,N_21350);
xor U23269 (N_23269,N_22371,N_22357);
nand U23270 (N_23270,N_21286,N_22339);
xor U23271 (N_23271,N_22295,N_21522);
and U23272 (N_23272,N_22364,N_21510);
nand U23273 (N_23273,N_21522,N_21728);
xor U23274 (N_23274,N_22044,N_21338);
and U23275 (N_23275,N_21587,N_22006);
and U23276 (N_23276,N_21513,N_21961);
nor U23277 (N_23277,N_21591,N_22494);
or U23278 (N_23278,N_21833,N_21582);
or U23279 (N_23279,N_22347,N_22127);
nand U23280 (N_23280,N_21415,N_22074);
or U23281 (N_23281,N_21594,N_22408);
and U23282 (N_23282,N_22433,N_21690);
nor U23283 (N_23283,N_21373,N_21495);
and U23284 (N_23284,N_21649,N_22367);
nor U23285 (N_23285,N_21451,N_21317);
or U23286 (N_23286,N_21664,N_21962);
nand U23287 (N_23287,N_21404,N_22058);
and U23288 (N_23288,N_21954,N_21854);
or U23289 (N_23289,N_22033,N_21615);
nor U23290 (N_23290,N_22410,N_21510);
nor U23291 (N_23291,N_21846,N_22419);
or U23292 (N_23292,N_21636,N_22319);
and U23293 (N_23293,N_21718,N_21664);
nand U23294 (N_23294,N_21266,N_22482);
and U23295 (N_23295,N_21551,N_21584);
or U23296 (N_23296,N_21474,N_22344);
nand U23297 (N_23297,N_21369,N_22404);
xnor U23298 (N_23298,N_21764,N_21821);
and U23299 (N_23299,N_22363,N_21869);
nand U23300 (N_23300,N_21966,N_21984);
or U23301 (N_23301,N_22133,N_21508);
nand U23302 (N_23302,N_21839,N_21417);
nor U23303 (N_23303,N_21438,N_22069);
nand U23304 (N_23304,N_21259,N_21747);
xor U23305 (N_23305,N_22112,N_21754);
or U23306 (N_23306,N_21271,N_21939);
nand U23307 (N_23307,N_22269,N_21945);
and U23308 (N_23308,N_21941,N_21321);
xor U23309 (N_23309,N_21699,N_21462);
xor U23310 (N_23310,N_21634,N_21981);
and U23311 (N_23311,N_22323,N_21766);
nand U23312 (N_23312,N_21418,N_22241);
nor U23313 (N_23313,N_21652,N_21355);
nor U23314 (N_23314,N_22068,N_21286);
xor U23315 (N_23315,N_21530,N_21479);
nand U23316 (N_23316,N_22257,N_21811);
nor U23317 (N_23317,N_21943,N_22296);
and U23318 (N_23318,N_21667,N_21803);
nand U23319 (N_23319,N_22201,N_21283);
nand U23320 (N_23320,N_22175,N_22382);
or U23321 (N_23321,N_21697,N_22074);
or U23322 (N_23322,N_22276,N_21493);
and U23323 (N_23323,N_22040,N_22470);
xnor U23324 (N_23324,N_22433,N_21991);
nand U23325 (N_23325,N_21434,N_21562);
xor U23326 (N_23326,N_22291,N_22488);
nor U23327 (N_23327,N_21619,N_21961);
nand U23328 (N_23328,N_21358,N_22263);
and U23329 (N_23329,N_22076,N_21577);
and U23330 (N_23330,N_22333,N_21988);
nor U23331 (N_23331,N_21786,N_22008);
nor U23332 (N_23332,N_22432,N_21703);
xnor U23333 (N_23333,N_22049,N_21403);
xnor U23334 (N_23334,N_21745,N_22172);
nor U23335 (N_23335,N_21841,N_22464);
xnor U23336 (N_23336,N_22470,N_21530);
nor U23337 (N_23337,N_22385,N_21316);
xnor U23338 (N_23338,N_22448,N_21657);
and U23339 (N_23339,N_21844,N_21521);
xnor U23340 (N_23340,N_21435,N_21553);
or U23341 (N_23341,N_22096,N_22380);
or U23342 (N_23342,N_21887,N_21807);
and U23343 (N_23343,N_21566,N_21737);
or U23344 (N_23344,N_22185,N_21740);
and U23345 (N_23345,N_21951,N_21675);
or U23346 (N_23346,N_21446,N_22291);
nor U23347 (N_23347,N_21865,N_22204);
nand U23348 (N_23348,N_21894,N_21772);
and U23349 (N_23349,N_21898,N_21589);
and U23350 (N_23350,N_21951,N_21661);
xor U23351 (N_23351,N_21829,N_21756);
or U23352 (N_23352,N_21965,N_22170);
xnor U23353 (N_23353,N_21317,N_22084);
and U23354 (N_23354,N_22045,N_21381);
or U23355 (N_23355,N_21292,N_22389);
or U23356 (N_23356,N_22183,N_21351);
nor U23357 (N_23357,N_22110,N_21972);
xor U23358 (N_23358,N_21807,N_21827);
xnor U23359 (N_23359,N_22471,N_21785);
and U23360 (N_23360,N_21662,N_21578);
nand U23361 (N_23361,N_21750,N_22152);
and U23362 (N_23362,N_21823,N_22305);
or U23363 (N_23363,N_22176,N_22306);
or U23364 (N_23364,N_22204,N_21988);
or U23365 (N_23365,N_21780,N_21956);
nor U23366 (N_23366,N_21465,N_22328);
nor U23367 (N_23367,N_21286,N_21844);
nand U23368 (N_23368,N_22317,N_21779);
nand U23369 (N_23369,N_21283,N_22418);
nand U23370 (N_23370,N_22394,N_21710);
or U23371 (N_23371,N_22204,N_21776);
and U23372 (N_23372,N_21747,N_21695);
nand U23373 (N_23373,N_22096,N_21692);
nand U23374 (N_23374,N_21460,N_22389);
and U23375 (N_23375,N_21814,N_21859);
xnor U23376 (N_23376,N_22156,N_21888);
and U23377 (N_23377,N_22136,N_21439);
xor U23378 (N_23378,N_22414,N_21756);
nor U23379 (N_23379,N_21726,N_21627);
and U23380 (N_23380,N_22340,N_21522);
or U23381 (N_23381,N_21526,N_22158);
nand U23382 (N_23382,N_21487,N_22265);
nor U23383 (N_23383,N_21306,N_22318);
and U23384 (N_23384,N_22332,N_21832);
and U23385 (N_23385,N_22131,N_21360);
or U23386 (N_23386,N_21878,N_21548);
and U23387 (N_23387,N_22188,N_21698);
and U23388 (N_23388,N_21622,N_22156);
nand U23389 (N_23389,N_21966,N_21769);
or U23390 (N_23390,N_21367,N_22378);
or U23391 (N_23391,N_21348,N_22210);
nand U23392 (N_23392,N_21371,N_21948);
or U23393 (N_23393,N_21413,N_22270);
or U23394 (N_23394,N_21250,N_21691);
nor U23395 (N_23395,N_22256,N_21631);
and U23396 (N_23396,N_21899,N_21340);
nor U23397 (N_23397,N_22027,N_21424);
xnor U23398 (N_23398,N_21536,N_22089);
xor U23399 (N_23399,N_21844,N_22318);
nor U23400 (N_23400,N_22373,N_21905);
or U23401 (N_23401,N_22188,N_22032);
nor U23402 (N_23402,N_21728,N_21518);
nor U23403 (N_23403,N_21933,N_22064);
xnor U23404 (N_23404,N_21624,N_21665);
and U23405 (N_23405,N_22166,N_21598);
xnor U23406 (N_23406,N_22046,N_22037);
nand U23407 (N_23407,N_22094,N_22177);
and U23408 (N_23408,N_21711,N_21382);
and U23409 (N_23409,N_21788,N_22000);
or U23410 (N_23410,N_22031,N_21737);
and U23411 (N_23411,N_21580,N_22124);
or U23412 (N_23412,N_21874,N_22153);
or U23413 (N_23413,N_22087,N_21252);
nor U23414 (N_23414,N_22039,N_21753);
nand U23415 (N_23415,N_21345,N_21343);
nor U23416 (N_23416,N_22140,N_21437);
xnor U23417 (N_23417,N_21526,N_21946);
and U23418 (N_23418,N_21700,N_22427);
or U23419 (N_23419,N_21666,N_21617);
or U23420 (N_23420,N_21603,N_21843);
xnor U23421 (N_23421,N_21498,N_22255);
and U23422 (N_23422,N_22028,N_22055);
nor U23423 (N_23423,N_22109,N_21892);
or U23424 (N_23424,N_22492,N_21942);
and U23425 (N_23425,N_21359,N_22245);
and U23426 (N_23426,N_21829,N_22033);
and U23427 (N_23427,N_22434,N_22166);
xnor U23428 (N_23428,N_22366,N_21463);
and U23429 (N_23429,N_22179,N_21799);
and U23430 (N_23430,N_21258,N_21601);
and U23431 (N_23431,N_22111,N_21837);
or U23432 (N_23432,N_21962,N_22002);
nor U23433 (N_23433,N_21997,N_22091);
xnor U23434 (N_23434,N_21533,N_22293);
nand U23435 (N_23435,N_22357,N_22233);
nor U23436 (N_23436,N_22228,N_22208);
and U23437 (N_23437,N_21727,N_21710);
and U23438 (N_23438,N_22236,N_22108);
xor U23439 (N_23439,N_21970,N_22057);
xor U23440 (N_23440,N_21586,N_22395);
or U23441 (N_23441,N_21440,N_22374);
or U23442 (N_23442,N_21573,N_22073);
nand U23443 (N_23443,N_21782,N_21564);
or U23444 (N_23444,N_21906,N_22474);
xor U23445 (N_23445,N_21429,N_22064);
nor U23446 (N_23446,N_22471,N_22376);
nand U23447 (N_23447,N_22194,N_21645);
and U23448 (N_23448,N_22202,N_21664);
nand U23449 (N_23449,N_21832,N_21528);
nand U23450 (N_23450,N_21937,N_21598);
nand U23451 (N_23451,N_22401,N_22309);
and U23452 (N_23452,N_22319,N_21556);
or U23453 (N_23453,N_21880,N_21429);
nand U23454 (N_23454,N_22135,N_21296);
nand U23455 (N_23455,N_21305,N_21978);
xnor U23456 (N_23456,N_21497,N_21669);
nand U23457 (N_23457,N_22190,N_21257);
and U23458 (N_23458,N_22498,N_21756);
xor U23459 (N_23459,N_21656,N_22471);
or U23460 (N_23460,N_21471,N_21921);
xnor U23461 (N_23461,N_21455,N_22105);
xor U23462 (N_23462,N_22246,N_22179);
nand U23463 (N_23463,N_21730,N_21690);
and U23464 (N_23464,N_21738,N_22436);
xnor U23465 (N_23465,N_21717,N_21532);
nand U23466 (N_23466,N_21788,N_21521);
nand U23467 (N_23467,N_22061,N_22433);
nand U23468 (N_23468,N_21651,N_21411);
xnor U23469 (N_23469,N_21589,N_21728);
nor U23470 (N_23470,N_21483,N_22497);
xor U23471 (N_23471,N_21340,N_22113);
nor U23472 (N_23472,N_21890,N_21557);
or U23473 (N_23473,N_21529,N_22442);
xnor U23474 (N_23474,N_22252,N_22019);
xor U23475 (N_23475,N_21492,N_21574);
or U23476 (N_23476,N_21809,N_21650);
and U23477 (N_23477,N_22467,N_22113);
and U23478 (N_23478,N_21934,N_21266);
nor U23479 (N_23479,N_21821,N_21378);
nor U23480 (N_23480,N_22308,N_22137);
nand U23481 (N_23481,N_21656,N_21922);
or U23482 (N_23482,N_21734,N_21986);
or U23483 (N_23483,N_22478,N_22241);
nor U23484 (N_23484,N_21337,N_22101);
nor U23485 (N_23485,N_21437,N_21893);
nand U23486 (N_23486,N_22295,N_22202);
xnor U23487 (N_23487,N_21595,N_21670);
nand U23488 (N_23488,N_22138,N_22214);
and U23489 (N_23489,N_22027,N_22036);
nor U23490 (N_23490,N_21385,N_21754);
and U23491 (N_23491,N_21492,N_21802);
nor U23492 (N_23492,N_22161,N_21883);
or U23493 (N_23493,N_21306,N_21252);
and U23494 (N_23494,N_21958,N_21970);
and U23495 (N_23495,N_22077,N_21964);
and U23496 (N_23496,N_21574,N_22010);
and U23497 (N_23497,N_21274,N_21938);
nor U23498 (N_23498,N_21367,N_22261);
or U23499 (N_23499,N_22158,N_21665);
nand U23500 (N_23500,N_21878,N_21412);
nand U23501 (N_23501,N_21549,N_21692);
or U23502 (N_23502,N_22087,N_21713);
or U23503 (N_23503,N_22137,N_21423);
nor U23504 (N_23504,N_22040,N_21866);
nor U23505 (N_23505,N_22426,N_21755);
xor U23506 (N_23506,N_22391,N_21884);
nand U23507 (N_23507,N_21484,N_22146);
and U23508 (N_23508,N_21697,N_22281);
and U23509 (N_23509,N_22034,N_21798);
nor U23510 (N_23510,N_21888,N_21700);
and U23511 (N_23511,N_22195,N_22285);
nand U23512 (N_23512,N_21258,N_21643);
nor U23513 (N_23513,N_21603,N_21735);
nand U23514 (N_23514,N_21690,N_22366);
nor U23515 (N_23515,N_21893,N_21814);
nand U23516 (N_23516,N_22261,N_21262);
and U23517 (N_23517,N_22396,N_22354);
nor U23518 (N_23518,N_21555,N_21492);
or U23519 (N_23519,N_21546,N_21443);
and U23520 (N_23520,N_21638,N_22234);
xor U23521 (N_23521,N_22000,N_21362);
and U23522 (N_23522,N_21459,N_22337);
and U23523 (N_23523,N_21321,N_22136);
xor U23524 (N_23524,N_21845,N_21364);
xnor U23525 (N_23525,N_22449,N_21564);
nor U23526 (N_23526,N_22357,N_22034);
xnor U23527 (N_23527,N_22425,N_21478);
nor U23528 (N_23528,N_22469,N_21642);
and U23529 (N_23529,N_22170,N_21602);
xor U23530 (N_23530,N_22311,N_22183);
or U23531 (N_23531,N_22032,N_21534);
and U23532 (N_23532,N_21678,N_21280);
nand U23533 (N_23533,N_21868,N_21415);
and U23534 (N_23534,N_21994,N_21373);
xor U23535 (N_23535,N_22138,N_21380);
xor U23536 (N_23536,N_21773,N_22107);
nand U23537 (N_23537,N_22289,N_22313);
or U23538 (N_23538,N_21744,N_22219);
and U23539 (N_23539,N_21276,N_22445);
nor U23540 (N_23540,N_21956,N_21774);
nand U23541 (N_23541,N_21290,N_22205);
and U23542 (N_23542,N_22287,N_22325);
and U23543 (N_23543,N_21303,N_21366);
nand U23544 (N_23544,N_21910,N_22031);
and U23545 (N_23545,N_22259,N_22178);
xor U23546 (N_23546,N_21678,N_21889);
or U23547 (N_23547,N_21269,N_22356);
nor U23548 (N_23548,N_21392,N_21648);
and U23549 (N_23549,N_21769,N_22170);
xnor U23550 (N_23550,N_21253,N_21759);
xor U23551 (N_23551,N_22112,N_21584);
nand U23552 (N_23552,N_21301,N_22102);
nand U23553 (N_23553,N_21494,N_22355);
and U23554 (N_23554,N_21413,N_22015);
or U23555 (N_23555,N_22228,N_21528);
and U23556 (N_23556,N_22240,N_21583);
xor U23557 (N_23557,N_21456,N_22202);
xnor U23558 (N_23558,N_21895,N_22499);
and U23559 (N_23559,N_22431,N_21425);
xor U23560 (N_23560,N_22327,N_21514);
xnor U23561 (N_23561,N_21599,N_22322);
or U23562 (N_23562,N_21391,N_22391);
or U23563 (N_23563,N_21493,N_22212);
and U23564 (N_23564,N_21376,N_21604);
and U23565 (N_23565,N_22305,N_21558);
nand U23566 (N_23566,N_22254,N_22034);
nor U23567 (N_23567,N_21854,N_22087);
and U23568 (N_23568,N_21725,N_22418);
xnor U23569 (N_23569,N_22159,N_21548);
or U23570 (N_23570,N_22253,N_21548);
nand U23571 (N_23571,N_21474,N_21540);
and U23572 (N_23572,N_21252,N_22499);
nand U23573 (N_23573,N_21597,N_21838);
nand U23574 (N_23574,N_21801,N_22173);
and U23575 (N_23575,N_21848,N_21796);
or U23576 (N_23576,N_22438,N_21399);
and U23577 (N_23577,N_21639,N_21265);
and U23578 (N_23578,N_21757,N_22485);
xor U23579 (N_23579,N_22114,N_21344);
or U23580 (N_23580,N_21911,N_21990);
and U23581 (N_23581,N_22456,N_21886);
xnor U23582 (N_23582,N_21279,N_21679);
xor U23583 (N_23583,N_22339,N_22035);
nand U23584 (N_23584,N_22484,N_21861);
or U23585 (N_23585,N_21710,N_21951);
or U23586 (N_23586,N_22237,N_22002);
xor U23587 (N_23587,N_21662,N_21751);
or U23588 (N_23588,N_22230,N_22256);
or U23589 (N_23589,N_21748,N_22485);
nand U23590 (N_23590,N_22317,N_22313);
and U23591 (N_23591,N_21941,N_22439);
or U23592 (N_23592,N_21489,N_21388);
nand U23593 (N_23593,N_21982,N_21749);
or U23594 (N_23594,N_21726,N_21486);
and U23595 (N_23595,N_22103,N_22202);
and U23596 (N_23596,N_22284,N_22391);
nand U23597 (N_23597,N_22289,N_22031);
and U23598 (N_23598,N_22410,N_21928);
nand U23599 (N_23599,N_21581,N_21345);
or U23600 (N_23600,N_21497,N_22359);
nand U23601 (N_23601,N_21871,N_21846);
and U23602 (N_23602,N_21557,N_22143);
or U23603 (N_23603,N_22401,N_22113);
or U23604 (N_23604,N_21708,N_22162);
nor U23605 (N_23605,N_22342,N_21301);
nor U23606 (N_23606,N_21913,N_22215);
or U23607 (N_23607,N_21882,N_21318);
or U23608 (N_23608,N_21576,N_22152);
and U23609 (N_23609,N_22443,N_21262);
xnor U23610 (N_23610,N_22395,N_22130);
nor U23611 (N_23611,N_22077,N_22216);
nand U23612 (N_23612,N_21261,N_21821);
xor U23613 (N_23613,N_21628,N_21689);
or U23614 (N_23614,N_22412,N_21752);
nand U23615 (N_23615,N_21309,N_21904);
or U23616 (N_23616,N_21534,N_21514);
or U23617 (N_23617,N_22053,N_21302);
nor U23618 (N_23618,N_22084,N_21592);
nand U23619 (N_23619,N_22155,N_22011);
xnor U23620 (N_23620,N_22088,N_21368);
and U23621 (N_23621,N_21922,N_21324);
xor U23622 (N_23622,N_22012,N_21748);
nor U23623 (N_23623,N_21356,N_21899);
xor U23624 (N_23624,N_21353,N_22397);
nor U23625 (N_23625,N_22184,N_21695);
xor U23626 (N_23626,N_21269,N_21514);
and U23627 (N_23627,N_21310,N_22006);
xor U23628 (N_23628,N_22453,N_22262);
nand U23629 (N_23629,N_21781,N_21375);
xor U23630 (N_23630,N_21957,N_22391);
nand U23631 (N_23631,N_21692,N_21759);
and U23632 (N_23632,N_21773,N_22418);
or U23633 (N_23633,N_21613,N_22030);
xor U23634 (N_23634,N_22192,N_22180);
nor U23635 (N_23635,N_21617,N_22162);
xnor U23636 (N_23636,N_21666,N_22018);
nor U23637 (N_23637,N_21388,N_22446);
xnor U23638 (N_23638,N_22046,N_22228);
or U23639 (N_23639,N_21455,N_21460);
or U23640 (N_23640,N_22081,N_21327);
and U23641 (N_23641,N_21862,N_21316);
xor U23642 (N_23642,N_21630,N_21536);
and U23643 (N_23643,N_22497,N_21831);
nand U23644 (N_23644,N_22186,N_22061);
nand U23645 (N_23645,N_22096,N_22025);
or U23646 (N_23646,N_21342,N_21417);
nand U23647 (N_23647,N_21427,N_22271);
nand U23648 (N_23648,N_21534,N_22258);
xor U23649 (N_23649,N_22125,N_21866);
nor U23650 (N_23650,N_22371,N_21695);
nand U23651 (N_23651,N_22243,N_22177);
xnor U23652 (N_23652,N_21888,N_21496);
and U23653 (N_23653,N_21760,N_22018);
and U23654 (N_23654,N_21758,N_21572);
xor U23655 (N_23655,N_21956,N_21989);
nor U23656 (N_23656,N_21652,N_21801);
nor U23657 (N_23657,N_22333,N_21817);
and U23658 (N_23658,N_21696,N_21995);
nor U23659 (N_23659,N_22433,N_21892);
xor U23660 (N_23660,N_21268,N_21664);
nand U23661 (N_23661,N_21906,N_21566);
nand U23662 (N_23662,N_22385,N_22233);
xnor U23663 (N_23663,N_21490,N_22327);
and U23664 (N_23664,N_21661,N_22276);
nor U23665 (N_23665,N_21951,N_21380);
nor U23666 (N_23666,N_21307,N_22331);
nor U23667 (N_23667,N_21476,N_21934);
nor U23668 (N_23668,N_22339,N_21873);
and U23669 (N_23669,N_21769,N_21678);
nand U23670 (N_23670,N_21738,N_22341);
xnor U23671 (N_23671,N_21975,N_21712);
xor U23672 (N_23672,N_21617,N_21349);
xnor U23673 (N_23673,N_21880,N_22333);
nor U23674 (N_23674,N_22095,N_21467);
xnor U23675 (N_23675,N_22196,N_21357);
xor U23676 (N_23676,N_22059,N_22485);
nand U23677 (N_23677,N_21475,N_22365);
nor U23678 (N_23678,N_21445,N_22376);
xor U23679 (N_23679,N_21644,N_21342);
xnor U23680 (N_23680,N_21256,N_21461);
nand U23681 (N_23681,N_21628,N_21859);
nor U23682 (N_23682,N_22437,N_21488);
nand U23683 (N_23683,N_21412,N_21307);
nand U23684 (N_23684,N_22092,N_22360);
xnor U23685 (N_23685,N_21392,N_21339);
or U23686 (N_23686,N_21349,N_22049);
or U23687 (N_23687,N_22430,N_21717);
and U23688 (N_23688,N_21984,N_21480);
xnor U23689 (N_23689,N_21392,N_21525);
nor U23690 (N_23690,N_21786,N_21403);
or U23691 (N_23691,N_21764,N_21493);
and U23692 (N_23692,N_21742,N_21317);
nand U23693 (N_23693,N_21312,N_21757);
nand U23694 (N_23694,N_22388,N_21837);
and U23695 (N_23695,N_21730,N_21764);
xnor U23696 (N_23696,N_21930,N_21823);
xor U23697 (N_23697,N_22345,N_21816);
nor U23698 (N_23698,N_21902,N_21645);
or U23699 (N_23699,N_22480,N_21295);
nor U23700 (N_23700,N_21432,N_21307);
and U23701 (N_23701,N_21421,N_21503);
nand U23702 (N_23702,N_21688,N_21686);
xor U23703 (N_23703,N_21460,N_21711);
nand U23704 (N_23704,N_22284,N_21325);
or U23705 (N_23705,N_21983,N_22333);
and U23706 (N_23706,N_22179,N_21814);
or U23707 (N_23707,N_22050,N_22457);
and U23708 (N_23708,N_21631,N_22147);
or U23709 (N_23709,N_22443,N_22274);
nand U23710 (N_23710,N_22417,N_21857);
nand U23711 (N_23711,N_21682,N_21650);
nand U23712 (N_23712,N_21328,N_22336);
and U23713 (N_23713,N_21621,N_22094);
or U23714 (N_23714,N_22099,N_21315);
and U23715 (N_23715,N_22395,N_21849);
xor U23716 (N_23716,N_21291,N_22053);
nand U23717 (N_23717,N_21688,N_22036);
nor U23718 (N_23718,N_21925,N_22139);
xor U23719 (N_23719,N_22357,N_22167);
xor U23720 (N_23720,N_21278,N_22113);
or U23721 (N_23721,N_21856,N_22363);
or U23722 (N_23722,N_22353,N_21689);
or U23723 (N_23723,N_22205,N_21282);
xnor U23724 (N_23724,N_21918,N_21942);
or U23725 (N_23725,N_22247,N_21519);
and U23726 (N_23726,N_22273,N_21976);
or U23727 (N_23727,N_21626,N_21958);
xor U23728 (N_23728,N_21514,N_21342);
nor U23729 (N_23729,N_22120,N_21506);
xor U23730 (N_23730,N_21949,N_22143);
and U23731 (N_23731,N_22408,N_21849);
nor U23732 (N_23732,N_22153,N_21972);
xor U23733 (N_23733,N_21771,N_21951);
nand U23734 (N_23734,N_22166,N_21525);
or U23735 (N_23735,N_21621,N_21382);
nor U23736 (N_23736,N_22161,N_21943);
nor U23737 (N_23737,N_21700,N_21562);
nor U23738 (N_23738,N_21988,N_22322);
nor U23739 (N_23739,N_21921,N_22310);
nor U23740 (N_23740,N_22421,N_21346);
nand U23741 (N_23741,N_21312,N_22167);
xor U23742 (N_23742,N_21945,N_21852);
nand U23743 (N_23743,N_22482,N_22385);
nand U23744 (N_23744,N_22384,N_22129);
xor U23745 (N_23745,N_22323,N_21747);
nand U23746 (N_23746,N_22464,N_21918);
and U23747 (N_23747,N_21708,N_21784);
and U23748 (N_23748,N_21539,N_21973);
xor U23749 (N_23749,N_22023,N_21336);
xnor U23750 (N_23750,N_22924,N_22958);
nand U23751 (N_23751,N_22621,N_22540);
and U23752 (N_23752,N_23097,N_22663);
or U23753 (N_23753,N_22956,N_23143);
xnor U23754 (N_23754,N_22604,N_23559);
nor U23755 (N_23755,N_23413,N_22821);
xnor U23756 (N_23756,N_22874,N_22984);
xor U23757 (N_23757,N_23366,N_23256);
nand U23758 (N_23758,N_23354,N_22925);
nor U23759 (N_23759,N_23241,N_23575);
nor U23760 (N_23760,N_22862,N_23006);
nor U23761 (N_23761,N_22989,N_22948);
nor U23762 (N_23762,N_23152,N_22839);
xor U23763 (N_23763,N_23258,N_23374);
xnor U23764 (N_23764,N_22784,N_23588);
xor U23765 (N_23765,N_23333,N_23730);
xnor U23766 (N_23766,N_23326,N_23236);
or U23767 (N_23767,N_23500,N_23502);
xor U23768 (N_23768,N_23721,N_23393);
xor U23769 (N_23769,N_22754,N_23069);
and U23770 (N_23770,N_23388,N_23586);
nand U23771 (N_23771,N_23112,N_22899);
or U23772 (N_23772,N_23117,N_23705);
and U23773 (N_23773,N_22666,N_23528);
nor U23774 (N_23774,N_22584,N_23075);
nor U23775 (N_23775,N_22701,N_23183);
nand U23776 (N_23776,N_23059,N_23283);
nor U23777 (N_23777,N_23430,N_23179);
nand U23778 (N_23778,N_23564,N_22528);
nor U23779 (N_23779,N_23661,N_23002);
or U23780 (N_23780,N_22959,N_23450);
xor U23781 (N_23781,N_22826,N_22801);
nor U23782 (N_23782,N_22803,N_22601);
nor U23783 (N_23783,N_23307,N_23552);
xnor U23784 (N_23784,N_23154,N_23512);
nor U23785 (N_23785,N_22947,N_23306);
nor U23786 (N_23786,N_23071,N_23194);
or U23787 (N_23787,N_22673,N_23579);
and U23788 (N_23788,N_23297,N_23580);
or U23789 (N_23789,N_22976,N_23402);
nor U23790 (N_23790,N_23682,N_23554);
nand U23791 (N_23791,N_23400,N_23358);
xnor U23792 (N_23792,N_22715,N_23298);
nand U23793 (N_23793,N_23477,N_22648);
nand U23794 (N_23794,N_23475,N_22992);
nand U23795 (N_23795,N_23079,N_22689);
or U23796 (N_23796,N_22697,N_23033);
or U23797 (N_23797,N_23271,N_23234);
xor U23798 (N_23798,N_23441,N_23448);
nor U23799 (N_23799,N_22906,N_23318);
xor U23800 (N_23800,N_22572,N_23418);
and U23801 (N_23801,N_22664,N_23521);
xor U23802 (N_23802,N_22587,N_23092);
or U23803 (N_23803,N_22879,N_23699);
nor U23804 (N_23804,N_22716,N_23639);
nand U23805 (N_23805,N_23224,N_23733);
nand U23806 (N_23806,N_23381,N_22917);
nor U23807 (N_23807,N_23574,N_22990);
or U23808 (N_23808,N_23556,N_22759);
nand U23809 (N_23809,N_23540,N_23080);
nor U23810 (N_23810,N_22692,N_23166);
nor U23811 (N_23811,N_23604,N_23544);
xnor U23812 (N_23812,N_23195,N_23188);
xor U23813 (N_23813,N_22966,N_23596);
nor U23814 (N_23814,N_23395,N_22570);
xor U23815 (N_23815,N_22977,N_23009);
and U23816 (N_23816,N_22852,N_22964);
xor U23817 (N_23817,N_22619,N_23459);
xor U23818 (N_23818,N_22986,N_23683);
xnor U23819 (N_23819,N_23022,N_23165);
nand U23820 (N_23820,N_23669,N_23511);
nand U23821 (N_23821,N_22921,N_23386);
nand U23822 (N_23822,N_22571,N_22516);
and U23823 (N_23823,N_22972,N_22554);
and U23824 (N_23824,N_23200,N_23024);
xnor U23825 (N_23825,N_23504,N_23695);
nand U23826 (N_23826,N_22645,N_23285);
nor U23827 (N_23827,N_23626,N_23478);
xnor U23828 (N_23828,N_23222,N_22809);
nor U23829 (N_23829,N_22591,N_23676);
and U23830 (N_23830,N_23090,N_22951);
xor U23831 (N_23831,N_23719,N_23157);
nand U23832 (N_23832,N_22856,N_23207);
nand U23833 (N_23833,N_22789,N_23401);
or U23834 (N_23834,N_23199,N_22600);
xor U23835 (N_23835,N_23387,N_23688);
or U23836 (N_23836,N_22950,N_22548);
nor U23837 (N_23837,N_23738,N_22779);
xor U23838 (N_23838,N_23175,N_23216);
xnor U23839 (N_23839,N_23427,N_22647);
and U23840 (N_23840,N_22565,N_22502);
and U23841 (N_23841,N_23189,N_22883);
or U23842 (N_23842,N_22617,N_23264);
xor U23843 (N_23843,N_22919,N_22876);
nor U23844 (N_23844,N_23634,N_23573);
and U23845 (N_23845,N_23037,N_22740);
or U23846 (N_23846,N_23254,N_23398);
and U23847 (N_23847,N_23276,N_23630);
or U23848 (N_23848,N_23671,N_23220);
xnor U23849 (N_23849,N_22655,N_22892);
or U23850 (N_23850,N_22598,N_22590);
xor U23851 (N_23851,N_22824,N_22529);
nand U23852 (N_23852,N_23549,N_23693);
and U23853 (N_23853,N_22633,N_23225);
nand U23854 (N_23854,N_23066,N_22946);
xor U23855 (N_23855,N_22694,N_23308);
xnor U23856 (N_23856,N_22551,N_22806);
xor U23857 (N_23857,N_22967,N_23319);
nand U23858 (N_23858,N_23052,N_23168);
and U23859 (N_23859,N_22635,N_23729);
or U23860 (N_23860,N_23568,N_22653);
xor U23861 (N_23861,N_22766,N_23440);
nor U23862 (N_23862,N_23550,N_22707);
or U23863 (N_23863,N_23193,N_22684);
and U23864 (N_23864,N_23600,N_22616);
or U23865 (N_23865,N_23057,N_23660);
xor U23866 (N_23866,N_23372,N_23129);
nand U23867 (N_23867,N_23133,N_23042);
or U23868 (N_23868,N_23289,N_23268);
xnor U23869 (N_23869,N_23598,N_22912);
xor U23870 (N_23870,N_23299,N_23049);
nand U23871 (N_23871,N_23293,N_23063);
nand U23872 (N_23872,N_23023,N_23491);
and U23873 (N_23873,N_23359,N_22953);
xor U23874 (N_23874,N_22525,N_23313);
nor U23875 (N_23875,N_23294,N_23741);
xnor U23876 (N_23876,N_23192,N_22945);
nor U23877 (N_23877,N_22804,N_23247);
nor U23878 (N_23878,N_23099,N_22888);
or U23879 (N_23879,N_23583,N_23458);
and U23880 (N_23880,N_23235,N_22615);
nor U23881 (N_23881,N_22629,N_23186);
nor U23882 (N_23882,N_23601,N_22890);
and U23883 (N_23883,N_23507,N_22935);
and U23884 (N_23884,N_23499,N_23347);
nand U23885 (N_23885,N_22574,N_23217);
nor U23886 (N_23886,N_22726,N_22939);
xor U23887 (N_23887,N_23451,N_23173);
or U23888 (N_23888,N_22805,N_23396);
and U23889 (N_23889,N_23594,N_23365);
or U23890 (N_23890,N_23290,N_23265);
or U23891 (N_23891,N_23340,N_23134);
nor U23892 (N_23892,N_23467,N_23288);
and U23893 (N_23893,N_23013,N_22652);
and U23894 (N_23894,N_23722,N_23447);
or U23895 (N_23895,N_22886,N_23518);
or U23896 (N_23896,N_22911,N_23565);
xor U23897 (N_23897,N_22513,N_22757);
nor U23898 (N_23898,N_22781,N_22717);
nand U23899 (N_23899,N_22631,N_23085);
and U23900 (N_23900,N_23355,N_23102);
and U23901 (N_23901,N_22868,N_22792);
nor U23902 (N_23902,N_23370,N_23566);
nand U23903 (N_23903,N_23460,N_23449);
or U23904 (N_23904,N_23390,N_23015);
nand U23905 (N_23905,N_23261,N_22651);
nand U23906 (N_23906,N_23674,N_23132);
nor U23907 (N_23907,N_23690,N_23468);
and U23908 (N_23908,N_23051,N_23205);
xor U23909 (N_23909,N_23380,N_22910);
or U23910 (N_23910,N_22918,N_23602);
and U23911 (N_23911,N_23537,N_22749);
and U23912 (N_23912,N_22968,N_23481);
nor U23913 (N_23913,N_22987,N_22503);
or U23914 (N_23914,N_22567,N_23303);
nand U23915 (N_23915,N_23076,N_23629);
nand U23916 (N_23916,N_22535,N_22895);
and U23917 (N_23917,N_23399,N_22593);
nand U23918 (N_23918,N_23105,N_22931);
xor U23919 (N_23919,N_23487,N_23296);
xor U23920 (N_23920,N_23334,N_22514);
nand U23921 (N_23921,N_23167,N_23169);
or U23922 (N_23922,N_22793,N_23603);
or U23923 (N_23923,N_22699,N_23558);
nor U23924 (N_23924,N_22996,N_23182);
nor U23925 (N_23925,N_22705,N_22656);
nand U23926 (N_23926,N_22698,N_23109);
and U23927 (N_23927,N_22538,N_22864);
nor U23928 (N_23928,N_22612,N_23613);
nor U23929 (N_23929,N_22830,N_23520);
nor U23930 (N_23930,N_23532,N_23275);
and U23931 (N_23931,N_22929,N_22597);
nor U23932 (N_23932,N_23078,N_23489);
nor U23933 (N_23933,N_22880,N_23642);
xor U23934 (N_23934,N_22702,N_22547);
nor U23935 (N_23935,N_23198,N_22928);
nand U23936 (N_23936,N_22532,N_23170);
nand U23937 (N_23937,N_23547,N_22898);
or U23938 (N_23938,N_22873,N_22997);
and U23939 (N_23939,N_23280,N_22800);
and U23940 (N_23940,N_22506,N_22669);
nor U23941 (N_23941,N_23068,N_23171);
xor U23942 (N_23942,N_23151,N_22831);
or U23943 (N_23943,N_22797,N_23587);
or U23944 (N_23944,N_23245,N_23045);
and U23945 (N_23945,N_23464,N_22727);
and U23946 (N_23946,N_22802,N_23329);
and U23947 (N_23947,N_23272,N_22678);
nand U23948 (N_23948,N_23701,N_23067);
or U23949 (N_23949,N_23680,N_23437);
and U23950 (N_23950,N_23578,N_22933);
or U23951 (N_23951,N_22578,N_22541);
xnor U23952 (N_23952,N_22676,N_23367);
or U23953 (N_23953,N_23576,N_23316);
and U23954 (N_23954,N_22519,N_23715);
and U23955 (N_23955,N_23569,N_23727);
nor U23956 (N_23956,N_23230,N_23163);
and U23957 (N_23957,N_23156,N_23221);
nand U23958 (N_23958,N_22988,N_22739);
nand U23959 (N_23959,N_23332,N_23328);
and U23960 (N_23960,N_23710,N_22900);
xor U23961 (N_23961,N_23597,N_23726);
xor U23962 (N_23962,N_23589,N_22536);
and U23963 (N_23963,N_23043,N_22636);
or U23964 (N_23964,N_23346,N_22835);
xnor U23965 (N_23965,N_22552,N_23593);
nor U23966 (N_23966,N_23125,N_22782);
nand U23967 (N_23967,N_23749,N_23124);
and U23968 (N_23968,N_22825,N_22796);
and U23969 (N_23969,N_23608,N_22704);
or U23970 (N_23970,N_23331,N_23620);
or U23971 (N_23971,N_23214,N_22508);
nor U23972 (N_23972,N_22644,N_22575);
nor U23973 (N_23973,N_23571,N_22773);
nand U23974 (N_23974,N_22588,N_22654);
nor U23975 (N_23975,N_22668,N_22788);
or U23976 (N_23976,N_22563,N_23208);
xnor U23977 (N_23977,N_23716,N_22827);
nand U23978 (N_23978,N_22811,N_23403);
nand U23979 (N_23979,N_23177,N_23000);
or U23980 (N_23980,N_22973,N_23257);
or U23981 (N_23981,N_22559,N_23029);
nand U23982 (N_23982,N_23535,N_23591);
nand U23983 (N_23983,N_23570,N_23356);
or U23984 (N_23984,N_22776,N_23160);
nor U23985 (N_23985,N_22914,N_22661);
or U23986 (N_23986,N_22812,N_23384);
xnor U23987 (N_23987,N_22582,N_22542);
xnor U23988 (N_23988,N_22708,N_23667);
or U23989 (N_23989,N_23005,N_23628);
nand U23990 (N_23990,N_23582,N_22869);
xor U23991 (N_23991,N_23153,N_23496);
nand U23992 (N_23992,N_22814,N_23127);
xnor U23993 (N_23993,N_22557,N_22614);
xor U23994 (N_23994,N_23323,N_23229);
nand U23995 (N_23995,N_23697,N_23414);
nor U23996 (N_23996,N_22837,N_23244);
nor U23997 (N_23997,N_23243,N_22760);
and U23998 (N_23998,N_23662,N_22863);
or U23999 (N_23999,N_23016,N_23083);
and U24000 (N_24000,N_22738,N_23126);
nand U24001 (N_24001,N_23149,N_23300);
nand U24002 (N_24002,N_23344,N_22768);
nand U24003 (N_24003,N_23562,N_23702);
nand U24004 (N_24004,N_23108,N_22683);
and U24005 (N_24005,N_23203,N_22783);
and U24006 (N_24006,N_23526,N_22944);
or U24007 (N_24007,N_23546,N_23618);
or U24008 (N_24008,N_23514,N_23737);
nor U24009 (N_24009,N_23648,N_22954);
nand U24010 (N_24010,N_22670,N_22596);
nor U24011 (N_24011,N_23379,N_23336);
and U24012 (N_24012,N_22696,N_23302);
and U24013 (N_24013,N_22628,N_22555);
or U24014 (N_24014,N_23641,N_22808);
nor U24015 (N_24015,N_23227,N_22969);
nor U24016 (N_24016,N_22905,N_22690);
nor U24017 (N_24017,N_23627,N_22936);
xor U24018 (N_24018,N_23426,N_23098);
and U24019 (N_24019,N_23010,N_23349);
and U24020 (N_24020,N_22657,N_23653);
and U24021 (N_24021,N_23656,N_23461);
xnor U24022 (N_24022,N_23025,N_23056);
nor U24023 (N_24023,N_23508,N_22855);
or U24024 (N_24024,N_23250,N_23073);
nor U24025 (N_24025,N_22703,N_22624);
or U24026 (N_24026,N_23012,N_22734);
nor U24027 (N_24027,N_22832,N_23538);
nand U24028 (N_24028,N_22998,N_23455);
nor U24029 (N_24029,N_22724,N_23158);
and U24030 (N_24030,N_23407,N_22711);
xnor U24031 (N_24031,N_23541,N_23637);
and U24032 (N_24032,N_23736,N_23095);
or U24033 (N_24033,N_23425,N_23341);
or U24034 (N_24034,N_23077,N_22840);
and U24035 (N_24035,N_23020,N_23466);
xnor U24036 (N_24036,N_22938,N_23647);
and U24037 (N_24037,N_23338,N_22626);
nor U24038 (N_24038,N_22706,N_22592);
nand U24039 (N_24039,N_23436,N_22751);
nand U24040 (N_24040,N_22957,N_22609);
and U24041 (N_24041,N_23592,N_23144);
nor U24042 (N_24042,N_22995,N_23429);
nor U24043 (N_24043,N_22822,N_23301);
or U24044 (N_24044,N_22819,N_22842);
xnor U24045 (N_24045,N_23501,N_22980);
and U24046 (N_24046,N_23219,N_23457);
nor U24047 (N_24047,N_23226,N_23633);
or U24048 (N_24048,N_22518,N_23120);
nor U24049 (N_24049,N_22870,N_23021);
nor U24050 (N_24050,N_22630,N_23202);
xnor U24051 (N_24051,N_23050,N_23419);
and U24052 (N_24052,N_23040,N_22894);
or U24053 (N_24053,N_22583,N_22564);
or U24054 (N_24054,N_23411,N_23624);
or U24055 (N_24055,N_23585,N_23255);
or U24056 (N_24056,N_22786,N_23492);
nand U24057 (N_24057,N_22533,N_23664);
nand U24058 (N_24058,N_22772,N_23391);
xor U24059 (N_24059,N_22861,N_22737);
nand U24060 (N_24060,N_23516,N_22896);
nand U24061 (N_24061,N_23339,N_23452);
or U24062 (N_24062,N_23191,N_22560);
nand U24063 (N_24063,N_22658,N_23375);
and U24064 (N_24064,N_22878,N_23704);
and U24065 (N_24065,N_22985,N_23612);
nor U24066 (N_24066,N_23616,N_23121);
nor U24067 (N_24067,N_23545,N_23432);
xnor U24068 (N_24068,N_23348,N_22761);
or U24069 (N_24069,N_22610,N_22817);
xnor U24070 (N_24070,N_22623,N_22723);
nand U24071 (N_24071,N_22775,N_23420);
nor U24072 (N_24072,N_23231,N_23096);
or U24073 (N_24073,N_23657,N_23228);
nor U24074 (N_24074,N_23482,N_23111);
nor U24075 (N_24075,N_22790,N_23707);
nor U24076 (N_24076,N_23542,N_23130);
nand U24077 (N_24077,N_23712,N_22764);
xor U24078 (N_24078,N_22729,N_22885);
or U24079 (N_24079,N_22753,N_22765);
and U24080 (N_24080,N_23438,N_22882);
nor U24081 (N_24081,N_23135,N_23287);
or U24082 (N_24082,N_23714,N_22643);
or U24083 (N_24083,N_22746,N_22889);
and U24084 (N_24084,N_22660,N_23061);
and U24085 (N_24085,N_23717,N_23211);
and U24086 (N_24086,N_23510,N_23665);
and U24087 (N_24087,N_23617,N_22970);
or U24088 (N_24088,N_22904,N_22755);
and U24089 (N_24089,N_23421,N_22915);
xor U24090 (N_24090,N_22920,N_23252);
or U24091 (N_24091,N_23406,N_22770);
nor U24092 (N_24092,N_22829,N_22975);
or U24093 (N_24093,N_22665,N_22569);
nand U24094 (N_24094,N_22586,N_22530);
or U24095 (N_24095,N_23218,N_23162);
and U24096 (N_24096,N_22730,N_23453);
nor U24097 (N_24097,N_23164,N_23089);
xor U24098 (N_24098,N_23343,N_23679);
nand U24099 (N_24099,N_22688,N_22700);
nand U24100 (N_24100,N_23476,N_23509);
xor U24101 (N_24101,N_22558,N_23035);
nor U24102 (N_24102,N_23106,N_23497);
xor U24103 (N_24103,N_22620,N_23039);
and U24104 (N_24104,N_23248,N_23531);
nand U24105 (N_24105,N_22504,N_22748);
and U24106 (N_24106,N_23315,N_22510);
nand U24107 (N_24107,N_22544,N_23139);
nor U24108 (N_24108,N_22871,N_23495);
or U24109 (N_24109,N_22679,N_22599);
xor U24110 (N_24110,N_23732,N_22983);
nor U24111 (N_24111,N_23394,N_22712);
nand U24112 (N_24112,N_23110,N_22934);
nor U24113 (N_24113,N_22971,N_23373);
nand U24114 (N_24114,N_23262,N_23278);
nand U24115 (N_24115,N_23734,N_23397);
xor U24116 (N_24116,N_22627,N_23524);
nor U24117 (N_24117,N_23743,N_22930);
nor U24118 (N_24118,N_23181,N_22500);
xnor U24119 (N_24119,N_23595,N_23353);
or U24120 (N_24120,N_23696,N_22941);
or U24121 (N_24121,N_23610,N_22763);
or U24122 (N_24122,N_22686,N_23655);
nor U24123 (N_24123,N_23363,N_23465);
nor U24124 (N_24124,N_22791,N_23703);
and U24125 (N_24125,N_23525,N_23041);
or U24126 (N_24126,N_22750,N_22999);
and U24127 (N_24127,N_22756,N_23515);
nor U24128 (N_24128,N_22893,N_23146);
xnor U24129 (N_24129,N_23176,N_23213);
xor U24130 (N_24130,N_23215,N_23074);
nor U24131 (N_24131,N_23150,N_23197);
and U24132 (N_24132,N_22642,N_22854);
and U24133 (N_24133,N_23141,N_22622);
xor U24134 (N_24134,N_23240,N_23223);
and U24135 (N_24135,N_23072,N_22675);
and U24136 (N_24136,N_23357,N_23654);
nor U24137 (N_24137,N_23590,N_23282);
nand U24138 (N_24138,N_23201,N_23113);
nor U24139 (N_24139,N_23027,N_23644);
or U24140 (N_24140,N_23560,N_23032);
nor U24141 (N_24141,N_23454,N_23003);
xnor U24142 (N_24142,N_22709,N_23337);
xnor U24143 (N_24143,N_23055,N_23670);
and U24144 (N_24144,N_22762,N_22795);
nand U24145 (N_24145,N_22594,N_23269);
xnor U24146 (N_24146,N_22522,N_23529);
xnor U24147 (N_24147,N_22877,N_23434);
nor U24148 (N_24148,N_23030,N_22962);
nor U24149 (N_24149,N_22866,N_23615);
nand U24150 (N_24150,N_23115,N_23431);
and U24151 (N_24151,N_23614,N_23446);
nor U24152 (N_24152,N_22807,N_23739);
nor U24153 (N_24153,N_23369,N_23048);
nor U24154 (N_24154,N_22942,N_23658);
and U24155 (N_24155,N_22539,N_22505);
xor U24156 (N_24156,N_23292,N_22721);
or U24157 (N_24157,N_23324,N_23607);
nand U24158 (N_24158,N_23118,N_22838);
and U24159 (N_24159,N_22521,N_22747);
and U24160 (N_24160,N_22847,N_22816);
nor U24161 (N_24161,N_22974,N_22515);
nor U24162 (N_24162,N_23563,N_22741);
and U24163 (N_24163,N_22507,N_23718);
or U24164 (N_24164,N_22693,N_23631);
or U24165 (N_24165,N_23327,N_22613);
or U24166 (N_24166,N_23689,N_23174);
xnor U24167 (N_24167,N_22566,N_22736);
or U24168 (N_24168,N_23038,N_23433);
xnor U24169 (N_24169,N_23577,N_23019);
nor U24170 (N_24170,N_23137,N_23708);
or U24171 (N_24171,N_22713,N_23103);
nand U24172 (N_24172,N_22537,N_23463);
and U24173 (N_24173,N_23304,N_23456);
or U24174 (N_24174,N_22672,N_23044);
nor U24175 (N_24175,N_23505,N_23543);
xor U24176 (N_24176,N_23686,N_23107);
xor U24177 (N_24177,N_23145,N_23249);
xor U24178 (N_24178,N_22843,N_23410);
xnor U24179 (N_24179,N_23081,N_23498);
or U24180 (N_24180,N_23483,N_23405);
nand U24181 (N_24181,N_22511,N_23101);
xor U24182 (N_24182,N_22714,N_23291);
and U24183 (N_24183,N_23148,N_23212);
or U24184 (N_24184,N_23709,N_22758);
xnor U24185 (N_24185,N_23747,N_22955);
or U24186 (N_24186,N_22733,N_23004);
and U24187 (N_24187,N_22602,N_22965);
xnor U24188 (N_24188,N_22815,N_22573);
or U24189 (N_24189,N_23321,N_22909);
nor U24190 (N_24190,N_23371,N_23428);
or U24191 (N_24191,N_23735,N_23519);
nor U24192 (N_24192,N_22891,N_22778);
and U24193 (N_24193,N_22650,N_23470);
nor U24194 (N_24194,N_23486,N_23204);
nand U24195 (N_24195,N_22674,N_23060);
and U24196 (N_24196,N_23530,N_23622);
nand U24197 (N_24197,N_23155,N_23746);
nand U24198 (N_24198,N_23485,N_22982);
and U24199 (N_24199,N_22677,N_23368);
or U24200 (N_24200,N_23522,N_22932);
nor U24201 (N_24201,N_23281,N_23311);
nor U24202 (N_24202,N_22794,N_23599);
and U24203 (N_24203,N_22682,N_23360);
xnor U24204 (N_24204,N_23691,N_23180);
nor U24205 (N_24205,N_22527,N_22845);
nand U24206 (N_24206,N_23026,N_23415);
and U24207 (N_24207,N_23266,N_23178);
and U24208 (N_24208,N_23445,N_23335);
nand U24209 (N_24209,N_23650,N_23422);
nand U24210 (N_24210,N_23377,N_23100);
xnor U24211 (N_24211,N_23136,N_23036);
xor U24212 (N_24212,N_22828,N_22545);
nand U24213 (N_24213,N_22785,N_23270);
xor U24214 (N_24214,N_22742,N_23123);
or U24215 (N_24215,N_22605,N_23645);
nor U24216 (N_24216,N_23493,N_23314);
and U24217 (N_24217,N_23251,N_22851);
nor U24218 (N_24218,N_23253,N_23484);
or U24219 (N_24219,N_23190,N_23273);
or U24220 (N_24220,N_23551,N_23416);
nand U24221 (N_24221,N_23104,N_23744);
or U24222 (N_24222,N_22625,N_23286);
and U24223 (N_24223,N_23533,N_23687);
and U24224 (N_24224,N_22952,N_22787);
and U24225 (N_24225,N_22848,N_22960);
xor U24226 (N_24226,N_23513,N_23119);
and U24227 (N_24227,N_22769,N_23084);
nor U24228 (N_24228,N_23128,N_22774);
nand U24229 (N_24229,N_23309,N_23404);
or U24230 (N_24230,N_22659,N_23122);
and U24231 (N_24231,N_23443,N_23675);
nand U24232 (N_24232,N_22908,N_22646);
or U24233 (N_24233,N_23088,N_23196);
xnor U24234 (N_24234,N_23317,N_22979);
nor U24235 (N_24235,N_23138,N_23720);
nor U24236 (N_24236,N_23014,N_23320);
or U24237 (N_24237,N_23635,N_22526);
or U24238 (N_24238,N_22901,N_23742);
and U24239 (N_24239,N_23274,N_23007);
xnor U24240 (N_24240,N_23330,N_23046);
and U24241 (N_24241,N_23444,N_22836);
nor U24242 (N_24242,N_23581,N_23408);
nor U24243 (N_24243,N_23263,N_22745);
nand U24244 (N_24244,N_23503,N_22581);
and U24245 (N_24245,N_22940,N_22813);
or U24246 (N_24246,N_23646,N_23527);
nand U24247 (N_24247,N_22720,N_22512);
nor U24248 (N_24248,N_23062,N_22534);
xnor U24249 (N_24249,N_23091,N_22833);
and U24250 (N_24250,N_23677,N_22916);
xnor U24251 (N_24251,N_23672,N_22860);
nand U24252 (N_24252,N_23439,N_22517);
nand U24253 (N_24253,N_22556,N_23724);
nor U24254 (N_24254,N_22608,N_22799);
or U24255 (N_24255,N_23116,N_22922);
nor U24256 (N_24256,N_23362,N_22949);
nor U24257 (N_24257,N_22913,N_22585);
xor U24258 (N_24258,N_23001,N_23442);
or U24259 (N_24259,N_22857,N_22927);
and U24260 (N_24260,N_22710,N_23536);
xor U24261 (N_24261,N_23094,N_22926);
or U24262 (N_24262,N_22577,N_23070);
nor U24263 (N_24263,N_22767,N_22897);
nand U24264 (N_24264,N_22872,N_22561);
nand U24265 (N_24265,N_22501,N_22991);
nand U24266 (N_24266,N_23553,N_23539);
nor U24267 (N_24267,N_23322,N_23623);
nand U24268 (N_24268,N_23206,N_22553);
nor U24269 (N_24269,N_23233,N_23728);
and U24270 (N_24270,N_22576,N_22865);
nor U24271 (N_24271,N_22725,N_23011);
xnor U24272 (N_24272,N_22743,N_23534);
nor U24273 (N_24273,N_22691,N_23209);
and U24274 (N_24274,N_22667,N_22771);
nor U24275 (N_24275,N_23567,N_22695);
or U24276 (N_24276,N_22637,N_23523);
or U24277 (N_24277,N_23047,N_22963);
nand U24278 (N_24278,N_22744,N_23706);
or U24279 (N_24279,N_22978,N_22632);
and U24280 (N_24280,N_23605,N_22606);
xnor U24281 (N_24281,N_22579,N_23008);
or U24282 (N_24282,N_22943,N_23424);
or U24283 (N_24283,N_23572,N_23711);
nand U24284 (N_24284,N_23259,N_23673);
nand U24285 (N_24285,N_23412,N_23018);
or U24286 (N_24286,N_22618,N_22640);
or U24287 (N_24287,N_22902,N_23237);
or U24288 (N_24288,N_23625,N_23017);
or U24289 (N_24289,N_23474,N_22611);
xor U24290 (N_24290,N_23694,N_22649);
and U24291 (N_24291,N_23409,N_23640);
nor U24292 (N_24292,N_22884,N_23611);
xor U24293 (N_24293,N_23305,N_23364);
xor U24294 (N_24294,N_23479,N_22719);
nor U24295 (N_24295,N_23246,N_23462);
nand U24296 (N_24296,N_23086,N_23668);
nand U24297 (N_24297,N_23494,N_23632);
or U24298 (N_24298,N_23636,N_23382);
nor U24299 (N_24299,N_23260,N_22728);
and U24300 (N_24300,N_23034,N_23725);
or U24301 (N_24301,N_23638,N_22685);
or U24302 (N_24302,N_23185,N_22858);
nand U24303 (N_24303,N_23184,N_23376);
xnor U24304 (N_24304,N_23417,N_23279);
nand U24305 (N_24305,N_23684,N_22820);
and U24306 (N_24306,N_23392,N_22607);
nand U24307 (N_24307,N_23093,N_22993);
nor U24308 (N_24308,N_22680,N_23389);
nand U24309 (N_24309,N_22994,N_23473);
xnor U24310 (N_24310,N_23748,N_22546);
or U24311 (N_24311,N_22589,N_22846);
xor U24312 (N_24312,N_23698,N_22881);
or U24313 (N_24313,N_22562,N_23685);
xor U24314 (N_24314,N_22735,N_23142);
or U24315 (N_24315,N_23385,N_22887);
and U24316 (N_24316,N_22777,N_23561);
nand U24317 (N_24317,N_23488,N_23310);
or U24318 (N_24318,N_22543,N_23210);
xnor U24319 (N_24319,N_23352,N_22523);
nor U24320 (N_24320,N_23147,N_23649);
nor U24321 (N_24321,N_22639,N_23350);
and U24322 (N_24322,N_23140,N_22752);
and U24323 (N_24323,N_23053,N_23490);
nand U24324 (N_24324,N_22520,N_22903);
nand U24325 (N_24325,N_23517,N_23740);
xor U24326 (N_24326,N_23471,N_22641);
xor U24327 (N_24327,N_22981,N_22687);
nand U24328 (N_24328,N_22844,N_23031);
nand U24329 (N_24329,N_23239,N_23087);
nand U24330 (N_24330,N_22731,N_23435);
or U24331 (N_24331,N_23383,N_23159);
and U24332 (N_24332,N_23284,N_22550);
xor U24333 (N_24333,N_23584,N_23663);
xor U24334 (N_24334,N_23342,N_23643);
and U24335 (N_24335,N_22722,N_23745);
nand U24336 (N_24336,N_23238,N_23609);
or U24337 (N_24337,N_23692,N_22849);
or U24338 (N_24338,N_22634,N_23713);
nand U24339 (N_24339,N_23666,N_22798);
and U24340 (N_24340,N_23506,N_23731);
nand U24341 (N_24341,N_23606,N_23351);
xor U24342 (N_24342,N_22638,N_23378);
nor U24343 (N_24343,N_22853,N_23555);
nand U24344 (N_24344,N_22671,N_22531);
and U24345 (N_24345,N_22732,N_22937);
nand U24346 (N_24346,N_22867,N_23082);
nand U24347 (N_24347,N_22875,N_23681);
nor U24348 (N_24348,N_23295,N_23557);
and U24349 (N_24349,N_22524,N_23423);
and U24350 (N_24350,N_22923,N_22841);
nand U24351 (N_24351,N_23131,N_23700);
xor U24352 (N_24352,N_23172,N_23054);
nor U24353 (N_24353,N_23469,N_23678);
and U24354 (N_24354,N_22603,N_22718);
or U24355 (N_24355,N_23345,N_22549);
or U24356 (N_24356,N_23277,N_23114);
xnor U24357 (N_24357,N_22823,N_23065);
nand U24358 (N_24358,N_23312,N_23472);
and U24359 (N_24359,N_22850,N_22595);
nand U24360 (N_24360,N_22818,N_23480);
and U24361 (N_24361,N_23058,N_23242);
or U24362 (N_24362,N_22859,N_23267);
and U24363 (N_24363,N_22580,N_22780);
and U24364 (N_24364,N_23361,N_22907);
and U24365 (N_24365,N_23028,N_22834);
nand U24366 (N_24366,N_22681,N_23325);
nand U24367 (N_24367,N_23619,N_22961);
or U24368 (N_24368,N_23232,N_23621);
or U24369 (N_24369,N_22810,N_23161);
nor U24370 (N_24370,N_23652,N_22568);
nand U24371 (N_24371,N_23723,N_22662);
and U24372 (N_24372,N_23064,N_23659);
nor U24373 (N_24373,N_23548,N_23187);
xnor U24374 (N_24374,N_22509,N_23651);
or U24375 (N_24375,N_23012,N_23276);
and U24376 (N_24376,N_23261,N_22660);
and U24377 (N_24377,N_23303,N_23601);
xor U24378 (N_24378,N_22958,N_22710);
and U24379 (N_24379,N_23120,N_23205);
xnor U24380 (N_24380,N_23089,N_23533);
nand U24381 (N_24381,N_23549,N_22679);
nor U24382 (N_24382,N_22658,N_22663);
nor U24383 (N_24383,N_23158,N_22594);
or U24384 (N_24384,N_23619,N_22534);
xnor U24385 (N_24385,N_23269,N_22590);
and U24386 (N_24386,N_23291,N_23586);
xnor U24387 (N_24387,N_23289,N_22859);
nand U24388 (N_24388,N_23073,N_22729);
or U24389 (N_24389,N_22956,N_23716);
xor U24390 (N_24390,N_23711,N_22712);
or U24391 (N_24391,N_23168,N_22554);
and U24392 (N_24392,N_22628,N_22812);
and U24393 (N_24393,N_23079,N_22707);
nand U24394 (N_24394,N_22559,N_22664);
nor U24395 (N_24395,N_23233,N_22651);
or U24396 (N_24396,N_22666,N_22793);
nand U24397 (N_24397,N_23207,N_22675);
xor U24398 (N_24398,N_23467,N_22634);
and U24399 (N_24399,N_23055,N_23323);
nor U24400 (N_24400,N_22909,N_23688);
nor U24401 (N_24401,N_22800,N_23419);
nor U24402 (N_24402,N_23461,N_23395);
xor U24403 (N_24403,N_23424,N_22983);
nor U24404 (N_24404,N_23613,N_23467);
nor U24405 (N_24405,N_22578,N_22627);
xnor U24406 (N_24406,N_22789,N_23174);
nand U24407 (N_24407,N_22612,N_23627);
xnor U24408 (N_24408,N_22920,N_22761);
or U24409 (N_24409,N_22870,N_23721);
or U24410 (N_24410,N_23070,N_22874);
or U24411 (N_24411,N_22629,N_23143);
or U24412 (N_24412,N_23325,N_23622);
xnor U24413 (N_24413,N_22509,N_23747);
xor U24414 (N_24414,N_22803,N_22755);
nor U24415 (N_24415,N_22803,N_22566);
xnor U24416 (N_24416,N_22968,N_23192);
and U24417 (N_24417,N_23025,N_22612);
nor U24418 (N_24418,N_23411,N_23332);
and U24419 (N_24419,N_23403,N_23566);
or U24420 (N_24420,N_23313,N_22888);
nand U24421 (N_24421,N_22695,N_22996);
and U24422 (N_24422,N_23287,N_23422);
and U24423 (N_24423,N_23515,N_22532);
and U24424 (N_24424,N_23546,N_22917);
xor U24425 (N_24425,N_22692,N_23310);
nor U24426 (N_24426,N_22812,N_22622);
or U24427 (N_24427,N_22745,N_23181);
nand U24428 (N_24428,N_23340,N_22814);
xnor U24429 (N_24429,N_23099,N_23280);
or U24430 (N_24430,N_22579,N_23303);
xnor U24431 (N_24431,N_23269,N_23017);
xnor U24432 (N_24432,N_22938,N_23479);
nor U24433 (N_24433,N_23187,N_23490);
or U24434 (N_24434,N_22519,N_23499);
xor U24435 (N_24435,N_23094,N_23476);
or U24436 (N_24436,N_23281,N_23749);
nand U24437 (N_24437,N_23159,N_22760);
and U24438 (N_24438,N_23584,N_23662);
or U24439 (N_24439,N_22945,N_22795);
and U24440 (N_24440,N_23028,N_23036);
and U24441 (N_24441,N_23422,N_22752);
nand U24442 (N_24442,N_23323,N_23538);
nor U24443 (N_24443,N_23493,N_22574);
xnor U24444 (N_24444,N_22723,N_23303);
xor U24445 (N_24445,N_23246,N_22851);
or U24446 (N_24446,N_23665,N_23501);
xor U24447 (N_24447,N_23239,N_23361);
xnor U24448 (N_24448,N_23649,N_23492);
or U24449 (N_24449,N_23444,N_23477);
and U24450 (N_24450,N_23512,N_23723);
or U24451 (N_24451,N_23436,N_22989);
or U24452 (N_24452,N_22603,N_23133);
or U24453 (N_24453,N_23386,N_23198);
and U24454 (N_24454,N_23295,N_23745);
and U24455 (N_24455,N_22830,N_23713);
nand U24456 (N_24456,N_23278,N_23495);
xnor U24457 (N_24457,N_23410,N_23442);
nor U24458 (N_24458,N_23150,N_23282);
or U24459 (N_24459,N_22808,N_22900);
xnor U24460 (N_24460,N_23298,N_23458);
xnor U24461 (N_24461,N_22947,N_23458);
xnor U24462 (N_24462,N_23192,N_22603);
nor U24463 (N_24463,N_22502,N_22870);
or U24464 (N_24464,N_23072,N_23098);
and U24465 (N_24465,N_23157,N_23438);
or U24466 (N_24466,N_22825,N_23022);
and U24467 (N_24467,N_22566,N_23592);
xor U24468 (N_24468,N_22784,N_23529);
nand U24469 (N_24469,N_23504,N_23421);
xor U24470 (N_24470,N_22698,N_23631);
xnor U24471 (N_24471,N_23085,N_23036);
and U24472 (N_24472,N_23511,N_23234);
or U24473 (N_24473,N_23664,N_23617);
xor U24474 (N_24474,N_22589,N_22758);
nor U24475 (N_24475,N_23069,N_23280);
and U24476 (N_24476,N_23140,N_23385);
and U24477 (N_24477,N_22635,N_22555);
and U24478 (N_24478,N_23029,N_23664);
or U24479 (N_24479,N_23697,N_23279);
xnor U24480 (N_24480,N_22513,N_23164);
xor U24481 (N_24481,N_22846,N_23068);
or U24482 (N_24482,N_22682,N_23313);
and U24483 (N_24483,N_22639,N_22629);
nor U24484 (N_24484,N_22741,N_22757);
and U24485 (N_24485,N_23520,N_22953);
xnor U24486 (N_24486,N_22724,N_23322);
or U24487 (N_24487,N_22801,N_22571);
xor U24488 (N_24488,N_23414,N_23367);
and U24489 (N_24489,N_22763,N_22639);
nor U24490 (N_24490,N_23310,N_22931);
nor U24491 (N_24491,N_23386,N_23689);
nor U24492 (N_24492,N_22891,N_23235);
nand U24493 (N_24493,N_22548,N_22631);
xnor U24494 (N_24494,N_23316,N_23230);
and U24495 (N_24495,N_23568,N_23631);
nor U24496 (N_24496,N_23162,N_23052);
nand U24497 (N_24497,N_23629,N_22525);
nand U24498 (N_24498,N_23654,N_22883);
nor U24499 (N_24499,N_23568,N_22745);
nor U24500 (N_24500,N_22547,N_23747);
nand U24501 (N_24501,N_23512,N_22588);
nand U24502 (N_24502,N_23356,N_23136);
nand U24503 (N_24503,N_23541,N_23318);
nor U24504 (N_24504,N_23000,N_23209);
xnor U24505 (N_24505,N_23720,N_23577);
nand U24506 (N_24506,N_23239,N_22504);
or U24507 (N_24507,N_23120,N_22637);
and U24508 (N_24508,N_23007,N_23302);
nor U24509 (N_24509,N_23114,N_23288);
and U24510 (N_24510,N_22930,N_22676);
and U24511 (N_24511,N_23618,N_22906);
or U24512 (N_24512,N_23712,N_22955);
or U24513 (N_24513,N_23554,N_23479);
nor U24514 (N_24514,N_23417,N_22729);
or U24515 (N_24515,N_22792,N_22556);
or U24516 (N_24516,N_23285,N_23522);
nand U24517 (N_24517,N_22950,N_23573);
nand U24518 (N_24518,N_23105,N_23576);
xor U24519 (N_24519,N_23106,N_23733);
nor U24520 (N_24520,N_22843,N_23433);
nor U24521 (N_24521,N_22591,N_23654);
or U24522 (N_24522,N_22675,N_23681);
or U24523 (N_24523,N_23482,N_23528);
nor U24524 (N_24524,N_23489,N_23053);
or U24525 (N_24525,N_22619,N_23392);
xnor U24526 (N_24526,N_23155,N_23430);
xor U24527 (N_24527,N_23608,N_23480);
and U24528 (N_24528,N_22669,N_22952);
xnor U24529 (N_24529,N_23427,N_22988);
nor U24530 (N_24530,N_22666,N_23224);
or U24531 (N_24531,N_23091,N_23557);
nand U24532 (N_24532,N_23501,N_23111);
or U24533 (N_24533,N_23165,N_23735);
nand U24534 (N_24534,N_23529,N_22715);
or U24535 (N_24535,N_23449,N_22646);
or U24536 (N_24536,N_22955,N_23334);
and U24537 (N_24537,N_23069,N_23569);
nor U24538 (N_24538,N_22960,N_23702);
xnor U24539 (N_24539,N_22679,N_23236);
and U24540 (N_24540,N_23157,N_23591);
or U24541 (N_24541,N_23465,N_23053);
and U24542 (N_24542,N_23603,N_23677);
xnor U24543 (N_24543,N_22531,N_23117);
or U24544 (N_24544,N_23638,N_23377);
nor U24545 (N_24545,N_22737,N_22924);
and U24546 (N_24546,N_22854,N_23204);
xor U24547 (N_24547,N_23061,N_23717);
or U24548 (N_24548,N_22708,N_22969);
nand U24549 (N_24549,N_23038,N_23260);
xor U24550 (N_24550,N_23380,N_23140);
nand U24551 (N_24551,N_22970,N_23682);
and U24552 (N_24552,N_23169,N_22722);
xnor U24553 (N_24553,N_23255,N_23308);
nand U24554 (N_24554,N_23469,N_23243);
xor U24555 (N_24555,N_23507,N_23108);
and U24556 (N_24556,N_23083,N_22598);
or U24557 (N_24557,N_23586,N_23456);
or U24558 (N_24558,N_23496,N_22624);
nand U24559 (N_24559,N_22725,N_22764);
or U24560 (N_24560,N_22568,N_23170);
nor U24561 (N_24561,N_23126,N_22862);
xor U24562 (N_24562,N_23274,N_22706);
and U24563 (N_24563,N_22617,N_23223);
xor U24564 (N_24564,N_22721,N_23657);
and U24565 (N_24565,N_22930,N_23121);
or U24566 (N_24566,N_22848,N_23432);
xnor U24567 (N_24567,N_22913,N_23159);
nand U24568 (N_24568,N_22524,N_22982);
and U24569 (N_24569,N_22831,N_22734);
nor U24570 (N_24570,N_23487,N_23600);
nand U24571 (N_24571,N_23569,N_23527);
or U24572 (N_24572,N_23061,N_23102);
or U24573 (N_24573,N_23525,N_23608);
nand U24574 (N_24574,N_22609,N_23269);
xor U24575 (N_24575,N_22657,N_23111);
or U24576 (N_24576,N_22584,N_23650);
and U24577 (N_24577,N_23302,N_23713);
or U24578 (N_24578,N_23058,N_23713);
nor U24579 (N_24579,N_23636,N_23152);
nor U24580 (N_24580,N_22890,N_22738);
or U24581 (N_24581,N_23562,N_23485);
nor U24582 (N_24582,N_22527,N_22618);
and U24583 (N_24583,N_23718,N_23264);
nor U24584 (N_24584,N_22710,N_22944);
xor U24585 (N_24585,N_23202,N_23748);
and U24586 (N_24586,N_22943,N_23705);
and U24587 (N_24587,N_23672,N_22681);
nor U24588 (N_24588,N_22525,N_23093);
xor U24589 (N_24589,N_22797,N_23385);
nand U24590 (N_24590,N_23658,N_23664);
or U24591 (N_24591,N_22639,N_23364);
xor U24592 (N_24592,N_23719,N_22690);
nor U24593 (N_24593,N_23302,N_22752);
and U24594 (N_24594,N_23002,N_23331);
and U24595 (N_24595,N_23197,N_22878);
nor U24596 (N_24596,N_23181,N_23274);
xnor U24597 (N_24597,N_23180,N_23656);
nor U24598 (N_24598,N_23599,N_22798);
and U24599 (N_24599,N_23292,N_22905);
nor U24600 (N_24600,N_22666,N_22579);
xnor U24601 (N_24601,N_23355,N_22832);
and U24602 (N_24602,N_23581,N_23318);
xnor U24603 (N_24603,N_23139,N_23276);
nor U24604 (N_24604,N_22553,N_23558);
and U24605 (N_24605,N_23338,N_23006);
nor U24606 (N_24606,N_23209,N_22636);
and U24607 (N_24607,N_23210,N_22508);
and U24608 (N_24608,N_22580,N_22838);
and U24609 (N_24609,N_23150,N_23058);
nor U24610 (N_24610,N_23038,N_22567);
nor U24611 (N_24611,N_23110,N_23280);
nand U24612 (N_24612,N_23155,N_23513);
nor U24613 (N_24613,N_23160,N_23195);
or U24614 (N_24614,N_22647,N_23399);
xnor U24615 (N_24615,N_22623,N_22914);
nand U24616 (N_24616,N_22903,N_23474);
or U24617 (N_24617,N_22561,N_22624);
nand U24618 (N_24618,N_22685,N_23382);
and U24619 (N_24619,N_23509,N_23626);
and U24620 (N_24620,N_23734,N_22552);
nor U24621 (N_24621,N_23214,N_22769);
nand U24622 (N_24622,N_22653,N_22893);
nand U24623 (N_24623,N_23228,N_23255);
nor U24624 (N_24624,N_22574,N_23344);
and U24625 (N_24625,N_22838,N_23342);
nor U24626 (N_24626,N_23369,N_23586);
or U24627 (N_24627,N_23110,N_23702);
xnor U24628 (N_24628,N_22892,N_22893);
nand U24629 (N_24629,N_23029,N_23584);
nand U24630 (N_24630,N_22569,N_23576);
or U24631 (N_24631,N_22953,N_22733);
nand U24632 (N_24632,N_23246,N_23393);
or U24633 (N_24633,N_22686,N_22558);
nand U24634 (N_24634,N_22928,N_23311);
nor U24635 (N_24635,N_23274,N_23361);
nor U24636 (N_24636,N_23461,N_22501);
nor U24637 (N_24637,N_23653,N_22533);
and U24638 (N_24638,N_22765,N_23351);
nand U24639 (N_24639,N_23519,N_22569);
or U24640 (N_24640,N_22631,N_22661);
nand U24641 (N_24641,N_22741,N_23617);
nor U24642 (N_24642,N_23597,N_23292);
or U24643 (N_24643,N_23480,N_23564);
or U24644 (N_24644,N_22949,N_22805);
and U24645 (N_24645,N_22968,N_23725);
or U24646 (N_24646,N_23175,N_23636);
nor U24647 (N_24647,N_23484,N_23307);
nor U24648 (N_24648,N_23587,N_22517);
nand U24649 (N_24649,N_23498,N_23159);
and U24650 (N_24650,N_23626,N_22525);
and U24651 (N_24651,N_23588,N_23608);
and U24652 (N_24652,N_23273,N_23428);
nand U24653 (N_24653,N_22608,N_23560);
and U24654 (N_24654,N_22779,N_23723);
or U24655 (N_24655,N_22506,N_23329);
and U24656 (N_24656,N_22948,N_23418);
nor U24657 (N_24657,N_22591,N_23222);
and U24658 (N_24658,N_22978,N_23410);
or U24659 (N_24659,N_22524,N_23140);
nor U24660 (N_24660,N_22820,N_23305);
and U24661 (N_24661,N_22703,N_23307);
nand U24662 (N_24662,N_23402,N_22848);
xor U24663 (N_24663,N_22541,N_23526);
and U24664 (N_24664,N_22672,N_23643);
or U24665 (N_24665,N_22823,N_23069);
xor U24666 (N_24666,N_23742,N_23457);
or U24667 (N_24667,N_22883,N_22688);
xnor U24668 (N_24668,N_23094,N_23661);
xnor U24669 (N_24669,N_22613,N_22501);
and U24670 (N_24670,N_23191,N_22982);
or U24671 (N_24671,N_23705,N_22960);
and U24672 (N_24672,N_23076,N_23033);
and U24673 (N_24673,N_22575,N_23316);
xnor U24674 (N_24674,N_23059,N_23159);
or U24675 (N_24675,N_22837,N_23665);
xor U24676 (N_24676,N_23256,N_22624);
xnor U24677 (N_24677,N_23366,N_22791);
and U24678 (N_24678,N_23376,N_22863);
nand U24679 (N_24679,N_22927,N_23658);
and U24680 (N_24680,N_22947,N_22950);
and U24681 (N_24681,N_23204,N_23019);
nor U24682 (N_24682,N_23511,N_23252);
or U24683 (N_24683,N_22735,N_23421);
or U24684 (N_24684,N_23420,N_23017);
nor U24685 (N_24685,N_23105,N_23648);
nand U24686 (N_24686,N_23159,N_22949);
nor U24687 (N_24687,N_22895,N_23481);
or U24688 (N_24688,N_22615,N_22890);
xnor U24689 (N_24689,N_23235,N_23368);
nand U24690 (N_24690,N_23630,N_23295);
and U24691 (N_24691,N_23476,N_23589);
or U24692 (N_24692,N_23418,N_23178);
nor U24693 (N_24693,N_23697,N_23430);
xor U24694 (N_24694,N_22570,N_23205);
or U24695 (N_24695,N_23237,N_22807);
nand U24696 (N_24696,N_22945,N_23585);
xnor U24697 (N_24697,N_23489,N_22889);
nor U24698 (N_24698,N_23011,N_23377);
nor U24699 (N_24699,N_23083,N_23310);
xnor U24700 (N_24700,N_23134,N_22945);
or U24701 (N_24701,N_23628,N_23206);
and U24702 (N_24702,N_22961,N_23643);
xnor U24703 (N_24703,N_23404,N_23244);
or U24704 (N_24704,N_22881,N_23524);
nand U24705 (N_24705,N_23157,N_22776);
and U24706 (N_24706,N_23015,N_22503);
and U24707 (N_24707,N_23502,N_23609);
nor U24708 (N_24708,N_23088,N_23110);
xnor U24709 (N_24709,N_23185,N_23440);
and U24710 (N_24710,N_22873,N_23654);
and U24711 (N_24711,N_22901,N_23718);
and U24712 (N_24712,N_23113,N_23404);
nand U24713 (N_24713,N_23660,N_22688);
or U24714 (N_24714,N_22725,N_22643);
and U24715 (N_24715,N_23308,N_23073);
nor U24716 (N_24716,N_22711,N_22843);
and U24717 (N_24717,N_23023,N_22771);
xor U24718 (N_24718,N_23299,N_22911);
and U24719 (N_24719,N_22694,N_22686);
xor U24720 (N_24720,N_23110,N_23151);
or U24721 (N_24721,N_23181,N_22908);
nand U24722 (N_24722,N_23229,N_22812);
nor U24723 (N_24723,N_22671,N_23104);
or U24724 (N_24724,N_22721,N_23320);
nor U24725 (N_24725,N_23342,N_23318);
nand U24726 (N_24726,N_22654,N_22842);
nor U24727 (N_24727,N_23268,N_23605);
nor U24728 (N_24728,N_23139,N_23225);
xor U24729 (N_24729,N_22887,N_22945);
xnor U24730 (N_24730,N_22957,N_23342);
and U24731 (N_24731,N_22709,N_22954);
or U24732 (N_24732,N_22527,N_22860);
xor U24733 (N_24733,N_23400,N_23090);
or U24734 (N_24734,N_23262,N_22794);
and U24735 (N_24735,N_22934,N_22878);
nand U24736 (N_24736,N_23131,N_23029);
nor U24737 (N_24737,N_23204,N_23507);
or U24738 (N_24738,N_22728,N_23324);
nand U24739 (N_24739,N_23595,N_22715);
xnor U24740 (N_24740,N_23690,N_22780);
nand U24741 (N_24741,N_23593,N_23518);
nor U24742 (N_24742,N_22907,N_22793);
or U24743 (N_24743,N_23470,N_23224);
xnor U24744 (N_24744,N_23353,N_23149);
xor U24745 (N_24745,N_23250,N_23461);
xor U24746 (N_24746,N_22980,N_23482);
nor U24747 (N_24747,N_22879,N_23187);
nor U24748 (N_24748,N_23597,N_23287);
and U24749 (N_24749,N_23325,N_22961);
and U24750 (N_24750,N_23447,N_23483);
nand U24751 (N_24751,N_22560,N_23341);
xor U24752 (N_24752,N_23744,N_23550);
nor U24753 (N_24753,N_22896,N_23084);
xnor U24754 (N_24754,N_23424,N_22787);
nand U24755 (N_24755,N_23230,N_22854);
and U24756 (N_24756,N_22978,N_23480);
and U24757 (N_24757,N_23522,N_22848);
nor U24758 (N_24758,N_23054,N_23692);
nand U24759 (N_24759,N_22600,N_23400);
xor U24760 (N_24760,N_23183,N_23375);
or U24761 (N_24761,N_23049,N_22749);
nor U24762 (N_24762,N_22785,N_23507);
and U24763 (N_24763,N_22823,N_23014);
nor U24764 (N_24764,N_23633,N_23396);
nand U24765 (N_24765,N_23318,N_23547);
nand U24766 (N_24766,N_23306,N_23731);
nand U24767 (N_24767,N_22685,N_23372);
xnor U24768 (N_24768,N_23692,N_22794);
xnor U24769 (N_24769,N_22579,N_22611);
xor U24770 (N_24770,N_22506,N_22763);
xor U24771 (N_24771,N_23686,N_23484);
nor U24772 (N_24772,N_23466,N_23139);
nor U24773 (N_24773,N_23013,N_23328);
nand U24774 (N_24774,N_22537,N_22582);
xor U24775 (N_24775,N_23067,N_23139);
or U24776 (N_24776,N_22549,N_23086);
nand U24777 (N_24777,N_23570,N_23223);
and U24778 (N_24778,N_22870,N_23716);
or U24779 (N_24779,N_23370,N_22952);
xor U24780 (N_24780,N_22644,N_22712);
nand U24781 (N_24781,N_23048,N_22699);
xor U24782 (N_24782,N_22788,N_22710);
xnor U24783 (N_24783,N_23315,N_23707);
or U24784 (N_24784,N_23647,N_23380);
xor U24785 (N_24785,N_23513,N_23116);
xnor U24786 (N_24786,N_23744,N_23745);
nor U24787 (N_24787,N_22897,N_23118);
nand U24788 (N_24788,N_22762,N_23544);
and U24789 (N_24789,N_23199,N_23227);
and U24790 (N_24790,N_23520,N_22640);
nor U24791 (N_24791,N_22924,N_22596);
or U24792 (N_24792,N_23324,N_23282);
or U24793 (N_24793,N_23661,N_23225);
and U24794 (N_24794,N_23490,N_23247);
nand U24795 (N_24795,N_22841,N_23147);
nand U24796 (N_24796,N_23411,N_23466);
or U24797 (N_24797,N_22527,N_22588);
and U24798 (N_24798,N_23258,N_22906);
nor U24799 (N_24799,N_22734,N_23681);
nor U24800 (N_24800,N_23415,N_23117);
or U24801 (N_24801,N_22981,N_23233);
nor U24802 (N_24802,N_23227,N_23412);
xor U24803 (N_24803,N_23411,N_22614);
nand U24804 (N_24804,N_23160,N_23545);
and U24805 (N_24805,N_23096,N_22621);
or U24806 (N_24806,N_23579,N_23724);
and U24807 (N_24807,N_22780,N_23691);
or U24808 (N_24808,N_22963,N_22841);
or U24809 (N_24809,N_22939,N_23452);
and U24810 (N_24810,N_22837,N_23463);
or U24811 (N_24811,N_22550,N_23490);
and U24812 (N_24812,N_23398,N_23447);
xnor U24813 (N_24813,N_23747,N_23236);
nor U24814 (N_24814,N_23114,N_22503);
xor U24815 (N_24815,N_22697,N_23580);
nor U24816 (N_24816,N_22963,N_23552);
xnor U24817 (N_24817,N_23213,N_23695);
and U24818 (N_24818,N_23478,N_23365);
xor U24819 (N_24819,N_22886,N_23093);
nand U24820 (N_24820,N_23195,N_22884);
nand U24821 (N_24821,N_23253,N_22597);
or U24822 (N_24822,N_23621,N_23492);
nand U24823 (N_24823,N_22539,N_22936);
nor U24824 (N_24824,N_23464,N_23605);
and U24825 (N_24825,N_23068,N_22745);
and U24826 (N_24826,N_22663,N_22711);
xor U24827 (N_24827,N_23095,N_23301);
nand U24828 (N_24828,N_23346,N_22867);
nand U24829 (N_24829,N_23467,N_23408);
xor U24830 (N_24830,N_22842,N_23277);
nor U24831 (N_24831,N_22931,N_22782);
nor U24832 (N_24832,N_22896,N_22914);
nor U24833 (N_24833,N_23022,N_23172);
or U24834 (N_24834,N_23072,N_23219);
nand U24835 (N_24835,N_22573,N_23226);
or U24836 (N_24836,N_22515,N_23712);
or U24837 (N_24837,N_22947,N_22846);
or U24838 (N_24838,N_23309,N_22838);
or U24839 (N_24839,N_22578,N_23613);
nor U24840 (N_24840,N_22667,N_22660);
xor U24841 (N_24841,N_22787,N_23641);
and U24842 (N_24842,N_22694,N_22950);
nor U24843 (N_24843,N_23625,N_23251);
and U24844 (N_24844,N_22792,N_22763);
xor U24845 (N_24845,N_23191,N_22765);
nand U24846 (N_24846,N_22855,N_23045);
or U24847 (N_24847,N_22770,N_22678);
nand U24848 (N_24848,N_23413,N_22721);
nand U24849 (N_24849,N_22627,N_22671);
nor U24850 (N_24850,N_23576,N_22785);
nand U24851 (N_24851,N_23597,N_23325);
or U24852 (N_24852,N_23626,N_23057);
nor U24853 (N_24853,N_23193,N_23460);
nor U24854 (N_24854,N_23253,N_23597);
nand U24855 (N_24855,N_23457,N_22742);
nor U24856 (N_24856,N_23000,N_22578);
xor U24857 (N_24857,N_23747,N_22894);
nand U24858 (N_24858,N_23154,N_22971);
and U24859 (N_24859,N_23192,N_22904);
and U24860 (N_24860,N_23157,N_23734);
nand U24861 (N_24861,N_22698,N_23718);
nor U24862 (N_24862,N_23000,N_23604);
xnor U24863 (N_24863,N_22864,N_23226);
xor U24864 (N_24864,N_23584,N_23287);
nand U24865 (N_24865,N_23715,N_23491);
or U24866 (N_24866,N_22516,N_22954);
and U24867 (N_24867,N_23733,N_23054);
nor U24868 (N_24868,N_23357,N_22782);
or U24869 (N_24869,N_22969,N_23559);
nor U24870 (N_24870,N_23528,N_23161);
or U24871 (N_24871,N_23214,N_22987);
and U24872 (N_24872,N_23685,N_22704);
or U24873 (N_24873,N_22799,N_22531);
or U24874 (N_24874,N_23083,N_23597);
xor U24875 (N_24875,N_23016,N_23033);
nor U24876 (N_24876,N_22986,N_23057);
nand U24877 (N_24877,N_23704,N_22975);
nand U24878 (N_24878,N_23350,N_22732);
or U24879 (N_24879,N_22506,N_23639);
nor U24880 (N_24880,N_23106,N_23441);
and U24881 (N_24881,N_23115,N_22505);
nor U24882 (N_24882,N_22694,N_22997);
xnor U24883 (N_24883,N_23474,N_22569);
or U24884 (N_24884,N_23426,N_23149);
xnor U24885 (N_24885,N_22742,N_22821);
and U24886 (N_24886,N_22984,N_22816);
or U24887 (N_24887,N_23273,N_23040);
and U24888 (N_24888,N_22624,N_23173);
or U24889 (N_24889,N_23495,N_22596);
and U24890 (N_24890,N_23263,N_23308);
nand U24891 (N_24891,N_23339,N_23013);
xnor U24892 (N_24892,N_22508,N_23315);
nand U24893 (N_24893,N_23680,N_23486);
or U24894 (N_24894,N_23237,N_23284);
or U24895 (N_24895,N_23091,N_23634);
or U24896 (N_24896,N_23714,N_22573);
nor U24897 (N_24897,N_23434,N_23667);
nor U24898 (N_24898,N_23083,N_23693);
nor U24899 (N_24899,N_23525,N_23679);
and U24900 (N_24900,N_23695,N_23421);
xnor U24901 (N_24901,N_23252,N_22883);
nand U24902 (N_24902,N_23723,N_22778);
nor U24903 (N_24903,N_23396,N_23063);
or U24904 (N_24904,N_22979,N_22914);
or U24905 (N_24905,N_23171,N_22863);
and U24906 (N_24906,N_22787,N_23695);
nand U24907 (N_24907,N_22576,N_23200);
xor U24908 (N_24908,N_22556,N_23281);
or U24909 (N_24909,N_23330,N_22758);
xor U24910 (N_24910,N_23182,N_23151);
nor U24911 (N_24911,N_23725,N_23691);
xor U24912 (N_24912,N_22512,N_22993);
or U24913 (N_24913,N_23693,N_22716);
and U24914 (N_24914,N_23454,N_22740);
or U24915 (N_24915,N_23000,N_23666);
nand U24916 (N_24916,N_22624,N_22591);
nor U24917 (N_24917,N_23130,N_23039);
or U24918 (N_24918,N_22581,N_23526);
or U24919 (N_24919,N_23251,N_23741);
nor U24920 (N_24920,N_23001,N_23375);
xor U24921 (N_24921,N_22952,N_22548);
nand U24922 (N_24922,N_22696,N_23360);
nand U24923 (N_24923,N_23277,N_23318);
nor U24924 (N_24924,N_23722,N_22848);
and U24925 (N_24925,N_22589,N_23112);
or U24926 (N_24926,N_22636,N_22977);
nand U24927 (N_24927,N_23314,N_23206);
xor U24928 (N_24928,N_23181,N_22906);
xnor U24929 (N_24929,N_23359,N_23163);
nor U24930 (N_24930,N_23586,N_23023);
nor U24931 (N_24931,N_22651,N_23238);
or U24932 (N_24932,N_23226,N_23258);
or U24933 (N_24933,N_23549,N_23069);
or U24934 (N_24934,N_22574,N_22862);
nand U24935 (N_24935,N_23690,N_22821);
xor U24936 (N_24936,N_23462,N_23727);
nand U24937 (N_24937,N_22630,N_23006);
and U24938 (N_24938,N_22808,N_23518);
xnor U24939 (N_24939,N_23182,N_23450);
and U24940 (N_24940,N_23587,N_22973);
and U24941 (N_24941,N_23087,N_23645);
and U24942 (N_24942,N_23557,N_23586);
or U24943 (N_24943,N_22900,N_23525);
nor U24944 (N_24944,N_22903,N_23301);
nor U24945 (N_24945,N_23261,N_23511);
and U24946 (N_24946,N_23036,N_23213);
and U24947 (N_24947,N_23181,N_23162);
and U24948 (N_24948,N_22988,N_23051);
nor U24949 (N_24949,N_22972,N_23323);
xor U24950 (N_24950,N_23594,N_22828);
and U24951 (N_24951,N_22944,N_23718);
nand U24952 (N_24952,N_23593,N_22895);
or U24953 (N_24953,N_22822,N_23739);
nor U24954 (N_24954,N_23579,N_22984);
xor U24955 (N_24955,N_23077,N_23235);
nor U24956 (N_24956,N_22540,N_22824);
or U24957 (N_24957,N_23008,N_23229);
or U24958 (N_24958,N_23496,N_22562);
or U24959 (N_24959,N_22860,N_23589);
xnor U24960 (N_24960,N_23169,N_23356);
or U24961 (N_24961,N_23645,N_22575);
xor U24962 (N_24962,N_23713,N_22602);
xor U24963 (N_24963,N_23521,N_23537);
nand U24964 (N_24964,N_23262,N_22711);
xor U24965 (N_24965,N_23110,N_23366);
nand U24966 (N_24966,N_23022,N_22832);
nand U24967 (N_24967,N_23621,N_23723);
and U24968 (N_24968,N_22951,N_23478);
nand U24969 (N_24969,N_22791,N_22916);
and U24970 (N_24970,N_23182,N_23212);
xnor U24971 (N_24971,N_22739,N_22788);
and U24972 (N_24972,N_23030,N_23022);
and U24973 (N_24973,N_22757,N_23495);
nand U24974 (N_24974,N_22558,N_23396);
nand U24975 (N_24975,N_22881,N_23728);
xor U24976 (N_24976,N_23710,N_23260);
nand U24977 (N_24977,N_22570,N_22580);
xnor U24978 (N_24978,N_22769,N_22841);
nand U24979 (N_24979,N_22808,N_22745);
nand U24980 (N_24980,N_23607,N_22892);
nand U24981 (N_24981,N_23404,N_23538);
and U24982 (N_24982,N_23070,N_23473);
xor U24983 (N_24983,N_22965,N_22883);
or U24984 (N_24984,N_23605,N_22560);
and U24985 (N_24985,N_22888,N_23385);
xor U24986 (N_24986,N_23329,N_22795);
and U24987 (N_24987,N_22808,N_23547);
or U24988 (N_24988,N_23382,N_23536);
xor U24989 (N_24989,N_22512,N_22513);
and U24990 (N_24990,N_22664,N_22837);
nand U24991 (N_24991,N_23653,N_23362);
and U24992 (N_24992,N_23679,N_23159);
nor U24993 (N_24993,N_23117,N_22704);
xor U24994 (N_24994,N_22713,N_23444);
or U24995 (N_24995,N_23055,N_23627);
or U24996 (N_24996,N_23711,N_22950);
and U24997 (N_24997,N_23115,N_22724);
nand U24998 (N_24998,N_23276,N_22577);
or U24999 (N_24999,N_23316,N_23094);
nor UO_0 (O_0,N_24221,N_24093);
nand UO_1 (O_1,N_23980,N_24012);
nand UO_2 (O_2,N_24806,N_24094);
nor UO_3 (O_3,N_24827,N_24575);
or UO_4 (O_4,N_24549,N_24264);
or UO_5 (O_5,N_24725,N_24112);
xnor UO_6 (O_6,N_24638,N_24371);
and UO_7 (O_7,N_24572,N_23785);
xor UO_8 (O_8,N_24483,N_23811);
nand UO_9 (O_9,N_24916,N_24228);
or UO_10 (O_10,N_24266,N_24678);
nor UO_11 (O_11,N_24867,N_24988);
nor UO_12 (O_12,N_24679,N_24664);
xnor UO_13 (O_13,N_24615,N_23891);
or UO_14 (O_14,N_23775,N_24895);
xnor UO_15 (O_15,N_24713,N_24558);
xnor UO_16 (O_16,N_23765,N_24170);
nand UO_17 (O_17,N_23834,N_24121);
nor UO_18 (O_18,N_24577,N_24402);
nor UO_19 (O_19,N_24650,N_24687);
nor UO_20 (O_20,N_24798,N_24835);
nand UO_21 (O_21,N_23977,N_24858);
xor UO_22 (O_22,N_24699,N_24801);
or UO_23 (O_23,N_24669,N_24810);
nand UO_24 (O_24,N_24846,N_24611);
nand UO_25 (O_25,N_24028,N_24641);
nor UO_26 (O_26,N_24367,N_23781);
nand UO_27 (O_27,N_23852,N_23955);
and UO_28 (O_28,N_24720,N_24978);
nand UO_29 (O_29,N_24844,N_24658);
nand UO_30 (O_30,N_24301,N_24239);
nor UO_31 (O_31,N_24491,N_24388);
nor UO_32 (O_32,N_24532,N_23944);
and UO_33 (O_33,N_24114,N_24142);
nand UO_34 (O_34,N_23936,N_24585);
and UO_35 (O_35,N_24697,N_24994);
or UO_36 (O_36,N_24597,N_24890);
and UO_37 (O_37,N_24152,N_24771);
or UO_38 (O_38,N_24631,N_24764);
or UO_39 (O_39,N_24602,N_24681);
xnor UO_40 (O_40,N_24352,N_23880);
or UO_41 (O_41,N_24546,N_24870);
and UO_42 (O_42,N_23892,N_24282);
or UO_43 (O_43,N_24928,N_24325);
nor UO_44 (O_44,N_24969,N_24022);
xor UO_45 (O_45,N_24355,N_23905);
and UO_46 (O_46,N_24131,N_23992);
xnor UO_47 (O_47,N_24195,N_24876);
xor UO_48 (O_48,N_24494,N_24904);
and UO_49 (O_49,N_23913,N_24097);
nand UO_50 (O_50,N_24811,N_24020);
nor UO_51 (O_51,N_24008,N_23832);
and UO_52 (O_52,N_24832,N_24898);
nor UO_53 (O_53,N_24481,N_24484);
xnor UO_54 (O_54,N_24790,N_24618);
and UO_55 (O_55,N_24182,N_24884);
xnor UO_56 (O_56,N_24622,N_23814);
xor UO_57 (O_57,N_24940,N_24249);
and UO_58 (O_58,N_24099,N_24290);
nand UO_59 (O_59,N_24214,N_24854);
and UO_60 (O_60,N_24981,N_24018);
or UO_61 (O_61,N_23789,N_24626);
and UO_62 (O_62,N_23750,N_24710);
nor UO_63 (O_63,N_24410,N_23876);
and UO_64 (O_64,N_24750,N_24505);
xnor UO_65 (O_65,N_23879,N_24184);
nor UO_66 (O_66,N_24507,N_24468);
and UO_67 (O_67,N_24158,N_24574);
xor UO_68 (O_68,N_24077,N_24103);
or UO_69 (O_69,N_24747,N_24145);
nand UO_70 (O_70,N_23760,N_23885);
and UO_71 (O_71,N_24005,N_24021);
or UO_72 (O_72,N_23886,N_24144);
and UO_73 (O_73,N_24691,N_24236);
nor UO_74 (O_74,N_23815,N_24438);
xor UO_75 (O_75,N_23889,N_24939);
xnor UO_76 (O_76,N_23822,N_24224);
nor UO_77 (O_77,N_24253,N_24983);
or UO_78 (O_78,N_24035,N_24081);
xor UO_79 (O_79,N_24490,N_24902);
xnor UO_80 (O_80,N_24318,N_24670);
xor UO_81 (O_81,N_23973,N_23870);
nand UO_82 (O_82,N_24361,N_24384);
nand UO_83 (O_83,N_23954,N_23989);
nand UO_84 (O_84,N_24124,N_23873);
and UO_85 (O_85,N_24760,N_24470);
nor UO_86 (O_86,N_24376,N_24275);
nor UO_87 (O_87,N_23917,N_24113);
and UO_88 (O_88,N_23969,N_23847);
nor UO_89 (O_89,N_24584,N_24444);
or UO_90 (O_90,N_23755,N_24581);
nand UO_91 (O_91,N_24339,N_24565);
or UO_92 (O_92,N_24996,N_24905);
nand UO_93 (O_93,N_23807,N_24377);
xnor UO_94 (O_94,N_24954,N_24447);
nand UO_95 (O_95,N_24054,N_23831);
nand UO_96 (O_96,N_24536,N_24774);
nor UO_97 (O_97,N_24989,N_24218);
or UO_98 (O_98,N_24949,N_24831);
nand UO_99 (O_99,N_24010,N_23777);
or UO_100 (O_100,N_24515,N_24425);
nor UO_101 (O_101,N_24231,N_24960);
nor UO_102 (O_102,N_24467,N_24935);
and UO_103 (O_103,N_24098,N_24823);
or UO_104 (O_104,N_23940,N_24766);
and UO_105 (O_105,N_23768,N_24837);
and UO_106 (O_106,N_23896,N_24030);
and UO_107 (O_107,N_24952,N_24364);
xnor UO_108 (O_108,N_24762,N_23862);
nand UO_109 (O_109,N_24213,N_24399);
and UO_110 (O_110,N_24134,N_24965);
and UO_111 (O_111,N_24219,N_24987);
or UO_112 (O_112,N_24476,N_24143);
and UO_113 (O_113,N_24270,N_23962);
and UO_114 (O_114,N_24118,N_24633);
and UO_115 (O_115,N_24729,N_24707);
nand UO_116 (O_116,N_23829,N_24544);
xnor UO_117 (O_117,N_24921,N_24526);
nand UO_118 (O_118,N_24997,N_23872);
nor UO_119 (O_119,N_24272,N_24652);
and UO_120 (O_120,N_24246,N_24179);
nor UO_121 (O_121,N_24995,N_24576);
or UO_122 (O_122,N_23945,N_24892);
or UO_123 (O_123,N_24086,N_24464);
xor UO_124 (O_124,N_24688,N_24976);
nor UO_125 (O_125,N_23849,N_24190);
xnor UO_126 (O_126,N_24812,N_23758);
or UO_127 (O_127,N_24853,N_24451);
and UO_128 (O_128,N_23900,N_24485);
nor UO_129 (O_129,N_24802,N_24692);
nand UO_130 (O_130,N_24937,N_24535);
nor UO_131 (O_131,N_23937,N_24828);
or UO_132 (O_132,N_24662,N_24409);
and UO_133 (O_133,N_24059,N_24958);
or UO_134 (O_134,N_24871,N_24616);
or UO_135 (O_135,N_24672,N_23909);
nor UO_136 (O_136,N_24242,N_24323);
nor UO_137 (O_137,N_24724,N_23804);
nor UO_138 (O_138,N_24529,N_24805);
nand UO_139 (O_139,N_24786,N_24265);
or UO_140 (O_140,N_24941,N_23828);
and UO_141 (O_141,N_24233,N_24357);
nor UO_142 (O_142,N_24522,N_24078);
nor UO_143 (O_143,N_23767,N_24075);
nor UO_144 (O_144,N_24421,N_24962);
nor UO_145 (O_145,N_24732,N_23802);
and UO_146 (O_146,N_24723,N_24082);
and UO_147 (O_147,N_23761,N_23943);
or UO_148 (O_148,N_24792,N_24189);
nor UO_149 (O_149,N_24552,N_24226);
xor UO_150 (O_150,N_24069,N_24503);
and UO_151 (O_151,N_24406,N_24986);
and UO_152 (O_152,N_24469,N_24934);
nor UO_153 (O_153,N_24668,N_24701);
nor UO_154 (O_154,N_24684,N_24188);
or UO_155 (O_155,N_24562,N_24915);
nand UO_156 (O_156,N_24795,N_24130);
or UO_157 (O_157,N_24966,N_24207);
nor UO_158 (O_158,N_24051,N_24480);
and UO_159 (O_159,N_23827,N_23839);
xor UO_160 (O_160,N_24197,N_23867);
and UO_161 (O_161,N_24770,N_24560);
nand UO_162 (O_162,N_24778,N_24177);
and UO_163 (O_163,N_23919,N_24926);
nor UO_164 (O_164,N_24977,N_24959);
and UO_165 (O_165,N_24389,N_24003);
or UO_166 (O_166,N_24337,N_23887);
nor UO_167 (O_167,N_23800,N_24610);
or UO_168 (O_168,N_24527,N_24340);
or UO_169 (O_169,N_24247,N_24769);
and UO_170 (O_170,N_24925,N_24164);
and UO_171 (O_171,N_24818,N_23841);
xor UO_172 (O_172,N_24841,N_23949);
and UO_173 (O_173,N_24859,N_23821);
nor UO_174 (O_174,N_24454,N_24386);
nor UO_175 (O_175,N_24079,N_23899);
xnor UO_176 (O_176,N_24504,N_24525);
xnor UO_177 (O_177,N_24624,N_23995);
nand UO_178 (O_178,N_24437,N_24726);
and UO_179 (O_179,N_24794,N_23825);
or UO_180 (O_180,N_24807,N_24412);
xor UO_181 (O_181,N_24336,N_24160);
and UO_182 (O_182,N_24609,N_23788);
nor UO_183 (O_183,N_23942,N_24696);
or UO_184 (O_184,N_24788,N_23983);
or UO_185 (O_185,N_24605,N_24136);
nand UO_186 (O_186,N_24394,N_24791);
xnor UO_187 (O_187,N_24924,N_24666);
xnor UO_188 (O_188,N_24580,N_24975);
and UO_189 (O_189,N_24300,N_24127);
xor UO_190 (O_190,N_24324,N_24055);
nand UO_191 (O_191,N_24209,N_24024);
or UO_192 (O_192,N_24070,N_24327);
nand UO_193 (O_193,N_24334,N_24542);
nor UO_194 (O_194,N_24023,N_24284);
and UO_195 (O_195,N_23911,N_24745);
nor UO_196 (O_196,N_24053,N_24202);
and UO_197 (O_197,N_24196,N_24872);
or UO_198 (O_198,N_24563,N_24200);
xnor UO_199 (O_199,N_24653,N_24155);
nor UO_200 (O_200,N_24319,N_24091);
nand UO_201 (O_201,N_23810,N_24919);
xor UO_202 (O_202,N_23966,N_23986);
xnor UO_203 (O_203,N_24623,N_23895);
xor UO_204 (O_204,N_23897,N_24401);
xnor UO_205 (O_205,N_24755,N_24080);
xnor UO_206 (O_206,N_24248,N_24799);
and UO_207 (O_207,N_24839,N_23857);
and UO_208 (O_208,N_24632,N_23791);
and UO_209 (O_209,N_24974,N_24273);
and UO_210 (O_210,N_24101,N_24946);
xnor UO_211 (O_211,N_24932,N_24443);
nand UO_212 (O_212,N_24417,N_24117);
and UO_213 (O_213,N_24474,N_24048);
nand UO_214 (O_214,N_24243,N_23948);
and UO_215 (O_215,N_24822,N_24141);
xnor UO_216 (O_216,N_23923,N_24911);
nor UO_217 (O_217,N_24353,N_24917);
nor UO_218 (O_218,N_24088,N_24703);
and UO_219 (O_219,N_24660,N_23799);
or UO_220 (O_220,N_24104,N_24220);
nand UO_221 (O_221,N_23796,N_23903);
and UO_222 (O_222,N_24448,N_24592);
xor UO_223 (O_223,N_23812,N_24608);
nand UO_224 (O_224,N_24201,N_24735);
nor UO_225 (O_225,N_24604,N_24737);
xnor UO_226 (O_226,N_23907,N_24797);
xnor UO_227 (O_227,N_24711,N_24899);
nor UO_228 (O_228,N_24475,N_23865);
xnor UO_229 (O_229,N_23974,N_24174);
nor UO_230 (O_230,N_24889,N_24132);
xnor UO_231 (O_231,N_24217,N_24716);
nand UO_232 (O_232,N_24739,N_24199);
or UO_233 (O_233,N_24756,N_23787);
and UO_234 (O_234,N_24524,N_24366);
xor UO_235 (O_235,N_24495,N_24175);
nand UO_236 (O_236,N_24619,N_24682);
xnor UO_237 (O_237,N_23939,N_24385);
nor UO_238 (O_238,N_24204,N_24167);
nor UO_239 (O_239,N_24316,N_24759);
nor UO_240 (O_240,N_24335,N_24800);
xor UO_241 (O_241,N_24803,N_24543);
or UO_242 (O_242,N_23764,N_24383);
xor UO_243 (O_243,N_24076,N_24740);
nor UO_244 (O_244,N_24087,N_23931);
and UO_245 (O_245,N_24721,N_23993);
xor UO_246 (O_246,N_24489,N_24743);
nand UO_247 (O_247,N_24773,N_24044);
or UO_248 (O_248,N_24727,N_24450);
xor UO_249 (O_249,N_24063,N_24000);
xor UO_250 (O_250,N_24520,N_24550);
or UO_251 (O_251,N_24135,N_24478);
nor UO_252 (O_252,N_24493,N_24897);
nand UO_253 (O_253,N_24458,N_24257);
nor UO_254 (O_254,N_24040,N_24646);
nand UO_255 (O_255,N_24110,N_24856);
xnor UO_256 (O_256,N_23902,N_24173);
xor UO_257 (O_257,N_24434,N_23926);
xnor UO_258 (O_258,N_24255,N_24556);
nand UO_259 (O_259,N_23778,N_23972);
xnor UO_260 (O_260,N_24838,N_23874);
and UO_261 (O_261,N_24582,N_24185);
or UO_262 (O_262,N_24782,N_24322);
xnor UO_263 (O_263,N_24548,N_23774);
nand UO_264 (O_264,N_24569,N_23990);
xnor UO_265 (O_265,N_24751,N_24393);
nand UO_266 (O_266,N_24930,N_24479);
nor UO_267 (O_267,N_23752,N_23965);
nor UO_268 (O_268,N_24288,N_24815);
and UO_269 (O_269,N_24629,N_24279);
or UO_270 (O_270,N_24900,N_24901);
nor UO_271 (O_271,N_24292,N_24100);
and UO_272 (O_272,N_23784,N_23920);
nor UO_273 (O_273,N_24089,N_24878);
or UO_274 (O_274,N_24061,N_24886);
and UO_275 (O_275,N_23753,N_24305);
nand UO_276 (O_276,N_23845,N_23918);
and UO_277 (O_277,N_24208,N_24639);
xnor UO_278 (O_278,N_24068,N_23816);
or UO_279 (O_279,N_24861,N_24980);
or UO_280 (O_280,N_24095,N_23871);
or UO_281 (O_281,N_24547,N_24763);
xnor UO_282 (O_282,N_24765,N_24212);
and UO_283 (O_283,N_23757,N_24165);
or UO_284 (O_284,N_24445,N_24768);
or UO_285 (O_285,N_24293,N_24833);
nor UO_286 (O_286,N_23754,N_24378);
xor UO_287 (O_287,N_24950,N_24809);
xnor UO_288 (O_288,N_24671,N_24187);
and UO_289 (O_289,N_24391,N_24936);
nor UO_290 (O_290,N_23859,N_24488);
nor UO_291 (O_291,N_23792,N_24056);
and UO_292 (O_292,N_23877,N_24403);
nor UO_293 (O_293,N_24758,N_24487);
and UO_294 (O_294,N_24348,N_24347);
and UO_295 (O_295,N_24627,N_23964);
xnor UO_296 (O_296,N_24566,N_24883);
and UO_297 (O_297,N_23963,N_24829);
or UO_298 (O_298,N_24230,N_24382);
xnor UO_299 (O_299,N_24304,N_23795);
and UO_300 (O_300,N_23952,N_24256);
and UO_301 (O_301,N_23894,N_24037);
or UO_302 (O_302,N_24840,N_24085);
nand UO_303 (O_303,N_23836,N_24090);
or UO_304 (O_304,N_24129,N_23971);
nor UO_305 (O_305,N_24302,N_24343);
nor UO_306 (O_306,N_24423,N_24455);
xor UO_307 (O_307,N_24634,N_24492);
xor UO_308 (O_308,N_24426,N_24011);
or UO_309 (O_309,N_23884,N_23994);
nand UO_310 (O_310,N_24531,N_24240);
nor UO_311 (O_311,N_23869,N_23898);
nor UO_312 (O_312,N_24241,N_23801);
nor UO_313 (O_313,N_24712,N_24731);
or UO_314 (O_314,N_24122,N_24499);
or UO_315 (O_315,N_24049,N_24599);
nand UO_316 (O_316,N_24014,N_24990);
nand UO_317 (O_317,N_24392,N_23805);
nand UO_318 (O_318,N_24414,N_23766);
or UO_319 (O_319,N_24295,N_24320);
and UO_320 (O_320,N_24294,N_24636);
or UO_321 (O_321,N_24850,N_24001);
nor UO_322 (O_322,N_24612,N_24595);
and UO_323 (O_323,N_24780,N_24864);
nand UO_324 (O_324,N_24262,N_24620);
and UO_325 (O_325,N_24693,N_24172);
nand UO_326 (O_326,N_24258,N_24181);
or UO_327 (O_327,N_24530,N_24553);
xor UO_328 (O_328,N_23863,N_24757);
xnor UO_329 (O_329,N_23979,N_24073);
nand UO_330 (O_330,N_24123,N_23916);
nor UO_331 (O_331,N_24004,N_24910);
nand UO_332 (O_332,N_23762,N_23947);
xnor UO_333 (O_333,N_23881,N_24052);
nand UO_334 (O_334,N_23958,N_24108);
xnor UO_335 (O_335,N_24276,N_23912);
nand UO_336 (O_336,N_24852,N_24642);
or UO_337 (O_337,N_24358,N_24914);
xor UO_338 (O_338,N_24706,N_24111);
nand UO_339 (O_339,N_24374,N_24545);
xor UO_340 (O_340,N_24999,N_24497);
xor UO_341 (O_341,N_23860,N_23783);
nor UO_342 (O_342,N_24036,N_24120);
or UO_343 (O_343,N_24453,N_24923);
nor UO_344 (O_344,N_24779,N_23826);
or UO_345 (O_345,N_24150,N_23813);
and UO_346 (O_346,N_24222,N_24362);
nand UO_347 (O_347,N_23961,N_24907);
or UO_348 (O_348,N_24533,N_24863);
nor UO_349 (O_349,N_23835,N_24722);
xnor UO_350 (O_350,N_23866,N_24156);
xor UO_351 (O_351,N_24689,N_24537);
xor UO_352 (O_352,N_24065,N_23779);
and UO_353 (O_353,N_24311,N_23803);
nand UO_354 (O_354,N_24083,N_24128);
nor UO_355 (O_355,N_24702,N_23893);
xnor UO_356 (O_356,N_23953,N_24342);
nand UO_357 (O_357,N_24661,N_24808);
nand UO_358 (O_358,N_24953,N_24951);
nor UO_359 (O_359,N_24397,N_24793);
or UO_360 (O_360,N_24704,N_24269);
or UO_361 (O_361,N_24223,N_24881);
or UO_362 (O_362,N_24486,N_23794);
nor UO_363 (O_363,N_24422,N_24888);
nor UO_364 (O_364,N_24673,N_24598);
and UO_365 (O_365,N_24328,N_24695);
xnor UO_366 (O_366,N_24513,N_23858);
and UO_367 (O_367,N_24922,N_24587);
xor UO_368 (O_368,N_23987,N_24459);
and UO_369 (O_369,N_24578,N_24719);
or UO_370 (O_370,N_24521,N_24819);
or UO_371 (O_371,N_24506,N_24814);
nand UO_372 (O_372,N_24590,N_24643);
or UO_373 (O_373,N_24153,N_24432);
nor UO_374 (O_374,N_24429,N_23956);
and UO_375 (O_375,N_24215,N_24512);
xor UO_376 (O_376,N_24390,N_24178);
nand UO_377 (O_377,N_24903,N_24875);
nor UO_378 (O_378,N_24216,N_24657);
nor UO_379 (O_379,N_24440,N_24171);
and UO_380 (O_380,N_23856,N_24970);
and UO_381 (O_381,N_24163,N_24009);
or UO_382 (O_382,N_24945,N_24194);
or UO_383 (O_383,N_24462,N_24349);
and UO_384 (O_384,N_24787,N_24109);
xnor UO_385 (O_385,N_24395,N_24205);
and UO_386 (O_386,N_24733,N_24998);
or UO_387 (O_387,N_24596,N_24250);
and UO_388 (O_388,N_24331,N_24449);
or UO_389 (O_389,N_24857,N_24730);
nand UO_390 (O_390,N_24192,N_24271);
nand UO_391 (O_391,N_24571,N_24614);
and UO_392 (O_392,N_24717,N_24237);
or UO_393 (O_393,N_24379,N_23854);
and UO_394 (O_394,N_24728,N_24849);
or UO_395 (O_395,N_23967,N_24594);
nor UO_396 (O_396,N_24238,N_24140);
nor UO_397 (O_397,N_24541,N_24415);
nor UO_398 (O_398,N_24784,N_24982);
or UO_399 (O_399,N_24452,N_24625);
nand UO_400 (O_400,N_24084,N_24516);
and UO_401 (O_401,N_23759,N_24166);
nor UO_402 (O_402,N_24232,N_24748);
and UO_403 (O_403,N_24551,N_24607);
nand UO_404 (O_404,N_24909,N_24789);
nor UO_405 (O_405,N_23855,N_24956);
and UO_406 (O_406,N_24830,N_24058);
nor UO_407 (O_407,N_23818,N_24064);
nand UO_408 (O_408,N_24102,N_24312);
nor UO_409 (O_409,N_24498,N_24979);
and UO_410 (O_410,N_24938,N_24225);
or UO_411 (O_411,N_24873,N_24777);
nand UO_412 (O_412,N_24333,N_24655);
xor UO_413 (O_413,N_24685,N_24973);
xnor UO_414 (O_414,N_24927,N_24433);
xor UO_415 (O_415,N_24033,N_24738);
nor UO_416 (O_416,N_24473,N_23808);
xnor UO_417 (O_417,N_23751,N_23793);
or UO_418 (O_418,N_24540,N_24775);
xnor UO_419 (O_419,N_24570,N_23850);
and UO_420 (O_420,N_24420,N_24583);
nand UO_421 (O_421,N_24435,N_24557);
and UO_422 (O_422,N_24894,N_24038);
and UO_423 (O_423,N_24006,N_24330);
or UO_424 (O_424,N_24176,N_24539);
xnor UO_425 (O_425,N_23819,N_24427);
nor UO_426 (O_426,N_23846,N_24880);
nor UO_427 (O_427,N_24635,N_24025);
or UO_428 (O_428,N_24317,N_24676);
xnor UO_429 (O_429,N_24326,N_23776);
and UO_430 (O_430,N_24050,N_24193);
nor UO_431 (O_431,N_24133,N_24667);
and UO_432 (O_432,N_24026,N_24621);
nor UO_433 (O_433,N_24229,N_24509);
nand UO_434 (O_434,N_24523,N_24306);
nor UO_435 (O_435,N_24408,N_24561);
xor UO_436 (O_436,N_24183,N_23985);
and UO_437 (O_437,N_23960,N_24442);
xnor UO_438 (O_438,N_23769,N_23934);
and UO_439 (O_439,N_24428,N_24254);
or UO_440 (O_440,N_24508,N_24862);
and UO_441 (O_441,N_24252,N_23763);
nor UO_442 (O_442,N_24466,N_24105);
and UO_443 (O_443,N_24234,N_24308);
nand UO_444 (O_444,N_24119,N_24929);
nand UO_445 (O_445,N_23838,N_24041);
nor UO_446 (O_446,N_24511,N_24984);
nand UO_447 (O_447,N_24744,N_23817);
xnor UO_448 (O_448,N_24694,N_24148);
nand UO_449 (O_449,N_24341,N_24971);
nand UO_450 (O_450,N_24617,N_23924);
nor UO_451 (O_451,N_24869,N_24502);
or UO_452 (O_452,N_23842,N_23997);
xnor UO_453 (O_453,N_24912,N_23976);
nand UO_454 (O_454,N_24820,N_23782);
and UO_455 (O_455,N_24244,N_24715);
and UO_456 (O_456,N_24972,N_24821);
and UO_457 (O_457,N_24675,N_24307);
nor UO_458 (O_458,N_23998,N_24465);
xnor UO_459 (O_459,N_23908,N_24845);
nor UO_460 (O_460,N_24138,N_24877);
nand UO_461 (O_461,N_24783,N_24601);
nor UO_462 (O_462,N_24968,N_24992);
xor UO_463 (O_463,N_24168,N_24588);
and UO_464 (O_464,N_24332,N_24879);
xnor UO_465 (O_465,N_24329,N_24380);
and UO_466 (O_466,N_24203,N_24640);
nor UO_467 (O_467,N_24297,N_23991);
or UO_468 (O_468,N_24648,N_23843);
nor UO_469 (O_469,N_23786,N_24649);
nor UO_470 (O_470,N_24781,N_24991);
nand UO_471 (O_471,N_23833,N_24709);
or UO_472 (O_472,N_24874,N_24344);
nor UO_473 (O_473,N_24017,N_23820);
nand UO_474 (O_474,N_23910,N_24263);
or UO_475 (O_475,N_24683,N_24651);
nor UO_476 (O_476,N_23844,N_24834);
and UO_477 (O_477,N_24211,N_24125);
nor UO_478 (O_478,N_24235,N_24031);
nand UO_479 (O_479,N_23780,N_24198);
nor UO_480 (O_480,N_24045,N_24955);
nand UO_481 (O_481,N_23929,N_23906);
nand UO_482 (O_482,N_24993,N_24287);
nor UO_483 (O_483,N_24002,N_24538);
and UO_484 (O_484,N_24137,N_24591);
nand UO_485 (O_485,N_24314,N_24510);
or UO_486 (O_486,N_24149,N_23951);
or UO_487 (O_487,N_24375,N_23875);
nor UO_488 (O_488,N_24776,N_24500);
or UO_489 (O_489,N_24654,N_24013);
or UO_490 (O_490,N_24372,N_24816);
xnor UO_491 (O_491,N_24370,N_24644);
nor UO_492 (O_492,N_24043,N_24659);
nand UO_493 (O_493,N_24436,N_24942);
or UO_494 (O_494,N_23950,N_23837);
xnor UO_495 (O_495,N_24274,N_23888);
nand UO_496 (O_496,N_24461,N_24554);
nand UO_497 (O_497,N_24047,N_24107);
or UO_498 (O_498,N_24457,N_24456);
or UO_499 (O_499,N_24072,N_24472);
xnor UO_500 (O_500,N_24303,N_24291);
nand UO_501 (O_501,N_23982,N_24656);
xor UO_502 (O_502,N_24865,N_24847);
xor UO_503 (O_503,N_24191,N_24754);
xor UO_504 (O_504,N_23790,N_24411);
or UO_505 (O_505,N_24964,N_24586);
xor UO_506 (O_506,N_24268,N_24365);
xnor UO_507 (O_507,N_23959,N_24825);
nor UO_508 (O_508,N_23864,N_24589);
and UO_509 (O_509,N_23984,N_24753);
and UO_510 (O_510,N_24039,N_23851);
nor UO_511 (O_511,N_24154,N_23922);
and UO_512 (O_512,N_24891,N_24804);
xor UO_513 (O_513,N_24032,N_24439);
nand UO_514 (O_514,N_24407,N_23930);
nand UO_515 (O_515,N_23914,N_24663);
and UO_516 (O_516,N_24933,N_24882);
and UO_517 (O_517,N_23770,N_24680);
and UO_518 (O_518,N_24665,N_24848);
or UO_519 (O_519,N_24034,N_23809);
and UO_520 (O_520,N_23806,N_24593);
nand UO_521 (O_521,N_24564,N_24967);
or UO_522 (O_522,N_23878,N_24700);
nand UO_523 (O_523,N_24360,N_24742);
nand UO_524 (O_524,N_23798,N_24315);
nand UO_525 (O_525,N_24363,N_24029);
nand UO_526 (O_526,N_24943,N_24431);
xnor UO_527 (O_527,N_23848,N_24368);
or UO_528 (O_528,N_24046,N_24906);
nor UO_529 (O_529,N_24772,N_24947);
xnor UO_530 (O_530,N_23773,N_24151);
nor UO_531 (O_531,N_23756,N_24734);
xor UO_532 (O_532,N_24245,N_24842);
and UO_533 (O_533,N_24060,N_24637);
and UO_534 (O_534,N_24813,N_24855);
nand UO_535 (O_535,N_24277,N_23823);
xnor UO_536 (O_536,N_23861,N_23938);
or UO_537 (O_537,N_24309,N_23824);
and UO_538 (O_538,N_24096,N_23840);
or UO_539 (O_539,N_24517,N_24918);
nor UO_540 (O_540,N_24957,N_24396);
and UO_541 (O_541,N_24603,N_23890);
xor UO_542 (O_542,N_23933,N_24161);
and UO_543 (O_543,N_23797,N_24345);
xnor UO_544 (O_544,N_24299,N_24628);
nor UO_545 (O_545,N_24868,N_24413);
xor UO_546 (O_546,N_24338,N_24369);
or UO_547 (O_547,N_23771,N_24206);
xnor UO_548 (O_548,N_24824,N_24027);
or UO_549 (O_549,N_24162,N_23996);
nor UO_550 (O_550,N_24416,N_24836);
nor UO_551 (O_551,N_24893,N_23830);
xor UO_552 (O_552,N_24139,N_23883);
or UO_553 (O_553,N_24630,N_24126);
and UO_554 (O_554,N_24767,N_24645);
and UO_555 (O_555,N_24157,N_24261);
xor UO_556 (O_556,N_23901,N_23925);
and UO_557 (O_557,N_24746,N_24573);
and UO_558 (O_558,N_24920,N_24259);
nand UO_559 (O_559,N_24647,N_24400);
xor UO_560 (O_560,N_24346,N_23868);
or UO_561 (O_561,N_24686,N_24528);
or UO_562 (O_562,N_24948,N_23981);
xnor UO_563 (O_563,N_24534,N_23853);
and UO_564 (O_564,N_24356,N_23935);
or UO_565 (O_565,N_24718,N_24698);
nand UO_566 (O_566,N_23968,N_24736);
nor UO_567 (O_567,N_24714,N_24600);
xnor UO_568 (O_568,N_24146,N_23946);
and UO_569 (O_569,N_24321,N_24514);
nor UO_570 (O_570,N_23970,N_24286);
nand UO_571 (O_571,N_24613,N_24042);
or UO_572 (O_572,N_24705,N_24016);
nand UO_573 (O_573,N_24741,N_24579);
and UO_574 (O_574,N_24885,N_24285);
nand UO_575 (O_575,N_24354,N_23988);
and UO_576 (O_576,N_24460,N_24398);
xor UO_577 (O_577,N_23772,N_23882);
xor UO_578 (O_578,N_24278,N_23904);
nand UO_579 (O_579,N_24186,N_23915);
or UO_580 (O_580,N_24674,N_24430);
nor UO_581 (O_581,N_24985,N_23927);
nand UO_582 (O_582,N_24260,N_24761);
nor UO_583 (O_583,N_24866,N_24463);
xor UO_584 (O_584,N_24350,N_24913);
and UO_585 (O_585,N_23978,N_24057);
nand UO_586 (O_586,N_24471,N_24351);
and UO_587 (O_587,N_24067,N_24071);
and UO_588 (O_588,N_24298,N_24296);
nor UO_589 (O_589,N_24843,N_24251);
or UO_590 (O_590,N_24169,N_24961);
or UO_591 (O_591,N_24310,N_24568);
or UO_592 (O_592,N_24281,N_24690);
or UO_593 (O_593,N_24405,N_24373);
and UO_594 (O_594,N_24501,N_24147);
xnor UO_595 (O_595,N_24092,N_24931);
nand UO_596 (O_596,N_24555,N_24062);
xnor UO_597 (O_597,N_24606,N_24404);
or UO_598 (O_598,N_24210,N_24441);
xor UO_599 (O_599,N_24785,N_24908);
nand UO_600 (O_600,N_24860,N_24019);
xnor UO_601 (O_601,N_23928,N_24267);
nand UO_602 (O_602,N_24159,N_24944);
nand UO_603 (O_603,N_24708,N_24896);
and UO_604 (O_604,N_24283,N_24007);
nor UO_605 (O_605,N_24116,N_24749);
and UO_606 (O_606,N_24963,N_24851);
nand UO_607 (O_607,N_24677,N_24496);
and UO_608 (O_608,N_24518,N_23975);
nand UO_609 (O_609,N_23957,N_24387);
xnor UO_610 (O_610,N_24752,N_24559);
or UO_611 (O_611,N_23932,N_24280);
nand UO_612 (O_612,N_24313,N_24817);
or UO_613 (O_613,N_24359,N_24227);
or UO_614 (O_614,N_23921,N_23999);
xnor UO_615 (O_615,N_24826,N_23941);
xnor UO_616 (O_616,N_24289,N_24519);
nor UO_617 (O_617,N_24446,N_24015);
or UO_618 (O_618,N_24381,N_24567);
nor UO_619 (O_619,N_24074,N_24115);
or UO_620 (O_620,N_24796,N_24180);
nand UO_621 (O_621,N_24482,N_24424);
xnor UO_622 (O_622,N_24106,N_24887);
or UO_623 (O_623,N_24477,N_24418);
nand UO_624 (O_624,N_24066,N_24419);
xnor UO_625 (O_625,N_24469,N_24100);
nor UO_626 (O_626,N_24909,N_24560);
xnor UO_627 (O_627,N_24191,N_23974);
xor UO_628 (O_628,N_23909,N_24749);
xor UO_629 (O_629,N_24618,N_23899);
xnor UO_630 (O_630,N_24009,N_24253);
nor UO_631 (O_631,N_24065,N_24001);
or UO_632 (O_632,N_24225,N_23997);
xor UO_633 (O_633,N_24564,N_23992);
nor UO_634 (O_634,N_23871,N_23968);
or UO_635 (O_635,N_24527,N_24600);
and UO_636 (O_636,N_24287,N_24678);
nor UO_637 (O_637,N_24595,N_24150);
nor UO_638 (O_638,N_24745,N_23941);
nor UO_639 (O_639,N_24139,N_24304);
xor UO_640 (O_640,N_24572,N_24146);
nand UO_641 (O_641,N_24606,N_24240);
or UO_642 (O_642,N_24791,N_24671);
nand UO_643 (O_643,N_24761,N_24844);
or UO_644 (O_644,N_24271,N_24450);
and UO_645 (O_645,N_24303,N_24156);
and UO_646 (O_646,N_24386,N_24150);
or UO_647 (O_647,N_24841,N_24996);
and UO_648 (O_648,N_24823,N_24423);
and UO_649 (O_649,N_24220,N_23776);
and UO_650 (O_650,N_24503,N_24907);
nor UO_651 (O_651,N_24332,N_24369);
or UO_652 (O_652,N_24797,N_23805);
nand UO_653 (O_653,N_24358,N_24141);
xor UO_654 (O_654,N_24419,N_24617);
and UO_655 (O_655,N_24514,N_24375);
and UO_656 (O_656,N_24386,N_24868);
or UO_657 (O_657,N_24449,N_23870);
nand UO_658 (O_658,N_24647,N_24681);
or UO_659 (O_659,N_24912,N_23890);
or UO_660 (O_660,N_24394,N_23946);
or UO_661 (O_661,N_24518,N_24354);
and UO_662 (O_662,N_24643,N_24982);
and UO_663 (O_663,N_24759,N_24719);
xor UO_664 (O_664,N_24636,N_24467);
or UO_665 (O_665,N_23986,N_24471);
nor UO_666 (O_666,N_24947,N_24210);
nor UO_667 (O_667,N_24516,N_24497);
or UO_668 (O_668,N_24492,N_24384);
nand UO_669 (O_669,N_24860,N_24985);
nand UO_670 (O_670,N_24132,N_24381);
nand UO_671 (O_671,N_24789,N_24525);
nor UO_672 (O_672,N_24835,N_24561);
nand UO_673 (O_673,N_24200,N_24670);
nor UO_674 (O_674,N_24016,N_24936);
and UO_675 (O_675,N_24884,N_24593);
nand UO_676 (O_676,N_24590,N_24833);
nand UO_677 (O_677,N_24083,N_24542);
nand UO_678 (O_678,N_24476,N_24017);
nor UO_679 (O_679,N_24604,N_24707);
xnor UO_680 (O_680,N_24294,N_24589);
xnor UO_681 (O_681,N_24404,N_24684);
xor UO_682 (O_682,N_24123,N_23993);
xor UO_683 (O_683,N_24145,N_24683);
or UO_684 (O_684,N_24453,N_24498);
and UO_685 (O_685,N_24263,N_23985);
nor UO_686 (O_686,N_24699,N_24994);
nor UO_687 (O_687,N_24638,N_24193);
xnor UO_688 (O_688,N_24952,N_24114);
xor UO_689 (O_689,N_24844,N_23752);
nor UO_690 (O_690,N_24869,N_23835);
and UO_691 (O_691,N_24123,N_23906);
or UO_692 (O_692,N_23923,N_24453);
nor UO_693 (O_693,N_23988,N_24058);
or UO_694 (O_694,N_24980,N_23951);
or UO_695 (O_695,N_24960,N_23796);
nor UO_696 (O_696,N_23877,N_23886);
xor UO_697 (O_697,N_24072,N_24160);
or UO_698 (O_698,N_24306,N_24355);
and UO_699 (O_699,N_24604,N_24490);
and UO_700 (O_700,N_24723,N_23925);
or UO_701 (O_701,N_24541,N_24696);
or UO_702 (O_702,N_24511,N_24626);
nor UO_703 (O_703,N_24306,N_24556);
nand UO_704 (O_704,N_24385,N_24221);
xor UO_705 (O_705,N_24021,N_24728);
nor UO_706 (O_706,N_24945,N_24948);
xnor UO_707 (O_707,N_24012,N_24207);
xor UO_708 (O_708,N_24541,N_24031);
or UO_709 (O_709,N_24772,N_24545);
xor UO_710 (O_710,N_23867,N_24980);
and UO_711 (O_711,N_24125,N_23910);
nand UO_712 (O_712,N_24437,N_24446);
xor UO_713 (O_713,N_24306,N_24934);
and UO_714 (O_714,N_24667,N_24392);
or UO_715 (O_715,N_24532,N_24645);
nand UO_716 (O_716,N_24953,N_23908);
and UO_717 (O_717,N_24327,N_24722);
nand UO_718 (O_718,N_24647,N_23839);
nor UO_719 (O_719,N_24624,N_24060);
nand UO_720 (O_720,N_24711,N_24529);
and UO_721 (O_721,N_24604,N_24588);
and UO_722 (O_722,N_23968,N_23829);
nor UO_723 (O_723,N_24289,N_23857);
or UO_724 (O_724,N_24925,N_23857);
nor UO_725 (O_725,N_23825,N_24399);
and UO_726 (O_726,N_24004,N_23990);
or UO_727 (O_727,N_24865,N_24215);
and UO_728 (O_728,N_24240,N_24042);
and UO_729 (O_729,N_24090,N_24763);
nand UO_730 (O_730,N_23807,N_23972);
nand UO_731 (O_731,N_24450,N_24683);
nand UO_732 (O_732,N_24567,N_24370);
or UO_733 (O_733,N_24090,N_24035);
xor UO_734 (O_734,N_24214,N_24897);
nand UO_735 (O_735,N_23947,N_24496);
nand UO_736 (O_736,N_24571,N_24459);
nand UO_737 (O_737,N_24818,N_24126);
nand UO_738 (O_738,N_24769,N_23867);
nand UO_739 (O_739,N_24837,N_23956);
or UO_740 (O_740,N_24653,N_24826);
nand UO_741 (O_741,N_24374,N_23816);
nand UO_742 (O_742,N_24161,N_24955);
or UO_743 (O_743,N_24284,N_24119);
or UO_744 (O_744,N_24536,N_24927);
nor UO_745 (O_745,N_24192,N_24020);
and UO_746 (O_746,N_24823,N_24356);
and UO_747 (O_747,N_24297,N_23774);
nor UO_748 (O_748,N_24768,N_24794);
xnor UO_749 (O_749,N_24658,N_24029);
xnor UO_750 (O_750,N_24234,N_24445);
or UO_751 (O_751,N_23864,N_24172);
or UO_752 (O_752,N_24831,N_24979);
nand UO_753 (O_753,N_24225,N_23792);
xor UO_754 (O_754,N_24105,N_23911);
or UO_755 (O_755,N_24112,N_24073);
or UO_756 (O_756,N_24853,N_24573);
nor UO_757 (O_757,N_23803,N_23955);
and UO_758 (O_758,N_24138,N_23864);
nor UO_759 (O_759,N_24652,N_24728);
nor UO_760 (O_760,N_24349,N_24572);
or UO_761 (O_761,N_23942,N_24426);
nand UO_762 (O_762,N_23755,N_24669);
or UO_763 (O_763,N_24269,N_24522);
and UO_764 (O_764,N_23977,N_24333);
and UO_765 (O_765,N_24519,N_23834);
and UO_766 (O_766,N_24420,N_23843);
xor UO_767 (O_767,N_24420,N_24708);
nand UO_768 (O_768,N_24461,N_24804);
nand UO_769 (O_769,N_24739,N_24871);
xnor UO_770 (O_770,N_23845,N_24206);
or UO_771 (O_771,N_24084,N_23762);
nand UO_772 (O_772,N_24895,N_24515);
xnor UO_773 (O_773,N_24630,N_24349);
xor UO_774 (O_774,N_24078,N_24971);
nor UO_775 (O_775,N_23994,N_24061);
xor UO_776 (O_776,N_23906,N_24501);
nand UO_777 (O_777,N_24343,N_24577);
and UO_778 (O_778,N_24418,N_24876);
xor UO_779 (O_779,N_24377,N_24790);
or UO_780 (O_780,N_24765,N_24285);
nor UO_781 (O_781,N_24840,N_24145);
xor UO_782 (O_782,N_24785,N_24692);
or UO_783 (O_783,N_24555,N_23824);
and UO_784 (O_784,N_24600,N_24929);
or UO_785 (O_785,N_24532,N_24845);
and UO_786 (O_786,N_24020,N_24783);
nor UO_787 (O_787,N_24468,N_24377);
nand UO_788 (O_788,N_23943,N_24832);
xnor UO_789 (O_789,N_24153,N_23902);
or UO_790 (O_790,N_24233,N_24612);
xor UO_791 (O_791,N_24832,N_24745);
nor UO_792 (O_792,N_24472,N_24120);
or UO_793 (O_793,N_24619,N_24853);
nor UO_794 (O_794,N_23969,N_24061);
or UO_795 (O_795,N_24059,N_23856);
nand UO_796 (O_796,N_24019,N_24804);
xnor UO_797 (O_797,N_24800,N_24812);
or UO_798 (O_798,N_23790,N_24403);
and UO_799 (O_799,N_24523,N_24318);
nor UO_800 (O_800,N_24689,N_24292);
xor UO_801 (O_801,N_24794,N_24881);
and UO_802 (O_802,N_24845,N_24485);
and UO_803 (O_803,N_24038,N_24328);
or UO_804 (O_804,N_23837,N_24122);
or UO_805 (O_805,N_24304,N_24552);
xor UO_806 (O_806,N_24352,N_24199);
or UO_807 (O_807,N_24232,N_24966);
nor UO_808 (O_808,N_23958,N_23977);
nand UO_809 (O_809,N_24623,N_24758);
xnor UO_810 (O_810,N_24076,N_23911);
xor UO_811 (O_811,N_23973,N_24707);
or UO_812 (O_812,N_24635,N_24683);
or UO_813 (O_813,N_24537,N_24329);
and UO_814 (O_814,N_23809,N_24089);
or UO_815 (O_815,N_24429,N_24518);
xor UO_816 (O_816,N_24500,N_24205);
and UO_817 (O_817,N_23992,N_24226);
nand UO_818 (O_818,N_24673,N_24341);
nor UO_819 (O_819,N_24109,N_24476);
nand UO_820 (O_820,N_24017,N_24991);
nand UO_821 (O_821,N_24067,N_23806);
nand UO_822 (O_822,N_24874,N_23971);
xor UO_823 (O_823,N_24018,N_24170);
nor UO_824 (O_824,N_23773,N_24710);
nand UO_825 (O_825,N_23815,N_24459);
or UO_826 (O_826,N_24671,N_23874);
nor UO_827 (O_827,N_24780,N_24737);
nor UO_828 (O_828,N_24436,N_24903);
or UO_829 (O_829,N_23931,N_24503);
nor UO_830 (O_830,N_24875,N_24709);
xor UO_831 (O_831,N_24907,N_24115);
nand UO_832 (O_832,N_24848,N_24797);
nand UO_833 (O_833,N_24103,N_24219);
or UO_834 (O_834,N_24296,N_24720);
nand UO_835 (O_835,N_24612,N_23905);
or UO_836 (O_836,N_23994,N_24765);
and UO_837 (O_837,N_23934,N_23762);
nand UO_838 (O_838,N_24826,N_24450);
nand UO_839 (O_839,N_24132,N_23863);
xor UO_840 (O_840,N_24658,N_24779);
nand UO_841 (O_841,N_24898,N_23911);
nor UO_842 (O_842,N_23965,N_24568);
nand UO_843 (O_843,N_24854,N_23849);
xnor UO_844 (O_844,N_24708,N_24250);
and UO_845 (O_845,N_23968,N_24202);
nor UO_846 (O_846,N_24893,N_23753);
nand UO_847 (O_847,N_23917,N_24242);
or UO_848 (O_848,N_24662,N_24342);
and UO_849 (O_849,N_24983,N_24317);
nor UO_850 (O_850,N_24600,N_24653);
or UO_851 (O_851,N_24747,N_24203);
and UO_852 (O_852,N_24575,N_24195);
nor UO_853 (O_853,N_24936,N_24377);
nor UO_854 (O_854,N_24990,N_24276);
or UO_855 (O_855,N_23783,N_24447);
nor UO_856 (O_856,N_24375,N_23881);
nor UO_857 (O_857,N_24492,N_24597);
and UO_858 (O_858,N_24472,N_24757);
nand UO_859 (O_859,N_24264,N_23849);
and UO_860 (O_860,N_24437,N_24673);
nor UO_861 (O_861,N_23986,N_24864);
nor UO_862 (O_862,N_24704,N_24555);
or UO_863 (O_863,N_24347,N_24579);
nor UO_864 (O_864,N_24269,N_24177);
or UO_865 (O_865,N_24771,N_24247);
nand UO_866 (O_866,N_23870,N_24854);
nor UO_867 (O_867,N_24242,N_24931);
or UO_868 (O_868,N_24573,N_24663);
and UO_869 (O_869,N_24522,N_24842);
and UO_870 (O_870,N_23908,N_24387);
nor UO_871 (O_871,N_24490,N_24735);
nand UO_872 (O_872,N_23931,N_24843);
nor UO_873 (O_873,N_24859,N_24925);
nor UO_874 (O_874,N_24283,N_24089);
xnor UO_875 (O_875,N_24276,N_24455);
or UO_876 (O_876,N_24458,N_23990);
or UO_877 (O_877,N_24832,N_24565);
nor UO_878 (O_878,N_24897,N_24482);
and UO_879 (O_879,N_24692,N_23756);
xnor UO_880 (O_880,N_24621,N_24287);
or UO_881 (O_881,N_24421,N_24431);
nor UO_882 (O_882,N_24976,N_24899);
xor UO_883 (O_883,N_24438,N_24649);
xnor UO_884 (O_884,N_23805,N_24479);
nor UO_885 (O_885,N_24879,N_24898);
and UO_886 (O_886,N_24110,N_24506);
nor UO_887 (O_887,N_24235,N_24341);
nand UO_888 (O_888,N_24342,N_24985);
nand UO_889 (O_889,N_24290,N_24876);
nand UO_890 (O_890,N_24310,N_24492);
xnor UO_891 (O_891,N_24853,N_24426);
and UO_892 (O_892,N_24666,N_24280);
and UO_893 (O_893,N_24948,N_24411);
nand UO_894 (O_894,N_24846,N_24865);
xnor UO_895 (O_895,N_24633,N_24716);
nor UO_896 (O_896,N_23773,N_24688);
or UO_897 (O_897,N_24261,N_24671);
nor UO_898 (O_898,N_24220,N_24801);
or UO_899 (O_899,N_24885,N_24663);
and UO_900 (O_900,N_23891,N_24739);
nor UO_901 (O_901,N_24392,N_24090);
or UO_902 (O_902,N_24192,N_24952);
and UO_903 (O_903,N_24108,N_23890);
nand UO_904 (O_904,N_24836,N_23882);
nand UO_905 (O_905,N_24512,N_24609);
xnor UO_906 (O_906,N_24511,N_24390);
nand UO_907 (O_907,N_23808,N_23991);
and UO_908 (O_908,N_24520,N_24877);
or UO_909 (O_909,N_24621,N_24025);
nor UO_910 (O_910,N_24826,N_24439);
nand UO_911 (O_911,N_24037,N_24150);
and UO_912 (O_912,N_24650,N_24377);
nand UO_913 (O_913,N_24691,N_24283);
nor UO_914 (O_914,N_23885,N_23789);
or UO_915 (O_915,N_24379,N_23880);
or UO_916 (O_916,N_23876,N_24858);
and UO_917 (O_917,N_24395,N_24369);
nand UO_918 (O_918,N_24578,N_23826);
nand UO_919 (O_919,N_24292,N_24377);
xor UO_920 (O_920,N_24784,N_24099);
nand UO_921 (O_921,N_23756,N_24705);
nor UO_922 (O_922,N_24421,N_24320);
xnor UO_923 (O_923,N_23794,N_23833);
nor UO_924 (O_924,N_24886,N_24696);
xnor UO_925 (O_925,N_24639,N_24858);
and UO_926 (O_926,N_23975,N_24846);
nor UO_927 (O_927,N_24030,N_23778);
nor UO_928 (O_928,N_24805,N_24001);
nand UO_929 (O_929,N_24368,N_24046);
nand UO_930 (O_930,N_23951,N_23940);
nor UO_931 (O_931,N_24112,N_24330);
and UO_932 (O_932,N_23903,N_23994);
xor UO_933 (O_933,N_24255,N_24789);
nand UO_934 (O_934,N_24898,N_24250);
and UO_935 (O_935,N_23771,N_23820);
and UO_936 (O_936,N_23837,N_24549);
nand UO_937 (O_937,N_24665,N_24286);
and UO_938 (O_938,N_23869,N_24672);
and UO_939 (O_939,N_24663,N_24984);
or UO_940 (O_940,N_24145,N_24123);
nand UO_941 (O_941,N_24449,N_24889);
and UO_942 (O_942,N_23963,N_23899);
and UO_943 (O_943,N_24191,N_24343);
and UO_944 (O_944,N_24934,N_24927);
and UO_945 (O_945,N_24172,N_24143);
or UO_946 (O_946,N_23848,N_24749);
nand UO_947 (O_947,N_24528,N_24508);
xor UO_948 (O_948,N_23777,N_24972);
nor UO_949 (O_949,N_23975,N_24831);
nor UO_950 (O_950,N_23966,N_24634);
or UO_951 (O_951,N_24853,N_24896);
nor UO_952 (O_952,N_24916,N_24932);
nand UO_953 (O_953,N_24716,N_24318);
and UO_954 (O_954,N_24593,N_23997);
nand UO_955 (O_955,N_24004,N_24417);
or UO_956 (O_956,N_24502,N_24414);
or UO_957 (O_957,N_24237,N_23842);
nor UO_958 (O_958,N_24389,N_23858);
nor UO_959 (O_959,N_24146,N_24475);
xnor UO_960 (O_960,N_24013,N_24988);
and UO_961 (O_961,N_24655,N_24742);
or UO_962 (O_962,N_23814,N_23905);
and UO_963 (O_963,N_24701,N_23936);
nor UO_964 (O_964,N_24366,N_23952);
or UO_965 (O_965,N_24051,N_24356);
nor UO_966 (O_966,N_24628,N_24865);
nor UO_967 (O_967,N_24710,N_24108);
and UO_968 (O_968,N_24320,N_24922);
nor UO_969 (O_969,N_24656,N_24361);
nand UO_970 (O_970,N_24037,N_24351);
or UO_971 (O_971,N_23878,N_24433);
or UO_972 (O_972,N_24241,N_24296);
nand UO_973 (O_973,N_24282,N_24091);
nor UO_974 (O_974,N_24596,N_23881);
nor UO_975 (O_975,N_24275,N_24280);
nor UO_976 (O_976,N_24481,N_24901);
nor UO_977 (O_977,N_23975,N_24300);
nor UO_978 (O_978,N_24489,N_23984);
xnor UO_979 (O_979,N_23911,N_24265);
nor UO_980 (O_980,N_24943,N_24799);
nor UO_981 (O_981,N_24960,N_24629);
nor UO_982 (O_982,N_24242,N_24795);
and UO_983 (O_983,N_23802,N_24583);
xor UO_984 (O_984,N_24567,N_24534);
xor UO_985 (O_985,N_24290,N_24781);
nor UO_986 (O_986,N_24793,N_24945);
or UO_987 (O_987,N_24506,N_24230);
and UO_988 (O_988,N_23924,N_23804);
xor UO_989 (O_989,N_24687,N_24048);
nor UO_990 (O_990,N_23921,N_24543);
and UO_991 (O_991,N_23915,N_24430);
xor UO_992 (O_992,N_24368,N_24124);
nor UO_993 (O_993,N_24654,N_23792);
nand UO_994 (O_994,N_23896,N_24340);
and UO_995 (O_995,N_24875,N_24234);
nor UO_996 (O_996,N_24487,N_24659);
xnor UO_997 (O_997,N_24803,N_24419);
nor UO_998 (O_998,N_23927,N_24252);
xor UO_999 (O_999,N_24068,N_24123);
xor UO_1000 (O_1000,N_23957,N_24658);
xor UO_1001 (O_1001,N_24757,N_23979);
and UO_1002 (O_1002,N_24505,N_24381);
nor UO_1003 (O_1003,N_24764,N_24897);
or UO_1004 (O_1004,N_24269,N_24945);
or UO_1005 (O_1005,N_24756,N_24178);
xnor UO_1006 (O_1006,N_24391,N_24914);
and UO_1007 (O_1007,N_24986,N_24231);
xor UO_1008 (O_1008,N_24213,N_23933);
or UO_1009 (O_1009,N_24534,N_24993);
xor UO_1010 (O_1010,N_24721,N_24110);
nand UO_1011 (O_1011,N_24443,N_23771);
nor UO_1012 (O_1012,N_24077,N_24425);
nor UO_1013 (O_1013,N_24506,N_24858);
nor UO_1014 (O_1014,N_24979,N_23945);
or UO_1015 (O_1015,N_23973,N_24076);
nor UO_1016 (O_1016,N_24718,N_24903);
nor UO_1017 (O_1017,N_24027,N_24706);
nand UO_1018 (O_1018,N_24496,N_23824);
and UO_1019 (O_1019,N_23790,N_24824);
and UO_1020 (O_1020,N_24292,N_24879);
or UO_1021 (O_1021,N_23942,N_23969);
nand UO_1022 (O_1022,N_24874,N_24953);
and UO_1023 (O_1023,N_24694,N_24431);
nand UO_1024 (O_1024,N_23827,N_23893);
nand UO_1025 (O_1025,N_24972,N_24951);
nor UO_1026 (O_1026,N_24090,N_24665);
nand UO_1027 (O_1027,N_24105,N_24692);
nand UO_1028 (O_1028,N_24842,N_24904);
xnor UO_1029 (O_1029,N_24561,N_23927);
nand UO_1030 (O_1030,N_24436,N_24460);
or UO_1031 (O_1031,N_24877,N_24279);
nand UO_1032 (O_1032,N_23986,N_24965);
or UO_1033 (O_1033,N_23763,N_23822);
nand UO_1034 (O_1034,N_24415,N_24955);
nand UO_1035 (O_1035,N_24263,N_24726);
or UO_1036 (O_1036,N_24837,N_24094);
or UO_1037 (O_1037,N_23966,N_24959);
xnor UO_1038 (O_1038,N_24212,N_24959);
nand UO_1039 (O_1039,N_24942,N_24160);
or UO_1040 (O_1040,N_23813,N_24796);
or UO_1041 (O_1041,N_24325,N_23876);
xnor UO_1042 (O_1042,N_24714,N_24952);
or UO_1043 (O_1043,N_24418,N_24530);
and UO_1044 (O_1044,N_24191,N_24990);
or UO_1045 (O_1045,N_24612,N_24483);
or UO_1046 (O_1046,N_24245,N_24127);
or UO_1047 (O_1047,N_24934,N_24713);
nor UO_1048 (O_1048,N_24844,N_24421);
nor UO_1049 (O_1049,N_24051,N_24628);
or UO_1050 (O_1050,N_24025,N_24372);
and UO_1051 (O_1051,N_24078,N_23836);
nand UO_1052 (O_1052,N_24937,N_24194);
or UO_1053 (O_1053,N_24218,N_24937);
nand UO_1054 (O_1054,N_23768,N_24656);
or UO_1055 (O_1055,N_24773,N_23975);
or UO_1056 (O_1056,N_24228,N_24632);
or UO_1057 (O_1057,N_24976,N_24724);
or UO_1058 (O_1058,N_24548,N_23940);
xnor UO_1059 (O_1059,N_24785,N_24130);
or UO_1060 (O_1060,N_24647,N_24838);
nand UO_1061 (O_1061,N_24388,N_24853);
xor UO_1062 (O_1062,N_24927,N_24732);
nand UO_1063 (O_1063,N_24808,N_24722);
nand UO_1064 (O_1064,N_24762,N_24991);
and UO_1065 (O_1065,N_24878,N_23923);
xor UO_1066 (O_1066,N_24822,N_24872);
nor UO_1067 (O_1067,N_24466,N_24399);
nand UO_1068 (O_1068,N_23833,N_23813);
xor UO_1069 (O_1069,N_24397,N_24185);
nand UO_1070 (O_1070,N_24609,N_24331);
xor UO_1071 (O_1071,N_24174,N_24801);
or UO_1072 (O_1072,N_24868,N_24200);
nor UO_1073 (O_1073,N_24980,N_24282);
nand UO_1074 (O_1074,N_24885,N_24426);
nor UO_1075 (O_1075,N_24868,N_24469);
xnor UO_1076 (O_1076,N_24568,N_24830);
and UO_1077 (O_1077,N_23765,N_24475);
or UO_1078 (O_1078,N_23757,N_24170);
xnor UO_1079 (O_1079,N_24230,N_24968);
xor UO_1080 (O_1080,N_23875,N_23993);
nor UO_1081 (O_1081,N_23769,N_24232);
nand UO_1082 (O_1082,N_24169,N_24443);
xor UO_1083 (O_1083,N_24486,N_23965);
nand UO_1084 (O_1084,N_24200,N_24408);
and UO_1085 (O_1085,N_23754,N_24404);
xnor UO_1086 (O_1086,N_23812,N_24411);
or UO_1087 (O_1087,N_24528,N_24099);
or UO_1088 (O_1088,N_24120,N_24772);
and UO_1089 (O_1089,N_23995,N_24434);
and UO_1090 (O_1090,N_24484,N_24401);
nor UO_1091 (O_1091,N_24390,N_24793);
nand UO_1092 (O_1092,N_24740,N_24458);
xor UO_1093 (O_1093,N_24994,N_24512);
xnor UO_1094 (O_1094,N_24480,N_23956);
and UO_1095 (O_1095,N_24493,N_24139);
xor UO_1096 (O_1096,N_24025,N_24991);
nand UO_1097 (O_1097,N_23937,N_24303);
nor UO_1098 (O_1098,N_24516,N_24871);
nor UO_1099 (O_1099,N_24061,N_23797);
or UO_1100 (O_1100,N_24165,N_24863);
and UO_1101 (O_1101,N_23954,N_24539);
xor UO_1102 (O_1102,N_24318,N_24236);
nand UO_1103 (O_1103,N_23926,N_24030);
xor UO_1104 (O_1104,N_24956,N_23986);
nor UO_1105 (O_1105,N_23906,N_23783);
or UO_1106 (O_1106,N_23781,N_24871);
and UO_1107 (O_1107,N_24074,N_24588);
nor UO_1108 (O_1108,N_24545,N_24857);
xnor UO_1109 (O_1109,N_24573,N_24020);
and UO_1110 (O_1110,N_24176,N_24235);
nand UO_1111 (O_1111,N_24479,N_24079);
and UO_1112 (O_1112,N_24658,N_24723);
or UO_1113 (O_1113,N_24757,N_24389);
xor UO_1114 (O_1114,N_23904,N_24641);
nand UO_1115 (O_1115,N_24301,N_23929);
xnor UO_1116 (O_1116,N_23931,N_24457);
nor UO_1117 (O_1117,N_24550,N_23853);
and UO_1118 (O_1118,N_24896,N_24078);
nand UO_1119 (O_1119,N_24154,N_24216);
nor UO_1120 (O_1120,N_23884,N_24044);
nor UO_1121 (O_1121,N_23772,N_23867);
nor UO_1122 (O_1122,N_24961,N_24026);
and UO_1123 (O_1123,N_24078,N_24583);
xor UO_1124 (O_1124,N_24304,N_24411);
nor UO_1125 (O_1125,N_23979,N_24580);
nor UO_1126 (O_1126,N_24488,N_23937);
or UO_1127 (O_1127,N_23766,N_24852);
nand UO_1128 (O_1128,N_24010,N_24641);
and UO_1129 (O_1129,N_24026,N_24201);
nand UO_1130 (O_1130,N_24218,N_24249);
nand UO_1131 (O_1131,N_24054,N_24398);
nor UO_1132 (O_1132,N_24754,N_24023);
nand UO_1133 (O_1133,N_24261,N_24560);
or UO_1134 (O_1134,N_24321,N_23751);
xnor UO_1135 (O_1135,N_23772,N_24279);
xor UO_1136 (O_1136,N_24838,N_24148);
xor UO_1137 (O_1137,N_23918,N_24493);
xnor UO_1138 (O_1138,N_23921,N_24346);
nor UO_1139 (O_1139,N_24072,N_24760);
or UO_1140 (O_1140,N_24584,N_24284);
and UO_1141 (O_1141,N_24325,N_24114);
and UO_1142 (O_1142,N_23890,N_24154);
or UO_1143 (O_1143,N_23948,N_23822);
nand UO_1144 (O_1144,N_24194,N_24230);
or UO_1145 (O_1145,N_23810,N_24267);
and UO_1146 (O_1146,N_24420,N_24198);
nor UO_1147 (O_1147,N_24337,N_24151);
xor UO_1148 (O_1148,N_24650,N_24409);
nor UO_1149 (O_1149,N_24197,N_24846);
or UO_1150 (O_1150,N_24248,N_23751);
nor UO_1151 (O_1151,N_24484,N_24082);
and UO_1152 (O_1152,N_24957,N_24115);
or UO_1153 (O_1153,N_23940,N_24731);
nand UO_1154 (O_1154,N_24855,N_23982);
nand UO_1155 (O_1155,N_24468,N_24575);
nor UO_1156 (O_1156,N_23870,N_24045);
or UO_1157 (O_1157,N_24470,N_24853);
nand UO_1158 (O_1158,N_24926,N_24478);
and UO_1159 (O_1159,N_24655,N_24162);
and UO_1160 (O_1160,N_23878,N_24146);
and UO_1161 (O_1161,N_24321,N_24022);
or UO_1162 (O_1162,N_23773,N_24701);
or UO_1163 (O_1163,N_24056,N_23857);
nand UO_1164 (O_1164,N_24002,N_24047);
or UO_1165 (O_1165,N_24437,N_24631);
and UO_1166 (O_1166,N_24163,N_24347);
or UO_1167 (O_1167,N_24336,N_24916);
nand UO_1168 (O_1168,N_24828,N_24017);
xnor UO_1169 (O_1169,N_24554,N_24553);
xor UO_1170 (O_1170,N_23847,N_24151);
nand UO_1171 (O_1171,N_24335,N_24443);
nand UO_1172 (O_1172,N_23802,N_24381);
nor UO_1173 (O_1173,N_24435,N_23930);
or UO_1174 (O_1174,N_24782,N_23784);
and UO_1175 (O_1175,N_24690,N_24911);
or UO_1176 (O_1176,N_24980,N_24036);
and UO_1177 (O_1177,N_24100,N_24352);
and UO_1178 (O_1178,N_24244,N_24208);
nand UO_1179 (O_1179,N_24081,N_24594);
nor UO_1180 (O_1180,N_24757,N_24802);
nand UO_1181 (O_1181,N_24035,N_23862);
nand UO_1182 (O_1182,N_24721,N_23790);
or UO_1183 (O_1183,N_24792,N_24111);
xnor UO_1184 (O_1184,N_24393,N_24664);
nand UO_1185 (O_1185,N_24562,N_24075);
and UO_1186 (O_1186,N_24525,N_24482);
or UO_1187 (O_1187,N_24349,N_24023);
and UO_1188 (O_1188,N_24520,N_24036);
nand UO_1189 (O_1189,N_23881,N_24729);
or UO_1190 (O_1190,N_24983,N_24083);
xnor UO_1191 (O_1191,N_23836,N_24051);
nor UO_1192 (O_1192,N_24447,N_24373);
nor UO_1193 (O_1193,N_24112,N_24724);
nand UO_1194 (O_1194,N_24976,N_23852);
nor UO_1195 (O_1195,N_24829,N_24815);
nand UO_1196 (O_1196,N_24452,N_24142);
and UO_1197 (O_1197,N_24230,N_24517);
nand UO_1198 (O_1198,N_24188,N_24346);
nor UO_1199 (O_1199,N_24710,N_24660);
nor UO_1200 (O_1200,N_24299,N_23970);
or UO_1201 (O_1201,N_24020,N_24999);
nand UO_1202 (O_1202,N_23993,N_24217);
and UO_1203 (O_1203,N_23841,N_24207);
or UO_1204 (O_1204,N_24328,N_24314);
xor UO_1205 (O_1205,N_24363,N_24689);
and UO_1206 (O_1206,N_24864,N_24211);
and UO_1207 (O_1207,N_24515,N_24341);
nor UO_1208 (O_1208,N_23903,N_23776);
or UO_1209 (O_1209,N_24457,N_24696);
or UO_1210 (O_1210,N_24248,N_24567);
xnor UO_1211 (O_1211,N_23799,N_24425);
xor UO_1212 (O_1212,N_24955,N_23930);
nor UO_1213 (O_1213,N_24598,N_24419);
nand UO_1214 (O_1214,N_24106,N_24077);
nand UO_1215 (O_1215,N_24053,N_24162);
and UO_1216 (O_1216,N_24115,N_23754);
and UO_1217 (O_1217,N_23968,N_24440);
nand UO_1218 (O_1218,N_24355,N_24423);
nand UO_1219 (O_1219,N_24913,N_24932);
or UO_1220 (O_1220,N_24648,N_24358);
or UO_1221 (O_1221,N_23775,N_24851);
nand UO_1222 (O_1222,N_23883,N_24323);
nor UO_1223 (O_1223,N_24421,N_24567);
and UO_1224 (O_1224,N_24833,N_23912);
xnor UO_1225 (O_1225,N_24330,N_24765);
nor UO_1226 (O_1226,N_24713,N_23959);
and UO_1227 (O_1227,N_24177,N_24948);
nand UO_1228 (O_1228,N_24800,N_24033);
nor UO_1229 (O_1229,N_24890,N_24031);
and UO_1230 (O_1230,N_24413,N_24222);
nor UO_1231 (O_1231,N_24268,N_24207);
nand UO_1232 (O_1232,N_23926,N_24879);
nand UO_1233 (O_1233,N_24384,N_23912);
nor UO_1234 (O_1234,N_23805,N_24035);
nand UO_1235 (O_1235,N_24459,N_24406);
and UO_1236 (O_1236,N_24989,N_23875);
xnor UO_1237 (O_1237,N_24706,N_24959);
or UO_1238 (O_1238,N_24358,N_24684);
nand UO_1239 (O_1239,N_24460,N_24529);
nor UO_1240 (O_1240,N_24965,N_24670);
xor UO_1241 (O_1241,N_24105,N_24086);
and UO_1242 (O_1242,N_23909,N_24702);
and UO_1243 (O_1243,N_24772,N_24174);
nor UO_1244 (O_1244,N_24470,N_24563);
and UO_1245 (O_1245,N_24757,N_24171);
or UO_1246 (O_1246,N_24658,N_24587);
nor UO_1247 (O_1247,N_24600,N_24896);
or UO_1248 (O_1248,N_24932,N_24985);
xnor UO_1249 (O_1249,N_24311,N_24267);
nand UO_1250 (O_1250,N_24999,N_24755);
nor UO_1251 (O_1251,N_23962,N_24779);
xor UO_1252 (O_1252,N_24814,N_24435);
nor UO_1253 (O_1253,N_23944,N_24067);
and UO_1254 (O_1254,N_24388,N_24633);
xor UO_1255 (O_1255,N_24975,N_24912);
or UO_1256 (O_1256,N_24196,N_24565);
and UO_1257 (O_1257,N_23913,N_24991);
nor UO_1258 (O_1258,N_23794,N_24766);
or UO_1259 (O_1259,N_24308,N_24972);
nand UO_1260 (O_1260,N_24255,N_24731);
xor UO_1261 (O_1261,N_23983,N_24315);
and UO_1262 (O_1262,N_24784,N_24004);
nand UO_1263 (O_1263,N_24865,N_24805);
and UO_1264 (O_1264,N_23812,N_24554);
nor UO_1265 (O_1265,N_23940,N_24873);
xor UO_1266 (O_1266,N_24381,N_24546);
xnor UO_1267 (O_1267,N_24397,N_24421);
and UO_1268 (O_1268,N_24818,N_24772);
and UO_1269 (O_1269,N_24546,N_23874);
xor UO_1270 (O_1270,N_24286,N_23788);
and UO_1271 (O_1271,N_24784,N_24216);
or UO_1272 (O_1272,N_24702,N_24661);
or UO_1273 (O_1273,N_24761,N_23986);
nor UO_1274 (O_1274,N_24984,N_24810);
nor UO_1275 (O_1275,N_24930,N_24744);
and UO_1276 (O_1276,N_24326,N_23934);
nor UO_1277 (O_1277,N_24279,N_24491);
and UO_1278 (O_1278,N_23832,N_24131);
or UO_1279 (O_1279,N_24473,N_24753);
and UO_1280 (O_1280,N_24217,N_23910);
and UO_1281 (O_1281,N_24566,N_24455);
xor UO_1282 (O_1282,N_24294,N_24122);
nor UO_1283 (O_1283,N_24644,N_24634);
xnor UO_1284 (O_1284,N_24499,N_24495);
nand UO_1285 (O_1285,N_23839,N_24928);
xnor UO_1286 (O_1286,N_23922,N_24621);
nor UO_1287 (O_1287,N_24510,N_24037);
xor UO_1288 (O_1288,N_23791,N_24548);
nand UO_1289 (O_1289,N_24598,N_24301);
or UO_1290 (O_1290,N_24227,N_24924);
nand UO_1291 (O_1291,N_24556,N_24171);
xor UO_1292 (O_1292,N_23936,N_23945);
and UO_1293 (O_1293,N_24479,N_23938);
nand UO_1294 (O_1294,N_24307,N_24855);
nor UO_1295 (O_1295,N_24316,N_24285);
nor UO_1296 (O_1296,N_24968,N_23923);
xnor UO_1297 (O_1297,N_24323,N_24739);
xnor UO_1298 (O_1298,N_24077,N_24434);
xnor UO_1299 (O_1299,N_24730,N_24007);
nand UO_1300 (O_1300,N_23986,N_23892);
xnor UO_1301 (O_1301,N_24255,N_24796);
xor UO_1302 (O_1302,N_24658,N_24623);
and UO_1303 (O_1303,N_24383,N_24405);
and UO_1304 (O_1304,N_24401,N_24872);
or UO_1305 (O_1305,N_24535,N_23809);
nor UO_1306 (O_1306,N_24689,N_24247);
nor UO_1307 (O_1307,N_24115,N_24997);
or UO_1308 (O_1308,N_23800,N_24661);
nand UO_1309 (O_1309,N_24514,N_24251);
xor UO_1310 (O_1310,N_24201,N_24734);
and UO_1311 (O_1311,N_23968,N_23800);
nand UO_1312 (O_1312,N_24383,N_24753);
nor UO_1313 (O_1313,N_24085,N_24784);
and UO_1314 (O_1314,N_23945,N_24800);
nand UO_1315 (O_1315,N_24829,N_24286);
xor UO_1316 (O_1316,N_24125,N_24187);
nor UO_1317 (O_1317,N_24456,N_24041);
nand UO_1318 (O_1318,N_23962,N_24610);
xor UO_1319 (O_1319,N_24535,N_24484);
and UO_1320 (O_1320,N_24622,N_24544);
xor UO_1321 (O_1321,N_23899,N_24109);
nor UO_1322 (O_1322,N_24892,N_24660);
and UO_1323 (O_1323,N_24576,N_24755);
nand UO_1324 (O_1324,N_24209,N_24223);
xor UO_1325 (O_1325,N_24510,N_24399);
nor UO_1326 (O_1326,N_24823,N_23869);
or UO_1327 (O_1327,N_24002,N_23946);
or UO_1328 (O_1328,N_23936,N_24822);
nand UO_1329 (O_1329,N_24352,N_24492);
or UO_1330 (O_1330,N_24629,N_24004);
and UO_1331 (O_1331,N_24686,N_24960);
or UO_1332 (O_1332,N_24861,N_24406);
xor UO_1333 (O_1333,N_24519,N_23852);
xnor UO_1334 (O_1334,N_24372,N_24264);
and UO_1335 (O_1335,N_24418,N_24707);
nor UO_1336 (O_1336,N_24185,N_24972);
or UO_1337 (O_1337,N_24200,N_24618);
nand UO_1338 (O_1338,N_23990,N_24662);
nor UO_1339 (O_1339,N_24225,N_24840);
xnor UO_1340 (O_1340,N_24886,N_24773);
and UO_1341 (O_1341,N_24486,N_23790);
or UO_1342 (O_1342,N_24255,N_24849);
or UO_1343 (O_1343,N_24860,N_23767);
nor UO_1344 (O_1344,N_24523,N_24599);
xor UO_1345 (O_1345,N_23884,N_24142);
and UO_1346 (O_1346,N_24310,N_24212);
or UO_1347 (O_1347,N_23952,N_24439);
nand UO_1348 (O_1348,N_24845,N_24936);
xnor UO_1349 (O_1349,N_24584,N_24470);
or UO_1350 (O_1350,N_24178,N_24068);
nand UO_1351 (O_1351,N_24096,N_24847);
nor UO_1352 (O_1352,N_24274,N_24830);
nor UO_1353 (O_1353,N_24656,N_24378);
xnor UO_1354 (O_1354,N_24514,N_24884);
or UO_1355 (O_1355,N_23798,N_24311);
and UO_1356 (O_1356,N_23974,N_23867);
nor UO_1357 (O_1357,N_24558,N_24999);
nor UO_1358 (O_1358,N_24954,N_24891);
and UO_1359 (O_1359,N_24357,N_24074);
xor UO_1360 (O_1360,N_24500,N_24078);
nand UO_1361 (O_1361,N_24980,N_24850);
nand UO_1362 (O_1362,N_24663,N_24980);
and UO_1363 (O_1363,N_24235,N_24434);
xnor UO_1364 (O_1364,N_24381,N_24548);
nand UO_1365 (O_1365,N_24020,N_24669);
or UO_1366 (O_1366,N_24703,N_24147);
nor UO_1367 (O_1367,N_24817,N_24178);
xor UO_1368 (O_1368,N_24781,N_24679);
and UO_1369 (O_1369,N_24469,N_23791);
and UO_1370 (O_1370,N_23969,N_24290);
xor UO_1371 (O_1371,N_24715,N_24287);
nor UO_1372 (O_1372,N_24873,N_24745);
xor UO_1373 (O_1373,N_24331,N_23921);
nand UO_1374 (O_1374,N_23810,N_24453);
nor UO_1375 (O_1375,N_24825,N_24769);
or UO_1376 (O_1376,N_24828,N_24404);
nor UO_1377 (O_1377,N_24229,N_24468);
nor UO_1378 (O_1378,N_24984,N_24061);
nor UO_1379 (O_1379,N_24432,N_24233);
nor UO_1380 (O_1380,N_24291,N_23976);
or UO_1381 (O_1381,N_24824,N_24684);
nand UO_1382 (O_1382,N_24216,N_24419);
or UO_1383 (O_1383,N_24071,N_24639);
nor UO_1384 (O_1384,N_24867,N_24420);
and UO_1385 (O_1385,N_24507,N_24157);
nor UO_1386 (O_1386,N_24217,N_23846);
or UO_1387 (O_1387,N_24793,N_24563);
nor UO_1388 (O_1388,N_24066,N_24487);
nor UO_1389 (O_1389,N_24468,N_23767);
and UO_1390 (O_1390,N_24153,N_23888);
nor UO_1391 (O_1391,N_24109,N_24052);
xor UO_1392 (O_1392,N_24871,N_23860);
xnor UO_1393 (O_1393,N_24324,N_24440);
nor UO_1394 (O_1394,N_24587,N_24908);
and UO_1395 (O_1395,N_24172,N_24655);
xor UO_1396 (O_1396,N_24198,N_24595);
nand UO_1397 (O_1397,N_24691,N_24035);
xor UO_1398 (O_1398,N_24279,N_24190);
nor UO_1399 (O_1399,N_24599,N_23761);
xor UO_1400 (O_1400,N_23814,N_24633);
and UO_1401 (O_1401,N_24960,N_24053);
xor UO_1402 (O_1402,N_23957,N_24414);
xnor UO_1403 (O_1403,N_24862,N_24529);
nand UO_1404 (O_1404,N_23917,N_24103);
nand UO_1405 (O_1405,N_24403,N_23857);
and UO_1406 (O_1406,N_24968,N_24769);
or UO_1407 (O_1407,N_24072,N_24151);
or UO_1408 (O_1408,N_24591,N_24717);
nand UO_1409 (O_1409,N_24988,N_24846);
nor UO_1410 (O_1410,N_24280,N_24068);
nor UO_1411 (O_1411,N_24890,N_24820);
nor UO_1412 (O_1412,N_24784,N_23923);
or UO_1413 (O_1413,N_24288,N_24183);
nand UO_1414 (O_1414,N_24158,N_24400);
xnor UO_1415 (O_1415,N_24038,N_24767);
nor UO_1416 (O_1416,N_23864,N_24393);
nor UO_1417 (O_1417,N_23750,N_23831);
xnor UO_1418 (O_1418,N_24381,N_24700);
and UO_1419 (O_1419,N_24626,N_24518);
and UO_1420 (O_1420,N_23907,N_24834);
xnor UO_1421 (O_1421,N_23861,N_23829);
nand UO_1422 (O_1422,N_24714,N_24678);
or UO_1423 (O_1423,N_23995,N_24847);
or UO_1424 (O_1424,N_24912,N_24357);
or UO_1425 (O_1425,N_24252,N_24049);
or UO_1426 (O_1426,N_24036,N_24369);
and UO_1427 (O_1427,N_23789,N_24704);
xor UO_1428 (O_1428,N_23900,N_24838);
xor UO_1429 (O_1429,N_23871,N_24940);
xnor UO_1430 (O_1430,N_24881,N_24631);
xnor UO_1431 (O_1431,N_23971,N_24612);
nor UO_1432 (O_1432,N_24310,N_24979);
xor UO_1433 (O_1433,N_24822,N_24315);
xor UO_1434 (O_1434,N_23760,N_24484);
and UO_1435 (O_1435,N_24418,N_24538);
nor UO_1436 (O_1436,N_24049,N_24384);
nand UO_1437 (O_1437,N_24825,N_23829);
xor UO_1438 (O_1438,N_24809,N_24054);
nand UO_1439 (O_1439,N_24913,N_24303);
xnor UO_1440 (O_1440,N_23806,N_24242);
nor UO_1441 (O_1441,N_24959,N_24369);
or UO_1442 (O_1442,N_23946,N_24092);
or UO_1443 (O_1443,N_24936,N_24440);
nor UO_1444 (O_1444,N_23976,N_24963);
nand UO_1445 (O_1445,N_24691,N_23885);
xnor UO_1446 (O_1446,N_23848,N_24287);
and UO_1447 (O_1447,N_24328,N_24023);
nor UO_1448 (O_1448,N_24851,N_24474);
or UO_1449 (O_1449,N_24043,N_24259);
and UO_1450 (O_1450,N_24202,N_24631);
xnor UO_1451 (O_1451,N_23783,N_24538);
nand UO_1452 (O_1452,N_24996,N_24219);
nand UO_1453 (O_1453,N_24214,N_23924);
nor UO_1454 (O_1454,N_23945,N_23821);
and UO_1455 (O_1455,N_24980,N_24184);
nor UO_1456 (O_1456,N_24296,N_23998);
xnor UO_1457 (O_1457,N_24289,N_24016);
or UO_1458 (O_1458,N_23891,N_24600);
nor UO_1459 (O_1459,N_24139,N_24234);
or UO_1460 (O_1460,N_24775,N_24552);
xor UO_1461 (O_1461,N_24090,N_24555);
or UO_1462 (O_1462,N_24861,N_24035);
nand UO_1463 (O_1463,N_23920,N_24678);
or UO_1464 (O_1464,N_24919,N_23834);
xor UO_1465 (O_1465,N_24454,N_24711);
xnor UO_1466 (O_1466,N_24383,N_24588);
nand UO_1467 (O_1467,N_24966,N_24270);
and UO_1468 (O_1468,N_24195,N_24320);
xor UO_1469 (O_1469,N_24323,N_24106);
and UO_1470 (O_1470,N_24758,N_23781);
or UO_1471 (O_1471,N_24486,N_24159);
nand UO_1472 (O_1472,N_23989,N_24341);
and UO_1473 (O_1473,N_24749,N_24362);
or UO_1474 (O_1474,N_24809,N_24693);
nand UO_1475 (O_1475,N_24042,N_24995);
or UO_1476 (O_1476,N_24500,N_23996);
and UO_1477 (O_1477,N_23920,N_24483);
nor UO_1478 (O_1478,N_24787,N_24886);
nand UO_1479 (O_1479,N_24126,N_24000);
nor UO_1480 (O_1480,N_24614,N_24400);
nor UO_1481 (O_1481,N_24408,N_24871);
nand UO_1482 (O_1482,N_24035,N_24784);
or UO_1483 (O_1483,N_24981,N_24394);
or UO_1484 (O_1484,N_24009,N_24963);
and UO_1485 (O_1485,N_24066,N_24359);
or UO_1486 (O_1486,N_24679,N_24267);
nor UO_1487 (O_1487,N_24059,N_24258);
or UO_1488 (O_1488,N_24081,N_24098);
nand UO_1489 (O_1489,N_24854,N_24683);
xnor UO_1490 (O_1490,N_24364,N_24935);
nand UO_1491 (O_1491,N_24605,N_24273);
and UO_1492 (O_1492,N_24431,N_24216);
or UO_1493 (O_1493,N_24241,N_24537);
nand UO_1494 (O_1494,N_23854,N_24665);
nand UO_1495 (O_1495,N_24782,N_23774);
and UO_1496 (O_1496,N_24310,N_24675);
nor UO_1497 (O_1497,N_24423,N_24593);
nand UO_1498 (O_1498,N_24490,N_24786);
nand UO_1499 (O_1499,N_24944,N_24060);
nor UO_1500 (O_1500,N_24580,N_24422);
xor UO_1501 (O_1501,N_24465,N_23918);
and UO_1502 (O_1502,N_23799,N_24005);
nor UO_1503 (O_1503,N_23866,N_24716);
nand UO_1504 (O_1504,N_24165,N_24720);
nand UO_1505 (O_1505,N_24863,N_24410);
xor UO_1506 (O_1506,N_24582,N_24894);
or UO_1507 (O_1507,N_23814,N_23754);
nor UO_1508 (O_1508,N_23777,N_23889);
or UO_1509 (O_1509,N_24650,N_23812);
xor UO_1510 (O_1510,N_24387,N_23885);
nor UO_1511 (O_1511,N_24275,N_23859);
and UO_1512 (O_1512,N_23751,N_24468);
or UO_1513 (O_1513,N_24321,N_24714);
and UO_1514 (O_1514,N_24682,N_24264);
xor UO_1515 (O_1515,N_23966,N_23776);
nor UO_1516 (O_1516,N_23754,N_24319);
and UO_1517 (O_1517,N_24967,N_24283);
and UO_1518 (O_1518,N_24427,N_23964);
xnor UO_1519 (O_1519,N_24419,N_24125);
or UO_1520 (O_1520,N_24845,N_24333);
nand UO_1521 (O_1521,N_24434,N_24362);
xnor UO_1522 (O_1522,N_24937,N_24052);
and UO_1523 (O_1523,N_24177,N_24333);
xor UO_1524 (O_1524,N_24684,N_23821);
and UO_1525 (O_1525,N_24252,N_23826);
nor UO_1526 (O_1526,N_24550,N_24731);
nor UO_1527 (O_1527,N_24795,N_23869);
and UO_1528 (O_1528,N_24437,N_23766);
or UO_1529 (O_1529,N_24193,N_24087);
nor UO_1530 (O_1530,N_24666,N_24138);
nor UO_1531 (O_1531,N_24276,N_24255);
nor UO_1532 (O_1532,N_23764,N_24216);
nor UO_1533 (O_1533,N_24552,N_23824);
and UO_1534 (O_1534,N_24606,N_24895);
nand UO_1535 (O_1535,N_24437,N_24881);
nand UO_1536 (O_1536,N_23965,N_24611);
nand UO_1537 (O_1537,N_24699,N_24625);
and UO_1538 (O_1538,N_23768,N_24968);
nand UO_1539 (O_1539,N_24131,N_24687);
or UO_1540 (O_1540,N_23966,N_24442);
nor UO_1541 (O_1541,N_24444,N_24943);
and UO_1542 (O_1542,N_23859,N_24098);
nand UO_1543 (O_1543,N_23817,N_24178);
and UO_1544 (O_1544,N_23985,N_23832);
or UO_1545 (O_1545,N_24666,N_23896);
and UO_1546 (O_1546,N_24906,N_24789);
nand UO_1547 (O_1547,N_24846,N_24431);
nand UO_1548 (O_1548,N_24579,N_24952);
nor UO_1549 (O_1549,N_24529,N_23836);
and UO_1550 (O_1550,N_24344,N_24216);
or UO_1551 (O_1551,N_24534,N_24152);
nor UO_1552 (O_1552,N_24406,N_24240);
or UO_1553 (O_1553,N_24160,N_24869);
xnor UO_1554 (O_1554,N_24223,N_24362);
nand UO_1555 (O_1555,N_24126,N_24580);
and UO_1556 (O_1556,N_24456,N_24278);
nand UO_1557 (O_1557,N_24767,N_23761);
nand UO_1558 (O_1558,N_23810,N_24110);
or UO_1559 (O_1559,N_23798,N_23898);
nand UO_1560 (O_1560,N_24658,N_23797);
and UO_1561 (O_1561,N_24787,N_24757);
and UO_1562 (O_1562,N_24236,N_24593);
or UO_1563 (O_1563,N_24231,N_24054);
xnor UO_1564 (O_1564,N_24945,N_24365);
xor UO_1565 (O_1565,N_24631,N_23797);
or UO_1566 (O_1566,N_24911,N_24295);
and UO_1567 (O_1567,N_24269,N_24476);
nand UO_1568 (O_1568,N_24428,N_24681);
nor UO_1569 (O_1569,N_24265,N_24879);
nand UO_1570 (O_1570,N_24334,N_23808);
or UO_1571 (O_1571,N_23941,N_24073);
nor UO_1572 (O_1572,N_23794,N_24699);
nor UO_1573 (O_1573,N_24091,N_24657);
or UO_1574 (O_1574,N_24348,N_24206);
xnor UO_1575 (O_1575,N_24230,N_23804);
nand UO_1576 (O_1576,N_24202,N_24882);
xnor UO_1577 (O_1577,N_24032,N_24279);
nor UO_1578 (O_1578,N_24701,N_24472);
xor UO_1579 (O_1579,N_24605,N_24382);
nand UO_1580 (O_1580,N_24451,N_24371);
nand UO_1581 (O_1581,N_24456,N_23903);
and UO_1582 (O_1582,N_24257,N_23776);
nand UO_1583 (O_1583,N_23780,N_23954);
and UO_1584 (O_1584,N_24002,N_24355);
or UO_1585 (O_1585,N_23996,N_24527);
or UO_1586 (O_1586,N_24173,N_24762);
and UO_1587 (O_1587,N_24139,N_24254);
xnor UO_1588 (O_1588,N_24134,N_24409);
nand UO_1589 (O_1589,N_24389,N_24781);
nor UO_1590 (O_1590,N_24750,N_23939);
and UO_1591 (O_1591,N_24006,N_24217);
or UO_1592 (O_1592,N_23861,N_24430);
nor UO_1593 (O_1593,N_24835,N_23760);
nor UO_1594 (O_1594,N_24341,N_24943);
and UO_1595 (O_1595,N_24678,N_24244);
nor UO_1596 (O_1596,N_24906,N_24029);
or UO_1597 (O_1597,N_23966,N_23944);
or UO_1598 (O_1598,N_24508,N_23873);
xor UO_1599 (O_1599,N_24615,N_24034);
and UO_1600 (O_1600,N_24769,N_24049);
or UO_1601 (O_1601,N_24420,N_24463);
xor UO_1602 (O_1602,N_24302,N_24934);
xnor UO_1603 (O_1603,N_23808,N_24879);
nor UO_1604 (O_1604,N_24636,N_24537);
and UO_1605 (O_1605,N_24973,N_24578);
and UO_1606 (O_1606,N_24286,N_24379);
nand UO_1607 (O_1607,N_24545,N_23881);
and UO_1608 (O_1608,N_24004,N_24425);
or UO_1609 (O_1609,N_24452,N_24810);
and UO_1610 (O_1610,N_24767,N_24286);
nor UO_1611 (O_1611,N_24005,N_24561);
xor UO_1612 (O_1612,N_24124,N_24152);
nand UO_1613 (O_1613,N_24943,N_24629);
nor UO_1614 (O_1614,N_24321,N_24060);
xor UO_1615 (O_1615,N_23986,N_24193);
or UO_1616 (O_1616,N_24714,N_24544);
xnor UO_1617 (O_1617,N_24006,N_24861);
nor UO_1618 (O_1618,N_24691,N_24442);
xor UO_1619 (O_1619,N_23851,N_24166);
or UO_1620 (O_1620,N_24137,N_24246);
nor UO_1621 (O_1621,N_24808,N_24051);
nand UO_1622 (O_1622,N_24413,N_24854);
or UO_1623 (O_1623,N_23893,N_24558);
nor UO_1624 (O_1624,N_24687,N_24155);
xor UO_1625 (O_1625,N_24440,N_23879);
and UO_1626 (O_1626,N_23981,N_24347);
or UO_1627 (O_1627,N_24543,N_24761);
nor UO_1628 (O_1628,N_24571,N_24474);
nor UO_1629 (O_1629,N_24003,N_24661);
nor UO_1630 (O_1630,N_24817,N_24308);
xnor UO_1631 (O_1631,N_23942,N_24302);
nor UO_1632 (O_1632,N_24136,N_24187);
and UO_1633 (O_1633,N_23912,N_24736);
or UO_1634 (O_1634,N_24558,N_24000);
and UO_1635 (O_1635,N_24883,N_24834);
xnor UO_1636 (O_1636,N_24442,N_24505);
nor UO_1637 (O_1637,N_24368,N_24701);
xnor UO_1638 (O_1638,N_24600,N_24993);
and UO_1639 (O_1639,N_24612,N_24516);
nand UO_1640 (O_1640,N_24244,N_24059);
or UO_1641 (O_1641,N_24344,N_24705);
xnor UO_1642 (O_1642,N_24550,N_24773);
xnor UO_1643 (O_1643,N_24919,N_23805);
and UO_1644 (O_1644,N_24734,N_24635);
and UO_1645 (O_1645,N_24156,N_24957);
nand UO_1646 (O_1646,N_24851,N_24796);
nand UO_1647 (O_1647,N_24412,N_24381);
nor UO_1648 (O_1648,N_24341,N_24967);
nand UO_1649 (O_1649,N_24710,N_24608);
or UO_1650 (O_1650,N_24799,N_24290);
or UO_1651 (O_1651,N_24781,N_24025);
nor UO_1652 (O_1652,N_24686,N_24692);
xnor UO_1653 (O_1653,N_24394,N_23921);
xnor UO_1654 (O_1654,N_23762,N_24517);
and UO_1655 (O_1655,N_23966,N_24513);
or UO_1656 (O_1656,N_24512,N_24460);
nand UO_1657 (O_1657,N_23753,N_24382);
and UO_1658 (O_1658,N_24109,N_24295);
nor UO_1659 (O_1659,N_23938,N_23990);
or UO_1660 (O_1660,N_24351,N_24396);
and UO_1661 (O_1661,N_23902,N_24414);
nor UO_1662 (O_1662,N_23964,N_24455);
nor UO_1663 (O_1663,N_24621,N_24724);
and UO_1664 (O_1664,N_24972,N_24018);
or UO_1665 (O_1665,N_24648,N_24644);
or UO_1666 (O_1666,N_24660,N_24330);
and UO_1667 (O_1667,N_24577,N_24323);
or UO_1668 (O_1668,N_24863,N_24063);
nand UO_1669 (O_1669,N_24459,N_24279);
and UO_1670 (O_1670,N_24506,N_24112);
or UO_1671 (O_1671,N_24480,N_23959);
nor UO_1672 (O_1672,N_23864,N_24997);
xor UO_1673 (O_1673,N_24896,N_24534);
and UO_1674 (O_1674,N_23901,N_24075);
xnor UO_1675 (O_1675,N_23850,N_23799);
and UO_1676 (O_1676,N_24733,N_23820);
xnor UO_1677 (O_1677,N_24091,N_23766);
nand UO_1678 (O_1678,N_24996,N_24939);
and UO_1679 (O_1679,N_24369,N_24805);
and UO_1680 (O_1680,N_23914,N_23835);
nand UO_1681 (O_1681,N_24885,N_23784);
xnor UO_1682 (O_1682,N_23777,N_24903);
xnor UO_1683 (O_1683,N_24584,N_24767);
and UO_1684 (O_1684,N_24226,N_23841);
nor UO_1685 (O_1685,N_23974,N_24440);
and UO_1686 (O_1686,N_24060,N_23772);
nor UO_1687 (O_1687,N_24286,N_24639);
or UO_1688 (O_1688,N_23855,N_24021);
nor UO_1689 (O_1689,N_24221,N_24209);
and UO_1690 (O_1690,N_24943,N_24772);
and UO_1691 (O_1691,N_24352,N_24759);
nand UO_1692 (O_1692,N_24277,N_23968);
and UO_1693 (O_1693,N_24962,N_24291);
and UO_1694 (O_1694,N_24653,N_24854);
nand UO_1695 (O_1695,N_24993,N_24271);
xnor UO_1696 (O_1696,N_24582,N_24296);
xor UO_1697 (O_1697,N_24987,N_24964);
xor UO_1698 (O_1698,N_24449,N_24535);
or UO_1699 (O_1699,N_24921,N_23922);
nor UO_1700 (O_1700,N_23836,N_24531);
xor UO_1701 (O_1701,N_23807,N_24707);
nand UO_1702 (O_1702,N_23757,N_24082);
and UO_1703 (O_1703,N_24490,N_24076);
nand UO_1704 (O_1704,N_24204,N_24023);
xnor UO_1705 (O_1705,N_24283,N_23759);
or UO_1706 (O_1706,N_24226,N_24537);
nand UO_1707 (O_1707,N_23925,N_23943);
nor UO_1708 (O_1708,N_24174,N_24589);
xor UO_1709 (O_1709,N_24818,N_24722);
xnor UO_1710 (O_1710,N_24393,N_24960);
and UO_1711 (O_1711,N_24742,N_24579);
nor UO_1712 (O_1712,N_24159,N_24093);
and UO_1713 (O_1713,N_24574,N_24286);
nand UO_1714 (O_1714,N_24616,N_24516);
and UO_1715 (O_1715,N_24573,N_23966);
xor UO_1716 (O_1716,N_24960,N_24057);
or UO_1717 (O_1717,N_24816,N_24112);
nand UO_1718 (O_1718,N_24849,N_24529);
xor UO_1719 (O_1719,N_24678,N_23889);
and UO_1720 (O_1720,N_24753,N_24138);
nand UO_1721 (O_1721,N_24279,N_24017);
and UO_1722 (O_1722,N_23832,N_24960);
and UO_1723 (O_1723,N_23876,N_24137);
or UO_1724 (O_1724,N_24208,N_24051);
or UO_1725 (O_1725,N_23765,N_23914);
or UO_1726 (O_1726,N_24598,N_24776);
xor UO_1727 (O_1727,N_24020,N_24510);
nand UO_1728 (O_1728,N_24180,N_24531);
nor UO_1729 (O_1729,N_24153,N_24057);
and UO_1730 (O_1730,N_24925,N_24582);
or UO_1731 (O_1731,N_24839,N_23905);
or UO_1732 (O_1732,N_23770,N_24470);
and UO_1733 (O_1733,N_24225,N_24619);
xnor UO_1734 (O_1734,N_24886,N_24684);
xnor UO_1735 (O_1735,N_23806,N_24370);
nor UO_1736 (O_1736,N_23991,N_24311);
nand UO_1737 (O_1737,N_24029,N_23824);
and UO_1738 (O_1738,N_24143,N_24915);
xnor UO_1739 (O_1739,N_24819,N_24720);
xor UO_1740 (O_1740,N_24035,N_24016);
nand UO_1741 (O_1741,N_24358,N_24505);
nand UO_1742 (O_1742,N_24997,N_24778);
xnor UO_1743 (O_1743,N_24479,N_24257);
xor UO_1744 (O_1744,N_23758,N_24819);
and UO_1745 (O_1745,N_23922,N_23796);
nand UO_1746 (O_1746,N_24684,N_24379);
nand UO_1747 (O_1747,N_24559,N_24981);
xor UO_1748 (O_1748,N_23923,N_23840);
xor UO_1749 (O_1749,N_24299,N_23884);
nand UO_1750 (O_1750,N_24787,N_24300);
or UO_1751 (O_1751,N_24143,N_24422);
xor UO_1752 (O_1752,N_24182,N_24272);
nor UO_1753 (O_1753,N_24994,N_23760);
or UO_1754 (O_1754,N_24627,N_24223);
nand UO_1755 (O_1755,N_24166,N_24871);
nor UO_1756 (O_1756,N_24294,N_23970);
xnor UO_1757 (O_1757,N_23915,N_24959);
nand UO_1758 (O_1758,N_24754,N_24498);
nor UO_1759 (O_1759,N_24821,N_24093);
nand UO_1760 (O_1760,N_23855,N_24108);
or UO_1761 (O_1761,N_24618,N_24520);
nor UO_1762 (O_1762,N_23767,N_24088);
and UO_1763 (O_1763,N_24369,N_24026);
and UO_1764 (O_1764,N_23978,N_24705);
xnor UO_1765 (O_1765,N_24480,N_24892);
and UO_1766 (O_1766,N_24738,N_23930);
or UO_1767 (O_1767,N_24688,N_24024);
nor UO_1768 (O_1768,N_24607,N_24962);
xnor UO_1769 (O_1769,N_24181,N_24362);
nor UO_1770 (O_1770,N_24313,N_24209);
xnor UO_1771 (O_1771,N_24464,N_24982);
nor UO_1772 (O_1772,N_24151,N_23969);
xor UO_1773 (O_1773,N_24896,N_24965);
or UO_1774 (O_1774,N_24866,N_24593);
or UO_1775 (O_1775,N_24724,N_24323);
nor UO_1776 (O_1776,N_24824,N_24081);
xnor UO_1777 (O_1777,N_23979,N_24371);
xnor UO_1778 (O_1778,N_24490,N_24070);
and UO_1779 (O_1779,N_24710,N_24328);
or UO_1780 (O_1780,N_24526,N_24337);
or UO_1781 (O_1781,N_24904,N_24618);
and UO_1782 (O_1782,N_24046,N_23769);
or UO_1783 (O_1783,N_24691,N_24715);
and UO_1784 (O_1784,N_24551,N_24137);
nand UO_1785 (O_1785,N_24536,N_23837);
nand UO_1786 (O_1786,N_24366,N_24665);
nand UO_1787 (O_1787,N_24403,N_24195);
xor UO_1788 (O_1788,N_24239,N_24100);
nor UO_1789 (O_1789,N_23978,N_24138);
nand UO_1790 (O_1790,N_24824,N_24904);
xor UO_1791 (O_1791,N_24376,N_24649);
nand UO_1792 (O_1792,N_24190,N_24305);
or UO_1793 (O_1793,N_24525,N_23979);
or UO_1794 (O_1794,N_24281,N_24527);
or UO_1795 (O_1795,N_24275,N_24992);
nor UO_1796 (O_1796,N_23977,N_24376);
nand UO_1797 (O_1797,N_24465,N_23979);
or UO_1798 (O_1798,N_24721,N_24884);
nor UO_1799 (O_1799,N_24777,N_24162);
and UO_1800 (O_1800,N_24560,N_23956);
nor UO_1801 (O_1801,N_24248,N_24711);
xor UO_1802 (O_1802,N_24874,N_24415);
or UO_1803 (O_1803,N_24107,N_24326);
xor UO_1804 (O_1804,N_23894,N_24663);
xnor UO_1805 (O_1805,N_24101,N_24266);
and UO_1806 (O_1806,N_24880,N_24086);
or UO_1807 (O_1807,N_24512,N_24834);
nor UO_1808 (O_1808,N_24414,N_24962);
or UO_1809 (O_1809,N_24502,N_23926);
nand UO_1810 (O_1810,N_24238,N_24273);
nand UO_1811 (O_1811,N_24030,N_24146);
nor UO_1812 (O_1812,N_24015,N_23898);
nand UO_1813 (O_1813,N_24891,N_24238);
and UO_1814 (O_1814,N_24873,N_24039);
nand UO_1815 (O_1815,N_24894,N_23824);
xor UO_1816 (O_1816,N_24530,N_24537);
or UO_1817 (O_1817,N_24669,N_23770);
nand UO_1818 (O_1818,N_24897,N_24710);
xor UO_1819 (O_1819,N_24044,N_24368);
nand UO_1820 (O_1820,N_24941,N_24270);
and UO_1821 (O_1821,N_24724,N_24385);
xor UO_1822 (O_1822,N_24879,N_24711);
and UO_1823 (O_1823,N_24169,N_24902);
nand UO_1824 (O_1824,N_23770,N_24187);
and UO_1825 (O_1825,N_24918,N_23856);
or UO_1826 (O_1826,N_24107,N_24479);
and UO_1827 (O_1827,N_24635,N_24327);
xnor UO_1828 (O_1828,N_24385,N_23874);
nand UO_1829 (O_1829,N_23987,N_24811);
and UO_1830 (O_1830,N_23856,N_24314);
nand UO_1831 (O_1831,N_24426,N_24057);
nand UO_1832 (O_1832,N_23912,N_24805);
xor UO_1833 (O_1833,N_24432,N_24421);
and UO_1834 (O_1834,N_24707,N_24071);
and UO_1835 (O_1835,N_23969,N_24282);
nor UO_1836 (O_1836,N_24576,N_24597);
or UO_1837 (O_1837,N_24690,N_23964);
xor UO_1838 (O_1838,N_23803,N_23757);
xor UO_1839 (O_1839,N_24610,N_24176);
or UO_1840 (O_1840,N_23954,N_23753);
xor UO_1841 (O_1841,N_23929,N_24307);
xnor UO_1842 (O_1842,N_24906,N_24997);
nand UO_1843 (O_1843,N_23814,N_24703);
or UO_1844 (O_1844,N_24373,N_24860);
nor UO_1845 (O_1845,N_24352,N_24304);
and UO_1846 (O_1846,N_24874,N_23854);
and UO_1847 (O_1847,N_24506,N_23903);
nand UO_1848 (O_1848,N_24072,N_24829);
nor UO_1849 (O_1849,N_23778,N_24967);
and UO_1850 (O_1850,N_24430,N_24176);
xnor UO_1851 (O_1851,N_24343,N_24785);
nor UO_1852 (O_1852,N_24562,N_24766);
or UO_1853 (O_1853,N_24310,N_23928);
nand UO_1854 (O_1854,N_24690,N_24556);
nand UO_1855 (O_1855,N_24392,N_24678);
xnor UO_1856 (O_1856,N_24329,N_24249);
or UO_1857 (O_1857,N_24246,N_24359);
nand UO_1858 (O_1858,N_24670,N_24489);
nor UO_1859 (O_1859,N_24179,N_24398);
nor UO_1860 (O_1860,N_24001,N_24864);
xor UO_1861 (O_1861,N_23876,N_24117);
xor UO_1862 (O_1862,N_24574,N_24836);
and UO_1863 (O_1863,N_24882,N_24971);
or UO_1864 (O_1864,N_24338,N_24849);
xor UO_1865 (O_1865,N_24776,N_23753);
and UO_1866 (O_1866,N_24480,N_24856);
nor UO_1867 (O_1867,N_24026,N_23968);
xnor UO_1868 (O_1868,N_23934,N_23936);
or UO_1869 (O_1869,N_24134,N_24957);
or UO_1870 (O_1870,N_23902,N_23801);
or UO_1871 (O_1871,N_24315,N_23974);
nand UO_1872 (O_1872,N_23818,N_23753);
nor UO_1873 (O_1873,N_24219,N_24022);
and UO_1874 (O_1874,N_24375,N_24344);
xnor UO_1875 (O_1875,N_24891,N_24305);
nor UO_1876 (O_1876,N_24472,N_24828);
nand UO_1877 (O_1877,N_24300,N_23798);
nor UO_1878 (O_1878,N_24256,N_24316);
and UO_1879 (O_1879,N_24807,N_24800);
xnor UO_1880 (O_1880,N_23790,N_24193);
nand UO_1881 (O_1881,N_24844,N_24511);
or UO_1882 (O_1882,N_24453,N_24564);
nor UO_1883 (O_1883,N_24688,N_24025);
and UO_1884 (O_1884,N_24550,N_24598);
xnor UO_1885 (O_1885,N_24178,N_24094);
and UO_1886 (O_1886,N_24703,N_24229);
and UO_1887 (O_1887,N_24568,N_24270);
nand UO_1888 (O_1888,N_24399,N_24899);
xor UO_1889 (O_1889,N_24771,N_24568);
nand UO_1890 (O_1890,N_24267,N_24703);
nand UO_1891 (O_1891,N_23949,N_24301);
nand UO_1892 (O_1892,N_24147,N_23764);
or UO_1893 (O_1893,N_23777,N_24377);
nand UO_1894 (O_1894,N_24363,N_24170);
nand UO_1895 (O_1895,N_24408,N_24864);
nand UO_1896 (O_1896,N_24416,N_24371);
and UO_1897 (O_1897,N_24711,N_24222);
nor UO_1898 (O_1898,N_24508,N_24292);
nand UO_1899 (O_1899,N_24133,N_23863);
xnor UO_1900 (O_1900,N_24268,N_23919);
and UO_1901 (O_1901,N_23806,N_24919);
nand UO_1902 (O_1902,N_23787,N_24675);
xor UO_1903 (O_1903,N_24901,N_24872);
xor UO_1904 (O_1904,N_24999,N_24841);
nor UO_1905 (O_1905,N_24623,N_24302);
or UO_1906 (O_1906,N_24182,N_24143);
and UO_1907 (O_1907,N_24235,N_24549);
nand UO_1908 (O_1908,N_24874,N_23789);
nor UO_1909 (O_1909,N_23970,N_24316);
or UO_1910 (O_1910,N_24113,N_24804);
nor UO_1911 (O_1911,N_24049,N_24072);
or UO_1912 (O_1912,N_24533,N_23853);
xor UO_1913 (O_1913,N_23760,N_24760);
and UO_1914 (O_1914,N_24117,N_24356);
and UO_1915 (O_1915,N_23792,N_23901);
nor UO_1916 (O_1916,N_24573,N_24677);
nand UO_1917 (O_1917,N_23838,N_23889);
and UO_1918 (O_1918,N_23918,N_23977);
nor UO_1919 (O_1919,N_24117,N_24445);
nor UO_1920 (O_1920,N_24779,N_24812);
nor UO_1921 (O_1921,N_24370,N_24896);
nor UO_1922 (O_1922,N_24160,N_23791);
nor UO_1923 (O_1923,N_23754,N_24716);
or UO_1924 (O_1924,N_24623,N_24648);
nor UO_1925 (O_1925,N_24231,N_24113);
xnor UO_1926 (O_1926,N_24959,N_24090);
nor UO_1927 (O_1927,N_24331,N_24389);
and UO_1928 (O_1928,N_24008,N_24294);
or UO_1929 (O_1929,N_24485,N_23953);
and UO_1930 (O_1930,N_23956,N_24488);
xnor UO_1931 (O_1931,N_24250,N_23856);
and UO_1932 (O_1932,N_24740,N_24401);
nand UO_1933 (O_1933,N_24305,N_24653);
or UO_1934 (O_1934,N_24255,N_23962);
or UO_1935 (O_1935,N_24109,N_24198);
nand UO_1936 (O_1936,N_24899,N_24001);
nand UO_1937 (O_1937,N_23886,N_23804);
xor UO_1938 (O_1938,N_24641,N_24061);
xnor UO_1939 (O_1939,N_23804,N_24109);
nand UO_1940 (O_1940,N_24261,N_23788);
or UO_1941 (O_1941,N_23871,N_24502);
or UO_1942 (O_1942,N_23927,N_24496);
nand UO_1943 (O_1943,N_24851,N_24700);
and UO_1944 (O_1944,N_23844,N_23793);
nor UO_1945 (O_1945,N_24026,N_24476);
xor UO_1946 (O_1946,N_24677,N_24910);
and UO_1947 (O_1947,N_24925,N_23963);
or UO_1948 (O_1948,N_23786,N_24549);
or UO_1949 (O_1949,N_24787,N_24345);
or UO_1950 (O_1950,N_24747,N_23759);
nor UO_1951 (O_1951,N_24384,N_24216);
and UO_1952 (O_1952,N_23920,N_24736);
or UO_1953 (O_1953,N_24579,N_24190);
nor UO_1954 (O_1954,N_24072,N_23909);
nor UO_1955 (O_1955,N_23990,N_24663);
and UO_1956 (O_1956,N_24739,N_23954);
or UO_1957 (O_1957,N_24849,N_24753);
xnor UO_1958 (O_1958,N_24258,N_23873);
nand UO_1959 (O_1959,N_24891,N_23793);
nand UO_1960 (O_1960,N_24308,N_24320);
or UO_1961 (O_1961,N_23892,N_24003);
xnor UO_1962 (O_1962,N_24275,N_24822);
and UO_1963 (O_1963,N_24920,N_24062);
and UO_1964 (O_1964,N_24680,N_24021);
or UO_1965 (O_1965,N_24621,N_24893);
and UO_1966 (O_1966,N_24696,N_23814);
or UO_1967 (O_1967,N_24919,N_24770);
nand UO_1968 (O_1968,N_24207,N_23930);
nand UO_1969 (O_1969,N_23773,N_24561);
xnor UO_1970 (O_1970,N_24896,N_23821);
and UO_1971 (O_1971,N_24661,N_24626);
and UO_1972 (O_1972,N_24129,N_24446);
xor UO_1973 (O_1973,N_24217,N_24236);
or UO_1974 (O_1974,N_24675,N_23778);
xor UO_1975 (O_1975,N_23815,N_24906);
nand UO_1976 (O_1976,N_24458,N_24577);
or UO_1977 (O_1977,N_23983,N_24106);
xor UO_1978 (O_1978,N_24334,N_24567);
xor UO_1979 (O_1979,N_24453,N_24651);
nor UO_1980 (O_1980,N_24984,N_24489);
xor UO_1981 (O_1981,N_24300,N_24903);
or UO_1982 (O_1982,N_24621,N_23891);
xor UO_1983 (O_1983,N_24077,N_24003);
nand UO_1984 (O_1984,N_24609,N_24754);
or UO_1985 (O_1985,N_23773,N_24022);
xnor UO_1986 (O_1986,N_24165,N_24311);
nand UO_1987 (O_1987,N_24698,N_24259);
xor UO_1988 (O_1988,N_24351,N_24558);
nand UO_1989 (O_1989,N_24234,N_23760);
and UO_1990 (O_1990,N_24031,N_24814);
and UO_1991 (O_1991,N_24899,N_24521);
xnor UO_1992 (O_1992,N_24443,N_24451);
or UO_1993 (O_1993,N_24681,N_24149);
or UO_1994 (O_1994,N_24232,N_24388);
nand UO_1995 (O_1995,N_24349,N_24664);
xor UO_1996 (O_1996,N_23789,N_24993);
and UO_1997 (O_1997,N_24038,N_24517);
and UO_1998 (O_1998,N_24972,N_24061);
nor UO_1999 (O_1999,N_24006,N_23955);
or UO_2000 (O_2000,N_24399,N_23927);
and UO_2001 (O_2001,N_23799,N_24985);
and UO_2002 (O_2002,N_24443,N_23841);
xnor UO_2003 (O_2003,N_24810,N_24787);
or UO_2004 (O_2004,N_24811,N_24014);
or UO_2005 (O_2005,N_24200,N_24686);
xor UO_2006 (O_2006,N_24534,N_23874);
and UO_2007 (O_2007,N_24533,N_24270);
nor UO_2008 (O_2008,N_24500,N_24047);
nand UO_2009 (O_2009,N_24878,N_24301);
and UO_2010 (O_2010,N_24917,N_24362);
nor UO_2011 (O_2011,N_24234,N_24028);
nor UO_2012 (O_2012,N_23988,N_24745);
or UO_2013 (O_2013,N_24796,N_24651);
nand UO_2014 (O_2014,N_24465,N_24898);
and UO_2015 (O_2015,N_24180,N_24633);
and UO_2016 (O_2016,N_24445,N_24265);
xor UO_2017 (O_2017,N_24336,N_24241);
or UO_2018 (O_2018,N_24512,N_24794);
or UO_2019 (O_2019,N_23819,N_24178);
or UO_2020 (O_2020,N_24606,N_23911);
and UO_2021 (O_2021,N_23841,N_24732);
and UO_2022 (O_2022,N_24182,N_24377);
or UO_2023 (O_2023,N_24405,N_23822);
xnor UO_2024 (O_2024,N_24661,N_24856);
or UO_2025 (O_2025,N_24034,N_24966);
and UO_2026 (O_2026,N_24030,N_24878);
or UO_2027 (O_2027,N_24408,N_24564);
nor UO_2028 (O_2028,N_24558,N_24693);
xor UO_2029 (O_2029,N_24936,N_24864);
or UO_2030 (O_2030,N_24500,N_24041);
nor UO_2031 (O_2031,N_24717,N_24199);
nand UO_2032 (O_2032,N_23763,N_24241);
nor UO_2033 (O_2033,N_24985,N_24061);
xor UO_2034 (O_2034,N_23801,N_24900);
xnor UO_2035 (O_2035,N_23997,N_24883);
or UO_2036 (O_2036,N_24015,N_23838);
xor UO_2037 (O_2037,N_24974,N_23877);
nor UO_2038 (O_2038,N_23850,N_23838);
xnor UO_2039 (O_2039,N_24546,N_24511);
or UO_2040 (O_2040,N_24554,N_24644);
and UO_2041 (O_2041,N_24865,N_24027);
and UO_2042 (O_2042,N_23765,N_23931);
xnor UO_2043 (O_2043,N_24883,N_24186);
or UO_2044 (O_2044,N_23800,N_24551);
nor UO_2045 (O_2045,N_24009,N_24833);
nand UO_2046 (O_2046,N_23974,N_24065);
nor UO_2047 (O_2047,N_24124,N_24267);
or UO_2048 (O_2048,N_24552,N_24989);
nor UO_2049 (O_2049,N_24210,N_24344);
and UO_2050 (O_2050,N_23967,N_23949);
or UO_2051 (O_2051,N_23931,N_24473);
nand UO_2052 (O_2052,N_24992,N_24512);
and UO_2053 (O_2053,N_23937,N_23954);
nor UO_2054 (O_2054,N_24861,N_24929);
and UO_2055 (O_2055,N_24628,N_24872);
nand UO_2056 (O_2056,N_23770,N_24014);
nand UO_2057 (O_2057,N_23884,N_24688);
xor UO_2058 (O_2058,N_24022,N_24080);
xnor UO_2059 (O_2059,N_24217,N_24119);
and UO_2060 (O_2060,N_24989,N_24071);
nor UO_2061 (O_2061,N_24537,N_24278);
or UO_2062 (O_2062,N_24568,N_24945);
nand UO_2063 (O_2063,N_24338,N_24003);
nor UO_2064 (O_2064,N_24837,N_24131);
nor UO_2065 (O_2065,N_24001,N_24530);
or UO_2066 (O_2066,N_24433,N_24877);
xnor UO_2067 (O_2067,N_24945,N_24890);
and UO_2068 (O_2068,N_24831,N_24883);
nor UO_2069 (O_2069,N_24852,N_24725);
and UO_2070 (O_2070,N_24133,N_23994);
nor UO_2071 (O_2071,N_24754,N_24020);
xor UO_2072 (O_2072,N_24681,N_23974);
or UO_2073 (O_2073,N_24484,N_24594);
nor UO_2074 (O_2074,N_24745,N_23756);
or UO_2075 (O_2075,N_24685,N_24120);
or UO_2076 (O_2076,N_23893,N_24408);
xnor UO_2077 (O_2077,N_24379,N_24770);
nand UO_2078 (O_2078,N_24414,N_24357);
xnor UO_2079 (O_2079,N_24451,N_24895);
nor UO_2080 (O_2080,N_24368,N_23839);
nor UO_2081 (O_2081,N_24732,N_24112);
nor UO_2082 (O_2082,N_23975,N_23869);
xnor UO_2083 (O_2083,N_24901,N_24322);
nand UO_2084 (O_2084,N_24793,N_24448);
nand UO_2085 (O_2085,N_24932,N_24702);
or UO_2086 (O_2086,N_24777,N_23911);
nand UO_2087 (O_2087,N_24210,N_24634);
nor UO_2088 (O_2088,N_24839,N_24427);
nand UO_2089 (O_2089,N_24052,N_24392);
nand UO_2090 (O_2090,N_24028,N_24943);
nand UO_2091 (O_2091,N_24610,N_24196);
nor UO_2092 (O_2092,N_24714,N_24571);
and UO_2093 (O_2093,N_24347,N_24018);
or UO_2094 (O_2094,N_24629,N_23787);
and UO_2095 (O_2095,N_23788,N_24251);
or UO_2096 (O_2096,N_23822,N_24594);
xnor UO_2097 (O_2097,N_24129,N_24093);
nor UO_2098 (O_2098,N_24468,N_24392);
nor UO_2099 (O_2099,N_24209,N_24401);
nand UO_2100 (O_2100,N_24862,N_24502);
nand UO_2101 (O_2101,N_23770,N_24143);
nor UO_2102 (O_2102,N_24431,N_24436);
nor UO_2103 (O_2103,N_23916,N_23988);
nor UO_2104 (O_2104,N_24717,N_24381);
nand UO_2105 (O_2105,N_24660,N_24803);
xnor UO_2106 (O_2106,N_24235,N_23921);
nor UO_2107 (O_2107,N_24302,N_24635);
xor UO_2108 (O_2108,N_23799,N_24803);
nor UO_2109 (O_2109,N_24205,N_24161);
or UO_2110 (O_2110,N_24851,N_23947);
xor UO_2111 (O_2111,N_24096,N_24636);
and UO_2112 (O_2112,N_24975,N_24457);
and UO_2113 (O_2113,N_23769,N_24693);
nor UO_2114 (O_2114,N_23757,N_24544);
nor UO_2115 (O_2115,N_24228,N_24852);
xnor UO_2116 (O_2116,N_24223,N_24071);
nor UO_2117 (O_2117,N_24286,N_23779);
and UO_2118 (O_2118,N_24286,N_23842);
or UO_2119 (O_2119,N_24979,N_24660);
or UO_2120 (O_2120,N_24527,N_23980);
and UO_2121 (O_2121,N_24986,N_24555);
xnor UO_2122 (O_2122,N_24313,N_24280);
and UO_2123 (O_2123,N_23902,N_24643);
xor UO_2124 (O_2124,N_24158,N_24396);
nand UO_2125 (O_2125,N_24143,N_24175);
nor UO_2126 (O_2126,N_24368,N_24424);
nor UO_2127 (O_2127,N_24026,N_24255);
xnor UO_2128 (O_2128,N_23758,N_23838);
and UO_2129 (O_2129,N_24226,N_24971);
or UO_2130 (O_2130,N_23775,N_24002);
nand UO_2131 (O_2131,N_23953,N_24082);
nor UO_2132 (O_2132,N_23951,N_24835);
xnor UO_2133 (O_2133,N_24265,N_24491);
and UO_2134 (O_2134,N_24727,N_24206);
and UO_2135 (O_2135,N_24618,N_24340);
nor UO_2136 (O_2136,N_23820,N_24481);
nand UO_2137 (O_2137,N_24441,N_24514);
nor UO_2138 (O_2138,N_24611,N_24066);
nand UO_2139 (O_2139,N_24519,N_24791);
nor UO_2140 (O_2140,N_24908,N_24623);
nor UO_2141 (O_2141,N_23897,N_24552);
nand UO_2142 (O_2142,N_24625,N_24439);
or UO_2143 (O_2143,N_24806,N_24692);
and UO_2144 (O_2144,N_23802,N_23945);
xor UO_2145 (O_2145,N_24114,N_23968);
xnor UO_2146 (O_2146,N_24520,N_24410);
and UO_2147 (O_2147,N_24920,N_24100);
and UO_2148 (O_2148,N_24029,N_24564);
xnor UO_2149 (O_2149,N_24265,N_24765);
nor UO_2150 (O_2150,N_24035,N_24737);
nand UO_2151 (O_2151,N_24820,N_24962);
xnor UO_2152 (O_2152,N_24595,N_24950);
and UO_2153 (O_2153,N_24818,N_24977);
nor UO_2154 (O_2154,N_24000,N_23770);
and UO_2155 (O_2155,N_24968,N_24514);
and UO_2156 (O_2156,N_24348,N_24055);
nor UO_2157 (O_2157,N_24011,N_24579);
or UO_2158 (O_2158,N_24553,N_24594);
xor UO_2159 (O_2159,N_23980,N_23905);
nor UO_2160 (O_2160,N_24382,N_23862);
or UO_2161 (O_2161,N_24461,N_24886);
xnor UO_2162 (O_2162,N_23889,N_24087);
nand UO_2163 (O_2163,N_23901,N_23880);
xor UO_2164 (O_2164,N_24329,N_24834);
or UO_2165 (O_2165,N_24819,N_24673);
and UO_2166 (O_2166,N_24171,N_23876);
nand UO_2167 (O_2167,N_24097,N_24954);
nand UO_2168 (O_2168,N_24243,N_23965);
nand UO_2169 (O_2169,N_24956,N_24870);
and UO_2170 (O_2170,N_24903,N_24057);
xor UO_2171 (O_2171,N_24735,N_24104);
xor UO_2172 (O_2172,N_24493,N_23970);
or UO_2173 (O_2173,N_24363,N_24627);
and UO_2174 (O_2174,N_24976,N_24059);
or UO_2175 (O_2175,N_24865,N_24018);
xor UO_2176 (O_2176,N_24851,N_24078);
nor UO_2177 (O_2177,N_24540,N_24126);
or UO_2178 (O_2178,N_24087,N_23902);
xnor UO_2179 (O_2179,N_24882,N_24122);
or UO_2180 (O_2180,N_24267,N_24556);
nor UO_2181 (O_2181,N_24926,N_23924);
nand UO_2182 (O_2182,N_24253,N_24994);
xor UO_2183 (O_2183,N_24969,N_24052);
or UO_2184 (O_2184,N_23935,N_24725);
and UO_2185 (O_2185,N_24094,N_24292);
or UO_2186 (O_2186,N_24506,N_23982);
xor UO_2187 (O_2187,N_24193,N_24157);
and UO_2188 (O_2188,N_23826,N_24048);
xnor UO_2189 (O_2189,N_24772,N_24901);
or UO_2190 (O_2190,N_24939,N_24977);
nand UO_2191 (O_2191,N_24206,N_23873);
nor UO_2192 (O_2192,N_23879,N_24424);
or UO_2193 (O_2193,N_24842,N_24402);
nor UO_2194 (O_2194,N_23766,N_24050);
nor UO_2195 (O_2195,N_23993,N_24920);
or UO_2196 (O_2196,N_24629,N_24544);
and UO_2197 (O_2197,N_24308,N_24458);
nand UO_2198 (O_2198,N_24033,N_24637);
nand UO_2199 (O_2199,N_24203,N_24351);
or UO_2200 (O_2200,N_24448,N_24919);
nand UO_2201 (O_2201,N_24245,N_24720);
and UO_2202 (O_2202,N_24656,N_23867);
nand UO_2203 (O_2203,N_24258,N_23864);
or UO_2204 (O_2204,N_24935,N_24575);
nand UO_2205 (O_2205,N_24638,N_23969);
nand UO_2206 (O_2206,N_24584,N_24238);
and UO_2207 (O_2207,N_24679,N_23843);
and UO_2208 (O_2208,N_23834,N_24460);
or UO_2209 (O_2209,N_24840,N_24209);
nand UO_2210 (O_2210,N_24859,N_24927);
nand UO_2211 (O_2211,N_24177,N_24672);
or UO_2212 (O_2212,N_24616,N_24340);
and UO_2213 (O_2213,N_24384,N_24925);
nor UO_2214 (O_2214,N_24263,N_24118);
or UO_2215 (O_2215,N_24870,N_24478);
nand UO_2216 (O_2216,N_24478,N_24058);
nor UO_2217 (O_2217,N_24695,N_24990);
nor UO_2218 (O_2218,N_24423,N_24441);
nor UO_2219 (O_2219,N_24575,N_24546);
and UO_2220 (O_2220,N_24634,N_24003);
xor UO_2221 (O_2221,N_24738,N_24674);
nand UO_2222 (O_2222,N_24456,N_24798);
xnor UO_2223 (O_2223,N_24892,N_23790);
nand UO_2224 (O_2224,N_24439,N_23768);
or UO_2225 (O_2225,N_24299,N_24105);
or UO_2226 (O_2226,N_24399,N_23900);
or UO_2227 (O_2227,N_24374,N_24119);
and UO_2228 (O_2228,N_23833,N_23850);
nand UO_2229 (O_2229,N_24190,N_24526);
nor UO_2230 (O_2230,N_24587,N_24253);
nand UO_2231 (O_2231,N_24560,N_24732);
or UO_2232 (O_2232,N_24081,N_24578);
and UO_2233 (O_2233,N_23840,N_24453);
and UO_2234 (O_2234,N_24472,N_24523);
nor UO_2235 (O_2235,N_24542,N_24961);
nand UO_2236 (O_2236,N_24534,N_24688);
xnor UO_2237 (O_2237,N_24105,N_24829);
xor UO_2238 (O_2238,N_24507,N_24024);
nor UO_2239 (O_2239,N_24320,N_24583);
and UO_2240 (O_2240,N_24136,N_24903);
nor UO_2241 (O_2241,N_23817,N_24802);
nand UO_2242 (O_2242,N_23868,N_24351);
xnor UO_2243 (O_2243,N_24867,N_24969);
nand UO_2244 (O_2244,N_23788,N_23897);
nand UO_2245 (O_2245,N_24005,N_24246);
xor UO_2246 (O_2246,N_23778,N_24660);
xnor UO_2247 (O_2247,N_24299,N_24231);
nor UO_2248 (O_2248,N_24761,N_24092);
and UO_2249 (O_2249,N_24634,N_23846);
or UO_2250 (O_2250,N_24018,N_24122);
nand UO_2251 (O_2251,N_24181,N_24648);
or UO_2252 (O_2252,N_23856,N_24797);
and UO_2253 (O_2253,N_24335,N_24353);
nor UO_2254 (O_2254,N_23966,N_23980);
nor UO_2255 (O_2255,N_24034,N_24710);
xnor UO_2256 (O_2256,N_24561,N_24031);
nor UO_2257 (O_2257,N_23968,N_24715);
nor UO_2258 (O_2258,N_24698,N_23754);
xor UO_2259 (O_2259,N_23903,N_23976);
nand UO_2260 (O_2260,N_24966,N_24956);
or UO_2261 (O_2261,N_24608,N_24741);
nor UO_2262 (O_2262,N_24444,N_24257);
nand UO_2263 (O_2263,N_24008,N_24254);
and UO_2264 (O_2264,N_24765,N_24107);
nand UO_2265 (O_2265,N_24188,N_24960);
and UO_2266 (O_2266,N_23905,N_24475);
or UO_2267 (O_2267,N_24374,N_24881);
or UO_2268 (O_2268,N_23955,N_24280);
and UO_2269 (O_2269,N_24682,N_24912);
nand UO_2270 (O_2270,N_24966,N_24130);
xor UO_2271 (O_2271,N_24757,N_23832);
nand UO_2272 (O_2272,N_23958,N_24075);
or UO_2273 (O_2273,N_24389,N_24480);
xnor UO_2274 (O_2274,N_24841,N_24461);
nand UO_2275 (O_2275,N_24468,N_24424);
xnor UO_2276 (O_2276,N_24406,N_23845);
or UO_2277 (O_2277,N_24899,N_24610);
and UO_2278 (O_2278,N_24764,N_24028);
nand UO_2279 (O_2279,N_24358,N_23761);
nor UO_2280 (O_2280,N_24133,N_23911);
and UO_2281 (O_2281,N_24920,N_24957);
nand UO_2282 (O_2282,N_24498,N_24015);
and UO_2283 (O_2283,N_23881,N_24888);
nor UO_2284 (O_2284,N_24066,N_23924);
xor UO_2285 (O_2285,N_24743,N_24150);
nand UO_2286 (O_2286,N_24432,N_23975);
or UO_2287 (O_2287,N_24812,N_24940);
nand UO_2288 (O_2288,N_24970,N_24176);
or UO_2289 (O_2289,N_24264,N_24403);
nand UO_2290 (O_2290,N_24904,N_24136);
and UO_2291 (O_2291,N_23799,N_23897);
xor UO_2292 (O_2292,N_24485,N_24875);
xnor UO_2293 (O_2293,N_24519,N_24530);
xnor UO_2294 (O_2294,N_24935,N_24901);
or UO_2295 (O_2295,N_23993,N_24173);
nor UO_2296 (O_2296,N_23835,N_24864);
nor UO_2297 (O_2297,N_24221,N_24331);
nand UO_2298 (O_2298,N_23986,N_23947);
nand UO_2299 (O_2299,N_24684,N_24119);
xor UO_2300 (O_2300,N_23866,N_24166);
or UO_2301 (O_2301,N_24102,N_24079);
nor UO_2302 (O_2302,N_24751,N_23910);
or UO_2303 (O_2303,N_24228,N_24272);
or UO_2304 (O_2304,N_23803,N_24909);
or UO_2305 (O_2305,N_24352,N_24232);
or UO_2306 (O_2306,N_24384,N_23786);
and UO_2307 (O_2307,N_24282,N_24646);
nor UO_2308 (O_2308,N_23808,N_24978);
nor UO_2309 (O_2309,N_24888,N_24046);
nor UO_2310 (O_2310,N_24552,N_24531);
nand UO_2311 (O_2311,N_24462,N_24530);
nor UO_2312 (O_2312,N_24680,N_24711);
nand UO_2313 (O_2313,N_24654,N_23802);
and UO_2314 (O_2314,N_24823,N_24709);
and UO_2315 (O_2315,N_24724,N_24408);
or UO_2316 (O_2316,N_23814,N_24321);
nor UO_2317 (O_2317,N_24370,N_24740);
nor UO_2318 (O_2318,N_24216,N_24291);
or UO_2319 (O_2319,N_23772,N_24730);
and UO_2320 (O_2320,N_24240,N_24473);
nor UO_2321 (O_2321,N_24929,N_24578);
xor UO_2322 (O_2322,N_23998,N_23902);
or UO_2323 (O_2323,N_23850,N_24359);
nand UO_2324 (O_2324,N_24969,N_24671);
nor UO_2325 (O_2325,N_24374,N_24045);
xor UO_2326 (O_2326,N_24067,N_24910);
and UO_2327 (O_2327,N_23948,N_24534);
or UO_2328 (O_2328,N_23822,N_23823);
nand UO_2329 (O_2329,N_24931,N_24609);
nor UO_2330 (O_2330,N_24303,N_23903);
xor UO_2331 (O_2331,N_24323,N_24627);
xor UO_2332 (O_2332,N_24136,N_24687);
nand UO_2333 (O_2333,N_24421,N_24746);
xor UO_2334 (O_2334,N_24277,N_24983);
and UO_2335 (O_2335,N_24406,N_24409);
or UO_2336 (O_2336,N_23936,N_24428);
and UO_2337 (O_2337,N_23830,N_23752);
nor UO_2338 (O_2338,N_24471,N_23892);
and UO_2339 (O_2339,N_24620,N_24700);
nor UO_2340 (O_2340,N_23822,N_24171);
and UO_2341 (O_2341,N_24456,N_24360);
or UO_2342 (O_2342,N_24001,N_24263);
nor UO_2343 (O_2343,N_24486,N_24393);
or UO_2344 (O_2344,N_24909,N_23991);
or UO_2345 (O_2345,N_24331,N_24141);
or UO_2346 (O_2346,N_24118,N_24516);
or UO_2347 (O_2347,N_24832,N_24624);
nor UO_2348 (O_2348,N_23874,N_24942);
nor UO_2349 (O_2349,N_24749,N_23776);
or UO_2350 (O_2350,N_23980,N_24318);
and UO_2351 (O_2351,N_24458,N_24647);
nand UO_2352 (O_2352,N_24920,N_24263);
xor UO_2353 (O_2353,N_24826,N_24201);
and UO_2354 (O_2354,N_24635,N_24392);
xor UO_2355 (O_2355,N_24901,N_24018);
xnor UO_2356 (O_2356,N_24220,N_24335);
and UO_2357 (O_2357,N_23757,N_23985);
xor UO_2358 (O_2358,N_24300,N_24548);
nor UO_2359 (O_2359,N_24264,N_24301);
nor UO_2360 (O_2360,N_24931,N_24364);
or UO_2361 (O_2361,N_24042,N_24540);
xor UO_2362 (O_2362,N_23872,N_24923);
nor UO_2363 (O_2363,N_24863,N_24299);
nor UO_2364 (O_2364,N_24263,N_24757);
xnor UO_2365 (O_2365,N_24325,N_24428);
or UO_2366 (O_2366,N_24973,N_24310);
nand UO_2367 (O_2367,N_24158,N_23751);
xor UO_2368 (O_2368,N_24341,N_23942);
xnor UO_2369 (O_2369,N_24579,N_23976);
nor UO_2370 (O_2370,N_24155,N_23755);
or UO_2371 (O_2371,N_23873,N_24378);
xor UO_2372 (O_2372,N_24698,N_24210);
and UO_2373 (O_2373,N_24159,N_23803);
nand UO_2374 (O_2374,N_24960,N_24298);
or UO_2375 (O_2375,N_24445,N_24083);
or UO_2376 (O_2376,N_24713,N_24949);
nor UO_2377 (O_2377,N_23872,N_24215);
and UO_2378 (O_2378,N_24790,N_24171);
nand UO_2379 (O_2379,N_24744,N_24435);
nor UO_2380 (O_2380,N_23762,N_23979);
nand UO_2381 (O_2381,N_24604,N_24354);
and UO_2382 (O_2382,N_24014,N_23915);
xnor UO_2383 (O_2383,N_23828,N_24362);
xnor UO_2384 (O_2384,N_24626,N_24433);
or UO_2385 (O_2385,N_24665,N_24624);
and UO_2386 (O_2386,N_24325,N_24328);
or UO_2387 (O_2387,N_24346,N_24806);
or UO_2388 (O_2388,N_24133,N_24023);
and UO_2389 (O_2389,N_24750,N_24379);
and UO_2390 (O_2390,N_24386,N_24399);
nor UO_2391 (O_2391,N_24623,N_24807);
xor UO_2392 (O_2392,N_24541,N_24447);
or UO_2393 (O_2393,N_24582,N_23943);
and UO_2394 (O_2394,N_24642,N_24215);
xor UO_2395 (O_2395,N_24972,N_24563);
nor UO_2396 (O_2396,N_24922,N_23957);
nand UO_2397 (O_2397,N_24614,N_24676);
or UO_2398 (O_2398,N_24378,N_24002);
nand UO_2399 (O_2399,N_24607,N_24747);
nor UO_2400 (O_2400,N_24607,N_24440);
nor UO_2401 (O_2401,N_24092,N_23884);
xnor UO_2402 (O_2402,N_24243,N_24425);
and UO_2403 (O_2403,N_23870,N_24063);
and UO_2404 (O_2404,N_24623,N_24319);
or UO_2405 (O_2405,N_24721,N_23914);
xor UO_2406 (O_2406,N_24956,N_24070);
xor UO_2407 (O_2407,N_24141,N_24222);
xor UO_2408 (O_2408,N_24129,N_24437);
and UO_2409 (O_2409,N_24017,N_24878);
and UO_2410 (O_2410,N_24833,N_24559);
and UO_2411 (O_2411,N_24178,N_24511);
or UO_2412 (O_2412,N_24993,N_23992);
and UO_2413 (O_2413,N_24795,N_23765);
nor UO_2414 (O_2414,N_24212,N_24832);
or UO_2415 (O_2415,N_24652,N_23980);
and UO_2416 (O_2416,N_23906,N_24080);
xnor UO_2417 (O_2417,N_24868,N_23846);
xor UO_2418 (O_2418,N_24394,N_24311);
nand UO_2419 (O_2419,N_23972,N_24875);
or UO_2420 (O_2420,N_24870,N_23767);
or UO_2421 (O_2421,N_24363,N_24260);
xor UO_2422 (O_2422,N_24145,N_24046);
nand UO_2423 (O_2423,N_24858,N_24067);
and UO_2424 (O_2424,N_24860,N_24589);
nand UO_2425 (O_2425,N_24403,N_24254);
nor UO_2426 (O_2426,N_24967,N_24086);
and UO_2427 (O_2427,N_24818,N_23968);
or UO_2428 (O_2428,N_23882,N_24511);
nor UO_2429 (O_2429,N_23849,N_23933);
nand UO_2430 (O_2430,N_24064,N_24257);
nor UO_2431 (O_2431,N_23879,N_23987);
nand UO_2432 (O_2432,N_24407,N_24580);
xnor UO_2433 (O_2433,N_24146,N_23772);
or UO_2434 (O_2434,N_24812,N_23856);
and UO_2435 (O_2435,N_23775,N_24938);
or UO_2436 (O_2436,N_24882,N_24801);
xor UO_2437 (O_2437,N_24485,N_24005);
or UO_2438 (O_2438,N_23985,N_24974);
or UO_2439 (O_2439,N_24964,N_24906);
xnor UO_2440 (O_2440,N_24361,N_24956);
nand UO_2441 (O_2441,N_23900,N_24017);
nor UO_2442 (O_2442,N_23816,N_24246);
and UO_2443 (O_2443,N_24868,N_24489);
nand UO_2444 (O_2444,N_24635,N_23795);
xnor UO_2445 (O_2445,N_24076,N_24252);
and UO_2446 (O_2446,N_23768,N_24295);
nand UO_2447 (O_2447,N_23817,N_23826);
xor UO_2448 (O_2448,N_23920,N_24241);
xor UO_2449 (O_2449,N_24623,N_24504);
or UO_2450 (O_2450,N_24916,N_24262);
and UO_2451 (O_2451,N_24523,N_23839);
or UO_2452 (O_2452,N_24095,N_24298);
or UO_2453 (O_2453,N_24276,N_24671);
nor UO_2454 (O_2454,N_24859,N_24880);
and UO_2455 (O_2455,N_24749,N_23806);
and UO_2456 (O_2456,N_24255,N_24059);
xnor UO_2457 (O_2457,N_24040,N_23884);
nor UO_2458 (O_2458,N_24894,N_24758);
xor UO_2459 (O_2459,N_23909,N_23833);
or UO_2460 (O_2460,N_24447,N_24126);
xor UO_2461 (O_2461,N_24660,N_24812);
and UO_2462 (O_2462,N_24746,N_24512);
xnor UO_2463 (O_2463,N_24438,N_23912);
nor UO_2464 (O_2464,N_23926,N_23880);
and UO_2465 (O_2465,N_24838,N_24829);
or UO_2466 (O_2466,N_24585,N_24395);
and UO_2467 (O_2467,N_23777,N_24901);
and UO_2468 (O_2468,N_23898,N_24283);
xor UO_2469 (O_2469,N_24723,N_24688);
nand UO_2470 (O_2470,N_24669,N_24061);
nand UO_2471 (O_2471,N_24747,N_24059);
and UO_2472 (O_2472,N_24289,N_24424);
xnor UO_2473 (O_2473,N_24165,N_24201);
or UO_2474 (O_2474,N_24639,N_24377);
nand UO_2475 (O_2475,N_24266,N_24340);
and UO_2476 (O_2476,N_24360,N_24890);
nor UO_2477 (O_2477,N_23932,N_24785);
nor UO_2478 (O_2478,N_24959,N_23986);
or UO_2479 (O_2479,N_24641,N_24894);
and UO_2480 (O_2480,N_23896,N_24454);
xnor UO_2481 (O_2481,N_24074,N_24403);
or UO_2482 (O_2482,N_24946,N_24943);
nor UO_2483 (O_2483,N_24099,N_24598);
nand UO_2484 (O_2484,N_24594,N_24804);
or UO_2485 (O_2485,N_24693,N_24334);
nor UO_2486 (O_2486,N_24106,N_24813);
or UO_2487 (O_2487,N_23788,N_24453);
and UO_2488 (O_2488,N_24010,N_23872);
nand UO_2489 (O_2489,N_24854,N_24804);
and UO_2490 (O_2490,N_23884,N_24488);
and UO_2491 (O_2491,N_23896,N_24938);
xnor UO_2492 (O_2492,N_24966,N_24982);
and UO_2493 (O_2493,N_24373,N_24770);
xor UO_2494 (O_2494,N_23813,N_24260);
and UO_2495 (O_2495,N_23859,N_24163);
and UO_2496 (O_2496,N_24276,N_24490);
xor UO_2497 (O_2497,N_24411,N_24709);
nor UO_2498 (O_2498,N_24779,N_23902);
and UO_2499 (O_2499,N_24659,N_24886);
or UO_2500 (O_2500,N_24444,N_23896);
nand UO_2501 (O_2501,N_24553,N_23989);
and UO_2502 (O_2502,N_24141,N_23790);
xnor UO_2503 (O_2503,N_24616,N_24525);
or UO_2504 (O_2504,N_24845,N_24905);
or UO_2505 (O_2505,N_23919,N_24912);
xor UO_2506 (O_2506,N_24228,N_24793);
or UO_2507 (O_2507,N_24711,N_24872);
and UO_2508 (O_2508,N_24025,N_24987);
xor UO_2509 (O_2509,N_24521,N_24378);
and UO_2510 (O_2510,N_23785,N_24789);
nor UO_2511 (O_2511,N_24937,N_24465);
xnor UO_2512 (O_2512,N_24151,N_24418);
xnor UO_2513 (O_2513,N_24620,N_24040);
or UO_2514 (O_2514,N_24304,N_24142);
or UO_2515 (O_2515,N_24040,N_24996);
xor UO_2516 (O_2516,N_24882,N_24559);
and UO_2517 (O_2517,N_23930,N_23895);
nor UO_2518 (O_2518,N_24009,N_24680);
and UO_2519 (O_2519,N_24049,N_24985);
nor UO_2520 (O_2520,N_24894,N_23957);
and UO_2521 (O_2521,N_24919,N_24663);
nand UO_2522 (O_2522,N_23974,N_24026);
and UO_2523 (O_2523,N_23907,N_24633);
and UO_2524 (O_2524,N_23938,N_24252);
xor UO_2525 (O_2525,N_24147,N_24582);
nand UO_2526 (O_2526,N_24575,N_24535);
nor UO_2527 (O_2527,N_23935,N_23956);
or UO_2528 (O_2528,N_24715,N_24054);
or UO_2529 (O_2529,N_24518,N_24433);
nand UO_2530 (O_2530,N_24262,N_23959);
nand UO_2531 (O_2531,N_24771,N_24159);
nor UO_2532 (O_2532,N_24360,N_24937);
nor UO_2533 (O_2533,N_24151,N_24273);
nand UO_2534 (O_2534,N_24709,N_24747);
nor UO_2535 (O_2535,N_24153,N_24303);
nor UO_2536 (O_2536,N_24587,N_23754);
nand UO_2537 (O_2537,N_23780,N_24120);
nor UO_2538 (O_2538,N_24709,N_24335);
nor UO_2539 (O_2539,N_24427,N_24878);
or UO_2540 (O_2540,N_24962,N_23752);
or UO_2541 (O_2541,N_24858,N_24326);
nand UO_2542 (O_2542,N_23987,N_23989);
or UO_2543 (O_2543,N_24968,N_24751);
nand UO_2544 (O_2544,N_23843,N_24404);
nand UO_2545 (O_2545,N_24739,N_24406);
xnor UO_2546 (O_2546,N_23811,N_23750);
xor UO_2547 (O_2547,N_24883,N_24198);
nand UO_2548 (O_2548,N_24546,N_24492);
nand UO_2549 (O_2549,N_24297,N_24951);
and UO_2550 (O_2550,N_23864,N_24044);
nor UO_2551 (O_2551,N_24739,N_23971);
nor UO_2552 (O_2552,N_24040,N_24462);
nor UO_2553 (O_2553,N_24016,N_23849);
nand UO_2554 (O_2554,N_24413,N_23800);
or UO_2555 (O_2555,N_23782,N_23945);
or UO_2556 (O_2556,N_24378,N_24743);
xor UO_2557 (O_2557,N_23921,N_24649);
or UO_2558 (O_2558,N_24341,N_24769);
or UO_2559 (O_2559,N_24025,N_24595);
or UO_2560 (O_2560,N_24903,N_23976);
nor UO_2561 (O_2561,N_24466,N_24653);
xnor UO_2562 (O_2562,N_23869,N_24306);
xnor UO_2563 (O_2563,N_24926,N_23911);
xor UO_2564 (O_2564,N_24111,N_24385);
and UO_2565 (O_2565,N_24869,N_23867);
and UO_2566 (O_2566,N_24587,N_24527);
nand UO_2567 (O_2567,N_23778,N_24450);
nand UO_2568 (O_2568,N_24877,N_24394);
nand UO_2569 (O_2569,N_23952,N_24014);
or UO_2570 (O_2570,N_24603,N_23976);
nand UO_2571 (O_2571,N_24051,N_24761);
nor UO_2572 (O_2572,N_24715,N_24115);
nand UO_2573 (O_2573,N_24440,N_24117);
nor UO_2574 (O_2574,N_24022,N_24863);
nand UO_2575 (O_2575,N_24310,N_24228);
nor UO_2576 (O_2576,N_24682,N_24177);
nor UO_2577 (O_2577,N_24394,N_24604);
nor UO_2578 (O_2578,N_23768,N_24094);
or UO_2579 (O_2579,N_24734,N_23938);
xor UO_2580 (O_2580,N_24400,N_24066);
nor UO_2581 (O_2581,N_24031,N_24257);
and UO_2582 (O_2582,N_24362,N_24372);
xor UO_2583 (O_2583,N_24771,N_24040);
nor UO_2584 (O_2584,N_24261,N_24969);
nand UO_2585 (O_2585,N_23816,N_24826);
xnor UO_2586 (O_2586,N_24356,N_24813);
nor UO_2587 (O_2587,N_24495,N_24064);
and UO_2588 (O_2588,N_24404,N_24862);
xor UO_2589 (O_2589,N_24762,N_24760);
xnor UO_2590 (O_2590,N_23856,N_24951);
and UO_2591 (O_2591,N_23873,N_23945);
or UO_2592 (O_2592,N_24863,N_24836);
and UO_2593 (O_2593,N_23948,N_24617);
and UO_2594 (O_2594,N_23750,N_24900);
and UO_2595 (O_2595,N_24977,N_24716);
nor UO_2596 (O_2596,N_24823,N_24394);
nand UO_2597 (O_2597,N_24318,N_23799);
nand UO_2598 (O_2598,N_23960,N_24465);
and UO_2599 (O_2599,N_24699,N_24690);
and UO_2600 (O_2600,N_23884,N_23910);
or UO_2601 (O_2601,N_24503,N_24457);
nand UO_2602 (O_2602,N_24812,N_24585);
nor UO_2603 (O_2603,N_24454,N_24807);
nor UO_2604 (O_2604,N_24372,N_24877);
xnor UO_2605 (O_2605,N_23880,N_23881);
or UO_2606 (O_2606,N_24228,N_23990);
and UO_2607 (O_2607,N_24012,N_24449);
nand UO_2608 (O_2608,N_23929,N_24090);
or UO_2609 (O_2609,N_24208,N_23792);
nor UO_2610 (O_2610,N_24476,N_24774);
and UO_2611 (O_2611,N_24560,N_24601);
or UO_2612 (O_2612,N_24291,N_24154);
or UO_2613 (O_2613,N_24632,N_24554);
nor UO_2614 (O_2614,N_24149,N_23954);
or UO_2615 (O_2615,N_24131,N_24333);
and UO_2616 (O_2616,N_24924,N_24667);
nor UO_2617 (O_2617,N_24287,N_24724);
and UO_2618 (O_2618,N_24083,N_23922);
nor UO_2619 (O_2619,N_24208,N_24608);
xnor UO_2620 (O_2620,N_24980,N_24667);
nand UO_2621 (O_2621,N_24190,N_24322);
and UO_2622 (O_2622,N_24710,N_24162);
nand UO_2623 (O_2623,N_24007,N_24468);
or UO_2624 (O_2624,N_24203,N_23896);
and UO_2625 (O_2625,N_23891,N_24616);
and UO_2626 (O_2626,N_24718,N_24765);
and UO_2627 (O_2627,N_24307,N_24699);
and UO_2628 (O_2628,N_24551,N_24692);
nor UO_2629 (O_2629,N_24934,N_24853);
or UO_2630 (O_2630,N_24040,N_24225);
and UO_2631 (O_2631,N_24683,N_24423);
nor UO_2632 (O_2632,N_24585,N_24898);
or UO_2633 (O_2633,N_24192,N_24577);
or UO_2634 (O_2634,N_24192,N_23804);
and UO_2635 (O_2635,N_24194,N_24630);
nand UO_2636 (O_2636,N_24486,N_24290);
xnor UO_2637 (O_2637,N_23757,N_24455);
and UO_2638 (O_2638,N_24314,N_24344);
and UO_2639 (O_2639,N_24412,N_24553);
xor UO_2640 (O_2640,N_24398,N_24334);
and UO_2641 (O_2641,N_23929,N_24940);
or UO_2642 (O_2642,N_23908,N_24477);
xnor UO_2643 (O_2643,N_23970,N_24656);
nand UO_2644 (O_2644,N_24077,N_23879);
nor UO_2645 (O_2645,N_24312,N_24074);
or UO_2646 (O_2646,N_24879,N_23912);
xor UO_2647 (O_2647,N_24171,N_24076);
nor UO_2648 (O_2648,N_24818,N_23762);
nor UO_2649 (O_2649,N_24427,N_24190);
nor UO_2650 (O_2650,N_23867,N_23884);
nor UO_2651 (O_2651,N_24832,N_24434);
nor UO_2652 (O_2652,N_24379,N_23847);
and UO_2653 (O_2653,N_24577,N_24697);
xnor UO_2654 (O_2654,N_24397,N_23868);
nand UO_2655 (O_2655,N_23939,N_24270);
nor UO_2656 (O_2656,N_24539,N_23884);
or UO_2657 (O_2657,N_24375,N_24373);
nor UO_2658 (O_2658,N_24220,N_24630);
xor UO_2659 (O_2659,N_24430,N_23822);
nor UO_2660 (O_2660,N_24883,N_23791);
nor UO_2661 (O_2661,N_24679,N_24633);
or UO_2662 (O_2662,N_24764,N_24221);
nor UO_2663 (O_2663,N_24771,N_23819);
or UO_2664 (O_2664,N_24529,N_24582);
or UO_2665 (O_2665,N_24550,N_24817);
or UO_2666 (O_2666,N_24740,N_24708);
and UO_2667 (O_2667,N_24141,N_24608);
nand UO_2668 (O_2668,N_24439,N_24378);
xnor UO_2669 (O_2669,N_24899,N_24405);
nor UO_2670 (O_2670,N_24028,N_24993);
or UO_2671 (O_2671,N_24724,N_24930);
nor UO_2672 (O_2672,N_23753,N_24670);
and UO_2673 (O_2673,N_24826,N_23955);
nand UO_2674 (O_2674,N_24685,N_23782);
and UO_2675 (O_2675,N_24724,N_23994);
and UO_2676 (O_2676,N_24979,N_24526);
or UO_2677 (O_2677,N_24552,N_23782);
and UO_2678 (O_2678,N_24682,N_24523);
or UO_2679 (O_2679,N_24310,N_24778);
or UO_2680 (O_2680,N_24260,N_23768);
or UO_2681 (O_2681,N_24703,N_24467);
or UO_2682 (O_2682,N_24062,N_24907);
nor UO_2683 (O_2683,N_24651,N_24998);
and UO_2684 (O_2684,N_24750,N_23903);
xor UO_2685 (O_2685,N_24632,N_24661);
and UO_2686 (O_2686,N_24029,N_24359);
nor UO_2687 (O_2687,N_23985,N_24218);
xnor UO_2688 (O_2688,N_23842,N_24611);
nor UO_2689 (O_2689,N_24264,N_24431);
xor UO_2690 (O_2690,N_24537,N_24922);
nand UO_2691 (O_2691,N_24575,N_24959);
xor UO_2692 (O_2692,N_24885,N_24887);
xnor UO_2693 (O_2693,N_24878,N_23804);
nor UO_2694 (O_2694,N_24151,N_24456);
nand UO_2695 (O_2695,N_24265,N_24321);
nor UO_2696 (O_2696,N_24876,N_24292);
or UO_2697 (O_2697,N_24314,N_24829);
and UO_2698 (O_2698,N_24086,N_23766);
nor UO_2699 (O_2699,N_24516,N_23849);
nor UO_2700 (O_2700,N_23977,N_24742);
and UO_2701 (O_2701,N_24190,N_24387);
or UO_2702 (O_2702,N_24359,N_24759);
nor UO_2703 (O_2703,N_24983,N_24434);
nand UO_2704 (O_2704,N_24423,N_24856);
nor UO_2705 (O_2705,N_24182,N_23754);
xnor UO_2706 (O_2706,N_24336,N_24214);
or UO_2707 (O_2707,N_24547,N_24037);
nor UO_2708 (O_2708,N_23849,N_23874);
or UO_2709 (O_2709,N_24886,N_24494);
and UO_2710 (O_2710,N_24777,N_24940);
xnor UO_2711 (O_2711,N_24872,N_24758);
nand UO_2712 (O_2712,N_23982,N_24782);
or UO_2713 (O_2713,N_24665,N_24282);
xnor UO_2714 (O_2714,N_24785,N_24372);
xnor UO_2715 (O_2715,N_23851,N_24836);
nor UO_2716 (O_2716,N_24154,N_23844);
and UO_2717 (O_2717,N_24975,N_24301);
nand UO_2718 (O_2718,N_24311,N_23988);
or UO_2719 (O_2719,N_24664,N_24857);
nand UO_2720 (O_2720,N_23908,N_24782);
nand UO_2721 (O_2721,N_24913,N_23839);
xor UO_2722 (O_2722,N_24589,N_23755);
nor UO_2723 (O_2723,N_24007,N_23760);
xnor UO_2724 (O_2724,N_24399,N_24853);
nand UO_2725 (O_2725,N_24817,N_24591);
and UO_2726 (O_2726,N_23906,N_23891);
or UO_2727 (O_2727,N_24530,N_24302);
or UO_2728 (O_2728,N_24373,N_24761);
nor UO_2729 (O_2729,N_24998,N_24939);
or UO_2730 (O_2730,N_24634,N_23781);
nand UO_2731 (O_2731,N_24800,N_23803);
xor UO_2732 (O_2732,N_24171,N_24064);
xnor UO_2733 (O_2733,N_24644,N_24199);
and UO_2734 (O_2734,N_24736,N_24226);
xnor UO_2735 (O_2735,N_24701,N_24222);
nor UO_2736 (O_2736,N_24701,N_24620);
xor UO_2737 (O_2737,N_24931,N_24643);
xor UO_2738 (O_2738,N_24909,N_23872);
xnor UO_2739 (O_2739,N_24467,N_24341);
nand UO_2740 (O_2740,N_24823,N_24490);
xnor UO_2741 (O_2741,N_24581,N_24114);
nand UO_2742 (O_2742,N_23874,N_24308);
xnor UO_2743 (O_2743,N_23973,N_24908);
xnor UO_2744 (O_2744,N_24856,N_24154);
and UO_2745 (O_2745,N_24645,N_23946);
xor UO_2746 (O_2746,N_24957,N_24714);
nor UO_2747 (O_2747,N_24634,N_24459);
nor UO_2748 (O_2748,N_23953,N_23993);
and UO_2749 (O_2749,N_24334,N_24775);
nand UO_2750 (O_2750,N_24211,N_24698);
xor UO_2751 (O_2751,N_24557,N_23850);
xor UO_2752 (O_2752,N_23784,N_24361);
nor UO_2753 (O_2753,N_24631,N_23814);
xor UO_2754 (O_2754,N_24552,N_24804);
nand UO_2755 (O_2755,N_23982,N_23835);
xnor UO_2756 (O_2756,N_24544,N_24819);
nand UO_2757 (O_2757,N_24447,N_24956);
xor UO_2758 (O_2758,N_24077,N_24314);
and UO_2759 (O_2759,N_24393,N_24157);
or UO_2760 (O_2760,N_24198,N_23788);
and UO_2761 (O_2761,N_24854,N_24727);
nor UO_2762 (O_2762,N_24940,N_24922);
nor UO_2763 (O_2763,N_24171,N_24617);
and UO_2764 (O_2764,N_23915,N_23919);
nor UO_2765 (O_2765,N_23875,N_24717);
nand UO_2766 (O_2766,N_23989,N_24627);
nand UO_2767 (O_2767,N_24760,N_24728);
xor UO_2768 (O_2768,N_24850,N_23779);
xnor UO_2769 (O_2769,N_24431,N_23758);
nand UO_2770 (O_2770,N_24472,N_24314);
or UO_2771 (O_2771,N_24119,N_24577);
and UO_2772 (O_2772,N_24835,N_24617);
or UO_2773 (O_2773,N_24925,N_23791);
or UO_2774 (O_2774,N_24360,N_24790);
nor UO_2775 (O_2775,N_24059,N_24333);
nor UO_2776 (O_2776,N_24221,N_24361);
nor UO_2777 (O_2777,N_24197,N_24760);
and UO_2778 (O_2778,N_24968,N_23999);
or UO_2779 (O_2779,N_24496,N_24126);
nand UO_2780 (O_2780,N_23802,N_24890);
xnor UO_2781 (O_2781,N_24857,N_24818);
or UO_2782 (O_2782,N_24900,N_23760);
and UO_2783 (O_2783,N_24277,N_24507);
nand UO_2784 (O_2784,N_24869,N_24681);
and UO_2785 (O_2785,N_23983,N_24935);
or UO_2786 (O_2786,N_24740,N_24227);
nand UO_2787 (O_2787,N_23754,N_24934);
xnor UO_2788 (O_2788,N_24302,N_24907);
and UO_2789 (O_2789,N_24104,N_24118);
or UO_2790 (O_2790,N_23793,N_24579);
xnor UO_2791 (O_2791,N_23831,N_24705);
and UO_2792 (O_2792,N_24585,N_24878);
nand UO_2793 (O_2793,N_24661,N_24810);
nand UO_2794 (O_2794,N_24475,N_24897);
and UO_2795 (O_2795,N_23947,N_24294);
or UO_2796 (O_2796,N_23887,N_24757);
xnor UO_2797 (O_2797,N_23810,N_24109);
or UO_2798 (O_2798,N_24659,N_23840);
nor UO_2799 (O_2799,N_24701,N_23918);
and UO_2800 (O_2800,N_24937,N_24860);
nand UO_2801 (O_2801,N_23906,N_23947);
and UO_2802 (O_2802,N_24139,N_24877);
nor UO_2803 (O_2803,N_23843,N_24476);
nand UO_2804 (O_2804,N_23968,N_23930);
and UO_2805 (O_2805,N_24315,N_24955);
xnor UO_2806 (O_2806,N_24832,N_24990);
nand UO_2807 (O_2807,N_24828,N_24977);
nor UO_2808 (O_2808,N_24948,N_23771);
and UO_2809 (O_2809,N_23883,N_24155);
nand UO_2810 (O_2810,N_24197,N_24390);
xor UO_2811 (O_2811,N_24810,N_24806);
nand UO_2812 (O_2812,N_24111,N_24055);
and UO_2813 (O_2813,N_24270,N_24056);
and UO_2814 (O_2814,N_23909,N_23963);
nor UO_2815 (O_2815,N_24212,N_24782);
or UO_2816 (O_2816,N_24639,N_24832);
nand UO_2817 (O_2817,N_24580,N_23840);
nor UO_2818 (O_2818,N_24490,N_24885);
or UO_2819 (O_2819,N_24346,N_24746);
nand UO_2820 (O_2820,N_24317,N_24899);
nor UO_2821 (O_2821,N_24945,N_24523);
or UO_2822 (O_2822,N_24739,N_24914);
and UO_2823 (O_2823,N_24087,N_24062);
and UO_2824 (O_2824,N_24459,N_24854);
nor UO_2825 (O_2825,N_24746,N_23984);
nor UO_2826 (O_2826,N_24012,N_24289);
and UO_2827 (O_2827,N_24258,N_24173);
or UO_2828 (O_2828,N_24307,N_24925);
nor UO_2829 (O_2829,N_24880,N_24440);
nor UO_2830 (O_2830,N_23936,N_24502);
xnor UO_2831 (O_2831,N_24029,N_24813);
or UO_2832 (O_2832,N_24314,N_24942);
xor UO_2833 (O_2833,N_23902,N_24180);
nor UO_2834 (O_2834,N_24436,N_24319);
xor UO_2835 (O_2835,N_24391,N_24941);
nand UO_2836 (O_2836,N_23975,N_23858);
nand UO_2837 (O_2837,N_24136,N_24775);
and UO_2838 (O_2838,N_24963,N_23968);
and UO_2839 (O_2839,N_24789,N_24722);
and UO_2840 (O_2840,N_24386,N_24475);
or UO_2841 (O_2841,N_24372,N_24294);
xor UO_2842 (O_2842,N_24928,N_24149);
and UO_2843 (O_2843,N_23891,N_24306);
and UO_2844 (O_2844,N_24295,N_24802);
or UO_2845 (O_2845,N_24784,N_23828);
or UO_2846 (O_2846,N_24100,N_24718);
nand UO_2847 (O_2847,N_24221,N_24190);
nand UO_2848 (O_2848,N_24974,N_24746);
nor UO_2849 (O_2849,N_24852,N_24338);
nand UO_2850 (O_2850,N_24478,N_24704);
and UO_2851 (O_2851,N_24926,N_23956);
or UO_2852 (O_2852,N_24467,N_24108);
or UO_2853 (O_2853,N_24996,N_24704);
nand UO_2854 (O_2854,N_24913,N_24536);
nand UO_2855 (O_2855,N_23941,N_23834);
nor UO_2856 (O_2856,N_24747,N_23890);
or UO_2857 (O_2857,N_24838,N_24758);
or UO_2858 (O_2858,N_24955,N_24753);
nand UO_2859 (O_2859,N_24408,N_23992);
xnor UO_2860 (O_2860,N_24559,N_23970);
xor UO_2861 (O_2861,N_24734,N_24066);
or UO_2862 (O_2862,N_23911,N_24307);
or UO_2863 (O_2863,N_24202,N_24890);
and UO_2864 (O_2864,N_24716,N_24256);
nor UO_2865 (O_2865,N_24543,N_24928);
nor UO_2866 (O_2866,N_24582,N_24012);
xnor UO_2867 (O_2867,N_24890,N_24920);
xnor UO_2868 (O_2868,N_24356,N_24508);
xor UO_2869 (O_2869,N_24324,N_24229);
nor UO_2870 (O_2870,N_24112,N_24066);
or UO_2871 (O_2871,N_24977,N_24549);
and UO_2872 (O_2872,N_24100,N_24348);
or UO_2873 (O_2873,N_24963,N_24775);
nor UO_2874 (O_2874,N_23759,N_24712);
nand UO_2875 (O_2875,N_24974,N_24715);
nor UO_2876 (O_2876,N_24635,N_24403);
or UO_2877 (O_2877,N_24484,N_24774);
and UO_2878 (O_2878,N_24185,N_24374);
nand UO_2879 (O_2879,N_23884,N_24098);
nand UO_2880 (O_2880,N_24768,N_24659);
nor UO_2881 (O_2881,N_24300,N_24261);
xnor UO_2882 (O_2882,N_24015,N_24137);
nor UO_2883 (O_2883,N_24247,N_24901);
nor UO_2884 (O_2884,N_23984,N_24009);
and UO_2885 (O_2885,N_24049,N_24689);
and UO_2886 (O_2886,N_24445,N_24499);
xor UO_2887 (O_2887,N_24175,N_24122);
or UO_2888 (O_2888,N_23794,N_24840);
xnor UO_2889 (O_2889,N_24691,N_23951);
nor UO_2890 (O_2890,N_24186,N_24135);
xor UO_2891 (O_2891,N_24859,N_24531);
xor UO_2892 (O_2892,N_24885,N_24469);
and UO_2893 (O_2893,N_24715,N_24576);
nand UO_2894 (O_2894,N_23910,N_23788);
nand UO_2895 (O_2895,N_24410,N_24905);
or UO_2896 (O_2896,N_24926,N_23994);
nor UO_2897 (O_2897,N_24607,N_23883);
nand UO_2898 (O_2898,N_23864,N_24218);
and UO_2899 (O_2899,N_24674,N_24910);
nor UO_2900 (O_2900,N_24728,N_24050);
nor UO_2901 (O_2901,N_23789,N_23806);
or UO_2902 (O_2902,N_23761,N_24265);
and UO_2903 (O_2903,N_24709,N_24627);
nand UO_2904 (O_2904,N_24162,N_24569);
nor UO_2905 (O_2905,N_24830,N_24025);
nand UO_2906 (O_2906,N_24508,N_24249);
xor UO_2907 (O_2907,N_24787,N_24923);
xor UO_2908 (O_2908,N_24801,N_24347);
or UO_2909 (O_2909,N_24571,N_23983);
nor UO_2910 (O_2910,N_24764,N_24281);
and UO_2911 (O_2911,N_23751,N_24620);
or UO_2912 (O_2912,N_24621,N_24943);
and UO_2913 (O_2913,N_24527,N_24145);
xor UO_2914 (O_2914,N_24546,N_24991);
nand UO_2915 (O_2915,N_24931,N_24266);
nor UO_2916 (O_2916,N_24968,N_24453);
nor UO_2917 (O_2917,N_24587,N_24440);
or UO_2918 (O_2918,N_24902,N_24677);
nor UO_2919 (O_2919,N_24267,N_24804);
nand UO_2920 (O_2920,N_24557,N_24782);
and UO_2921 (O_2921,N_24181,N_24226);
xnor UO_2922 (O_2922,N_24483,N_24444);
or UO_2923 (O_2923,N_24561,N_24669);
and UO_2924 (O_2924,N_24866,N_24209);
nand UO_2925 (O_2925,N_23993,N_24354);
xnor UO_2926 (O_2926,N_24596,N_24048);
xor UO_2927 (O_2927,N_24291,N_24879);
nand UO_2928 (O_2928,N_24779,N_23855);
xor UO_2929 (O_2929,N_24515,N_24519);
xnor UO_2930 (O_2930,N_24684,N_23760);
or UO_2931 (O_2931,N_24768,N_24416);
and UO_2932 (O_2932,N_23925,N_24034);
xor UO_2933 (O_2933,N_24285,N_24479);
or UO_2934 (O_2934,N_24911,N_24649);
xnor UO_2935 (O_2935,N_24822,N_24305);
nor UO_2936 (O_2936,N_23941,N_23751);
nand UO_2937 (O_2937,N_23933,N_23814);
and UO_2938 (O_2938,N_24018,N_24198);
nand UO_2939 (O_2939,N_24737,N_24516);
or UO_2940 (O_2940,N_24339,N_24909);
or UO_2941 (O_2941,N_24180,N_24031);
nand UO_2942 (O_2942,N_24023,N_24912);
or UO_2943 (O_2943,N_24973,N_23872);
and UO_2944 (O_2944,N_24615,N_24956);
or UO_2945 (O_2945,N_24244,N_24779);
and UO_2946 (O_2946,N_24440,N_24351);
and UO_2947 (O_2947,N_24267,N_24590);
nand UO_2948 (O_2948,N_24721,N_24801);
nor UO_2949 (O_2949,N_24393,N_23779);
nor UO_2950 (O_2950,N_24125,N_24032);
and UO_2951 (O_2951,N_24042,N_24457);
nor UO_2952 (O_2952,N_23759,N_24128);
xor UO_2953 (O_2953,N_23998,N_24636);
or UO_2954 (O_2954,N_23804,N_23860);
xnor UO_2955 (O_2955,N_24831,N_23961);
or UO_2956 (O_2956,N_23839,N_23868);
or UO_2957 (O_2957,N_24366,N_23978);
xnor UO_2958 (O_2958,N_24825,N_24630);
xor UO_2959 (O_2959,N_24667,N_24420);
xnor UO_2960 (O_2960,N_23980,N_24666);
nor UO_2961 (O_2961,N_24500,N_23926);
and UO_2962 (O_2962,N_24125,N_24813);
nand UO_2963 (O_2963,N_24819,N_24184);
nor UO_2964 (O_2964,N_24546,N_24130);
or UO_2965 (O_2965,N_24598,N_23922);
nor UO_2966 (O_2966,N_23983,N_24778);
nor UO_2967 (O_2967,N_23796,N_24731);
xor UO_2968 (O_2968,N_23796,N_24654);
nor UO_2969 (O_2969,N_23817,N_24740);
or UO_2970 (O_2970,N_24659,N_23879);
or UO_2971 (O_2971,N_24374,N_23813);
nor UO_2972 (O_2972,N_24278,N_23931);
nor UO_2973 (O_2973,N_24400,N_23931);
or UO_2974 (O_2974,N_24602,N_24148);
xor UO_2975 (O_2975,N_24583,N_24493);
and UO_2976 (O_2976,N_24528,N_24909);
or UO_2977 (O_2977,N_24813,N_23799);
and UO_2978 (O_2978,N_23781,N_23852);
nand UO_2979 (O_2979,N_24602,N_23851);
xnor UO_2980 (O_2980,N_24802,N_24376);
nor UO_2981 (O_2981,N_24926,N_24486);
xnor UO_2982 (O_2982,N_24236,N_24838);
or UO_2983 (O_2983,N_24402,N_24514);
xnor UO_2984 (O_2984,N_24044,N_23765);
xor UO_2985 (O_2985,N_23882,N_24140);
xor UO_2986 (O_2986,N_24496,N_24581);
nor UO_2987 (O_2987,N_24184,N_24885);
nand UO_2988 (O_2988,N_24780,N_24490);
nand UO_2989 (O_2989,N_24975,N_23782);
and UO_2990 (O_2990,N_24590,N_23841);
nand UO_2991 (O_2991,N_23855,N_24316);
and UO_2992 (O_2992,N_24720,N_24801);
nor UO_2993 (O_2993,N_23862,N_24411);
or UO_2994 (O_2994,N_24903,N_24808);
or UO_2995 (O_2995,N_23821,N_24223);
xnor UO_2996 (O_2996,N_23847,N_23810);
and UO_2997 (O_2997,N_24437,N_24918);
and UO_2998 (O_2998,N_24847,N_24806);
xnor UO_2999 (O_2999,N_24198,N_24448);
endmodule