module basic_500_3000_500_3_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_90,In_368);
nand U1 (N_1,In_347,In_47);
and U2 (N_2,In_92,In_498);
or U3 (N_3,In_73,In_12);
and U4 (N_4,In_230,In_176);
and U5 (N_5,In_252,In_345);
xnor U6 (N_6,In_100,In_476);
or U7 (N_7,In_406,In_223);
nor U8 (N_8,In_56,In_53);
xor U9 (N_9,In_114,In_281);
nor U10 (N_10,In_13,In_83);
nand U11 (N_11,In_191,In_208);
and U12 (N_12,In_175,In_210);
nand U13 (N_13,In_106,In_153);
and U14 (N_14,In_243,In_299);
nor U15 (N_15,In_264,In_438);
nor U16 (N_16,In_415,In_456);
or U17 (N_17,In_34,In_387);
or U18 (N_18,In_18,In_494);
nand U19 (N_19,In_475,In_414);
xor U20 (N_20,In_481,In_474);
nand U21 (N_21,In_420,In_152);
nor U22 (N_22,In_473,In_333);
xnor U23 (N_23,In_180,In_0);
and U24 (N_24,In_36,In_313);
nor U25 (N_25,In_284,In_91);
or U26 (N_26,In_156,In_198);
and U27 (N_27,In_188,In_460);
and U28 (N_28,In_427,In_261);
nand U29 (N_29,In_104,In_331);
and U30 (N_30,In_364,In_317);
xnor U31 (N_31,In_40,In_51);
and U32 (N_32,In_351,In_170);
xor U33 (N_33,In_404,In_55);
or U34 (N_34,In_386,In_107);
xnor U35 (N_35,In_214,In_298);
or U36 (N_36,In_183,In_88);
or U37 (N_37,In_256,In_209);
xnor U38 (N_38,In_353,In_161);
nor U39 (N_39,In_461,In_126);
and U40 (N_40,In_325,In_362);
xor U41 (N_41,In_479,In_242);
nor U42 (N_42,In_365,In_162);
and U43 (N_43,In_154,In_105);
nand U44 (N_44,In_16,In_169);
xor U45 (N_45,In_94,In_167);
and U46 (N_46,In_292,In_289);
or U47 (N_47,In_430,In_269);
or U48 (N_48,In_311,In_149);
and U49 (N_49,In_371,In_488);
xor U50 (N_50,In_22,In_428);
xnor U51 (N_51,In_57,In_446);
or U52 (N_52,In_140,In_141);
and U53 (N_53,In_369,In_463);
nand U54 (N_54,In_440,In_253);
and U55 (N_55,In_426,In_128);
and U56 (N_56,In_423,In_268);
nand U57 (N_57,In_86,In_118);
xor U58 (N_58,In_168,In_410);
nand U59 (N_59,In_95,In_472);
nor U60 (N_60,In_31,In_335);
or U61 (N_61,In_151,In_424);
xnor U62 (N_62,In_236,In_246);
or U63 (N_63,In_412,In_316);
nor U64 (N_64,In_379,In_108);
and U65 (N_65,In_30,In_159);
nand U66 (N_66,In_113,In_134);
nand U67 (N_67,In_482,In_224);
nand U68 (N_68,In_186,In_480);
nand U69 (N_69,In_244,In_164);
and U70 (N_70,In_355,In_288);
nand U71 (N_71,In_382,In_41);
nor U72 (N_72,In_499,In_258);
and U73 (N_73,In_150,In_119);
or U74 (N_74,In_181,In_241);
and U75 (N_75,In_346,In_21);
nand U76 (N_76,In_489,In_216);
nand U77 (N_77,In_24,In_367);
or U78 (N_78,In_323,In_303);
and U79 (N_79,In_177,In_235);
and U80 (N_80,In_458,In_229);
and U81 (N_81,In_96,In_321);
nand U82 (N_82,In_37,In_413);
nor U83 (N_83,In_130,In_206);
or U84 (N_84,In_68,In_77);
nand U85 (N_85,In_334,In_308);
and U86 (N_86,In_343,In_304);
nand U87 (N_87,In_464,In_495);
and U88 (N_88,In_459,In_467);
or U89 (N_89,In_129,In_99);
nor U90 (N_90,In_207,In_190);
nor U91 (N_91,In_219,In_221);
nor U92 (N_92,In_44,In_434);
and U93 (N_93,In_120,In_443);
or U94 (N_94,In_338,In_43);
nand U95 (N_95,In_396,In_60);
and U96 (N_96,In_436,In_136);
xor U97 (N_97,In_417,In_80);
and U98 (N_98,In_232,In_14);
and U99 (N_99,In_419,In_293);
and U100 (N_100,In_337,In_237);
nand U101 (N_101,In_283,In_455);
nand U102 (N_102,In_145,In_266);
nor U103 (N_103,In_416,In_380);
nand U104 (N_104,In_381,In_447);
nor U105 (N_105,In_182,In_227);
or U106 (N_106,In_75,In_296);
and U107 (N_107,In_211,In_32);
nand U108 (N_108,In_233,In_245);
and U109 (N_109,In_318,In_69);
or U110 (N_110,In_139,In_354);
nand U111 (N_111,In_437,In_59);
or U112 (N_112,In_231,In_9);
nor U113 (N_113,In_360,In_263);
nand U114 (N_114,In_247,In_204);
and U115 (N_115,In_148,In_271);
and U116 (N_116,In_179,In_195);
and U117 (N_117,In_6,In_225);
nand U118 (N_118,In_84,In_407);
and U119 (N_119,In_307,In_185);
nor U120 (N_120,In_262,In_490);
and U121 (N_121,In_276,In_110);
nand U122 (N_122,In_52,In_117);
nand U123 (N_123,In_8,In_385);
nand U124 (N_124,In_444,In_294);
nand U125 (N_125,In_121,In_295);
or U126 (N_126,In_312,In_297);
or U127 (N_127,In_131,In_239);
xor U128 (N_128,In_402,In_485);
or U129 (N_129,In_255,In_89);
and U130 (N_130,In_222,In_497);
or U131 (N_131,In_138,In_193);
or U132 (N_132,In_265,In_187);
nor U133 (N_133,In_7,In_341);
and U134 (N_134,In_42,In_274);
and U135 (N_135,In_314,In_425);
xnor U136 (N_136,In_1,In_226);
or U137 (N_137,In_445,In_278);
xor U138 (N_138,In_248,In_192);
and U139 (N_139,In_286,In_363);
and U140 (N_140,In_109,In_122);
nor U141 (N_141,In_282,In_123);
nand U142 (N_142,In_127,In_330);
nor U143 (N_143,In_372,In_442);
nor U144 (N_144,In_116,In_431);
nand U145 (N_145,In_93,In_78);
xnor U146 (N_146,In_384,In_54);
or U147 (N_147,In_433,In_63);
nand U148 (N_148,In_377,In_3);
and U149 (N_149,In_39,In_273);
nor U150 (N_150,In_102,In_391);
nor U151 (N_151,In_189,In_422);
nand U152 (N_152,In_328,In_234);
or U153 (N_153,In_409,In_394);
nor U154 (N_154,In_142,In_260);
xor U155 (N_155,In_215,In_212);
or U156 (N_156,In_393,In_220);
or U157 (N_157,In_270,In_49);
nand U158 (N_158,In_315,In_203);
or U159 (N_159,In_174,In_395);
nor U160 (N_160,In_309,In_448);
nor U161 (N_161,In_132,In_249);
and U162 (N_162,In_101,In_115);
and U163 (N_163,In_429,In_33);
nand U164 (N_164,In_327,In_85);
xor U165 (N_165,In_398,In_125);
and U166 (N_166,In_238,In_111);
xnor U167 (N_167,In_202,In_124);
xnor U168 (N_168,In_137,In_392);
nand U169 (N_169,In_79,In_435);
nor U170 (N_170,In_285,In_25);
nor U171 (N_171,In_82,In_477);
nand U172 (N_172,In_135,In_366);
and U173 (N_173,In_72,In_452);
xnor U174 (N_174,In_155,In_103);
nand U175 (N_175,In_98,In_38);
nand U176 (N_176,In_378,In_173);
and U177 (N_177,In_466,In_342);
xnor U178 (N_178,In_450,In_487);
and U179 (N_179,In_171,In_35);
and U180 (N_180,In_10,In_287);
xor U181 (N_181,In_205,In_468);
or U182 (N_182,In_201,In_301);
and U183 (N_183,In_496,In_71);
and U184 (N_184,In_352,In_336);
or U185 (N_185,In_199,In_484);
and U186 (N_186,In_228,In_441);
nand U187 (N_187,In_184,In_340);
and U188 (N_188,In_250,In_449);
xor U189 (N_189,In_370,In_324);
nor U190 (N_190,In_357,In_401);
nor U191 (N_191,In_26,In_350);
nor U192 (N_192,In_251,In_418);
or U193 (N_193,In_397,In_112);
and U194 (N_194,In_310,In_462);
nand U195 (N_195,In_15,In_359);
or U196 (N_196,In_302,In_196);
or U197 (N_197,In_451,In_218);
nand U198 (N_198,In_405,In_17);
or U199 (N_199,In_348,In_290);
xor U200 (N_200,In_11,In_332);
nand U201 (N_201,In_46,In_453);
nor U202 (N_202,In_27,In_160);
nor U203 (N_203,In_383,In_454);
nand U204 (N_204,In_469,In_326);
or U205 (N_205,In_439,In_471);
and U206 (N_206,In_319,In_158);
or U207 (N_207,In_388,In_144);
nand U208 (N_208,In_279,In_66);
nor U209 (N_209,In_305,In_48);
or U210 (N_210,In_5,In_165);
and U211 (N_211,In_376,In_257);
or U212 (N_212,In_259,In_28);
nand U213 (N_213,In_374,In_19);
and U214 (N_214,In_349,In_87);
nor U215 (N_215,In_163,In_329);
and U216 (N_216,In_178,In_361);
or U217 (N_217,In_465,In_493);
nor U218 (N_218,In_356,In_2);
nand U219 (N_219,In_23,In_166);
or U220 (N_220,In_217,In_344);
or U221 (N_221,In_20,In_146);
xnor U222 (N_222,In_50,In_200);
or U223 (N_223,In_4,In_277);
nor U224 (N_224,In_29,In_390);
nand U225 (N_225,In_81,In_291);
or U226 (N_226,In_70,In_280);
nor U227 (N_227,In_45,In_400);
xor U228 (N_228,In_143,In_97);
or U229 (N_229,In_61,In_254);
and U230 (N_230,In_457,In_421);
nand U231 (N_231,In_375,In_403);
and U232 (N_232,In_62,In_76);
nand U233 (N_233,In_74,In_483);
nor U234 (N_234,In_432,In_373);
and U235 (N_235,In_147,In_470);
or U236 (N_236,In_399,In_320);
nand U237 (N_237,In_65,In_492);
or U238 (N_238,In_300,In_358);
or U239 (N_239,In_486,In_64);
or U240 (N_240,In_411,In_58);
and U241 (N_241,In_389,In_408);
xor U242 (N_242,In_157,In_197);
or U243 (N_243,In_267,In_213);
nand U244 (N_244,In_322,In_194);
nand U245 (N_245,In_478,In_172);
nor U246 (N_246,In_240,In_272);
nor U247 (N_247,In_275,In_133);
or U248 (N_248,In_339,In_306);
nand U249 (N_249,In_491,In_67);
nor U250 (N_250,In_13,In_414);
or U251 (N_251,In_122,In_459);
xnor U252 (N_252,In_257,In_1);
nor U253 (N_253,In_51,In_461);
nand U254 (N_254,In_440,In_404);
nor U255 (N_255,In_68,In_228);
nand U256 (N_256,In_68,In_339);
or U257 (N_257,In_203,In_18);
and U258 (N_258,In_292,In_74);
or U259 (N_259,In_472,In_434);
nand U260 (N_260,In_247,In_398);
and U261 (N_261,In_499,In_371);
nor U262 (N_262,In_296,In_369);
nor U263 (N_263,In_381,In_428);
and U264 (N_264,In_93,In_279);
xnor U265 (N_265,In_123,In_188);
nand U266 (N_266,In_260,In_252);
or U267 (N_267,In_23,In_12);
and U268 (N_268,In_134,In_163);
nand U269 (N_269,In_72,In_249);
and U270 (N_270,In_128,In_451);
nor U271 (N_271,In_399,In_278);
and U272 (N_272,In_215,In_267);
nand U273 (N_273,In_55,In_338);
and U274 (N_274,In_112,In_455);
or U275 (N_275,In_482,In_463);
nand U276 (N_276,In_465,In_56);
and U277 (N_277,In_492,In_348);
and U278 (N_278,In_81,In_406);
or U279 (N_279,In_78,In_225);
or U280 (N_280,In_145,In_488);
and U281 (N_281,In_213,In_106);
or U282 (N_282,In_262,In_264);
and U283 (N_283,In_340,In_317);
or U284 (N_284,In_411,In_231);
nand U285 (N_285,In_41,In_490);
nor U286 (N_286,In_461,In_107);
nand U287 (N_287,In_226,In_421);
and U288 (N_288,In_242,In_328);
nor U289 (N_289,In_380,In_113);
nor U290 (N_290,In_320,In_448);
nand U291 (N_291,In_211,In_431);
nand U292 (N_292,In_82,In_374);
or U293 (N_293,In_455,In_244);
xnor U294 (N_294,In_155,In_270);
and U295 (N_295,In_232,In_70);
and U296 (N_296,In_18,In_294);
and U297 (N_297,In_101,In_178);
and U298 (N_298,In_271,In_390);
or U299 (N_299,In_234,In_495);
xnor U300 (N_300,In_19,In_391);
nor U301 (N_301,In_431,In_185);
or U302 (N_302,In_449,In_196);
xnor U303 (N_303,In_246,In_168);
nor U304 (N_304,In_14,In_308);
nand U305 (N_305,In_236,In_336);
or U306 (N_306,In_48,In_304);
or U307 (N_307,In_326,In_262);
xnor U308 (N_308,In_273,In_429);
nand U309 (N_309,In_66,In_108);
nand U310 (N_310,In_73,In_396);
nor U311 (N_311,In_194,In_318);
nor U312 (N_312,In_170,In_418);
nor U313 (N_313,In_195,In_41);
xnor U314 (N_314,In_178,In_482);
and U315 (N_315,In_180,In_420);
or U316 (N_316,In_292,In_244);
nor U317 (N_317,In_290,In_341);
and U318 (N_318,In_16,In_218);
and U319 (N_319,In_258,In_273);
xor U320 (N_320,In_81,In_38);
and U321 (N_321,In_381,In_294);
nand U322 (N_322,In_218,In_422);
nor U323 (N_323,In_380,In_409);
and U324 (N_324,In_356,In_206);
nand U325 (N_325,In_162,In_255);
nand U326 (N_326,In_304,In_453);
and U327 (N_327,In_409,In_82);
nor U328 (N_328,In_87,In_462);
or U329 (N_329,In_341,In_393);
or U330 (N_330,In_7,In_100);
nand U331 (N_331,In_425,In_354);
or U332 (N_332,In_348,In_150);
or U333 (N_333,In_167,In_118);
and U334 (N_334,In_152,In_305);
nand U335 (N_335,In_303,In_64);
nand U336 (N_336,In_459,In_177);
nor U337 (N_337,In_472,In_378);
nor U338 (N_338,In_231,In_35);
nand U339 (N_339,In_377,In_38);
or U340 (N_340,In_251,In_465);
or U341 (N_341,In_296,In_371);
nor U342 (N_342,In_394,In_246);
nor U343 (N_343,In_257,In_218);
nor U344 (N_344,In_362,In_478);
nand U345 (N_345,In_143,In_330);
nand U346 (N_346,In_63,In_323);
nand U347 (N_347,In_199,In_407);
nor U348 (N_348,In_351,In_442);
nand U349 (N_349,In_353,In_135);
nand U350 (N_350,In_423,In_474);
nand U351 (N_351,In_61,In_428);
and U352 (N_352,In_181,In_422);
and U353 (N_353,In_21,In_343);
xnor U354 (N_354,In_14,In_475);
nor U355 (N_355,In_352,In_431);
nand U356 (N_356,In_370,In_304);
nand U357 (N_357,In_464,In_316);
or U358 (N_358,In_106,In_121);
nor U359 (N_359,In_128,In_342);
and U360 (N_360,In_474,In_459);
nand U361 (N_361,In_389,In_472);
nor U362 (N_362,In_368,In_238);
xor U363 (N_363,In_187,In_221);
or U364 (N_364,In_253,In_22);
and U365 (N_365,In_327,In_411);
nand U366 (N_366,In_197,In_283);
and U367 (N_367,In_111,In_320);
nor U368 (N_368,In_206,In_192);
nor U369 (N_369,In_223,In_237);
nand U370 (N_370,In_466,In_301);
nor U371 (N_371,In_195,In_408);
nor U372 (N_372,In_46,In_255);
nor U373 (N_373,In_284,In_344);
xor U374 (N_374,In_462,In_480);
or U375 (N_375,In_396,In_66);
nand U376 (N_376,In_294,In_449);
nor U377 (N_377,In_316,In_296);
nand U378 (N_378,In_29,In_77);
nor U379 (N_379,In_348,In_147);
or U380 (N_380,In_18,In_14);
nor U381 (N_381,In_118,In_307);
and U382 (N_382,In_392,In_290);
nand U383 (N_383,In_29,In_158);
nor U384 (N_384,In_291,In_83);
and U385 (N_385,In_332,In_25);
and U386 (N_386,In_267,In_175);
xor U387 (N_387,In_345,In_261);
or U388 (N_388,In_204,In_276);
nor U389 (N_389,In_447,In_369);
or U390 (N_390,In_40,In_61);
xnor U391 (N_391,In_58,In_414);
nor U392 (N_392,In_337,In_183);
nor U393 (N_393,In_459,In_478);
and U394 (N_394,In_38,In_375);
and U395 (N_395,In_463,In_480);
or U396 (N_396,In_72,In_354);
or U397 (N_397,In_376,In_321);
and U398 (N_398,In_390,In_241);
or U399 (N_399,In_423,In_17);
and U400 (N_400,In_306,In_234);
or U401 (N_401,In_115,In_482);
nor U402 (N_402,In_92,In_81);
nand U403 (N_403,In_47,In_61);
and U404 (N_404,In_438,In_443);
and U405 (N_405,In_410,In_38);
nor U406 (N_406,In_263,In_219);
nor U407 (N_407,In_124,In_491);
nand U408 (N_408,In_331,In_62);
and U409 (N_409,In_303,In_482);
or U410 (N_410,In_385,In_179);
and U411 (N_411,In_430,In_96);
and U412 (N_412,In_295,In_246);
or U413 (N_413,In_378,In_423);
xnor U414 (N_414,In_16,In_455);
and U415 (N_415,In_129,In_202);
xor U416 (N_416,In_168,In_19);
xor U417 (N_417,In_445,In_81);
xnor U418 (N_418,In_213,In_44);
nor U419 (N_419,In_498,In_347);
nand U420 (N_420,In_452,In_138);
and U421 (N_421,In_38,In_110);
xnor U422 (N_422,In_15,In_160);
and U423 (N_423,In_333,In_381);
and U424 (N_424,In_263,In_260);
xor U425 (N_425,In_33,In_213);
nand U426 (N_426,In_269,In_300);
or U427 (N_427,In_7,In_379);
or U428 (N_428,In_404,In_411);
and U429 (N_429,In_9,In_276);
xnor U430 (N_430,In_431,In_180);
and U431 (N_431,In_289,In_71);
nand U432 (N_432,In_290,In_243);
and U433 (N_433,In_37,In_275);
nor U434 (N_434,In_383,In_243);
and U435 (N_435,In_308,In_361);
nor U436 (N_436,In_201,In_328);
and U437 (N_437,In_491,In_207);
nor U438 (N_438,In_192,In_356);
nand U439 (N_439,In_378,In_488);
or U440 (N_440,In_348,In_347);
or U441 (N_441,In_309,In_362);
and U442 (N_442,In_155,In_313);
and U443 (N_443,In_180,In_353);
or U444 (N_444,In_83,In_362);
nand U445 (N_445,In_402,In_238);
and U446 (N_446,In_466,In_133);
nor U447 (N_447,In_475,In_67);
or U448 (N_448,In_393,In_106);
and U449 (N_449,In_85,In_484);
nand U450 (N_450,In_66,In_6);
or U451 (N_451,In_308,In_88);
or U452 (N_452,In_366,In_107);
xor U453 (N_453,In_163,In_351);
nand U454 (N_454,In_134,In_47);
and U455 (N_455,In_16,In_479);
or U456 (N_456,In_371,In_437);
nand U457 (N_457,In_494,In_320);
nand U458 (N_458,In_226,In_133);
nor U459 (N_459,In_406,In_246);
nor U460 (N_460,In_405,In_250);
nand U461 (N_461,In_453,In_272);
nor U462 (N_462,In_442,In_132);
nor U463 (N_463,In_220,In_216);
nor U464 (N_464,In_176,In_90);
xnor U465 (N_465,In_274,In_73);
nand U466 (N_466,In_11,In_206);
or U467 (N_467,In_368,In_57);
and U468 (N_468,In_358,In_123);
nand U469 (N_469,In_73,In_394);
nand U470 (N_470,In_306,In_262);
or U471 (N_471,In_282,In_107);
xor U472 (N_472,In_5,In_232);
and U473 (N_473,In_111,In_28);
nor U474 (N_474,In_490,In_325);
nand U475 (N_475,In_90,In_125);
nor U476 (N_476,In_286,In_285);
or U477 (N_477,In_359,In_43);
xor U478 (N_478,In_156,In_277);
nor U479 (N_479,In_216,In_129);
nor U480 (N_480,In_173,In_326);
or U481 (N_481,In_216,In_53);
nand U482 (N_482,In_268,In_477);
nor U483 (N_483,In_97,In_336);
and U484 (N_484,In_281,In_8);
nand U485 (N_485,In_336,In_403);
and U486 (N_486,In_345,In_323);
and U487 (N_487,In_130,In_186);
nor U488 (N_488,In_5,In_290);
or U489 (N_489,In_1,In_272);
nand U490 (N_490,In_41,In_310);
nor U491 (N_491,In_94,In_183);
and U492 (N_492,In_496,In_0);
nor U493 (N_493,In_169,In_422);
nor U494 (N_494,In_479,In_212);
nand U495 (N_495,In_166,In_271);
nand U496 (N_496,In_246,In_60);
or U497 (N_497,In_499,In_458);
or U498 (N_498,In_447,In_65);
or U499 (N_499,In_221,In_286);
nor U500 (N_500,In_220,In_242);
and U501 (N_501,In_456,In_49);
or U502 (N_502,In_367,In_9);
or U503 (N_503,In_347,In_483);
or U504 (N_504,In_435,In_245);
and U505 (N_505,In_38,In_58);
nand U506 (N_506,In_462,In_412);
and U507 (N_507,In_31,In_441);
nand U508 (N_508,In_280,In_277);
nand U509 (N_509,In_304,In_435);
nor U510 (N_510,In_295,In_467);
and U511 (N_511,In_270,In_165);
and U512 (N_512,In_246,In_114);
and U513 (N_513,In_66,In_281);
xor U514 (N_514,In_234,In_412);
nand U515 (N_515,In_322,In_127);
nand U516 (N_516,In_453,In_56);
or U517 (N_517,In_29,In_225);
nor U518 (N_518,In_110,In_61);
nor U519 (N_519,In_285,In_117);
and U520 (N_520,In_369,In_166);
nand U521 (N_521,In_133,In_475);
xnor U522 (N_522,In_448,In_55);
or U523 (N_523,In_65,In_185);
and U524 (N_524,In_441,In_332);
and U525 (N_525,In_459,In_361);
or U526 (N_526,In_361,In_322);
nand U527 (N_527,In_424,In_259);
nand U528 (N_528,In_387,In_325);
and U529 (N_529,In_14,In_151);
nand U530 (N_530,In_159,In_243);
and U531 (N_531,In_412,In_145);
and U532 (N_532,In_2,In_462);
and U533 (N_533,In_391,In_226);
nor U534 (N_534,In_195,In_175);
nand U535 (N_535,In_101,In_150);
or U536 (N_536,In_134,In_240);
and U537 (N_537,In_212,In_288);
and U538 (N_538,In_370,In_317);
nand U539 (N_539,In_397,In_275);
nand U540 (N_540,In_357,In_66);
and U541 (N_541,In_367,In_385);
nand U542 (N_542,In_361,In_384);
or U543 (N_543,In_82,In_482);
and U544 (N_544,In_388,In_206);
nand U545 (N_545,In_496,In_189);
nand U546 (N_546,In_14,In_155);
nand U547 (N_547,In_210,In_226);
or U548 (N_548,In_302,In_318);
nand U549 (N_549,In_217,In_484);
nand U550 (N_550,In_115,In_243);
xor U551 (N_551,In_237,In_56);
nand U552 (N_552,In_400,In_103);
nor U553 (N_553,In_424,In_291);
and U554 (N_554,In_407,In_360);
and U555 (N_555,In_150,In_461);
or U556 (N_556,In_161,In_275);
and U557 (N_557,In_429,In_313);
xor U558 (N_558,In_49,In_296);
nor U559 (N_559,In_69,In_342);
or U560 (N_560,In_155,In_68);
xor U561 (N_561,In_145,In_76);
or U562 (N_562,In_357,In_153);
or U563 (N_563,In_407,In_480);
and U564 (N_564,In_80,In_262);
nand U565 (N_565,In_76,In_443);
nor U566 (N_566,In_163,In_347);
nor U567 (N_567,In_194,In_56);
nor U568 (N_568,In_80,In_116);
nand U569 (N_569,In_94,In_232);
xnor U570 (N_570,In_494,In_64);
nand U571 (N_571,In_110,In_157);
and U572 (N_572,In_19,In_393);
nor U573 (N_573,In_337,In_248);
or U574 (N_574,In_324,In_289);
and U575 (N_575,In_486,In_456);
or U576 (N_576,In_113,In_254);
nand U577 (N_577,In_165,In_350);
nand U578 (N_578,In_53,In_249);
and U579 (N_579,In_164,In_104);
nor U580 (N_580,In_340,In_57);
xnor U581 (N_581,In_87,In_212);
and U582 (N_582,In_237,In_150);
nor U583 (N_583,In_28,In_70);
nand U584 (N_584,In_149,In_448);
nor U585 (N_585,In_390,In_57);
or U586 (N_586,In_24,In_34);
nor U587 (N_587,In_8,In_13);
xnor U588 (N_588,In_236,In_331);
and U589 (N_589,In_322,In_122);
and U590 (N_590,In_348,In_66);
xor U591 (N_591,In_307,In_268);
nand U592 (N_592,In_150,In_323);
or U593 (N_593,In_305,In_148);
or U594 (N_594,In_228,In_298);
nand U595 (N_595,In_109,In_44);
and U596 (N_596,In_356,In_130);
or U597 (N_597,In_448,In_78);
nor U598 (N_598,In_155,In_478);
nand U599 (N_599,In_281,In_33);
xor U600 (N_600,In_80,In_402);
nand U601 (N_601,In_391,In_198);
nor U602 (N_602,In_8,In_40);
nor U603 (N_603,In_167,In_392);
nor U604 (N_604,In_313,In_102);
or U605 (N_605,In_254,In_152);
or U606 (N_606,In_145,In_21);
nand U607 (N_607,In_312,In_98);
xor U608 (N_608,In_409,In_30);
and U609 (N_609,In_498,In_276);
and U610 (N_610,In_474,In_394);
nor U611 (N_611,In_91,In_136);
and U612 (N_612,In_0,In_440);
and U613 (N_613,In_401,In_264);
nand U614 (N_614,In_74,In_407);
nor U615 (N_615,In_200,In_266);
nor U616 (N_616,In_181,In_304);
or U617 (N_617,In_68,In_121);
and U618 (N_618,In_380,In_381);
or U619 (N_619,In_23,In_291);
xor U620 (N_620,In_73,In_346);
or U621 (N_621,In_473,In_223);
or U622 (N_622,In_287,In_121);
nor U623 (N_623,In_230,In_155);
nand U624 (N_624,In_35,In_261);
nand U625 (N_625,In_478,In_170);
and U626 (N_626,In_307,In_208);
nand U627 (N_627,In_22,In_195);
and U628 (N_628,In_149,In_64);
and U629 (N_629,In_66,In_89);
nor U630 (N_630,In_121,In_416);
or U631 (N_631,In_372,In_125);
and U632 (N_632,In_482,In_250);
nor U633 (N_633,In_393,In_97);
nor U634 (N_634,In_102,In_342);
nand U635 (N_635,In_354,In_66);
or U636 (N_636,In_363,In_93);
nand U637 (N_637,In_416,In_264);
and U638 (N_638,In_38,In_361);
and U639 (N_639,In_4,In_243);
or U640 (N_640,In_310,In_186);
nor U641 (N_641,In_494,In_78);
nand U642 (N_642,In_137,In_450);
or U643 (N_643,In_487,In_103);
nor U644 (N_644,In_457,In_331);
nand U645 (N_645,In_365,In_386);
and U646 (N_646,In_342,In_84);
or U647 (N_647,In_202,In_100);
xor U648 (N_648,In_18,In_427);
nand U649 (N_649,In_131,In_318);
or U650 (N_650,In_361,In_219);
and U651 (N_651,In_114,In_276);
or U652 (N_652,In_418,In_412);
nor U653 (N_653,In_176,In_259);
nor U654 (N_654,In_427,In_251);
and U655 (N_655,In_466,In_472);
xor U656 (N_656,In_406,In_402);
and U657 (N_657,In_208,In_59);
xnor U658 (N_658,In_85,In_101);
and U659 (N_659,In_313,In_58);
nor U660 (N_660,In_161,In_446);
or U661 (N_661,In_285,In_48);
nor U662 (N_662,In_167,In_71);
or U663 (N_663,In_300,In_261);
nor U664 (N_664,In_50,In_116);
nand U665 (N_665,In_292,In_99);
nor U666 (N_666,In_379,In_287);
or U667 (N_667,In_499,In_497);
nor U668 (N_668,In_398,In_8);
nor U669 (N_669,In_151,In_310);
nand U670 (N_670,In_33,In_377);
or U671 (N_671,In_68,In_207);
nor U672 (N_672,In_251,In_328);
nand U673 (N_673,In_56,In_164);
nand U674 (N_674,In_323,In_348);
and U675 (N_675,In_293,In_308);
and U676 (N_676,In_147,In_354);
nor U677 (N_677,In_459,In_60);
or U678 (N_678,In_244,In_279);
and U679 (N_679,In_141,In_241);
nand U680 (N_680,In_18,In_345);
and U681 (N_681,In_479,In_373);
nor U682 (N_682,In_413,In_90);
nor U683 (N_683,In_321,In_469);
or U684 (N_684,In_33,In_243);
nand U685 (N_685,In_49,In_279);
nand U686 (N_686,In_109,In_76);
or U687 (N_687,In_125,In_97);
xnor U688 (N_688,In_71,In_73);
nand U689 (N_689,In_197,In_484);
nor U690 (N_690,In_207,In_25);
or U691 (N_691,In_498,In_75);
nor U692 (N_692,In_43,In_445);
or U693 (N_693,In_59,In_246);
and U694 (N_694,In_365,In_208);
xor U695 (N_695,In_497,In_424);
nand U696 (N_696,In_107,In_449);
and U697 (N_697,In_220,In_404);
xor U698 (N_698,In_70,In_416);
nor U699 (N_699,In_401,In_74);
or U700 (N_700,In_453,In_177);
and U701 (N_701,In_350,In_340);
or U702 (N_702,In_190,In_169);
or U703 (N_703,In_330,In_393);
nor U704 (N_704,In_168,In_298);
and U705 (N_705,In_368,In_433);
and U706 (N_706,In_195,In_201);
xor U707 (N_707,In_245,In_337);
or U708 (N_708,In_119,In_418);
nor U709 (N_709,In_200,In_291);
and U710 (N_710,In_270,In_75);
and U711 (N_711,In_355,In_114);
nor U712 (N_712,In_119,In_265);
nand U713 (N_713,In_81,In_33);
and U714 (N_714,In_481,In_209);
and U715 (N_715,In_336,In_10);
nor U716 (N_716,In_417,In_453);
nand U717 (N_717,In_274,In_235);
and U718 (N_718,In_298,In_83);
or U719 (N_719,In_64,In_459);
nor U720 (N_720,In_286,In_99);
nor U721 (N_721,In_13,In_166);
nand U722 (N_722,In_180,In_484);
nand U723 (N_723,In_220,In_283);
nand U724 (N_724,In_490,In_232);
nand U725 (N_725,In_132,In_488);
and U726 (N_726,In_290,In_120);
nor U727 (N_727,In_294,In_300);
xnor U728 (N_728,In_162,In_130);
or U729 (N_729,In_429,In_106);
nand U730 (N_730,In_222,In_215);
nor U731 (N_731,In_106,In_206);
or U732 (N_732,In_55,In_130);
nor U733 (N_733,In_369,In_198);
and U734 (N_734,In_449,In_136);
and U735 (N_735,In_227,In_170);
xnor U736 (N_736,In_340,In_269);
or U737 (N_737,In_157,In_76);
and U738 (N_738,In_92,In_0);
xnor U739 (N_739,In_456,In_423);
and U740 (N_740,In_232,In_323);
nand U741 (N_741,In_79,In_485);
and U742 (N_742,In_27,In_58);
xnor U743 (N_743,In_105,In_70);
nand U744 (N_744,In_219,In_30);
nand U745 (N_745,In_104,In_114);
and U746 (N_746,In_234,In_93);
nand U747 (N_747,In_252,In_284);
nor U748 (N_748,In_255,In_450);
and U749 (N_749,In_267,In_194);
or U750 (N_750,In_398,In_475);
and U751 (N_751,In_2,In_475);
or U752 (N_752,In_39,In_367);
xor U753 (N_753,In_267,In_252);
and U754 (N_754,In_229,In_275);
and U755 (N_755,In_313,In_124);
or U756 (N_756,In_251,In_93);
nand U757 (N_757,In_211,In_374);
or U758 (N_758,In_447,In_89);
xnor U759 (N_759,In_51,In_73);
or U760 (N_760,In_23,In_430);
nor U761 (N_761,In_39,In_461);
and U762 (N_762,In_186,In_335);
nand U763 (N_763,In_322,In_493);
nor U764 (N_764,In_273,In_476);
nor U765 (N_765,In_142,In_404);
nor U766 (N_766,In_104,In_410);
nand U767 (N_767,In_297,In_229);
nand U768 (N_768,In_475,In_4);
and U769 (N_769,In_345,In_183);
or U770 (N_770,In_3,In_257);
and U771 (N_771,In_136,In_166);
nor U772 (N_772,In_26,In_164);
and U773 (N_773,In_350,In_150);
nand U774 (N_774,In_418,In_11);
or U775 (N_775,In_322,In_98);
nand U776 (N_776,In_119,In_342);
nor U777 (N_777,In_239,In_397);
nor U778 (N_778,In_370,In_488);
xor U779 (N_779,In_311,In_65);
nand U780 (N_780,In_272,In_294);
or U781 (N_781,In_18,In_413);
nor U782 (N_782,In_117,In_112);
nor U783 (N_783,In_217,In_434);
nand U784 (N_784,In_127,In_378);
and U785 (N_785,In_8,In_14);
nand U786 (N_786,In_473,In_444);
xor U787 (N_787,In_397,In_249);
nand U788 (N_788,In_264,In_76);
xor U789 (N_789,In_369,In_137);
and U790 (N_790,In_149,In_420);
nand U791 (N_791,In_442,In_29);
xor U792 (N_792,In_146,In_213);
or U793 (N_793,In_474,In_112);
or U794 (N_794,In_193,In_488);
nor U795 (N_795,In_486,In_77);
and U796 (N_796,In_138,In_328);
nand U797 (N_797,In_434,In_216);
or U798 (N_798,In_350,In_175);
or U799 (N_799,In_460,In_399);
nand U800 (N_800,In_344,In_32);
xnor U801 (N_801,In_395,In_330);
nor U802 (N_802,In_242,In_182);
and U803 (N_803,In_436,In_204);
and U804 (N_804,In_195,In_185);
xnor U805 (N_805,In_116,In_2);
and U806 (N_806,In_20,In_195);
xor U807 (N_807,In_322,In_228);
or U808 (N_808,In_469,In_250);
xor U809 (N_809,In_60,In_323);
nand U810 (N_810,In_25,In_90);
nor U811 (N_811,In_358,In_7);
or U812 (N_812,In_73,In_267);
nor U813 (N_813,In_372,In_2);
and U814 (N_814,In_35,In_223);
nor U815 (N_815,In_425,In_385);
nand U816 (N_816,In_254,In_242);
nand U817 (N_817,In_48,In_396);
or U818 (N_818,In_324,In_435);
nand U819 (N_819,In_9,In_33);
nand U820 (N_820,In_1,In_167);
and U821 (N_821,In_179,In_193);
or U822 (N_822,In_178,In_131);
and U823 (N_823,In_351,In_133);
or U824 (N_824,In_475,In_313);
and U825 (N_825,In_237,In_256);
and U826 (N_826,In_365,In_223);
nand U827 (N_827,In_447,In_494);
and U828 (N_828,In_355,In_431);
nand U829 (N_829,In_90,In_108);
nand U830 (N_830,In_371,In_355);
or U831 (N_831,In_53,In_309);
and U832 (N_832,In_134,In_417);
and U833 (N_833,In_370,In_144);
nor U834 (N_834,In_90,In_164);
or U835 (N_835,In_104,In_436);
and U836 (N_836,In_358,In_488);
or U837 (N_837,In_332,In_357);
and U838 (N_838,In_159,In_148);
or U839 (N_839,In_384,In_284);
nand U840 (N_840,In_355,In_405);
nand U841 (N_841,In_220,In_232);
nor U842 (N_842,In_141,In_384);
and U843 (N_843,In_42,In_480);
and U844 (N_844,In_285,In_180);
nor U845 (N_845,In_198,In_197);
or U846 (N_846,In_324,In_113);
xor U847 (N_847,In_241,In_92);
or U848 (N_848,In_202,In_410);
xor U849 (N_849,In_234,In_5);
and U850 (N_850,In_312,In_480);
nand U851 (N_851,In_217,In_384);
xor U852 (N_852,In_406,In_257);
nand U853 (N_853,In_72,In_207);
nor U854 (N_854,In_12,In_463);
and U855 (N_855,In_266,In_331);
nor U856 (N_856,In_101,In_36);
nand U857 (N_857,In_417,In_280);
or U858 (N_858,In_166,In_52);
and U859 (N_859,In_474,In_428);
or U860 (N_860,In_427,In_474);
nand U861 (N_861,In_193,In_89);
and U862 (N_862,In_332,In_429);
or U863 (N_863,In_450,In_69);
or U864 (N_864,In_185,In_41);
nor U865 (N_865,In_224,In_345);
and U866 (N_866,In_257,In_263);
nand U867 (N_867,In_147,In_293);
or U868 (N_868,In_5,In_315);
nor U869 (N_869,In_27,In_103);
and U870 (N_870,In_427,In_307);
nand U871 (N_871,In_67,In_216);
nor U872 (N_872,In_387,In_152);
nor U873 (N_873,In_44,In_336);
xor U874 (N_874,In_339,In_277);
and U875 (N_875,In_46,In_312);
and U876 (N_876,In_242,In_71);
or U877 (N_877,In_231,In_73);
or U878 (N_878,In_0,In_327);
and U879 (N_879,In_110,In_220);
nand U880 (N_880,In_2,In_292);
or U881 (N_881,In_201,In_81);
or U882 (N_882,In_374,In_404);
and U883 (N_883,In_157,In_254);
and U884 (N_884,In_82,In_44);
and U885 (N_885,In_194,In_166);
nor U886 (N_886,In_118,In_13);
nand U887 (N_887,In_251,In_130);
nand U888 (N_888,In_42,In_207);
nor U889 (N_889,In_390,In_379);
nand U890 (N_890,In_100,In_200);
nand U891 (N_891,In_73,In_342);
and U892 (N_892,In_129,In_107);
or U893 (N_893,In_162,In_405);
nand U894 (N_894,In_97,In_433);
and U895 (N_895,In_455,In_226);
or U896 (N_896,In_160,In_46);
nor U897 (N_897,In_236,In_164);
nor U898 (N_898,In_48,In_115);
xnor U899 (N_899,In_202,In_101);
and U900 (N_900,In_126,In_18);
nor U901 (N_901,In_124,In_427);
and U902 (N_902,In_232,In_112);
or U903 (N_903,In_49,In_483);
and U904 (N_904,In_283,In_83);
nand U905 (N_905,In_162,In_106);
nand U906 (N_906,In_365,In_280);
nor U907 (N_907,In_174,In_223);
nor U908 (N_908,In_475,In_28);
or U909 (N_909,In_8,In_389);
and U910 (N_910,In_231,In_268);
or U911 (N_911,In_4,In_175);
and U912 (N_912,In_319,In_40);
and U913 (N_913,In_137,In_2);
or U914 (N_914,In_127,In_122);
and U915 (N_915,In_35,In_457);
and U916 (N_916,In_316,In_216);
nor U917 (N_917,In_18,In_125);
xnor U918 (N_918,In_448,In_201);
or U919 (N_919,In_85,In_284);
and U920 (N_920,In_345,In_122);
xor U921 (N_921,In_295,In_493);
and U922 (N_922,In_399,In_131);
and U923 (N_923,In_459,In_443);
xor U924 (N_924,In_17,In_222);
or U925 (N_925,In_248,In_485);
or U926 (N_926,In_242,In_388);
or U927 (N_927,In_414,In_156);
nor U928 (N_928,In_28,In_152);
nand U929 (N_929,In_314,In_282);
or U930 (N_930,In_154,In_334);
nand U931 (N_931,In_204,In_354);
nor U932 (N_932,In_444,In_269);
or U933 (N_933,In_440,In_96);
nor U934 (N_934,In_334,In_332);
nand U935 (N_935,In_91,In_487);
xnor U936 (N_936,In_461,In_413);
and U937 (N_937,In_275,In_268);
and U938 (N_938,In_62,In_431);
and U939 (N_939,In_269,In_342);
or U940 (N_940,In_163,In_266);
xor U941 (N_941,In_327,In_368);
nand U942 (N_942,In_175,In_459);
and U943 (N_943,In_96,In_105);
nor U944 (N_944,In_226,In_67);
or U945 (N_945,In_198,In_492);
or U946 (N_946,In_41,In_284);
nor U947 (N_947,In_422,In_115);
or U948 (N_948,In_349,In_227);
nand U949 (N_949,In_32,In_154);
xor U950 (N_950,In_67,In_492);
and U951 (N_951,In_299,In_98);
xor U952 (N_952,In_461,In_492);
or U953 (N_953,In_145,In_197);
nand U954 (N_954,In_274,In_215);
nor U955 (N_955,In_133,In_488);
and U956 (N_956,In_194,In_355);
nand U957 (N_957,In_56,In_496);
and U958 (N_958,In_215,In_487);
and U959 (N_959,In_108,In_278);
or U960 (N_960,In_355,In_417);
nand U961 (N_961,In_376,In_101);
nor U962 (N_962,In_201,In_406);
nand U963 (N_963,In_216,In_458);
nand U964 (N_964,In_365,In_427);
and U965 (N_965,In_26,In_299);
and U966 (N_966,In_90,In_280);
and U967 (N_967,In_178,In_129);
or U968 (N_968,In_488,In_208);
nand U969 (N_969,In_8,In_117);
nand U970 (N_970,In_211,In_167);
and U971 (N_971,In_392,In_176);
xnor U972 (N_972,In_128,In_159);
nor U973 (N_973,In_348,In_70);
xnor U974 (N_974,In_226,In_151);
nor U975 (N_975,In_191,In_218);
nor U976 (N_976,In_285,In_489);
or U977 (N_977,In_373,In_330);
nor U978 (N_978,In_88,In_496);
or U979 (N_979,In_213,In_331);
nand U980 (N_980,In_4,In_405);
xnor U981 (N_981,In_241,In_101);
xnor U982 (N_982,In_246,In_294);
nor U983 (N_983,In_410,In_83);
and U984 (N_984,In_198,In_389);
nand U985 (N_985,In_407,In_164);
and U986 (N_986,In_414,In_216);
nand U987 (N_987,In_195,In_168);
and U988 (N_988,In_80,In_77);
nor U989 (N_989,In_293,In_431);
nand U990 (N_990,In_56,In_337);
nor U991 (N_991,In_114,In_28);
nand U992 (N_992,In_497,In_344);
nor U993 (N_993,In_257,In_188);
and U994 (N_994,In_320,In_173);
nor U995 (N_995,In_390,In_79);
nand U996 (N_996,In_360,In_247);
xor U997 (N_997,In_154,In_219);
nor U998 (N_998,In_438,In_244);
and U999 (N_999,In_190,In_144);
nor U1000 (N_1000,N_204,N_96);
or U1001 (N_1001,N_636,N_86);
nand U1002 (N_1002,N_252,N_883);
nor U1003 (N_1003,N_786,N_348);
or U1004 (N_1004,N_500,N_908);
or U1005 (N_1005,N_360,N_964);
or U1006 (N_1006,N_587,N_205);
or U1007 (N_1007,N_757,N_231);
nand U1008 (N_1008,N_826,N_877);
or U1009 (N_1009,N_197,N_857);
or U1010 (N_1010,N_916,N_933);
nor U1011 (N_1011,N_974,N_407);
and U1012 (N_1012,N_732,N_842);
or U1013 (N_1013,N_542,N_195);
and U1014 (N_1014,N_919,N_42);
nand U1015 (N_1015,N_101,N_927);
and U1016 (N_1016,N_169,N_488);
nor U1017 (N_1017,N_520,N_991);
or U1018 (N_1018,N_453,N_679);
nand U1019 (N_1019,N_869,N_705);
nand U1020 (N_1020,N_621,N_954);
and U1021 (N_1021,N_394,N_380);
nor U1022 (N_1022,N_812,N_736);
and U1023 (N_1023,N_317,N_618);
or U1024 (N_1024,N_836,N_474);
nand U1025 (N_1025,N_35,N_619);
nand U1026 (N_1026,N_65,N_498);
nor U1027 (N_1027,N_814,N_67);
nor U1028 (N_1028,N_129,N_238);
nor U1029 (N_1029,N_177,N_439);
xor U1030 (N_1030,N_476,N_239);
or U1031 (N_1031,N_638,N_492);
and U1032 (N_1032,N_354,N_11);
nand U1033 (N_1033,N_456,N_191);
nor U1034 (N_1034,N_668,N_574);
nor U1035 (N_1035,N_213,N_134);
and U1036 (N_1036,N_540,N_811);
or U1037 (N_1037,N_772,N_401);
or U1038 (N_1038,N_405,N_17);
and U1039 (N_1039,N_450,N_9);
nor U1040 (N_1040,N_894,N_925);
or U1041 (N_1041,N_700,N_104);
or U1042 (N_1042,N_607,N_704);
nor U1043 (N_1043,N_54,N_23);
and U1044 (N_1044,N_733,N_852);
or U1045 (N_1045,N_897,N_534);
nor U1046 (N_1046,N_575,N_988);
nand U1047 (N_1047,N_863,N_751);
nor U1048 (N_1048,N_14,N_831);
nand U1049 (N_1049,N_721,N_263);
nor U1050 (N_1050,N_911,N_510);
or U1051 (N_1051,N_907,N_63);
and U1052 (N_1052,N_557,N_385);
nand U1053 (N_1053,N_47,N_291);
nand U1054 (N_1054,N_81,N_313);
xor U1055 (N_1055,N_146,N_411);
or U1056 (N_1056,N_701,N_100);
or U1057 (N_1057,N_403,N_16);
nand U1058 (N_1058,N_79,N_840);
nor U1059 (N_1059,N_678,N_387);
nand U1060 (N_1060,N_523,N_102);
nand U1061 (N_1061,N_130,N_222);
xnor U1062 (N_1062,N_578,N_622);
or U1063 (N_1063,N_981,N_612);
and U1064 (N_1064,N_0,N_650);
xor U1065 (N_1065,N_284,N_475);
xor U1066 (N_1066,N_57,N_333);
xor U1067 (N_1067,N_369,N_583);
xor U1068 (N_1068,N_83,N_173);
or U1069 (N_1069,N_703,N_861);
or U1070 (N_1070,N_508,N_396);
nand U1071 (N_1071,N_410,N_151);
or U1072 (N_1072,N_315,N_659);
or U1073 (N_1073,N_189,N_968);
nor U1074 (N_1074,N_242,N_804);
or U1075 (N_1075,N_728,N_642);
nor U1076 (N_1076,N_725,N_752);
nor U1077 (N_1077,N_902,N_764);
nor U1078 (N_1078,N_867,N_122);
and U1079 (N_1079,N_53,N_368);
nor U1080 (N_1080,N_643,N_494);
nor U1081 (N_1081,N_942,N_967);
and U1082 (N_1082,N_422,N_546);
nor U1083 (N_1083,N_228,N_879);
nand U1084 (N_1084,N_871,N_107);
nand U1085 (N_1085,N_92,N_20);
and U1086 (N_1086,N_535,N_309);
nand U1087 (N_1087,N_155,N_278);
and U1088 (N_1088,N_271,N_485);
or U1089 (N_1089,N_289,N_549);
nand U1090 (N_1090,N_604,N_428);
nand U1091 (N_1091,N_353,N_175);
nor U1092 (N_1092,N_32,N_606);
or U1093 (N_1093,N_215,N_435);
nand U1094 (N_1094,N_868,N_441);
nor U1095 (N_1095,N_221,N_64);
nand U1096 (N_1096,N_331,N_567);
nor U1097 (N_1097,N_220,N_691);
xor U1098 (N_1098,N_795,N_749);
xor U1099 (N_1099,N_468,N_406);
nand U1100 (N_1100,N_181,N_525);
nor U1101 (N_1101,N_998,N_59);
and U1102 (N_1102,N_750,N_71);
or U1103 (N_1103,N_595,N_298);
nand U1104 (N_1104,N_979,N_936);
nand U1105 (N_1105,N_266,N_891);
or U1106 (N_1106,N_788,N_293);
nor U1107 (N_1107,N_496,N_243);
xnor U1108 (N_1108,N_73,N_610);
and U1109 (N_1109,N_671,N_423);
or U1110 (N_1110,N_192,N_794);
or U1111 (N_1111,N_276,N_361);
nand U1112 (N_1112,N_737,N_677);
or U1113 (N_1113,N_778,N_288);
nor U1114 (N_1114,N_538,N_760);
or U1115 (N_1115,N_487,N_835);
and U1116 (N_1116,N_225,N_945);
xnor U1117 (N_1117,N_944,N_247);
xor U1118 (N_1118,N_304,N_766);
or U1119 (N_1119,N_947,N_440);
nor U1120 (N_1120,N_420,N_8);
and U1121 (N_1121,N_555,N_438);
or U1122 (N_1122,N_923,N_543);
and U1123 (N_1123,N_808,N_913);
or U1124 (N_1124,N_886,N_952);
nor U1125 (N_1125,N_996,N_109);
or U1126 (N_1126,N_875,N_388);
nand U1127 (N_1127,N_881,N_273);
or U1128 (N_1128,N_655,N_731);
nor U1129 (N_1129,N_72,N_254);
nand U1130 (N_1130,N_519,N_370);
nor U1131 (N_1131,N_69,N_341);
nand U1132 (N_1132,N_588,N_885);
and U1133 (N_1133,N_183,N_589);
or U1134 (N_1134,N_392,N_218);
and U1135 (N_1135,N_335,N_187);
or U1136 (N_1136,N_290,N_36);
nand U1137 (N_1137,N_38,N_295);
nor U1138 (N_1138,N_268,N_644);
and U1139 (N_1139,N_563,N_532);
and U1140 (N_1140,N_434,N_825);
or U1141 (N_1141,N_142,N_145);
nand U1142 (N_1142,N_929,N_179);
xor U1143 (N_1143,N_900,N_775);
and U1144 (N_1144,N_522,N_623);
nand U1145 (N_1145,N_397,N_986);
and U1146 (N_1146,N_934,N_745);
or U1147 (N_1147,N_161,N_85);
and U1148 (N_1148,N_459,N_157);
and U1149 (N_1149,N_277,N_336);
nor U1150 (N_1150,N_320,N_666);
xnor U1151 (N_1151,N_199,N_648);
nand U1152 (N_1152,N_481,N_138);
or U1153 (N_1153,N_471,N_470);
nand U1154 (N_1154,N_505,N_417);
and U1155 (N_1155,N_915,N_890);
nand U1156 (N_1156,N_372,N_358);
or U1157 (N_1157,N_251,N_553);
nor U1158 (N_1158,N_926,N_383);
xnor U1159 (N_1159,N_51,N_373);
nand U1160 (N_1160,N_586,N_314);
nand U1161 (N_1161,N_973,N_870);
nor U1162 (N_1162,N_250,N_377);
or U1163 (N_1163,N_46,N_174);
or U1164 (N_1164,N_31,N_558);
and U1165 (N_1165,N_139,N_105);
nor U1166 (N_1166,N_918,N_939);
and U1167 (N_1167,N_854,N_948);
nor U1168 (N_1168,N_217,N_489);
nor U1169 (N_1169,N_108,N_582);
and U1170 (N_1170,N_620,N_741);
nand U1171 (N_1171,N_693,N_975);
nor U1172 (N_1172,N_327,N_874);
or U1173 (N_1173,N_796,N_949);
nor U1174 (N_1174,N_303,N_924);
and U1175 (N_1175,N_608,N_374);
xnor U1176 (N_1176,N_33,N_625);
nor U1177 (N_1177,N_119,N_355);
nor U1178 (N_1178,N_415,N_740);
nor U1179 (N_1179,N_882,N_329);
nor U1180 (N_1180,N_371,N_922);
nand U1181 (N_1181,N_163,N_713);
nor U1182 (N_1182,N_779,N_340);
xor U1183 (N_1183,N_91,N_511);
and U1184 (N_1184,N_236,N_860);
and U1185 (N_1185,N_465,N_647);
nor U1186 (N_1186,N_497,N_707);
nor U1187 (N_1187,N_389,N_849);
nand U1188 (N_1188,N_955,N_180);
nand U1189 (N_1189,N_951,N_632);
nand U1190 (N_1190,N_229,N_112);
nor U1191 (N_1191,N_657,N_244);
nand U1192 (N_1192,N_305,N_711);
xor U1193 (N_1193,N_230,N_89);
or U1194 (N_1194,N_483,N_717);
nor U1195 (N_1195,N_531,N_381);
nand U1196 (N_1196,N_363,N_602);
and U1197 (N_1197,N_712,N_654);
or U1198 (N_1198,N_834,N_503);
nand U1199 (N_1199,N_859,N_421);
nor U1200 (N_1200,N_123,N_432);
nor U1201 (N_1201,N_95,N_524);
nor U1202 (N_1202,N_1,N_953);
or U1203 (N_1203,N_302,N_30);
nor U1204 (N_1204,N_253,N_564);
or U1205 (N_1205,N_256,N_568);
or U1206 (N_1206,N_629,N_635);
nor U1207 (N_1207,N_889,N_528);
or U1208 (N_1208,N_837,N_773);
nor U1209 (N_1209,N_708,N_364);
and U1210 (N_1210,N_424,N_530);
or U1211 (N_1211,N_801,N_166);
nor U1212 (N_1212,N_754,N_744);
and U1213 (N_1213,N_670,N_120);
nand U1214 (N_1214,N_444,N_841);
nand U1215 (N_1215,N_93,N_798);
or U1216 (N_1216,N_339,N_790);
nor U1217 (N_1217,N_715,N_547);
xor U1218 (N_1218,N_573,N_910);
nand U1219 (N_1219,N_966,N_656);
nand U1220 (N_1220,N_661,N_997);
or U1221 (N_1221,N_4,N_993);
or U1222 (N_1222,N_90,N_651);
or U1223 (N_1223,N_345,N_931);
nor U1224 (N_1224,N_426,N_819);
nor U1225 (N_1225,N_233,N_560);
or U1226 (N_1226,N_149,N_84);
nand U1227 (N_1227,N_527,N_628);
xor U1228 (N_1228,N_507,N_914);
nor U1229 (N_1229,N_235,N_682);
nand U1230 (N_1230,N_738,N_472);
and U1231 (N_1231,N_807,N_504);
nand U1232 (N_1232,N_594,N_70);
nand U1233 (N_1233,N_198,N_855);
and U1234 (N_1234,N_689,N_137);
nor U1235 (N_1235,N_203,N_714);
and U1236 (N_1236,N_80,N_730);
or U1237 (N_1237,N_539,N_310);
and U1238 (N_1238,N_627,N_709);
nand U1239 (N_1239,N_978,N_941);
nor U1240 (N_1240,N_743,N_828);
or U1241 (N_1241,N_675,N_599);
or U1242 (N_1242,N_436,N_950);
nor U1243 (N_1243,N_280,N_584);
nand U1244 (N_1244,N_696,N_49);
nor U1245 (N_1245,N_958,N_402);
or U1246 (N_1246,N_735,N_272);
and U1247 (N_1247,N_178,N_478);
xor U1248 (N_1248,N_971,N_264);
or U1249 (N_1249,N_851,N_763);
or U1250 (N_1250,N_74,N_660);
nand U1251 (N_1251,N_185,N_147);
or U1252 (N_1252,N_884,N_452);
nand U1253 (N_1253,N_113,N_140);
and U1254 (N_1254,N_495,N_631);
or U1255 (N_1255,N_550,N_316);
nand U1256 (N_1256,N_409,N_159);
and U1257 (N_1257,N_809,N_816);
nor U1258 (N_1258,N_328,N_126);
and U1259 (N_1259,N_210,N_455);
and U1260 (N_1260,N_824,N_769);
and U1261 (N_1261,N_202,N_899);
nand U1262 (N_1262,N_698,N_433);
nand U1263 (N_1263,N_722,N_379);
and U1264 (N_1264,N_541,N_529);
and U1265 (N_1265,N_226,N_269);
and U1266 (N_1266,N_58,N_301);
nor U1267 (N_1267,N_847,N_274);
or U1268 (N_1268,N_992,N_641);
nor U1269 (N_1269,N_308,N_771);
or U1270 (N_1270,N_398,N_937);
and U1271 (N_1271,N_548,N_330);
nor U1272 (N_1272,N_756,N_512);
nand U1273 (N_1273,N_556,N_959);
and U1274 (N_1274,N_674,N_294);
nand U1275 (N_1275,N_633,N_190);
nor U1276 (N_1276,N_904,N_262);
nand U1277 (N_1277,N_160,N_344);
or U1278 (N_1278,N_995,N_878);
nor U1279 (N_1279,N_898,N_820);
or U1280 (N_1280,N_774,N_224);
nand U1281 (N_1281,N_956,N_792);
nor U1282 (N_1282,N_404,N_427);
nand U1283 (N_1283,N_111,N_676);
nand U1284 (N_1284,N_850,N_509);
or U1285 (N_1285,N_591,N_695);
nor U1286 (N_1286,N_117,N_352);
nor U1287 (N_1287,N_357,N_780);
or U1288 (N_1288,N_386,N_818);
and U1289 (N_1289,N_260,N_200);
nand U1290 (N_1290,N_862,N_457);
or U1291 (N_1291,N_152,N_680);
nand U1292 (N_1292,N_480,N_283);
nand U1293 (N_1293,N_34,N_571);
and U1294 (N_1294,N_150,N_227);
or U1295 (N_1295,N_56,N_75);
nand U1296 (N_1296,N_653,N_626);
or U1297 (N_1297,N_990,N_52);
and U1298 (N_1298,N_346,N_3);
xnor U1299 (N_1299,N_669,N_296);
xnor U1300 (N_1300,N_22,N_62);
nor U1301 (N_1301,N_19,N_133);
nand U1302 (N_1302,N_892,N_601);
xnor U1303 (N_1303,N_617,N_630);
and U1304 (N_1304,N_473,N_781);
nand U1305 (N_1305,N_337,N_989);
and U1306 (N_1306,N_148,N_982);
or U1307 (N_1307,N_917,N_935);
and U1308 (N_1308,N_41,N_300);
nor U1309 (N_1309,N_833,N_943);
xnor U1310 (N_1310,N_970,N_580);
nor U1311 (N_1311,N_10,N_103);
xnor U1312 (N_1312,N_901,N_165);
xor U1313 (N_1313,N_141,N_976);
nand U1314 (N_1314,N_613,N_611);
or U1315 (N_1315,N_864,N_526);
nor U1316 (N_1316,N_13,N_603);
nor U1317 (N_1317,N_68,N_797);
nor U1318 (N_1318,N_219,N_464);
nor U1319 (N_1319,N_125,N_482);
or U1320 (N_1320,N_21,N_267);
xor U1321 (N_1321,N_282,N_765);
or U1322 (N_1322,N_24,N_193);
nor U1323 (N_1323,N_762,N_286);
or U1324 (N_1324,N_326,N_645);
nand U1325 (N_1325,N_43,N_7);
or U1326 (N_1326,N_920,N_872);
or U1327 (N_1327,N_961,N_697);
or U1328 (N_1328,N_437,N_376);
nor U1329 (N_1329,N_592,N_318);
nand U1330 (N_1330,N_261,N_516);
and U1331 (N_1331,N_930,N_742);
and U1332 (N_1332,N_776,N_972);
or U1333 (N_1333,N_206,N_249);
nor U1334 (N_1334,N_817,N_856);
and U1335 (N_1335,N_727,N_395);
or U1336 (N_1336,N_170,N_158);
or U1337 (N_1337,N_66,N_969);
or U1338 (N_1338,N_431,N_977);
or U1339 (N_1339,N_739,N_581);
and U1340 (N_1340,N_815,N_28);
xnor U1341 (N_1341,N_806,N_297);
nor U1342 (N_1342,N_755,N_813);
nor U1343 (N_1343,N_895,N_240);
nand U1344 (N_1344,N_466,N_40);
or U1345 (N_1345,N_685,N_597);
and U1346 (N_1346,N_803,N_999);
or U1347 (N_1347,N_590,N_26);
nor U1348 (N_1348,N_419,N_609);
or U1349 (N_1349,N_131,N_848);
or U1350 (N_1350,N_462,N_706);
or U1351 (N_1351,N_365,N_367);
or U1352 (N_1352,N_843,N_39);
nand U1353 (N_1353,N_502,N_552);
and U1354 (N_1354,N_248,N_658);
nor U1355 (N_1355,N_164,N_275);
or U1356 (N_1356,N_957,N_561);
nor U1357 (N_1357,N_454,N_127);
nand U1358 (N_1358,N_829,N_646);
nand U1359 (N_1359,N_167,N_533);
nand U1360 (N_1360,N_97,N_2);
or U1361 (N_1361,N_723,N_292);
and U1362 (N_1362,N_873,N_888);
nor U1363 (N_1363,N_514,N_614);
or U1364 (N_1364,N_176,N_279);
xnor U1365 (N_1365,N_694,N_784);
and U1366 (N_1366,N_799,N_938);
xnor U1367 (N_1367,N_839,N_234);
or U1368 (N_1368,N_5,N_810);
nor U1369 (N_1369,N_416,N_446);
or U1370 (N_1370,N_463,N_299);
nand U1371 (N_1371,N_338,N_866);
or U1372 (N_1372,N_325,N_761);
nor U1373 (N_1373,N_585,N_838);
xnor U1374 (N_1374,N_12,N_445);
or U1375 (N_1375,N_342,N_285);
xnor U1376 (N_1376,N_307,N_201);
or U1377 (N_1377,N_237,N_55);
and U1378 (N_1378,N_759,N_827);
nand U1379 (N_1379,N_566,N_334);
nand U1380 (N_1380,N_29,N_212);
xnor U1381 (N_1381,N_718,N_517);
nor U1382 (N_1382,N_724,N_281);
nor U1383 (N_1383,N_893,N_600);
and U1384 (N_1384,N_257,N_570);
nand U1385 (N_1385,N_143,N_50);
or U1386 (N_1386,N_323,N_734);
or U1387 (N_1387,N_903,N_664);
or U1388 (N_1388,N_746,N_132);
or U1389 (N_1389,N_171,N_683);
and U1390 (N_1390,N_121,N_115);
nand U1391 (N_1391,N_182,N_593);
xnor U1392 (N_1392,N_110,N_906);
and U1393 (N_1393,N_758,N_425);
nand U1394 (N_1394,N_479,N_783);
nor U1395 (N_1395,N_60,N_554);
nand U1396 (N_1396,N_702,N_76);
nor U1397 (N_1397,N_576,N_493);
nand U1398 (N_1398,N_259,N_965);
nand U1399 (N_1399,N_545,N_412);
nor U1400 (N_1400,N_767,N_27);
nand U1401 (N_1401,N_865,N_486);
nor U1402 (N_1402,N_88,N_399);
nand U1403 (N_1403,N_324,N_306);
or U1404 (N_1404,N_681,N_467);
xnor U1405 (N_1405,N_544,N_82);
xnor U1406 (N_1406,N_846,N_343);
nand U1407 (N_1407,N_18,N_673);
and U1408 (N_1408,N_747,N_984);
and U1409 (N_1409,N_805,N_499);
nor U1410 (N_1410,N_241,N_729);
nor U1411 (N_1411,N_753,N_429);
nor U1412 (N_1412,N_114,N_946);
or U1413 (N_1413,N_87,N_572);
or U1414 (N_1414,N_985,N_687);
nor U1415 (N_1415,N_214,N_6);
or U1416 (N_1416,N_665,N_559);
or U1417 (N_1417,N_932,N_94);
xnor U1418 (N_1418,N_186,N_216);
and U1419 (N_1419,N_782,N_359);
and U1420 (N_1420,N_321,N_366);
and U1421 (N_1421,N_506,N_270);
nand U1422 (N_1422,N_347,N_640);
or U1423 (N_1423,N_15,N_853);
and U1424 (N_1424,N_245,N_800);
and U1425 (N_1425,N_598,N_414);
nor U1426 (N_1426,N_537,N_255);
and U1427 (N_1427,N_719,N_390);
and U1428 (N_1428,N_77,N_802);
or U1429 (N_1429,N_789,N_960);
nor U1430 (N_1430,N_172,N_188);
nand U1431 (N_1431,N_349,N_624);
nor U1432 (N_1432,N_876,N_461);
xor U1433 (N_1433,N_562,N_686);
xor U1434 (N_1434,N_135,N_44);
or U1435 (N_1435,N_61,N_136);
or U1436 (N_1436,N_209,N_513);
or U1437 (N_1437,N_484,N_393);
nor U1438 (N_1438,N_144,N_37);
or U1439 (N_1439,N_994,N_663);
nor U1440 (N_1440,N_196,N_375);
xnor U1441 (N_1441,N_912,N_726);
nand U1442 (N_1442,N_720,N_116);
and U1443 (N_1443,N_211,N_830);
or U1444 (N_1444,N_905,N_319);
nor U1445 (N_1445,N_447,N_350);
and U1446 (N_1446,N_787,N_928);
nand U1447 (N_1447,N_154,N_822);
or U1448 (N_1448,N_362,N_962);
nand U1449 (N_1449,N_246,N_652);
or U1450 (N_1450,N_987,N_832);
or U1451 (N_1451,N_418,N_521);
and U1452 (N_1452,N_106,N_312);
nand U1453 (N_1453,N_845,N_356);
nand U1454 (N_1454,N_615,N_637);
nor U1455 (N_1455,N_207,N_551);
xnor U1456 (N_1456,N_844,N_983);
and U1457 (N_1457,N_690,N_791);
nand U1458 (N_1458,N_400,N_672);
nor U1459 (N_1459,N_963,N_569);
nor U1460 (N_1460,N_184,N_258);
or U1461 (N_1461,N_515,N_48);
or U1462 (N_1462,N_684,N_477);
or U1463 (N_1463,N_382,N_710);
or U1464 (N_1464,N_768,N_491);
nand U1465 (N_1465,N_980,N_332);
or U1466 (N_1466,N_823,N_748);
nor U1467 (N_1467,N_408,N_577);
nor U1468 (N_1468,N_858,N_265);
nand U1469 (N_1469,N_98,N_909);
nand U1470 (N_1470,N_777,N_469);
or U1471 (N_1471,N_458,N_194);
and U1472 (N_1472,N_692,N_351);
nor U1473 (N_1473,N_448,N_162);
nand U1474 (N_1474,N_785,N_716);
xnor U1475 (N_1475,N_311,N_770);
nand U1476 (N_1476,N_384,N_605);
nor U1477 (N_1477,N_880,N_156);
and U1478 (N_1478,N_793,N_649);
nand U1479 (N_1479,N_634,N_391);
and U1480 (N_1480,N_118,N_662);
xnor U1481 (N_1481,N_443,N_518);
or U1482 (N_1482,N_639,N_78);
xnor U1483 (N_1483,N_128,N_223);
nor U1484 (N_1484,N_501,N_168);
or U1485 (N_1485,N_887,N_699);
nor U1486 (N_1486,N_667,N_25);
or U1487 (N_1487,N_460,N_821);
nor U1488 (N_1488,N_287,N_536);
nand U1489 (N_1489,N_378,N_896);
and U1490 (N_1490,N_451,N_940);
or U1491 (N_1491,N_430,N_208);
or U1492 (N_1492,N_565,N_153);
nor U1493 (N_1493,N_490,N_616);
and U1494 (N_1494,N_688,N_579);
or U1495 (N_1495,N_442,N_322);
or U1496 (N_1496,N_99,N_45);
nor U1497 (N_1497,N_124,N_413);
xnor U1498 (N_1498,N_921,N_596);
nor U1499 (N_1499,N_232,N_449);
or U1500 (N_1500,N_70,N_859);
nor U1501 (N_1501,N_496,N_579);
nand U1502 (N_1502,N_387,N_219);
and U1503 (N_1503,N_333,N_74);
nor U1504 (N_1504,N_806,N_428);
nand U1505 (N_1505,N_296,N_996);
nor U1506 (N_1506,N_227,N_386);
nor U1507 (N_1507,N_789,N_558);
and U1508 (N_1508,N_589,N_981);
nor U1509 (N_1509,N_76,N_443);
xor U1510 (N_1510,N_655,N_286);
nor U1511 (N_1511,N_962,N_672);
or U1512 (N_1512,N_346,N_202);
nor U1513 (N_1513,N_205,N_534);
or U1514 (N_1514,N_807,N_626);
and U1515 (N_1515,N_380,N_305);
xnor U1516 (N_1516,N_32,N_978);
or U1517 (N_1517,N_488,N_142);
nor U1518 (N_1518,N_380,N_114);
nand U1519 (N_1519,N_788,N_10);
xor U1520 (N_1520,N_457,N_445);
xnor U1521 (N_1521,N_885,N_661);
nor U1522 (N_1522,N_281,N_900);
xnor U1523 (N_1523,N_516,N_279);
nand U1524 (N_1524,N_456,N_102);
nand U1525 (N_1525,N_597,N_716);
nand U1526 (N_1526,N_594,N_632);
nor U1527 (N_1527,N_220,N_647);
or U1528 (N_1528,N_544,N_445);
and U1529 (N_1529,N_3,N_997);
and U1530 (N_1530,N_716,N_137);
and U1531 (N_1531,N_19,N_706);
nand U1532 (N_1532,N_248,N_663);
or U1533 (N_1533,N_841,N_654);
or U1534 (N_1534,N_677,N_695);
or U1535 (N_1535,N_184,N_19);
or U1536 (N_1536,N_134,N_265);
xor U1537 (N_1537,N_409,N_407);
nor U1538 (N_1538,N_936,N_720);
nor U1539 (N_1539,N_224,N_223);
or U1540 (N_1540,N_51,N_358);
xnor U1541 (N_1541,N_64,N_200);
nand U1542 (N_1542,N_890,N_398);
or U1543 (N_1543,N_843,N_510);
nand U1544 (N_1544,N_661,N_901);
nand U1545 (N_1545,N_642,N_381);
nor U1546 (N_1546,N_883,N_980);
nor U1547 (N_1547,N_965,N_600);
and U1548 (N_1548,N_235,N_156);
nor U1549 (N_1549,N_531,N_521);
or U1550 (N_1550,N_968,N_760);
nand U1551 (N_1551,N_661,N_194);
and U1552 (N_1552,N_427,N_653);
xor U1553 (N_1553,N_327,N_316);
nand U1554 (N_1554,N_895,N_822);
nor U1555 (N_1555,N_216,N_563);
nand U1556 (N_1556,N_700,N_976);
and U1557 (N_1557,N_993,N_113);
and U1558 (N_1558,N_61,N_793);
or U1559 (N_1559,N_503,N_351);
nor U1560 (N_1560,N_4,N_549);
and U1561 (N_1561,N_250,N_537);
nand U1562 (N_1562,N_143,N_565);
nand U1563 (N_1563,N_458,N_130);
and U1564 (N_1564,N_690,N_73);
nand U1565 (N_1565,N_761,N_467);
nor U1566 (N_1566,N_829,N_61);
xor U1567 (N_1567,N_918,N_176);
xor U1568 (N_1568,N_266,N_990);
nand U1569 (N_1569,N_410,N_920);
or U1570 (N_1570,N_677,N_333);
nor U1571 (N_1571,N_368,N_839);
and U1572 (N_1572,N_760,N_919);
and U1573 (N_1573,N_651,N_219);
nor U1574 (N_1574,N_488,N_986);
nand U1575 (N_1575,N_650,N_43);
nand U1576 (N_1576,N_447,N_433);
or U1577 (N_1577,N_792,N_945);
nand U1578 (N_1578,N_285,N_740);
and U1579 (N_1579,N_957,N_103);
nand U1580 (N_1580,N_311,N_240);
nand U1581 (N_1581,N_168,N_432);
nand U1582 (N_1582,N_133,N_320);
nor U1583 (N_1583,N_709,N_970);
and U1584 (N_1584,N_578,N_376);
or U1585 (N_1585,N_322,N_99);
and U1586 (N_1586,N_413,N_465);
and U1587 (N_1587,N_510,N_317);
and U1588 (N_1588,N_301,N_841);
and U1589 (N_1589,N_352,N_423);
nor U1590 (N_1590,N_399,N_250);
nand U1591 (N_1591,N_319,N_888);
or U1592 (N_1592,N_682,N_168);
nor U1593 (N_1593,N_493,N_212);
and U1594 (N_1594,N_32,N_902);
nor U1595 (N_1595,N_709,N_899);
and U1596 (N_1596,N_765,N_175);
and U1597 (N_1597,N_887,N_228);
xor U1598 (N_1598,N_794,N_590);
and U1599 (N_1599,N_79,N_954);
and U1600 (N_1600,N_899,N_696);
or U1601 (N_1601,N_510,N_102);
or U1602 (N_1602,N_3,N_97);
or U1603 (N_1603,N_969,N_988);
or U1604 (N_1604,N_656,N_705);
or U1605 (N_1605,N_144,N_513);
nor U1606 (N_1606,N_817,N_458);
nand U1607 (N_1607,N_573,N_484);
nand U1608 (N_1608,N_168,N_724);
and U1609 (N_1609,N_898,N_27);
xnor U1610 (N_1610,N_498,N_943);
nor U1611 (N_1611,N_839,N_185);
xnor U1612 (N_1612,N_171,N_858);
nor U1613 (N_1613,N_629,N_781);
and U1614 (N_1614,N_39,N_361);
nor U1615 (N_1615,N_831,N_535);
and U1616 (N_1616,N_371,N_770);
or U1617 (N_1617,N_597,N_653);
and U1618 (N_1618,N_887,N_362);
or U1619 (N_1619,N_786,N_982);
and U1620 (N_1620,N_118,N_885);
and U1621 (N_1621,N_569,N_974);
and U1622 (N_1622,N_719,N_599);
and U1623 (N_1623,N_377,N_758);
and U1624 (N_1624,N_393,N_667);
nor U1625 (N_1625,N_45,N_994);
nor U1626 (N_1626,N_513,N_115);
nand U1627 (N_1627,N_554,N_763);
or U1628 (N_1628,N_850,N_99);
and U1629 (N_1629,N_768,N_791);
or U1630 (N_1630,N_43,N_953);
xor U1631 (N_1631,N_827,N_961);
or U1632 (N_1632,N_364,N_596);
nor U1633 (N_1633,N_957,N_579);
xnor U1634 (N_1634,N_353,N_303);
nand U1635 (N_1635,N_124,N_395);
nand U1636 (N_1636,N_259,N_413);
nor U1637 (N_1637,N_515,N_626);
nor U1638 (N_1638,N_990,N_914);
nand U1639 (N_1639,N_906,N_446);
nor U1640 (N_1640,N_989,N_519);
and U1641 (N_1641,N_527,N_407);
or U1642 (N_1642,N_622,N_612);
xor U1643 (N_1643,N_793,N_694);
and U1644 (N_1644,N_113,N_583);
nand U1645 (N_1645,N_312,N_507);
nand U1646 (N_1646,N_11,N_457);
nor U1647 (N_1647,N_495,N_999);
or U1648 (N_1648,N_535,N_501);
nand U1649 (N_1649,N_930,N_107);
and U1650 (N_1650,N_197,N_12);
nor U1651 (N_1651,N_212,N_552);
nand U1652 (N_1652,N_197,N_644);
and U1653 (N_1653,N_169,N_639);
and U1654 (N_1654,N_166,N_926);
xor U1655 (N_1655,N_594,N_978);
nor U1656 (N_1656,N_779,N_428);
and U1657 (N_1657,N_298,N_664);
nor U1658 (N_1658,N_672,N_0);
and U1659 (N_1659,N_264,N_639);
and U1660 (N_1660,N_795,N_107);
and U1661 (N_1661,N_417,N_822);
nor U1662 (N_1662,N_284,N_894);
and U1663 (N_1663,N_541,N_893);
or U1664 (N_1664,N_684,N_261);
and U1665 (N_1665,N_223,N_74);
nand U1666 (N_1666,N_672,N_854);
and U1667 (N_1667,N_396,N_393);
and U1668 (N_1668,N_384,N_621);
or U1669 (N_1669,N_461,N_256);
xnor U1670 (N_1670,N_556,N_243);
xnor U1671 (N_1671,N_293,N_486);
or U1672 (N_1672,N_632,N_758);
and U1673 (N_1673,N_938,N_218);
nand U1674 (N_1674,N_210,N_385);
xnor U1675 (N_1675,N_943,N_496);
and U1676 (N_1676,N_567,N_427);
or U1677 (N_1677,N_88,N_245);
or U1678 (N_1678,N_214,N_769);
nor U1679 (N_1679,N_267,N_992);
nand U1680 (N_1680,N_167,N_466);
and U1681 (N_1681,N_861,N_450);
nand U1682 (N_1682,N_688,N_545);
nand U1683 (N_1683,N_55,N_570);
nand U1684 (N_1684,N_851,N_301);
nor U1685 (N_1685,N_692,N_377);
or U1686 (N_1686,N_58,N_552);
nand U1687 (N_1687,N_5,N_946);
xor U1688 (N_1688,N_165,N_32);
nand U1689 (N_1689,N_694,N_586);
nor U1690 (N_1690,N_896,N_540);
nor U1691 (N_1691,N_257,N_863);
and U1692 (N_1692,N_907,N_590);
and U1693 (N_1693,N_905,N_892);
and U1694 (N_1694,N_577,N_696);
nor U1695 (N_1695,N_588,N_776);
nand U1696 (N_1696,N_726,N_590);
nand U1697 (N_1697,N_639,N_811);
or U1698 (N_1698,N_684,N_64);
nor U1699 (N_1699,N_228,N_531);
nand U1700 (N_1700,N_962,N_96);
nand U1701 (N_1701,N_310,N_138);
nand U1702 (N_1702,N_440,N_667);
or U1703 (N_1703,N_506,N_841);
nor U1704 (N_1704,N_787,N_615);
or U1705 (N_1705,N_635,N_562);
or U1706 (N_1706,N_573,N_616);
xnor U1707 (N_1707,N_6,N_566);
nand U1708 (N_1708,N_65,N_676);
and U1709 (N_1709,N_20,N_141);
nand U1710 (N_1710,N_933,N_766);
and U1711 (N_1711,N_281,N_222);
and U1712 (N_1712,N_536,N_186);
or U1713 (N_1713,N_24,N_167);
or U1714 (N_1714,N_368,N_585);
xor U1715 (N_1715,N_217,N_267);
and U1716 (N_1716,N_264,N_841);
nor U1717 (N_1717,N_877,N_196);
or U1718 (N_1718,N_276,N_86);
xor U1719 (N_1719,N_771,N_550);
nand U1720 (N_1720,N_60,N_584);
xnor U1721 (N_1721,N_89,N_556);
and U1722 (N_1722,N_425,N_828);
or U1723 (N_1723,N_372,N_794);
nor U1724 (N_1724,N_835,N_272);
xor U1725 (N_1725,N_912,N_49);
nor U1726 (N_1726,N_589,N_50);
and U1727 (N_1727,N_515,N_621);
or U1728 (N_1728,N_216,N_925);
or U1729 (N_1729,N_506,N_27);
nor U1730 (N_1730,N_436,N_442);
or U1731 (N_1731,N_884,N_673);
or U1732 (N_1732,N_366,N_815);
nor U1733 (N_1733,N_88,N_972);
nand U1734 (N_1734,N_309,N_556);
nor U1735 (N_1735,N_282,N_357);
or U1736 (N_1736,N_767,N_849);
nor U1737 (N_1737,N_686,N_843);
and U1738 (N_1738,N_490,N_356);
or U1739 (N_1739,N_989,N_653);
and U1740 (N_1740,N_557,N_774);
nand U1741 (N_1741,N_344,N_227);
xor U1742 (N_1742,N_312,N_594);
xor U1743 (N_1743,N_760,N_59);
nor U1744 (N_1744,N_15,N_827);
nand U1745 (N_1745,N_743,N_742);
and U1746 (N_1746,N_503,N_652);
and U1747 (N_1747,N_737,N_282);
xnor U1748 (N_1748,N_748,N_67);
nand U1749 (N_1749,N_537,N_25);
or U1750 (N_1750,N_651,N_831);
xnor U1751 (N_1751,N_203,N_512);
and U1752 (N_1752,N_345,N_550);
nand U1753 (N_1753,N_188,N_253);
or U1754 (N_1754,N_827,N_435);
nor U1755 (N_1755,N_14,N_546);
xnor U1756 (N_1756,N_147,N_657);
nor U1757 (N_1757,N_756,N_344);
or U1758 (N_1758,N_219,N_922);
nand U1759 (N_1759,N_666,N_203);
and U1760 (N_1760,N_933,N_5);
nor U1761 (N_1761,N_672,N_980);
nand U1762 (N_1762,N_496,N_769);
nand U1763 (N_1763,N_173,N_111);
nand U1764 (N_1764,N_122,N_131);
nor U1765 (N_1765,N_172,N_454);
or U1766 (N_1766,N_479,N_757);
xor U1767 (N_1767,N_438,N_527);
or U1768 (N_1768,N_636,N_317);
nor U1769 (N_1769,N_818,N_539);
nor U1770 (N_1770,N_139,N_158);
nand U1771 (N_1771,N_483,N_341);
xnor U1772 (N_1772,N_353,N_448);
or U1773 (N_1773,N_421,N_932);
or U1774 (N_1774,N_720,N_980);
nor U1775 (N_1775,N_662,N_70);
nand U1776 (N_1776,N_909,N_561);
and U1777 (N_1777,N_206,N_676);
nor U1778 (N_1778,N_852,N_541);
nand U1779 (N_1779,N_364,N_382);
and U1780 (N_1780,N_341,N_871);
and U1781 (N_1781,N_45,N_543);
and U1782 (N_1782,N_259,N_681);
nand U1783 (N_1783,N_522,N_592);
and U1784 (N_1784,N_537,N_942);
nor U1785 (N_1785,N_664,N_377);
xnor U1786 (N_1786,N_4,N_814);
or U1787 (N_1787,N_155,N_626);
nand U1788 (N_1788,N_185,N_139);
nor U1789 (N_1789,N_250,N_678);
or U1790 (N_1790,N_954,N_155);
nand U1791 (N_1791,N_942,N_511);
and U1792 (N_1792,N_372,N_752);
nor U1793 (N_1793,N_273,N_621);
nor U1794 (N_1794,N_54,N_996);
and U1795 (N_1795,N_952,N_341);
nor U1796 (N_1796,N_586,N_216);
and U1797 (N_1797,N_65,N_142);
nor U1798 (N_1798,N_374,N_650);
and U1799 (N_1799,N_363,N_199);
or U1800 (N_1800,N_240,N_106);
or U1801 (N_1801,N_958,N_701);
nor U1802 (N_1802,N_190,N_460);
nand U1803 (N_1803,N_648,N_133);
xor U1804 (N_1804,N_434,N_856);
nor U1805 (N_1805,N_652,N_883);
and U1806 (N_1806,N_783,N_437);
nor U1807 (N_1807,N_236,N_311);
nand U1808 (N_1808,N_767,N_208);
or U1809 (N_1809,N_462,N_14);
nand U1810 (N_1810,N_222,N_376);
nor U1811 (N_1811,N_380,N_466);
or U1812 (N_1812,N_129,N_398);
nand U1813 (N_1813,N_215,N_540);
and U1814 (N_1814,N_769,N_43);
or U1815 (N_1815,N_402,N_128);
nand U1816 (N_1816,N_735,N_907);
nand U1817 (N_1817,N_848,N_451);
or U1818 (N_1818,N_674,N_450);
or U1819 (N_1819,N_550,N_254);
and U1820 (N_1820,N_449,N_625);
and U1821 (N_1821,N_844,N_904);
xnor U1822 (N_1822,N_163,N_466);
or U1823 (N_1823,N_294,N_650);
nand U1824 (N_1824,N_94,N_913);
or U1825 (N_1825,N_820,N_743);
nor U1826 (N_1826,N_978,N_982);
or U1827 (N_1827,N_876,N_119);
nand U1828 (N_1828,N_715,N_801);
and U1829 (N_1829,N_651,N_393);
xor U1830 (N_1830,N_439,N_979);
or U1831 (N_1831,N_761,N_831);
and U1832 (N_1832,N_449,N_601);
nand U1833 (N_1833,N_707,N_17);
nor U1834 (N_1834,N_524,N_568);
nor U1835 (N_1835,N_466,N_72);
nor U1836 (N_1836,N_882,N_610);
nand U1837 (N_1837,N_321,N_142);
nand U1838 (N_1838,N_186,N_134);
and U1839 (N_1839,N_343,N_774);
or U1840 (N_1840,N_748,N_546);
nor U1841 (N_1841,N_702,N_315);
nor U1842 (N_1842,N_186,N_870);
xor U1843 (N_1843,N_469,N_379);
xor U1844 (N_1844,N_595,N_578);
nor U1845 (N_1845,N_396,N_262);
or U1846 (N_1846,N_973,N_846);
nor U1847 (N_1847,N_18,N_819);
nand U1848 (N_1848,N_533,N_320);
nor U1849 (N_1849,N_467,N_765);
or U1850 (N_1850,N_53,N_471);
and U1851 (N_1851,N_670,N_288);
nor U1852 (N_1852,N_535,N_51);
and U1853 (N_1853,N_954,N_449);
xnor U1854 (N_1854,N_225,N_260);
nand U1855 (N_1855,N_935,N_211);
and U1856 (N_1856,N_34,N_354);
xnor U1857 (N_1857,N_97,N_176);
or U1858 (N_1858,N_391,N_750);
nor U1859 (N_1859,N_815,N_377);
and U1860 (N_1860,N_488,N_79);
nand U1861 (N_1861,N_538,N_576);
or U1862 (N_1862,N_596,N_861);
nand U1863 (N_1863,N_122,N_13);
or U1864 (N_1864,N_971,N_929);
or U1865 (N_1865,N_91,N_683);
or U1866 (N_1866,N_825,N_598);
nand U1867 (N_1867,N_778,N_257);
nor U1868 (N_1868,N_895,N_573);
and U1869 (N_1869,N_158,N_799);
nor U1870 (N_1870,N_488,N_290);
xor U1871 (N_1871,N_731,N_777);
nor U1872 (N_1872,N_565,N_278);
and U1873 (N_1873,N_712,N_929);
xnor U1874 (N_1874,N_679,N_277);
and U1875 (N_1875,N_613,N_655);
nor U1876 (N_1876,N_876,N_411);
nor U1877 (N_1877,N_801,N_432);
nor U1878 (N_1878,N_931,N_551);
and U1879 (N_1879,N_168,N_121);
nor U1880 (N_1880,N_405,N_732);
and U1881 (N_1881,N_689,N_59);
and U1882 (N_1882,N_851,N_421);
xor U1883 (N_1883,N_188,N_880);
and U1884 (N_1884,N_646,N_83);
and U1885 (N_1885,N_925,N_554);
nand U1886 (N_1886,N_729,N_418);
and U1887 (N_1887,N_930,N_255);
nand U1888 (N_1888,N_770,N_68);
nor U1889 (N_1889,N_201,N_633);
nand U1890 (N_1890,N_375,N_148);
xor U1891 (N_1891,N_627,N_567);
nor U1892 (N_1892,N_142,N_995);
xor U1893 (N_1893,N_695,N_797);
or U1894 (N_1894,N_373,N_198);
and U1895 (N_1895,N_83,N_917);
or U1896 (N_1896,N_858,N_457);
or U1897 (N_1897,N_654,N_880);
and U1898 (N_1898,N_594,N_243);
nor U1899 (N_1899,N_714,N_712);
nor U1900 (N_1900,N_674,N_381);
or U1901 (N_1901,N_848,N_569);
and U1902 (N_1902,N_656,N_333);
nand U1903 (N_1903,N_486,N_468);
xnor U1904 (N_1904,N_964,N_595);
and U1905 (N_1905,N_115,N_435);
nand U1906 (N_1906,N_278,N_794);
nand U1907 (N_1907,N_333,N_43);
nor U1908 (N_1908,N_374,N_933);
nand U1909 (N_1909,N_844,N_49);
and U1910 (N_1910,N_276,N_957);
nand U1911 (N_1911,N_935,N_426);
or U1912 (N_1912,N_198,N_451);
or U1913 (N_1913,N_915,N_274);
nor U1914 (N_1914,N_674,N_406);
nand U1915 (N_1915,N_364,N_257);
nor U1916 (N_1916,N_819,N_680);
and U1917 (N_1917,N_362,N_922);
nand U1918 (N_1918,N_564,N_466);
nand U1919 (N_1919,N_762,N_977);
nand U1920 (N_1920,N_291,N_659);
or U1921 (N_1921,N_181,N_855);
nand U1922 (N_1922,N_667,N_146);
nand U1923 (N_1923,N_104,N_747);
and U1924 (N_1924,N_636,N_65);
nand U1925 (N_1925,N_88,N_6);
nand U1926 (N_1926,N_564,N_871);
and U1927 (N_1927,N_55,N_225);
nor U1928 (N_1928,N_284,N_810);
or U1929 (N_1929,N_130,N_121);
or U1930 (N_1930,N_952,N_300);
nand U1931 (N_1931,N_633,N_228);
nor U1932 (N_1932,N_733,N_881);
nand U1933 (N_1933,N_576,N_571);
nand U1934 (N_1934,N_751,N_297);
or U1935 (N_1935,N_990,N_655);
nor U1936 (N_1936,N_998,N_566);
or U1937 (N_1937,N_353,N_593);
and U1938 (N_1938,N_521,N_357);
and U1939 (N_1939,N_778,N_95);
and U1940 (N_1940,N_571,N_134);
nor U1941 (N_1941,N_552,N_618);
nor U1942 (N_1942,N_376,N_753);
or U1943 (N_1943,N_478,N_204);
nand U1944 (N_1944,N_729,N_806);
and U1945 (N_1945,N_294,N_52);
nor U1946 (N_1946,N_429,N_107);
nand U1947 (N_1947,N_84,N_566);
xor U1948 (N_1948,N_732,N_841);
nand U1949 (N_1949,N_501,N_714);
and U1950 (N_1950,N_160,N_432);
xor U1951 (N_1951,N_84,N_948);
nand U1952 (N_1952,N_436,N_532);
and U1953 (N_1953,N_151,N_652);
or U1954 (N_1954,N_133,N_313);
xor U1955 (N_1955,N_957,N_552);
and U1956 (N_1956,N_48,N_47);
or U1957 (N_1957,N_610,N_624);
or U1958 (N_1958,N_872,N_287);
and U1959 (N_1959,N_809,N_794);
or U1960 (N_1960,N_662,N_632);
xor U1961 (N_1961,N_9,N_329);
and U1962 (N_1962,N_265,N_144);
or U1963 (N_1963,N_666,N_847);
nor U1964 (N_1964,N_178,N_601);
nor U1965 (N_1965,N_606,N_224);
or U1966 (N_1966,N_74,N_36);
nor U1967 (N_1967,N_781,N_699);
nor U1968 (N_1968,N_475,N_958);
and U1969 (N_1969,N_375,N_737);
nand U1970 (N_1970,N_456,N_117);
or U1971 (N_1971,N_896,N_683);
and U1972 (N_1972,N_255,N_523);
or U1973 (N_1973,N_706,N_852);
and U1974 (N_1974,N_326,N_574);
and U1975 (N_1975,N_0,N_448);
or U1976 (N_1976,N_782,N_121);
and U1977 (N_1977,N_151,N_533);
or U1978 (N_1978,N_915,N_466);
or U1979 (N_1979,N_696,N_144);
nor U1980 (N_1980,N_512,N_160);
nor U1981 (N_1981,N_715,N_285);
and U1982 (N_1982,N_197,N_398);
nor U1983 (N_1983,N_527,N_697);
nor U1984 (N_1984,N_974,N_851);
nor U1985 (N_1985,N_670,N_798);
nor U1986 (N_1986,N_621,N_884);
nor U1987 (N_1987,N_815,N_612);
or U1988 (N_1988,N_881,N_230);
nand U1989 (N_1989,N_210,N_610);
nor U1990 (N_1990,N_724,N_321);
or U1991 (N_1991,N_311,N_108);
and U1992 (N_1992,N_957,N_92);
nor U1993 (N_1993,N_754,N_114);
and U1994 (N_1994,N_180,N_377);
or U1995 (N_1995,N_825,N_903);
or U1996 (N_1996,N_146,N_245);
or U1997 (N_1997,N_872,N_948);
nand U1998 (N_1998,N_652,N_540);
and U1999 (N_1999,N_49,N_492);
and U2000 (N_2000,N_1341,N_1099);
nand U2001 (N_2001,N_1582,N_1411);
and U2002 (N_2002,N_1236,N_1635);
or U2003 (N_2003,N_1401,N_1052);
and U2004 (N_2004,N_1436,N_1804);
xnor U2005 (N_2005,N_1239,N_1329);
and U2006 (N_2006,N_1038,N_1039);
or U2007 (N_2007,N_1233,N_1928);
nor U2008 (N_2008,N_1667,N_1805);
or U2009 (N_2009,N_1322,N_1979);
nand U2010 (N_2010,N_1083,N_1189);
nand U2011 (N_2011,N_1725,N_1969);
and U2012 (N_2012,N_1927,N_1556);
nor U2013 (N_2013,N_1658,N_1656);
or U2014 (N_2014,N_1823,N_1109);
and U2015 (N_2015,N_1758,N_1707);
and U2016 (N_2016,N_1946,N_1594);
and U2017 (N_2017,N_1032,N_1248);
or U2018 (N_2018,N_1954,N_1179);
or U2019 (N_2019,N_1832,N_1220);
nor U2020 (N_2020,N_1947,N_1950);
xnor U2021 (N_2021,N_1791,N_1546);
or U2022 (N_2022,N_1394,N_1535);
and U2023 (N_2023,N_1747,N_1173);
and U2024 (N_2024,N_1020,N_1323);
nor U2025 (N_2025,N_1042,N_1757);
xnor U2026 (N_2026,N_1112,N_1653);
nand U2027 (N_2027,N_1922,N_1122);
nand U2028 (N_2028,N_1751,N_1129);
or U2029 (N_2029,N_1944,N_1466);
and U2030 (N_2030,N_1385,N_1524);
nor U2031 (N_2031,N_1822,N_1696);
nand U2032 (N_2032,N_1160,N_1448);
nor U2033 (N_2033,N_1602,N_1544);
or U2034 (N_2034,N_1313,N_1028);
nand U2035 (N_2035,N_1593,N_1507);
or U2036 (N_2036,N_1825,N_1506);
nor U2037 (N_2037,N_1100,N_1939);
nor U2038 (N_2038,N_1429,N_1228);
nand U2039 (N_2039,N_1999,N_1242);
nand U2040 (N_2040,N_1205,N_1362);
or U2041 (N_2041,N_1257,N_1246);
or U2042 (N_2042,N_1186,N_1365);
or U2043 (N_2043,N_1345,N_1245);
and U2044 (N_2044,N_1679,N_1421);
nand U2045 (N_2045,N_1354,N_1631);
nand U2046 (N_2046,N_1607,N_1624);
or U2047 (N_2047,N_1292,N_1533);
nand U2048 (N_2048,N_1244,N_1495);
and U2049 (N_2049,N_1647,N_1092);
nor U2050 (N_2050,N_1929,N_1131);
nand U2051 (N_2051,N_1991,N_1031);
nor U2052 (N_2052,N_1847,N_1215);
nand U2053 (N_2053,N_1876,N_1618);
xor U2054 (N_2054,N_1837,N_1234);
xor U2055 (N_2055,N_1386,N_1782);
xor U2056 (N_2056,N_1063,N_1152);
and U2057 (N_2057,N_1278,N_1579);
xor U2058 (N_2058,N_1843,N_1216);
and U2059 (N_2059,N_1114,N_1407);
and U2060 (N_2060,N_1255,N_1285);
or U2061 (N_2061,N_1680,N_1017);
nand U2062 (N_2062,N_1360,N_1460);
nor U2063 (N_2063,N_1865,N_1930);
or U2064 (N_2064,N_1718,N_1363);
nand U2065 (N_2065,N_1261,N_1397);
or U2066 (N_2066,N_1300,N_1437);
or U2067 (N_2067,N_1128,N_1968);
and U2068 (N_2068,N_1826,N_1254);
or U2069 (N_2069,N_1056,N_1351);
nand U2070 (N_2070,N_1457,N_1761);
nand U2071 (N_2071,N_1540,N_1730);
nand U2072 (N_2072,N_1277,N_1859);
and U2073 (N_2073,N_1095,N_1797);
and U2074 (N_2074,N_1461,N_1167);
and U2075 (N_2075,N_1860,N_1990);
and U2076 (N_2076,N_1796,N_1101);
and U2077 (N_2077,N_1952,N_1549);
or U2078 (N_2078,N_1497,N_1170);
nor U2079 (N_2079,N_1404,N_1955);
nand U2080 (N_2080,N_1472,N_1755);
or U2081 (N_2081,N_1502,N_1270);
nand U2082 (N_2082,N_1456,N_1494);
xnor U2083 (N_2083,N_1318,N_1268);
nand U2084 (N_2084,N_1985,N_1102);
and U2085 (N_2085,N_1945,N_1288);
nor U2086 (N_2086,N_1282,N_1334);
or U2087 (N_2087,N_1193,N_1789);
nand U2088 (N_2088,N_1879,N_1200);
nor U2089 (N_2089,N_1511,N_1941);
nand U2090 (N_2090,N_1603,N_1724);
nor U2091 (N_2091,N_1516,N_1088);
xnor U2092 (N_2092,N_1813,N_1652);
nand U2093 (N_2093,N_1606,N_1116);
xor U2094 (N_2094,N_1640,N_1190);
and U2095 (N_2095,N_1742,N_1306);
and U2096 (N_2096,N_1575,N_1044);
or U2097 (N_2097,N_1195,N_1184);
nor U2098 (N_2098,N_1011,N_1552);
and U2099 (N_2099,N_1975,N_1223);
xnor U2100 (N_2100,N_1415,N_1512);
or U2101 (N_2101,N_1849,N_1621);
xor U2102 (N_2102,N_1368,N_1445);
nand U2103 (N_2103,N_1956,N_1733);
xor U2104 (N_2104,N_1885,N_1441);
or U2105 (N_2105,N_1286,N_1830);
nor U2106 (N_2106,N_1387,N_1355);
nor U2107 (N_2107,N_1417,N_1633);
or U2108 (N_2108,N_1086,N_1105);
and U2109 (N_2109,N_1882,N_1382);
or U2110 (N_2110,N_1523,N_1339);
xnor U2111 (N_2111,N_1644,N_1046);
or U2112 (N_2112,N_1887,N_1886);
or U2113 (N_2113,N_1779,N_1366);
and U2114 (N_2114,N_1219,N_1821);
nand U2115 (N_2115,N_1439,N_1615);
xnor U2116 (N_2116,N_1539,N_1126);
and U2117 (N_2117,N_1094,N_1522);
nand U2118 (N_2118,N_1921,N_1869);
nor U2119 (N_2119,N_1636,N_1375);
nand U2120 (N_2120,N_1935,N_1080);
or U2121 (N_2121,N_1914,N_1295);
nor U2122 (N_2122,N_1358,N_1474);
nor U2123 (N_2123,N_1263,N_1156);
nor U2124 (N_2124,N_1915,N_1484);
and U2125 (N_2125,N_1024,N_1290);
and U2126 (N_2126,N_1150,N_1060);
or U2127 (N_2127,N_1340,N_1663);
nor U2128 (N_2128,N_1369,N_1192);
or U2129 (N_2129,N_1049,N_1058);
nand U2130 (N_2130,N_1934,N_1344);
nand U2131 (N_2131,N_1580,N_1949);
nor U2132 (N_2132,N_1061,N_1289);
nor U2133 (N_2133,N_1159,N_1325);
or U2134 (N_2134,N_1891,N_1564);
and U2135 (N_2135,N_1671,N_1576);
nand U2136 (N_2136,N_1180,N_1875);
xnor U2137 (N_2137,N_1650,N_1877);
nor U2138 (N_2138,N_1670,N_1807);
nor U2139 (N_2139,N_1222,N_1809);
or U2140 (N_2140,N_1786,N_1047);
or U2141 (N_2141,N_1224,N_1316);
or U2142 (N_2142,N_1002,N_1710);
xnor U2143 (N_2143,N_1940,N_1019);
or U2144 (N_2144,N_1878,N_1588);
and U2145 (N_2145,N_1583,N_1297);
nand U2146 (N_2146,N_1706,N_1326);
nor U2147 (N_2147,N_1854,N_1722);
nor U2148 (N_2148,N_1605,N_1501);
and U2149 (N_2149,N_1816,N_1734);
nand U2150 (N_2150,N_1266,N_1701);
nor U2151 (N_2151,N_1685,N_1151);
nor U2152 (N_2152,N_1759,N_1719);
nor U2153 (N_2153,N_1335,N_1899);
nor U2154 (N_2154,N_1136,N_1957);
nor U2155 (N_2155,N_1550,N_1642);
xor U2156 (N_2156,N_1127,N_1463);
and U2157 (N_2157,N_1760,N_1695);
xor U2158 (N_2158,N_1364,N_1983);
and U2159 (N_2159,N_1515,N_1767);
and U2160 (N_2160,N_1021,N_1978);
xnor U2161 (N_2161,N_1469,N_1165);
nand U2162 (N_2162,N_1059,N_1555);
and U2163 (N_2163,N_1093,N_1487);
and U2164 (N_2164,N_1924,N_1121);
nor U2165 (N_2165,N_1634,N_1256);
nand U2166 (N_2166,N_1569,N_1824);
nand U2167 (N_2167,N_1856,N_1206);
nor U2168 (N_2168,N_1962,N_1571);
and U2169 (N_2169,N_1850,N_1681);
nor U2170 (N_2170,N_1905,N_1451);
or U2171 (N_2171,N_1545,N_1135);
xnor U2172 (N_2172,N_1752,N_1661);
nand U2173 (N_2173,N_1800,N_1444);
nand U2174 (N_2174,N_1691,N_1853);
nor U2175 (N_2175,N_1775,N_1053);
nand U2176 (N_2176,N_1327,N_1848);
nor U2177 (N_2177,N_1177,N_1209);
nor U2178 (N_2178,N_1932,N_1532);
nor U2179 (N_2179,N_1458,N_1374);
xnor U2180 (N_2180,N_1835,N_1519);
nor U2181 (N_2181,N_1995,N_1777);
nand U2182 (N_2182,N_1526,N_1008);
and U2183 (N_2183,N_1740,N_1713);
or U2184 (N_2184,N_1446,N_1284);
nand U2185 (N_2185,N_1303,N_1328);
or U2186 (N_2186,N_1513,N_1072);
nand U2187 (N_2187,N_1692,N_1089);
xnor U2188 (N_2188,N_1378,N_1475);
nor U2189 (N_2189,N_1980,N_1669);
and U2190 (N_2190,N_1243,N_1400);
nand U2191 (N_2191,N_1308,N_1525);
or U2192 (N_2192,N_1183,N_1735);
or U2193 (N_2193,N_1015,N_1542);
nor U2194 (N_2194,N_1736,N_1396);
and U2195 (N_2195,N_1863,N_1925);
nor U2196 (N_2196,N_1960,N_1953);
nand U2197 (N_2197,N_1174,N_1162);
and U2198 (N_2198,N_1204,N_1611);
and U2199 (N_2199,N_1070,N_1793);
and U2200 (N_2200,N_1749,N_1637);
nor U2201 (N_2201,N_1504,N_1666);
or U2202 (N_2202,N_1182,N_1645);
or U2203 (N_2203,N_1732,N_1874);
and U2204 (N_2204,N_1349,N_1408);
nand U2205 (N_2205,N_1918,N_1449);
and U2206 (N_2206,N_1076,N_1589);
or U2207 (N_2207,N_1563,N_1443);
nor U2208 (N_2208,N_1842,N_1125);
or U2209 (N_2209,N_1772,N_1132);
and U2210 (N_2210,N_1997,N_1210);
or U2211 (N_2211,N_1855,N_1269);
and U2212 (N_2212,N_1778,N_1614);
nand U2213 (N_2213,N_1188,N_1438);
nand U2214 (N_2214,N_1007,N_1572);
nor U2215 (N_2215,N_1534,N_1901);
or U2216 (N_2216,N_1373,N_1062);
nand U2217 (N_2217,N_1919,N_1794);
and U2218 (N_2218,N_1144,N_1252);
or U2219 (N_2219,N_1166,N_1766);
or U2220 (N_2220,N_1500,N_1221);
or U2221 (N_2221,N_1912,N_1683);
xor U2222 (N_2222,N_1176,N_1178);
nor U2223 (N_2223,N_1505,N_1381);
or U2224 (N_2224,N_1699,N_1479);
and U2225 (N_2225,N_1851,N_1483);
or U2226 (N_2226,N_1304,N_1689);
and U2227 (N_2227,N_1181,N_1187);
nor U2228 (N_2228,N_1802,N_1768);
and U2229 (N_2229,N_1998,N_1194);
nand U2230 (N_2230,N_1447,N_1149);
nand U2231 (N_2231,N_1541,N_1389);
or U2232 (N_2232,N_1048,N_1147);
nand U2233 (N_2233,N_1490,N_1091);
nor U2234 (N_2234,N_1130,N_1764);
or U2235 (N_2235,N_1016,N_1291);
nand U2236 (N_2236,N_1276,N_1867);
xnor U2237 (N_2237,N_1283,N_1037);
or U2238 (N_2238,N_1081,N_1141);
nor U2239 (N_2239,N_1967,N_1069);
or U2240 (N_2240,N_1774,N_1419);
nor U2241 (N_2241,N_1597,N_1586);
nand U2242 (N_2242,N_1330,N_1423);
nor U2243 (N_2243,N_1858,N_1004);
nand U2244 (N_2244,N_1888,N_1737);
nor U2245 (N_2245,N_1521,N_1414);
nor U2246 (N_2246,N_1529,N_1391);
nor U2247 (N_2247,N_1079,N_1894);
or U2248 (N_2248,N_1350,N_1903);
and U2249 (N_2249,N_1973,N_1909);
nor U2250 (N_2250,N_1343,N_1829);
nor U2251 (N_2251,N_1342,N_1320);
nand U2252 (N_2252,N_1942,N_1119);
nand U2253 (N_2253,N_1841,N_1982);
nor U2254 (N_2254,N_1230,N_1030);
nor U2255 (N_2255,N_1727,N_1551);
nor U2256 (N_2256,N_1298,N_1009);
and U2257 (N_2257,N_1705,N_1452);
nor U2258 (N_2258,N_1834,N_1025);
nor U2259 (N_2259,N_1811,N_1933);
nand U2260 (N_2260,N_1820,N_1347);
or U2261 (N_2261,N_1638,N_1591);
or U2262 (N_2262,N_1668,N_1976);
nand U2263 (N_2263,N_1574,N_1034);
and U2264 (N_2264,N_1473,N_1208);
or U2265 (N_2265,N_1106,N_1784);
nor U2266 (N_2266,N_1068,N_1662);
or U2267 (N_2267,N_1258,N_1074);
nor U2268 (N_2268,N_1197,N_1754);
nand U2269 (N_2269,N_1274,N_1570);
nor U2270 (N_2270,N_1338,N_1943);
nand U2271 (N_2271,N_1309,N_1623);
xor U2272 (N_2272,N_1674,N_1371);
nand U2273 (N_2273,N_1198,N_1169);
or U2274 (N_2274,N_1965,N_1299);
or U2275 (N_2275,N_1711,N_1138);
and U2276 (N_2276,N_1043,N_1087);
or U2277 (N_2277,N_1164,N_1155);
xor U2278 (N_2278,N_1410,N_1686);
nor U2279 (N_2279,N_1161,N_1476);
nor U2280 (N_2280,N_1280,N_1708);
or U2281 (N_2281,N_1085,N_1632);
nand U2282 (N_2282,N_1346,N_1936);
nand U2283 (N_2283,N_1014,N_1720);
and U2284 (N_2284,N_1993,N_1241);
xnor U2285 (N_2285,N_1600,N_1664);
and U2286 (N_2286,N_1917,N_1311);
and U2287 (N_2287,N_1773,N_1787);
or U2288 (N_2288,N_1665,N_1413);
and U2289 (N_2289,N_1045,N_1265);
nor U2290 (N_2290,N_1433,N_1498);
or U2291 (N_2291,N_1753,N_1050);
nor U2292 (N_2292,N_1154,N_1310);
nor U2293 (N_2293,N_1022,N_1981);
and U2294 (N_2294,N_1873,N_1026);
and U2295 (N_2295,N_1920,N_1424);
nand U2296 (N_2296,N_1431,N_1577);
nor U2297 (N_2297,N_1649,N_1465);
xnor U2298 (N_2298,N_1785,N_1312);
and U2299 (N_2299,N_1726,N_1229);
or U2300 (N_2300,N_1432,N_1157);
or U2301 (N_2301,N_1817,N_1040);
xor U2302 (N_2302,N_1913,N_1697);
xnor U2303 (N_2303,N_1616,N_1225);
nand U2304 (N_2304,N_1808,N_1840);
or U2305 (N_2305,N_1171,N_1247);
nor U2306 (N_2306,N_1884,N_1054);
or U2307 (N_2307,N_1321,N_1868);
nand U2308 (N_2308,N_1491,N_1987);
nor U2309 (N_2309,N_1510,N_1251);
and U2310 (N_2310,N_1527,N_1281);
xnor U2311 (N_2311,N_1622,N_1937);
and U2312 (N_2312,N_1051,N_1124);
and U2313 (N_2313,N_1972,N_1133);
or U2314 (N_2314,N_1994,N_1682);
or U2315 (N_2315,N_1827,N_1035);
xnor U2316 (N_2316,N_1911,N_1609);
nand U2317 (N_2317,N_1212,N_1238);
nor U2318 (N_2318,N_1693,N_1619);
and U2319 (N_2319,N_1450,N_1818);
nor U2320 (N_2320,N_1815,N_1464);
or U2321 (N_2321,N_1348,N_1839);
nor U2322 (N_2322,N_1420,N_1426);
nor U2323 (N_2323,N_1199,N_1771);
and U2324 (N_2324,N_1561,N_1958);
nor U2325 (N_2325,N_1769,N_1931);
xor U2326 (N_2326,N_1357,N_1567);
nor U2327 (N_2327,N_1393,N_1900);
and U2328 (N_2328,N_1890,N_1963);
nor U2329 (N_2329,N_1961,N_1333);
and U2330 (N_2330,N_1536,N_1977);
or U2331 (N_2331,N_1585,N_1250);
or U2332 (N_2332,N_1118,N_1573);
xor U2333 (N_2333,N_1639,N_1648);
or U2334 (N_2334,N_1036,N_1454);
and U2335 (N_2335,N_1499,N_1906);
nand U2336 (N_2336,N_1264,N_1989);
or U2337 (N_2337,N_1714,N_1646);
nor U2338 (N_2338,N_1746,N_1425);
nand U2339 (N_2339,N_1379,N_1356);
or U2340 (N_2340,N_1996,N_1684);
nand U2341 (N_2341,N_1898,N_1055);
and U2342 (N_2342,N_1459,N_1831);
xnor U2343 (N_2343,N_1202,N_1294);
or U2344 (N_2344,N_1213,N_1324);
or U2345 (N_2345,N_1677,N_1140);
and U2346 (N_2346,N_1845,N_1590);
or U2347 (N_2347,N_1717,N_1629);
nand U2348 (N_2348,N_1496,N_1148);
and U2349 (N_2349,N_1814,N_1275);
and U2350 (N_2350,N_1559,N_1592);
nor U2351 (N_2351,N_1272,N_1383);
and U2352 (N_2352,N_1380,N_1599);
or U2353 (N_2353,N_1795,N_1974);
and U2354 (N_2354,N_1598,N_1001);
or U2355 (N_2355,N_1568,N_1731);
or U2356 (N_2356,N_1077,N_1738);
or U2357 (N_2357,N_1478,N_1553);
nor U2358 (N_2358,N_1812,N_1010);
and U2359 (N_2359,N_1715,N_1548);
and U2360 (N_2360,N_1331,N_1883);
xnor U2361 (N_2361,N_1279,N_1608);
and U2362 (N_2362,N_1123,N_1704);
nand U2363 (N_2363,N_1792,N_1703);
nor U2364 (N_2364,N_1938,N_1314);
nor U2365 (N_2365,N_1493,N_1626);
and U2366 (N_2366,N_1728,N_1517);
and U2367 (N_2367,N_1406,N_1872);
and U2368 (N_2368,N_1405,N_1700);
or U2369 (N_2369,N_1078,N_1442);
nor U2370 (N_2370,N_1687,N_1897);
and U2371 (N_2371,N_1006,N_1104);
nor U2372 (N_2372,N_1688,N_1352);
and U2373 (N_2373,N_1508,N_1399);
nand U2374 (N_2374,N_1240,N_1833);
nor U2375 (N_2375,N_1110,N_1470);
nand U2376 (N_2376,N_1108,N_1332);
nor U2377 (N_2377,N_1145,N_1596);
nor U2378 (N_2378,N_1057,N_1153);
or U2379 (N_2379,N_1492,N_1852);
and U2380 (N_2380,N_1218,N_1232);
xor U2381 (N_2381,N_1528,N_1163);
nor U2382 (N_2382,N_1412,N_1485);
nor U2383 (N_2383,N_1065,N_1509);
nand U2384 (N_2384,N_1617,N_1075);
nand U2385 (N_2385,N_1870,N_1741);
and U2386 (N_2386,N_1096,N_1226);
nor U2387 (N_2387,N_1098,N_1262);
nor U2388 (N_2388,N_1107,N_1395);
xnor U2389 (N_2389,N_1971,N_1227);
or U2390 (N_2390,N_1783,N_1547);
or U2391 (N_2391,N_1203,N_1828);
or U2392 (N_2392,N_1090,N_1146);
or U2393 (N_2393,N_1578,N_1798);
or U2394 (N_2394,N_1750,N_1595);
or U2395 (N_2395,N_1709,N_1889);
nand U2396 (N_2396,N_1115,N_1013);
nand U2397 (N_2397,N_1673,N_1482);
nor U2398 (N_2398,N_1235,N_1970);
xor U2399 (N_2399,N_1370,N_1111);
nand U2400 (N_2400,N_1520,N_1214);
and U2401 (N_2401,N_1336,N_1744);
xor U2402 (N_2402,N_1904,N_1988);
or U2403 (N_2403,N_1803,N_1073);
nor U2404 (N_2404,N_1029,N_1293);
nor U2405 (N_2405,N_1185,N_1315);
and U2406 (N_2406,N_1984,N_1003);
nor U2407 (N_2407,N_1601,N_1537);
xnor U2408 (N_2408,N_1353,N_1033);
nand U2409 (N_2409,N_1158,N_1403);
and U2410 (N_2410,N_1846,N_1103);
and U2411 (N_2411,N_1558,N_1455);
nor U2412 (N_2412,N_1267,N_1630);
nor U2413 (N_2413,N_1430,N_1628);
nor U2414 (N_2414,N_1702,N_1120);
nand U2415 (N_2415,N_1672,N_1748);
and U2416 (N_2416,N_1388,N_1908);
xnor U2417 (N_2417,N_1005,N_1895);
nor U2418 (N_2418,N_1207,N_1319);
nand U2419 (N_2419,N_1142,N_1531);
nand U2420 (N_2420,N_1806,N_1296);
or U2421 (N_2421,N_1892,N_1756);
nand U2422 (N_2422,N_1620,N_1543);
nor U2423 (N_2423,N_1468,N_1907);
or U2424 (N_2424,N_1675,N_1367);
nand U2425 (N_2425,N_1012,N_1770);
or U2426 (N_2426,N_1518,N_1866);
xor U2427 (N_2427,N_1402,N_1307);
and U2428 (N_2428,N_1819,N_1948);
nor U2429 (N_2429,N_1657,N_1776);
or U2430 (N_2430,N_1966,N_1416);
nor U2431 (N_2431,N_1390,N_1844);
and U2432 (N_2432,N_1765,N_1762);
and U2433 (N_2433,N_1838,N_1467);
xor U2434 (N_2434,N_1880,N_1857);
and U2435 (N_2435,N_1302,N_1790);
xor U2436 (N_2436,N_1651,N_1959);
xor U2437 (N_2437,N_1613,N_1721);
or U2438 (N_2438,N_1698,N_1986);
or U2439 (N_2439,N_1643,N_1139);
nor U2440 (N_2440,N_1196,N_1557);
nor U2441 (N_2441,N_1538,N_1253);
and U2442 (N_2442,N_1862,N_1951);
and U2443 (N_2443,N_1694,N_1716);
and U2444 (N_2444,N_1260,N_1745);
xor U2445 (N_2445,N_1064,N_1678);
nand U2446 (N_2446,N_1896,N_1627);
and U2447 (N_2447,N_1398,N_1836);
nor U2448 (N_2448,N_1259,N_1271);
nand U2449 (N_2449,N_1641,N_1249);
or U2450 (N_2450,N_1409,N_1560);
and U2451 (N_2451,N_1788,N_1881);
or U2452 (N_2452,N_1376,N_1916);
and U2453 (N_2453,N_1992,N_1810);
nor U2454 (N_2454,N_1372,N_1902);
nor U2455 (N_2455,N_1359,N_1712);
xnor U2456 (N_2456,N_1301,N_1581);
nand U2457 (N_2457,N_1201,N_1137);
nor U2458 (N_2458,N_1625,N_1018);
nor U2459 (N_2459,N_1554,N_1067);
nand U2460 (N_2460,N_1584,N_1477);
and U2461 (N_2461,N_1097,N_1799);
and U2462 (N_2462,N_1428,N_1440);
nand U2463 (N_2463,N_1041,N_1660);
or U2464 (N_2464,N_1175,N_1612);
xnor U2465 (N_2465,N_1071,N_1143);
nor U2466 (N_2466,N_1117,N_1763);
nand U2467 (N_2467,N_1000,N_1893);
and U2468 (N_2468,N_1676,N_1113);
and U2469 (N_2469,N_1729,N_1871);
nor U2470 (N_2470,N_1435,N_1723);
or U2471 (N_2471,N_1743,N_1481);
and U2472 (N_2472,N_1659,N_1514);
or U2473 (N_2473,N_1462,N_1305);
nor U2474 (N_2474,N_1211,N_1486);
or U2475 (N_2475,N_1023,N_1191);
or U2476 (N_2476,N_1418,N_1066);
nor U2477 (N_2477,N_1655,N_1801);
or U2478 (N_2478,N_1434,N_1780);
nand U2479 (N_2479,N_1084,N_1923);
or U2480 (N_2480,N_1082,N_1377);
or U2481 (N_2481,N_1317,N_1361);
or U2482 (N_2482,N_1861,N_1566);
and U2483 (N_2483,N_1910,N_1530);
or U2484 (N_2484,N_1384,N_1587);
or U2485 (N_2485,N_1168,N_1654);
nand U2486 (N_2486,N_1427,N_1610);
and U2487 (N_2487,N_1565,N_1237);
and U2488 (N_2488,N_1453,N_1562);
or U2489 (N_2489,N_1503,N_1471);
nor U2490 (N_2490,N_1690,N_1781);
and U2491 (N_2491,N_1489,N_1392);
nand U2492 (N_2492,N_1480,N_1488);
nand U2493 (N_2493,N_1231,N_1337);
nand U2494 (N_2494,N_1926,N_1964);
or U2495 (N_2495,N_1172,N_1864);
and U2496 (N_2496,N_1027,N_1422);
and U2497 (N_2497,N_1273,N_1739);
nand U2498 (N_2498,N_1217,N_1287);
nor U2499 (N_2499,N_1134,N_1604);
nand U2500 (N_2500,N_1606,N_1933);
and U2501 (N_2501,N_1957,N_1821);
nand U2502 (N_2502,N_1716,N_1846);
or U2503 (N_2503,N_1253,N_1613);
and U2504 (N_2504,N_1065,N_1999);
and U2505 (N_2505,N_1756,N_1486);
and U2506 (N_2506,N_1748,N_1222);
and U2507 (N_2507,N_1192,N_1952);
nand U2508 (N_2508,N_1545,N_1228);
and U2509 (N_2509,N_1460,N_1892);
nor U2510 (N_2510,N_1190,N_1312);
or U2511 (N_2511,N_1296,N_1531);
or U2512 (N_2512,N_1481,N_1180);
nand U2513 (N_2513,N_1454,N_1326);
nand U2514 (N_2514,N_1877,N_1017);
nand U2515 (N_2515,N_1669,N_1663);
nor U2516 (N_2516,N_1677,N_1935);
xnor U2517 (N_2517,N_1892,N_1328);
and U2518 (N_2518,N_1676,N_1290);
xnor U2519 (N_2519,N_1302,N_1863);
nand U2520 (N_2520,N_1813,N_1074);
nor U2521 (N_2521,N_1792,N_1599);
nand U2522 (N_2522,N_1823,N_1468);
nor U2523 (N_2523,N_1703,N_1663);
and U2524 (N_2524,N_1260,N_1446);
and U2525 (N_2525,N_1164,N_1138);
nor U2526 (N_2526,N_1673,N_1519);
and U2527 (N_2527,N_1289,N_1330);
and U2528 (N_2528,N_1975,N_1263);
nor U2529 (N_2529,N_1235,N_1416);
and U2530 (N_2530,N_1907,N_1357);
and U2531 (N_2531,N_1794,N_1282);
and U2532 (N_2532,N_1192,N_1253);
and U2533 (N_2533,N_1231,N_1115);
nand U2534 (N_2534,N_1084,N_1277);
nor U2535 (N_2535,N_1616,N_1329);
and U2536 (N_2536,N_1033,N_1014);
nor U2537 (N_2537,N_1149,N_1474);
or U2538 (N_2538,N_1814,N_1315);
and U2539 (N_2539,N_1012,N_1815);
or U2540 (N_2540,N_1794,N_1782);
xor U2541 (N_2541,N_1699,N_1491);
and U2542 (N_2542,N_1466,N_1377);
and U2543 (N_2543,N_1892,N_1480);
nor U2544 (N_2544,N_1145,N_1954);
nand U2545 (N_2545,N_1564,N_1518);
or U2546 (N_2546,N_1752,N_1512);
and U2547 (N_2547,N_1256,N_1894);
and U2548 (N_2548,N_1802,N_1212);
nor U2549 (N_2549,N_1854,N_1293);
xnor U2550 (N_2550,N_1391,N_1461);
xnor U2551 (N_2551,N_1860,N_1312);
and U2552 (N_2552,N_1651,N_1522);
nand U2553 (N_2553,N_1879,N_1342);
xor U2554 (N_2554,N_1092,N_1195);
and U2555 (N_2555,N_1028,N_1306);
nand U2556 (N_2556,N_1201,N_1386);
xnor U2557 (N_2557,N_1347,N_1926);
nand U2558 (N_2558,N_1773,N_1025);
nor U2559 (N_2559,N_1448,N_1161);
or U2560 (N_2560,N_1721,N_1009);
nor U2561 (N_2561,N_1164,N_1810);
nor U2562 (N_2562,N_1110,N_1189);
and U2563 (N_2563,N_1360,N_1010);
nor U2564 (N_2564,N_1367,N_1059);
nor U2565 (N_2565,N_1289,N_1807);
nand U2566 (N_2566,N_1167,N_1868);
and U2567 (N_2567,N_1484,N_1739);
nand U2568 (N_2568,N_1582,N_1431);
xnor U2569 (N_2569,N_1186,N_1173);
or U2570 (N_2570,N_1624,N_1743);
or U2571 (N_2571,N_1490,N_1204);
nand U2572 (N_2572,N_1209,N_1565);
and U2573 (N_2573,N_1349,N_1841);
nor U2574 (N_2574,N_1953,N_1318);
or U2575 (N_2575,N_1708,N_1287);
nand U2576 (N_2576,N_1678,N_1128);
nor U2577 (N_2577,N_1253,N_1227);
and U2578 (N_2578,N_1111,N_1750);
or U2579 (N_2579,N_1956,N_1095);
or U2580 (N_2580,N_1677,N_1463);
and U2581 (N_2581,N_1818,N_1569);
nor U2582 (N_2582,N_1897,N_1929);
nand U2583 (N_2583,N_1251,N_1976);
and U2584 (N_2584,N_1513,N_1210);
and U2585 (N_2585,N_1546,N_1648);
xor U2586 (N_2586,N_1965,N_1016);
or U2587 (N_2587,N_1802,N_1039);
nand U2588 (N_2588,N_1531,N_1844);
and U2589 (N_2589,N_1966,N_1928);
nor U2590 (N_2590,N_1267,N_1858);
nand U2591 (N_2591,N_1117,N_1824);
nor U2592 (N_2592,N_1018,N_1293);
and U2593 (N_2593,N_1377,N_1306);
and U2594 (N_2594,N_1707,N_1332);
or U2595 (N_2595,N_1394,N_1487);
and U2596 (N_2596,N_1938,N_1552);
and U2597 (N_2597,N_1755,N_1860);
or U2598 (N_2598,N_1127,N_1103);
or U2599 (N_2599,N_1585,N_1889);
nor U2600 (N_2600,N_1842,N_1074);
nand U2601 (N_2601,N_1592,N_1631);
or U2602 (N_2602,N_1654,N_1836);
and U2603 (N_2603,N_1860,N_1390);
and U2604 (N_2604,N_1819,N_1125);
nand U2605 (N_2605,N_1399,N_1860);
nor U2606 (N_2606,N_1284,N_1747);
nand U2607 (N_2607,N_1465,N_1388);
nand U2608 (N_2608,N_1282,N_1469);
or U2609 (N_2609,N_1533,N_1213);
nor U2610 (N_2610,N_1197,N_1630);
and U2611 (N_2611,N_1669,N_1691);
or U2612 (N_2612,N_1414,N_1844);
nor U2613 (N_2613,N_1689,N_1422);
nand U2614 (N_2614,N_1729,N_1160);
and U2615 (N_2615,N_1545,N_1124);
nor U2616 (N_2616,N_1756,N_1666);
or U2617 (N_2617,N_1377,N_1187);
and U2618 (N_2618,N_1862,N_1726);
nor U2619 (N_2619,N_1318,N_1331);
and U2620 (N_2620,N_1990,N_1314);
nor U2621 (N_2621,N_1813,N_1173);
or U2622 (N_2622,N_1053,N_1460);
nand U2623 (N_2623,N_1892,N_1647);
and U2624 (N_2624,N_1708,N_1194);
and U2625 (N_2625,N_1092,N_1999);
nand U2626 (N_2626,N_1795,N_1807);
and U2627 (N_2627,N_1023,N_1960);
nor U2628 (N_2628,N_1844,N_1309);
or U2629 (N_2629,N_1490,N_1518);
and U2630 (N_2630,N_1092,N_1648);
or U2631 (N_2631,N_1202,N_1679);
nor U2632 (N_2632,N_1435,N_1247);
xor U2633 (N_2633,N_1777,N_1030);
and U2634 (N_2634,N_1218,N_1205);
or U2635 (N_2635,N_1515,N_1686);
nand U2636 (N_2636,N_1017,N_1367);
and U2637 (N_2637,N_1061,N_1158);
or U2638 (N_2638,N_1198,N_1377);
and U2639 (N_2639,N_1543,N_1182);
nor U2640 (N_2640,N_1470,N_1588);
and U2641 (N_2641,N_1807,N_1203);
nand U2642 (N_2642,N_1751,N_1977);
and U2643 (N_2643,N_1834,N_1307);
and U2644 (N_2644,N_1444,N_1676);
xnor U2645 (N_2645,N_1848,N_1902);
nand U2646 (N_2646,N_1960,N_1501);
nand U2647 (N_2647,N_1573,N_1934);
nor U2648 (N_2648,N_1901,N_1073);
or U2649 (N_2649,N_1290,N_1730);
nor U2650 (N_2650,N_1864,N_1578);
xor U2651 (N_2651,N_1458,N_1860);
nand U2652 (N_2652,N_1442,N_1106);
nor U2653 (N_2653,N_1795,N_1408);
nor U2654 (N_2654,N_1368,N_1825);
nor U2655 (N_2655,N_1632,N_1702);
or U2656 (N_2656,N_1472,N_1264);
or U2657 (N_2657,N_1943,N_1069);
and U2658 (N_2658,N_1839,N_1192);
or U2659 (N_2659,N_1261,N_1284);
and U2660 (N_2660,N_1073,N_1951);
and U2661 (N_2661,N_1227,N_1862);
nand U2662 (N_2662,N_1021,N_1154);
and U2663 (N_2663,N_1594,N_1821);
nor U2664 (N_2664,N_1244,N_1985);
or U2665 (N_2665,N_1169,N_1302);
or U2666 (N_2666,N_1975,N_1589);
nor U2667 (N_2667,N_1224,N_1082);
and U2668 (N_2668,N_1737,N_1759);
and U2669 (N_2669,N_1234,N_1058);
nand U2670 (N_2670,N_1354,N_1019);
and U2671 (N_2671,N_1342,N_1091);
xor U2672 (N_2672,N_1474,N_1586);
and U2673 (N_2673,N_1674,N_1953);
nand U2674 (N_2674,N_1687,N_1590);
xor U2675 (N_2675,N_1339,N_1610);
nor U2676 (N_2676,N_1408,N_1257);
and U2677 (N_2677,N_1229,N_1037);
nand U2678 (N_2678,N_1763,N_1356);
or U2679 (N_2679,N_1153,N_1545);
xor U2680 (N_2680,N_1083,N_1935);
nor U2681 (N_2681,N_1400,N_1584);
nand U2682 (N_2682,N_1894,N_1064);
or U2683 (N_2683,N_1199,N_1679);
or U2684 (N_2684,N_1042,N_1874);
xor U2685 (N_2685,N_1399,N_1668);
nand U2686 (N_2686,N_1170,N_1545);
nor U2687 (N_2687,N_1390,N_1157);
and U2688 (N_2688,N_1281,N_1560);
or U2689 (N_2689,N_1627,N_1299);
nand U2690 (N_2690,N_1002,N_1012);
and U2691 (N_2691,N_1755,N_1139);
and U2692 (N_2692,N_1308,N_1956);
or U2693 (N_2693,N_1361,N_1697);
or U2694 (N_2694,N_1595,N_1862);
nor U2695 (N_2695,N_1409,N_1613);
nand U2696 (N_2696,N_1517,N_1791);
nand U2697 (N_2697,N_1585,N_1155);
nor U2698 (N_2698,N_1618,N_1772);
xnor U2699 (N_2699,N_1662,N_1484);
xnor U2700 (N_2700,N_1658,N_1308);
nand U2701 (N_2701,N_1282,N_1326);
nor U2702 (N_2702,N_1472,N_1663);
or U2703 (N_2703,N_1395,N_1330);
nor U2704 (N_2704,N_1353,N_1373);
and U2705 (N_2705,N_1674,N_1476);
and U2706 (N_2706,N_1662,N_1316);
nor U2707 (N_2707,N_1714,N_1286);
nand U2708 (N_2708,N_1333,N_1425);
nand U2709 (N_2709,N_1999,N_1302);
and U2710 (N_2710,N_1006,N_1253);
and U2711 (N_2711,N_1571,N_1697);
and U2712 (N_2712,N_1548,N_1850);
or U2713 (N_2713,N_1042,N_1626);
and U2714 (N_2714,N_1966,N_1386);
xor U2715 (N_2715,N_1546,N_1880);
nand U2716 (N_2716,N_1541,N_1657);
nand U2717 (N_2717,N_1575,N_1019);
and U2718 (N_2718,N_1878,N_1578);
or U2719 (N_2719,N_1747,N_1749);
nand U2720 (N_2720,N_1884,N_1863);
and U2721 (N_2721,N_1093,N_1789);
nor U2722 (N_2722,N_1469,N_1001);
nand U2723 (N_2723,N_1553,N_1654);
and U2724 (N_2724,N_1475,N_1783);
or U2725 (N_2725,N_1824,N_1099);
nor U2726 (N_2726,N_1868,N_1292);
or U2727 (N_2727,N_1014,N_1103);
nand U2728 (N_2728,N_1491,N_1938);
nor U2729 (N_2729,N_1123,N_1996);
xnor U2730 (N_2730,N_1135,N_1747);
nor U2731 (N_2731,N_1016,N_1306);
or U2732 (N_2732,N_1549,N_1080);
nor U2733 (N_2733,N_1465,N_1592);
nand U2734 (N_2734,N_1836,N_1743);
nand U2735 (N_2735,N_1852,N_1921);
xnor U2736 (N_2736,N_1597,N_1432);
xnor U2737 (N_2737,N_1115,N_1976);
or U2738 (N_2738,N_1530,N_1421);
and U2739 (N_2739,N_1728,N_1874);
nand U2740 (N_2740,N_1297,N_1313);
nand U2741 (N_2741,N_1316,N_1186);
and U2742 (N_2742,N_1965,N_1591);
or U2743 (N_2743,N_1905,N_1662);
xnor U2744 (N_2744,N_1346,N_1853);
nand U2745 (N_2745,N_1360,N_1932);
nor U2746 (N_2746,N_1955,N_1673);
or U2747 (N_2747,N_1075,N_1080);
nor U2748 (N_2748,N_1297,N_1335);
and U2749 (N_2749,N_1785,N_1081);
or U2750 (N_2750,N_1556,N_1771);
nor U2751 (N_2751,N_1378,N_1958);
nand U2752 (N_2752,N_1466,N_1162);
xor U2753 (N_2753,N_1789,N_1986);
or U2754 (N_2754,N_1650,N_1264);
xor U2755 (N_2755,N_1215,N_1095);
or U2756 (N_2756,N_1296,N_1566);
nor U2757 (N_2757,N_1110,N_1859);
nor U2758 (N_2758,N_1179,N_1533);
nand U2759 (N_2759,N_1901,N_1581);
and U2760 (N_2760,N_1848,N_1693);
nor U2761 (N_2761,N_1905,N_1856);
and U2762 (N_2762,N_1947,N_1898);
and U2763 (N_2763,N_1562,N_1194);
nor U2764 (N_2764,N_1768,N_1436);
xor U2765 (N_2765,N_1553,N_1545);
or U2766 (N_2766,N_1617,N_1215);
nor U2767 (N_2767,N_1104,N_1018);
nor U2768 (N_2768,N_1094,N_1569);
nand U2769 (N_2769,N_1182,N_1239);
nor U2770 (N_2770,N_1918,N_1445);
nand U2771 (N_2771,N_1318,N_1590);
and U2772 (N_2772,N_1248,N_1278);
nor U2773 (N_2773,N_1588,N_1144);
nor U2774 (N_2774,N_1298,N_1969);
nand U2775 (N_2775,N_1992,N_1056);
nand U2776 (N_2776,N_1081,N_1075);
nand U2777 (N_2777,N_1236,N_1511);
nor U2778 (N_2778,N_1146,N_1166);
nand U2779 (N_2779,N_1377,N_1790);
xnor U2780 (N_2780,N_1677,N_1711);
or U2781 (N_2781,N_1904,N_1869);
nor U2782 (N_2782,N_1543,N_1281);
nand U2783 (N_2783,N_1015,N_1932);
nand U2784 (N_2784,N_1371,N_1868);
or U2785 (N_2785,N_1046,N_1761);
nand U2786 (N_2786,N_1846,N_1848);
nand U2787 (N_2787,N_1756,N_1340);
nor U2788 (N_2788,N_1578,N_1292);
and U2789 (N_2789,N_1969,N_1900);
nand U2790 (N_2790,N_1839,N_1366);
nand U2791 (N_2791,N_1709,N_1140);
nand U2792 (N_2792,N_1027,N_1721);
and U2793 (N_2793,N_1780,N_1636);
and U2794 (N_2794,N_1442,N_1474);
or U2795 (N_2795,N_1567,N_1756);
nor U2796 (N_2796,N_1413,N_1180);
and U2797 (N_2797,N_1994,N_1661);
or U2798 (N_2798,N_1645,N_1270);
or U2799 (N_2799,N_1463,N_1036);
nand U2800 (N_2800,N_1931,N_1038);
nor U2801 (N_2801,N_1273,N_1872);
and U2802 (N_2802,N_1327,N_1102);
nor U2803 (N_2803,N_1224,N_1775);
or U2804 (N_2804,N_1299,N_1804);
or U2805 (N_2805,N_1229,N_1556);
nor U2806 (N_2806,N_1411,N_1331);
xor U2807 (N_2807,N_1297,N_1507);
or U2808 (N_2808,N_1167,N_1853);
nand U2809 (N_2809,N_1188,N_1572);
nor U2810 (N_2810,N_1629,N_1565);
and U2811 (N_2811,N_1360,N_1762);
and U2812 (N_2812,N_1517,N_1257);
or U2813 (N_2813,N_1443,N_1060);
nand U2814 (N_2814,N_1101,N_1877);
nand U2815 (N_2815,N_1059,N_1535);
or U2816 (N_2816,N_1692,N_1332);
or U2817 (N_2817,N_1401,N_1635);
nor U2818 (N_2818,N_1398,N_1696);
nand U2819 (N_2819,N_1400,N_1879);
nand U2820 (N_2820,N_1694,N_1709);
nor U2821 (N_2821,N_1165,N_1744);
and U2822 (N_2822,N_1001,N_1031);
nor U2823 (N_2823,N_1202,N_1920);
or U2824 (N_2824,N_1750,N_1669);
nor U2825 (N_2825,N_1358,N_1415);
nor U2826 (N_2826,N_1957,N_1387);
nor U2827 (N_2827,N_1805,N_1331);
nand U2828 (N_2828,N_1387,N_1207);
and U2829 (N_2829,N_1801,N_1735);
and U2830 (N_2830,N_1774,N_1906);
nor U2831 (N_2831,N_1708,N_1113);
nand U2832 (N_2832,N_1137,N_1030);
nor U2833 (N_2833,N_1608,N_1986);
xor U2834 (N_2834,N_1221,N_1450);
nor U2835 (N_2835,N_1449,N_1737);
or U2836 (N_2836,N_1076,N_1851);
or U2837 (N_2837,N_1031,N_1500);
or U2838 (N_2838,N_1748,N_1816);
nand U2839 (N_2839,N_1767,N_1189);
and U2840 (N_2840,N_1971,N_1339);
nor U2841 (N_2841,N_1504,N_1170);
nor U2842 (N_2842,N_1577,N_1320);
or U2843 (N_2843,N_1016,N_1862);
nor U2844 (N_2844,N_1935,N_1914);
and U2845 (N_2845,N_1018,N_1037);
xor U2846 (N_2846,N_1562,N_1110);
or U2847 (N_2847,N_1472,N_1178);
and U2848 (N_2848,N_1236,N_1515);
and U2849 (N_2849,N_1241,N_1818);
and U2850 (N_2850,N_1863,N_1202);
nor U2851 (N_2851,N_1662,N_1774);
nor U2852 (N_2852,N_1823,N_1151);
xor U2853 (N_2853,N_1061,N_1202);
nor U2854 (N_2854,N_1810,N_1905);
or U2855 (N_2855,N_1253,N_1784);
xor U2856 (N_2856,N_1374,N_1159);
nand U2857 (N_2857,N_1608,N_1521);
or U2858 (N_2858,N_1468,N_1040);
nand U2859 (N_2859,N_1995,N_1248);
nor U2860 (N_2860,N_1416,N_1751);
and U2861 (N_2861,N_1908,N_1881);
nor U2862 (N_2862,N_1397,N_1103);
nand U2863 (N_2863,N_1105,N_1264);
nor U2864 (N_2864,N_1989,N_1834);
and U2865 (N_2865,N_1522,N_1108);
or U2866 (N_2866,N_1821,N_1893);
or U2867 (N_2867,N_1093,N_1715);
or U2868 (N_2868,N_1186,N_1065);
xnor U2869 (N_2869,N_1500,N_1590);
or U2870 (N_2870,N_1846,N_1365);
nand U2871 (N_2871,N_1659,N_1328);
and U2872 (N_2872,N_1958,N_1369);
nand U2873 (N_2873,N_1023,N_1899);
nand U2874 (N_2874,N_1172,N_1973);
and U2875 (N_2875,N_1101,N_1572);
nand U2876 (N_2876,N_1727,N_1642);
xnor U2877 (N_2877,N_1734,N_1471);
nand U2878 (N_2878,N_1415,N_1759);
xnor U2879 (N_2879,N_1552,N_1929);
nor U2880 (N_2880,N_1524,N_1531);
nand U2881 (N_2881,N_1824,N_1747);
or U2882 (N_2882,N_1407,N_1901);
nand U2883 (N_2883,N_1362,N_1663);
nand U2884 (N_2884,N_1848,N_1027);
or U2885 (N_2885,N_1391,N_1641);
nand U2886 (N_2886,N_1813,N_1759);
nor U2887 (N_2887,N_1339,N_1330);
and U2888 (N_2888,N_1968,N_1817);
or U2889 (N_2889,N_1870,N_1233);
nor U2890 (N_2890,N_1308,N_1269);
and U2891 (N_2891,N_1517,N_1369);
nor U2892 (N_2892,N_1707,N_1305);
xnor U2893 (N_2893,N_1466,N_1424);
nor U2894 (N_2894,N_1018,N_1238);
nand U2895 (N_2895,N_1512,N_1326);
and U2896 (N_2896,N_1124,N_1530);
or U2897 (N_2897,N_1035,N_1112);
or U2898 (N_2898,N_1688,N_1116);
nand U2899 (N_2899,N_1874,N_1779);
xnor U2900 (N_2900,N_1220,N_1610);
nor U2901 (N_2901,N_1535,N_1685);
or U2902 (N_2902,N_1600,N_1082);
or U2903 (N_2903,N_1198,N_1284);
or U2904 (N_2904,N_1877,N_1630);
nand U2905 (N_2905,N_1782,N_1437);
and U2906 (N_2906,N_1816,N_1574);
or U2907 (N_2907,N_1483,N_1431);
nor U2908 (N_2908,N_1153,N_1026);
and U2909 (N_2909,N_1525,N_1084);
xnor U2910 (N_2910,N_1703,N_1604);
nor U2911 (N_2911,N_1259,N_1964);
nor U2912 (N_2912,N_1679,N_1713);
xnor U2913 (N_2913,N_1965,N_1613);
nor U2914 (N_2914,N_1799,N_1410);
and U2915 (N_2915,N_1285,N_1322);
nand U2916 (N_2916,N_1520,N_1390);
nand U2917 (N_2917,N_1691,N_1164);
nor U2918 (N_2918,N_1470,N_1181);
and U2919 (N_2919,N_1058,N_1797);
and U2920 (N_2920,N_1009,N_1735);
nand U2921 (N_2921,N_1769,N_1274);
or U2922 (N_2922,N_1552,N_1547);
and U2923 (N_2923,N_1855,N_1443);
and U2924 (N_2924,N_1368,N_1191);
or U2925 (N_2925,N_1593,N_1698);
nor U2926 (N_2926,N_1378,N_1761);
nand U2927 (N_2927,N_1279,N_1486);
and U2928 (N_2928,N_1928,N_1603);
and U2929 (N_2929,N_1478,N_1464);
nand U2930 (N_2930,N_1185,N_1856);
nand U2931 (N_2931,N_1919,N_1801);
nand U2932 (N_2932,N_1243,N_1778);
and U2933 (N_2933,N_1900,N_1327);
or U2934 (N_2934,N_1789,N_1240);
nand U2935 (N_2935,N_1803,N_1996);
nor U2936 (N_2936,N_1571,N_1626);
nor U2937 (N_2937,N_1750,N_1934);
and U2938 (N_2938,N_1213,N_1689);
nor U2939 (N_2939,N_1051,N_1771);
nor U2940 (N_2940,N_1018,N_1265);
nor U2941 (N_2941,N_1699,N_1235);
or U2942 (N_2942,N_1000,N_1973);
nor U2943 (N_2943,N_1859,N_1824);
nand U2944 (N_2944,N_1749,N_1211);
nor U2945 (N_2945,N_1346,N_1171);
or U2946 (N_2946,N_1363,N_1980);
xnor U2947 (N_2947,N_1231,N_1091);
or U2948 (N_2948,N_1668,N_1375);
nor U2949 (N_2949,N_1797,N_1325);
and U2950 (N_2950,N_1727,N_1878);
xnor U2951 (N_2951,N_1868,N_1298);
nand U2952 (N_2952,N_1913,N_1001);
or U2953 (N_2953,N_1387,N_1810);
nor U2954 (N_2954,N_1586,N_1845);
nor U2955 (N_2955,N_1248,N_1270);
nor U2956 (N_2956,N_1647,N_1673);
nand U2957 (N_2957,N_1489,N_1074);
nor U2958 (N_2958,N_1052,N_1950);
xnor U2959 (N_2959,N_1895,N_1337);
nor U2960 (N_2960,N_1216,N_1165);
or U2961 (N_2961,N_1528,N_1278);
xnor U2962 (N_2962,N_1288,N_1792);
or U2963 (N_2963,N_1344,N_1996);
nor U2964 (N_2964,N_1085,N_1049);
xor U2965 (N_2965,N_1053,N_1817);
or U2966 (N_2966,N_1314,N_1100);
nand U2967 (N_2967,N_1482,N_1117);
and U2968 (N_2968,N_1264,N_1564);
nand U2969 (N_2969,N_1685,N_1442);
nor U2970 (N_2970,N_1995,N_1853);
nor U2971 (N_2971,N_1607,N_1528);
or U2972 (N_2972,N_1264,N_1864);
and U2973 (N_2973,N_1750,N_1488);
nand U2974 (N_2974,N_1093,N_1187);
or U2975 (N_2975,N_1261,N_1953);
or U2976 (N_2976,N_1694,N_1662);
nand U2977 (N_2977,N_1337,N_1013);
or U2978 (N_2978,N_1430,N_1653);
xor U2979 (N_2979,N_1440,N_1478);
xnor U2980 (N_2980,N_1782,N_1340);
nand U2981 (N_2981,N_1424,N_1066);
nor U2982 (N_2982,N_1744,N_1495);
and U2983 (N_2983,N_1946,N_1633);
nand U2984 (N_2984,N_1485,N_1683);
nor U2985 (N_2985,N_1700,N_1027);
and U2986 (N_2986,N_1991,N_1853);
or U2987 (N_2987,N_1341,N_1338);
nand U2988 (N_2988,N_1018,N_1611);
nand U2989 (N_2989,N_1666,N_1846);
nor U2990 (N_2990,N_1547,N_1752);
nand U2991 (N_2991,N_1531,N_1922);
nand U2992 (N_2992,N_1707,N_1588);
or U2993 (N_2993,N_1739,N_1745);
nor U2994 (N_2994,N_1747,N_1143);
or U2995 (N_2995,N_1142,N_1040);
nor U2996 (N_2996,N_1957,N_1050);
and U2997 (N_2997,N_1412,N_1874);
and U2998 (N_2998,N_1413,N_1124);
nand U2999 (N_2999,N_1386,N_1647);
nand UO_0 (O_0,N_2840,N_2029);
or UO_1 (O_1,N_2101,N_2978);
and UO_2 (O_2,N_2828,N_2086);
and UO_3 (O_3,N_2410,N_2125);
nand UO_4 (O_4,N_2194,N_2306);
nand UO_5 (O_5,N_2476,N_2129);
xor UO_6 (O_6,N_2654,N_2708);
nor UO_7 (O_7,N_2287,N_2366);
and UO_8 (O_8,N_2383,N_2648);
nand UO_9 (O_9,N_2594,N_2509);
xnor UO_10 (O_10,N_2701,N_2007);
nand UO_11 (O_11,N_2760,N_2847);
nand UO_12 (O_12,N_2770,N_2661);
nand UO_13 (O_13,N_2347,N_2564);
nand UO_14 (O_14,N_2791,N_2051);
nor UO_15 (O_15,N_2527,N_2518);
and UO_16 (O_16,N_2923,N_2266);
or UO_17 (O_17,N_2519,N_2486);
or UO_18 (O_18,N_2653,N_2581);
and UO_19 (O_19,N_2852,N_2424);
nor UO_20 (O_20,N_2352,N_2888);
nand UO_21 (O_21,N_2827,N_2530);
xor UO_22 (O_22,N_2612,N_2599);
nor UO_23 (O_23,N_2872,N_2679);
nand UO_24 (O_24,N_2765,N_2388);
nand UO_25 (O_25,N_2319,N_2451);
nand UO_26 (O_26,N_2664,N_2467);
and UO_27 (O_27,N_2878,N_2951);
nor UO_28 (O_28,N_2326,N_2589);
or UO_29 (O_29,N_2365,N_2456);
nor UO_30 (O_30,N_2292,N_2091);
or UO_31 (O_31,N_2503,N_2056);
and UO_32 (O_32,N_2914,N_2290);
nor UO_33 (O_33,N_2850,N_2845);
and UO_34 (O_34,N_2475,N_2186);
or UO_35 (O_35,N_2110,N_2587);
or UO_36 (O_36,N_2882,N_2187);
xnor UO_37 (O_37,N_2991,N_2277);
nand UO_38 (O_38,N_2686,N_2657);
nor UO_39 (O_39,N_2211,N_2085);
and UO_40 (O_40,N_2099,N_2736);
and UO_41 (O_41,N_2331,N_2485);
or UO_42 (O_42,N_2321,N_2283);
xor UO_43 (O_43,N_2514,N_2919);
xor UO_44 (O_44,N_2180,N_2055);
nand UO_45 (O_45,N_2258,N_2360);
or UO_46 (O_46,N_2675,N_2504);
and UO_47 (O_47,N_2119,N_2027);
and UO_48 (O_48,N_2846,N_2245);
or UO_49 (O_49,N_2979,N_2320);
nand UO_50 (O_50,N_2309,N_2651);
and UO_51 (O_51,N_2553,N_2566);
or UO_52 (O_52,N_2896,N_2870);
nor UO_53 (O_53,N_2899,N_2992);
or UO_54 (O_54,N_2148,N_2133);
nand UO_55 (O_55,N_2555,N_2502);
and UO_56 (O_56,N_2719,N_2976);
or UO_57 (O_57,N_2733,N_2989);
or UO_58 (O_58,N_2229,N_2384);
nor UO_59 (O_59,N_2756,N_2173);
nor UO_60 (O_60,N_2794,N_2439);
and UO_61 (O_61,N_2833,N_2655);
or UO_62 (O_62,N_2047,N_2274);
and UO_63 (O_63,N_2449,N_2551);
or UO_64 (O_64,N_2997,N_2821);
and UO_65 (O_65,N_2251,N_2677);
nand UO_66 (O_66,N_2061,N_2597);
and UO_67 (O_67,N_2787,N_2582);
and UO_68 (O_68,N_2220,N_2069);
and UO_69 (O_69,N_2167,N_2005);
and UO_70 (O_70,N_2205,N_2407);
nor UO_71 (O_71,N_2049,N_2912);
or UO_72 (O_72,N_2834,N_2721);
nand UO_73 (O_73,N_2592,N_2171);
or UO_74 (O_74,N_2925,N_2644);
nor UO_75 (O_75,N_2779,N_2482);
and UO_76 (O_76,N_2747,N_2958);
nor UO_77 (O_77,N_2906,N_2818);
nor UO_78 (O_78,N_2716,N_2073);
and UO_79 (O_79,N_2829,N_2843);
and UO_80 (O_80,N_2610,N_2370);
or UO_81 (O_81,N_2307,N_2971);
nor UO_82 (O_82,N_2869,N_2798);
nor UO_83 (O_83,N_2092,N_2973);
nor UO_84 (O_84,N_2448,N_2304);
and UO_85 (O_85,N_2533,N_2017);
nor UO_86 (O_86,N_2100,N_2473);
nor UO_87 (O_87,N_2134,N_2639);
nor UO_88 (O_88,N_2190,N_2605);
or UO_89 (O_89,N_2534,N_2087);
nand UO_90 (O_90,N_2621,N_2106);
nand UO_91 (O_91,N_2506,N_2334);
nand UO_92 (O_92,N_2253,N_2928);
xor UO_93 (O_93,N_2004,N_2738);
and UO_94 (O_94,N_2408,N_2294);
and UO_95 (O_95,N_2768,N_2668);
or UO_96 (O_96,N_2762,N_2404);
nor UO_97 (O_97,N_2315,N_2214);
or UO_98 (O_98,N_2436,N_2557);
and UO_99 (O_99,N_2584,N_2030);
or UO_100 (O_100,N_2426,N_2987);
and UO_101 (O_101,N_2702,N_2993);
or UO_102 (O_102,N_2396,N_2411);
or UO_103 (O_103,N_2662,N_2616);
nand UO_104 (O_104,N_2392,N_2132);
nand UO_105 (O_105,N_2837,N_2666);
nor UO_106 (O_106,N_2217,N_2570);
and UO_107 (O_107,N_2959,N_2545);
and UO_108 (O_108,N_2728,N_2720);
nor UO_109 (O_109,N_2505,N_2603);
xor UO_110 (O_110,N_2921,N_2308);
and UO_111 (O_111,N_2002,N_2062);
xnor UO_112 (O_112,N_2703,N_2905);
nor UO_113 (O_113,N_2795,N_2851);
and UO_114 (O_114,N_2036,N_2957);
or UO_115 (O_115,N_2683,N_2685);
or UO_116 (O_116,N_2389,N_2942);
or UO_117 (O_117,N_2113,N_2913);
or UO_118 (O_118,N_2001,N_2147);
and UO_119 (O_119,N_2611,N_2885);
or UO_120 (O_120,N_2579,N_2780);
nand UO_121 (O_121,N_2151,N_2907);
nor UO_122 (O_122,N_2363,N_2465);
nor UO_123 (O_123,N_2994,N_2397);
or UO_124 (O_124,N_2523,N_2715);
or UO_125 (O_125,N_2037,N_2096);
nand UO_126 (O_126,N_2706,N_2182);
nand UO_127 (O_127,N_2313,N_2983);
and UO_128 (O_128,N_2831,N_2452);
nor UO_129 (O_129,N_2781,N_2725);
or UO_130 (O_130,N_2117,N_2267);
xnor UO_131 (O_131,N_2749,N_2016);
and UO_132 (O_132,N_2230,N_2572);
or UO_133 (O_133,N_2883,N_2803);
nor UO_134 (O_134,N_2927,N_2481);
or UO_135 (O_135,N_2947,N_2961);
xnor UO_136 (O_136,N_2717,N_2350);
and UO_137 (O_137,N_2429,N_2077);
nand UO_138 (O_138,N_2734,N_2197);
nor UO_139 (O_139,N_2676,N_2494);
nand UO_140 (O_140,N_2246,N_2152);
nand UO_141 (O_141,N_2338,N_2866);
and UO_142 (O_142,N_2932,N_2632);
and UO_143 (O_143,N_2689,N_2364);
nor UO_144 (O_144,N_2713,N_2568);
nand UO_145 (O_145,N_2788,N_2757);
and UO_146 (O_146,N_2012,N_2554);
nand UO_147 (O_147,N_2335,N_2876);
nor UO_148 (O_148,N_2945,N_2224);
nand UO_149 (O_149,N_2743,N_2415);
nand UO_150 (O_150,N_2826,N_2346);
xor UO_151 (O_151,N_2937,N_2751);
nor UO_152 (O_152,N_2140,N_2446);
or UO_153 (O_153,N_2636,N_2412);
xor UO_154 (O_154,N_2512,N_2430);
or UO_155 (O_155,N_2115,N_2952);
nor UO_156 (O_156,N_2969,N_2295);
nand UO_157 (O_157,N_2875,N_2520);
and UO_158 (O_158,N_2238,N_2684);
nor UO_159 (O_159,N_2272,N_2312);
or UO_160 (O_160,N_2785,N_2416);
and UO_161 (O_161,N_2059,N_2041);
nor UO_162 (O_162,N_2874,N_2460);
and UO_163 (O_163,N_2348,N_2967);
nand UO_164 (O_164,N_2130,N_2019);
nor UO_165 (O_165,N_2394,N_2243);
or UO_166 (O_166,N_2578,N_2832);
xor UO_167 (O_167,N_2081,N_2746);
or UO_168 (O_168,N_2709,N_2879);
xnor UO_169 (O_169,N_2844,N_2417);
or UO_170 (O_170,N_2790,N_2641);
or UO_171 (O_171,N_2585,N_2042);
nand UO_172 (O_172,N_2468,N_2435);
or UO_173 (O_173,N_2470,N_2647);
and UO_174 (O_174,N_2811,N_2381);
and UO_175 (O_175,N_2445,N_2303);
nor UO_176 (O_176,N_2006,N_2195);
xnor UO_177 (O_177,N_2786,N_2842);
nand UO_178 (O_178,N_2362,N_2332);
nor UO_179 (O_179,N_2420,N_2172);
nor UO_180 (O_180,N_2228,N_2154);
and UO_181 (O_181,N_2998,N_2783);
and UO_182 (O_182,N_2903,N_2282);
and UO_183 (O_183,N_2910,N_2109);
nand UO_184 (O_184,N_2139,N_2240);
and UO_185 (O_185,N_2218,N_2595);
and UO_186 (O_186,N_2179,N_2204);
nand UO_187 (O_187,N_2529,N_2457);
and UO_188 (O_188,N_2672,N_2718);
and UO_189 (O_189,N_2089,N_2082);
or UO_190 (O_190,N_2400,N_2206);
xnor UO_191 (O_191,N_2618,N_2965);
nand UO_192 (O_192,N_2271,N_2886);
nor UO_193 (O_193,N_2273,N_2090);
or UO_194 (O_194,N_2447,N_2895);
nor UO_195 (O_195,N_2543,N_2023);
and UO_196 (O_196,N_2576,N_2963);
nor UO_197 (O_197,N_2337,N_2669);
nand UO_198 (O_198,N_2469,N_2276);
and UO_199 (O_199,N_2136,N_2462);
or UO_200 (O_200,N_2966,N_2854);
xnor UO_201 (O_201,N_2804,N_2120);
or UO_202 (O_202,N_2615,N_2072);
nor UO_203 (O_203,N_2614,N_2990);
or UO_204 (O_204,N_2065,N_2114);
nor UO_205 (O_205,N_2285,N_2466);
or UO_206 (O_206,N_2499,N_2269);
and UO_207 (O_207,N_2155,N_2962);
nor UO_208 (O_208,N_2975,N_2542);
nand UO_209 (O_209,N_2691,N_2488);
and UO_210 (O_210,N_2627,N_2707);
xnor UO_211 (O_211,N_2898,N_2053);
or UO_212 (O_212,N_2112,N_2191);
and UO_213 (O_213,N_2633,N_2095);
and UO_214 (O_214,N_2122,N_2442);
or UO_215 (O_215,N_2735,N_2193);
or UO_216 (O_216,N_2613,N_2261);
nor UO_217 (O_217,N_2111,N_2617);
nand UO_218 (O_218,N_2043,N_2038);
or UO_219 (O_219,N_2311,N_2225);
nand UO_220 (O_220,N_2200,N_2208);
and UO_221 (O_221,N_2789,N_2301);
nor UO_222 (O_222,N_2263,N_2353);
and UO_223 (O_223,N_2729,N_2014);
nor UO_224 (O_224,N_2860,N_2935);
and UO_225 (O_225,N_2142,N_2897);
and UO_226 (O_226,N_2950,N_2265);
or UO_227 (O_227,N_2700,N_2593);
xor UO_228 (O_228,N_2867,N_2284);
nand UO_229 (O_229,N_2464,N_2825);
nor UO_230 (O_230,N_2813,N_2423);
nand UO_231 (O_231,N_2637,N_2547);
nor UO_232 (O_232,N_2541,N_2894);
or UO_233 (O_233,N_2591,N_2936);
or UO_234 (O_234,N_2540,N_2819);
nor UO_235 (O_235,N_2538,N_2583);
or UO_236 (O_236,N_2500,N_2257);
nand UO_237 (O_237,N_2419,N_2450);
or UO_238 (O_238,N_2046,N_2810);
nand UO_239 (O_239,N_2045,N_2640);
or UO_240 (O_240,N_2628,N_2558);
nor UO_241 (O_241,N_2658,N_2076);
and UO_242 (O_242,N_2836,N_2344);
and UO_243 (O_243,N_2477,N_2774);
nand UO_244 (O_244,N_2358,N_2562);
or UO_245 (O_245,N_2431,N_2455);
nand UO_246 (O_246,N_2807,N_2674);
nor UO_247 (O_247,N_2242,N_2501);
or UO_248 (O_248,N_2255,N_2724);
nand UO_249 (O_249,N_2682,N_2093);
nor UO_250 (O_250,N_2699,N_2079);
xor UO_251 (O_251,N_2608,N_2490);
nand UO_252 (O_252,N_2646,N_2176);
and UO_253 (O_253,N_2175,N_2623);
xnor UO_254 (O_254,N_2580,N_2345);
nand UO_255 (O_255,N_2479,N_2239);
and UO_256 (O_256,N_2213,N_2880);
and UO_257 (O_257,N_2607,N_2008);
or UO_258 (O_258,N_2575,N_2696);
and UO_259 (O_259,N_2857,N_2153);
nand UO_260 (O_260,N_2946,N_2234);
nand UO_261 (O_261,N_2454,N_2126);
or UO_262 (O_262,N_2569,N_2472);
or UO_263 (O_263,N_2236,N_2066);
and UO_264 (O_264,N_2216,N_2740);
xnor UO_265 (O_265,N_2385,N_2552);
and UO_266 (O_266,N_2441,N_2609);
and UO_267 (O_267,N_2517,N_2356);
and UO_268 (O_268,N_2972,N_2567);
or UO_269 (O_269,N_2943,N_2643);
nand UO_270 (O_270,N_2281,N_2944);
and UO_271 (O_271,N_2414,N_2771);
nor UO_272 (O_272,N_2799,N_2088);
nand UO_273 (O_273,N_2496,N_2980);
nor UO_274 (O_274,N_2219,N_2968);
nor UO_275 (O_275,N_2302,N_2138);
nor UO_276 (O_276,N_2393,N_2704);
xnor UO_277 (O_277,N_2891,N_2964);
and UO_278 (O_278,N_2022,N_2590);
xnor UO_279 (O_279,N_2052,N_2838);
xnor UO_280 (O_280,N_2098,N_2550);
nor UO_281 (O_281,N_2080,N_2177);
or UO_282 (O_282,N_2560,N_2020);
nand UO_283 (O_283,N_2291,N_2814);
nand UO_284 (O_284,N_2600,N_2588);
and UO_285 (O_285,N_2071,N_2940);
or UO_286 (O_286,N_2050,N_2954);
or UO_287 (O_287,N_2250,N_2687);
or UO_288 (O_288,N_2830,N_2443);
nand UO_289 (O_289,N_2268,N_2889);
nor UO_290 (O_290,N_2298,N_2726);
or UO_291 (O_291,N_2296,N_2275);
nand UO_292 (O_292,N_2861,N_2596);
nand UO_293 (O_293,N_2625,N_2920);
nand UO_294 (O_294,N_2556,N_2714);
or UO_295 (O_295,N_2432,N_2440);
and UO_296 (O_296,N_2824,N_2528);
nor UO_297 (O_297,N_2395,N_2336);
xor UO_298 (O_298,N_2808,N_2698);
and UO_299 (O_299,N_2561,N_2372);
nor UO_300 (O_300,N_2314,N_2170);
nor UO_301 (O_301,N_2802,N_2150);
or UO_302 (O_302,N_2157,N_2453);
or UO_303 (O_303,N_2996,N_2280);
nand UO_304 (O_304,N_2160,N_2759);
xnor UO_305 (O_305,N_2650,N_2163);
and UO_306 (O_306,N_2985,N_2137);
nor UO_307 (O_307,N_2782,N_2398);
xnor UO_308 (O_308,N_2031,N_2820);
nand UO_309 (O_309,N_2901,N_2801);
or UO_310 (O_310,N_2342,N_2333);
nor UO_311 (O_311,N_2670,N_2577);
or UO_312 (O_312,N_2156,N_2425);
or UO_313 (O_313,N_2855,N_2800);
and UO_314 (O_314,N_2340,N_2645);
and UO_315 (O_315,N_2428,N_2723);
nor UO_316 (O_316,N_2009,N_2471);
xor UO_317 (O_317,N_2767,N_2955);
and UO_318 (O_318,N_2339,N_2680);
and UO_319 (O_319,N_2097,N_2249);
xnor UO_320 (O_320,N_2769,N_2498);
nand UO_321 (O_321,N_2681,N_2739);
or UO_322 (O_322,N_2330,N_2262);
nand UO_323 (O_323,N_2916,N_2034);
nand UO_324 (O_324,N_2635,N_2158);
nand UO_325 (O_325,N_2908,N_2382);
or UO_326 (O_326,N_2209,N_2174);
and UO_327 (O_327,N_2816,N_2652);
or UO_328 (O_328,N_2571,N_2131);
nand UO_329 (O_329,N_2018,N_2143);
or UO_330 (O_330,N_2981,N_2537);
nor UO_331 (O_331,N_2660,N_2598);
and UO_332 (O_332,N_2507,N_2904);
or UO_333 (O_333,N_2753,N_2183);
nand UO_334 (O_334,N_2064,N_2162);
or UO_335 (O_335,N_2865,N_2378);
or UO_336 (O_336,N_2493,N_2233);
nor UO_337 (O_337,N_2323,N_2159);
nor UO_338 (O_338,N_2437,N_2070);
and UO_339 (O_339,N_2033,N_2227);
nor UO_340 (O_340,N_2401,N_2178);
nor UO_341 (O_341,N_2862,N_2619);
nor UO_342 (O_342,N_2970,N_2902);
and UO_343 (O_343,N_2232,N_2710);
or UO_344 (O_344,N_2754,N_2237);
xnor UO_345 (O_345,N_2806,N_2145);
and UO_346 (O_346,N_2484,N_2548);
xnor UO_347 (O_347,N_2094,N_2602);
or UO_348 (O_348,N_2761,N_2565);
nand UO_349 (O_349,N_2438,N_2796);
nand UO_350 (O_350,N_2241,N_2522);
xor UO_351 (O_351,N_2631,N_2368);
or UO_352 (O_352,N_2013,N_2773);
nor UO_353 (O_353,N_2659,N_2999);
xnor UO_354 (O_354,N_2524,N_2003);
xnor UO_355 (O_355,N_2642,N_2793);
nor UO_356 (O_356,N_2201,N_2848);
or UO_357 (O_357,N_2202,N_2930);
xor UO_358 (O_358,N_2858,N_2293);
nor UO_359 (O_359,N_2521,N_2058);
nor UO_360 (O_360,N_2688,N_2692);
nor UO_361 (O_361,N_2722,N_2135);
or UO_362 (O_362,N_2297,N_2075);
nand UO_363 (O_363,N_2549,N_2244);
nand UO_364 (O_364,N_2764,N_2629);
nand UO_365 (O_365,N_2601,N_2856);
nand UO_366 (O_366,N_2165,N_2511);
nor UO_367 (O_367,N_2532,N_2254);
or UO_368 (O_368,N_2695,N_2712);
nor UO_369 (O_369,N_2673,N_2116);
and UO_370 (O_370,N_2744,N_2264);
or UO_371 (O_371,N_2784,N_2421);
or UO_372 (O_372,N_2525,N_2938);
nor UO_373 (O_373,N_2638,N_2104);
nand UO_374 (O_374,N_2982,N_2573);
or UO_375 (O_375,N_2387,N_2391);
nor UO_376 (O_376,N_2349,N_2948);
or UO_377 (O_377,N_2461,N_2300);
or UO_378 (O_378,N_2044,N_2102);
and UO_379 (O_379,N_2226,N_2068);
or UO_380 (O_380,N_2354,N_2977);
and UO_381 (O_381,N_2288,N_2057);
nor UO_382 (O_382,N_2063,N_2375);
and UO_383 (O_383,N_2040,N_2871);
or UO_384 (O_384,N_2402,N_2986);
or UO_385 (O_385,N_2752,N_2103);
and UO_386 (O_386,N_2915,N_2536);
nand UO_387 (O_387,N_2409,N_2203);
nor UO_388 (O_388,N_2161,N_2327);
or UO_389 (O_389,N_2900,N_2483);
or UO_390 (O_390,N_2355,N_2497);
nor UO_391 (O_391,N_2210,N_2054);
xnor UO_392 (O_392,N_2823,N_2060);
nor UO_393 (O_393,N_2015,N_2359);
nand UO_394 (O_394,N_2864,N_2222);
nor UO_395 (O_395,N_2667,N_2390);
nor UO_396 (O_396,N_2247,N_2763);
or UO_397 (O_397,N_2199,N_2035);
and UO_398 (O_398,N_2189,N_2922);
and UO_399 (O_399,N_2805,N_2166);
xnor UO_400 (O_400,N_2931,N_2678);
nand UO_401 (O_401,N_2748,N_2325);
nand UO_402 (O_402,N_2877,N_2956);
or UO_403 (O_403,N_2539,N_2289);
and UO_404 (O_404,N_2192,N_2149);
and UO_405 (O_405,N_2491,N_2474);
nor UO_406 (O_406,N_2656,N_2422);
or UO_407 (O_407,N_2750,N_2124);
nand UO_408 (O_408,N_2995,N_2960);
and UO_409 (O_409,N_2141,N_2386);
nor UO_410 (O_410,N_2884,N_2926);
nor UO_411 (O_411,N_2809,N_2766);
nor UO_412 (O_412,N_2403,N_2367);
and UO_413 (O_413,N_2373,N_2917);
and UO_414 (O_414,N_2286,N_2604);
or UO_415 (O_415,N_2444,N_2513);
nor UO_416 (O_416,N_2169,N_2406);
and UO_417 (O_417,N_2705,N_2893);
or UO_418 (O_418,N_2732,N_2776);
or UO_419 (O_419,N_2316,N_2624);
nand UO_420 (O_420,N_2563,N_2011);
or UO_421 (O_421,N_2433,N_2121);
or UO_422 (O_422,N_2934,N_2881);
or UO_423 (O_423,N_2853,N_2817);
or UO_424 (O_424,N_2622,N_2742);
and UO_425 (O_425,N_2074,N_2252);
or UO_426 (O_426,N_2863,N_2778);
or UO_427 (O_427,N_2418,N_2039);
nand UO_428 (O_428,N_2480,N_2510);
xnor UO_429 (O_429,N_2026,N_2317);
and UO_430 (O_430,N_2634,N_2105);
and UO_431 (O_431,N_2815,N_2574);
xor UO_432 (O_432,N_2489,N_2181);
nor UO_433 (O_433,N_2299,N_2164);
and UO_434 (O_434,N_2207,N_2758);
xor UO_435 (O_435,N_2949,N_2278);
nor UO_436 (O_436,N_2792,N_2361);
nor UO_437 (O_437,N_2626,N_2478);
or UO_438 (O_438,N_2371,N_2797);
or UO_439 (O_439,N_2777,N_2405);
or UO_440 (O_440,N_2427,N_2188);
and UO_441 (O_441,N_2835,N_2526);
nand UO_442 (O_442,N_2492,N_2487);
and UO_443 (O_443,N_2730,N_2841);
or UO_444 (O_444,N_2535,N_2463);
nor UO_445 (O_445,N_2516,N_2918);
nor UO_446 (O_446,N_2909,N_2663);
and UO_447 (O_447,N_2887,N_2310);
and UO_448 (O_448,N_2671,N_2546);
or UO_449 (O_449,N_2184,N_2873);
nand UO_450 (O_450,N_2256,N_2231);
nand UO_451 (O_451,N_2067,N_2495);
nand UO_452 (O_452,N_2939,N_2731);
and UO_453 (O_453,N_2775,N_2032);
nor UO_454 (O_454,N_2048,N_2849);
or UO_455 (O_455,N_2127,N_2221);
nand UO_456 (O_456,N_2941,N_2697);
nor UO_457 (O_457,N_2118,N_2399);
or UO_458 (O_458,N_2305,N_2128);
and UO_459 (O_459,N_2343,N_2694);
or UO_460 (O_460,N_2329,N_2434);
or UO_461 (O_461,N_2168,N_2021);
nand UO_462 (O_462,N_2146,N_2380);
nor UO_463 (O_463,N_2318,N_2260);
or UO_464 (O_464,N_2531,N_2185);
or UO_465 (O_465,N_2737,N_2812);
or UO_466 (O_466,N_2078,N_2198);
or UO_467 (O_467,N_2000,N_2459);
nand UO_468 (O_468,N_2351,N_2357);
or UO_469 (O_469,N_2620,N_2279);
or UO_470 (O_470,N_2322,N_2515);
and UO_471 (O_471,N_2868,N_2988);
nor UO_472 (O_472,N_2377,N_2693);
xor UO_473 (O_473,N_2328,N_2508);
and UO_474 (O_474,N_2711,N_2107);
or UO_475 (O_475,N_2690,N_2544);
nor UO_476 (O_476,N_2248,N_2974);
nand UO_477 (O_477,N_2374,N_2822);
and UO_478 (O_478,N_2376,N_2324);
nor UO_479 (O_479,N_2123,N_2586);
and UO_480 (O_480,N_2755,N_2379);
nand UO_481 (O_481,N_2745,N_2606);
or UO_482 (O_482,N_2929,N_2215);
and UO_483 (O_483,N_2270,N_2144);
nand UO_484 (O_484,N_2665,N_2010);
nor UO_485 (O_485,N_2933,N_2772);
or UO_486 (O_486,N_2839,N_2084);
nand UO_487 (O_487,N_2196,N_2235);
nor UO_488 (O_488,N_2259,N_2028);
nor UO_489 (O_489,N_2341,N_2727);
nor UO_490 (O_490,N_2924,N_2890);
nor UO_491 (O_491,N_2413,N_2024);
or UO_492 (O_492,N_2741,N_2212);
nand UO_493 (O_493,N_2025,N_2892);
and UO_494 (O_494,N_2911,N_2369);
or UO_495 (O_495,N_2083,N_2223);
or UO_496 (O_496,N_2630,N_2458);
and UO_497 (O_497,N_2108,N_2649);
nor UO_498 (O_498,N_2953,N_2859);
nor UO_499 (O_499,N_2559,N_2984);
endmodule