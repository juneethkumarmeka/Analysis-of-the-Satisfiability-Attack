module basic_750_5000_1000_10_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
xor U0 (N_0,In_335,In_165);
nor U1 (N_1,In_138,In_734);
and U2 (N_2,In_281,In_403);
nand U3 (N_3,In_436,In_314);
and U4 (N_4,In_354,In_192);
nor U5 (N_5,In_630,In_680);
or U6 (N_6,In_116,In_455);
xnor U7 (N_7,In_329,In_157);
xnor U8 (N_8,In_635,In_568);
nand U9 (N_9,In_23,In_505);
or U10 (N_10,In_544,In_285);
nand U11 (N_11,In_200,In_178);
nand U12 (N_12,In_631,In_690);
nand U13 (N_13,In_91,In_357);
or U14 (N_14,In_307,In_208);
nor U15 (N_15,In_124,In_209);
or U16 (N_16,In_614,In_684);
nor U17 (N_17,In_168,In_177);
xor U18 (N_18,In_400,In_601);
or U19 (N_19,In_180,In_310);
xor U20 (N_20,In_615,In_741);
nor U21 (N_21,In_462,In_582);
nand U22 (N_22,In_540,In_569);
nor U23 (N_23,In_426,In_437);
nand U24 (N_24,In_340,In_586);
and U25 (N_25,In_243,In_632);
or U26 (N_26,In_146,In_244);
nand U27 (N_27,In_738,In_578);
and U28 (N_28,In_351,In_583);
or U29 (N_29,In_737,In_464);
and U30 (N_30,In_317,In_451);
nor U31 (N_31,In_654,In_519);
nor U32 (N_32,In_158,In_383);
nor U33 (N_33,In_644,In_401);
and U34 (N_34,In_167,In_486);
and U35 (N_35,In_723,In_139);
and U36 (N_36,In_12,In_114);
or U37 (N_37,In_602,In_597);
nand U38 (N_38,In_106,In_82);
or U39 (N_39,In_699,In_604);
and U40 (N_40,In_560,In_298);
nor U41 (N_41,In_217,In_66);
or U42 (N_42,In_274,In_236);
or U43 (N_43,In_56,In_170);
nand U44 (N_44,In_350,In_34);
nand U45 (N_45,In_683,In_725);
nand U46 (N_46,In_358,In_223);
or U47 (N_47,In_376,In_360);
nor U48 (N_48,In_619,In_598);
nor U49 (N_49,In_570,In_131);
or U50 (N_50,In_364,In_29);
xor U51 (N_51,In_117,In_469);
or U52 (N_52,In_641,In_506);
and U53 (N_53,In_443,In_390);
and U54 (N_54,In_704,In_380);
or U55 (N_55,In_160,In_149);
or U56 (N_56,In_190,In_304);
nor U57 (N_57,In_674,In_418);
xnor U58 (N_58,In_42,In_64);
or U59 (N_59,In_458,In_435);
and U60 (N_60,In_652,In_130);
or U61 (N_61,In_471,In_466);
xnor U62 (N_62,In_341,In_36);
nand U63 (N_63,In_522,In_457);
or U64 (N_64,In_148,In_186);
or U65 (N_65,In_361,In_521);
or U66 (N_66,In_487,In_71);
or U67 (N_67,In_573,In_20);
nand U68 (N_68,In_97,In_491);
or U69 (N_69,In_474,In_103);
nand U70 (N_70,In_219,In_156);
and U71 (N_71,In_293,In_695);
nor U72 (N_72,In_502,In_470);
nand U73 (N_73,In_442,In_323);
nand U74 (N_74,In_107,In_255);
nor U75 (N_75,In_639,In_137);
nand U76 (N_76,In_567,In_580);
and U77 (N_77,In_83,In_254);
xor U78 (N_78,In_332,In_478);
nor U79 (N_79,In_270,In_536);
nor U80 (N_80,In_9,In_104);
and U81 (N_81,In_239,In_182);
and U82 (N_82,In_133,In_689);
xnor U83 (N_83,In_269,In_155);
or U84 (N_84,In_425,In_265);
xor U85 (N_85,In_11,In_444);
and U86 (N_86,In_539,In_296);
nand U87 (N_87,In_241,In_132);
nor U88 (N_88,In_245,In_108);
nor U89 (N_89,In_185,In_111);
and U90 (N_90,In_678,In_234);
nand U91 (N_91,In_144,In_284);
nor U92 (N_92,In_414,In_685);
or U93 (N_93,In_187,In_735);
or U94 (N_94,In_384,In_183);
nor U95 (N_95,In_608,In_375);
nand U96 (N_96,In_480,In_694);
nor U97 (N_97,In_647,In_159);
and U98 (N_98,In_365,In_371);
nor U99 (N_99,In_579,In_93);
or U100 (N_100,In_589,In_413);
nor U101 (N_101,In_657,In_55);
and U102 (N_102,In_382,In_69);
nor U103 (N_103,In_113,In_295);
nor U104 (N_104,In_74,In_460);
nand U105 (N_105,In_336,In_507);
nor U106 (N_106,In_433,In_525);
xor U107 (N_107,In_634,In_423);
nor U108 (N_108,In_417,In_710);
and U109 (N_109,In_542,In_653);
nand U110 (N_110,In_261,In_708);
nor U111 (N_111,In_465,In_247);
or U112 (N_112,In_687,In_575);
and U113 (N_113,In_272,In_89);
or U114 (N_114,In_225,In_297);
nor U115 (N_115,In_421,In_19);
or U116 (N_116,In_289,In_98);
or U117 (N_117,In_729,In_529);
or U118 (N_118,In_370,In_587);
and U119 (N_119,In_576,In_603);
and U120 (N_120,In_324,In_612);
or U121 (N_121,In_744,In_681);
and U122 (N_122,In_299,In_260);
nor U123 (N_123,In_745,In_176);
nand U124 (N_124,In_720,In_659);
nor U125 (N_125,In_327,In_218);
and U126 (N_126,In_456,In_326);
nand U127 (N_127,In_22,In_488);
nand U128 (N_128,In_196,In_584);
or U129 (N_129,In_268,In_682);
nor U130 (N_130,In_292,In_562);
nand U131 (N_131,In_731,In_303);
nand U132 (N_132,In_571,In_651);
and U133 (N_133,In_238,In_668);
or U134 (N_134,In_367,In_495);
or U135 (N_135,In_319,In_422);
and U136 (N_136,In_10,In_445);
nand U137 (N_137,In_4,In_408);
and U138 (N_138,In_724,In_561);
nand U139 (N_139,In_730,In_161);
xnor U140 (N_140,In_275,In_102);
nand U141 (N_141,In_393,In_179);
nor U142 (N_142,In_482,In_429);
and U143 (N_143,In_728,In_153);
or U144 (N_144,In_688,In_496);
or U145 (N_145,In_59,In_483);
or U146 (N_146,In_88,In_100);
nor U147 (N_147,In_169,In_8);
nand U148 (N_148,In_16,In_611);
xnor U149 (N_149,In_325,In_676);
nor U150 (N_150,In_534,In_385);
xor U151 (N_151,In_701,In_171);
nand U152 (N_152,In_337,In_191);
xor U153 (N_153,In_472,In_321);
nand U154 (N_154,In_650,In_527);
or U155 (N_155,In_373,In_347);
nor U156 (N_156,In_151,In_585);
nand U157 (N_157,In_553,In_546);
and U158 (N_158,In_248,In_44);
xor U159 (N_159,In_342,In_645);
or U160 (N_160,In_428,In_447);
nor U161 (N_161,In_606,In_99);
or U162 (N_162,In_345,In_147);
nand U163 (N_163,In_212,In_92);
or U164 (N_164,In_353,In_748);
nor U165 (N_165,In_698,In_621);
nor U166 (N_166,In_391,In_713);
or U167 (N_167,In_90,In_705);
or U168 (N_168,In_467,In_476);
xnor U169 (N_169,In_600,In_162);
or U170 (N_170,In_312,In_714);
and U171 (N_171,In_438,In_60);
nand U172 (N_172,In_271,In_202);
nor U173 (N_173,In_520,In_221);
nand U174 (N_174,In_331,In_294);
xnor U175 (N_175,In_649,In_381);
nand U176 (N_176,In_38,In_564);
or U177 (N_177,In_5,In_508);
nand U178 (N_178,In_446,In_229);
nor U179 (N_179,In_677,In_172);
and U180 (N_180,In_660,In_300);
nand U181 (N_181,In_78,In_95);
and U182 (N_182,In_646,In_626);
and U183 (N_183,In_552,In_70);
nor U184 (N_184,In_313,In_510);
nand U185 (N_185,In_454,In_712);
xor U186 (N_186,In_87,In_431);
nor U187 (N_187,In_302,In_369);
and U188 (N_188,In_112,In_715);
or U189 (N_189,In_427,In_374);
and U190 (N_190,In_96,In_493);
or U191 (N_191,In_499,In_45);
nor U192 (N_192,In_625,In_49);
nor U193 (N_193,In_85,In_3);
nor U194 (N_194,In_35,In_81);
nor U195 (N_195,In_204,In_309);
and U196 (N_196,In_105,In_581);
nand U197 (N_197,In_194,In_363);
nor U198 (N_198,In_51,In_258);
nor U199 (N_199,In_13,In_516);
and U200 (N_200,In_63,In_226);
nand U201 (N_201,In_407,In_339);
or U202 (N_202,In_419,In_173);
nor U203 (N_203,In_14,In_605);
nand U204 (N_204,In_711,In_101);
and U205 (N_205,In_287,In_57);
or U206 (N_206,In_262,In_468);
nor U207 (N_207,In_230,In_152);
and U208 (N_208,In_749,In_432);
and U209 (N_209,In_637,In_322);
or U210 (N_210,In_727,In_141);
and U211 (N_211,In_648,In_420);
and U212 (N_212,In_37,In_150);
nand U213 (N_213,In_256,In_532);
or U214 (N_214,In_566,In_500);
and U215 (N_215,In_206,In_18);
xnor U216 (N_216,In_479,In_662);
and U217 (N_217,In_28,In_592);
nor U218 (N_218,In_237,In_41);
or U219 (N_219,In_665,In_377);
nand U220 (N_220,In_477,In_747);
nand U221 (N_221,In_278,In_291);
or U222 (N_222,In_80,In_618);
or U223 (N_223,In_555,In_328);
nand U224 (N_224,In_609,In_216);
and U225 (N_225,In_207,In_15);
or U226 (N_226,In_263,In_617);
nor U227 (N_227,In_128,In_246);
nor U228 (N_228,In_175,In_655);
or U229 (N_229,In_40,In_693);
nand U230 (N_230,In_283,In_633);
nor U231 (N_231,In_355,In_197);
nor U232 (N_232,In_249,In_214);
nand U233 (N_233,In_61,In_703);
nand U234 (N_234,In_242,In_231);
or U235 (N_235,In_228,In_2);
and U236 (N_236,In_671,In_742);
nand U237 (N_237,In_475,In_181);
or U238 (N_238,In_453,In_76);
and U239 (N_239,In_675,In_664);
nand U240 (N_240,In_352,In_129);
or U241 (N_241,In_563,In_115);
and U242 (N_242,In_174,In_697);
nand U243 (N_243,In_613,In_308);
or U244 (N_244,In_0,In_473);
or U245 (N_245,In_679,In_515);
nand U246 (N_246,In_222,In_94);
nor U247 (N_247,In_389,In_590);
nand U248 (N_248,In_395,In_224);
nand U249 (N_249,In_514,In_315);
and U250 (N_250,In_538,In_122);
and U251 (N_251,In_548,In_557);
or U252 (N_252,In_610,In_667);
nor U253 (N_253,In_349,In_253);
nand U254 (N_254,In_193,In_378);
and U255 (N_255,In_398,In_526);
nor U256 (N_256,In_368,In_485);
or U257 (N_257,In_338,In_392);
and U258 (N_258,In_346,In_53);
nand U259 (N_259,In_556,In_356);
and U260 (N_260,In_732,In_558);
or U261 (N_261,In_402,In_50);
or U262 (N_262,In_524,In_490);
nand U263 (N_263,In_84,In_448);
and U264 (N_264,In_692,In_276);
or U265 (N_265,In_424,In_541);
nand U266 (N_266,In_73,In_623);
nor U267 (N_267,In_233,In_545);
xor U268 (N_268,In_673,In_52);
nor U269 (N_269,In_142,In_127);
xor U270 (N_270,In_547,In_126);
nand U271 (N_271,In_559,In_288);
nor U272 (N_272,In_17,In_620);
xor U273 (N_273,In_593,In_210);
or U274 (N_274,In_492,In_517);
nor U275 (N_275,In_565,In_27);
and U276 (N_276,In_594,In_627);
xor U277 (N_277,In_201,In_643);
nor U278 (N_278,In_1,In_449);
xor U279 (N_279,In_706,In_717);
nand U280 (N_280,In_386,In_109);
and U281 (N_281,In_533,In_195);
or U282 (N_282,In_461,In_79);
nor U283 (N_283,In_595,In_397);
nand U284 (N_284,In_316,In_118);
or U285 (N_285,In_740,In_415);
and U286 (N_286,In_250,In_77);
nand U287 (N_287,In_504,In_509);
xor U288 (N_288,In_702,In_251);
and U289 (N_289,In_722,In_199);
nor U290 (N_290,In_232,In_333);
or U291 (N_291,In_188,In_743);
or U292 (N_292,In_718,In_624);
nor U293 (N_293,In_136,In_434);
and U294 (N_294,In_135,In_26);
nand U295 (N_295,In_394,In_640);
nand U296 (N_296,In_362,In_588);
or U297 (N_297,In_72,In_290);
xor U298 (N_298,In_24,In_119);
and U299 (N_299,In_43,In_489);
nand U300 (N_300,In_387,In_622);
and U301 (N_301,In_301,In_551);
and U302 (N_302,In_707,In_372);
or U303 (N_303,In_543,In_359);
nor U304 (N_304,In_240,In_198);
and U305 (N_305,In_279,In_125);
nand U306 (N_306,In_33,In_535);
or U307 (N_307,In_670,In_320);
nand U308 (N_308,In_145,In_691);
xor U309 (N_309,In_518,In_86);
nand U310 (N_310,In_220,In_409);
nand U311 (N_311,In_48,In_215);
nand U312 (N_312,In_656,In_379);
or U313 (N_313,In_334,In_596);
or U314 (N_314,In_628,In_512);
nand U315 (N_315,In_528,In_503);
nand U316 (N_316,In_58,In_235);
nand U317 (N_317,In_54,In_67);
and U318 (N_318,In_366,In_252);
xnor U319 (N_319,In_412,In_616);
or U320 (N_320,In_348,In_638);
xnor U321 (N_321,In_75,In_497);
nor U322 (N_322,In_266,In_163);
and U323 (N_323,In_642,In_746);
nor U324 (N_324,In_666,In_31);
nand U325 (N_325,In_7,In_134);
and U326 (N_326,In_411,In_405);
nor U327 (N_327,In_452,In_531);
nor U328 (N_328,In_550,In_166);
xnor U329 (N_329,In_62,In_410);
xnor U330 (N_330,In_513,In_661);
nand U331 (N_331,In_65,In_591);
xnor U332 (N_332,In_574,In_629);
nand U333 (N_333,In_343,In_686);
nor U334 (N_334,In_481,In_404);
nor U335 (N_335,In_273,In_154);
nand U336 (N_336,In_733,In_277);
nand U337 (N_337,In_709,In_416);
and U338 (N_338,In_306,In_396);
and U339 (N_339,In_32,In_399);
nor U340 (N_340,In_439,In_484);
nor U341 (N_341,In_719,In_658);
nand U342 (N_342,In_110,In_184);
or U343 (N_343,In_311,In_120);
nand U344 (N_344,In_523,In_286);
nand U345 (N_345,In_47,In_282);
nor U346 (N_346,In_121,In_39);
and U347 (N_347,In_463,In_46);
xor U348 (N_348,In_68,In_736);
or U349 (N_349,In_259,In_123);
or U350 (N_350,In_318,In_721);
nor U351 (N_351,In_267,In_501);
nor U352 (N_352,In_388,In_498);
and U353 (N_353,In_672,In_599);
or U354 (N_354,In_305,In_636);
nor U355 (N_355,In_450,In_164);
nand U356 (N_356,In_21,In_537);
nor U357 (N_357,In_494,In_716);
or U358 (N_358,In_572,In_6);
nor U359 (N_359,In_430,In_440);
or U360 (N_360,In_280,In_663);
nand U361 (N_361,In_143,In_203);
or U362 (N_362,In_739,In_607);
and U363 (N_363,In_577,In_140);
and U364 (N_364,In_511,In_549);
nor U365 (N_365,In_257,In_696);
nor U366 (N_366,In_669,In_406);
nor U367 (N_367,In_530,In_30);
xnor U368 (N_368,In_264,In_205);
nor U369 (N_369,In_211,In_700);
xor U370 (N_370,In_25,In_441);
xnor U371 (N_371,In_189,In_726);
xnor U372 (N_372,In_344,In_213);
nand U373 (N_373,In_330,In_554);
nor U374 (N_374,In_227,In_459);
or U375 (N_375,In_626,In_513);
nand U376 (N_376,In_107,In_303);
or U377 (N_377,In_263,In_476);
or U378 (N_378,In_118,In_240);
nor U379 (N_379,In_193,In_698);
or U380 (N_380,In_465,In_128);
or U381 (N_381,In_717,In_452);
or U382 (N_382,In_249,In_5);
nor U383 (N_383,In_103,In_570);
nand U384 (N_384,In_605,In_457);
xor U385 (N_385,In_474,In_414);
or U386 (N_386,In_287,In_117);
nor U387 (N_387,In_211,In_360);
nand U388 (N_388,In_563,In_519);
and U389 (N_389,In_289,In_609);
or U390 (N_390,In_389,In_319);
nor U391 (N_391,In_88,In_134);
and U392 (N_392,In_684,In_202);
or U393 (N_393,In_613,In_79);
and U394 (N_394,In_111,In_434);
nor U395 (N_395,In_599,In_734);
and U396 (N_396,In_167,In_603);
xor U397 (N_397,In_742,In_110);
nand U398 (N_398,In_709,In_507);
nand U399 (N_399,In_289,In_85);
xnor U400 (N_400,In_553,In_267);
or U401 (N_401,In_649,In_41);
nand U402 (N_402,In_75,In_384);
and U403 (N_403,In_586,In_425);
and U404 (N_404,In_181,In_410);
nor U405 (N_405,In_695,In_386);
nor U406 (N_406,In_597,In_5);
nand U407 (N_407,In_455,In_359);
and U408 (N_408,In_450,In_144);
or U409 (N_409,In_56,In_270);
and U410 (N_410,In_154,In_97);
nand U411 (N_411,In_727,In_748);
nor U412 (N_412,In_743,In_538);
and U413 (N_413,In_411,In_292);
and U414 (N_414,In_695,In_127);
and U415 (N_415,In_328,In_36);
or U416 (N_416,In_60,In_336);
or U417 (N_417,In_295,In_397);
nand U418 (N_418,In_47,In_248);
and U419 (N_419,In_364,In_315);
xor U420 (N_420,In_512,In_190);
nor U421 (N_421,In_742,In_309);
nand U422 (N_422,In_471,In_650);
nand U423 (N_423,In_169,In_667);
nor U424 (N_424,In_225,In_561);
and U425 (N_425,In_395,In_239);
or U426 (N_426,In_495,In_65);
xnor U427 (N_427,In_548,In_37);
nor U428 (N_428,In_697,In_260);
nor U429 (N_429,In_317,In_450);
nand U430 (N_430,In_650,In_688);
nor U431 (N_431,In_361,In_267);
and U432 (N_432,In_398,In_375);
nor U433 (N_433,In_282,In_663);
or U434 (N_434,In_735,In_33);
nor U435 (N_435,In_421,In_202);
nor U436 (N_436,In_394,In_391);
or U437 (N_437,In_229,In_37);
and U438 (N_438,In_274,In_611);
nand U439 (N_439,In_435,In_702);
and U440 (N_440,In_346,In_676);
nor U441 (N_441,In_325,In_174);
nor U442 (N_442,In_664,In_243);
nand U443 (N_443,In_313,In_509);
and U444 (N_444,In_586,In_578);
nor U445 (N_445,In_546,In_607);
nand U446 (N_446,In_328,In_258);
xor U447 (N_447,In_554,In_729);
nand U448 (N_448,In_28,In_17);
nor U449 (N_449,In_675,In_635);
nand U450 (N_450,In_499,In_253);
or U451 (N_451,In_50,In_407);
nor U452 (N_452,In_699,In_215);
and U453 (N_453,In_407,In_576);
or U454 (N_454,In_92,In_522);
nand U455 (N_455,In_563,In_15);
nand U456 (N_456,In_542,In_544);
xor U457 (N_457,In_371,In_668);
nand U458 (N_458,In_698,In_611);
nand U459 (N_459,In_12,In_361);
xnor U460 (N_460,In_607,In_14);
or U461 (N_461,In_370,In_581);
xnor U462 (N_462,In_440,In_583);
nand U463 (N_463,In_566,In_625);
xor U464 (N_464,In_27,In_485);
and U465 (N_465,In_583,In_565);
and U466 (N_466,In_582,In_647);
nand U467 (N_467,In_644,In_5);
nand U468 (N_468,In_108,In_438);
nand U469 (N_469,In_51,In_683);
nor U470 (N_470,In_120,In_264);
nor U471 (N_471,In_454,In_13);
nor U472 (N_472,In_242,In_169);
nor U473 (N_473,In_682,In_222);
nor U474 (N_474,In_151,In_524);
nand U475 (N_475,In_451,In_252);
nand U476 (N_476,In_439,In_524);
nor U477 (N_477,In_175,In_341);
xnor U478 (N_478,In_282,In_172);
nand U479 (N_479,In_386,In_669);
and U480 (N_480,In_413,In_416);
and U481 (N_481,In_220,In_469);
and U482 (N_482,In_675,In_32);
nand U483 (N_483,In_741,In_127);
nand U484 (N_484,In_593,In_731);
nand U485 (N_485,In_243,In_565);
xor U486 (N_486,In_338,In_346);
nor U487 (N_487,In_606,In_707);
nand U488 (N_488,In_206,In_558);
and U489 (N_489,In_464,In_354);
or U490 (N_490,In_338,In_361);
and U491 (N_491,In_703,In_336);
nor U492 (N_492,In_287,In_515);
and U493 (N_493,In_514,In_438);
and U494 (N_494,In_159,In_477);
xor U495 (N_495,In_84,In_14);
nand U496 (N_496,In_237,In_691);
and U497 (N_497,In_259,In_622);
nor U498 (N_498,In_554,In_268);
nor U499 (N_499,In_253,In_563);
nor U500 (N_500,N_476,N_461);
nor U501 (N_501,N_363,N_224);
or U502 (N_502,N_244,N_340);
nand U503 (N_503,N_339,N_129);
xor U504 (N_504,N_283,N_300);
nand U505 (N_505,N_118,N_59);
nand U506 (N_506,N_314,N_178);
nand U507 (N_507,N_425,N_409);
and U508 (N_508,N_215,N_307);
or U509 (N_509,N_234,N_305);
nand U510 (N_510,N_399,N_445);
nor U511 (N_511,N_172,N_334);
xnor U512 (N_512,N_5,N_127);
or U513 (N_513,N_359,N_406);
or U514 (N_514,N_130,N_405);
and U515 (N_515,N_472,N_190);
xnor U516 (N_516,N_8,N_96);
and U517 (N_517,N_411,N_344);
nor U518 (N_518,N_140,N_350);
nor U519 (N_519,N_120,N_413);
and U520 (N_520,N_138,N_100);
nor U521 (N_521,N_349,N_122);
or U522 (N_522,N_163,N_309);
nand U523 (N_523,N_115,N_391);
nor U524 (N_524,N_70,N_203);
nand U525 (N_525,N_225,N_210);
and U526 (N_526,N_422,N_331);
and U527 (N_527,N_471,N_173);
nand U528 (N_528,N_449,N_368);
and U529 (N_529,N_12,N_437);
and U530 (N_530,N_328,N_342);
nor U531 (N_531,N_117,N_250);
or U532 (N_532,N_369,N_407);
or U533 (N_533,N_373,N_160);
and U534 (N_534,N_237,N_183);
xnor U535 (N_535,N_343,N_306);
and U536 (N_536,N_86,N_470);
or U537 (N_537,N_231,N_92);
xor U538 (N_538,N_208,N_410);
or U539 (N_539,N_91,N_3);
nor U540 (N_540,N_474,N_47);
and U541 (N_541,N_150,N_416);
and U542 (N_542,N_301,N_321);
or U543 (N_543,N_319,N_477);
nand U544 (N_544,N_311,N_2);
xor U545 (N_545,N_49,N_459);
nor U546 (N_546,N_336,N_93);
or U547 (N_547,N_146,N_226);
nand U548 (N_548,N_73,N_443);
or U549 (N_549,N_255,N_191);
nor U550 (N_550,N_478,N_176);
nor U551 (N_551,N_356,N_290);
or U552 (N_552,N_25,N_376);
nand U553 (N_553,N_98,N_281);
nand U554 (N_554,N_389,N_168);
nor U555 (N_555,N_157,N_372);
nand U556 (N_556,N_317,N_392);
and U557 (N_557,N_132,N_291);
and U558 (N_558,N_421,N_209);
nor U559 (N_559,N_415,N_324);
and U560 (N_560,N_345,N_329);
and U561 (N_561,N_29,N_180);
nand U562 (N_562,N_486,N_24);
nand U563 (N_563,N_397,N_35);
and U564 (N_564,N_384,N_196);
and U565 (N_565,N_377,N_275);
and U566 (N_566,N_143,N_412);
nand U567 (N_567,N_76,N_54);
and U568 (N_568,N_362,N_17);
and U569 (N_569,N_94,N_89);
or U570 (N_570,N_465,N_246);
and U571 (N_571,N_330,N_403);
nor U572 (N_572,N_490,N_285);
nand U573 (N_573,N_303,N_77);
and U574 (N_574,N_232,N_274);
and U575 (N_575,N_469,N_82);
nand U576 (N_576,N_308,N_261);
nor U577 (N_577,N_253,N_134);
nor U578 (N_578,N_186,N_39);
and U579 (N_579,N_279,N_154);
nor U580 (N_580,N_189,N_236);
nor U581 (N_581,N_361,N_245);
and U582 (N_582,N_327,N_87);
nand U583 (N_583,N_6,N_464);
or U584 (N_584,N_144,N_105);
nor U585 (N_585,N_444,N_83);
or U586 (N_586,N_278,N_95);
or U587 (N_587,N_165,N_48);
nand U588 (N_588,N_11,N_164);
nor U589 (N_589,N_200,N_45);
nor U590 (N_590,N_346,N_90);
nor U591 (N_591,N_457,N_229);
nor U592 (N_592,N_58,N_204);
nor U593 (N_593,N_55,N_171);
nand U594 (N_594,N_396,N_0);
xnor U595 (N_595,N_153,N_68);
nand U596 (N_596,N_241,N_36);
and U597 (N_597,N_379,N_194);
xor U598 (N_598,N_467,N_254);
and U599 (N_599,N_398,N_7);
nand U600 (N_600,N_33,N_61);
and U601 (N_601,N_497,N_395);
xnor U602 (N_602,N_51,N_71);
nand U603 (N_603,N_66,N_390);
or U604 (N_604,N_259,N_152);
or U605 (N_605,N_431,N_248);
or U606 (N_606,N_142,N_207);
xnor U607 (N_607,N_299,N_374);
nand U608 (N_608,N_136,N_30);
nand U609 (N_609,N_197,N_423);
or U610 (N_610,N_364,N_417);
or U611 (N_611,N_298,N_304);
or U612 (N_612,N_205,N_97);
and U613 (N_613,N_332,N_104);
xnor U614 (N_614,N_460,N_335);
nor U615 (N_615,N_133,N_263);
nand U616 (N_616,N_31,N_62);
nand U617 (N_617,N_267,N_230);
nor U618 (N_618,N_494,N_109);
nand U619 (N_619,N_216,N_260);
nand U620 (N_620,N_108,N_269);
nor U621 (N_621,N_473,N_84);
nor U622 (N_622,N_270,N_318);
nand U623 (N_623,N_13,N_27);
nor U624 (N_624,N_126,N_125);
or U625 (N_625,N_258,N_155);
nor U626 (N_626,N_402,N_135);
and U627 (N_627,N_434,N_371);
nand U628 (N_628,N_74,N_326);
xnor U629 (N_629,N_447,N_441);
nor U630 (N_630,N_139,N_206);
nor U631 (N_631,N_193,N_147);
nand U632 (N_632,N_420,N_440);
nand U633 (N_633,N_316,N_148);
and U634 (N_634,N_375,N_455);
nor U635 (N_635,N_107,N_352);
and U636 (N_636,N_26,N_20);
xnor U637 (N_637,N_401,N_247);
nand U638 (N_638,N_448,N_320);
nor U639 (N_639,N_488,N_22);
or U640 (N_640,N_432,N_454);
or U641 (N_641,N_370,N_427);
or U642 (N_642,N_99,N_9);
or U643 (N_643,N_111,N_60);
nor U644 (N_644,N_498,N_466);
or U645 (N_645,N_458,N_385);
or U646 (N_646,N_158,N_37);
and U647 (N_647,N_451,N_400);
and U648 (N_648,N_348,N_184);
nand U649 (N_649,N_19,N_233);
and U650 (N_650,N_430,N_289);
or U651 (N_651,N_495,N_201);
nor U652 (N_652,N_151,N_264);
nor U653 (N_653,N_212,N_404);
xor U654 (N_654,N_1,N_387);
nand U655 (N_655,N_272,N_10);
and U656 (N_656,N_65,N_337);
nand U657 (N_657,N_295,N_450);
nand U658 (N_658,N_428,N_78);
and U659 (N_659,N_169,N_79);
nor U660 (N_660,N_288,N_195);
nor U661 (N_661,N_333,N_322);
and U662 (N_662,N_42,N_439);
nand U663 (N_663,N_175,N_141);
nor U664 (N_664,N_463,N_475);
nor U665 (N_665,N_192,N_338);
or U666 (N_666,N_75,N_182);
and U667 (N_667,N_214,N_43);
nor U668 (N_668,N_493,N_88);
nor U669 (N_669,N_199,N_102);
nand U670 (N_670,N_491,N_67);
nand U671 (N_671,N_360,N_174);
nor U672 (N_672,N_456,N_185);
xor U673 (N_673,N_177,N_161);
and U674 (N_674,N_251,N_365);
nand U675 (N_675,N_44,N_277);
or U676 (N_676,N_149,N_357);
nand U677 (N_677,N_81,N_103);
nor U678 (N_678,N_284,N_483);
nand U679 (N_679,N_38,N_221);
nand U680 (N_680,N_121,N_57);
nor U681 (N_681,N_46,N_426);
and U682 (N_682,N_114,N_63);
nor U683 (N_683,N_280,N_293);
nor U684 (N_684,N_489,N_167);
or U685 (N_685,N_266,N_452);
or U686 (N_686,N_315,N_419);
or U687 (N_687,N_156,N_367);
nand U688 (N_688,N_162,N_499);
or U689 (N_689,N_496,N_223);
or U690 (N_690,N_468,N_113);
and U691 (N_691,N_145,N_380);
xnor U692 (N_692,N_313,N_128);
nor U693 (N_693,N_242,N_179);
nand U694 (N_694,N_323,N_124);
or U695 (N_695,N_249,N_28);
nand U696 (N_696,N_351,N_282);
or U697 (N_697,N_383,N_453);
nand U698 (N_698,N_442,N_238);
nor U699 (N_699,N_462,N_424);
and U700 (N_700,N_271,N_482);
or U701 (N_701,N_85,N_41);
nor U702 (N_702,N_481,N_292);
nor U703 (N_703,N_227,N_235);
and U704 (N_704,N_276,N_408);
nor U705 (N_705,N_492,N_256);
or U706 (N_706,N_378,N_265);
nand U707 (N_707,N_435,N_56);
nor U708 (N_708,N_222,N_341);
nand U709 (N_709,N_50,N_72);
nand U710 (N_710,N_347,N_418);
or U711 (N_711,N_257,N_294);
and U712 (N_712,N_262,N_312);
xor U713 (N_713,N_297,N_446);
nand U714 (N_714,N_388,N_53);
or U715 (N_715,N_188,N_170);
nand U716 (N_716,N_4,N_112);
or U717 (N_717,N_394,N_252);
nand U718 (N_718,N_101,N_52);
and U719 (N_719,N_286,N_21);
or U720 (N_720,N_220,N_198);
nor U721 (N_721,N_433,N_310);
nand U722 (N_722,N_273,N_354);
or U723 (N_723,N_382,N_381);
xnor U724 (N_724,N_302,N_64);
and U725 (N_725,N_479,N_243);
nand U726 (N_726,N_355,N_80);
or U727 (N_727,N_18,N_32);
and U728 (N_728,N_218,N_484);
or U729 (N_729,N_429,N_386);
or U730 (N_730,N_202,N_119);
nand U731 (N_731,N_110,N_34);
and U732 (N_732,N_123,N_287);
nand U733 (N_733,N_213,N_181);
nand U734 (N_734,N_228,N_296);
or U735 (N_735,N_106,N_487);
nor U736 (N_736,N_436,N_240);
nand U737 (N_737,N_353,N_217);
or U738 (N_738,N_485,N_366);
nor U739 (N_739,N_480,N_116);
xor U740 (N_740,N_16,N_393);
nor U741 (N_741,N_137,N_358);
and U742 (N_742,N_187,N_15);
or U743 (N_743,N_325,N_219);
nand U744 (N_744,N_414,N_40);
or U745 (N_745,N_14,N_159);
xor U746 (N_746,N_131,N_166);
nor U747 (N_747,N_69,N_23);
and U748 (N_748,N_211,N_438);
nand U749 (N_749,N_268,N_239);
or U750 (N_750,N_481,N_82);
nor U751 (N_751,N_358,N_240);
and U752 (N_752,N_465,N_99);
or U753 (N_753,N_454,N_427);
and U754 (N_754,N_206,N_348);
or U755 (N_755,N_274,N_469);
and U756 (N_756,N_18,N_363);
xnor U757 (N_757,N_271,N_287);
or U758 (N_758,N_285,N_311);
nor U759 (N_759,N_444,N_319);
or U760 (N_760,N_199,N_52);
or U761 (N_761,N_276,N_361);
nand U762 (N_762,N_309,N_227);
nand U763 (N_763,N_41,N_213);
nand U764 (N_764,N_64,N_55);
nand U765 (N_765,N_221,N_20);
xor U766 (N_766,N_235,N_315);
and U767 (N_767,N_452,N_10);
or U768 (N_768,N_168,N_220);
and U769 (N_769,N_172,N_335);
nand U770 (N_770,N_154,N_345);
xor U771 (N_771,N_212,N_27);
xnor U772 (N_772,N_405,N_411);
or U773 (N_773,N_132,N_335);
nor U774 (N_774,N_68,N_62);
nor U775 (N_775,N_128,N_295);
nor U776 (N_776,N_434,N_103);
or U777 (N_777,N_9,N_392);
xor U778 (N_778,N_81,N_75);
or U779 (N_779,N_365,N_157);
xnor U780 (N_780,N_375,N_287);
nor U781 (N_781,N_228,N_125);
nor U782 (N_782,N_131,N_194);
or U783 (N_783,N_344,N_193);
or U784 (N_784,N_463,N_148);
nor U785 (N_785,N_89,N_201);
nor U786 (N_786,N_171,N_204);
and U787 (N_787,N_391,N_313);
or U788 (N_788,N_288,N_381);
and U789 (N_789,N_415,N_493);
nand U790 (N_790,N_337,N_173);
nand U791 (N_791,N_251,N_136);
and U792 (N_792,N_5,N_73);
and U793 (N_793,N_355,N_359);
nor U794 (N_794,N_475,N_277);
and U795 (N_795,N_397,N_136);
or U796 (N_796,N_213,N_239);
or U797 (N_797,N_198,N_7);
or U798 (N_798,N_464,N_96);
or U799 (N_799,N_90,N_109);
or U800 (N_800,N_246,N_112);
or U801 (N_801,N_446,N_178);
nand U802 (N_802,N_303,N_177);
nand U803 (N_803,N_385,N_481);
nor U804 (N_804,N_88,N_105);
and U805 (N_805,N_67,N_236);
nor U806 (N_806,N_469,N_10);
nor U807 (N_807,N_191,N_155);
nor U808 (N_808,N_98,N_400);
and U809 (N_809,N_187,N_97);
nor U810 (N_810,N_27,N_234);
or U811 (N_811,N_124,N_153);
or U812 (N_812,N_361,N_201);
or U813 (N_813,N_256,N_211);
nor U814 (N_814,N_40,N_234);
nor U815 (N_815,N_8,N_476);
nand U816 (N_816,N_7,N_368);
nor U817 (N_817,N_140,N_105);
and U818 (N_818,N_146,N_114);
or U819 (N_819,N_486,N_246);
nand U820 (N_820,N_316,N_305);
nor U821 (N_821,N_445,N_289);
nand U822 (N_822,N_274,N_298);
and U823 (N_823,N_319,N_338);
and U824 (N_824,N_237,N_420);
nor U825 (N_825,N_306,N_450);
and U826 (N_826,N_427,N_135);
or U827 (N_827,N_8,N_144);
nand U828 (N_828,N_313,N_212);
nor U829 (N_829,N_292,N_61);
nor U830 (N_830,N_261,N_298);
nor U831 (N_831,N_298,N_468);
and U832 (N_832,N_221,N_336);
xnor U833 (N_833,N_116,N_217);
and U834 (N_834,N_48,N_423);
nor U835 (N_835,N_263,N_11);
and U836 (N_836,N_353,N_9);
nand U837 (N_837,N_297,N_67);
or U838 (N_838,N_33,N_282);
or U839 (N_839,N_480,N_86);
nand U840 (N_840,N_69,N_288);
xnor U841 (N_841,N_69,N_115);
or U842 (N_842,N_76,N_258);
nor U843 (N_843,N_365,N_413);
nor U844 (N_844,N_326,N_139);
nand U845 (N_845,N_142,N_126);
and U846 (N_846,N_101,N_192);
nand U847 (N_847,N_179,N_8);
nand U848 (N_848,N_433,N_165);
and U849 (N_849,N_143,N_36);
and U850 (N_850,N_268,N_489);
nor U851 (N_851,N_28,N_181);
and U852 (N_852,N_319,N_2);
nand U853 (N_853,N_466,N_164);
nand U854 (N_854,N_304,N_129);
and U855 (N_855,N_474,N_453);
nand U856 (N_856,N_274,N_426);
and U857 (N_857,N_56,N_286);
nor U858 (N_858,N_107,N_445);
xor U859 (N_859,N_164,N_307);
nand U860 (N_860,N_116,N_375);
nor U861 (N_861,N_396,N_365);
nor U862 (N_862,N_336,N_341);
nor U863 (N_863,N_182,N_290);
xnor U864 (N_864,N_316,N_274);
nor U865 (N_865,N_397,N_43);
nand U866 (N_866,N_63,N_150);
xor U867 (N_867,N_70,N_349);
or U868 (N_868,N_292,N_97);
nor U869 (N_869,N_106,N_19);
xnor U870 (N_870,N_431,N_212);
xor U871 (N_871,N_282,N_461);
xor U872 (N_872,N_146,N_402);
xnor U873 (N_873,N_69,N_199);
or U874 (N_874,N_223,N_414);
nand U875 (N_875,N_110,N_345);
nor U876 (N_876,N_135,N_208);
nor U877 (N_877,N_32,N_159);
and U878 (N_878,N_110,N_112);
xor U879 (N_879,N_28,N_376);
nand U880 (N_880,N_299,N_444);
or U881 (N_881,N_281,N_471);
or U882 (N_882,N_72,N_4);
or U883 (N_883,N_237,N_60);
nand U884 (N_884,N_174,N_37);
and U885 (N_885,N_455,N_364);
nand U886 (N_886,N_229,N_123);
or U887 (N_887,N_241,N_231);
nand U888 (N_888,N_363,N_427);
xor U889 (N_889,N_370,N_335);
nor U890 (N_890,N_113,N_85);
nor U891 (N_891,N_319,N_479);
nand U892 (N_892,N_353,N_83);
and U893 (N_893,N_56,N_256);
nand U894 (N_894,N_486,N_92);
and U895 (N_895,N_350,N_40);
nand U896 (N_896,N_329,N_348);
and U897 (N_897,N_173,N_193);
nand U898 (N_898,N_455,N_3);
xnor U899 (N_899,N_267,N_470);
and U900 (N_900,N_336,N_487);
and U901 (N_901,N_355,N_286);
xnor U902 (N_902,N_434,N_152);
or U903 (N_903,N_397,N_37);
and U904 (N_904,N_230,N_346);
nor U905 (N_905,N_495,N_274);
nand U906 (N_906,N_43,N_186);
or U907 (N_907,N_47,N_346);
nor U908 (N_908,N_497,N_363);
and U909 (N_909,N_46,N_437);
and U910 (N_910,N_200,N_254);
or U911 (N_911,N_177,N_457);
xor U912 (N_912,N_418,N_157);
nor U913 (N_913,N_377,N_204);
nand U914 (N_914,N_422,N_90);
or U915 (N_915,N_195,N_399);
nor U916 (N_916,N_374,N_26);
or U917 (N_917,N_205,N_401);
or U918 (N_918,N_142,N_362);
xor U919 (N_919,N_345,N_289);
nand U920 (N_920,N_77,N_325);
nand U921 (N_921,N_377,N_125);
or U922 (N_922,N_98,N_250);
or U923 (N_923,N_176,N_103);
and U924 (N_924,N_298,N_493);
and U925 (N_925,N_28,N_256);
xnor U926 (N_926,N_253,N_271);
xnor U927 (N_927,N_417,N_424);
and U928 (N_928,N_50,N_194);
nor U929 (N_929,N_111,N_216);
nand U930 (N_930,N_424,N_0);
xor U931 (N_931,N_346,N_449);
nand U932 (N_932,N_347,N_282);
xnor U933 (N_933,N_224,N_161);
nand U934 (N_934,N_2,N_86);
and U935 (N_935,N_487,N_115);
and U936 (N_936,N_256,N_209);
and U937 (N_937,N_195,N_294);
and U938 (N_938,N_373,N_449);
or U939 (N_939,N_448,N_300);
and U940 (N_940,N_451,N_316);
nand U941 (N_941,N_416,N_282);
and U942 (N_942,N_416,N_149);
nand U943 (N_943,N_191,N_210);
or U944 (N_944,N_356,N_422);
and U945 (N_945,N_99,N_497);
and U946 (N_946,N_140,N_108);
or U947 (N_947,N_86,N_476);
nor U948 (N_948,N_262,N_210);
xor U949 (N_949,N_53,N_220);
or U950 (N_950,N_361,N_280);
nand U951 (N_951,N_267,N_114);
xnor U952 (N_952,N_113,N_121);
and U953 (N_953,N_154,N_465);
and U954 (N_954,N_300,N_110);
nand U955 (N_955,N_28,N_111);
or U956 (N_956,N_326,N_24);
and U957 (N_957,N_367,N_251);
nor U958 (N_958,N_120,N_34);
or U959 (N_959,N_65,N_279);
nand U960 (N_960,N_187,N_469);
or U961 (N_961,N_125,N_288);
nand U962 (N_962,N_272,N_217);
and U963 (N_963,N_47,N_405);
nand U964 (N_964,N_68,N_390);
nor U965 (N_965,N_201,N_459);
nand U966 (N_966,N_350,N_247);
nand U967 (N_967,N_429,N_84);
or U968 (N_968,N_339,N_199);
xor U969 (N_969,N_296,N_414);
and U970 (N_970,N_174,N_227);
nor U971 (N_971,N_289,N_121);
nand U972 (N_972,N_132,N_490);
and U973 (N_973,N_378,N_114);
or U974 (N_974,N_158,N_374);
nor U975 (N_975,N_373,N_89);
or U976 (N_976,N_1,N_441);
xnor U977 (N_977,N_95,N_32);
xor U978 (N_978,N_175,N_286);
nor U979 (N_979,N_473,N_478);
or U980 (N_980,N_286,N_402);
and U981 (N_981,N_119,N_121);
and U982 (N_982,N_78,N_303);
xnor U983 (N_983,N_474,N_356);
xnor U984 (N_984,N_43,N_128);
and U985 (N_985,N_157,N_258);
or U986 (N_986,N_178,N_208);
and U987 (N_987,N_318,N_451);
and U988 (N_988,N_290,N_479);
nand U989 (N_989,N_256,N_422);
and U990 (N_990,N_103,N_184);
nand U991 (N_991,N_382,N_329);
nor U992 (N_992,N_409,N_499);
or U993 (N_993,N_388,N_10);
xnor U994 (N_994,N_1,N_286);
nand U995 (N_995,N_319,N_78);
nor U996 (N_996,N_103,N_427);
nor U997 (N_997,N_498,N_14);
and U998 (N_998,N_36,N_412);
xnor U999 (N_999,N_455,N_408);
or U1000 (N_1000,N_705,N_711);
or U1001 (N_1001,N_893,N_670);
nand U1002 (N_1002,N_708,N_923);
nor U1003 (N_1003,N_867,N_552);
nor U1004 (N_1004,N_803,N_807);
nor U1005 (N_1005,N_640,N_943);
or U1006 (N_1006,N_706,N_891);
nand U1007 (N_1007,N_641,N_997);
nand U1008 (N_1008,N_725,N_908);
and U1009 (N_1009,N_782,N_650);
nand U1010 (N_1010,N_609,N_700);
or U1011 (N_1011,N_579,N_666);
xnor U1012 (N_1012,N_516,N_993);
and U1013 (N_1013,N_956,N_871);
nand U1014 (N_1014,N_851,N_998);
or U1015 (N_1015,N_716,N_749);
nand U1016 (N_1016,N_944,N_904);
nand U1017 (N_1017,N_620,N_907);
nand U1018 (N_1018,N_755,N_726);
xnor U1019 (N_1019,N_506,N_878);
or U1020 (N_1020,N_563,N_933);
nor U1021 (N_1021,N_550,N_853);
and U1022 (N_1022,N_630,N_963);
xor U1023 (N_1023,N_996,N_827);
nand U1024 (N_1024,N_844,N_614);
nand U1025 (N_1025,N_929,N_764);
nor U1026 (N_1026,N_843,N_890);
and U1027 (N_1027,N_680,N_549);
or U1028 (N_1028,N_837,N_575);
and U1029 (N_1029,N_877,N_611);
nor U1030 (N_1030,N_814,N_570);
nor U1031 (N_1031,N_758,N_813);
nand U1032 (N_1032,N_791,N_790);
xnor U1033 (N_1033,N_863,N_538);
or U1034 (N_1034,N_903,N_581);
or U1035 (N_1035,N_615,N_584);
nor U1036 (N_1036,N_553,N_777);
nand U1037 (N_1037,N_905,N_687);
and U1038 (N_1038,N_509,N_539);
xnor U1039 (N_1039,N_828,N_528);
or U1040 (N_1040,N_534,N_564);
and U1041 (N_1041,N_602,N_595);
nor U1042 (N_1042,N_840,N_653);
and U1043 (N_1043,N_888,N_503);
or U1044 (N_1044,N_601,N_635);
nand U1045 (N_1045,N_838,N_899);
nor U1046 (N_1046,N_809,N_709);
and U1047 (N_1047,N_642,N_942);
and U1048 (N_1048,N_554,N_675);
nand U1049 (N_1049,N_874,N_722);
or U1050 (N_1050,N_808,N_622);
nor U1051 (N_1051,N_823,N_946);
xnor U1052 (N_1052,N_770,N_805);
xnor U1053 (N_1053,N_517,N_834);
or U1054 (N_1054,N_662,N_735);
nand U1055 (N_1055,N_589,N_574);
nand U1056 (N_1056,N_859,N_619);
nand U1057 (N_1057,N_717,N_772);
or U1058 (N_1058,N_961,N_846);
nor U1059 (N_1059,N_737,N_594);
and U1060 (N_1060,N_776,N_537);
or U1061 (N_1061,N_951,N_606);
nor U1062 (N_1062,N_625,N_804);
or U1063 (N_1063,N_991,N_992);
nor U1064 (N_1064,N_559,N_718);
or U1065 (N_1065,N_600,N_565);
and U1066 (N_1066,N_707,N_898);
nand U1067 (N_1067,N_748,N_751);
nand U1068 (N_1068,N_861,N_616);
nor U1069 (N_1069,N_817,N_521);
or U1070 (N_1070,N_924,N_762);
nand U1071 (N_1071,N_848,N_701);
and U1072 (N_1072,N_543,N_511);
nand U1073 (N_1073,N_637,N_518);
nor U1074 (N_1074,N_881,N_866);
or U1075 (N_1075,N_824,N_842);
xor U1076 (N_1076,N_730,N_679);
xnor U1077 (N_1077,N_761,N_832);
and U1078 (N_1078,N_750,N_608);
and U1079 (N_1079,N_887,N_788);
and U1080 (N_1080,N_533,N_994);
nand U1081 (N_1081,N_932,N_884);
nor U1082 (N_1082,N_970,N_671);
or U1083 (N_1083,N_958,N_535);
or U1084 (N_1084,N_959,N_703);
nor U1085 (N_1085,N_667,N_811);
nor U1086 (N_1086,N_693,N_794);
nand U1087 (N_1087,N_967,N_987);
and U1088 (N_1088,N_646,N_856);
nor U1089 (N_1089,N_775,N_855);
nand U1090 (N_1090,N_598,N_950);
nand U1091 (N_1091,N_826,N_919);
xnor U1092 (N_1092,N_681,N_806);
or U1093 (N_1093,N_800,N_973);
nand U1094 (N_1094,N_659,N_548);
or U1095 (N_1095,N_953,N_732);
or U1096 (N_1096,N_948,N_854);
nand U1097 (N_1097,N_918,N_572);
and U1098 (N_1098,N_603,N_763);
and U1099 (N_1099,N_911,N_519);
or U1100 (N_1100,N_873,N_986);
or U1101 (N_1101,N_765,N_927);
or U1102 (N_1102,N_779,N_741);
xor U1103 (N_1103,N_939,N_704);
and U1104 (N_1104,N_580,N_822);
or U1105 (N_1105,N_810,N_566);
nor U1106 (N_1106,N_930,N_885);
nand U1107 (N_1107,N_781,N_812);
nor U1108 (N_1108,N_985,N_829);
xor U1109 (N_1109,N_696,N_604);
and U1110 (N_1110,N_644,N_922);
and U1111 (N_1111,N_815,N_767);
nand U1112 (N_1112,N_510,N_720);
nand U1113 (N_1113,N_523,N_949);
nand U1114 (N_1114,N_545,N_597);
or U1115 (N_1115,N_917,N_870);
nand U1116 (N_1116,N_724,N_821);
and U1117 (N_1117,N_520,N_974);
nand U1118 (N_1118,N_547,N_652);
nand U1119 (N_1119,N_864,N_744);
nand U1120 (N_1120,N_561,N_968);
nand U1121 (N_1121,N_906,N_654);
nor U1122 (N_1122,N_660,N_979);
and U1123 (N_1123,N_629,N_995);
nor U1124 (N_1124,N_663,N_558);
and U1125 (N_1125,N_895,N_818);
and U1126 (N_1126,N_728,N_556);
nor U1127 (N_1127,N_698,N_965);
or U1128 (N_1128,N_583,N_976);
nor U1129 (N_1129,N_978,N_540);
or U1130 (N_1130,N_682,N_868);
and U1131 (N_1131,N_766,N_592);
nand U1132 (N_1132,N_971,N_684);
and U1133 (N_1133,N_689,N_771);
nand U1134 (N_1134,N_673,N_512);
or U1135 (N_1135,N_757,N_988);
nand U1136 (N_1136,N_957,N_880);
or U1137 (N_1137,N_714,N_505);
and U1138 (N_1138,N_555,N_731);
nand U1139 (N_1139,N_723,N_613);
and U1140 (N_1140,N_785,N_882);
xnor U1141 (N_1141,N_801,N_876);
nand U1142 (N_1142,N_835,N_799);
nor U1143 (N_1143,N_894,N_531);
nor U1144 (N_1144,N_819,N_754);
xnor U1145 (N_1145,N_648,N_530);
and U1146 (N_1146,N_590,N_909);
nor U1147 (N_1147,N_672,N_802);
xor U1148 (N_1148,N_743,N_872);
nand U1149 (N_1149,N_591,N_984);
nand U1150 (N_1150,N_627,N_669);
nand U1151 (N_1151,N_536,N_830);
nor U1152 (N_1152,N_685,N_862);
nand U1153 (N_1153,N_768,N_686);
nand U1154 (N_1154,N_710,N_839);
and U1155 (N_1155,N_634,N_831);
nand U1156 (N_1156,N_526,N_721);
nand U1157 (N_1157,N_975,N_977);
nand U1158 (N_1158,N_712,N_850);
or U1159 (N_1159,N_631,N_784);
nor U1160 (N_1160,N_941,N_610);
nor U1161 (N_1161,N_524,N_527);
or U1162 (N_1162,N_739,N_797);
and U1163 (N_1163,N_639,N_841);
or U1164 (N_1164,N_585,N_621);
or U1165 (N_1165,N_665,N_734);
nand U1166 (N_1166,N_656,N_982);
nand U1167 (N_1167,N_643,N_966);
nor U1168 (N_1168,N_715,N_542);
and U1169 (N_1169,N_912,N_668);
nand U1170 (N_1170,N_798,N_915);
nand U1171 (N_1171,N_921,N_578);
or U1172 (N_1172,N_945,N_981);
and U1173 (N_1173,N_658,N_789);
nand U1174 (N_1174,N_889,N_618);
or U1175 (N_1175,N_820,N_759);
or U1176 (N_1176,N_914,N_568);
and U1177 (N_1177,N_661,N_936);
xnor U1178 (N_1178,N_916,N_931);
nand U1179 (N_1179,N_733,N_736);
nand U1180 (N_1180,N_576,N_753);
nand U1181 (N_1181,N_514,N_857);
nor U1182 (N_1182,N_746,N_883);
or U1183 (N_1183,N_623,N_532);
and U1184 (N_1184,N_901,N_886);
nand U1185 (N_1185,N_964,N_617);
and U1186 (N_1186,N_586,N_677);
or U1187 (N_1187,N_962,N_729);
xnor U1188 (N_1188,N_502,N_980);
nor U1189 (N_1189,N_596,N_719);
and U1190 (N_1190,N_571,N_501);
nand U1191 (N_1191,N_865,N_825);
nand U1192 (N_1192,N_849,N_875);
and U1193 (N_1193,N_560,N_633);
or U1194 (N_1194,N_969,N_773);
nand U1195 (N_1195,N_508,N_683);
or U1196 (N_1196,N_507,N_938);
nor U1197 (N_1197,N_638,N_836);
nor U1198 (N_1198,N_740,N_624);
nand U1199 (N_1199,N_541,N_632);
nand U1200 (N_1200,N_816,N_910);
nand U1201 (N_1201,N_674,N_989);
and U1202 (N_1202,N_664,N_972);
or U1203 (N_1203,N_588,N_522);
nand U1204 (N_1204,N_504,N_599);
or U1205 (N_1205,N_902,N_934);
or U1206 (N_1206,N_960,N_896);
nand U1207 (N_1207,N_792,N_845);
and U1208 (N_1208,N_587,N_645);
or U1209 (N_1209,N_573,N_940);
nand U1210 (N_1210,N_702,N_699);
or U1211 (N_1211,N_852,N_795);
nand U1212 (N_1212,N_892,N_612);
nor U1213 (N_1213,N_691,N_879);
nor U1214 (N_1214,N_858,N_947);
or U1215 (N_1215,N_954,N_694);
nand U1216 (N_1216,N_551,N_778);
xnor U1217 (N_1217,N_688,N_593);
or U1218 (N_1218,N_607,N_513);
nand U1219 (N_1219,N_738,N_655);
nand U1220 (N_1220,N_695,N_567);
nand U1221 (N_1221,N_780,N_742);
nor U1222 (N_1222,N_605,N_582);
or U1223 (N_1223,N_529,N_937);
xor U1224 (N_1224,N_713,N_727);
or U1225 (N_1225,N_525,N_678);
or U1226 (N_1226,N_833,N_897);
nor U1227 (N_1227,N_926,N_747);
nor U1228 (N_1228,N_626,N_783);
nand U1229 (N_1229,N_544,N_628);
nand U1230 (N_1230,N_649,N_999);
and U1231 (N_1231,N_697,N_752);
nor U1232 (N_1232,N_692,N_500);
nand U1233 (N_1233,N_636,N_793);
or U1234 (N_1234,N_847,N_925);
nand U1235 (N_1235,N_952,N_769);
nand U1236 (N_1236,N_869,N_955);
and U1237 (N_1237,N_676,N_787);
nor U1238 (N_1238,N_546,N_935);
nand U1239 (N_1239,N_651,N_983);
nor U1240 (N_1240,N_990,N_928);
nand U1241 (N_1241,N_577,N_690);
nand U1242 (N_1242,N_860,N_900);
or U1243 (N_1243,N_569,N_786);
and U1244 (N_1244,N_657,N_557);
or U1245 (N_1245,N_913,N_562);
or U1246 (N_1246,N_774,N_647);
or U1247 (N_1247,N_756,N_745);
or U1248 (N_1248,N_796,N_760);
xnor U1249 (N_1249,N_920,N_515);
nand U1250 (N_1250,N_836,N_719);
nand U1251 (N_1251,N_951,N_524);
and U1252 (N_1252,N_924,N_778);
nor U1253 (N_1253,N_904,N_714);
nand U1254 (N_1254,N_993,N_714);
and U1255 (N_1255,N_851,N_857);
and U1256 (N_1256,N_649,N_789);
and U1257 (N_1257,N_886,N_643);
nand U1258 (N_1258,N_939,N_994);
and U1259 (N_1259,N_775,N_870);
or U1260 (N_1260,N_785,N_572);
and U1261 (N_1261,N_594,N_714);
and U1262 (N_1262,N_660,N_912);
or U1263 (N_1263,N_684,N_745);
xnor U1264 (N_1264,N_577,N_835);
nor U1265 (N_1265,N_710,N_824);
nand U1266 (N_1266,N_818,N_561);
and U1267 (N_1267,N_709,N_572);
nand U1268 (N_1268,N_810,N_827);
xor U1269 (N_1269,N_613,N_831);
nor U1270 (N_1270,N_654,N_983);
and U1271 (N_1271,N_888,N_758);
or U1272 (N_1272,N_904,N_635);
nand U1273 (N_1273,N_572,N_802);
and U1274 (N_1274,N_915,N_578);
nor U1275 (N_1275,N_505,N_881);
and U1276 (N_1276,N_828,N_840);
nand U1277 (N_1277,N_696,N_780);
and U1278 (N_1278,N_850,N_503);
nand U1279 (N_1279,N_614,N_557);
and U1280 (N_1280,N_689,N_868);
nor U1281 (N_1281,N_642,N_605);
nor U1282 (N_1282,N_520,N_713);
xor U1283 (N_1283,N_664,N_656);
or U1284 (N_1284,N_654,N_860);
or U1285 (N_1285,N_848,N_854);
and U1286 (N_1286,N_897,N_924);
and U1287 (N_1287,N_583,N_509);
nand U1288 (N_1288,N_726,N_576);
nand U1289 (N_1289,N_828,N_554);
or U1290 (N_1290,N_978,N_988);
nand U1291 (N_1291,N_579,N_635);
nor U1292 (N_1292,N_532,N_834);
and U1293 (N_1293,N_617,N_997);
and U1294 (N_1294,N_746,N_523);
or U1295 (N_1295,N_903,N_542);
nand U1296 (N_1296,N_702,N_716);
nor U1297 (N_1297,N_650,N_759);
nor U1298 (N_1298,N_892,N_533);
nor U1299 (N_1299,N_722,N_914);
nand U1300 (N_1300,N_636,N_844);
and U1301 (N_1301,N_613,N_643);
xor U1302 (N_1302,N_610,N_857);
xnor U1303 (N_1303,N_889,N_544);
nand U1304 (N_1304,N_841,N_627);
xor U1305 (N_1305,N_613,N_981);
and U1306 (N_1306,N_991,N_916);
nor U1307 (N_1307,N_958,N_646);
nor U1308 (N_1308,N_899,N_751);
nand U1309 (N_1309,N_649,N_976);
nand U1310 (N_1310,N_682,N_537);
nand U1311 (N_1311,N_576,N_503);
nand U1312 (N_1312,N_611,N_788);
nor U1313 (N_1313,N_656,N_653);
xnor U1314 (N_1314,N_605,N_993);
and U1315 (N_1315,N_698,N_811);
and U1316 (N_1316,N_511,N_969);
nor U1317 (N_1317,N_918,N_772);
nand U1318 (N_1318,N_579,N_934);
xnor U1319 (N_1319,N_594,N_699);
xnor U1320 (N_1320,N_512,N_909);
and U1321 (N_1321,N_691,N_562);
xor U1322 (N_1322,N_647,N_782);
xnor U1323 (N_1323,N_850,N_840);
xor U1324 (N_1324,N_771,N_973);
nor U1325 (N_1325,N_851,N_805);
nand U1326 (N_1326,N_726,N_793);
nor U1327 (N_1327,N_808,N_902);
and U1328 (N_1328,N_603,N_753);
nand U1329 (N_1329,N_849,N_888);
xnor U1330 (N_1330,N_997,N_959);
xnor U1331 (N_1331,N_932,N_603);
or U1332 (N_1332,N_580,N_884);
nor U1333 (N_1333,N_623,N_555);
nand U1334 (N_1334,N_702,N_794);
and U1335 (N_1335,N_876,N_851);
nor U1336 (N_1336,N_732,N_822);
xnor U1337 (N_1337,N_717,N_848);
and U1338 (N_1338,N_549,N_578);
xnor U1339 (N_1339,N_644,N_997);
or U1340 (N_1340,N_760,N_603);
nand U1341 (N_1341,N_591,N_749);
and U1342 (N_1342,N_747,N_748);
and U1343 (N_1343,N_798,N_639);
xor U1344 (N_1344,N_512,N_844);
nand U1345 (N_1345,N_719,N_969);
or U1346 (N_1346,N_913,N_510);
xor U1347 (N_1347,N_588,N_865);
nand U1348 (N_1348,N_904,N_683);
and U1349 (N_1349,N_612,N_520);
or U1350 (N_1350,N_863,N_612);
or U1351 (N_1351,N_580,N_720);
and U1352 (N_1352,N_743,N_852);
nand U1353 (N_1353,N_903,N_942);
nand U1354 (N_1354,N_696,N_608);
nand U1355 (N_1355,N_882,N_510);
nand U1356 (N_1356,N_723,N_849);
or U1357 (N_1357,N_786,N_883);
nand U1358 (N_1358,N_769,N_863);
or U1359 (N_1359,N_997,N_891);
or U1360 (N_1360,N_668,N_729);
nor U1361 (N_1361,N_718,N_580);
and U1362 (N_1362,N_988,N_591);
and U1363 (N_1363,N_817,N_989);
nand U1364 (N_1364,N_609,N_844);
nor U1365 (N_1365,N_927,N_602);
nand U1366 (N_1366,N_711,N_887);
xnor U1367 (N_1367,N_567,N_580);
nand U1368 (N_1368,N_562,N_616);
or U1369 (N_1369,N_653,N_740);
nor U1370 (N_1370,N_946,N_691);
nor U1371 (N_1371,N_979,N_890);
nand U1372 (N_1372,N_914,N_607);
or U1373 (N_1373,N_587,N_789);
nor U1374 (N_1374,N_934,N_529);
or U1375 (N_1375,N_826,N_948);
xnor U1376 (N_1376,N_974,N_711);
and U1377 (N_1377,N_627,N_993);
nand U1378 (N_1378,N_744,N_881);
and U1379 (N_1379,N_871,N_719);
or U1380 (N_1380,N_517,N_817);
nand U1381 (N_1381,N_640,N_808);
nand U1382 (N_1382,N_721,N_612);
and U1383 (N_1383,N_660,N_881);
nand U1384 (N_1384,N_688,N_667);
nor U1385 (N_1385,N_652,N_520);
and U1386 (N_1386,N_675,N_642);
nand U1387 (N_1387,N_849,N_971);
nand U1388 (N_1388,N_764,N_972);
nand U1389 (N_1389,N_800,N_732);
nand U1390 (N_1390,N_589,N_931);
or U1391 (N_1391,N_802,N_973);
nor U1392 (N_1392,N_796,N_979);
or U1393 (N_1393,N_690,N_837);
nand U1394 (N_1394,N_806,N_514);
xor U1395 (N_1395,N_757,N_637);
nor U1396 (N_1396,N_605,N_661);
xor U1397 (N_1397,N_975,N_803);
xor U1398 (N_1398,N_985,N_675);
nor U1399 (N_1399,N_555,N_974);
nand U1400 (N_1400,N_758,N_833);
and U1401 (N_1401,N_620,N_506);
nand U1402 (N_1402,N_831,N_669);
and U1403 (N_1403,N_545,N_548);
nor U1404 (N_1404,N_632,N_798);
nor U1405 (N_1405,N_821,N_541);
nand U1406 (N_1406,N_555,N_938);
or U1407 (N_1407,N_942,N_875);
xor U1408 (N_1408,N_840,N_753);
or U1409 (N_1409,N_537,N_548);
or U1410 (N_1410,N_647,N_601);
nand U1411 (N_1411,N_642,N_641);
and U1412 (N_1412,N_575,N_616);
and U1413 (N_1413,N_667,N_981);
xor U1414 (N_1414,N_539,N_892);
and U1415 (N_1415,N_540,N_981);
or U1416 (N_1416,N_637,N_585);
xor U1417 (N_1417,N_954,N_750);
nor U1418 (N_1418,N_811,N_994);
or U1419 (N_1419,N_829,N_675);
or U1420 (N_1420,N_749,N_722);
nand U1421 (N_1421,N_887,N_961);
or U1422 (N_1422,N_634,N_758);
xor U1423 (N_1423,N_812,N_591);
xor U1424 (N_1424,N_892,N_615);
nor U1425 (N_1425,N_631,N_850);
and U1426 (N_1426,N_569,N_933);
and U1427 (N_1427,N_785,N_821);
or U1428 (N_1428,N_522,N_708);
nand U1429 (N_1429,N_774,N_990);
nand U1430 (N_1430,N_619,N_976);
and U1431 (N_1431,N_949,N_901);
xor U1432 (N_1432,N_812,N_593);
or U1433 (N_1433,N_967,N_605);
xnor U1434 (N_1434,N_515,N_797);
nand U1435 (N_1435,N_578,N_832);
and U1436 (N_1436,N_543,N_681);
and U1437 (N_1437,N_865,N_616);
or U1438 (N_1438,N_550,N_564);
nor U1439 (N_1439,N_804,N_593);
nand U1440 (N_1440,N_813,N_661);
nor U1441 (N_1441,N_758,N_777);
or U1442 (N_1442,N_592,N_877);
or U1443 (N_1443,N_754,N_573);
nand U1444 (N_1444,N_709,N_873);
nor U1445 (N_1445,N_883,N_891);
and U1446 (N_1446,N_816,N_800);
xor U1447 (N_1447,N_914,N_744);
and U1448 (N_1448,N_657,N_608);
nand U1449 (N_1449,N_714,N_721);
nor U1450 (N_1450,N_541,N_505);
and U1451 (N_1451,N_792,N_749);
and U1452 (N_1452,N_630,N_971);
or U1453 (N_1453,N_663,N_780);
nand U1454 (N_1454,N_777,N_587);
nor U1455 (N_1455,N_624,N_720);
nor U1456 (N_1456,N_610,N_502);
and U1457 (N_1457,N_956,N_906);
or U1458 (N_1458,N_837,N_856);
and U1459 (N_1459,N_643,N_707);
nand U1460 (N_1460,N_852,N_545);
nor U1461 (N_1461,N_701,N_897);
nand U1462 (N_1462,N_795,N_537);
nor U1463 (N_1463,N_784,N_556);
or U1464 (N_1464,N_652,N_805);
and U1465 (N_1465,N_962,N_699);
nand U1466 (N_1466,N_631,N_862);
nor U1467 (N_1467,N_695,N_774);
or U1468 (N_1468,N_980,N_597);
nand U1469 (N_1469,N_968,N_865);
and U1470 (N_1470,N_904,N_913);
nor U1471 (N_1471,N_812,N_972);
or U1472 (N_1472,N_546,N_897);
and U1473 (N_1473,N_778,N_754);
xor U1474 (N_1474,N_553,N_531);
nand U1475 (N_1475,N_826,N_795);
xor U1476 (N_1476,N_876,N_850);
and U1477 (N_1477,N_668,N_577);
or U1478 (N_1478,N_758,N_800);
xor U1479 (N_1479,N_765,N_730);
or U1480 (N_1480,N_619,N_878);
nor U1481 (N_1481,N_833,N_770);
or U1482 (N_1482,N_702,N_737);
and U1483 (N_1483,N_559,N_860);
and U1484 (N_1484,N_875,N_950);
nor U1485 (N_1485,N_566,N_562);
or U1486 (N_1486,N_513,N_880);
nand U1487 (N_1487,N_797,N_571);
nor U1488 (N_1488,N_539,N_727);
or U1489 (N_1489,N_529,N_990);
xor U1490 (N_1490,N_507,N_643);
or U1491 (N_1491,N_991,N_960);
and U1492 (N_1492,N_981,N_747);
or U1493 (N_1493,N_827,N_727);
and U1494 (N_1494,N_908,N_747);
and U1495 (N_1495,N_682,N_539);
xnor U1496 (N_1496,N_846,N_795);
or U1497 (N_1497,N_852,N_711);
nand U1498 (N_1498,N_704,N_560);
nor U1499 (N_1499,N_721,N_601);
nor U1500 (N_1500,N_1452,N_1474);
nand U1501 (N_1501,N_1027,N_1206);
nand U1502 (N_1502,N_1127,N_1009);
nor U1503 (N_1503,N_1349,N_1337);
nor U1504 (N_1504,N_1016,N_1306);
and U1505 (N_1505,N_1222,N_1445);
nand U1506 (N_1506,N_1096,N_1250);
or U1507 (N_1507,N_1091,N_1185);
and U1508 (N_1508,N_1438,N_1266);
and U1509 (N_1509,N_1208,N_1302);
xor U1510 (N_1510,N_1140,N_1097);
xor U1511 (N_1511,N_1259,N_1161);
nand U1512 (N_1512,N_1478,N_1340);
and U1513 (N_1513,N_1135,N_1022);
and U1514 (N_1514,N_1467,N_1450);
and U1515 (N_1515,N_1119,N_1498);
or U1516 (N_1516,N_1444,N_1138);
nor U1517 (N_1517,N_1032,N_1430);
or U1518 (N_1518,N_1439,N_1348);
and U1519 (N_1519,N_1333,N_1178);
nor U1520 (N_1520,N_1133,N_1416);
or U1521 (N_1521,N_1335,N_1093);
or U1522 (N_1522,N_1492,N_1146);
and U1523 (N_1523,N_1134,N_1220);
nand U1524 (N_1524,N_1285,N_1273);
and U1525 (N_1525,N_1103,N_1088);
nand U1526 (N_1526,N_1372,N_1287);
nor U1527 (N_1527,N_1375,N_1304);
nand U1528 (N_1528,N_1079,N_1351);
nand U1529 (N_1529,N_1459,N_1320);
nor U1530 (N_1530,N_1321,N_1184);
and U1531 (N_1531,N_1111,N_1479);
or U1532 (N_1532,N_1343,N_1473);
xnor U1533 (N_1533,N_1046,N_1130);
and U1534 (N_1534,N_1204,N_1368);
and U1535 (N_1535,N_1188,N_1485);
nor U1536 (N_1536,N_1165,N_1412);
xnor U1537 (N_1537,N_1442,N_1052);
xnor U1538 (N_1538,N_1158,N_1242);
and U1539 (N_1539,N_1326,N_1150);
nor U1540 (N_1540,N_1049,N_1075);
or U1541 (N_1541,N_1202,N_1328);
or U1542 (N_1542,N_1132,N_1290);
nor U1543 (N_1543,N_1128,N_1053);
or U1544 (N_1544,N_1436,N_1047);
nand U1545 (N_1545,N_1275,N_1059);
nand U1546 (N_1546,N_1175,N_1262);
and U1547 (N_1547,N_1226,N_1025);
and U1548 (N_1548,N_1354,N_1167);
or U1549 (N_1549,N_1115,N_1031);
and U1550 (N_1550,N_1044,N_1318);
nand U1551 (N_1551,N_1409,N_1051);
nand U1552 (N_1552,N_1179,N_1296);
nand U1553 (N_1553,N_1055,N_1311);
or U1554 (N_1554,N_1033,N_1376);
or U1555 (N_1555,N_1154,N_1398);
nor U1556 (N_1556,N_1141,N_1035);
or U1557 (N_1557,N_1377,N_1163);
nor U1558 (N_1558,N_1392,N_1070);
and U1559 (N_1559,N_1370,N_1000);
nor U1560 (N_1560,N_1252,N_1301);
nor U1561 (N_1561,N_1050,N_1063);
xor U1562 (N_1562,N_1282,N_1147);
or U1563 (N_1563,N_1008,N_1114);
nor U1564 (N_1564,N_1235,N_1057);
nand U1565 (N_1565,N_1257,N_1089);
nand U1566 (N_1566,N_1181,N_1383);
or U1567 (N_1567,N_1494,N_1207);
nand U1568 (N_1568,N_1477,N_1102);
or U1569 (N_1569,N_1469,N_1245);
and U1570 (N_1570,N_1329,N_1196);
and U1571 (N_1571,N_1325,N_1356);
xnor U1572 (N_1572,N_1232,N_1085);
nand U1573 (N_1573,N_1497,N_1263);
or U1574 (N_1574,N_1447,N_1371);
or U1575 (N_1575,N_1148,N_1194);
or U1576 (N_1576,N_1094,N_1172);
or U1577 (N_1577,N_1253,N_1122);
or U1578 (N_1578,N_1239,N_1421);
nand U1579 (N_1579,N_1401,N_1240);
nand U1580 (N_1580,N_1193,N_1411);
nand U1581 (N_1581,N_1312,N_1396);
xor U1582 (N_1582,N_1405,N_1344);
or U1583 (N_1583,N_1123,N_1422);
nand U1584 (N_1584,N_1299,N_1431);
and U1585 (N_1585,N_1261,N_1092);
nor U1586 (N_1586,N_1247,N_1381);
nand U1587 (N_1587,N_1455,N_1309);
and U1588 (N_1588,N_1030,N_1241);
xnor U1589 (N_1589,N_1342,N_1205);
nand U1590 (N_1590,N_1036,N_1365);
and U1591 (N_1591,N_1182,N_1308);
xnor U1592 (N_1592,N_1234,N_1034);
nand U1593 (N_1593,N_1280,N_1151);
nand U1594 (N_1594,N_1330,N_1180);
nand U1595 (N_1595,N_1095,N_1433);
nor U1596 (N_1596,N_1437,N_1106);
or U1597 (N_1597,N_1153,N_1112);
nor U1598 (N_1598,N_1471,N_1272);
nand U1599 (N_1599,N_1426,N_1144);
or U1600 (N_1600,N_1037,N_1389);
or U1601 (N_1601,N_1108,N_1026);
nor U1602 (N_1602,N_1197,N_1267);
or U1603 (N_1603,N_1137,N_1491);
and U1604 (N_1604,N_1129,N_1006);
and U1605 (N_1605,N_1440,N_1171);
and U1606 (N_1606,N_1294,N_1131);
nor U1607 (N_1607,N_1012,N_1260);
and U1608 (N_1608,N_1004,N_1039);
or U1609 (N_1609,N_1042,N_1427);
nor U1610 (N_1610,N_1105,N_1269);
nor U1611 (N_1611,N_1279,N_1305);
and U1612 (N_1612,N_1217,N_1200);
xor U1613 (N_1613,N_1230,N_1189);
and U1614 (N_1614,N_1339,N_1300);
nor U1615 (N_1615,N_1120,N_1186);
nand U1616 (N_1616,N_1005,N_1434);
nand U1617 (N_1617,N_1484,N_1454);
xnor U1618 (N_1618,N_1002,N_1238);
and U1619 (N_1619,N_1191,N_1314);
or U1620 (N_1620,N_1083,N_1216);
and U1621 (N_1621,N_1456,N_1378);
and U1622 (N_1622,N_1136,N_1227);
nand U1623 (N_1623,N_1319,N_1215);
or U1624 (N_1624,N_1203,N_1315);
nand U1625 (N_1625,N_1090,N_1283);
or U1626 (N_1626,N_1387,N_1080);
nand U1627 (N_1627,N_1391,N_1493);
or U1628 (N_1628,N_1323,N_1366);
nand U1629 (N_1629,N_1104,N_1110);
and U1630 (N_1630,N_1362,N_1380);
and U1631 (N_1631,N_1472,N_1461);
nand U1632 (N_1632,N_1345,N_1394);
nand U1633 (N_1633,N_1270,N_1069);
and U1634 (N_1634,N_1060,N_1384);
and U1635 (N_1635,N_1192,N_1099);
or U1636 (N_1636,N_1310,N_1143);
or U1637 (N_1637,N_1156,N_1303);
or U1638 (N_1638,N_1397,N_1201);
or U1639 (N_1639,N_1385,N_1449);
and U1640 (N_1640,N_1417,N_1152);
nand U1641 (N_1641,N_1068,N_1116);
or U1642 (N_1642,N_1019,N_1237);
nand U1643 (N_1643,N_1243,N_1198);
or U1644 (N_1644,N_1255,N_1404);
and U1645 (N_1645,N_1233,N_1334);
xor U1646 (N_1646,N_1281,N_1011);
nor U1647 (N_1647,N_1298,N_1064);
and U1648 (N_1648,N_1107,N_1221);
or U1649 (N_1649,N_1187,N_1499);
and U1650 (N_1650,N_1425,N_1407);
and U1651 (N_1651,N_1462,N_1061);
xor U1652 (N_1652,N_1468,N_1288);
or U1653 (N_1653,N_1278,N_1212);
and U1654 (N_1654,N_1256,N_1210);
or U1655 (N_1655,N_1361,N_1457);
and U1656 (N_1656,N_1023,N_1223);
nand U1657 (N_1657,N_1078,N_1015);
and U1658 (N_1658,N_1382,N_1169);
nand U1659 (N_1659,N_1084,N_1251);
or U1660 (N_1660,N_1065,N_1109);
nor U1661 (N_1661,N_1160,N_1359);
nand U1662 (N_1662,N_1423,N_1458);
or U1663 (N_1663,N_1347,N_1355);
nor U1664 (N_1664,N_1495,N_1415);
and U1665 (N_1665,N_1028,N_1066);
or U1666 (N_1666,N_1482,N_1435);
or U1667 (N_1667,N_1490,N_1475);
or U1668 (N_1668,N_1003,N_1463);
nor U1669 (N_1669,N_1327,N_1373);
or U1670 (N_1670,N_1341,N_1045);
nand U1671 (N_1671,N_1464,N_1386);
nor U1672 (N_1672,N_1211,N_1350);
and U1673 (N_1673,N_1038,N_1418);
and U1674 (N_1674,N_1199,N_1419);
and U1675 (N_1675,N_1214,N_1018);
nand U1676 (N_1676,N_1331,N_1324);
nand U1677 (N_1677,N_1056,N_1379);
nor U1678 (N_1678,N_1174,N_1124);
xnor U1679 (N_1679,N_1284,N_1399);
and U1680 (N_1680,N_1402,N_1408);
nand U1681 (N_1681,N_1480,N_1393);
or U1682 (N_1682,N_1390,N_1024);
or U1683 (N_1683,N_1013,N_1388);
xnor U1684 (N_1684,N_1077,N_1353);
nand U1685 (N_1685,N_1367,N_1338);
nor U1686 (N_1686,N_1357,N_1277);
nor U1687 (N_1687,N_1071,N_1168);
nor U1688 (N_1688,N_1358,N_1432);
nand U1689 (N_1689,N_1183,N_1265);
nand U1690 (N_1690,N_1336,N_1307);
and U1691 (N_1691,N_1224,N_1040);
nand U1692 (N_1692,N_1007,N_1489);
nor U1693 (N_1693,N_1414,N_1465);
nor U1694 (N_1694,N_1228,N_1086);
nor U1695 (N_1695,N_1476,N_1313);
or U1696 (N_1696,N_1451,N_1062);
nand U1697 (N_1697,N_1406,N_1352);
or U1698 (N_1698,N_1317,N_1496);
nand U1699 (N_1699,N_1369,N_1446);
or U1700 (N_1700,N_1121,N_1021);
and U1701 (N_1701,N_1048,N_1460);
xor U1702 (N_1702,N_1149,N_1441);
and U1703 (N_1703,N_1001,N_1043);
xor U1704 (N_1704,N_1072,N_1316);
or U1705 (N_1705,N_1213,N_1248);
and U1706 (N_1706,N_1470,N_1395);
xnor U1707 (N_1707,N_1264,N_1483);
or U1708 (N_1708,N_1249,N_1413);
or U1709 (N_1709,N_1410,N_1117);
nor U1710 (N_1710,N_1145,N_1297);
or U1711 (N_1711,N_1488,N_1443);
nand U1712 (N_1712,N_1157,N_1139);
and U1713 (N_1713,N_1020,N_1100);
nand U1714 (N_1714,N_1428,N_1058);
nor U1715 (N_1715,N_1177,N_1164);
or U1716 (N_1716,N_1014,N_1101);
and U1717 (N_1717,N_1292,N_1429);
nand U1718 (N_1718,N_1448,N_1170);
nand U1719 (N_1719,N_1173,N_1486);
nand U1720 (N_1720,N_1403,N_1159);
and U1721 (N_1721,N_1081,N_1400);
nand U1722 (N_1722,N_1087,N_1274);
and U1723 (N_1723,N_1125,N_1360);
or U1724 (N_1724,N_1225,N_1074);
nor U1725 (N_1725,N_1346,N_1082);
nand U1726 (N_1726,N_1209,N_1363);
and U1727 (N_1727,N_1322,N_1176);
or U1728 (N_1728,N_1118,N_1289);
or U1729 (N_1729,N_1113,N_1286);
nor U1730 (N_1730,N_1487,N_1017);
nor U1731 (N_1731,N_1246,N_1466);
and U1732 (N_1732,N_1166,N_1293);
or U1733 (N_1733,N_1010,N_1236);
xor U1734 (N_1734,N_1364,N_1041);
or U1735 (N_1735,N_1076,N_1054);
nand U1736 (N_1736,N_1276,N_1126);
nor U1737 (N_1737,N_1424,N_1332);
nand U1738 (N_1738,N_1190,N_1218);
and U1739 (N_1739,N_1142,N_1229);
and U1740 (N_1740,N_1073,N_1374);
nor U1741 (N_1741,N_1067,N_1258);
nand U1742 (N_1742,N_1420,N_1268);
xnor U1743 (N_1743,N_1029,N_1244);
xor U1744 (N_1744,N_1098,N_1155);
or U1745 (N_1745,N_1162,N_1291);
and U1746 (N_1746,N_1271,N_1231);
nand U1747 (N_1747,N_1481,N_1295);
nand U1748 (N_1748,N_1453,N_1254);
and U1749 (N_1749,N_1219,N_1195);
xnor U1750 (N_1750,N_1000,N_1031);
nand U1751 (N_1751,N_1271,N_1027);
xnor U1752 (N_1752,N_1091,N_1404);
nor U1753 (N_1753,N_1177,N_1027);
nor U1754 (N_1754,N_1170,N_1428);
nand U1755 (N_1755,N_1096,N_1353);
nand U1756 (N_1756,N_1044,N_1301);
or U1757 (N_1757,N_1020,N_1389);
and U1758 (N_1758,N_1101,N_1279);
and U1759 (N_1759,N_1248,N_1102);
nand U1760 (N_1760,N_1352,N_1362);
nand U1761 (N_1761,N_1334,N_1237);
and U1762 (N_1762,N_1205,N_1094);
or U1763 (N_1763,N_1096,N_1494);
nand U1764 (N_1764,N_1150,N_1434);
and U1765 (N_1765,N_1153,N_1009);
nand U1766 (N_1766,N_1156,N_1205);
nand U1767 (N_1767,N_1004,N_1107);
nand U1768 (N_1768,N_1362,N_1079);
and U1769 (N_1769,N_1495,N_1180);
nand U1770 (N_1770,N_1425,N_1246);
nor U1771 (N_1771,N_1247,N_1360);
or U1772 (N_1772,N_1370,N_1081);
xor U1773 (N_1773,N_1190,N_1373);
nor U1774 (N_1774,N_1334,N_1050);
nand U1775 (N_1775,N_1298,N_1296);
nor U1776 (N_1776,N_1199,N_1229);
and U1777 (N_1777,N_1099,N_1316);
nand U1778 (N_1778,N_1232,N_1211);
nand U1779 (N_1779,N_1071,N_1371);
or U1780 (N_1780,N_1083,N_1041);
or U1781 (N_1781,N_1126,N_1184);
nand U1782 (N_1782,N_1429,N_1275);
xor U1783 (N_1783,N_1039,N_1186);
or U1784 (N_1784,N_1119,N_1397);
or U1785 (N_1785,N_1149,N_1446);
or U1786 (N_1786,N_1317,N_1499);
nand U1787 (N_1787,N_1136,N_1443);
and U1788 (N_1788,N_1106,N_1187);
or U1789 (N_1789,N_1059,N_1202);
nand U1790 (N_1790,N_1295,N_1267);
xor U1791 (N_1791,N_1045,N_1411);
and U1792 (N_1792,N_1300,N_1375);
and U1793 (N_1793,N_1094,N_1448);
or U1794 (N_1794,N_1375,N_1484);
and U1795 (N_1795,N_1025,N_1393);
nand U1796 (N_1796,N_1212,N_1343);
and U1797 (N_1797,N_1418,N_1236);
nand U1798 (N_1798,N_1444,N_1238);
or U1799 (N_1799,N_1443,N_1217);
or U1800 (N_1800,N_1455,N_1025);
nor U1801 (N_1801,N_1113,N_1045);
nand U1802 (N_1802,N_1067,N_1056);
nor U1803 (N_1803,N_1421,N_1448);
nand U1804 (N_1804,N_1060,N_1445);
and U1805 (N_1805,N_1023,N_1469);
or U1806 (N_1806,N_1175,N_1239);
and U1807 (N_1807,N_1404,N_1221);
nor U1808 (N_1808,N_1058,N_1051);
nand U1809 (N_1809,N_1125,N_1396);
nor U1810 (N_1810,N_1240,N_1367);
nor U1811 (N_1811,N_1201,N_1011);
and U1812 (N_1812,N_1019,N_1399);
xor U1813 (N_1813,N_1018,N_1324);
nand U1814 (N_1814,N_1118,N_1392);
and U1815 (N_1815,N_1262,N_1088);
nor U1816 (N_1816,N_1132,N_1472);
nand U1817 (N_1817,N_1078,N_1112);
nand U1818 (N_1818,N_1199,N_1233);
nand U1819 (N_1819,N_1339,N_1469);
or U1820 (N_1820,N_1375,N_1356);
or U1821 (N_1821,N_1014,N_1030);
and U1822 (N_1822,N_1032,N_1061);
or U1823 (N_1823,N_1495,N_1399);
xnor U1824 (N_1824,N_1056,N_1098);
nand U1825 (N_1825,N_1303,N_1310);
nand U1826 (N_1826,N_1105,N_1444);
nand U1827 (N_1827,N_1087,N_1102);
or U1828 (N_1828,N_1311,N_1432);
nor U1829 (N_1829,N_1212,N_1431);
or U1830 (N_1830,N_1468,N_1301);
nand U1831 (N_1831,N_1192,N_1276);
and U1832 (N_1832,N_1183,N_1048);
nor U1833 (N_1833,N_1488,N_1156);
and U1834 (N_1834,N_1349,N_1314);
or U1835 (N_1835,N_1320,N_1366);
nor U1836 (N_1836,N_1166,N_1162);
or U1837 (N_1837,N_1206,N_1307);
or U1838 (N_1838,N_1415,N_1323);
and U1839 (N_1839,N_1379,N_1489);
nand U1840 (N_1840,N_1070,N_1378);
and U1841 (N_1841,N_1422,N_1006);
or U1842 (N_1842,N_1449,N_1063);
nand U1843 (N_1843,N_1081,N_1340);
or U1844 (N_1844,N_1040,N_1342);
and U1845 (N_1845,N_1127,N_1424);
or U1846 (N_1846,N_1298,N_1069);
and U1847 (N_1847,N_1079,N_1284);
or U1848 (N_1848,N_1209,N_1295);
xnor U1849 (N_1849,N_1320,N_1298);
and U1850 (N_1850,N_1214,N_1140);
nand U1851 (N_1851,N_1049,N_1114);
or U1852 (N_1852,N_1017,N_1425);
and U1853 (N_1853,N_1082,N_1396);
nand U1854 (N_1854,N_1272,N_1304);
nor U1855 (N_1855,N_1177,N_1041);
or U1856 (N_1856,N_1397,N_1012);
and U1857 (N_1857,N_1283,N_1352);
nor U1858 (N_1858,N_1029,N_1237);
and U1859 (N_1859,N_1294,N_1428);
nand U1860 (N_1860,N_1301,N_1480);
nand U1861 (N_1861,N_1272,N_1163);
and U1862 (N_1862,N_1018,N_1375);
or U1863 (N_1863,N_1277,N_1336);
or U1864 (N_1864,N_1012,N_1422);
nand U1865 (N_1865,N_1358,N_1109);
and U1866 (N_1866,N_1195,N_1229);
and U1867 (N_1867,N_1254,N_1127);
nor U1868 (N_1868,N_1324,N_1147);
nand U1869 (N_1869,N_1255,N_1239);
and U1870 (N_1870,N_1184,N_1380);
and U1871 (N_1871,N_1218,N_1461);
nor U1872 (N_1872,N_1462,N_1392);
nor U1873 (N_1873,N_1467,N_1087);
xor U1874 (N_1874,N_1054,N_1432);
and U1875 (N_1875,N_1021,N_1056);
or U1876 (N_1876,N_1472,N_1023);
nand U1877 (N_1877,N_1053,N_1077);
nand U1878 (N_1878,N_1003,N_1181);
xnor U1879 (N_1879,N_1013,N_1036);
or U1880 (N_1880,N_1333,N_1472);
and U1881 (N_1881,N_1064,N_1228);
nor U1882 (N_1882,N_1183,N_1282);
nor U1883 (N_1883,N_1243,N_1313);
nand U1884 (N_1884,N_1406,N_1431);
and U1885 (N_1885,N_1320,N_1423);
xor U1886 (N_1886,N_1106,N_1237);
or U1887 (N_1887,N_1078,N_1074);
and U1888 (N_1888,N_1130,N_1267);
nor U1889 (N_1889,N_1432,N_1388);
and U1890 (N_1890,N_1271,N_1280);
or U1891 (N_1891,N_1381,N_1073);
nor U1892 (N_1892,N_1321,N_1422);
nor U1893 (N_1893,N_1215,N_1492);
nand U1894 (N_1894,N_1259,N_1214);
nand U1895 (N_1895,N_1092,N_1252);
xnor U1896 (N_1896,N_1389,N_1301);
or U1897 (N_1897,N_1043,N_1183);
nand U1898 (N_1898,N_1288,N_1408);
nor U1899 (N_1899,N_1428,N_1163);
nand U1900 (N_1900,N_1011,N_1217);
and U1901 (N_1901,N_1289,N_1313);
and U1902 (N_1902,N_1198,N_1285);
and U1903 (N_1903,N_1272,N_1442);
nor U1904 (N_1904,N_1309,N_1439);
xor U1905 (N_1905,N_1180,N_1130);
nor U1906 (N_1906,N_1446,N_1184);
nand U1907 (N_1907,N_1439,N_1110);
xnor U1908 (N_1908,N_1071,N_1073);
nor U1909 (N_1909,N_1495,N_1367);
nor U1910 (N_1910,N_1160,N_1283);
nor U1911 (N_1911,N_1110,N_1404);
or U1912 (N_1912,N_1234,N_1121);
and U1913 (N_1913,N_1405,N_1156);
nand U1914 (N_1914,N_1041,N_1118);
nor U1915 (N_1915,N_1412,N_1456);
or U1916 (N_1916,N_1108,N_1458);
or U1917 (N_1917,N_1165,N_1439);
nand U1918 (N_1918,N_1149,N_1063);
xnor U1919 (N_1919,N_1023,N_1139);
and U1920 (N_1920,N_1355,N_1458);
and U1921 (N_1921,N_1209,N_1211);
nand U1922 (N_1922,N_1080,N_1484);
and U1923 (N_1923,N_1498,N_1166);
nand U1924 (N_1924,N_1152,N_1356);
nor U1925 (N_1925,N_1268,N_1314);
and U1926 (N_1926,N_1003,N_1063);
nand U1927 (N_1927,N_1381,N_1262);
and U1928 (N_1928,N_1206,N_1061);
and U1929 (N_1929,N_1109,N_1048);
xnor U1930 (N_1930,N_1253,N_1326);
or U1931 (N_1931,N_1238,N_1017);
nand U1932 (N_1932,N_1042,N_1073);
xnor U1933 (N_1933,N_1466,N_1294);
and U1934 (N_1934,N_1067,N_1134);
nor U1935 (N_1935,N_1190,N_1019);
nand U1936 (N_1936,N_1288,N_1435);
nand U1937 (N_1937,N_1018,N_1013);
or U1938 (N_1938,N_1242,N_1087);
nor U1939 (N_1939,N_1093,N_1485);
nand U1940 (N_1940,N_1081,N_1486);
nor U1941 (N_1941,N_1132,N_1222);
or U1942 (N_1942,N_1204,N_1490);
and U1943 (N_1943,N_1202,N_1045);
xor U1944 (N_1944,N_1494,N_1309);
and U1945 (N_1945,N_1480,N_1134);
and U1946 (N_1946,N_1492,N_1247);
or U1947 (N_1947,N_1228,N_1084);
and U1948 (N_1948,N_1371,N_1340);
and U1949 (N_1949,N_1419,N_1180);
and U1950 (N_1950,N_1073,N_1330);
nor U1951 (N_1951,N_1159,N_1232);
or U1952 (N_1952,N_1491,N_1376);
nand U1953 (N_1953,N_1292,N_1021);
or U1954 (N_1954,N_1427,N_1446);
xor U1955 (N_1955,N_1490,N_1299);
or U1956 (N_1956,N_1396,N_1280);
nor U1957 (N_1957,N_1231,N_1193);
nand U1958 (N_1958,N_1364,N_1137);
and U1959 (N_1959,N_1011,N_1381);
nor U1960 (N_1960,N_1356,N_1039);
nand U1961 (N_1961,N_1160,N_1300);
nor U1962 (N_1962,N_1110,N_1351);
nand U1963 (N_1963,N_1022,N_1112);
nand U1964 (N_1964,N_1006,N_1324);
nor U1965 (N_1965,N_1230,N_1043);
and U1966 (N_1966,N_1448,N_1278);
nor U1967 (N_1967,N_1221,N_1213);
nor U1968 (N_1968,N_1084,N_1359);
nand U1969 (N_1969,N_1225,N_1135);
xor U1970 (N_1970,N_1260,N_1296);
nand U1971 (N_1971,N_1133,N_1128);
or U1972 (N_1972,N_1352,N_1252);
nand U1973 (N_1973,N_1200,N_1384);
and U1974 (N_1974,N_1076,N_1117);
nor U1975 (N_1975,N_1118,N_1370);
or U1976 (N_1976,N_1102,N_1435);
nor U1977 (N_1977,N_1054,N_1279);
nor U1978 (N_1978,N_1310,N_1429);
nor U1979 (N_1979,N_1062,N_1145);
nand U1980 (N_1980,N_1490,N_1184);
nand U1981 (N_1981,N_1252,N_1074);
or U1982 (N_1982,N_1357,N_1035);
nand U1983 (N_1983,N_1104,N_1226);
and U1984 (N_1984,N_1321,N_1325);
nor U1985 (N_1985,N_1330,N_1367);
nor U1986 (N_1986,N_1460,N_1027);
nand U1987 (N_1987,N_1119,N_1311);
nand U1988 (N_1988,N_1185,N_1120);
nor U1989 (N_1989,N_1479,N_1075);
nor U1990 (N_1990,N_1363,N_1110);
nand U1991 (N_1991,N_1470,N_1022);
nand U1992 (N_1992,N_1159,N_1329);
and U1993 (N_1993,N_1381,N_1082);
nand U1994 (N_1994,N_1339,N_1457);
nand U1995 (N_1995,N_1392,N_1206);
nor U1996 (N_1996,N_1192,N_1038);
and U1997 (N_1997,N_1420,N_1480);
nor U1998 (N_1998,N_1250,N_1123);
nand U1999 (N_1999,N_1236,N_1129);
or U2000 (N_2000,N_1779,N_1870);
nand U2001 (N_2001,N_1880,N_1532);
or U2002 (N_2002,N_1616,N_1900);
nand U2003 (N_2003,N_1704,N_1890);
xor U2004 (N_2004,N_1978,N_1654);
nand U2005 (N_2005,N_1936,N_1850);
nor U2006 (N_2006,N_1662,N_1722);
or U2007 (N_2007,N_1904,N_1950);
nor U2008 (N_2008,N_1726,N_1983);
and U2009 (N_2009,N_1677,N_1928);
or U2010 (N_2010,N_1619,N_1982);
nand U2011 (N_2011,N_1559,N_1699);
nor U2012 (N_2012,N_1860,N_1872);
and U2013 (N_2013,N_1888,N_1683);
nand U2014 (N_2014,N_1750,N_1570);
nor U2015 (N_2015,N_1745,N_1641);
nand U2016 (N_2016,N_1709,N_1684);
or U2017 (N_2017,N_1583,N_1899);
and U2018 (N_2018,N_1985,N_1560);
nand U2019 (N_2019,N_1988,N_1887);
nor U2020 (N_2020,N_1925,N_1572);
and U2021 (N_2021,N_1891,N_1770);
nor U2022 (N_2022,N_1731,N_1550);
nand U2023 (N_2023,N_1640,N_1895);
or U2024 (N_2024,N_1916,N_1785);
or U2025 (N_2025,N_1674,N_1819);
nor U2026 (N_2026,N_1531,N_1682);
and U2027 (N_2027,N_1755,N_1869);
nor U2028 (N_2028,N_1644,N_1506);
nand U2029 (N_2029,N_1805,N_1664);
nand U2030 (N_2030,N_1517,N_1569);
or U2031 (N_2031,N_1837,N_1871);
nand U2032 (N_2032,N_1565,N_1702);
nand U2033 (N_2033,N_1839,N_1760);
and U2034 (N_2034,N_1799,N_1528);
nor U2035 (N_2035,N_1821,N_1715);
nor U2036 (N_2036,N_1545,N_1539);
and U2037 (N_2037,N_1812,N_1947);
nor U2038 (N_2038,N_1894,N_1633);
nor U2039 (N_2039,N_1929,N_1523);
or U2040 (N_2040,N_1769,N_1576);
nor U2041 (N_2041,N_1803,N_1518);
and U2042 (N_2042,N_1579,N_1575);
xor U2043 (N_2043,N_1730,N_1954);
xor U2044 (N_2044,N_1910,N_1938);
nor U2045 (N_2045,N_1658,N_1566);
nor U2046 (N_2046,N_1629,N_1663);
nand U2047 (N_2047,N_1774,N_1670);
and U2048 (N_2048,N_1949,N_1798);
nand U2049 (N_2049,N_1614,N_1541);
and U2050 (N_2050,N_1708,N_1653);
xor U2051 (N_2051,N_1697,N_1995);
xnor U2052 (N_2052,N_1747,N_1961);
or U2053 (N_2053,N_1649,N_1622);
xnor U2054 (N_2054,N_1739,N_1844);
xor U2055 (N_2055,N_1573,N_1940);
and U2056 (N_2056,N_1829,N_1973);
or U2057 (N_2057,N_1813,N_1868);
nor U2058 (N_2058,N_1848,N_1889);
nor U2059 (N_2059,N_1794,N_1881);
or U2060 (N_2060,N_1571,N_1934);
nand U2061 (N_2061,N_1533,N_1855);
nand U2062 (N_2062,N_1771,N_1919);
and U2063 (N_2063,N_1582,N_1909);
nand U2064 (N_2064,N_1707,N_1632);
and U2065 (N_2065,N_1841,N_1698);
or U2066 (N_2066,N_1943,N_1931);
nor U2067 (N_2067,N_1529,N_1547);
and U2068 (N_2068,N_1652,N_1519);
or U2069 (N_2069,N_1647,N_1555);
or U2070 (N_2070,N_1775,N_1937);
or U2071 (N_2071,N_1977,N_1723);
or U2072 (N_2072,N_1657,N_1721);
and U2073 (N_2073,N_1828,N_1751);
nand U2074 (N_2074,N_1503,N_1830);
nand U2075 (N_2075,N_1673,N_1941);
and U2076 (N_2076,N_1896,N_1603);
and U2077 (N_2077,N_1692,N_1907);
xnor U2078 (N_2078,N_1752,N_1686);
nand U2079 (N_2079,N_1924,N_1970);
and U2080 (N_2080,N_1962,N_1561);
or U2081 (N_2081,N_1676,N_1763);
xor U2082 (N_2082,N_1776,N_1668);
and U2083 (N_2083,N_1861,N_1557);
nand U2084 (N_2084,N_1631,N_1958);
nor U2085 (N_2085,N_1526,N_1567);
and U2086 (N_2086,N_1953,N_1678);
or U2087 (N_2087,N_1999,N_1511);
nor U2088 (N_2088,N_1994,N_1795);
nand U2089 (N_2089,N_1691,N_1955);
nand U2090 (N_2090,N_1585,N_1643);
and U2091 (N_2091,N_1717,N_1637);
or U2092 (N_2092,N_1784,N_1908);
nand U2093 (N_2093,N_1917,N_1987);
nand U2094 (N_2094,N_1898,N_1639);
or U2095 (N_2095,N_1588,N_1846);
and U2096 (N_2096,N_1690,N_1984);
and U2097 (N_2097,N_1744,N_1608);
nand U2098 (N_2098,N_1742,N_1661);
or U2099 (N_2099,N_1617,N_1666);
and U2100 (N_2100,N_1500,N_1655);
nand U2101 (N_2101,N_1823,N_1793);
nor U2102 (N_2102,N_1510,N_1766);
and U2103 (N_2103,N_1811,N_1724);
nor U2104 (N_2104,N_1710,N_1873);
nand U2105 (N_2105,N_1933,N_1515);
nand U2106 (N_2106,N_1551,N_1979);
or U2107 (N_2107,N_1612,N_1838);
or U2108 (N_2108,N_1866,N_1843);
and U2109 (N_2109,N_1832,N_1504);
nand U2110 (N_2110,N_1992,N_1563);
nor U2111 (N_2111,N_1544,N_1792);
and U2112 (N_2112,N_1607,N_1713);
nor U2113 (N_2113,N_1554,N_1712);
and U2114 (N_2114,N_1781,N_1758);
nand U2115 (N_2115,N_1728,N_1849);
nor U2116 (N_2116,N_1935,N_1802);
nor U2117 (N_2117,N_1630,N_1577);
and U2118 (N_2118,N_1867,N_1826);
and U2119 (N_2119,N_1578,N_1801);
and U2120 (N_2120,N_1820,N_1808);
nor U2121 (N_2121,N_1963,N_1853);
nor U2122 (N_2122,N_1535,N_1809);
and U2123 (N_2123,N_1736,N_1732);
nor U2124 (N_2124,N_1875,N_1615);
nand U2125 (N_2125,N_1759,N_1942);
nor U2126 (N_2126,N_1877,N_1972);
nor U2127 (N_2127,N_1773,N_1651);
xnor U2128 (N_2128,N_1915,N_1605);
nand U2129 (N_2129,N_1623,N_1748);
and U2130 (N_2130,N_1749,N_1705);
or U2131 (N_2131,N_1782,N_1549);
xor U2132 (N_2132,N_1635,N_1540);
nor U2133 (N_2133,N_1930,N_1680);
and U2134 (N_2134,N_1753,N_1834);
nand U2135 (N_2135,N_1521,N_1989);
nor U2136 (N_2136,N_1879,N_1513);
and U2137 (N_2137,N_1628,N_1672);
nor U2138 (N_2138,N_1636,N_1741);
nor U2139 (N_2139,N_1859,N_1610);
nor U2140 (N_2140,N_1642,N_1783);
nor U2141 (N_2141,N_1913,N_1778);
nand U2142 (N_2142,N_1911,N_1687);
xnor U2143 (N_2143,N_1800,N_1548);
nor U2144 (N_2144,N_1679,N_1991);
nand U2145 (N_2145,N_1822,N_1627);
xor U2146 (N_2146,N_1754,N_1516);
and U2147 (N_2147,N_1921,N_1886);
xnor U2148 (N_2148,N_1542,N_1905);
nor U2149 (N_2149,N_1606,N_1556);
and U2150 (N_2150,N_1893,N_1706);
nand U2151 (N_2151,N_1825,N_1638);
and U2152 (N_2152,N_1912,N_1599);
nor U2153 (N_2153,N_1719,N_1957);
nor U2154 (N_2154,N_1920,N_1788);
and U2155 (N_2155,N_1727,N_1787);
or U2156 (N_2156,N_1729,N_1827);
or U2157 (N_2157,N_1986,N_1512);
nand U2158 (N_2158,N_1592,N_1862);
and U2159 (N_2159,N_1927,N_1525);
nor U2160 (N_2160,N_1804,N_1976);
nand U2161 (N_2161,N_1740,N_1568);
nor U2162 (N_2162,N_1530,N_1842);
or U2163 (N_2163,N_1688,N_1586);
nor U2164 (N_2164,N_1669,N_1874);
nor U2165 (N_2165,N_1685,N_1946);
xnor U2166 (N_2166,N_1734,N_1743);
and U2167 (N_2167,N_1693,N_1903);
and U2168 (N_2168,N_1718,N_1836);
or U2169 (N_2169,N_1645,N_1847);
xnor U2170 (N_2170,N_1772,N_1611);
or U2171 (N_2171,N_1564,N_1854);
nor U2172 (N_2172,N_1667,N_1897);
nor U2173 (N_2173,N_1507,N_1501);
or U2174 (N_2174,N_1835,N_1509);
nor U2175 (N_2175,N_1815,N_1735);
or U2176 (N_2176,N_1971,N_1558);
nor U2177 (N_2177,N_1876,N_1914);
nand U2178 (N_2178,N_1789,N_1618);
and U2179 (N_2179,N_1951,N_1596);
xor U2180 (N_2180,N_1892,N_1967);
and U2181 (N_2181,N_1681,N_1598);
xor U2182 (N_2182,N_1725,N_1981);
or U2183 (N_2183,N_1944,N_1514);
nor U2184 (N_2184,N_1524,N_1546);
or U2185 (N_2185,N_1945,N_1602);
nor U2186 (N_2186,N_1502,N_1591);
nor U2187 (N_2187,N_1965,N_1952);
and U2188 (N_2188,N_1574,N_1594);
or U2189 (N_2189,N_1865,N_1714);
nand U2190 (N_2190,N_1765,N_1993);
or U2191 (N_2191,N_1768,N_1885);
or U2192 (N_2192,N_1543,N_1597);
nand U2193 (N_2193,N_1959,N_1878);
or U2194 (N_2194,N_1939,N_1918);
or U2195 (N_2195,N_1634,N_1580);
and U2196 (N_2196,N_1584,N_1716);
nand U2197 (N_2197,N_1650,N_1626);
nor U2198 (N_2198,N_1818,N_1780);
or U2199 (N_2199,N_1656,N_1620);
nand U2200 (N_2200,N_1536,N_1534);
nand U2201 (N_2201,N_1990,N_1522);
or U2202 (N_2202,N_1527,N_1817);
nor U2203 (N_2203,N_1665,N_1816);
xor U2204 (N_2204,N_1756,N_1767);
and U2205 (N_2205,N_1689,N_1857);
nand U2206 (N_2206,N_1840,N_1762);
nor U2207 (N_2207,N_1660,N_1701);
and U2208 (N_2208,N_1648,N_1587);
and U2209 (N_2209,N_1923,N_1595);
or U2210 (N_2210,N_1796,N_1508);
and U2211 (N_2211,N_1720,N_1864);
nor U2212 (N_2212,N_1552,N_1956);
nor U2213 (N_2213,N_1675,N_1998);
or U2214 (N_2214,N_1906,N_1902);
and U2215 (N_2215,N_1601,N_1593);
nor U2216 (N_2216,N_1806,N_1882);
nand U2217 (N_2217,N_1600,N_1797);
and U2218 (N_2218,N_1786,N_1858);
or U2219 (N_2219,N_1966,N_1926);
xnor U2220 (N_2220,N_1997,N_1703);
and U2221 (N_2221,N_1659,N_1621);
nor U2222 (N_2222,N_1700,N_1901);
nor U2223 (N_2223,N_1884,N_1757);
and U2224 (N_2224,N_1553,N_1833);
or U2225 (N_2225,N_1922,N_1761);
and U2226 (N_2226,N_1996,N_1746);
and U2227 (N_2227,N_1790,N_1791);
nand U2228 (N_2228,N_1505,N_1562);
and U2229 (N_2229,N_1738,N_1711);
and U2230 (N_2230,N_1814,N_1609);
nand U2231 (N_2231,N_1863,N_1777);
and U2232 (N_2232,N_1856,N_1646);
and U2233 (N_2233,N_1589,N_1831);
nor U2234 (N_2234,N_1625,N_1807);
and U2235 (N_2235,N_1537,N_1883);
or U2236 (N_2236,N_1980,N_1932);
nor U2237 (N_2237,N_1695,N_1696);
nand U2238 (N_2238,N_1974,N_1604);
nor U2239 (N_2239,N_1968,N_1960);
and U2240 (N_2240,N_1733,N_1810);
or U2241 (N_2241,N_1737,N_1969);
or U2242 (N_2242,N_1845,N_1694);
nand U2243 (N_2243,N_1851,N_1613);
and U2244 (N_2244,N_1624,N_1581);
nand U2245 (N_2245,N_1671,N_1590);
xnor U2246 (N_2246,N_1520,N_1948);
or U2247 (N_2247,N_1975,N_1964);
xor U2248 (N_2248,N_1824,N_1538);
xor U2249 (N_2249,N_1852,N_1764);
nand U2250 (N_2250,N_1522,N_1776);
or U2251 (N_2251,N_1963,N_1998);
and U2252 (N_2252,N_1829,N_1503);
nor U2253 (N_2253,N_1630,N_1846);
nor U2254 (N_2254,N_1864,N_1508);
or U2255 (N_2255,N_1815,N_1962);
nor U2256 (N_2256,N_1898,N_1828);
xnor U2257 (N_2257,N_1661,N_1505);
xor U2258 (N_2258,N_1534,N_1609);
and U2259 (N_2259,N_1626,N_1743);
or U2260 (N_2260,N_1582,N_1543);
or U2261 (N_2261,N_1927,N_1905);
nand U2262 (N_2262,N_1814,N_1568);
nand U2263 (N_2263,N_1993,N_1857);
or U2264 (N_2264,N_1581,N_1661);
or U2265 (N_2265,N_1631,N_1881);
nand U2266 (N_2266,N_1794,N_1969);
or U2267 (N_2267,N_1571,N_1992);
or U2268 (N_2268,N_1746,N_1812);
or U2269 (N_2269,N_1914,N_1960);
or U2270 (N_2270,N_1668,N_1940);
or U2271 (N_2271,N_1631,N_1638);
nand U2272 (N_2272,N_1781,N_1727);
and U2273 (N_2273,N_1999,N_1876);
nand U2274 (N_2274,N_1768,N_1857);
or U2275 (N_2275,N_1889,N_1824);
and U2276 (N_2276,N_1978,N_1960);
or U2277 (N_2277,N_1933,N_1865);
nor U2278 (N_2278,N_1562,N_1872);
and U2279 (N_2279,N_1538,N_1687);
and U2280 (N_2280,N_1727,N_1610);
xor U2281 (N_2281,N_1772,N_1717);
xnor U2282 (N_2282,N_1987,N_1794);
xor U2283 (N_2283,N_1987,N_1801);
or U2284 (N_2284,N_1611,N_1877);
nand U2285 (N_2285,N_1876,N_1735);
and U2286 (N_2286,N_1758,N_1767);
nor U2287 (N_2287,N_1728,N_1863);
or U2288 (N_2288,N_1999,N_1847);
and U2289 (N_2289,N_1626,N_1940);
and U2290 (N_2290,N_1991,N_1507);
nor U2291 (N_2291,N_1911,N_1733);
nor U2292 (N_2292,N_1917,N_1835);
nor U2293 (N_2293,N_1681,N_1966);
nor U2294 (N_2294,N_1957,N_1906);
nand U2295 (N_2295,N_1737,N_1772);
or U2296 (N_2296,N_1937,N_1678);
and U2297 (N_2297,N_1671,N_1917);
and U2298 (N_2298,N_1684,N_1865);
xor U2299 (N_2299,N_1726,N_1594);
xor U2300 (N_2300,N_1721,N_1829);
xor U2301 (N_2301,N_1564,N_1980);
or U2302 (N_2302,N_1698,N_1849);
xor U2303 (N_2303,N_1553,N_1583);
and U2304 (N_2304,N_1642,N_1562);
nor U2305 (N_2305,N_1929,N_1775);
and U2306 (N_2306,N_1925,N_1762);
and U2307 (N_2307,N_1770,N_1650);
nand U2308 (N_2308,N_1682,N_1509);
nand U2309 (N_2309,N_1670,N_1999);
nand U2310 (N_2310,N_1858,N_1662);
and U2311 (N_2311,N_1565,N_1632);
nand U2312 (N_2312,N_1745,N_1791);
or U2313 (N_2313,N_1581,N_1877);
or U2314 (N_2314,N_1580,N_1948);
or U2315 (N_2315,N_1687,N_1756);
or U2316 (N_2316,N_1813,N_1980);
and U2317 (N_2317,N_1724,N_1939);
nor U2318 (N_2318,N_1882,N_1983);
nor U2319 (N_2319,N_1576,N_1786);
and U2320 (N_2320,N_1897,N_1564);
or U2321 (N_2321,N_1536,N_1617);
xnor U2322 (N_2322,N_1824,N_1936);
nand U2323 (N_2323,N_1926,N_1847);
and U2324 (N_2324,N_1517,N_1806);
or U2325 (N_2325,N_1568,N_1911);
nand U2326 (N_2326,N_1874,N_1704);
nand U2327 (N_2327,N_1757,N_1891);
nor U2328 (N_2328,N_1624,N_1625);
nand U2329 (N_2329,N_1509,N_1782);
nor U2330 (N_2330,N_1860,N_1667);
nand U2331 (N_2331,N_1504,N_1979);
nand U2332 (N_2332,N_1915,N_1754);
nand U2333 (N_2333,N_1649,N_1899);
or U2334 (N_2334,N_1777,N_1753);
or U2335 (N_2335,N_1977,N_1892);
or U2336 (N_2336,N_1526,N_1603);
nand U2337 (N_2337,N_1650,N_1522);
or U2338 (N_2338,N_1816,N_1525);
xnor U2339 (N_2339,N_1661,N_1959);
xnor U2340 (N_2340,N_1868,N_1693);
nor U2341 (N_2341,N_1527,N_1705);
nor U2342 (N_2342,N_1917,N_1578);
or U2343 (N_2343,N_1609,N_1918);
and U2344 (N_2344,N_1724,N_1746);
or U2345 (N_2345,N_1946,N_1581);
or U2346 (N_2346,N_1873,N_1567);
and U2347 (N_2347,N_1633,N_1603);
nand U2348 (N_2348,N_1779,N_1566);
or U2349 (N_2349,N_1627,N_1525);
or U2350 (N_2350,N_1590,N_1809);
or U2351 (N_2351,N_1515,N_1819);
or U2352 (N_2352,N_1893,N_1971);
xnor U2353 (N_2353,N_1803,N_1777);
nor U2354 (N_2354,N_1547,N_1679);
nor U2355 (N_2355,N_1528,N_1678);
and U2356 (N_2356,N_1684,N_1525);
and U2357 (N_2357,N_1970,N_1601);
nor U2358 (N_2358,N_1665,N_1626);
nand U2359 (N_2359,N_1943,N_1750);
and U2360 (N_2360,N_1859,N_1869);
nor U2361 (N_2361,N_1601,N_1938);
nor U2362 (N_2362,N_1986,N_1619);
nand U2363 (N_2363,N_1549,N_1813);
and U2364 (N_2364,N_1627,N_1952);
xnor U2365 (N_2365,N_1590,N_1851);
or U2366 (N_2366,N_1617,N_1902);
or U2367 (N_2367,N_1541,N_1530);
or U2368 (N_2368,N_1601,N_1553);
and U2369 (N_2369,N_1874,N_1577);
or U2370 (N_2370,N_1848,N_1602);
nand U2371 (N_2371,N_1782,N_1648);
nand U2372 (N_2372,N_1542,N_1914);
and U2373 (N_2373,N_1675,N_1616);
or U2374 (N_2374,N_1567,N_1831);
nand U2375 (N_2375,N_1576,N_1876);
or U2376 (N_2376,N_1982,N_1861);
and U2377 (N_2377,N_1706,N_1683);
nor U2378 (N_2378,N_1647,N_1712);
nor U2379 (N_2379,N_1624,N_1994);
nor U2380 (N_2380,N_1831,N_1568);
xor U2381 (N_2381,N_1852,N_1670);
nor U2382 (N_2382,N_1975,N_1525);
nor U2383 (N_2383,N_1676,N_1853);
xnor U2384 (N_2384,N_1957,N_1520);
and U2385 (N_2385,N_1597,N_1971);
and U2386 (N_2386,N_1876,N_1746);
nor U2387 (N_2387,N_1714,N_1599);
or U2388 (N_2388,N_1987,N_1672);
xor U2389 (N_2389,N_1943,N_1653);
nand U2390 (N_2390,N_1589,N_1752);
or U2391 (N_2391,N_1974,N_1766);
nor U2392 (N_2392,N_1926,N_1998);
or U2393 (N_2393,N_1845,N_1905);
xnor U2394 (N_2394,N_1521,N_1831);
and U2395 (N_2395,N_1542,N_1764);
nand U2396 (N_2396,N_1703,N_1641);
or U2397 (N_2397,N_1703,N_1617);
nand U2398 (N_2398,N_1550,N_1693);
xor U2399 (N_2399,N_1855,N_1929);
nand U2400 (N_2400,N_1943,N_1954);
or U2401 (N_2401,N_1672,N_1618);
or U2402 (N_2402,N_1979,N_1881);
nand U2403 (N_2403,N_1821,N_1589);
nor U2404 (N_2404,N_1744,N_1981);
nor U2405 (N_2405,N_1599,N_1689);
or U2406 (N_2406,N_1502,N_1594);
or U2407 (N_2407,N_1620,N_1880);
or U2408 (N_2408,N_1850,N_1984);
or U2409 (N_2409,N_1899,N_1713);
nand U2410 (N_2410,N_1887,N_1537);
or U2411 (N_2411,N_1880,N_1622);
or U2412 (N_2412,N_1934,N_1702);
and U2413 (N_2413,N_1524,N_1581);
nand U2414 (N_2414,N_1929,N_1691);
nor U2415 (N_2415,N_1756,N_1778);
xnor U2416 (N_2416,N_1632,N_1705);
and U2417 (N_2417,N_1814,N_1974);
and U2418 (N_2418,N_1634,N_1597);
nand U2419 (N_2419,N_1703,N_1824);
nor U2420 (N_2420,N_1511,N_1635);
xnor U2421 (N_2421,N_1527,N_1794);
nand U2422 (N_2422,N_1747,N_1878);
nand U2423 (N_2423,N_1825,N_1941);
nor U2424 (N_2424,N_1822,N_1567);
nor U2425 (N_2425,N_1681,N_1587);
and U2426 (N_2426,N_1688,N_1810);
nand U2427 (N_2427,N_1567,N_1800);
nor U2428 (N_2428,N_1732,N_1616);
and U2429 (N_2429,N_1618,N_1517);
xnor U2430 (N_2430,N_1968,N_1811);
and U2431 (N_2431,N_1785,N_1807);
and U2432 (N_2432,N_1843,N_1982);
or U2433 (N_2433,N_1577,N_1631);
nand U2434 (N_2434,N_1865,N_1953);
nor U2435 (N_2435,N_1810,N_1778);
and U2436 (N_2436,N_1665,N_1606);
and U2437 (N_2437,N_1880,N_1825);
nor U2438 (N_2438,N_1764,N_1617);
xor U2439 (N_2439,N_1783,N_1511);
and U2440 (N_2440,N_1721,N_1933);
and U2441 (N_2441,N_1507,N_1780);
and U2442 (N_2442,N_1547,N_1743);
and U2443 (N_2443,N_1928,N_1723);
nor U2444 (N_2444,N_1604,N_1758);
or U2445 (N_2445,N_1504,N_1983);
nand U2446 (N_2446,N_1962,N_1798);
nand U2447 (N_2447,N_1512,N_1962);
and U2448 (N_2448,N_1832,N_1723);
and U2449 (N_2449,N_1977,N_1896);
nor U2450 (N_2450,N_1735,N_1603);
nor U2451 (N_2451,N_1752,N_1726);
or U2452 (N_2452,N_1716,N_1798);
and U2453 (N_2453,N_1542,N_1676);
and U2454 (N_2454,N_1791,N_1811);
or U2455 (N_2455,N_1897,N_1523);
and U2456 (N_2456,N_1628,N_1757);
nand U2457 (N_2457,N_1653,N_1647);
or U2458 (N_2458,N_1951,N_1858);
xor U2459 (N_2459,N_1854,N_1570);
or U2460 (N_2460,N_1906,N_1673);
and U2461 (N_2461,N_1922,N_1977);
or U2462 (N_2462,N_1521,N_1723);
nor U2463 (N_2463,N_1513,N_1728);
nand U2464 (N_2464,N_1891,N_1680);
nand U2465 (N_2465,N_1629,N_1827);
or U2466 (N_2466,N_1546,N_1993);
nor U2467 (N_2467,N_1579,N_1981);
or U2468 (N_2468,N_1731,N_1533);
xnor U2469 (N_2469,N_1517,N_1674);
xnor U2470 (N_2470,N_1799,N_1860);
and U2471 (N_2471,N_1617,N_1828);
nand U2472 (N_2472,N_1832,N_1909);
xnor U2473 (N_2473,N_1921,N_1919);
nor U2474 (N_2474,N_1680,N_1548);
or U2475 (N_2475,N_1949,N_1663);
nor U2476 (N_2476,N_1560,N_1722);
nand U2477 (N_2477,N_1681,N_1823);
or U2478 (N_2478,N_1963,N_1940);
nor U2479 (N_2479,N_1543,N_1998);
nand U2480 (N_2480,N_1967,N_1790);
and U2481 (N_2481,N_1683,N_1648);
and U2482 (N_2482,N_1571,N_1844);
and U2483 (N_2483,N_1595,N_1539);
nand U2484 (N_2484,N_1907,N_1606);
and U2485 (N_2485,N_1977,N_1971);
and U2486 (N_2486,N_1626,N_1868);
nand U2487 (N_2487,N_1643,N_1942);
or U2488 (N_2488,N_1666,N_1834);
and U2489 (N_2489,N_1965,N_1982);
or U2490 (N_2490,N_1548,N_1681);
or U2491 (N_2491,N_1688,N_1686);
and U2492 (N_2492,N_1984,N_1670);
nor U2493 (N_2493,N_1709,N_1746);
and U2494 (N_2494,N_1909,N_1661);
or U2495 (N_2495,N_1621,N_1733);
or U2496 (N_2496,N_1945,N_1508);
or U2497 (N_2497,N_1994,N_1515);
nand U2498 (N_2498,N_1993,N_1904);
and U2499 (N_2499,N_1810,N_1790);
nand U2500 (N_2500,N_2181,N_2097);
nand U2501 (N_2501,N_2083,N_2258);
or U2502 (N_2502,N_2367,N_2287);
nand U2503 (N_2503,N_2235,N_2248);
or U2504 (N_2504,N_2146,N_2392);
nor U2505 (N_2505,N_2124,N_2301);
or U2506 (N_2506,N_2055,N_2382);
nand U2507 (N_2507,N_2316,N_2034);
nor U2508 (N_2508,N_2335,N_2119);
nor U2509 (N_2509,N_2267,N_2195);
nand U2510 (N_2510,N_2458,N_2187);
nand U2511 (N_2511,N_2449,N_2320);
and U2512 (N_2512,N_2020,N_2385);
or U2513 (N_2513,N_2380,N_2089);
nor U2514 (N_2514,N_2217,N_2472);
and U2515 (N_2515,N_2305,N_2161);
nor U2516 (N_2516,N_2049,N_2017);
and U2517 (N_2517,N_2461,N_2384);
or U2518 (N_2518,N_2088,N_2370);
or U2519 (N_2519,N_2469,N_2206);
and U2520 (N_2520,N_2052,N_2318);
nand U2521 (N_2521,N_2118,N_2031);
nand U2522 (N_2522,N_2022,N_2252);
or U2523 (N_2523,N_2211,N_2349);
nor U2524 (N_2524,N_2149,N_2074);
nand U2525 (N_2525,N_2053,N_2369);
xor U2526 (N_2526,N_2038,N_2143);
xnor U2527 (N_2527,N_2485,N_2327);
and U2528 (N_2528,N_2404,N_2147);
or U2529 (N_2529,N_2168,N_2047);
xnor U2530 (N_2530,N_2006,N_2309);
or U2531 (N_2531,N_2304,N_2064);
nor U2532 (N_2532,N_2131,N_2105);
nor U2533 (N_2533,N_2411,N_2062);
and U2534 (N_2534,N_2448,N_2101);
xnor U2535 (N_2535,N_2428,N_2442);
xnor U2536 (N_2536,N_2078,N_2303);
nor U2537 (N_2537,N_2208,N_2390);
or U2538 (N_2538,N_2201,N_2160);
nor U2539 (N_2539,N_2285,N_2044);
nor U2540 (N_2540,N_2441,N_2003);
nor U2541 (N_2541,N_2165,N_2478);
or U2542 (N_2542,N_2107,N_2480);
nand U2543 (N_2543,N_2117,N_2266);
and U2544 (N_2544,N_2223,N_2154);
nand U2545 (N_2545,N_2346,N_2276);
nor U2546 (N_2546,N_2460,N_2113);
nand U2547 (N_2547,N_2256,N_2122);
and U2548 (N_2548,N_2210,N_2099);
xnor U2549 (N_2549,N_2462,N_2455);
xor U2550 (N_2550,N_2227,N_2274);
nor U2551 (N_2551,N_2130,N_2219);
and U2552 (N_2552,N_2232,N_2151);
nand U2553 (N_2553,N_2457,N_2126);
xor U2554 (N_2554,N_2324,N_2185);
and U2555 (N_2555,N_2467,N_2016);
nand U2556 (N_2556,N_2387,N_2395);
nand U2557 (N_2557,N_2138,N_2493);
nor U2558 (N_2558,N_2123,N_2296);
nand U2559 (N_2559,N_2239,N_2025);
nand U2560 (N_2560,N_2344,N_2036);
and U2561 (N_2561,N_2353,N_2262);
or U2562 (N_2562,N_2439,N_2333);
or U2563 (N_2563,N_2018,N_2070);
or U2564 (N_2564,N_2087,N_2269);
xnor U2565 (N_2565,N_2191,N_2365);
and U2566 (N_2566,N_2388,N_2121);
and U2567 (N_2567,N_2032,N_2495);
nand U2568 (N_2568,N_2104,N_2242);
nor U2569 (N_2569,N_2444,N_2141);
and U2570 (N_2570,N_2471,N_2278);
and U2571 (N_2571,N_2229,N_2090);
or U2572 (N_2572,N_2401,N_2356);
or U2573 (N_2573,N_2207,N_2376);
nand U2574 (N_2574,N_2215,N_2290);
and U2575 (N_2575,N_2407,N_2360);
nor U2576 (N_2576,N_2203,N_2076);
or U2577 (N_2577,N_2257,N_2073);
and U2578 (N_2578,N_2427,N_2486);
xnor U2579 (N_2579,N_2477,N_2354);
or U2580 (N_2580,N_2013,N_2081);
nand U2581 (N_2581,N_2204,N_2255);
nor U2582 (N_2582,N_2128,N_2222);
and U2583 (N_2583,N_2364,N_2288);
and U2584 (N_2584,N_2005,N_2422);
nand U2585 (N_2585,N_2112,N_2155);
nor U2586 (N_2586,N_2297,N_2093);
or U2587 (N_2587,N_2339,N_2129);
nor U2588 (N_2588,N_2136,N_2007);
and U2589 (N_2589,N_2426,N_2177);
or U2590 (N_2590,N_2280,N_2023);
or U2591 (N_2591,N_2043,N_2192);
and U2592 (N_2592,N_2412,N_2338);
and U2593 (N_2593,N_2092,N_2014);
and U2594 (N_2594,N_2035,N_2202);
or U2595 (N_2595,N_2488,N_2473);
nand U2596 (N_2596,N_2228,N_2051);
xor U2597 (N_2597,N_2283,N_2347);
nor U2598 (N_2598,N_2286,N_2205);
nand U2599 (N_2599,N_2487,N_2326);
nand U2600 (N_2600,N_2362,N_2132);
xnor U2601 (N_2601,N_2425,N_2402);
nor U2602 (N_2602,N_2348,N_2277);
nand U2603 (N_2603,N_2000,N_2225);
nand U2604 (N_2604,N_2397,N_2230);
nand U2605 (N_2605,N_2366,N_2321);
and U2606 (N_2606,N_2483,N_2340);
nand U2607 (N_2607,N_2443,N_2270);
nand U2608 (N_2608,N_2189,N_2220);
or U2609 (N_2609,N_2450,N_2259);
nand U2610 (N_2610,N_2357,N_2358);
nand U2611 (N_2611,N_2445,N_2419);
or U2612 (N_2612,N_2331,N_2307);
and U2613 (N_2613,N_2437,N_2153);
nand U2614 (N_2614,N_2102,N_2406);
and U2615 (N_2615,N_2260,N_2498);
or U2616 (N_2616,N_2332,N_2246);
or U2617 (N_2617,N_2325,N_2372);
nand U2618 (N_2618,N_2175,N_2075);
or U2619 (N_2619,N_2158,N_2001);
xnor U2620 (N_2620,N_2396,N_2250);
or U2621 (N_2621,N_2424,N_2183);
or U2622 (N_2622,N_2456,N_2135);
and U2623 (N_2623,N_2271,N_2436);
or U2624 (N_2624,N_2438,N_2150);
and U2625 (N_2625,N_2152,N_2253);
nor U2626 (N_2626,N_2029,N_2139);
or U2627 (N_2627,N_2383,N_2440);
or U2628 (N_2628,N_2039,N_2178);
xor U2629 (N_2629,N_2067,N_2140);
xnor U2630 (N_2630,N_2490,N_2243);
nor U2631 (N_2631,N_2176,N_2416);
nand U2632 (N_2632,N_2061,N_2080);
nor U2633 (N_2633,N_2468,N_2050);
nand U2634 (N_2634,N_2291,N_2209);
nand U2635 (N_2635,N_2447,N_2027);
nand U2636 (N_2636,N_2409,N_2096);
nor U2637 (N_2637,N_2275,N_2041);
or U2638 (N_2638,N_2342,N_2323);
nor U2639 (N_2639,N_2019,N_2085);
nand U2640 (N_2640,N_2294,N_2166);
and U2641 (N_2641,N_2106,N_2162);
or U2642 (N_2642,N_2476,N_2399);
nor U2643 (N_2643,N_2174,N_2184);
nor U2644 (N_2644,N_2079,N_2298);
nand U2645 (N_2645,N_2060,N_2116);
nand U2646 (N_2646,N_2247,N_2312);
nor U2647 (N_2647,N_2491,N_2418);
and U2648 (N_2648,N_2002,N_2351);
and U2649 (N_2649,N_2453,N_2413);
and U2650 (N_2650,N_2234,N_2337);
and U2651 (N_2651,N_2196,N_2224);
nand U2652 (N_2652,N_2361,N_2343);
or U2653 (N_2653,N_2492,N_2497);
or U2654 (N_2654,N_2499,N_2265);
nand U2655 (N_2655,N_2008,N_2310);
or U2656 (N_2656,N_2110,N_2408);
nor U2657 (N_2657,N_2058,N_2179);
or U2658 (N_2658,N_2186,N_2293);
or U2659 (N_2659,N_2355,N_2432);
nor U2660 (N_2660,N_2381,N_2496);
nor U2661 (N_2661,N_2459,N_2417);
nor U2662 (N_2662,N_2314,N_2420);
xnor U2663 (N_2663,N_2216,N_2302);
xor U2664 (N_2664,N_2429,N_2482);
nor U2665 (N_2665,N_2111,N_2386);
nand U2666 (N_2666,N_2197,N_2045);
nand U2667 (N_2667,N_2273,N_2170);
nand U2668 (N_2668,N_2172,N_2015);
or U2669 (N_2669,N_2193,N_2494);
or U2670 (N_2670,N_2137,N_2037);
or U2671 (N_2671,N_2198,N_2263);
and U2672 (N_2672,N_2048,N_2299);
and U2673 (N_2673,N_2466,N_2414);
and U2674 (N_2674,N_2133,N_2054);
or U2675 (N_2675,N_2373,N_2159);
nor U2676 (N_2676,N_2452,N_2200);
nor U2677 (N_2677,N_2245,N_2264);
and U2678 (N_2678,N_2268,N_2240);
nand U2679 (N_2679,N_2378,N_2095);
or U2680 (N_2680,N_2410,N_2328);
and U2681 (N_2681,N_2464,N_2394);
xor U2682 (N_2682,N_2292,N_2341);
nand U2683 (N_2683,N_2345,N_2167);
xor U2684 (N_2684,N_2134,N_2282);
nand U2685 (N_2685,N_2086,N_2156);
xnor U2686 (N_2686,N_2311,N_2330);
and U2687 (N_2687,N_2163,N_2470);
and U2688 (N_2688,N_2281,N_2180);
and U2689 (N_2689,N_2434,N_2094);
and U2690 (N_2690,N_2033,N_2212);
or U2691 (N_2691,N_2405,N_2415);
or U2692 (N_2692,N_2231,N_2463);
nor U2693 (N_2693,N_2423,N_2221);
or U2694 (N_2694,N_2289,N_2059);
nor U2695 (N_2695,N_2329,N_2254);
nand U2696 (N_2696,N_2238,N_2431);
or U2697 (N_2697,N_2421,N_2103);
or U2698 (N_2698,N_2433,N_2363);
xor U2699 (N_2699,N_2173,N_2479);
nor U2700 (N_2700,N_2249,N_2484);
nor U2701 (N_2701,N_2077,N_2115);
nor U2702 (N_2702,N_2352,N_2403);
or U2703 (N_2703,N_2114,N_2040);
or U2704 (N_2704,N_2319,N_2334);
and U2705 (N_2705,N_2371,N_2148);
or U2706 (N_2706,N_2030,N_2226);
nor U2707 (N_2707,N_2391,N_2157);
nand U2708 (N_2708,N_2308,N_2026);
and U2709 (N_2709,N_2481,N_2435);
and U2710 (N_2710,N_2084,N_2190);
nor U2711 (N_2711,N_2244,N_2489);
nor U2712 (N_2712,N_2199,N_2100);
or U2713 (N_2713,N_2272,N_2237);
and U2714 (N_2714,N_2295,N_2315);
or U2715 (N_2715,N_2400,N_2389);
and U2716 (N_2716,N_2012,N_2063);
and U2717 (N_2717,N_2214,N_2046);
nor U2718 (N_2718,N_2194,N_2024);
and U2719 (N_2719,N_2071,N_2474);
and U2720 (N_2720,N_2120,N_2375);
and U2721 (N_2721,N_2233,N_2313);
xor U2722 (N_2722,N_2475,N_2028);
or U2723 (N_2723,N_2236,N_2171);
or U2724 (N_2724,N_2454,N_2142);
nor U2725 (N_2725,N_2393,N_2068);
or U2726 (N_2726,N_2065,N_2336);
xor U2727 (N_2727,N_2057,N_2056);
xnor U2728 (N_2728,N_2377,N_2374);
or U2729 (N_2729,N_2451,N_2145);
and U2730 (N_2730,N_2010,N_2011);
xor U2731 (N_2731,N_2188,N_2359);
and U2732 (N_2732,N_2213,N_2430);
and U2733 (N_2733,N_2279,N_2368);
or U2734 (N_2734,N_2164,N_2398);
nand U2735 (N_2735,N_2379,N_2091);
nand U2736 (N_2736,N_2109,N_2322);
nor U2737 (N_2737,N_2021,N_2066);
nor U2738 (N_2738,N_2284,N_2306);
or U2739 (N_2739,N_2042,N_2218);
and U2740 (N_2740,N_2261,N_2108);
nor U2741 (N_2741,N_2098,N_2144);
nand U2742 (N_2742,N_2127,N_2125);
nand U2743 (N_2743,N_2465,N_2241);
nand U2744 (N_2744,N_2251,N_2317);
nand U2745 (N_2745,N_2300,N_2182);
xnor U2746 (N_2746,N_2069,N_2004);
or U2747 (N_2747,N_2009,N_2350);
nor U2748 (N_2748,N_2082,N_2446);
and U2749 (N_2749,N_2169,N_2072);
nor U2750 (N_2750,N_2120,N_2294);
or U2751 (N_2751,N_2425,N_2278);
nand U2752 (N_2752,N_2469,N_2373);
nand U2753 (N_2753,N_2244,N_2204);
and U2754 (N_2754,N_2462,N_2043);
nor U2755 (N_2755,N_2176,N_2274);
and U2756 (N_2756,N_2104,N_2071);
and U2757 (N_2757,N_2141,N_2137);
nand U2758 (N_2758,N_2313,N_2348);
and U2759 (N_2759,N_2483,N_2117);
and U2760 (N_2760,N_2042,N_2331);
nor U2761 (N_2761,N_2351,N_2306);
nor U2762 (N_2762,N_2379,N_2157);
nor U2763 (N_2763,N_2078,N_2464);
nand U2764 (N_2764,N_2448,N_2087);
or U2765 (N_2765,N_2487,N_2333);
xor U2766 (N_2766,N_2211,N_2327);
nand U2767 (N_2767,N_2474,N_2091);
xor U2768 (N_2768,N_2395,N_2057);
or U2769 (N_2769,N_2345,N_2101);
nand U2770 (N_2770,N_2463,N_2312);
nor U2771 (N_2771,N_2300,N_2140);
nand U2772 (N_2772,N_2233,N_2457);
nor U2773 (N_2773,N_2408,N_2415);
xor U2774 (N_2774,N_2427,N_2156);
or U2775 (N_2775,N_2315,N_2484);
or U2776 (N_2776,N_2357,N_2239);
and U2777 (N_2777,N_2384,N_2338);
nor U2778 (N_2778,N_2348,N_2298);
or U2779 (N_2779,N_2239,N_2165);
nand U2780 (N_2780,N_2437,N_2383);
or U2781 (N_2781,N_2144,N_2303);
nand U2782 (N_2782,N_2359,N_2248);
nand U2783 (N_2783,N_2364,N_2314);
xor U2784 (N_2784,N_2382,N_2330);
xnor U2785 (N_2785,N_2195,N_2191);
or U2786 (N_2786,N_2412,N_2109);
nand U2787 (N_2787,N_2498,N_2303);
and U2788 (N_2788,N_2021,N_2303);
xor U2789 (N_2789,N_2131,N_2179);
nand U2790 (N_2790,N_2171,N_2005);
or U2791 (N_2791,N_2108,N_2255);
nor U2792 (N_2792,N_2362,N_2216);
and U2793 (N_2793,N_2076,N_2089);
nor U2794 (N_2794,N_2014,N_2300);
nand U2795 (N_2795,N_2238,N_2401);
or U2796 (N_2796,N_2044,N_2309);
and U2797 (N_2797,N_2352,N_2413);
and U2798 (N_2798,N_2319,N_2423);
nor U2799 (N_2799,N_2037,N_2198);
nor U2800 (N_2800,N_2063,N_2444);
or U2801 (N_2801,N_2084,N_2436);
and U2802 (N_2802,N_2257,N_2330);
nor U2803 (N_2803,N_2015,N_2024);
nand U2804 (N_2804,N_2055,N_2317);
and U2805 (N_2805,N_2474,N_2350);
nand U2806 (N_2806,N_2318,N_2315);
and U2807 (N_2807,N_2459,N_2432);
nor U2808 (N_2808,N_2443,N_2087);
and U2809 (N_2809,N_2482,N_2176);
or U2810 (N_2810,N_2378,N_2110);
nand U2811 (N_2811,N_2034,N_2454);
and U2812 (N_2812,N_2206,N_2092);
and U2813 (N_2813,N_2439,N_2070);
xor U2814 (N_2814,N_2185,N_2147);
nand U2815 (N_2815,N_2301,N_2087);
xnor U2816 (N_2816,N_2178,N_2157);
xor U2817 (N_2817,N_2111,N_2225);
and U2818 (N_2818,N_2387,N_2235);
nor U2819 (N_2819,N_2175,N_2023);
nand U2820 (N_2820,N_2383,N_2091);
and U2821 (N_2821,N_2053,N_2046);
nand U2822 (N_2822,N_2076,N_2141);
nor U2823 (N_2823,N_2136,N_2241);
and U2824 (N_2824,N_2164,N_2062);
or U2825 (N_2825,N_2161,N_2139);
nor U2826 (N_2826,N_2496,N_2273);
xnor U2827 (N_2827,N_2046,N_2200);
and U2828 (N_2828,N_2104,N_2247);
nand U2829 (N_2829,N_2430,N_2169);
and U2830 (N_2830,N_2180,N_2159);
and U2831 (N_2831,N_2168,N_2465);
xnor U2832 (N_2832,N_2387,N_2025);
xnor U2833 (N_2833,N_2359,N_2144);
nor U2834 (N_2834,N_2243,N_2184);
or U2835 (N_2835,N_2028,N_2417);
nand U2836 (N_2836,N_2475,N_2027);
and U2837 (N_2837,N_2473,N_2346);
and U2838 (N_2838,N_2215,N_2285);
nor U2839 (N_2839,N_2308,N_2365);
and U2840 (N_2840,N_2149,N_2415);
nor U2841 (N_2841,N_2022,N_2225);
nor U2842 (N_2842,N_2016,N_2231);
nor U2843 (N_2843,N_2359,N_2355);
nand U2844 (N_2844,N_2307,N_2033);
or U2845 (N_2845,N_2380,N_2131);
nor U2846 (N_2846,N_2245,N_2192);
or U2847 (N_2847,N_2143,N_2056);
nor U2848 (N_2848,N_2224,N_2087);
and U2849 (N_2849,N_2389,N_2318);
nand U2850 (N_2850,N_2216,N_2259);
and U2851 (N_2851,N_2453,N_2042);
and U2852 (N_2852,N_2185,N_2019);
nor U2853 (N_2853,N_2463,N_2336);
or U2854 (N_2854,N_2224,N_2270);
and U2855 (N_2855,N_2309,N_2112);
and U2856 (N_2856,N_2028,N_2249);
nor U2857 (N_2857,N_2172,N_2016);
or U2858 (N_2858,N_2169,N_2167);
nand U2859 (N_2859,N_2120,N_2096);
nand U2860 (N_2860,N_2306,N_2368);
or U2861 (N_2861,N_2404,N_2434);
nor U2862 (N_2862,N_2148,N_2386);
and U2863 (N_2863,N_2411,N_2027);
nand U2864 (N_2864,N_2271,N_2301);
and U2865 (N_2865,N_2175,N_2177);
nand U2866 (N_2866,N_2164,N_2430);
nand U2867 (N_2867,N_2118,N_2300);
xor U2868 (N_2868,N_2294,N_2386);
nor U2869 (N_2869,N_2185,N_2440);
nor U2870 (N_2870,N_2070,N_2205);
nor U2871 (N_2871,N_2069,N_2243);
nor U2872 (N_2872,N_2292,N_2085);
and U2873 (N_2873,N_2180,N_2414);
and U2874 (N_2874,N_2389,N_2029);
and U2875 (N_2875,N_2487,N_2346);
xnor U2876 (N_2876,N_2104,N_2120);
or U2877 (N_2877,N_2415,N_2174);
and U2878 (N_2878,N_2060,N_2367);
or U2879 (N_2879,N_2069,N_2135);
or U2880 (N_2880,N_2314,N_2297);
and U2881 (N_2881,N_2280,N_2276);
or U2882 (N_2882,N_2335,N_2463);
nor U2883 (N_2883,N_2307,N_2382);
nand U2884 (N_2884,N_2432,N_2208);
nand U2885 (N_2885,N_2331,N_2257);
or U2886 (N_2886,N_2370,N_2135);
xnor U2887 (N_2887,N_2495,N_2379);
nand U2888 (N_2888,N_2090,N_2029);
nor U2889 (N_2889,N_2090,N_2428);
xnor U2890 (N_2890,N_2116,N_2343);
nor U2891 (N_2891,N_2033,N_2242);
nor U2892 (N_2892,N_2333,N_2132);
or U2893 (N_2893,N_2048,N_2249);
nand U2894 (N_2894,N_2148,N_2365);
nor U2895 (N_2895,N_2006,N_2287);
xor U2896 (N_2896,N_2035,N_2292);
nor U2897 (N_2897,N_2160,N_2367);
or U2898 (N_2898,N_2213,N_2196);
or U2899 (N_2899,N_2287,N_2123);
and U2900 (N_2900,N_2172,N_2391);
and U2901 (N_2901,N_2039,N_2494);
and U2902 (N_2902,N_2003,N_2345);
nor U2903 (N_2903,N_2453,N_2098);
and U2904 (N_2904,N_2494,N_2260);
nand U2905 (N_2905,N_2225,N_2430);
and U2906 (N_2906,N_2393,N_2094);
nand U2907 (N_2907,N_2401,N_2073);
nand U2908 (N_2908,N_2090,N_2486);
and U2909 (N_2909,N_2001,N_2498);
nor U2910 (N_2910,N_2483,N_2494);
and U2911 (N_2911,N_2336,N_2459);
nor U2912 (N_2912,N_2457,N_2395);
nor U2913 (N_2913,N_2387,N_2333);
nand U2914 (N_2914,N_2219,N_2109);
or U2915 (N_2915,N_2349,N_2056);
or U2916 (N_2916,N_2351,N_2036);
nand U2917 (N_2917,N_2421,N_2262);
nor U2918 (N_2918,N_2224,N_2350);
and U2919 (N_2919,N_2327,N_2105);
or U2920 (N_2920,N_2420,N_2258);
nand U2921 (N_2921,N_2321,N_2205);
and U2922 (N_2922,N_2268,N_2344);
and U2923 (N_2923,N_2307,N_2375);
or U2924 (N_2924,N_2330,N_2373);
and U2925 (N_2925,N_2391,N_2459);
nand U2926 (N_2926,N_2041,N_2050);
xor U2927 (N_2927,N_2025,N_2282);
nand U2928 (N_2928,N_2010,N_2115);
and U2929 (N_2929,N_2089,N_2472);
nor U2930 (N_2930,N_2325,N_2499);
or U2931 (N_2931,N_2092,N_2217);
xor U2932 (N_2932,N_2429,N_2100);
and U2933 (N_2933,N_2080,N_2001);
nand U2934 (N_2934,N_2115,N_2317);
xor U2935 (N_2935,N_2359,N_2311);
nand U2936 (N_2936,N_2300,N_2424);
nand U2937 (N_2937,N_2051,N_2439);
nor U2938 (N_2938,N_2318,N_2106);
and U2939 (N_2939,N_2441,N_2075);
and U2940 (N_2940,N_2294,N_2025);
or U2941 (N_2941,N_2494,N_2273);
nand U2942 (N_2942,N_2473,N_2031);
nand U2943 (N_2943,N_2114,N_2455);
or U2944 (N_2944,N_2244,N_2046);
nand U2945 (N_2945,N_2255,N_2132);
nand U2946 (N_2946,N_2012,N_2329);
and U2947 (N_2947,N_2401,N_2294);
or U2948 (N_2948,N_2296,N_2231);
nand U2949 (N_2949,N_2116,N_2082);
and U2950 (N_2950,N_2191,N_2316);
and U2951 (N_2951,N_2135,N_2348);
nand U2952 (N_2952,N_2113,N_2437);
or U2953 (N_2953,N_2260,N_2285);
nand U2954 (N_2954,N_2162,N_2374);
or U2955 (N_2955,N_2345,N_2189);
and U2956 (N_2956,N_2058,N_2115);
nand U2957 (N_2957,N_2450,N_2069);
and U2958 (N_2958,N_2199,N_2106);
nand U2959 (N_2959,N_2271,N_2177);
and U2960 (N_2960,N_2220,N_2481);
nand U2961 (N_2961,N_2317,N_2054);
or U2962 (N_2962,N_2246,N_2267);
or U2963 (N_2963,N_2066,N_2010);
nor U2964 (N_2964,N_2202,N_2203);
nor U2965 (N_2965,N_2429,N_2034);
or U2966 (N_2966,N_2169,N_2005);
nand U2967 (N_2967,N_2060,N_2115);
or U2968 (N_2968,N_2260,N_2368);
xnor U2969 (N_2969,N_2418,N_2228);
or U2970 (N_2970,N_2073,N_2332);
nand U2971 (N_2971,N_2146,N_2343);
or U2972 (N_2972,N_2214,N_2363);
and U2973 (N_2973,N_2317,N_2164);
or U2974 (N_2974,N_2128,N_2359);
xnor U2975 (N_2975,N_2454,N_2379);
nand U2976 (N_2976,N_2089,N_2318);
nand U2977 (N_2977,N_2486,N_2268);
nand U2978 (N_2978,N_2263,N_2404);
nand U2979 (N_2979,N_2243,N_2452);
or U2980 (N_2980,N_2495,N_2258);
or U2981 (N_2981,N_2015,N_2130);
nand U2982 (N_2982,N_2067,N_2157);
or U2983 (N_2983,N_2303,N_2107);
nand U2984 (N_2984,N_2050,N_2293);
and U2985 (N_2985,N_2052,N_2321);
nor U2986 (N_2986,N_2008,N_2485);
nor U2987 (N_2987,N_2178,N_2359);
or U2988 (N_2988,N_2490,N_2312);
nand U2989 (N_2989,N_2397,N_2033);
or U2990 (N_2990,N_2253,N_2486);
nand U2991 (N_2991,N_2077,N_2175);
nor U2992 (N_2992,N_2207,N_2322);
and U2993 (N_2993,N_2384,N_2041);
xor U2994 (N_2994,N_2251,N_2047);
and U2995 (N_2995,N_2150,N_2316);
and U2996 (N_2996,N_2160,N_2206);
and U2997 (N_2997,N_2074,N_2410);
nand U2998 (N_2998,N_2040,N_2498);
nor U2999 (N_2999,N_2000,N_2041);
and U3000 (N_3000,N_2641,N_2689);
nor U3001 (N_3001,N_2896,N_2968);
nor U3002 (N_3002,N_2540,N_2505);
or U3003 (N_3003,N_2745,N_2782);
nor U3004 (N_3004,N_2875,N_2506);
and U3005 (N_3005,N_2663,N_2788);
and U3006 (N_3006,N_2862,N_2572);
nand U3007 (N_3007,N_2747,N_2622);
nor U3008 (N_3008,N_2927,N_2885);
nor U3009 (N_3009,N_2691,N_2703);
nor U3010 (N_3010,N_2984,N_2701);
nand U3011 (N_3011,N_2762,N_2751);
nor U3012 (N_3012,N_2970,N_2864);
and U3013 (N_3013,N_2634,N_2675);
nand U3014 (N_3014,N_2738,N_2559);
or U3015 (N_3015,N_2633,N_2826);
or U3016 (N_3016,N_2833,N_2906);
nand U3017 (N_3017,N_2860,N_2585);
and U3018 (N_3018,N_2609,N_2538);
and U3019 (N_3019,N_2817,N_2525);
nor U3020 (N_3020,N_2658,N_2617);
or U3021 (N_3021,N_2953,N_2536);
or U3022 (N_3022,N_2792,N_2618);
nor U3023 (N_3023,N_2846,N_2805);
nor U3024 (N_3024,N_2734,N_2645);
nand U3025 (N_3025,N_2869,N_2892);
or U3026 (N_3026,N_2652,N_2661);
nand U3027 (N_3027,N_2774,N_2548);
and U3028 (N_3028,N_2537,N_2519);
xnor U3029 (N_3029,N_2996,N_2850);
nand U3030 (N_3030,N_2576,N_2770);
nand U3031 (N_3031,N_2898,N_2638);
or U3032 (N_3032,N_2657,N_2836);
nand U3033 (N_3033,N_2966,N_2752);
or U3034 (N_3034,N_2521,N_2640);
nor U3035 (N_3035,N_2508,N_2595);
and U3036 (N_3036,N_2730,N_2513);
or U3037 (N_3037,N_2951,N_2653);
xnor U3038 (N_3038,N_2727,N_2562);
xnor U3039 (N_3039,N_2929,N_2728);
nor U3040 (N_3040,N_2545,N_2676);
nand U3041 (N_3041,N_2733,N_2628);
xor U3042 (N_3042,N_2577,N_2811);
or U3043 (N_3043,N_2871,N_2878);
or U3044 (N_3044,N_2624,N_2565);
or U3045 (N_3045,N_2596,N_2724);
nand U3046 (N_3046,N_2590,N_2709);
or U3047 (N_3047,N_2606,N_2681);
and U3048 (N_3048,N_2771,N_2935);
nor U3049 (N_3049,N_2988,N_2554);
nor U3050 (N_3050,N_2589,N_2903);
and U3051 (N_3051,N_2563,N_2985);
nor U3052 (N_3052,N_2908,N_2720);
or U3053 (N_3053,N_2723,N_2717);
nand U3054 (N_3054,N_2603,N_2839);
nand U3055 (N_3055,N_2736,N_2804);
and U3056 (N_3056,N_2642,N_2821);
or U3057 (N_3057,N_2949,N_2791);
nand U3058 (N_3058,N_2761,N_2743);
nand U3059 (N_3059,N_2719,N_2764);
or U3060 (N_3060,N_2921,N_2650);
nor U3061 (N_3061,N_2810,N_2930);
nand U3062 (N_3062,N_2832,N_2979);
nor U3063 (N_3063,N_2760,N_2754);
nand U3064 (N_3064,N_2763,N_2844);
or U3065 (N_3065,N_2965,N_2943);
or U3066 (N_3066,N_2667,N_2647);
or U3067 (N_3067,N_2934,N_2830);
nand U3068 (N_3068,N_2831,N_2699);
xnor U3069 (N_3069,N_2694,N_2739);
xnor U3070 (N_3070,N_2961,N_2801);
or U3071 (N_3071,N_2907,N_2583);
and U3072 (N_3072,N_2981,N_2980);
nand U3073 (N_3073,N_2672,N_2888);
nand U3074 (N_3074,N_2651,N_2936);
or U3075 (N_3075,N_2722,N_2566);
nor U3076 (N_3076,N_2779,N_2767);
nand U3077 (N_3077,N_2776,N_2527);
nor U3078 (N_3078,N_2543,N_2992);
nand U3079 (N_3079,N_2790,N_2963);
xnor U3080 (N_3080,N_2796,N_2926);
nor U3081 (N_3081,N_2759,N_2911);
nor U3082 (N_3082,N_2948,N_2514);
xnor U3083 (N_3083,N_2999,N_2919);
nor U3084 (N_3084,N_2945,N_2847);
xor U3085 (N_3085,N_2837,N_2557);
and U3086 (N_3086,N_2858,N_2758);
nand U3087 (N_3087,N_2626,N_2815);
nor U3088 (N_3088,N_2808,N_2713);
or U3089 (N_3089,N_2838,N_2502);
xnor U3090 (N_3090,N_2881,N_2656);
and U3091 (N_3091,N_2889,N_2601);
nor U3092 (N_3092,N_2971,N_2662);
xnor U3093 (N_3093,N_2683,N_2855);
or U3094 (N_3094,N_2695,N_2978);
or U3095 (N_3095,N_2678,N_2620);
xor U3096 (N_3096,N_2615,N_2604);
nand U3097 (N_3097,N_2955,N_2795);
and U3098 (N_3098,N_2941,N_2768);
or U3099 (N_3099,N_2891,N_2664);
nand U3100 (N_3100,N_2588,N_2802);
nand U3101 (N_3101,N_2827,N_2500);
or U3102 (N_3102,N_2687,N_2915);
nor U3103 (N_3103,N_2825,N_2803);
or U3104 (N_3104,N_2928,N_2580);
or U3105 (N_3105,N_2535,N_2910);
nand U3106 (N_3106,N_2947,N_2977);
or U3107 (N_3107,N_2972,N_2732);
or U3108 (N_3108,N_2635,N_2600);
and U3109 (N_3109,N_2602,N_2964);
and U3110 (N_3110,N_2987,N_2772);
nor U3111 (N_3111,N_2507,N_2922);
xor U3112 (N_3112,N_2529,N_2567);
nand U3113 (N_3113,N_2784,N_2781);
and U3114 (N_3114,N_2637,N_2671);
nand U3115 (N_3115,N_2551,N_2581);
and U3116 (N_3116,N_2813,N_2986);
or U3117 (N_3117,N_2523,N_2900);
nor U3118 (N_3118,N_2940,N_2515);
nand U3119 (N_3119,N_2863,N_2917);
and U3120 (N_3120,N_2598,N_2693);
xor U3121 (N_3121,N_2913,N_2973);
and U3122 (N_3122,N_2621,N_2610);
nor U3123 (N_3123,N_2786,N_2669);
nor U3124 (N_3124,N_2872,N_2870);
nor U3125 (N_3125,N_2859,N_2544);
nand U3126 (N_3126,N_2599,N_2750);
xor U3127 (N_3127,N_2718,N_2841);
and U3128 (N_3128,N_2785,N_2522);
and U3129 (N_3129,N_2959,N_2503);
nor U3130 (N_3130,N_2655,N_2569);
and U3131 (N_3131,N_2818,N_2532);
nor U3132 (N_3132,N_2643,N_2904);
nand U3133 (N_3133,N_2840,N_2799);
xor U3134 (N_3134,N_2867,N_2704);
nand U3135 (N_3135,N_2578,N_2686);
nand U3136 (N_3136,N_2924,N_2593);
nor U3137 (N_3137,N_2794,N_2682);
nor U3138 (N_3138,N_2806,N_2614);
and U3139 (N_3139,N_2873,N_2773);
or U3140 (N_3140,N_2556,N_2866);
xor U3141 (N_3141,N_2616,N_2533);
xor U3142 (N_3142,N_2534,N_2688);
nand U3143 (N_3143,N_2909,N_2932);
and U3144 (N_3144,N_2636,N_2916);
or U3145 (N_3145,N_2712,N_2852);
and U3146 (N_3146,N_2542,N_2793);
or U3147 (N_3147,N_2937,N_2520);
or U3148 (N_3148,N_2550,N_2735);
or U3149 (N_3149,N_2778,N_2539);
nand U3150 (N_3150,N_2849,N_2510);
and U3151 (N_3151,N_2899,N_2920);
nor U3152 (N_3152,N_2822,N_2553);
nand U3153 (N_3153,N_2819,N_2777);
nand U3154 (N_3154,N_2974,N_2517);
xnor U3155 (N_3155,N_2625,N_2877);
and U3156 (N_3156,N_2708,N_2646);
and U3157 (N_3157,N_2748,N_2561);
and U3158 (N_3158,N_2879,N_2690);
nor U3159 (N_3159,N_2568,N_2518);
nand U3160 (N_3160,N_2611,N_2729);
nor U3161 (N_3161,N_2902,N_2575);
nor U3162 (N_3162,N_2757,N_2631);
and U3163 (N_3163,N_2876,N_2711);
nor U3164 (N_3164,N_2893,N_2956);
nor U3165 (N_3165,N_2853,N_2511);
nand U3166 (N_3166,N_2856,N_2942);
and U3167 (N_3167,N_2668,N_2512);
or U3168 (N_3168,N_2746,N_2605);
xnor U3169 (N_3169,N_2608,N_2887);
nor U3170 (N_3170,N_2528,N_2573);
nand U3171 (N_3171,N_2740,N_2714);
nand U3172 (N_3172,N_2680,N_2639);
nor U3173 (N_3173,N_2797,N_2737);
nor U3174 (N_3174,N_2659,N_2501);
or U3175 (N_3175,N_2787,N_2851);
xor U3176 (N_3176,N_2627,N_2912);
and U3177 (N_3177,N_2816,N_2555);
xnor U3178 (N_3178,N_2726,N_2597);
or U3179 (N_3179,N_2769,N_2731);
nor U3180 (N_3180,N_2882,N_2798);
nor U3181 (N_3181,N_2649,N_2696);
or U3182 (N_3182,N_2842,N_2905);
xnor U3183 (N_3183,N_2632,N_2541);
nor U3184 (N_3184,N_2571,N_2692);
or U3185 (N_3185,N_2939,N_2607);
nor U3186 (N_3186,N_2962,N_2957);
or U3187 (N_3187,N_2530,N_2861);
xnor U3188 (N_3188,N_2783,N_2812);
xor U3189 (N_3189,N_2946,N_2923);
nor U3190 (N_3190,N_2997,N_2716);
nand U3191 (N_3191,N_2698,N_2666);
or U3192 (N_3192,N_2775,N_2504);
nand U3193 (N_3193,N_2558,N_2587);
nand U3194 (N_3194,N_2976,N_2874);
nand U3195 (N_3195,N_2765,N_2612);
nor U3196 (N_3196,N_2592,N_2890);
or U3197 (N_3197,N_2613,N_2901);
nand U3198 (N_3198,N_2552,N_2660);
nand U3199 (N_3199,N_2549,N_2994);
nor U3200 (N_3200,N_2744,N_2800);
nand U3201 (N_3201,N_2829,N_2546);
nand U3202 (N_3202,N_2982,N_2789);
nand U3203 (N_3203,N_2702,N_2673);
nand U3204 (N_3204,N_2969,N_2574);
nor U3205 (N_3205,N_2938,N_2952);
nand U3206 (N_3206,N_2883,N_2895);
or U3207 (N_3207,N_2594,N_2848);
and U3208 (N_3208,N_2766,N_2880);
or U3209 (N_3209,N_2684,N_2547);
and U3210 (N_3210,N_2629,N_2700);
or U3211 (N_3211,N_2623,N_2654);
nor U3212 (N_3212,N_2706,N_2584);
nor U3213 (N_3213,N_2674,N_2807);
and U3214 (N_3214,N_2897,N_2998);
and U3215 (N_3215,N_2685,N_2989);
or U3216 (N_3216,N_2705,N_2967);
or U3217 (N_3217,N_2741,N_2619);
nand U3218 (N_3218,N_2835,N_2697);
and U3219 (N_3219,N_2509,N_2756);
xor U3220 (N_3220,N_2677,N_2828);
nor U3221 (N_3221,N_2990,N_2749);
and U3222 (N_3222,N_2886,N_2644);
or U3223 (N_3223,N_2931,N_2630);
or U3224 (N_3224,N_2665,N_2516);
nor U3225 (N_3225,N_2582,N_2991);
and U3226 (N_3226,N_2780,N_2983);
xor U3227 (N_3227,N_2526,N_2564);
nand U3228 (N_3228,N_2814,N_2679);
nand U3229 (N_3229,N_2958,N_2960);
and U3230 (N_3230,N_2823,N_2854);
xnor U3231 (N_3231,N_2914,N_2834);
or U3232 (N_3232,N_2884,N_2670);
and U3233 (N_3233,N_2954,N_2925);
xor U3234 (N_3234,N_2868,N_2531);
xor U3235 (N_3235,N_2570,N_2524);
nand U3236 (N_3236,N_2944,N_2753);
nand U3237 (N_3237,N_2707,N_2560);
nor U3238 (N_3238,N_2710,N_2715);
nor U3239 (N_3239,N_2843,N_2975);
nor U3240 (N_3240,N_2721,N_2894);
nand U3241 (N_3241,N_2865,N_2591);
or U3242 (N_3242,N_2933,N_2950);
and U3243 (N_3243,N_2995,N_2809);
or U3244 (N_3244,N_2820,N_2918);
nor U3245 (N_3245,N_2993,N_2742);
nand U3246 (N_3246,N_2755,N_2586);
or U3247 (N_3247,N_2857,N_2845);
nand U3248 (N_3248,N_2725,N_2579);
nor U3249 (N_3249,N_2824,N_2648);
nand U3250 (N_3250,N_2866,N_2790);
and U3251 (N_3251,N_2501,N_2601);
xor U3252 (N_3252,N_2668,N_2704);
or U3253 (N_3253,N_2607,N_2516);
and U3254 (N_3254,N_2574,N_2800);
or U3255 (N_3255,N_2854,N_2920);
and U3256 (N_3256,N_2753,N_2931);
and U3257 (N_3257,N_2513,N_2672);
and U3258 (N_3258,N_2561,N_2955);
xnor U3259 (N_3259,N_2544,N_2865);
nand U3260 (N_3260,N_2621,N_2738);
nor U3261 (N_3261,N_2556,N_2954);
nor U3262 (N_3262,N_2504,N_2782);
and U3263 (N_3263,N_2974,N_2629);
or U3264 (N_3264,N_2806,N_2825);
or U3265 (N_3265,N_2804,N_2992);
nand U3266 (N_3266,N_2508,N_2852);
and U3267 (N_3267,N_2840,N_2525);
xor U3268 (N_3268,N_2901,N_2953);
nand U3269 (N_3269,N_2984,N_2524);
and U3270 (N_3270,N_2714,N_2889);
or U3271 (N_3271,N_2846,N_2894);
nor U3272 (N_3272,N_2639,N_2953);
and U3273 (N_3273,N_2815,N_2585);
xnor U3274 (N_3274,N_2675,N_2912);
and U3275 (N_3275,N_2604,N_2922);
nor U3276 (N_3276,N_2993,N_2838);
nand U3277 (N_3277,N_2964,N_2980);
nand U3278 (N_3278,N_2539,N_2692);
nor U3279 (N_3279,N_2596,N_2982);
nand U3280 (N_3280,N_2957,N_2773);
or U3281 (N_3281,N_2986,N_2676);
xnor U3282 (N_3282,N_2899,N_2672);
nand U3283 (N_3283,N_2737,N_2823);
and U3284 (N_3284,N_2690,N_2872);
nand U3285 (N_3285,N_2649,N_2986);
and U3286 (N_3286,N_2963,N_2859);
or U3287 (N_3287,N_2546,N_2947);
nor U3288 (N_3288,N_2808,N_2811);
and U3289 (N_3289,N_2660,N_2721);
xor U3290 (N_3290,N_2914,N_2828);
and U3291 (N_3291,N_2681,N_2744);
or U3292 (N_3292,N_2762,N_2957);
nand U3293 (N_3293,N_2663,N_2656);
nand U3294 (N_3294,N_2941,N_2661);
or U3295 (N_3295,N_2505,N_2778);
nand U3296 (N_3296,N_2841,N_2688);
nor U3297 (N_3297,N_2924,N_2509);
nand U3298 (N_3298,N_2605,N_2513);
nand U3299 (N_3299,N_2714,N_2618);
or U3300 (N_3300,N_2685,N_2742);
and U3301 (N_3301,N_2652,N_2882);
or U3302 (N_3302,N_2953,N_2726);
nor U3303 (N_3303,N_2584,N_2896);
and U3304 (N_3304,N_2890,N_2976);
nand U3305 (N_3305,N_2854,N_2822);
or U3306 (N_3306,N_2931,N_2517);
or U3307 (N_3307,N_2745,N_2540);
and U3308 (N_3308,N_2521,N_2509);
or U3309 (N_3309,N_2534,N_2744);
or U3310 (N_3310,N_2609,N_2627);
nor U3311 (N_3311,N_2578,N_2558);
and U3312 (N_3312,N_2514,N_2728);
or U3313 (N_3313,N_2662,N_2773);
or U3314 (N_3314,N_2823,N_2688);
nand U3315 (N_3315,N_2664,N_2934);
or U3316 (N_3316,N_2888,N_2958);
and U3317 (N_3317,N_2629,N_2650);
nand U3318 (N_3318,N_2637,N_2665);
nor U3319 (N_3319,N_2539,N_2742);
nor U3320 (N_3320,N_2906,N_2884);
and U3321 (N_3321,N_2514,N_2819);
and U3322 (N_3322,N_2599,N_2954);
or U3323 (N_3323,N_2989,N_2868);
nor U3324 (N_3324,N_2803,N_2714);
or U3325 (N_3325,N_2650,N_2607);
nand U3326 (N_3326,N_2737,N_2770);
xnor U3327 (N_3327,N_2855,N_2801);
nor U3328 (N_3328,N_2516,N_2789);
nor U3329 (N_3329,N_2884,N_2933);
nand U3330 (N_3330,N_2920,N_2913);
nand U3331 (N_3331,N_2691,N_2663);
nand U3332 (N_3332,N_2555,N_2941);
nor U3333 (N_3333,N_2671,N_2830);
nand U3334 (N_3334,N_2657,N_2824);
and U3335 (N_3335,N_2795,N_2834);
or U3336 (N_3336,N_2833,N_2975);
or U3337 (N_3337,N_2849,N_2998);
or U3338 (N_3338,N_2699,N_2512);
nor U3339 (N_3339,N_2888,N_2996);
and U3340 (N_3340,N_2898,N_2561);
and U3341 (N_3341,N_2690,N_2747);
and U3342 (N_3342,N_2678,N_2888);
xor U3343 (N_3343,N_2724,N_2927);
or U3344 (N_3344,N_2825,N_2807);
nor U3345 (N_3345,N_2914,N_2821);
and U3346 (N_3346,N_2573,N_2588);
or U3347 (N_3347,N_2591,N_2879);
nand U3348 (N_3348,N_2721,N_2759);
and U3349 (N_3349,N_2876,N_2868);
nor U3350 (N_3350,N_2842,N_2729);
nand U3351 (N_3351,N_2901,N_2839);
or U3352 (N_3352,N_2986,N_2781);
nand U3353 (N_3353,N_2902,N_2562);
and U3354 (N_3354,N_2714,N_2762);
xor U3355 (N_3355,N_2802,N_2540);
nor U3356 (N_3356,N_2873,N_2669);
nor U3357 (N_3357,N_2594,N_2879);
nand U3358 (N_3358,N_2748,N_2932);
and U3359 (N_3359,N_2537,N_2644);
and U3360 (N_3360,N_2758,N_2734);
or U3361 (N_3361,N_2862,N_2509);
nor U3362 (N_3362,N_2797,N_2745);
and U3363 (N_3363,N_2537,N_2865);
nand U3364 (N_3364,N_2642,N_2860);
nor U3365 (N_3365,N_2847,N_2929);
and U3366 (N_3366,N_2741,N_2802);
nand U3367 (N_3367,N_2836,N_2930);
or U3368 (N_3368,N_2769,N_2579);
nor U3369 (N_3369,N_2963,N_2941);
and U3370 (N_3370,N_2606,N_2793);
or U3371 (N_3371,N_2501,N_2984);
nor U3372 (N_3372,N_2899,N_2935);
and U3373 (N_3373,N_2885,N_2705);
nand U3374 (N_3374,N_2989,N_2959);
and U3375 (N_3375,N_2867,N_2607);
and U3376 (N_3376,N_2779,N_2817);
nor U3377 (N_3377,N_2573,N_2993);
or U3378 (N_3378,N_2708,N_2928);
nor U3379 (N_3379,N_2947,N_2886);
or U3380 (N_3380,N_2777,N_2767);
nor U3381 (N_3381,N_2927,N_2792);
nor U3382 (N_3382,N_2606,N_2516);
nor U3383 (N_3383,N_2811,N_2628);
and U3384 (N_3384,N_2920,N_2647);
and U3385 (N_3385,N_2988,N_2671);
nor U3386 (N_3386,N_2881,N_2738);
or U3387 (N_3387,N_2865,N_2561);
and U3388 (N_3388,N_2542,N_2720);
or U3389 (N_3389,N_2618,N_2889);
or U3390 (N_3390,N_2670,N_2930);
or U3391 (N_3391,N_2715,N_2716);
and U3392 (N_3392,N_2647,N_2820);
and U3393 (N_3393,N_2619,N_2531);
or U3394 (N_3394,N_2645,N_2750);
or U3395 (N_3395,N_2656,N_2963);
or U3396 (N_3396,N_2949,N_2749);
nand U3397 (N_3397,N_2707,N_2747);
nor U3398 (N_3398,N_2566,N_2578);
and U3399 (N_3399,N_2909,N_2740);
nand U3400 (N_3400,N_2527,N_2553);
nor U3401 (N_3401,N_2504,N_2532);
and U3402 (N_3402,N_2600,N_2519);
xnor U3403 (N_3403,N_2568,N_2923);
nor U3404 (N_3404,N_2533,N_2886);
or U3405 (N_3405,N_2895,N_2733);
nand U3406 (N_3406,N_2666,N_2706);
nor U3407 (N_3407,N_2913,N_2722);
and U3408 (N_3408,N_2875,N_2885);
nor U3409 (N_3409,N_2765,N_2768);
and U3410 (N_3410,N_2849,N_2734);
and U3411 (N_3411,N_2617,N_2663);
nand U3412 (N_3412,N_2958,N_2804);
nand U3413 (N_3413,N_2525,N_2941);
nor U3414 (N_3414,N_2878,N_2742);
or U3415 (N_3415,N_2995,N_2771);
nor U3416 (N_3416,N_2863,N_2736);
nor U3417 (N_3417,N_2853,N_2908);
and U3418 (N_3418,N_2966,N_2631);
nand U3419 (N_3419,N_2642,N_2947);
xnor U3420 (N_3420,N_2615,N_2955);
and U3421 (N_3421,N_2720,N_2610);
nor U3422 (N_3422,N_2700,N_2540);
or U3423 (N_3423,N_2694,N_2566);
nor U3424 (N_3424,N_2592,N_2787);
or U3425 (N_3425,N_2789,N_2632);
xor U3426 (N_3426,N_2892,N_2593);
nand U3427 (N_3427,N_2507,N_2608);
nor U3428 (N_3428,N_2828,N_2682);
nand U3429 (N_3429,N_2560,N_2597);
nor U3430 (N_3430,N_2862,N_2810);
or U3431 (N_3431,N_2725,N_2524);
nor U3432 (N_3432,N_2929,N_2631);
and U3433 (N_3433,N_2646,N_2946);
or U3434 (N_3434,N_2607,N_2618);
xor U3435 (N_3435,N_2907,N_2680);
xnor U3436 (N_3436,N_2983,N_2811);
or U3437 (N_3437,N_2843,N_2592);
nor U3438 (N_3438,N_2704,N_2657);
nand U3439 (N_3439,N_2925,N_2986);
nor U3440 (N_3440,N_2880,N_2665);
and U3441 (N_3441,N_2561,N_2820);
and U3442 (N_3442,N_2527,N_2970);
xnor U3443 (N_3443,N_2589,N_2611);
and U3444 (N_3444,N_2584,N_2723);
and U3445 (N_3445,N_2807,N_2519);
xnor U3446 (N_3446,N_2605,N_2514);
and U3447 (N_3447,N_2807,N_2831);
xnor U3448 (N_3448,N_2589,N_2945);
or U3449 (N_3449,N_2665,N_2563);
or U3450 (N_3450,N_2541,N_2968);
or U3451 (N_3451,N_2842,N_2761);
nor U3452 (N_3452,N_2583,N_2910);
nor U3453 (N_3453,N_2899,N_2786);
nor U3454 (N_3454,N_2731,N_2925);
and U3455 (N_3455,N_2899,N_2732);
nor U3456 (N_3456,N_2502,N_2756);
xnor U3457 (N_3457,N_2824,N_2985);
nand U3458 (N_3458,N_2663,N_2944);
nor U3459 (N_3459,N_2594,N_2668);
nand U3460 (N_3460,N_2721,N_2749);
and U3461 (N_3461,N_2742,N_2805);
xnor U3462 (N_3462,N_2653,N_2801);
and U3463 (N_3463,N_2548,N_2885);
and U3464 (N_3464,N_2760,N_2612);
and U3465 (N_3465,N_2857,N_2834);
nor U3466 (N_3466,N_2736,N_2569);
xor U3467 (N_3467,N_2523,N_2708);
or U3468 (N_3468,N_2532,N_2811);
nor U3469 (N_3469,N_2729,N_2541);
nor U3470 (N_3470,N_2671,N_2992);
xor U3471 (N_3471,N_2572,N_2958);
xnor U3472 (N_3472,N_2825,N_2509);
and U3473 (N_3473,N_2720,N_2745);
nor U3474 (N_3474,N_2750,N_2639);
nand U3475 (N_3475,N_2990,N_2521);
or U3476 (N_3476,N_2913,N_2524);
nor U3477 (N_3477,N_2818,N_2688);
and U3478 (N_3478,N_2519,N_2591);
nand U3479 (N_3479,N_2554,N_2506);
nor U3480 (N_3480,N_2976,N_2705);
and U3481 (N_3481,N_2829,N_2664);
nand U3482 (N_3482,N_2686,N_2995);
nand U3483 (N_3483,N_2938,N_2715);
or U3484 (N_3484,N_2516,N_2561);
xor U3485 (N_3485,N_2794,N_2591);
nand U3486 (N_3486,N_2896,N_2711);
nand U3487 (N_3487,N_2546,N_2877);
nand U3488 (N_3488,N_2703,N_2710);
nand U3489 (N_3489,N_2867,N_2812);
and U3490 (N_3490,N_2719,N_2853);
or U3491 (N_3491,N_2930,N_2904);
and U3492 (N_3492,N_2613,N_2603);
xnor U3493 (N_3493,N_2594,N_2549);
or U3494 (N_3494,N_2871,N_2764);
or U3495 (N_3495,N_2894,N_2781);
or U3496 (N_3496,N_2908,N_2854);
nor U3497 (N_3497,N_2826,N_2853);
nor U3498 (N_3498,N_2762,N_2630);
nor U3499 (N_3499,N_2790,N_2869);
and U3500 (N_3500,N_3109,N_3251);
nand U3501 (N_3501,N_3355,N_3490);
and U3502 (N_3502,N_3450,N_3307);
nand U3503 (N_3503,N_3045,N_3051);
and U3504 (N_3504,N_3453,N_3137);
nor U3505 (N_3505,N_3023,N_3309);
nand U3506 (N_3506,N_3125,N_3236);
nand U3507 (N_3507,N_3310,N_3064);
or U3508 (N_3508,N_3448,N_3087);
and U3509 (N_3509,N_3094,N_3305);
nand U3510 (N_3510,N_3425,N_3092);
nor U3511 (N_3511,N_3267,N_3118);
nand U3512 (N_3512,N_3492,N_3391);
or U3513 (N_3513,N_3127,N_3122);
nand U3514 (N_3514,N_3286,N_3449);
nor U3515 (N_3515,N_3472,N_3046);
xor U3516 (N_3516,N_3254,N_3398);
nor U3517 (N_3517,N_3342,N_3083);
nand U3518 (N_3518,N_3006,N_3457);
nor U3519 (N_3519,N_3220,N_3435);
nor U3520 (N_3520,N_3481,N_3065);
xnor U3521 (N_3521,N_3404,N_3176);
xnor U3522 (N_3522,N_3390,N_3487);
nor U3523 (N_3523,N_3349,N_3119);
xor U3524 (N_3524,N_3243,N_3213);
and U3525 (N_3525,N_3356,N_3438);
and U3526 (N_3526,N_3173,N_3430);
xor U3527 (N_3527,N_3467,N_3299);
or U3528 (N_3528,N_3133,N_3460);
nor U3529 (N_3529,N_3334,N_3250);
and U3530 (N_3530,N_3016,N_3149);
or U3531 (N_3531,N_3145,N_3281);
or U3532 (N_3532,N_3297,N_3369);
and U3533 (N_3533,N_3190,N_3397);
and U3534 (N_3534,N_3270,N_3290);
nor U3535 (N_3535,N_3104,N_3249);
nor U3536 (N_3536,N_3107,N_3372);
and U3537 (N_3537,N_3429,N_3135);
nor U3538 (N_3538,N_3001,N_3382);
or U3539 (N_3539,N_3423,N_3366);
and U3540 (N_3540,N_3395,N_3204);
and U3541 (N_3541,N_3143,N_3141);
nor U3542 (N_3542,N_3099,N_3353);
xnor U3543 (N_3543,N_3072,N_3150);
or U3544 (N_3544,N_3033,N_3209);
or U3545 (N_3545,N_3496,N_3234);
nand U3546 (N_3546,N_3055,N_3217);
or U3547 (N_3547,N_3362,N_3185);
nand U3548 (N_3548,N_3462,N_3383);
and U3549 (N_3549,N_3428,N_3218);
nand U3550 (N_3550,N_3322,N_3073);
xnor U3551 (N_3551,N_3255,N_3017);
nand U3552 (N_3552,N_3455,N_3483);
or U3553 (N_3553,N_3189,N_3000);
nand U3554 (N_3554,N_3405,N_3288);
or U3555 (N_3555,N_3180,N_3028);
nor U3556 (N_3556,N_3002,N_3325);
nand U3557 (N_3557,N_3221,N_3205);
and U3558 (N_3558,N_3128,N_3308);
nor U3559 (N_3559,N_3193,N_3079);
xor U3560 (N_3560,N_3085,N_3163);
or U3561 (N_3561,N_3164,N_3203);
or U3562 (N_3562,N_3153,N_3461);
and U3563 (N_3563,N_3174,N_3178);
nand U3564 (N_3564,N_3371,N_3285);
nand U3565 (N_3565,N_3437,N_3088);
nand U3566 (N_3566,N_3486,N_3478);
and U3567 (N_3567,N_3054,N_3108);
nand U3568 (N_3568,N_3167,N_3413);
nand U3569 (N_3569,N_3060,N_3258);
or U3570 (N_3570,N_3191,N_3238);
and U3571 (N_3571,N_3129,N_3252);
nor U3572 (N_3572,N_3159,N_3080);
nor U3573 (N_3573,N_3186,N_3329);
nand U3574 (N_3574,N_3352,N_3420);
nor U3575 (N_3575,N_3379,N_3181);
nor U3576 (N_3576,N_3110,N_3296);
nand U3577 (N_3577,N_3284,N_3476);
nor U3578 (N_3578,N_3452,N_3412);
and U3579 (N_3579,N_3264,N_3009);
and U3580 (N_3580,N_3008,N_3061);
or U3581 (N_3581,N_3260,N_3302);
or U3582 (N_3582,N_3050,N_3123);
or U3583 (N_3583,N_3196,N_3484);
nor U3584 (N_3584,N_3120,N_3097);
or U3585 (N_3585,N_3439,N_3059);
nor U3586 (N_3586,N_3315,N_3426);
and U3587 (N_3587,N_3199,N_3084);
nand U3588 (N_3588,N_3364,N_3465);
xnor U3589 (N_3589,N_3126,N_3374);
or U3590 (N_3590,N_3078,N_3346);
nor U3591 (N_3591,N_3007,N_3049);
nor U3592 (N_3592,N_3134,N_3067);
and U3593 (N_3593,N_3479,N_3227);
nor U3594 (N_3594,N_3338,N_3081);
and U3595 (N_3595,N_3106,N_3259);
xnor U3596 (N_3596,N_3313,N_3187);
nand U3597 (N_3597,N_3222,N_3376);
nand U3598 (N_3598,N_3136,N_3231);
or U3599 (N_3599,N_3339,N_3406);
and U3600 (N_3600,N_3074,N_3387);
nand U3601 (N_3601,N_3032,N_3370);
and U3602 (N_3602,N_3410,N_3021);
nand U3603 (N_3603,N_3433,N_3330);
nor U3604 (N_3604,N_3161,N_3323);
nor U3605 (N_3605,N_3044,N_3424);
nand U3606 (N_3606,N_3361,N_3034);
nor U3607 (N_3607,N_3066,N_3399);
nor U3608 (N_3608,N_3321,N_3022);
xor U3609 (N_3609,N_3229,N_3169);
or U3610 (N_3610,N_3151,N_3377);
nor U3611 (N_3611,N_3202,N_3077);
nor U3612 (N_3612,N_3131,N_3152);
xnor U3613 (N_3613,N_3351,N_3058);
nand U3614 (N_3614,N_3068,N_3130);
or U3615 (N_3615,N_3183,N_3416);
nand U3616 (N_3616,N_3225,N_3385);
nand U3617 (N_3617,N_3324,N_3441);
nand U3618 (N_3618,N_3003,N_3272);
and U3619 (N_3619,N_3146,N_3027);
nand U3620 (N_3620,N_3367,N_3116);
nand U3621 (N_3621,N_3354,N_3473);
and U3622 (N_3622,N_3301,N_3115);
xnor U3623 (N_3623,N_3240,N_3262);
nand U3624 (N_3624,N_3417,N_3112);
nand U3625 (N_3625,N_3482,N_3400);
or U3626 (N_3626,N_3306,N_3172);
or U3627 (N_3627,N_3014,N_3314);
nor U3628 (N_3628,N_3101,N_3155);
nor U3629 (N_3629,N_3269,N_3341);
and U3630 (N_3630,N_3095,N_3247);
nor U3631 (N_3631,N_3018,N_3408);
or U3632 (N_3632,N_3442,N_3241);
and U3633 (N_3633,N_3117,N_3091);
nor U3634 (N_3634,N_3237,N_3257);
or U3635 (N_3635,N_3344,N_3293);
and U3636 (N_3636,N_3265,N_3019);
nor U3637 (N_3637,N_3015,N_3332);
nand U3638 (N_3638,N_3347,N_3147);
and U3639 (N_3639,N_3357,N_3327);
or U3640 (N_3640,N_3138,N_3188);
nand U3641 (N_3641,N_3440,N_3303);
nand U3642 (N_3642,N_3024,N_3421);
nand U3643 (N_3643,N_3333,N_3170);
nor U3644 (N_3644,N_3274,N_3025);
nor U3645 (N_3645,N_3069,N_3498);
nand U3646 (N_3646,N_3194,N_3200);
or U3647 (N_3647,N_3226,N_3463);
or U3648 (N_3648,N_3156,N_3335);
and U3649 (N_3649,N_3298,N_3171);
or U3650 (N_3650,N_3402,N_3013);
nor U3651 (N_3651,N_3211,N_3488);
nand U3652 (N_3652,N_3300,N_3278);
xnor U3653 (N_3653,N_3010,N_3456);
nand U3654 (N_3654,N_3090,N_3312);
or U3655 (N_3655,N_3446,N_3020);
nand U3656 (N_3656,N_3223,N_3041);
nor U3657 (N_3657,N_3148,N_3244);
nor U3658 (N_3658,N_3468,N_3388);
nor U3659 (N_3659,N_3411,N_3418);
or U3660 (N_3660,N_3140,N_3228);
and U3661 (N_3661,N_3444,N_3063);
and U3662 (N_3662,N_3328,N_3319);
nand U3663 (N_3663,N_3294,N_3037);
nor U3664 (N_3664,N_3434,N_3132);
and U3665 (N_3665,N_3105,N_3389);
nand U3666 (N_3666,N_3160,N_3005);
nor U3667 (N_3667,N_3062,N_3039);
nor U3668 (N_3668,N_3485,N_3415);
nor U3669 (N_3669,N_3215,N_3057);
nand U3670 (N_3670,N_3098,N_3480);
or U3671 (N_3671,N_3497,N_3394);
nor U3672 (N_3672,N_3358,N_3076);
and U3673 (N_3673,N_3144,N_3071);
nand U3674 (N_3674,N_3012,N_3287);
and U3675 (N_3675,N_3266,N_3165);
or U3676 (N_3676,N_3275,N_3230);
or U3677 (N_3677,N_3340,N_3124);
xor U3678 (N_3678,N_3179,N_3053);
or U3679 (N_3679,N_3380,N_3245);
nor U3680 (N_3680,N_3477,N_3317);
and U3681 (N_3681,N_3184,N_3337);
nand U3682 (N_3682,N_3102,N_3409);
or U3683 (N_3683,N_3035,N_3304);
and U3684 (N_3684,N_3386,N_3168);
nand U3685 (N_3685,N_3121,N_3432);
nand U3686 (N_3686,N_3336,N_3447);
nand U3687 (N_3687,N_3375,N_3427);
and U3688 (N_3688,N_3192,N_3182);
nand U3689 (N_3689,N_3162,N_3224);
and U3690 (N_3690,N_3082,N_3212);
or U3691 (N_3691,N_3111,N_3026);
or U3692 (N_3692,N_3154,N_3295);
or U3693 (N_3693,N_3316,N_3198);
or U3694 (N_3694,N_3454,N_3318);
nor U3695 (N_3695,N_3175,N_3177);
nand U3696 (N_3696,N_3253,N_3403);
nor U3697 (N_3697,N_3443,N_3248);
xnor U3698 (N_3698,N_3029,N_3422);
nand U3699 (N_3699,N_3292,N_3139);
and U3700 (N_3700,N_3048,N_3232);
nor U3701 (N_3701,N_3239,N_3279);
nor U3702 (N_3702,N_3373,N_3384);
and U3703 (N_3703,N_3256,N_3036);
nor U3704 (N_3704,N_3469,N_3277);
nor U3705 (N_3705,N_3392,N_3038);
nor U3706 (N_3706,N_3363,N_3086);
and U3707 (N_3707,N_3093,N_3075);
and U3708 (N_3708,N_3445,N_3491);
or U3709 (N_3709,N_3089,N_3393);
or U3710 (N_3710,N_3206,N_3291);
nand U3711 (N_3711,N_3378,N_3381);
or U3712 (N_3712,N_3011,N_3464);
xnor U3713 (N_3713,N_3216,N_3365);
and U3714 (N_3714,N_3419,N_3004);
and U3715 (N_3715,N_3268,N_3368);
nand U3716 (N_3716,N_3396,N_3242);
nor U3717 (N_3717,N_3096,N_3458);
nand U3718 (N_3718,N_3345,N_3350);
or U3719 (N_3719,N_3436,N_3052);
and U3720 (N_3720,N_3401,N_3195);
xnor U3721 (N_3721,N_3114,N_3207);
or U3722 (N_3722,N_3348,N_3047);
or U3723 (N_3723,N_3495,N_3494);
or U3724 (N_3724,N_3280,N_3466);
nand U3725 (N_3725,N_3359,N_3201);
nor U3726 (N_3726,N_3031,N_3276);
nand U3727 (N_3727,N_3489,N_3493);
nor U3728 (N_3728,N_3459,N_3210);
nor U3729 (N_3729,N_3040,N_3070);
nand U3730 (N_3730,N_3414,N_3475);
nor U3731 (N_3731,N_3208,N_3214);
nand U3732 (N_3732,N_3311,N_3158);
or U3733 (N_3733,N_3282,N_3343);
and U3734 (N_3734,N_3271,N_3142);
nand U3735 (N_3735,N_3407,N_3360);
or U3736 (N_3736,N_3320,N_3326);
or U3737 (N_3737,N_3470,N_3103);
nor U3738 (N_3738,N_3261,N_3233);
nand U3739 (N_3739,N_3157,N_3166);
nor U3740 (N_3740,N_3030,N_3043);
nor U3741 (N_3741,N_3263,N_3451);
and U3742 (N_3742,N_3283,N_3499);
nand U3743 (N_3743,N_3246,N_3100);
and U3744 (N_3744,N_3331,N_3474);
nand U3745 (N_3745,N_3273,N_3219);
nor U3746 (N_3746,N_3289,N_3431);
nor U3747 (N_3747,N_3235,N_3471);
nor U3748 (N_3748,N_3197,N_3042);
or U3749 (N_3749,N_3113,N_3056);
xor U3750 (N_3750,N_3045,N_3313);
or U3751 (N_3751,N_3144,N_3352);
nand U3752 (N_3752,N_3008,N_3264);
nor U3753 (N_3753,N_3255,N_3116);
xor U3754 (N_3754,N_3337,N_3362);
xor U3755 (N_3755,N_3335,N_3267);
nor U3756 (N_3756,N_3492,N_3299);
or U3757 (N_3757,N_3085,N_3213);
and U3758 (N_3758,N_3298,N_3033);
nor U3759 (N_3759,N_3375,N_3227);
or U3760 (N_3760,N_3168,N_3466);
and U3761 (N_3761,N_3399,N_3184);
nor U3762 (N_3762,N_3494,N_3486);
or U3763 (N_3763,N_3026,N_3117);
or U3764 (N_3764,N_3226,N_3340);
or U3765 (N_3765,N_3150,N_3308);
nor U3766 (N_3766,N_3141,N_3204);
xor U3767 (N_3767,N_3069,N_3367);
nand U3768 (N_3768,N_3166,N_3030);
or U3769 (N_3769,N_3162,N_3157);
or U3770 (N_3770,N_3076,N_3021);
nand U3771 (N_3771,N_3384,N_3409);
nand U3772 (N_3772,N_3387,N_3354);
nor U3773 (N_3773,N_3445,N_3003);
nand U3774 (N_3774,N_3193,N_3428);
and U3775 (N_3775,N_3228,N_3483);
or U3776 (N_3776,N_3236,N_3431);
and U3777 (N_3777,N_3100,N_3024);
nand U3778 (N_3778,N_3413,N_3172);
nand U3779 (N_3779,N_3492,N_3496);
nor U3780 (N_3780,N_3291,N_3377);
nand U3781 (N_3781,N_3445,N_3243);
and U3782 (N_3782,N_3439,N_3020);
and U3783 (N_3783,N_3060,N_3046);
nand U3784 (N_3784,N_3386,N_3485);
nand U3785 (N_3785,N_3487,N_3336);
or U3786 (N_3786,N_3052,N_3368);
or U3787 (N_3787,N_3321,N_3185);
and U3788 (N_3788,N_3278,N_3459);
and U3789 (N_3789,N_3102,N_3061);
or U3790 (N_3790,N_3488,N_3176);
and U3791 (N_3791,N_3226,N_3257);
nand U3792 (N_3792,N_3294,N_3286);
nand U3793 (N_3793,N_3379,N_3430);
xor U3794 (N_3794,N_3371,N_3217);
or U3795 (N_3795,N_3076,N_3473);
and U3796 (N_3796,N_3231,N_3013);
and U3797 (N_3797,N_3037,N_3247);
and U3798 (N_3798,N_3395,N_3045);
and U3799 (N_3799,N_3028,N_3269);
nand U3800 (N_3800,N_3017,N_3454);
and U3801 (N_3801,N_3466,N_3459);
nor U3802 (N_3802,N_3228,N_3083);
nand U3803 (N_3803,N_3084,N_3067);
nor U3804 (N_3804,N_3189,N_3210);
nand U3805 (N_3805,N_3337,N_3219);
and U3806 (N_3806,N_3145,N_3327);
nand U3807 (N_3807,N_3361,N_3370);
nand U3808 (N_3808,N_3007,N_3078);
nand U3809 (N_3809,N_3160,N_3188);
nor U3810 (N_3810,N_3419,N_3145);
and U3811 (N_3811,N_3159,N_3004);
and U3812 (N_3812,N_3117,N_3371);
nor U3813 (N_3813,N_3441,N_3207);
and U3814 (N_3814,N_3070,N_3318);
or U3815 (N_3815,N_3180,N_3034);
xnor U3816 (N_3816,N_3072,N_3207);
nor U3817 (N_3817,N_3481,N_3191);
nor U3818 (N_3818,N_3133,N_3127);
nand U3819 (N_3819,N_3056,N_3317);
nand U3820 (N_3820,N_3284,N_3299);
nor U3821 (N_3821,N_3048,N_3421);
nor U3822 (N_3822,N_3421,N_3153);
nor U3823 (N_3823,N_3075,N_3295);
nand U3824 (N_3824,N_3450,N_3036);
nor U3825 (N_3825,N_3218,N_3293);
nand U3826 (N_3826,N_3044,N_3031);
and U3827 (N_3827,N_3236,N_3368);
nand U3828 (N_3828,N_3145,N_3340);
nor U3829 (N_3829,N_3140,N_3119);
nand U3830 (N_3830,N_3026,N_3311);
and U3831 (N_3831,N_3116,N_3457);
or U3832 (N_3832,N_3389,N_3097);
nand U3833 (N_3833,N_3136,N_3293);
and U3834 (N_3834,N_3003,N_3461);
and U3835 (N_3835,N_3266,N_3091);
xnor U3836 (N_3836,N_3485,N_3296);
xor U3837 (N_3837,N_3414,N_3127);
nand U3838 (N_3838,N_3049,N_3130);
nor U3839 (N_3839,N_3425,N_3440);
nand U3840 (N_3840,N_3406,N_3462);
nor U3841 (N_3841,N_3060,N_3423);
and U3842 (N_3842,N_3159,N_3364);
nand U3843 (N_3843,N_3086,N_3426);
xnor U3844 (N_3844,N_3029,N_3296);
nand U3845 (N_3845,N_3073,N_3057);
or U3846 (N_3846,N_3339,N_3229);
or U3847 (N_3847,N_3130,N_3103);
and U3848 (N_3848,N_3326,N_3055);
or U3849 (N_3849,N_3286,N_3219);
and U3850 (N_3850,N_3057,N_3497);
or U3851 (N_3851,N_3306,N_3330);
nand U3852 (N_3852,N_3079,N_3187);
and U3853 (N_3853,N_3210,N_3336);
xor U3854 (N_3854,N_3244,N_3334);
nand U3855 (N_3855,N_3338,N_3454);
nand U3856 (N_3856,N_3409,N_3423);
or U3857 (N_3857,N_3395,N_3396);
nor U3858 (N_3858,N_3486,N_3463);
and U3859 (N_3859,N_3216,N_3165);
or U3860 (N_3860,N_3013,N_3285);
and U3861 (N_3861,N_3136,N_3131);
nor U3862 (N_3862,N_3123,N_3472);
or U3863 (N_3863,N_3354,N_3358);
nor U3864 (N_3864,N_3408,N_3470);
nor U3865 (N_3865,N_3078,N_3031);
or U3866 (N_3866,N_3041,N_3195);
nor U3867 (N_3867,N_3388,N_3240);
nand U3868 (N_3868,N_3446,N_3379);
nor U3869 (N_3869,N_3263,N_3494);
xor U3870 (N_3870,N_3117,N_3249);
and U3871 (N_3871,N_3115,N_3481);
nand U3872 (N_3872,N_3216,N_3076);
nand U3873 (N_3873,N_3165,N_3128);
nand U3874 (N_3874,N_3098,N_3269);
nand U3875 (N_3875,N_3439,N_3157);
or U3876 (N_3876,N_3209,N_3390);
and U3877 (N_3877,N_3393,N_3378);
nand U3878 (N_3878,N_3085,N_3403);
or U3879 (N_3879,N_3188,N_3174);
nor U3880 (N_3880,N_3128,N_3224);
nor U3881 (N_3881,N_3231,N_3456);
or U3882 (N_3882,N_3491,N_3192);
nand U3883 (N_3883,N_3426,N_3406);
nand U3884 (N_3884,N_3322,N_3282);
or U3885 (N_3885,N_3091,N_3201);
nand U3886 (N_3886,N_3195,N_3069);
or U3887 (N_3887,N_3274,N_3075);
or U3888 (N_3888,N_3210,N_3000);
and U3889 (N_3889,N_3319,N_3406);
xnor U3890 (N_3890,N_3195,N_3306);
xnor U3891 (N_3891,N_3353,N_3334);
nand U3892 (N_3892,N_3318,N_3365);
or U3893 (N_3893,N_3349,N_3309);
nor U3894 (N_3894,N_3042,N_3199);
nand U3895 (N_3895,N_3464,N_3496);
nor U3896 (N_3896,N_3046,N_3304);
nand U3897 (N_3897,N_3211,N_3214);
nand U3898 (N_3898,N_3103,N_3242);
or U3899 (N_3899,N_3491,N_3322);
and U3900 (N_3900,N_3121,N_3426);
or U3901 (N_3901,N_3409,N_3319);
or U3902 (N_3902,N_3290,N_3117);
or U3903 (N_3903,N_3014,N_3291);
nand U3904 (N_3904,N_3403,N_3298);
nor U3905 (N_3905,N_3037,N_3166);
and U3906 (N_3906,N_3111,N_3327);
or U3907 (N_3907,N_3486,N_3261);
or U3908 (N_3908,N_3100,N_3241);
or U3909 (N_3909,N_3135,N_3383);
nor U3910 (N_3910,N_3225,N_3084);
and U3911 (N_3911,N_3259,N_3286);
nor U3912 (N_3912,N_3152,N_3381);
nor U3913 (N_3913,N_3129,N_3361);
or U3914 (N_3914,N_3404,N_3030);
or U3915 (N_3915,N_3108,N_3069);
nor U3916 (N_3916,N_3078,N_3491);
or U3917 (N_3917,N_3369,N_3348);
nand U3918 (N_3918,N_3282,N_3223);
xor U3919 (N_3919,N_3374,N_3002);
or U3920 (N_3920,N_3338,N_3403);
nand U3921 (N_3921,N_3481,N_3175);
and U3922 (N_3922,N_3337,N_3307);
nor U3923 (N_3923,N_3055,N_3005);
and U3924 (N_3924,N_3115,N_3475);
and U3925 (N_3925,N_3012,N_3106);
nor U3926 (N_3926,N_3442,N_3164);
and U3927 (N_3927,N_3141,N_3479);
and U3928 (N_3928,N_3491,N_3304);
xnor U3929 (N_3929,N_3264,N_3303);
or U3930 (N_3930,N_3017,N_3124);
and U3931 (N_3931,N_3299,N_3460);
nand U3932 (N_3932,N_3228,N_3396);
nand U3933 (N_3933,N_3469,N_3112);
or U3934 (N_3934,N_3295,N_3318);
or U3935 (N_3935,N_3337,N_3196);
nor U3936 (N_3936,N_3275,N_3000);
and U3937 (N_3937,N_3451,N_3362);
and U3938 (N_3938,N_3320,N_3178);
or U3939 (N_3939,N_3247,N_3380);
nor U3940 (N_3940,N_3238,N_3464);
or U3941 (N_3941,N_3390,N_3004);
xor U3942 (N_3942,N_3346,N_3349);
or U3943 (N_3943,N_3386,N_3132);
nor U3944 (N_3944,N_3004,N_3391);
nand U3945 (N_3945,N_3478,N_3022);
and U3946 (N_3946,N_3221,N_3213);
and U3947 (N_3947,N_3307,N_3490);
nand U3948 (N_3948,N_3278,N_3372);
and U3949 (N_3949,N_3032,N_3173);
nand U3950 (N_3950,N_3219,N_3200);
nand U3951 (N_3951,N_3370,N_3377);
xnor U3952 (N_3952,N_3164,N_3272);
nand U3953 (N_3953,N_3403,N_3359);
and U3954 (N_3954,N_3277,N_3019);
or U3955 (N_3955,N_3468,N_3029);
xnor U3956 (N_3956,N_3306,N_3217);
or U3957 (N_3957,N_3262,N_3102);
nand U3958 (N_3958,N_3356,N_3330);
nor U3959 (N_3959,N_3255,N_3419);
nand U3960 (N_3960,N_3358,N_3339);
or U3961 (N_3961,N_3438,N_3118);
and U3962 (N_3962,N_3221,N_3232);
and U3963 (N_3963,N_3252,N_3024);
and U3964 (N_3964,N_3413,N_3226);
nor U3965 (N_3965,N_3260,N_3077);
nand U3966 (N_3966,N_3075,N_3184);
xnor U3967 (N_3967,N_3390,N_3326);
or U3968 (N_3968,N_3128,N_3269);
nor U3969 (N_3969,N_3402,N_3354);
or U3970 (N_3970,N_3021,N_3190);
or U3971 (N_3971,N_3122,N_3207);
nand U3972 (N_3972,N_3461,N_3146);
nor U3973 (N_3973,N_3006,N_3035);
nand U3974 (N_3974,N_3159,N_3398);
or U3975 (N_3975,N_3320,N_3148);
or U3976 (N_3976,N_3019,N_3031);
and U3977 (N_3977,N_3212,N_3200);
or U3978 (N_3978,N_3403,N_3344);
nand U3979 (N_3979,N_3333,N_3211);
nor U3980 (N_3980,N_3485,N_3171);
xnor U3981 (N_3981,N_3325,N_3206);
and U3982 (N_3982,N_3015,N_3058);
and U3983 (N_3983,N_3376,N_3231);
xnor U3984 (N_3984,N_3156,N_3350);
nor U3985 (N_3985,N_3375,N_3402);
nor U3986 (N_3986,N_3459,N_3024);
nor U3987 (N_3987,N_3155,N_3419);
nor U3988 (N_3988,N_3254,N_3363);
or U3989 (N_3989,N_3394,N_3253);
nand U3990 (N_3990,N_3237,N_3311);
and U3991 (N_3991,N_3124,N_3143);
nand U3992 (N_3992,N_3201,N_3398);
nor U3993 (N_3993,N_3336,N_3361);
or U3994 (N_3994,N_3371,N_3421);
and U3995 (N_3995,N_3279,N_3003);
nand U3996 (N_3996,N_3135,N_3086);
xor U3997 (N_3997,N_3027,N_3141);
or U3998 (N_3998,N_3282,N_3096);
nor U3999 (N_3999,N_3326,N_3309);
and U4000 (N_4000,N_3785,N_3834);
or U4001 (N_4001,N_3841,N_3822);
or U4002 (N_4002,N_3738,N_3883);
or U4003 (N_4003,N_3763,N_3908);
or U4004 (N_4004,N_3772,N_3682);
nor U4005 (N_4005,N_3629,N_3793);
or U4006 (N_4006,N_3791,N_3639);
nor U4007 (N_4007,N_3992,N_3511);
xor U4008 (N_4008,N_3860,N_3650);
or U4009 (N_4009,N_3741,N_3565);
nor U4010 (N_4010,N_3573,N_3951);
nor U4011 (N_4011,N_3576,N_3878);
nor U4012 (N_4012,N_3669,N_3646);
nand U4013 (N_4013,N_3588,N_3892);
nor U4014 (N_4014,N_3675,N_3854);
or U4015 (N_4015,N_3950,N_3911);
xor U4016 (N_4016,N_3631,N_3971);
xnor U4017 (N_4017,N_3527,N_3605);
nand U4018 (N_4018,N_3759,N_3616);
and U4019 (N_4019,N_3811,N_3641);
and U4020 (N_4020,N_3798,N_3945);
nand U4021 (N_4021,N_3940,N_3555);
or U4022 (N_4022,N_3550,N_3640);
nand U4023 (N_4023,N_3962,N_3916);
or U4024 (N_4024,N_3683,N_3899);
xnor U4025 (N_4025,N_3575,N_3517);
nor U4026 (N_4026,N_3836,N_3607);
nand U4027 (N_4027,N_3896,N_3634);
and U4028 (N_4028,N_3648,N_3967);
nand U4029 (N_4029,N_3999,N_3809);
and U4030 (N_4030,N_3920,N_3858);
and U4031 (N_4031,N_3826,N_3599);
and U4032 (N_4032,N_3747,N_3531);
and U4033 (N_4033,N_3571,N_3755);
or U4034 (N_4034,N_3996,N_3509);
nand U4035 (N_4035,N_3881,N_3699);
nand U4036 (N_4036,N_3898,N_3816);
nand U4037 (N_4037,N_3925,N_3937);
nor U4038 (N_4038,N_3824,N_3662);
nand U4039 (N_4039,N_3726,N_3503);
and U4040 (N_4040,N_3702,N_3514);
nand U4041 (N_4041,N_3621,N_3593);
nand U4042 (N_4042,N_3504,N_3594);
nand U4043 (N_4043,N_3723,N_3819);
nand U4044 (N_4044,N_3668,N_3815);
nor U4045 (N_4045,N_3852,N_3939);
nor U4046 (N_4046,N_3617,N_3606);
nand U4047 (N_4047,N_3773,N_3560);
or U4048 (N_4048,N_3863,N_3591);
xor U4049 (N_4049,N_3846,N_3724);
nor U4050 (N_4050,N_3540,N_3832);
xnor U4051 (N_4051,N_3960,N_3865);
nor U4052 (N_4052,N_3838,N_3895);
and U4053 (N_4053,N_3508,N_3830);
and U4054 (N_4054,N_3953,N_3601);
or U4055 (N_4055,N_3859,N_3615);
or U4056 (N_4056,N_3586,N_3988);
nor U4057 (N_4057,N_3567,N_3872);
or U4058 (N_4058,N_3913,N_3978);
or U4059 (N_4059,N_3882,N_3520);
nor U4060 (N_4060,N_3875,N_3611);
nor U4061 (N_4061,N_3928,N_3907);
xor U4062 (N_4062,N_3700,N_3544);
and U4063 (N_4063,N_3831,N_3628);
and U4064 (N_4064,N_3760,N_3614);
nor U4065 (N_4065,N_3966,N_3742);
nor U4066 (N_4066,N_3718,N_3526);
and U4067 (N_4067,N_3515,N_3532);
and U4068 (N_4068,N_3679,N_3703);
nor U4069 (N_4069,N_3769,N_3713);
nand U4070 (N_4070,N_3541,N_3968);
nand U4071 (N_4071,N_3549,N_3786);
and U4072 (N_4072,N_3918,N_3944);
nor U4073 (N_4073,N_3949,N_3589);
nand U4074 (N_4074,N_3891,N_3657);
xor U4075 (N_4075,N_3897,N_3754);
or U4076 (N_4076,N_3758,N_3731);
nand U4077 (N_4077,N_3947,N_3934);
or U4078 (N_4078,N_3991,N_3958);
or U4079 (N_4079,N_3692,N_3719);
and U4080 (N_4080,N_3709,N_3546);
xor U4081 (N_4081,N_3665,N_3554);
or U4082 (N_4082,N_3977,N_3516);
or U4083 (N_4083,N_3711,N_3817);
nor U4084 (N_4084,N_3551,N_3808);
and U4085 (N_4085,N_3630,N_3869);
and U4086 (N_4086,N_3562,N_3559);
nor U4087 (N_4087,N_3994,N_3855);
or U4088 (N_4088,N_3890,N_3833);
or U4089 (N_4089,N_3558,N_3697);
nand U4090 (N_4090,N_3510,N_3548);
and U4091 (N_4091,N_3998,N_3624);
xnor U4092 (N_4092,N_3847,N_3677);
and U4093 (N_4093,N_3670,N_3524);
and U4094 (N_4094,N_3535,N_3583);
and U4095 (N_4095,N_3579,N_3637);
and U4096 (N_4096,N_3587,N_3659);
or U4097 (N_4097,N_3904,N_3582);
and U4098 (N_4098,N_3935,N_3739);
xnor U4099 (N_4099,N_3885,N_3941);
nand U4100 (N_4100,N_3845,N_3955);
nand U4101 (N_4101,N_3625,N_3737);
nand U4102 (N_4102,N_3736,N_3705);
or U4103 (N_4103,N_3658,N_3919);
nor U4104 (N_4104,N_3656,N_3777);
and U4105 (N_4105,N_3704,N_3997);
and U4106 (N_4106,N_3686,N_3902);
nand U4107 (N_4107,N_3794,N_3647);
or U4108 (N_4108,N_3797,N_3735);
nor U4109 (N_4109,N_3782,N_3979);
nand U4110 (N_4110,N_3671,N_3609);
nor U4111 (N_4111,N_3730,N_3800);
or U4112 (N_4112,N_3954,N_3619);
or U4113 (N_4113,N_3814,N_3633);
nand U4114 (N_4114,N_3570,N_3751);
or U4115 (N_4115,N_3795,N_3871);
nor U4116 (N_4116,N_3672,N_3568);
nor U4117 (N_4117,N_3722,N_3712);
and U4118 (N_4118,N_3912,N_3687);
and U4119 (N_4119,N_3774,N_3884);
nand U4120 (N_4120,N_3923,N_3632);
nor U4121 (N_4121,N_3915,N_3693);
nand U4122 (N_4122,N_3602,N_3580);
xnor U4123 (N_4123,N_3856,N_3596);
xor U4124 (N_4124,N_3903,N_3645);
and U4125 (N_4125,N_3789,N_3876);
and U4126 (N_4126,N_3985,N_3973);
or U4127 (N_4127,N_3622,N_3661);
and U4128 (N_4128,N_3879,N_3542);
and U4129 (N_4129,N_3725,N_3528);
nor U4130 (N_4130,N_3706,N_3506);
xnor U4131 (N_4131,N_3710,N_3880);
or U4132 (N_4132,N_3837,N_3536);
nor U4133 (N_4133,N_3801,N_3849);
nor U4134 (N_4134,N_3783,N_3756);
and U4135 (N_4135,N_3539,N_3980);
nor U4136 (N_4136,N_3813,N_3969);
nand U4137 (N_4137,N_3715,N_3660);
or U4138 (N_4138,N_3975,N_3577);
and U4139 (N_4139,N_3956,N_3653);
nor U4140 (N_4140,N_3543,N_3500);
nand U4141 (N_4141,N_3851,N_3810);
nor U4142 (N_4142,N_3803,N_3917);
nor U4143 (N_4143,N_3748,N_3533);
and U4144 (N_4144,N_3853,N_3638);
nor U4145 (N_4145,N_3986,N_3750);
nor U4146 (N_4146,N_3924,N_3708);
nand U4147 (N_4147,N_3561,N_3820);
xor U4148 (N_4148,N_3821,N_3942);
or U4149 (N_4149,N_3696,N_3983);
xnor U4150 (N_4150,N_3825,N_3906);
and U4151 (N_4151,N_3770,N_3584);
nor U4152 (N_4152,N_3519,N_3936);
nor U4153 (N_4153,N_3525,N_3938);
nand U4154 (N_4154,N_3970,N_3512);
or U4155 (N_4155,N_3695,N_3557);
or U4156 (N_4156,N_3604,N_3595);
or U4157 (N_4157,N_3733,N_3778);
nor U4158 (N_4158,N_3578,N_3894);
nand U4159 (N_4159,N_3762,N_3620);
xor U4160 (N_4160,N_3707,N_3623);
xnor U4161 (N_4161,N_3959,N_3732);
nand U4162 (N_4162,N_3974,N_3804);
nand U4163 (N_4163,N_3775,N_3688);
nor U4164 (N_4164,N_3501,N_3600);
and U4165 (N_4165,N_3690,N_3745);
or U4166 (N_4166,N_3574,N_3921);
xor U4167 (N_4167,N_3654,N_3893);
xnor U4168 (N_4168,N_3530,N_3753);
or U4169 (N_4169,N_3943,N_3835);
nand U4170 (N_4170,N_3933,N_3910);
or U4171 (N_4171,N_3812,N_3744);
and U4172 (N_4172,N_3768,N_3868);
nand U4173 (N_4173,N_3929,N_3771);
and U4174 (N_4174,N_3909,N_3563);
nor U4175 (N_4175,N_3681,N_3537);
nor U4176 (N_4176,N_3684,N_3666);
nor U4177 (N_4177,N_3764,N_3721);
or U4178 (N_4178,N_3664,N_3674);
or U4179 (N_4179,N_3828,N_3781);
nor U4180 (N_4180,N_3635,N_3613);
and U4181 (N_4181,N_3521,N_3874);
nand U4182 (N_4182,N_3522,N_3870);
and U4183 (N_4183,N_3743,N_3610);
or U4184 (N_4184,N_3566,N_3716);
nand U4185 (N_4185,N_3673,N_3676);
nor U4186 (N_4186,N_3553,N_3839);
nor U4187 (N_4187,N_3678,N_3534);
and U4188 (N_4188,N_3757,N_3888);
nand U4189 (N_4189,N_3564,N_3848);
nor U4190 (N_4190,N_3972,N_3799);
or U4191 (N_4191,N_3842,N_3626);
xor U4192 (N_4192,N_3886,N_3698);
nand U4193 (N_4193,N_3765,N_3667);
and U4194 (N_4194,N_3779,N_3585);
xor U4195 (N_4195,N_3592,N_3729);
and U4196 (N_4196,N_3552,N_3952);
and U4197 (N_4197,N_3513,N_3900);
nor U4198 (N_4198,N_3734,N_3796);
nor U4199 (N_4199,N_3766,N_3598);
nand U4200 (N_4200,N_3685,N_3857);
nand U4201 (N_4201,N_3840,N_3627);
nor U4202 (N_4202,N_3538,N_3507);
nor U4203 (N_4203,N_3827,N_3850);
nand U4204 (N_4204,N_3818,N_3806);
nor U4205 (N_4205,N_3590,N_3761);
nor U4206 (N_4206,N_3752,N_3505);
and U4207 (N_4207,N_3502,N_3931);
nand U4208 (N_4208,N_3866,N_3663);
nand U4209 (N_4209,N_3989,N_3993);
xnor U4210 (N_4210,N_3926,N_3948);
and U4211 (N_4211,N_3694,N_3862);
nor U4212 (N_4212,N_3717,N_3914);
and U4213 (N_4213,N_3572,N_3901);
xor U4214 (N_4214,N_3649,N_3603);
or U4215 (N_4215,N_3689,N_3788);
and U4216 (N_4216,N_3981,N_3728);
nand U4217 (N_4217,N_3720,N_3877);
nand U4218 (N_4218,N_3691,N_3784);
nor U4219 (N_4219,N_3961,N_3652);
xnor U4220 (N_4220,N_3905,N_3965);
and U4221 (N_4221,N_3995,N_3829);
or U4222 (N_4222,N_3787,N_3608);
nand U4223 (N_4223,N_3957,N_3529);
or U4224 (N_4224,N_3643,N_3927);
nor U4225 (N_4225,N_3987,N_3597);
nand U4226 (N_4226,N_3746,N_3976);
or U4227 (N_4227,N_3727,N_3930);
nor U4228 (N_4228,N_3802,N_3932);
nand U4229 (N_4229,N_3776,N_3767);
or U4230 (N_4230,N_3523,N_3612);
nor U4231 (N_4231,N_3740,N_3873);
nor U4232 (N_4232,N_3636,N_3963);
nor U4233 (N_4233,N_3556,N_3807);
nor U4234 (N_4234,N_3581,N_3867);
xnor U4235 (N_4235,N_3680,N_3749);
nand U4236 (N_4236,N_3569,N_3982);
and U4237 (N_4237,N_3990,N_3547);
and U4238 (N_4238,N_3946,N_3780);
xnor U4239 (N_4239,N_3792,N_3843);
and U4240 (N_4240,N_3844,N_3823);
or U4241 (N_4241,N_3861,N_3964);
or U4242 (N_4242,N_3984,N_3864);
nor U4243 (N_4243,N_3644,N_3518);
nand U4244 (N_4244,N_3790,N_3714);
and U4245 (N_4245,N_3887,N_3655);
nand U4246 (N_4246,N_3618,N_3922);
nor U4247 (N_4247,N_3889,N_3651);
nand U4248 (N_4248,N_3805,N_3545);
and U4249 (N_4249,N_3642,N_3701);
and U4250 (N_4250,N_3695,N_3639);
nor U4251 (N_4251,N_3949,N_3957);
or U4252 (N_4252,N_3804,N_3696);
nor U4253 (N_4253,N_3929,N_3770);
and U4254 (N_4254,N_3667,N_3530);
and U4255 (N_4255,N_3896,N_3999);
xnor U4256 (N_4256,N_3723,N_3612);
nor U4257 (N_4257,N_3840,N_3509);
nor U4258 (N_4258,N_3538,N_3537);
nand U4259 (N_4259,N_3587,N_3503);
nand U4260 (N_4260,N_3698,N_3970);
xnor U4261 (N_4261,N_3698,N_3841);
nor U4262 (N_4262,N_3694,N_3907);
nor U4263 (N_4263,N_3720,N_3903);
or U4264 (N_4264,N_3959,N_3822);
nor U4265 (N_4265,N_3900,N_3727);
nand U4266 (N_4266,N_3939,N_3953);
xnor U4267 (N_4267,N_3584,N_3736);
or U4268 (N_4268,N_3695,N_3706);
or U4269 (N_4269,N_3561,N_3974);
and U4270 (N_4270,N_3974,N_3616);
nor U4271 (N_4271,N_3803,N_3935);
nand U4272 (N_4272,N_3954,N_3776);
xor U4273 (N_4273,N_3592,N_3565);
xor U4274 (N_4274,N_3654,N_3851);
nand U4275 (N_4275,N_3881,N_3869);
nor U4276 (N_4276,N_3748,N_3555);
or U4277 (N_4277,N_3865,N_3962);
and U4278 (N_4278,N_3848,N_3521);
xnor U4279 (N_4279,N_3721,N_3980);
nand U4280 (N_4280,N_3521,N_3881);
nor U4281 (N_4281,N_3997,N_3544);
and U4282 (N_4282,N_3862,N_3991);
or U4283 (N_4283,N_3548,N_3592);
and U4284 (N_4284,N_3728,N_3840);
nor U4285 (N_4285,N_3517,N_3885);
or U4286 (N_4286,N_3789,N_3532);
nand U4287 (N_4287,N_3550,N_3789);
nand U4288 (N_4288,N_3616,N_3848);
and U4289 (N_4289,N_3608,N_3507);
and U4290 (N_4290,N_3776,N_3615);
or U4291 (N_4291,N_3877,N_3876);
nor U4292 (N_4292,N_3882,N_3653);
and U4293 (N_4293,N_3589,N_3880);
nor U4294 (N_4294,N_3605,N_3775);
or U4295 (N_4295,N_3771,N_3796);
xor U4296 (N_4296,N_3679,N_3781);
xor U4297 (N_4297,N_3847,N_3919);
or U4298 (N_4298,N_3523,N_3828);
xnor U4299 (N_4299,N_3511,N_3564);
nor U4300 (N_4300,N_3667,N_3908);
nand U4301 (N_4301,N_3708,N_3981);
nor U4302 (N_4302,N_3551,N_3774);
nor U4303 (N_4303,N_3617,N_3674);
or U4304 (N_4304,N_3901,N_3696);
nand U4305 (N_4305,N_3716,N_3980);
and U4306 (N_4306,N_3552,N_3537);
nor U4307 (N_4307,N_3790,N_3862);
and U4308 (N_4308,N_3848,N_3986);
nor U4309 (N_4309,N_3736,N_3827);
and U4310 (N_4310,N_3805,N_3686);
and U4311 (N_4311,N_3816,N_3836);
nor U4312 (N_4312,N_3678,N_3689);
nor U4313 (N_4313,N_3789,N_3745);
or U4314 (N_4314,N_3946,N_3732);
xor U4315 (N_4315,N_3568,N_3819);
nand U4316 (N_4316,N_3799,N_3666);
and U4317 (N_4317,N_3705,N_3534);
nand U4318 (N_4318,N_3575,N_3638);
xor U4319 (N_4319,N_3689,N_3877);
nor U4320 (N_4320,N_3753,N_3689);
or U4321 (N_4321,N_3879,N_3871);
or U4322 (N_4322,N_3902,N_3694);
or U4323 (N_4323,N_3732,N_3870);
or U4324 (N_4324,N_3644,N_3735);
xnor U4325 (N_4325,N_3526,N_3701);
nand U4326 (N_4326,N_3528,N_3690);
and U4327 (N_4327,N_3790,N_3726);
and U4328 (N_4328,N_3904,N_3689);
nand U4329 (N_4329,N_3845,N_3806);
nor U4330 (N_4330,N_3767,N_3948);
nand U4331 (N_4331,N_3912,N_3749);
nand U4332 (N_4332,N_3949,N_3724);
xor U4333 (N_4333,N_3996,N_3745);
nor U4334 (N_4334,N_3912,N_3936);
and U4335 (N_4335,N_3638,N_3907);
nor U4336 (N_4336,N_3660,N_3808);
and U4337 (N_4337,N_3508,N_3921);
and U4338 (N_4338,N_3897,N_3981);
or U4339 (N_4339,N_3822,N_3630);
nand U4340 (N_4340,N_3650,N_3747);
or U4341 (N_4341,N_3863,N_3504);
nand U4342 (N_4342,N_3677,N_3573);
and U4343 (N_4343,N_3722,N_3776);
and U4344 (N_4344,N_3820,N_3537);
nand U4345 (N_4345,N_3515,N_3838);
xor U4346 (N_4346,N_3665,N_3827);
nand U4347 (N_4347,N_3856,N_3662);
xnor U4348 (N_4348,N_3832,N_3720);
nor U4349 (N_4349,N_3665,N_3766);
and U4350 (N_4350,N_3632,N_3711);
nor U4351 (N_4351,N_3533,N_3839);
or U4352 (N_4352,N_3685,N_3537);
and U4353 (N_4353,N_3739,N_3555);
xor U4354 (N_4354,N_3845,N_3956);
and U4355 (N_4355,N_3682,N_3584);
nand U4356 (N_4356,N_3804,N_3813);
and U4357 (N_4357,N_3703,N_3779);
or U4358 (N_4358,N_3570,N_3953);
and U4359 (N_4359,N_3540,N_3509);
xnor U4360 (N_4360,N_3607,N_3941);
or U4361 (N_4361,N_3590,N_3944);
nand U4362 (N_4362,N_3737,N_3789);
or U4363 (N_4363,N_3547,N_3940);
nor U4364 (N_4364,N_3974,N_3696);
or U4365 (N_4365,N_3592,N_3543);
or U4366 (N_4366,N_3801,N_3515);
nor U4367 (N_4367,N_3671,N_3891);
xnor U4368 (N_4368,N_3708,N_3626);
nand U4369 (N_4369,N_3694,N_3831);
and U4370 (N_4370,N_3855,N_3965);
and U4371 (N_4371,N_3641,N_3654);
nor U4372 (N_4372,N_3994,N_3552);
nand U4373 (N_4373,N_3666,N_3567);
or U4374 (N_4374,N_3959,N_3664);
or U4375 (N_4375,N_3670,N_3662);
nand U4376 (N_4376,N_3525,N_3701);
nand U4377 (N_4377,N_3998,N_3772);
nor U4378 (N_4378,N_3503,N_3591);
nor U4379 (N_4379,N_3616,N_3710);
xnor U4380 (N_4380,N_3647,N_3631);
xor U4381 (N_4381,N_3572,N_3567);
xor U4382 (N_4382,N_3850,N_3994);
nor U4383 (N_4383,N_3611,N_3526);
nand U4384 (N_4384,N_3660,N_3671);
nor U4385 (N_4385,N_3631,N_3895);
xnor U4386 (N_4386,N_3557,N_3884);
and U4387 (N_4387,N_3881,N_3612);
and U4388 (N_4388,N_3703,N_3715);
nor U4389 (N_4389,N_3832,N_3967);
xnor U4390 (N_4390,N_3637,N_3588);
nor U4391 (N_4391,N_3685,N_3588);
nor U4392 (N_4392,N_3924,N_3884);
or U4393 (N_4393,N_3579,N_3818);
nor U4394 (N_4394,N_3717,N_3882);
and U4395 (N_4395,N_3505,N_3942);
or U4396 (N_4396,N_3753,N_3938);
nand U4397 (N_4397,N_3624,N_3594);
xor U4398 (N_4398,N_3925,N_3977);
xor U4399 (N_4399,N_3793,N_3703);
and U4400 (N_4400,N_3719,N_3550);
nor U4401 (N_4401,N_3947,N_3535);
nand U4402 (N_4402,N_3835,N_3830);
nand U4403 (N_4403,N_3762,N_3701);
xor U4404 (N_4404,N_3949,N_3881);
or U4405 (N_4405,N_3861,N_3523);
nand U4406 (N_4406,N_3530,N_3881);
or U4407 (N_4407,N_3890,N_3651);
xor U4408 (N_4408,N_3626,N_3793);
nand U4409 (N_4409,N_3898,N_3868);
and U4410 (N_4410,N_3948,N_3582);
and U4411 (N_4411,N_3851,N_3637);
and U4412 (N_4412,N_3645,N_3977);
nor U4413 (N_4413,N_3688,N_3648);
nand U4414 (N_4414,N_3604,N_3511);
nand U4415 (N_4415,N_3566,N_3699);
nand U4416 (N_4416,N_3951,N_3637);
and U4417 (N_4417,N_3940,N_3647);
or U4418 (N_4418,N_3858,N_3946);
or U4419 (N_4419,N_3907,N_3724);
and U4420 (N_4420,N_3641,N_3727);
nor U4421 (N_4421,N_3907,N_3652);
and U4422 (N_4422,N_3516,N_3600);
or U4423 (N_4423,N_3891,N_3737);
nor U4424 (N_4424,N_3580,N_3906);
nand U4425 (N_4425,N_3753,N_3802);
xnor U4426 (N_4426,N_3837,N_3526);
nand U4427 (N_4427,N_3820,N_3925);
or U4428 (N_4428,N_3747,N_3603);
nand U4429 (N_4429,N_3692,N_3745);
nor U4430 (N_4430,N_3742,N_3802);
xor U4431 (N_4431,N_3512,N_3633);
nand U4432 (N_4432,N_3895,N_3636);
nor U4433 (N_4433,N_3974,N_3718);
nor U4434 (N_4434,N_3705,N_3750);
nand U4435 (N_4435,N_3943,N_3962);
and U4436 (N_4436,N_3750,N_3742);
and U4437 (N_4437,N_3599,N_3563);
or U4438 (N_4438,N_3892,N_3559);
or U4439 (N_4439,N_3503,N_3990);
nor U4440 (N_4440,N_3738,N_3838);
xnor U4441 (N_4441,N_3915,N_3701);
or U4442 (N_4442,N_3621,N_3511);
nand U4443 (N_4443,N_3945,N_3608);
nor U4444 (N_4444,N_3723,N_3652);
or U4445 (N_4445,N_3879,N_3723);
nand U4446 (N_4446,N_3736,N_3777);
or U4447 (N_4447,N_3815,N_3584);
nor U4448 (N_4448,N_3770,N_3850);
nand U4449 (N_4449,N_3753,N_3603);
nor U4450 (N_4450,N_3891,N_3896);
nand U4451 (N_4451,N_3798,N_3709);
xnor U4452 (N_4452,N_3612,N_3511);
and U4453 (N_4453,N_3579,N_3586);
nand U4454 (N_4454,N_3777,N_3578);
nor U4455 (N_4455,N_3823,N_3590);
or U4456 (N_4456,N_3685,N_3774);
nor U4457 (N_4457,N_3806,N_3990);
or U4458 (N_4458,N_3703,N_3664);
and U4459 (N_4459,N_3576,N_3936);
and U4460 (N_4460,N_3816,N_3644);
xnor U4461 (N_4461,N_3810,N_3698);
nor U4462 (N_4462,N_3508,N_3703);
xor U4463 (N_4463,N_3770,N_3604);
nand U4464 (N_4464,N_3512,N_3815);
or U4465 (N_4465,N_3604,N_3546);
nand U4466 (N_4466,N_3501,N_3537);
or U4467 (N_4467,N_3950,N_3767);
nor U4468 (N_4468,N_3549,N_3595);
and U4469 (N_4469,N_3676,N_3932);
and U4470 (N_4470,N_3711,N_3719);
or U4471 (N_4471,N_3914,N_3913);
and U4472 (N_4472,N_3705,N_3527);
nor U4473 (N_4473,N_3736,N_3587);
and U4474 (N_4474,N_3998,N_3629);
xor U4475 (N_4475,N_3652,N_3539);
or U4476 (N_4476,N_3973,N_3599);
nor U4477 (N_4477,N_3825,N_3750);
xor U4478 (N_4478,N_3894,N_3598);
nand U4479 (N_4479,N_3606,N_3510);
nor U4480 (N_4480,N_3910,N_3814);
nand U4481 (N_4481,N_3549,N_3558);
nand U4482 (N_4482,N_3843,N_3842);
or U4483 (N_4483,N_3669,N_3897);
or U4484 (N_4484,N_3586,N_3698);
xor U4485 (N_4485,N_3676,N_3808);
or U4486 (N_4486,N_3630,N_3852);
nor U4487 (N_4487,N_3916,N_3732);
nand U4488 (N_4488,N_3984,N_3680);
or U4489 (N_4489,N_3956,N_3957);
or U4490 (N_4490,N_3725,N_3848);
nand U4491 (N_4491,N_3621,N_3530);
and U4492 (N_4492,N_3991,N_3521);
or U4493 (N_4493,N_3640,N_3832);
nor U4494 (N_4494,N_3505,N_3880);
nand U4495 (N_4495,N_3743,N_3680);
and U4496 (N_4496,N_3975,N_3702);
nor U4497 (N_4497,N_3608,N_3744);
and U4498 (N_4498,N_3661,N_3541);
or U4499 (N_4499,N_3810,N_3648);
and U4500 (N_4500,N_4342,N_4149);
or U4501 (N_4501,N_4254,N_4016);
and U4502 (N_4502,N_4322,N_4439);
or U4503 (N_4503,N_4275,N_4328);
or U4504 (N_4504,N_4435,N_4233);
nand U4505 (N_4505,N_4413,N_4122);
or U4506 (N_4506,N_4491,N_4399);
nor U4507 (N_4507,N_4277,N_4177);
nand U4508 (N_4508,N_4118,N_4403);
nand U4509 (N_4509,N_4438,N_4467);
xnor U4510 (N_4510,N_4139,N_4428);
nor U4511 (N_4511,N_4338,N_4079);
and U4512 (N_4512,N_4488,N_4127);
and U4513 (N_4513,N_4462,N_4216);
nand U4514 (N_4514,N_4228,N_4286);
and U4515 (N_4515,N_4256,N_4384);
and U4516 (N_4516,N_4148,N_4451);
nor U4517 (N_4517,N_4238,N_4006);
and U4518 (N_4518,N_4013,N_4001);
or U4519 (N_4519,N_4408,N_4101);
nor U4520 (N_4520,N_4397,N_4489);
and U4521 (N_4521,N_4310,N_4221);
or U4522 (N_4522,N_4178,N_4250);
or U4523 (N_4523,N_4372,N_4436);
xnor U4524 (N_4524,N_4396,N_4158);
nand U4525 (N_4525,N_4093,N_4151);
xor U4526 (N_4526,N_4456,N_4214);
nor U4527 (N_4527,N_4077,N_4219);
nand U4528 (N_4528,N_4134,N_4272);
and U4529 (N_4529,N_4213,N_4369);
nand U4530 (N_4530,N_4363,N_4318);
nand U4531 (N_4531,N_4119,N_4291);
nand U4532 (N_4532,N_4131,N_4416);
and U4533 (N_4533,N_4374,N_4426);
nor U4534 (N_4534,N_4305,N_4126);
or U4535 (N_4535,N_4442,N_4311);
or U4536 (N_4536,N_4097,N_4031);
xnor U4537 (N_4537,N_4029,N_4080);
nand U4538 (N_4538,N_4303,N_4184);
or U4539 (N_4539,N_4162,N_4064);
nand U4540 (N_4540,N_4248,N_4479);
nand U4541 (N_4541,N_4030,N_4495);
and U4542 (N_4542,N_4483,N_4215);
nand U4543 (N_4543,N_4249,N_4446);
and U4544 (N_4544,N_4071,N_4498);
nand U4545 (N_4545,N_4344,N_4383);
and U4546 (N_4546,N_4279,N_4022);
and U4547 (N_4547,N_4458,N_4157);
nand U4548 (N_4548,N_4472,N_4058);
and U4549 (N_4549,N_4315,N_4251);
nor U4550 (N_4550,N_4468,N_4239);
nand U4551 (N_4551,N_4052,N_4260);
or U4552 (N_4552,N_4323,N_4181);
or U4553 (N_4553,N_4390,N_4459);
nor U4554 (N_4554,N_4194,N_4335);
and U4555 (N_4555,N_4032,N_4175);
nand U4556 (N_4556,N_4429,N_4469);
nor U4557 (N_4557,N_4120,N_4263);
and U4558 (N_4558,N_4350,N_4043);
nand U4559 (N_4559,N_4081,N_4227);
and U4560 (N_4560,N_4265,N_4018);
and U4561 (N_4561,N_4021,N_4146);
or U4562 (N_4562,N_4153,N_4395);
or U4563 (N_4563,N_4094,N_4267);
or U4564 (N_4564,N_4110,N_4357);
or U4565 (N_4565,N_4485,N_4351);
nor U4566 (N_4566,N_4476,N_4074);
nand U4567 (N_4567,N_4075,N_4063);
and U4568 (N_4568,N_4222,N_4261);
and U4569 (N_4569,N_4257,N_4060);
and U4570 (N_4570,N_4061,N_4172);
xnor U4571 (N_4571,N_4282,N_4044);
nand U4572 (N_4572,N_4378,N_4176);
or U4573 (N_4573,N_4220,N_4298);
and U4574 (N_4574,N_4053,N_4306);
nand U4575 (N_4575,N_4117,N_4202);
and U4576 (N_4576,N_4293,N_4288);
nand U4577 (N_4577,N_4147,N_4180);
or U4578 (N_4578,N_4155,N_4355);
nand U4579 (N_4579,N_4336,N_4089);
nor U4580 (N_4580,N_4103,N_4314);
and U4581 (N_4581,N_4448,N_4102);
xnor U4582 (N_4582,N_4169,N_4166);
and U4583 (N_4583,N_4112,N_4065);
xor U4584 (N_4584,N_4301,N_4240);
nand U4585 (N_4585,N_4133,N_4038);
nor U4586 (N_4586,N_4206,N_4212);
or U4587 (N_4587,N_4128,N_4003);
xor U4588 (N_4588,N_4391,N_4283);
or U4589 (N_4589,N_4193,N_4475);
and U4590 (N_4590,N_4247,N_4207);
nor U4591 (N_4591,N_4385,N_4224);
or U4592 (N_4592,N_4300,N_4269);
or U4593 (N_4593,N_4307,N_4072);
and U4594 (N_4594,N_4054,N_4360);
nor U4595 (N_4595,N_4009,N_4440);
nor U4596 (N_4596,N_4364,N_4258);
nor U4597 (N_4597,N_4441,N_4237);
nor U4598 (N_4598,N_4161,N_4020);
nand U4599 (N_4599,N_4368,N_4358);
nor U4600 (N_4600,N_4226,N_4411);
nor U4601 (N_4601,N_4142,N_4455);
xor U4602 (N_4602,N_4454,N_4199);
and U4603 (N_4603,N_4059,N_4168);
nor U4604 (N_4604,N_4015,N_4370);
or U4605 (N_4605,N_4473,N_4345);
and U4606 (N_4606,N_4235,N_4095);
or U4607 (N_4607,N_4167,N_4423);
or U4608 (N_4608,N_4105,N_4039);
nor U4609 (N_4609,N_4379,N_4409);
and U4610 (N_4610,N_4312,N_4460);
nand U4611 (N_4611,N_4490,N_4337);
and U4612 (N_4612,N_4088,N_4412);
and U4613 (N_4613,N_4244,N_4241);
or U4614 (N_4614,N_4218,N_4457);
and U4615 (N_4615,N_4253,N_4343);
nand U4616 (N_4616,N_4208,N_4185);
and U4617 (N_4617,N_4474,N_4203);
nand U4618 (N_4618,N_4477,N_4163);
nand U4619 (N_4619,N_4171,N_4047);
and U4620 (N_4620,N_4327,N_4091);
xnor U4621 (N_4621,N_4045,N_4245);
xor U4622 (N_4622,N_4443,N_4041);
nand U4623 (N_4623,N_4450,N_4452);
nor U4624 (N_4624,N_4154,N_4046);
or U4625 (N_4625,N_4414,N_4373);
nand U4626 (N_4626,N_4144,N_4198);
or U4627 (N_4627,N_4138,N_4406);
nand U4628 (N_4628,N_4324,N_4349);
and U4629 (N_4629,N_4422,N_4100);
or U4630 (N_4630,N_4129,N_4010);
or U4631 (N_4631,N_4280,N_4297);
nor U4632 (N_4632,N_4086,N_4421);
or U4633 (N_4633,N_4444,N_4090);
nand U4634 (N_4634,N_4493,N_4007);
or U4635 (N_4635,N_4114,N_4137);
xor U4636 (N_4636,N_4078,N_4353);
nand U4637 (N_4637,N_4434,N_4389);
and U4638 (N_4638,N_4376,N_4035);
and U4639 (N_4639,N_4432,N_4316);
xnor U4640 (N_4640,N_4197,N_4209);
and U4641 (N_4641,N_4140,N_4069);
nand U4642 (N_4642,N_4425,N_4024);
and U4643 (N_4643,N_4076,N_4321);
xor U4644 (N_4644,N_4330,N_4268);
and U4645 (N_4645,N_4229,N_4361);
and U4646 (N_4646,N_4381,N_4051);
and U4647 (N_4647,N_4463,N_4400);
nor U4648 (N_4648,N_4289,N_4070);
nor U4649 (N_4649,N_4281,N_4271);
nand U4650 (N_4650,N_4084,N_4073);
nand U4651 (N_4651,N_4099,N_4331);
nand U4652 (N_4652,N_4042,N_4002);
nor U4653 (N_4653,N_4200,N_4481);
nor U4654 (N_4654,N_4367,N_4023);
nand U4655 (N_4655,N_4453,N_4471);
and U4656 (N_4656,N_4055,N_4309);
nor U4657 (N_4657,N_4121,N_4132);
and U4658 (N_4658,N_4274,N_4496);
nand U4659 (N_4659,N_4332,N_4123);
or U4660 (N_4660,N_4417,N_4494);
nor U4661 (N_4661,N_4499,N_4296);
nor U4662 (N_4662,N_4401,N_4359);
xor U4663 (N_4663,N_4027,N_4050);
nor U4664 (N_4664,N_4375,N_4225);
xnor U4665 (N_4665,N_4415,N_4317);
or U4666 (N_4666,N_4246,N_4348);
xor U4667 (N_4667,N_4231,N_4266);
and U4668 (N_4668,N_4008,N_4033);
nor U4669 (N_4669,N_4326,N_4083);
and U4670 (N_4670,N_4124,N_4285);
or U4671 (N_4671,N_4325,N_4377);
nor U4672 (N_4672,N_4234,N_4273);
and U4673 (N_4673,N_4056,N_4341);
nand U4674 (N_4674,N_4201,N_4340);
nand U4675 (N_4675,N_4135,N_4160);
nor U4676 (N_4676,N_4111,N_4407);
nor U4677 (N_4677,N_4107,N_4017);
and U4678 (N_4678,N_4365,N_4294);
and U4679 (N_4679,N_4392,N_4427);
and U4680 (N_4680,N_4243,N_4262);
or U4681 (N_4681,N_4362,N_4026);
nor U4682 (N_4682,N_4182,N_4109);
nor U4683 (N_4683,N_4304,N_4388);
or U4684 (N_4684,N_4486,N_4048);
nor U4685 (N_4685,N_4386,N_4191);
nor U4686 (N_4686,N_4449,N_4085);
or U4687 (N_4687,N_4346,N_4196);
xor U4688 (N_4688,N_4040,N_4308);
or U4689 (N_4689,N_4366,N_4179);
and U4690 (N_4690,N_4082,N_4036);
nor U4691 (N_4691,N_4482,N_4394);
nand U4692 (N_4692,N_4313,N_4125);
nand U4693 (N_4693,N_4170,N_4431);
and U4694 (N_4694,N_4145,N_4393);
nand U4695 (N_4695,N_4329,N_4270);
or U4696 (N_4696,N_4188,N_4255);
xor U4697 (N_4697,N_4049,N_4419);
nand U4698 (N_4698,N_4264,N_4287);
nand U4699 (N_4699,N_4062,N_4497);
xor U4700 (N_4700,N_4424,N_4211);
nor U4701 (N_4701,N_4116,N_4217);
nand U4702 (N_4702,N_4130,N_4098);
nand U4703 (N_4703,N_4433,N_4339);
and U4704 (N_4704,N_4205,N_4164);
and U4705 (N_4705,N_4104,N_4096);
xnor U4706 (N_4706,N_4445,N_4106);
or U4707 (N_4707,N_4034,N_4405);
nor U4708 (N_4708,N_4470,N_4012);
and U4709 (N_4709,N_4011,N_4352);
and U4710 (N_4710,N_4210,N_4252);
nor U4711 (N_4711,N_4136,N_4320);
or U4712 (N_4712,N_4334,N_4156);
nand U4713 (N_4713,N_4230,N_4066);
or U4714 (N_4714,N_4382,N_4019);
nor U4715 (N_4715,N_4292,N_4420);
or U4716 (N_4716,N_4115,N_4430);
xnor U4717 (N_4717,N_4284,N_4152);
nor U4718 (N_4718,N_4478,N_4380);
or U4719 (N_4719,N_4242,N_4165);
xor U4720 (N_4720,N_4005,N_4067);
nor U4721 (N_4721,N_4025,N_4437);
nand U4722 (N_4722,N_4465,N_4186);
or U4723 (N_4723,N_4410,N_4387);
nor U4724 (N_4724,N_4232,N_4183);
nor U4725 (N_4725,N_4356,N_4190);
and U4726 (N_4726,N_4492,N_4299);
and U4727 (N_4727,N_4108,N_4159);
or U4728 (N_4728,N_4004,N_4347);
or U4729 (N_4729,N_4236,N_4173);
or U4730 (N_4730,N_4398,N_4259);
and U4731 (N_4731,N_4028,N_4087);
or U4732 (N_4732,N_4333,N_4014);
and U4733 (N_4733,N_4354,N_4402);
xor U4734 (N_4734,N_4278,N_4195);
and U4735 (N_4735,N_4487,N_4464);
or U4736 (N_4736,N_4404,N_4466);
or U4737 (N_4737,N_4092,N_4113);
or U4738 (N_4738,N_4057,N_4371);
nand U4739 (N_4739,N_4484,N_4000);
and U4740 (N_4740,N_4037,N_4174);
nand U4741 (N_4741,N_4480,N_4319);
and U4742 (N_4742,N_4143,N_4447);
nor U4743 (N_4743,N_4068,N_4461);
or U4744 (N_4744,N_4204,N_4295);
nand U4745 (N_4745,N_4187,N_4290);
or U4746 (N_4746,N_4276,N_4189);
nand U4747 (N_4747,N_4192,N_4302);
nor U4748 (N_4748,N_4141,N_4223);
and U4749 (N_4749,N_4418,N_4150);
nand U4750 (N_4750,N_4333,N_4097);
and U4751 (N_4751,N_4245,N_4326);
nand U4752 (N_4752,N_4366,N_4353);
xnor U4753 (N_4753,N_4385,N_4048);
nor U4754 (N_4754,N_4190,N_4475);
or U4755 (N_4755,N_4257,N_4258);
nand U4756 (N_4756,N_4057,N_4197);
nor U4757 (N_4757,N_4335,N_4221);
xnor U4758 (N_4758,N_4053,N_4201);
and U4759 (N_4759,N_4060,N_4227);
nor U4760 (N_4760,N_4105,N_4140);
or U4761 (N_4761,N_4479,N_4092);
nand U4762 (N_4762,N_4341,N_4496);
nor U4763 (N_4763,N_4259,N_4344);
nand U4764 (N_4764,N_4098,N_4485);
nand U4765 (N_4765,N_4252,N_4474);
nand U4766 (N_4766,N_4125,N_4016);
and U4767 (N_4767,N_4047,N_4149);
and U4768 (N_4768,N_4152,N_4389);
or U4769 (N_4769,N_4214,N_4015);
nand U4770 (N_4770,N_4497,N_4398);
or U4771 (N_4771,N_4047,N_4267);
xor U4772 (N_4772,N_4328,N_4495);
nand U4773 (N_4773,N_4245,N_4192);
nand U4774 (N_4774,N_4425,N_4342);
nand U4775 (N_4775,N_4203,N_4259);
and U4776 (N_4776,N_4201,N_4029);
nand U4777 (N_4777,N_4398,N_4335);
xor U4778 (N_4778,N_4013,N_4297);
or U4779 (N_4779,N_4465,N_4234);
xor U4780 (N_4780,N_4019,N_4150);
and U4781 (N_4781,N_4161,N_4012);
and U4782 (N_4782,N_4165,N_4120);
nor U4783 (N_4783,N_4110,N_4230);
and U4784 (N_4784,N_4119,N_4065);
and U4785 (N_4785,N_4232,N_4348);
and U4786 (N_4786,N_4424,N_4382);
xor U4787 (N_4787,N_4392,N_4017);
or U4788 (N_4788,N_4333,N_4479);
nand U4789 (N_4789,N_4127,N_4470);
nor U4790 (N_4790,N_4409,N_4469);
nand U4791 (N_4791,N_4207,N_4252);
nor U4792 (N_4792,N_4068,N_4240);
nand U4793 (N_4793,N_4324,N_4145);
and U4794 (N_4794,N_4190,N_4004);
nor U4795 (N_4795,N_4484,N_4319);
xor U4796 (N_4796,N_4008,N_4488);
or U4797 (N_4797,N_4300,N_4188);
nand U4798 (N_4798,N_4138,N_4314);
nor U4799 (N_4799,N_4485,N_4228);
nand U4800 (N_4800,N_4313,N_4272);
nor U4801 (N_4801,N_4394,N_4212);
and U4802 (N_4802,N_4329,N_4385);
nor U4803 (N_4803,N_4408,N_4284);
nor U4804 (N_4804,N_4262,N_4455);
and U4805 (N_4805,N_4258,N_4373);
and U4806 (N_4806,N_4087,N_4478);
and U4807 (N_4807,N_4094,N_4358);
or U4808 (N_4808,N_4215,N_4149);
and U4809 (N_4809,N_4478,N_4146);
and U4810 (N_4810,N_4122,N_4411);
and U4811 (N_4811,N_4345,N_4296);
nand U4812 (N_4812,N_4374,N_4092);
or U4813 (N_4813,N_4133,N_4475);
xor U4814 (N_4814,N_4456,N_4440);
nor U4815 (N_4815,N_4230,N_4462);
and U4816 (N_4816,N_4341,N_4243);
nor U4817 (N_4817,N_4107,N_4442);
and U4818 (N_4818,N_4335,N_4274);
nor U4819 (N_4819,N_4065,N_4427);
and U4820 (N_4820,N_4429,N_4016);
or U4821 (N_4821,N_4425,N_4347);
nand U4822 (N_4822,N_4364,N_4170);
and U4823 (N_4823,N_4195,N_4458);
nand U4824 (N_4824,N_4253,N_4478);
nand U4825 (N_4825,N_4140,N_4319);
nand U4826 (N_4826,N_4484,N_4441);
or U4827 (N_4827,N_4282,N_4398);
nand U4828 (N_4828,N_4104,N_4272);
and U4829 (N_4829,N_4383,N_4092);
nand U4830 (N_4830,N_4228,N_4167);
nand U4831 (N_4831,N_4386,N_4417);
and U4832 (N_4832,N_4475,N_4458);
or U4833 (N_4833,N_4139,N_4075);
nor U4834 (N_4834,N_4331,N_4091);
and U4835 (N_4835,N_4325,N_4098);
and U4836 (N_4836,N_4055,N_4202);
or U4837 (N_4837,N_4316,N_4257);
xnor U4838 (N_4838,N_4384,N_4433);
nor U4839 (N_4839,N_4237,N_4397);
nand U4840 (N_4840,N_4427,N_4447);
xor U4841 (N_4841,N_4465,N_4166);
or U4842 (N_4842,N_4219,N_4337);
nor U4843 (N_4843,N_4402,N_4474);
nand U4844 (N_4844,N_4345,N_4157);
xnor U4845 (N_4845,N_4038,N_4406);
nor U4846 (N_4846,N_4338,N_4205);
or U4847 (N_4847,N_4262,N_4334);
xnor U4848 (N_4848,N_4434,N_4317);
or U4849 (N_4849,N_4001,N_4378);
or U4850 (N_4850,N_4354,N_4006);
xor U4851 (N_4851,N_4471,N_4061);
or U4852 (N_4852,N_4462,N_4215);
xnor U4853 (N_4853,N_4322,N_4035);
nand U4854 (N_4854,N_4408,N_4486);
and U4855 (N_4855,N_4288,N_4316);
or U4856 (N_4856,N_4433,N_4066);
xor U4857 (N_4857,N_4040,N_4187);
nand U4858 (N_4858,N_4071,N_4151);
nor U4859 (N_4859,N_4130,N_4245);
or U4860 (N_4860,N_4142,N_4227);
or U4861 (N_4861,N_4271,N_4303);
and U4862 (N_4862,N_4499,N_4498);
nand U4863 (N_4863,N_4432,N_4364);
nor U4864 (N_4864,N_4348,N_4021);
nand U4865 (N_4865,N_4409,N_4027);
nand U4866 (N_4866,N_4474,N_4026);
nor U4867 (N_4867,N_4477,N_4013);
nor U4868 (N_4868,N_4401,N_4424);
and U4869 (N_4869,N_4345,N_4462);
nand U4870 (N_4870,N_4210,N_4249);
and U4871 (N_4871,N_4386,N_4465);
nand U4872 (N_4872,N_4382,N_4388);
and U4873 (N_4873,N_4242,N_4262);
nor U4874 (N_4874,N_4399,N_4306);
or U4875 (N_4875,N_4449,N_4146);
nor U4876 (N_4876,N_4197,N_4405);
or U4877 (N_4877,N_4115,N_4112);
or U4878 (N_4878,N_4173,N_4419);
nor U4879 (N_4879,N_4183,N_4246);
nand U4880 (N_4880,N_4277,N_4048);
and U4881 (N_4881,N_4271,N_4345);
or U4882 (N_4882,N_4420,N_4498);
nand U4883 (N_4883,N_4494,N_4053);
xnor U4884 (N_4884,N_4134,N_4371);
or U4885 (N_4885,N_4104,N_4244);
nor U4886 (N_4886,N_4453,N_4364);
nand U4887 (N_4887,N_4154,N_4448);
or U4888 (N_4888,N_4344,N_4293);
or U4889 (N_4889,N_4368,N_4083);
and U4890 (N_4890,N_4314,N_4407);
and U4891 (N_4891,N_4440,N_4204);
nand U4892 (N_4892,N_4373,N_4121);
nor U4893 (N_4893,N_4318,N_4273);
or U4894 (N_4894,N_4335,N_4271);
nor U4895 (N_4895,N_4361,N_4039);
nand U4896 (N_4896,N_4420,N_4017);
nand U4897 (N_4897,N_4105,N_4089);
or U4898 (N_4898,N_4014,N_4156);
nand U4899 (N_4899,N_4418,N_4282);
or U4900 (N_4900,N_4052,N_4241);
xnor U4901 (N_4901,N_4041,N_4375);
and U4902 (N_4902,N_4409,N_4048);
nand U4903 (N_4903,N_4435,N_4478);
nand U4904 (N_4904,N_4464,N_4150);
nand U4905 (N_4905,N_4441,N_4034);
nor U4906 (N_4906,N_4306,N_4192);
or U4907 (N_4907,N_4471,N_4338);
or U4908 (N_4908,N_4377,N_4013);
or U4909 (N_4909,N_4089,N_4213);
and U4910 (N_4910,N_4266,N_4475);
and U4911 (N_4911,N_4471,N_4390);
nor U4912 (N_4912,N_4266,N_4125);
nand U4913 (N_4913,N_4069,N_4004);
nor U4914 (N_4914,N_4248,N_4423);
and U4915 (N_4915,N_4171,N_4177);
nor U4916 (N_4916,N_4388,N_4008);
nand U4917 (N_4917,N_4011,N_4101);
nor U4918 (N_4918,N_4293,N_4046);
nor U4919 (N_4919,N_4486,N_4110);
or U4920 (N_4920,N_4249,N_4334);
nand U4921 (N_4921,N_4490,N_4175);
nand U4922 (N_4922,N_4024,N_4012);
nor U4923 (N_4923,N_4160,N_4167);
or U4924 (N_4924,N_4439,N_4070);
nor U4925 (N_4925,N_4303,N_4461);
nor U4926 (N_4926,N_4403,N_4333);
or U4927 (N_4927,N_4419,N_4152);
xnor U4928 (N_4928,N_4052,N_4072);
nor U4929 (N_4929,N_4009,N_4433);
xor U4930 (N_4930,N_4042,N_4229);
xnor U4931 (N_4931,N_4000,N_4102);
or U4932 (N_4932,N_4320,N_4048);
nor U4933 (N_4933,N_4246,N_4131);
xor U4934 (N_4934,N_4237,N_4277);
and U4935 (N_4935,N_4154,N_4334);
or U4936 (N_4936,N_4366,N_4142);
or U4937 (N_4937,N_4147,N_4415);
and U4938 (N_4938,N_4484,N_4007);
xor U4939 (N_4939,N_4200,N_4120);
or U4940 (N_4940,N_4221,N_4149);
or U4941 (N_4941,N_4333,N_4195);
xor U4942 (N_4942,N_4216,N_4001);
xnor U4943 (N_4943,N_4300,N_4367);
and U4944 (N_4944,N_4093,N_4485);
and U4945 (N_4945,N_4321,N_4249);
nand U4946 (N_4946,N_4133,N_4321);
nand U4947 (N_4947,N_4406,N_4388);
and U4948 (N_4948,N_4354,N_4406);
and U4949 (N_4949,N_4014,N_4062);
or U4950 (N_4950,N_4208,N_4463);
nor U4951 (N_4951,N_4222,N_4039);
and U4952 (N_4952,N_4371,N_4487);
or U4953 (N_4953,N_4047,N_4368);
nand U4954 (N_4954,N_4011,N_4118);
nor U4955 (N_4955,N_4175,N_4461);
and U4956 (N_4956,N_4193,N_4318);
nor U4957 (N_4957,N_4188,N_4488);
nor U4958 (N_4958,N_4404,N_4430);
nand U4959 (N_4959,N_4426,N_4266);
or U4960 (N_4960,N_4487,N_4014);
and U4961 (N_4961,N_4149,N_4006);
nor U4962 (N_4962,N_4235,N_4263);
nor U4963 (N_4963,N_4253,N_4288);
xor U4964 (N_4964,N_4231,N_4153);
or U4965 (N_4965,N_4215,N_4400);
xnor U4966 (N_4966,N_4268,N_4302);
nor U4967 (N_4967,N_4018,N_4038);
nor U4968 (N_4968,N_4018,N_4312);
and U4969 (N_4969,N_4132,N_4153);
and U4970 (N_4970,N_4423,N_4142);
nand U4971 (N_4971,N_4136,N_4242);
nor U4972 (N_4972,N_4014,N_4455);
xor U4973 (N_4973,N_4012,N_4164);
and U4974 (N_4974,N_4482,N_4409);
nand U4975 (N_4975,N_4348,N_4146);
and U4976 (N_4976,N_4277,N_4131);
nor U4977 (N_4977,N_4419,N_4094);
and U4978 (N_4978,N_4050,N_4057);
nor U4979 (N_4979,N_4195,N_4049);
nor U4980 (N_4980,N_4017,N_4461);
or U4981 (N_4981,N_4096,N_4394);
nand U4982 (N_4982,N_4088,N_4202);
and U4983 (N_4983,N_4245,N_4278);
or U4984 (N_4984,N_4186,N_4216);
xnor U4985 (N_4985,N_4074,N_4473);
or U4986 (N_4986,N_4350,N_4368);
nor U4987 (N_4987,N_4203,N_4274);
nor U4988 (N_4988,N_4157,N_4156);
or U4989 (N_4989,N_4289,N_4204);
nand U4990 (N_4990,N_4252,N_4341);
or U4991 (N_4991,N_4203,N_4284);
and U4992 (N_4992,N_4351,N_4304);
and U4993 (N_4993,N_4050,N_4326);
nor U4994 (N_4994,N_4085,N_4454);
or U4995 (N_4995,N_4145,N_4281);
or U4996 (N_4996,N_4329,N_4436);
nor U4997 (N_4997,N_4479,N_4148);
xor U4998 (N_4998,N_4467,N_4365);
nor U4999 (N_4999,N_4187,N_4233);
or UO_0 (O_0,N_4726,N_4811);
or UO_1 (O_1,N_4847,N_4630);
nor UO_2 (O_2,N_4517,N_4607);
or UO_3 (O_3,N_4547,N_4575);
or UO_4 (O_4,N_4609,N_4602);
nor UO_5 (O_5,N_4776,N_4754);
nand UO_6 (O_6,N_4694,N_4786);
nor UO_7 (O_7,N_4533,N_4621);
nor UO_8 (O_8,N_4833,N_4854);
or UO_9 (O_9,N_4532,N_4545);
nand UO_10 (O_10,N_4855,N_4873);
and UO_11 (O_11,N_4573,N_4821);
nor UO_12 (O_12,N_4942,N_4593);
xor UO_13 (O_13,N_4742,N_4586);
or UO_14 (O_14,N_4522,N_4973);
or UO_15 (O_15,N_4947,N_4616);
or UO_16 (O_16,N_4772,N_4600);
or UO_17 (O_17,N_4769,N_4709);
and UO_18 (O_18,N_4543,N_4687);
nand UO_19 (O_19,N_4552,N_4686);
nand UO_20 (O_20,N_4813,N_4800);
and UO_21 (O_21,N_4968,N_4915);
nor UO_22 (O_22,N_4967,N_4583);
nand UO_23 (O_23,N_4585,N_4566);
and UO_24 (O_24,N_4841,N_4713);
and UO_25 (O_25,N_4678,N_4738);
xnor UO_26 (O_26,N_4768,N_4832);
nand UO_27 (O_27,N_4749,N_4679);
and UO_28 (O_28,N_4682,N_4622);
nor UO_29 (O_29,N_4730,N_4565);
or UO_30 (O_30,N_4605,N_4712);
and UO_31 (O_31,N_4906,N_4657);
nand UO_32 (O_32,N_4755,N_4771);
xnor UO_33 (O_33,N_4893,N_4928);
and UO_34 (O_34,N_4684,N_4627);
xor UO_35 (O_35,N_4703,N_4674);
xnor UO_36 (O_36,N_4736,N_4719);
or UO_37 (O_37,N_4874,N_4676);
nand UO_38 (O_38,N_4564,N_4596);
nor UO_39 (O_39,N_4909,N_4704);
nand UO_40 (O_40,N_4670,N_4710);
nor UO_41 (O_41,N_4817,N_4628);
nand UO_42 (O_42,N_4883,N_4810);
nand UO_43 (O_43,N_4828,N_4639);
and UO_44 (O_44,N_4538,N_4519);
or UO_45 (O_45,N_4775,N_4721);
or UO_46 (O_46,N_4954,N_4509);
or UO_47 (O_47,N_4886,N_4572);
and UO_48 (O_48,N_4556,N_4830);
and UO_49 (O_49,N_4939,N_4969);
or UO_50 (O_50,N_4633,N_4515);
or UO_51 (O_51,N_4580,N_4912);
nor UO_52 (O_52,N_4598,N_4680);
and UO_53 (O_53,N_4534,N_4878);
nand UO_54 (O_54,N_4661,N_4784);
or UO_55 (O_55,N_4924,N_4945);
xor UO_56 (O_56,N_4812,N_4595);
nor UO_57 (O_57,N_4988,N_4646);
xor UO_58 (O_58,N_4570,N_4503);
nor UO_59 (O_59,N_4625,N_4783);
nand UO_60 (O_60,N_4880,N_4579);
nand UO_61 (O_61,N_4528,N_4706);
nand UO_62 (O_62,N_4508,N_4798);
nand UO_63 (O_63,N_4884,N_4727);
nor UO_64 (O_64,N_4871,N_4999);
and UO_65 (O_65,N_4685,N_4774);
nand UO_66 (O_66,N_4761,N_4864);
nor UO_67 (O_67,N_4756,N_4950);
or UO_68 (O_68,N_4904,N_4569);
nor UO_69 (O_69,N_4765,N_4737);
xnor UO_70 (O_70,N_4796,N_4531);
or UO_71 (O_71,N_4677,N_4716);
nor UO_72 (O_72,N_4663,N_4606);
xnor UO_73 (O_73,N_4699,N_4665);
nand UO_74 (O_74,N_4717,N_4513);
and UO_75 (O_75,N_4526,N_4914);
xor UO_76 (O_76,N_4599,N_4848);
nand UO_77 (O_77,N_4731,N_4695);
nand UO_78 (O_78,N_4501,N_4882);
or UO_79 (O_79,N_4591,N_4923);
nor UO_80 (O_80,N_4529,N_4707);
nor UO_81 (O_81,N_4885,N_4637);
xor UO_82 (O_82,N_4838,N_4766);
nor UO_83 (O_83,N_4753,N_4620);
or UO_84 (O_84,N_4908,N_4524);
nand UO_85 (O_85,N_4943,N_4782);
or UO_86 (O_86,N_4758,N_4669);
nand UO_87 (O_87,N_4649,N_4729);
or UO_88 (O_88,N_4732,N_4851);
and UO_89 (O_89,N_4842,N_4636);
nor UO_90 (O_90,N_4725,N_4525);
and UO_91 (O_91,N_4852,N_4592);
nand UO_92 (O_92,N_4807,N_4859);
and UO_93 (O_93,N_4617,N_4683);
nand UO_94 (O_94,N_4582,N_4613);
or UO_95 (O_95,N_4930,N_4819);
or UO_96 (O_96,N_4964,N_4597);
and UO_97 (O_97,N_4803,N_4820);
nand UO_98 (O_98,N_4963,N_4808);
nand UO_99 (O_99,N_4926,N_4751);
nor UO_100 (O_100,N_4916,N_4658);
and UO_101 (O_101,N_4589,N_4619);
nand UO_102 (O_102,N_4603,N_4972);
xnor UO_103 (O_103,N_4558,N_4922);
nor UO_104 (O_104,N_4938,N_4905);
nand UO_105 (O_105,N_4764,N_4568);
nand UO_106 (O_106,N_4701,N_4809);
or UO_107 (O_107,N_4601,N_4512);
and UO_108 (O_108,N_4734,N_4872);
nand UO_109 (O_109,N_4911,N_4890);
or UO_110 (O_110,N_4588,N_4994);
nand UO_111 (O_111,N_4790,N_4850);
or UO_112 (O_112,N_4671,N_4594);
nor UO_113 (O_113,N_4611,N_4961);
and UO_114 (O_114,N_4634,N_4535);
nor UO_115 (O_115,N_4760,N_4574);
and UO_116 (O_116,N_4971,N_4590);
nand UO_117 (O_117,N_4561,N_4826);
xnor UO_118 (O_118,N_4935,N_4577);
xor UO_119 (O_119,N_4741,N_4976);
xnor UO_120 (O_120,N_4921,N_4853);
or UO_121 (O_121,N_4759,N_4720);
nand UO_122 (O_122,N_4780,N_4693);
nand UO_123 (O_123,N_4511,N_4998);
nor UO_124 (O_124,N_4788,N_4949);
nand UO_125 (O_125,N_4844,N_4739);
and UO_126 (O_126,N_4746,N_4762);
nand UO_127 (O_127,N_4673,N_4527);
or UO_128 (O_128,N_4516,N_4974);
or UO_129 (O_129,N_4542,N_4696);
and UO_130 (O_130,N_4640,N_4518);
nand UO_131 (O_131,N_4691,N_4801);
nand UO_132 (O_132,N_4689,N_4551);
xor UO_133 (O_133,N_4578,N_4690);
nand UO_134 (O_134,N_4857,N_4668);
or UO_135 (O_135,N_4959,N_4692);
nand UO_136 (O_136,N_4925,N_4523);
or UO_137 (O_137,N_4814,N_4941);
and UO_138 (O_138,N_4645,N_4675);
nand UO_139 (O_139,N_4541,N_4553);
or UO_140 (O_140,N_4787,N_4555);
or UO_141 (O_141,N_4879,N_4867);
and UO_142 (O_142,N_4940,N_4934);
nor UO_143 (O_143,N_4987,N_4887);
nor UO_144 (O_144,N_4835,N_4724);
nor UO_145 (O_145,N_4910,N_4777);
or UO_146 (O_146,N_4650,N_4948);
and UO_147 (O_147,N_4608,N_4789);
nor UO_148 (O_148,N_4865,N_4818);
nand UO_149 (O_149,N_4979,N_4767);
or UO_150 (O_150,N_4831,N_4757);
nor UO_151 (O_151,N_4894,N_4791);
nand UO_152 (O_152,N_4951,N_4839);
and UO_153 (O_153,N_4986,N_4919);
nor UO_154 (O_154,N_4554,N_4576);
and UO_155 (O_155,N_4507,N_4795);
xnor UO_156 (O_156,N_4648,N_4877);
and UO_157 (O_157,N_4514,N_4697);
or UO_158 (O_158,N_4660,N_4846);
nor UO_159 (O_159,N_4824,N_4952);
nor UO_160 (O_160,N_4654,N_4953);
and UO_161 (O_161,N_4849,N_4980);
xnor UO_162 (O_162,N_4505,N_4977);
nor UO_163 (O_163,N_4891,N_4642);
or UO_164 (O_164,N_4702,N_4993);
nor UO_165 (O_165,N_4723,N_4546);
nor UO_166 (O_166,N_4632,N_4785);
or UO_167 (O_167,N_4700,N_4748);
or UO_168 (O_168,N_4770,N_4889);
and UO_169 (O_169,N_4548,N_4825);
nor UO_170 (O_170,N_4714,N_4705);
nor UO_171 (O_171,N_4792,N_4664);
or UO_172 (O_172,N_4781,N_4897);
nand UO_173 (O_173,N_4983,N_4900);
and UO_174 (O_174,N_4965,N_4957);
and UO_175 (O_175,N_4711,N_4866);
nand UO_176 (O_176,N_4823,N_4927);
nand UO_177 (O_177,N_4733,N_4614);
nor UO_178 (O_178,N_4740,N_4653);
nor UO_179 (O_179,N_4822,N_4918);
or UO_180 (O_180,N_4862,N_4985);
nor UO_181 (O_181,N_4715,N_4895);
nor UO_182 (O_182,N_4735,N_4802);
and UO_183 (O_183,N_4562,N_4837);
and UO_184 (O_184,N_4655,N_4989);
nor UO_185 (O_185,N_4946,N_4604);
or UO_186 (O_186,N_4991,N_4520);
nor UO_187 (O_187,N_4698,N_4500);
and UO_188 (O_188,N_4861,N_4662);
and UO_189 (O_189,N_4629,N_4920);
nor UO_190 (O_190,N_4995,N_4799);
xnor UO_191 (O_191,N_4840,N_4688);
or UO_192 (O_192,N_4647,N_4827);
nand UO_193 (O_193,N_4763,N_4931);
and UO_194 (O_194,N_4876,N_4936);
nand UO_195 (O_195,N_4960,N_4843);
xor UO_196 (O_196,N_4635,N_4610);
xor UO_197 (O_197,N_4681,N_4899);
nor UO_198 (O_198,N_4937,N_4978);
nand UO_199 (O_199,N_4745,N_4868);
nor UO_200 (O_200,N_4903,N_4997);
nor UO_201 (O_201,N_4863,N_4815);
or UO_202 (O_202,N_4656,N_4750);
or UO_203 (O_203,N_4990,N_4587);
nor UO_204 (O_204,N_4530,N_4536);
or UO_205 (O_205,N_4672,N_4956);
or UO_206 (O_206,N_4537,N_4521);
and UO_207 (O_207,N_4722,N_4626);
nor UO_208 (O_208,N_4506,N_4966);
and UO_209 (O_209,N_4917,N_4623);
and UO_210 (O_210,N_4984,N_4638);
and UO_211 (O_211,N_4631,N_4870);
and UO_212 (O_212,N_4540,N_4567);
or UO_213 (O_213,N_4896,N_4806);
nor UO_214 (O_214,N_4743,N_4902);
xor UO_215 (O_215,N_4718,N_4955);
or UO_216 (O_216,N_4571,N_4797);
xnor UO_217 (O_217,N_4652,N_4898);
and UO_218 (O_218,N_4641,N_4901);
nor UO_219 (O_219,N_4779,N_4982);
and UO_220 (O_220,N_4563,N_4856);
nor UO_221 (O_221,N_4667,N_4962);
and UO_222 (O_222,N_4612,N_4504);
or UO_223 (O_223,N_4744,N_4869);
or UO_224 (O_224,N_4581,N_4793);
and UO_225 (O_225,N_4958,N_4752);
or UO_226 (O_226,N_4996,N_4913);
nand UO_227 (O_227,N_4539,N_4549);
nor UO_228 (O_228,N_4666,N_4624);
xnor UO_229 (O_229,N_4975,N_4773);
or UO_230 (O_230,N_4805,N_4502);
nand UO_231 (O_231,N_4643,N_4659);
or UO_232 (O_232,N_4875,N_4615);
or UO_233 (O_233,N_4747,N_4584);
nor UO_234 (O_234,N_4860,N_4929);
nand UO_235 (O_235,N_4550,N_4944);
or UO_236 (O_236,N_4644,N_4892);
or UO_237 (O_237,N_4981,N_4933);
nand UO_238 (O_238,N_4510,N_4858);
or UO_239 (O_239,N_4794,N_4992);
or UO_240 (O_240,N_4932,N_4651);
and UO_241 (O_241,N_4829,N_4834);
and UO_242 (O_242,N_4708,N_4804);
and UO_243 (O_243,N_4559,N_4888);
xnor UO_244 (O_244,N_4557,N_4970);
and UO_245 (O_245,N_4560,N_4816);
and UO_246 (O_246,N_4881,N_4728);
nor UO_247 (O_247,N_4907,N_4778);
xor UO_248 (O_248,N_4618,N_4836);
or UO_249 (O_249,N_4544,N_4845);
or UO_250 (O_250,N_4599,N_4640);
and UO_251 (O_251,N_4664,N_4839);
xnor UO_252 (O_252,N_4807,N_4874);
nand UO_253 (O_253,N_4922,N_4935);
nand UO_254 (O_254,N_4911,N_4929);
nand UO_255 (O_255,N_4999,N_4795);
nor UO_256 (O_256,N_4805,N_4908);
and UO_257 (O_257,N_4867,N_4892);
nor UO_258 (O_258,N_4866,N_4699);
xnor UO_259 (O_259,N_4569,N_4633);
nand UO_260 (O_260,N_4900,N_4986);
nand UO_261 (O_261,N_4670,N_4743);
and UO_262 (O_262,N_4671,N_4721);
nand UO_263 (O_263,N_4821,N_4553);
nand UO_264 (O_264,N_4677,N_4604);
nand UO_265 (O_265,N_4696,N_4544);
or UO_266 (O_266,N_4596,N_4830);
or UO_267 (O_267,N_4941,N_4992);
nand UO_268 (O_268,N_4538,N_4656);
and UO_269 (O_269,N_4508,N_4584);
and UO_270 (O_270,N_4720,N_4527);
or UO_271 (O_271,N_4798,N_4943);
and UO_272 (O_272,N_4506,N_4525);
xor UO_273 (O_273,N_4539,N_4523);
or UO_274 (O_274,N_4726,N_4944);
xor UO_275 (O_275,N_4652,N_4582);
nand UO_276 (O_276,N_4606,N_4600);
xor UO_277 (O_277,N_4584,N_4511);
nor UO_278 (O_278,N_4658,N_4512);
nand UO_279 (O_279,N_4517,N_4769);
and UO_280 (O_280,N_4972,N_4783);
nor UO_281 (O_281,N_4505,N_4817);
nor UO_282 (O_282,N_4918,N_4777);
nand UO_283 (O_283,N_4545,N_4756);
nor UO_284 (O_284,N_4750,N_4773);
or UO_285 (O_285,N_4957,N_4775);
nor UO_286 (O_286,N_4645,N_4575);
nor UO_287 (O_287,N_4911,N_4829);
or UO_288 (O_288,N_4878,N_4782);
xnor UO_289 (O_289,N_4778,N_4623);
xor UO_290 (O_290,N_4621,N_4562);
nor UO_291 (O_291,N_4602,N_4752);
nand UO_292 (O_292,N_4555,N_4725);
or UO_293 (O_293,N_4616,N_4595);
nor UO_294 (O_294,N_4929,N_4505);
and UO_295 (O_295,N_4972,N_4797);
xnor UO_296 (O_296,N_4593,N_4813);
or UO_297 (O_297,N_4627,N_4736);
xor UO_298 (O_298,N_4959,N_4728);
nand UO_299 (O_299,N_4905,N_4961);
and UO_300 (O_300,N_4776,N_4769);
nand UO_301 (O_301,N_4611,N_4590);
nand UO_302 (O_302,N_4709,N_4535);
and UO_303 (O_303,N_4527,N_4630);
or UO_304 (O_304,N_4903,N_4841);
nand UO_305 (O_305,N_4500,N_4731);
or UO_306 (O_306,N_4737,N_4871);
and UO_307 (O_307,N_4917,N_4978);
nor UO_308 (O_308,N_4535,N_4658);
or UO_309 (O_309,N_4664,N_4969);
nor UO_310 (O_310,N_4529,N_4699);
nand UO_311 (O_311,N_4884,N_4869);
nor UO_312 (O_312,N_4832,N_4683);
nand UO_313 (O_313,N_4595,N_4631);
nand UO_314 (O_314,N_4826,N_4897);
xnor UO_315 (O_315,N_4500,N_4583);
or UO_316 (O_316,N_4991,N_4899);
nor UO_317 (O_317,N_4579,N_4517);
xnor UO_318 (O_318,N_4885,N_4583);
nor UO_319 (O_319,N_4981,N_4536);
nor UO_320 (O_320,N_4535,N_4594);
and UO_321 (O_321,N_4576,N_4689);
or UO_322 (O_322,N_4523,N_4624);
nand UO_323 (O_323,N_4538,N_4793);
and UO_324 (O_324,N_4620,N_4781);
or UO_325 (O_325,N_4550,N_4785);
or UO_326 (O_326,N_4924,N_4819);
or UO_327 (O_327,N_4773,N_4923);
nor UO_328 (O_328,N_4683,N_4922);
or UO_329 (O_329,N_4518,N_4561);
nor UO_330 (O_330,N_4914,N_4747);
or UO_331 (O_331,N_4833,N_4656);
nand UO_332 (O_332,N_4619,N_4780);
nor UO_333 (O_333,N_4799,N_4936);
nor UO_334 (O_334,N_4724,N_4738);
and UO_335 (O_335,N_4705,N_4918);
or UO_336 (O_336,N_4721,N_4922);
or UO_337 (O_337,N_4557,N_4890);
nand UO_338 (O_338,N_4865,N_4819);
or UO_339 (O_339,N_4663,N_4556);
or UO_340 (O_340,N_4962,N_4555);
nand UO_341 (O_341,N_4784,N_4643);
xor UO_342 (O_342,N_4940,N_4913);
or UO_343 (O_343,N_4776,N_4901);
and UO_344 (O_344,N_4622,N_4744);
xnor UO_345 (O_345,N_4700,N_4697);
and UO_346 (O_346,N_4587,N_4642);
and UO_347 (O_347,N_4634,N_4591);
or UO_348 (O_348,N_4532,N_4679);
and UO_349 (O_349,N_4658,N_4615);
and UO_350 (O_350,N_4690,N_4641);
nor UO_351 (O_351,N_4919,N_4514);
nand UO_352 (O_352,N_4740,N_4929);
nor UO_353 (O_353,N_4922,N_4830);
nand UO_354 (O_354,N_4552,N_4742);
nand UO_355 (O_355,N_4552,N_4584);
or UO_356 (O_356,N_4893,N_4876);
xnor UO_357 (O_357,N_4785,N_4847);
nand UO_358 (O_358,N_4777,N_4965);
and UO_359 (O_359,N_4974,N_4862);
or UO_360 (O_360,N_4943,N_4842);
nand UO_361 (O_361,N_4667,N_4615);
and UO_362 (O_362,N_4953,N_4946);
and UO_363 (O_363,N_4872,N_4740);
xnor UO_364 (O_364,N_4523,N_4867);
nand UO_365 (O_365,N_4875,N_4912);
and UO_366 (O_366,N_4577,N_4586);
nor UO_367 (O_367,N_4654,N_4901);
nor UO_368 (O_368,N_4599,N_4616);
and UO_369 (O_369,N_4778,N_4667);
xnor UO_370 (O_370,N_4774,N_4749);
nor UO_371 (O_371,N_4619,N_4541);
nor UO_372 (O_372,N_4834,N_4961);
nand UO_373 (O_373,N_4548,N_4900);
and UO_374 (O_374,N_4727,N_4789);
nand UO_375 (O_375,N_4921,N_4690);
nor UO_376 (O_376,N_4961,N_4908);
nor UO_377 (O_377,N_4523,N_4966);
xor UO_378 (O_378,N_4964,N_4640);
xnor UO_379 (O_379,N_4706,N_4786);
or UO_380 (O_380,N_4579,N_4560);
and UO_381 (O_381,N_4839,N_4548);
nand UO_382 (O_382,N_4867,N_4556);
nand UO_383 (O_383,N_4635,N_4876);
or UO_384 (O_384,N_4931,N_4687);
and UO_385 (O_385,N_4716,N_4500);
or UO_386 (O_386,N_4847,N_4659);
xor UO_387 (O_387,N_4566,N_4870);
nor UO_388 (O_388,N_4858,N_4544);
and UO_389 (O_389,N_4663,N_4584);
or UO_390 (O_390,N_4934,N_4535);
and UO_391 (O_391,N_4730,N_4503);
nor UO_392 (O_392,N_4707,N_4981);
and UO_393 (O_393,N_4520,N_4611);
or UO_394 (O_394,N_4780,N_4778);
or UO_395 (O_395,N_4915,N_4793);
and UO_396 (O_396,N_4512,N_4815);
and UO_397 (O_397,N_4617,N_4641);
nand UO_398 (O_398,N_4558,N_4686);
nor UO_399 (O_399,N_4868,N_4666);
xor UO_400 (O_400,N_4591,N_4750);
nor UO_401 (O_401,N_4623,N_4575);
and UO_402 (O_402,N_4694,N_4891);
nor UO_403 (O_403,N_4663,N_4505);
nand UO_404 (O_404,N_4686,N_4652);
or UO_405 (O_405,N_4937,N_4702);
and UO_406 (O_406,N_4808,N_4913);
xnor UO_407 (O_407,N_4807,N_4911);
nand UO_408 (O_408,N_4594,N_4540);
or UO_409 (O_409,N_4562,N_4965);
nand UO_410 (O_410,N_4592,N_4851);
nor UO_411 (O_411,N_4522,N_4511);
nor UO_412 (O_412,N_4623,N_4857);
nor UO_413 (O_413,N_4733,N_4926);
nor UO_414 (O_414,N_4656,N_4773);
or UO_415 (O_415,N_4866,N_4951);
and UO_416 (O_416,N_4822,N_4962);
and UO_417 (O_417,N_4614,N_4840);
nor UO_418 (O_418,N_4841,N_4833);
and UO_419 (O_419,N_4816,N_4550);
nand UO_420 (O_420,N_4514,N_4952);
or UO_421 (O_421,N_4715,N_4899);
nor UO_422 (O_422,N_4884,N_4766);
and UO_423 (O_423,N_4603,N_4635);
nor UO_424 (O_424,N_4838,N_4772);
and UO_425 (O_425,N_4555,N_4920);
nor UO_426 (O_426,N_4572,N_4878);
or UO_427 (O_427,N_4810,N_4893);
nor UO_428 (O_428,N_4571,N_4590);
nor UO_429 (O_429,N_4563,N_4669);
nor UO_430 (O_430,N_4633,N_4749);
xnor UO_431 (O_431,N_4680,N_4564);
or UO_432 (O_432,N_4640,N_4662);
nand UO_433 (O_433,N_4846,N_4778);
and UO_434 (O_434,N_4500,N_4825);
nor UO_435 (O_435,N_4819,N_4679);
nor UO_436 (O_436,N_4573,N_4926);
nand UO_437 (O_437,N_4538,N_4543);
nor UO_438 (O_438,N_4742,N_4584);
or UO_439 (O_439,N_4850,N_4854);
and UO_440 (O_440,N_4523,N_4720);
or UO_441 (O_441,N_4992,N_4688);
xor UO_442 (O_442,N_4681,N_4664);
and UO_443 (O_443,N_4590,N_4976);
nand UO_444 (O_444,N_4803,N_4832);
or UO_445 (O_445,N_4869,N_4672);
nand UO_446 (O_446,N_4817,N_4913);
nand UO_447 (O_447,N_4540,N_4608);
nand UO_448 (O_448,N_4708,N_4732);
nor UO_449 (O_449,N_4903,N_4515);
nand UO_450 (O_450,N_4692,N_4501);
or UO_451 (O_451,N_4690,N_4679);
xnor UO_452 (O_452,N_4507,N_4866);
nor UO_453 (O_453,N_4858,N_4603);
and UO_454 (O_454,N_4691,N_4757);
and UO_455 (O_455,N_4974,N_4547);
or UO_456 (O_456,N_4577,N_4849);
nand UO_457 (O_457,N_4976,N_4991);
nor UO_458 (O_458,N_4531,N_4766);
or UO_459 (O_459,N_4681,N_4507);
xnor UO_460 (O_460,N_4602,N_4687);
xnor UO_461 (O_461,N_4752,N_4504);
or UO_462 (O_462,N_4782,N_4883);
nand UO_463 (O_463,N_4855,N_4725);
and UO_464 (O_464,N_4789,N_4658);
or UO_465 (O_465,N_4669,N_4532);
xor UO_466 (O_466,N_4668,N_4579);
xnor UO_467 (O_467,N_4845,N_4694);
or UO_468 (O_468,N_4895,N_4722);
nand UO_469 (O_469,N_4790,N_4582);
and UO_470 (O_470,N_4906,N_4636);
nor UO_471 (O_471,N_4916,N_4621);
and UO_472 (O_472,N_4853,N_4634);
and UO_473 (O_473,N_4598,N_4900);
nand UO_474 (O_474,N_4903,N_4500);
and UO_475 (O_475,N_4596,N_4553);
or UO_476 (O_476,N_4796,N_4748);
nor UO_477 (O_477,N_4798,N_4832);
nor UO_478 (O_478,N_4603,N_4563);
nand UO_479 (O_479,N_4545,N_4675);
nand UO_480 (O_480,N_4908,N_4932);
nand UO_481 (O_481,N_4667,N_4675);
and UO_482 (O_482,N_4932,N_4757);
and UO_483 (O_483,N_4842,N_4731);
nand UO_484 (O_484,N_4930,N_4857);
xnor UO_485 (O_485,N_4923,N_4605);
and UO_486 (O_486,N_4544,N_4798);
and UO_487 (O_487,N_4633,N_4947);
and UO_488 (O_488,N_4890,N_4717);
or UO_489 (O_489,N_4936,N_4814);
or UO_490 (O_490,N_4637,N_4533);
or UO_491 (O_491,N_4985,N_4531);
and UO_492 (O_492,N_4872,N_4975);
xor UO_493 (O_493,N_4970,N_4778);
nand UO_494 (O_494,N_4634,N_4873);
nor UO_495 (O_495,N_4818,N_4508);
nor UO_496 (O_496,N_4593,N_4843);
or UO_497 (O_497,N_4845,N_4751);
and UO_498 (O_498,N_4542,N_4979);
xnor UO_499 (O_499,N_4635,N_4818);
or UO_500 (O_500,N_4505,N_4995);
and UO_501 (O_501,N_4683,N_4983);
nor UO_502 (O_502,N_4625,N_4948);
nor UO_503 (O_503,N_4578,N_4618);
nand UO_504 (O_504,N_4895,N_4505);
and UO_505 (O_505,N_4736,N_4544);
nor UO_506 (O_506,N_4901,N_4948);
or UO_507 (O_507,N_4594,N_4661);
and UO_508 (O_508,N_4748,N_4980);
nand UO_509 (O_509,N_4705,N_4921);
and UO_510 (O_510,N_4887,N_4833);
nand UO_511 (O_511,N_4725,N_4506);
nand UO_512 (O_512,N_4953,N_4564);
or UO_513 (O_513,N_4897,N_4685);
nand UO_514 (O_514,N_4705,N_4542);
nand UO_515 (O_515,N_4621,N_4585);
and UO_516 (O_516,N_4968,N_4801);
and UO_517 (O_517,N_4891,N_4977);
and UO_518 (O_518,N_4968,N_4725);
nand UO_519 (O_519,N_4824,N_4620);
or UO_520 (O_520,N_4962,N_4558);
and UO_521 (O_521,N_4902,N_4703);
and UO_522 (O_522,N_4807,N_4724);
nor UO_523 (O_523,N_4874,N_4526);
nor UO_524 (O_524,N_4814,N_4859);
nand UO_525 (O_525,N_4627,N_4614);
nand UO_526 (O_526,N_4935,N_4750);
xnor UO_527 (O_527,N_4645,N_4589);
nand UO_528 (O_528,N_4924,N_4533);
nand UO_529 (O_529,N_4965,N_4676);
or UO_530 (O_530,N_4653,N_4580);
nand UO_531 (O_531,N_4584,N_4514);
nand UO_532 (O_532,N_4855,N_4517);
nand UO_533 (O_533,N_4644,N_4757);
nor UO_534 (O_534,N_4999,N_4720);
or UO_535 (O_535,N_4584,N_4896);
and UO_536 (O_536,N_4932,N_4866);
xnor UO_537 (O_537,N_4720,N_4808);
or UO_538 (O_538,N_4857,N_4772);
nand UO_539 (O_539,N_4790,N_4856);
and UO_540 (O_540,N_4504,N_4746);
and UO_541 (O_541,N_4792,N_4966);
or UO_542 (O_542,N_4920,N_4615);
and UO_543 (O_543,N_4763,N_4814);
nor UO_544 (O_544,N_4662,N_4607);
xnor UO_545 (O_545,N_4738,N_4870);
nand UO_546 (O_546,N_4634,N_4625);
or UO_547 (O_547,N_4650,N_4708);
or UO_548 (O_548,N_4592,N_4528);
and UO_549 (O_549,N_4818,N_4676);
and UO_550 (O_550,N_4732,N_4650);
nor UO_551 (O_551,N_4648,N_4980);
nor UO_552 (O_552,N_4800,N_4865);
nand UO_553 (O_553,N_4870,N_4657);
nor UO_554 (O_554,N_4798,N_4937);
nor UO_555 (O_555,N_4977,N_4954);
xnor UO_556 (O_556,N_4579,N_4630);
nand UO_557 (O_557,N_4508,N_4937);
nand UO_558 (O_558,N_4558,N_4675);
and UO_559 (O_559,N_4711,N_4768);
xnor UO_560 (O_560,N_4615,N_4585);
and UO_561 (O_561,N_4552,N_4531);
nor UO_562 (O_562,N_4916,N_4735);
nor UO_563 (O_563,N_4702,N_4586);
or UO_564 (O_564,N_4643,N_4745);
nand UO_565 (O_565,N_4657,N_4889);
nand UO_566 (O_566,N_4828,N_4712);
or UO_567 (O_567,N_4540,N_4983);
and UO_568 (O_568,N_4628,N_4553);
nor UO_569 (O_569,N_4883,N_4974);
nand UO_570 (O_570,N_4568,N_4631);
nand UO_571 (O_571,N_4560,N_4621);
and UO_572 (O_572,N_4673,N_4754);
nand UO_573 (O_573,N_4902,N_4985);
nand UO_574 (O_574,N_4867,N_4878);
nand UO_575 (O_575,N_4880,N_4846);
nand UO_576 (O_576,N_4513,N_4719);
nand UO_577 (O_577,N_4585,N_4691);
or UO_578 (O_578,N_4733,N_4609);
nor UO_579 (O_579,N_4554,N_4780);
nand UO_580 (O_580,N_4587,N_4502);
or UO_581 (O_581,N_4630,N_4609);
nand UO_582 (O_582,N_4722,N_4511);
nor UO_583 (O_583,N_4732,N_4634);
or UO_584 (O_584,N_4574,N_4741);
or UO_585 (O_585,N_4657,N_4757);
xor UO_586 (O_586,N_4512,N_4913);
nand UO_587 (O_587,N_4579,N_4591);
nor UO_588 (O_588,N_4682,N_4649);
nor UO_589 (O_589,N_4942,N_4729);
nand UO_590 (O_590,N_4712,N_4769);
and UO_591 (O_591,N_4670,N_4779);
nor UO_592 (O_592,N_4793,N_4642);
nor UO_593 (O_593,N_4765,N_4920);
nor UO_594 (O_594,N_4678,N_4628);
nor UO_595 (O_595,N_4535,N_4691);
and UO_596 (O_596,N_4665,N_4527);
nand UO_597 (O_597,N_4538,N_4993);
and UO_598 (O_598,N_4759,N_4934);
nand UO_599 (O_599,N_4811,N_4604);
nor UO_600 (O_600,N_4531,N_4966);
and UO_601 (O_601,N_4968,N_4667);
and UO_602 (O_602,N_4767,N_4805);
or UO_603 (O_603,N_4640,N_4815);
and UO_604 (O_604,N_4809,N_4859);
nand UO_605 (O_605,N_4723,N_4539);
and UO_606 (O_606,N_4909,N_4652);
or UO_607 (O_607,N_4626,N_4582);
and UO_608 (O_608,N_4576,N_4962);
xor UO_609 (O_609,N_4879,N_4543);
nor UO_610 (O_610,N_4720,N_4671);
nor UO_611 (O_611,N_4894,N_4679);
and UO_612 (O_612,N_4976,N_4599);
and UO_613 (O_613,N_4763,N_4898);
nor UO_614 (O_614,N_4730,N_4534);
nand UO_615 (O_615,N_4540,N_4684);
xnor UO_616 (O_616,N_4542,N_4903);
nor UO_617 (O_617,N_4839,N_4960);
and UO_618 (O_618,N_4607,N_4614);
nor UO_619 (O_619,N_4810,N_4755);
and UO_620 (O_620,N_4844,N_4859);
or UO_621 (O_621,N_4974,N_4976);
xnor UO_622 (O_622,N_4904,N_4997);
nand UO_623 (O_623,N_4829,N_4885);
and UO_624 (O_624,N_4596,N_4688);
nor UO_625 (O_625,N_4677,N_4771);
nor UO_626 (O_626,N_4883,N_4674);
nor UO_627 (O_627,N_4544,N_4689);
nand UO_628 (O_628,N_4756,N_4873);
xor UO_629 (O_629,N_4513,N_4688);
or UO_630 (O_630,N_4867,N_4959);
and UO_631 (O_631,N_4622,N_4811);
nand UO_632 (O_632,N_4951,N_4925);
nand UO_633 (O_633,N_4965,N_4673);
or UO_634 (O_634,N_4974,N_4989);
or UO_635 (O_635,N_4862,N_4679);
nand UO_636 (O_636,N_4763,N_4768);
nand UO_637 (O_637,N_4531,N_4505);
xnor UO_638 (O_638,N_4558,N_4875);
nor UO_639 (O_639,N_4878,N_4981);
and UO_640 (O_640,N_4852,N_4762);
xnor UO_641 (O_641,N_4603,N_4765);
and UO_642 (O_642,N_4860,N_4840);
or UO_643 (O_643,N_4898,N_4638);
or UO_644 (O_644,N_4702,N_4687);
or UO_645 (O_645,N_4542,N_4516);
or UO_646 (O_646,N_4652,N_4562);
nand UO_647 (O_647,N_4764,N_4930);
xnor UO_648 (O_648,N_4686,N_4799);
nand UO_649 (O_649,N_4543,N_4760);
nor UO_650 (O_650,N_4683,N_4504);
or UO_651 (O_651,N_4697,N_4976);
and UO_652 (O_652,N_4942,N_4508);
nor UO_653 (O_653,N_4647,N_4522);
or UO_654 (O_654,N_4547,N_4861);
or UO_655 (O_655,N_4747,N_4620);
nand UO_656 (O_656,N_4593,N_4639);
or UO_657 (O_657,N_4664,N_4976);
xor UO_658 (O_658,N_4902,N_4511);
and UO_659 (O_659,N_4887,N_4801);
or UO_660 (O_660,N_4872,N_4507);
nor UO_661 (O_661,N_4625,N_4864);
xor UO_662 (O_662,N_4800,N_4799);
nor UO_663 (O_663,N_4958,N_4797);
nand UO_664 (O_664,N_4804,N_4903);
and UO_665 (O_665,N_4683,N_4916);
or UO_666 (O_666,N_4706,N_4556);
nand UO_667 (O_667,N_4675,N_4878);
and UO_668 (O_668,N_4707,N_4701);
and UO_669 (O_669,N_4618,N_4553);
nor UO_670 (O_670,N_4657,N_4604);
nor UO_671 (O_671,N_4747,N_4692);
and UO_672 (O_672,N_4524,N_4986);
or UO_673 (O_673,N_4950,N_4534);
xnor UO_674 (O_674,N_4829,N_4666);
and UO_675 (O_675,N_4895,N_4501);
nor UO_676 (O_676,N_4573,N_4765);
nor UO_677 (O_677,N_4596,N_4640);
or UO_678 (O_678,N_4701,N_4708);
nand UO_679 (O_679,N_4814,N_4576);
or UO_680 (O_680,N_4522,N_4978);
or UO_681 (O_681,N_4734,N_4927);
or UO_682 (O_682,N_4935,N_4597);
nand UO_683 (O_683,N_4538,N_4764);
or UO_684 (O_684,N_4789,N_4852);
or UO_685 (O_685,N_4526,N_4987);
nand UO_686 (O_686,N_4889,N_4692);
and UO_687 (O_687,N_4528,N_4860);
or UO_688 (O_688,N_4855,N_4632);
nand UO_689 (O_689,N_4530,N_4818);
and UO_690 (O_690,N_4963,N_4760);
and UO_691 (O_691,N_4593,N_4869);
or UO_692 (O_692,N_4980,N_4890);
or UO_693 (O_693,N_4569,N_4807);
nor UO_694 (O_694,N_4662,N_4803);
or UO_695 (O_695,N_4589,N_4521);
xnor UO_696 (O_696,N_4957,N_4977);
xnor UO_697 (O_697,N_4602,N_4875);
and UO_698 (O_698,N_4663,N_4753);
or UO_699 (O_699,N_4951,N_4995);
nand UO_700 (O_700,N_4898,N_4648);
nor UO_701 (O_701,N_4748,N_4586);
or UO_702 (O_702,N_4593,N_4808);
or UO_703 (O_703,N_4588,N_4635);
and UO_704 (O_704,N_4866,N_4827);
nand UO_705 (O_705,N_4990,N_4692);
or UO_706 (O_706,N_4699,N_4673);
nand UO_707 (O_707,N_4879,N_4779);
and UO_708 (O_708,N_4815,N_4529);
or UO_709 (O_709,N_4699,N_4770);
or UO_710 (O_710,N_4827,N_4779);
or UO_711 (O_711,N_4919,N_4761);
or UO_712 (O_712,N_4745,N_4810);
nor UO_713 (O_713,N_4681,N_4580);
and UO_714 (O_714,N_4850,N_4573);
nor UO_715 (O_715,N_4847,N_4517);
or UO_716 (O_716,N_4983,N_4965);
or UO_717 (O_717,N_4605,N_4717);
nand UO_718 (O_718,N_4865,N_4870);
and UO_719 (O_719,N_4834,N_4913);
or UO_720 (O_720,N_4597,N_4947);
and UO_721 (O_721,N_4899,N_4582);
nor UO_722 (O_722,N_4588,N_4701);
nand UO_723 (O_723,N_4881,N_4800);
nand UO_724 (O_724,N_4839,N_4554);
nand UO_725 (O_725,N_4835,N_4865);
nor UO_726 (O_726,N_4984,N_4795);
nor UO_727 (O_727,N_4741,N_4672);
or UO_728 (O_728,N_4562,N_4946);
nor UO_729 (O_729,N_4802,N_4767);
nor UO_730 (O_730,N_4767,N_4704);
nand UO_731 (O_731,N_4997,N_4806);
and UO_732 (O_732,N_4857,N_4718);
or UO_733 (O_733,N_4886,N_4623);
nor UO_734 (O_734,N_4549,N_4897);
or UO_735 (O_735,N_4614,N_4984);
or UO_736 (O_736,N_4699,N_4737);
nor UO_737 (O_737,N_4837,N_4723);
and UO_738 (O_738,N_4959,N_4890);
nand UO_739 (O_739,N_4982,N_4825);
or UO_740 (O_740,N_4941,N_4724);
nand UO_741 (O_741,N_4978,N_4703);
and UO_742 (O_742,N_4861,N_4794);
and UO_743 (O_743,N_4881,N_4622);
xor UO_744 (O_744,N_4553,N_4994);
nand UO_745 (O_745,N_4945,N_4526);
or UO_746 (O_746,N_4683,N_4820);
or UO_747 (O_747,N_4594,N_4666);
and UO_748 (O_748,N_4933,N_4605);
nor UO_749 (O_749,N_4664,N_4525);
nand UO_750 (O_750,N_4532,N_4647);
nor UO_751 (O_751,N_4722,N_4910);
and UO_752 (O_752,N_4649,N_4961);
nor UO_753 (O_753,N_4867,N_4707);
nand UO_754 (O_754,N_4815,N_4623);
nor UO_755 (O_755,N_4965,N_4534);
or UO_756 (O_756,N_4824,N_4700);
nor UO_757 (O_757,N_4557,N_4652);
and UO_758 (O_758,N_4630,N_4728);
or UO_759 (O_759,N_4984,N_4794);
nor UO_760 (O_760,N_4594,N_4737);
nand UO_761 (O_761,N_4548,N_4635);
or UO_762 (O_762,N_4953,N_4733);
nor UO_763 (O_763,N_4928,N_4508);
or UO_764 (O_764,N_4742,N_4676);
nor UO_765 (O_765,N_4709,N_4582);
nand UO_766 (O_766,N_4677,N_4744);
nand UO_767 (O_767,N_4792,N_4510);
or UO_768 (O_768,N_4776,N_4822);
or UO_769 (O_769,N_4796,N_4860);
and UO_770 (O_770,N_4959,N_4523);
and UO_771 (O_771,N_4760,N_4875);
nand UO_772 (O_772,N_4545,N_4997);
nor UO_773 (O_773,N_4781,N_4706);
or UO_774 (O_774,N_4996,N_4801);
nand UO_775 (O_775,N_4641,N_4586);
or UO_776 (O_776,N_4585,N_4623);
or UO_777 (O_777,N_4763,N_4584);
and UO_778 (O_778,N_4555,N_4738);
or UO_779 (O_779,N_4821,N_4711);
nor UO_780 (O_780,N_4537,N_4863);
and UO_781 (O_781,N_4599,N_4778);
and UO_782 (O_782,N_4984,N_4572);
nand UO_783 (O_783,N_4786,N_4538);
or UO_784 (O_784,N_4726,N_4744);
nor UO_785 (O_785,N_4823,N_4993);
or UO_786 (O_786,N_4986,N_4843);
and UO_787 (O_787,N_4509,N_4638);
xnor UO_788 (O_788,N_4811,N_4594);
or UO_789 (O_789,N_4811,N_4590);
or UO_790 (O_790,N_4842,N_4618);
nor UO_791 (O_791,N_4781,N_4687);
or UO_792 (O_792,N_4737,N_4703);
nand UO_793 (O_793,N_4980,N_4633);
nor UO_794 (O_794,N_4746,N_4533);
or UO_795 (O_795,N_4909,N_4760);
and UO_796 (O_796,N_4851,N_4803);
or UO_797 (O_797,N_4691,N_4655);
nand UO_798 (O_798,N_4852,N_4543);
nand UO_799 (O_799,N_4515,N_4503);
or UO_800 (O_800,N_4699,N_4723);
nand UO_801 (O_801,N_4589,N_4519);
and UO_802 (O_802,N_4835,N_4530);
xnor UO_803 (O_803,N_4578,N_4835);
nand UO_804 (O_804,N_4922,N_4977);
or UO_805 (O_805,N_4588,N_4874);
or UO_806 (O_806,N_4919,N_4881);
nand UO_807 (O_807,N_4507,N_4885);
nor UO_808 (O_808,N_4619,N_4656);
nand UO_809 (O_809,N_4562,N_4761);
or UO_810 (O_810,N_4739,N_4673);
nand UO_811 (O_811,N_4998,N_4981);
and UO_812 (O_812,N_4643,N_4503);
or UO_813 (O_813,N_4825,N_4559);
and UO_814 (O_814,N_4887,N_4981);
and UO_815 (O_815,N_4747,N_4843);
or UO_816 (O_816,N_4930,N_4893);
or UO_817 (O_817,N_4583,N_4739);
and UO_818 (O_818,N_4931,N_4741);
nor UO_819 (O_819,N_4847,N_4541);
or UO_820 (O_820,N_4799,N_4909);
nand UO_821 (O_821,N_4819,N_4806);
xor UO_822 (O_822,N_4643,N_4507);
xnor UO_823 (O_823,N_4707,N_4773);
or UO_824 (O_824,N_4502,N_4621);
and UO_825 (O_825,N_4615,N_4851);
nor UO_826 (O_826,N_4823,N_4753);
nand UO_827 (O_827,N_4937,N_4969);
and UO_828 (O_828,N_4584,N_4823);
nor UO_829 (O_829,N_4534,N_4634);
nand UO_830 (O_830,N_4762,N_4831);
nor UO_831 (O_831,N_4997,N_4678);
nand UO_832 (O_832,N_4553,N_4555);
nor UO_833 (O_833,N_4745,N_4503);
or UO_834 (O_834,N_4585,N_4684);
nor UO_835 (O_835,N_4876,N_4896);
or UO_836 (O_836,N_4832,N_4624);
or UO_837 (O_837,N_4782,N_4701);
or UO_838 (O_838,N_4959,N_4706);
nand UO_839 (O_839,N_4635,N_4901);
nor UO_840 (O_840,N_4924,N_4768);
nor UO_841 (O_841,N_4613,N_4893);
or UO_842 (O_842,N_4812,N_4677);
nor UO_843 (O_843,N_4684,N_4706);
or UO_844 (O_844,N_4523,N_4545);
or UO_845 (O_845,N_4549,N_4612);
nand UO_846 (O_846,N_4669,N_4864);
or UO_847 (O_847,N_4936,N_4708);
nand UO_848 (O_848,N_4561,N_4726);
or UO_849 (O_849,N_4982,N_4592);
and UO_850 (O_850,N_4880,N_4765);
or UO_851 (O_851,N_4943,N_4860);
nand UO_852 (O_852,N_4965,N_4538);
nor UO_853 (O_853,N_4562,N_4855);
or UO_854 (O_854,N_4689,N_4502);
or UO_855 (O_855,N_4506,N_4742);
or UO_856 (O_856,N_4694,N_4651);
xnor UO_857 (O_857,N_4668,N_4972);
nand UO_858 (O_858,N_4884,N_4601);
xnor UO_859 (O_859,N_4753,N_4891);
nor UO_860 (O_860,N_4899,N_4864);
and UO_861 (O_861,N_4691,N_4608);
or UO_862 (O_862,N_4888,N_4627);
nor UO_863 (O_863,N_4729,N_4944);
or UO_864 (O_864,N_4921,N_4621);
or UO_865 (O_865,N_4841,N_4924);
and UO_866 (O_866,N_4748,N_4613);
and UO_867 (O_867,N_4668,N_4911);
nand UO_868 (O_868,N_4650,N_4595);
or UO_869 (O_869,N_4749,N_4557);
nor UO_870 (O_870,N_4873,N_4572);
or UO_871 (O_871,N_4933,N_4793);
and UO_872 (O_872,N_4969,N_4572);
or UO_873 (O_873,N_4817,N_4619);
nor UO_874 (O_874,N_4839,N_4893);
or UO_875 (O_875,N_4947,N_4670);
or UO_876 (O_876,N_4818,N_4570);
nor UO_877 (O_877,N_4736,N_4607);
nor UO_878 (O_878,N_4585,N_4671);
nor UO_879 (O_879,N_4576,N_4781);
and UO_880 (O_880,N_4767,N_4594);
nand UO_881 (O_881,N_4816,N_4644);
xor UO_882 (O_882,N_4807,N_4712);
and UO_883 (O_883,N_4753,N_4838);
nor UO_884 (O_884,N_4902,N_4509);
and UO_885 (O_885,N_4759,N_4688);
or UO_886 (O_886,N_4949,N_4695);
nor UO_887 (O_887,N_4759,N_4663);
and UO_888 (O_888,N_4632,N_4935);
nor UO_889 (O_889,N_4685,N_4840);
nor UO_890 (O_890,N_4794,N_4681);
nand UO_891 (O_891,N_4601,N_4619);
or UO_892 (O_892,N_4913,N_4915);
nand UO_893 (O_893,N_4974,N_4998);
or UO_894 (O_894,N_4649,N_4533);
nor UO_895 (O_895,N_4994,N_4738);
nor UO_896 (O_896,N_4959,N_4820);
nand UO_897 (O_897,N_4999,N_4542);
and UO_898 (O_898,N_4632,N_4795);
and UO_899 (O_899,N_4555,N_4822);
or UO_900 (O_900,N_4932,N_4725);
nor UO_901 (O_901,N_4927,N_4536);
nand UO_902 (O_902,N_4528,N_4943);
nor UO_903 (O_903,N_4702,N_4994);
nand UO_904 (O_904,N_4601,N_4514);
and UO_905 (O_905,N_4692,N_4890);
nor UO_906 (O_906,N_4568,N_4730);
or UO_907 (O_907,N_4517,N_4768);
nor UO_908 (O_908,N_4670,N_4549);
nor UO_909 (O_909,N_4812,N_4744);
nor UO_910 (O_910,N_4916,N_4791);
or UO_911 (O_911,N_4571,N_4957);
nor UO_912 (O_912,N_4775,N_4684);
and UO_913 (O_913,N_4823,N_4570);
and UO_914 (O_914,N_4555,N_4743);
nand UO_915 (O_915,N_4650,N_4958);
nor UO_916 (O_916,N_4539,N_4839);
and UO_917 (O_917,N_4893,N_4805);
and UO_918 (O_918,N_4531,N_4762);
nand UO_919 (O_919,N_4569,N_4777);
or UO_920 (O_920,N_4935,N_4593);
and UO_921 (O_921,N_4770,N_4557);
and UO_922 (O_922,N_4631,N_4767);
and UO_923 (O_923,N_4758,N_4616);
and UO_924 (O_924,N_4736,N_4825);
and UO_925 (O_925,N_4946,N_4919);
and UO_926 (O_926,N_4862,N_4515);
or UO_927 (O_927,N_4839,N_4858);
xnor UO_928 (O_928,N_4940,N_4948);
or UO_929 (O_929,N_4808,N_4983);
and UO_930 (O_930,N_4666,N_4605);
xnor UO_931 (O_931,N_4874,N_4633);
and UO_932 (O_932,N_4793,N_4999);
nor UO_933 (O_933,N_4889,N_4779);
and UO_934 (O_934,N_4566,N_4722);
nand UO_935 (O_935,N_4944,N_4986);
xor UO_936 (O_936,N_4950,N_4657);
nor UO_937 (O_937,N_4876,N_4942);
and UO_938 (O_938,N_4853,N_4644);
nor UO_939 (O_939,N_4920,N_4767);
and UO_940 (O_940,N_4692,N_4594);
nor UO_941 (O_941,N_4937,N_4806);
or UO_942 (O_942,N_4925,N_4768);
xor UO_943 (O_943,N_4941,N_4530);
and UO_944 (O_944,N_4911,N_4779);
nor UO_945 (O_945,N_4660,N_4779);
nand UO_946 (O_946,N_4804,N_4888);
or UO_947 (O_947,N_4612,N_4948);
nand UO_948 (O_948,N_4945,N_4587);
and UO_949 (O_949,N_4783,N_4664);
xor UO_950 (O_950,N_4513,N_4538);
xnor UO_951 (O_951,N_4573,N_4533);
and UO_952 (O_952,N_4577,N_4984);
and UO_953 (O_953,N_4703,N_4742);
and UO_954 (O_954,N_4825,N_4579);
nor UO_955 (O_955,N_4631,N_4588);
nand UO_956 (O_956,N_4945,N_4782);
and UO_957 (O_957,N_4757,N_4737);
or UO_958 (O_958,N_4623,N_4516);
and UO_959 (O_959,N_4764,N_4664);
nand UO_960 (O_960,N_4995,N_4960);
nand UO_961 (O_961,N_4904,N_4658);
nor UO_962 (O_962,N_4781,N_4977);
nor UO_963 (O_963,N_4693,N_4699);
nand UO_964 (O_964,N_4566,N_4954);
nor UO_965 (O_965,N_4829,N_4884);
nand UO_966 (O_966,N_4814,N_4962);
and UO_967 (O_967,N_4813,N_4872);
nor UO_968 (O_968,N_4896,N_4729);
nand UO_969 (O_969,N_4586,N_4961);
nor UO_970 (O_970,N_4570,N_4853);
nor UO_971 (O_971,N_4636,N_4553);
and UO_972 (O_972,N_4761,N_4911);
or UO_973 (O_973,N_4977,N_4571);
or UO_974 (O_974,N_4538,N_4960);
or UO_975 (O_975,N_4558,N_4606);
nor UO_976 (O_976,N_4577,N_4973);
nor UO_977 (O_977,N_4538,N_4818);
nor UO_978 (O_978,N_4936,N_4932);
and UO_979 (O_979,N_4598,N_4573);
nor UO_980 (O_980,N_4530,N_4601);
xor UO_981 (O_981,N_4576,N_4515);
or UO_982 (O_982,N_4657,N_4798);
nor UO_983 (O_983,N_4604,N_4522);
and UO_984 (O_984,N_4953,N_4569);
nand UO_985 (O_985,N_4582,N_4634);
nor UO_986 (O_986,N_4536,N_4639);
nand UO_987 (O_987,N_4821,N_4896);
nand UO_988 (O_988,N_4562,N_4696);
nor UO_989 (O_989,N_4795,N_4819);
and UO_990 (O_990,N_4628,N_4891);
and UO_991 (O_991,N_4992,N_4850);
or UO_992 (O_992,N_4735,N_4933);
xor UO_993 (O_993,N_4779,N_4590);
and UO_994 (O_994,N_4908,N_4544);
nand UO_995 (O_995,N_4828,N_4853);
nand UO_996 (O_996,N_4772,N_4972);
and UO_997 (O_997,N_4994,N_4515);
xor UO_998 (O_998,N_4526,N_4907);
nor UO_999 (O_999,N_4561,N_4866);
endmodule