module basic_750_5000_1000_10_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_609,In_331);
nor U1 (N_1,In_326,In_391);
nand U2 (N_2,In_124,In_102);
or U3 (N_3,In_670,In_573);
nor U4 (N_4,In_691,In_168);
and U5 (N_5,In_27,In_625);
or U6 (N_6,In_730,In_103);
or U7 (N_7,In_117,In_685);
nor U8 (N_8,In_204,In_133);
nor U9 (N_9,In_218,In_402);
and U10 (N_10,In_570,In_151);
nand U11 (N_11,In_558,In_644);
nand U12 (N_12,In_296,In_422);
nor U13 (N_13,In_661,In_456);
and U14 (N_14,In_543,In_189);
nor U15 (N_15,In_426,In_455);
or U16 (N_16,In_598,In_370);
nand U17 (N_17,In_638,In_488);
and U18 (N_18,In_528,In_327);
nor U19 (N_19,In_735,In_413);
and U20 (N_20,In_78,In_385);
nand U21 (N_21,In_510,In_574);
nand U22 (N_22,In_449,In_509);
or U23 (N_23,In_744,In_224);
or U24 (N_24,In_722,In_375);
nor U25 (N_25,In_495,In_2);
nand U26 (N_26,In_489,In_277);
and U27 (N_27,In_677,In_442);
nand U28 (N_28,In_653,In_158);
nor U29 (N_29,In_155,In_95);
or U30 (N_30,In_259,In_494);
nor U31 (N_31,In_471,In_244);
nand U32 (N_32,In_746,In_154);
nor U33 (N_33,In_59,In_407);
nor U34 (N_34,In_553,In_294);
or U35 (N_35,In_39,In_212);
nand U36 (N_36,In_203,In_517);
and U37 (N_37,In_571,In_40);
or U38 (N_38,In_79,In_539);
nor U39 (N_39,In_80,In_160);
or U40 (N_40,In_374,In_431);
nand U41 (N_41,In_701,In_605);
or U42 (N_42,In_633,In_30);
and U43 (N_43,In_172,In_502);
and U44 (N_44,In_436,In_187);
and U45 (N_45,In_513,In_284);
nand U46 (N_46,In_740,In_292);
nand U47 (N_47,In_324,In_679);
or U48 (N_48,In_467,In_427);
nand U49 (N_49,In_287,In_611);
nand U50 (N_50,In_288,In_134);
and U51 (N_51,In_560,In_188);
and U52 (N_52,In_641,In_429);
nor U53 (N_53,In_659,In_579);
and U54 (N_54,In_351,In_314);
nor U55 (N_55,In_388,In_330);
nor U56 (N_56,In_359,In_478);
and U57 (N_57,In_137,In_62);
nand U58 (N_58,In_480,In_69);
nand U59 (N_59,In_438,In_736);
and U60 (N_60,In_556,In_248);
nor U61 (N_61,In_651,In_497);
nor U62 (N_62,In_643,In_577);
and U63 (N_63,In_209,In_684);
or U64 (N_64,In_298,In_106);
or U65 (N_65,In_369,In_197);
and U66 (N_66,In_715,In_71);
and U67 (N_67,In_460,In_153);
nand U68 (N_68,In_390,In_26);
and U69 (N_69,In_262,In_462);
nand U70 (N_70,In_15,In_228);
and U71 (N_71,In_210,In_24);
and U72 (N_72,In_648,In_148);
and U73 (N_73,In_46,In_113);
or U74 (N_74,In_589,In_563);
and U75 (N_75,In_175,In_184);
nand U76 (N_76,In_635,In_306);
nand U77 (N_77,In_672,In_163);
and U78 (N_78,In_88,In_665);
nor U79 (N_79,In_530,In_475);
nor U80 (N_80,In_315,In_512);
and U81 (N_81,In_724,In_166);
nand U82 (N_82,In_161,In_663);
and U83 (N_83,In_514,In_631);
or U84 (N_84,In_592,In_734);
and U85 (N_85,In_149,In_657);
nand U86 (N_86,In_333,In_87);
and U87 (N_87,In_485,In_405);
or U88 (N_88,In_465,In_237);
or U89 (N_89,In_608,In_575);
nor U90 (N_90,In_165,In_372);
nand U91 (N_91,In_299,In_96);
and U92 (N_92,In_297,In_423);
nor U93 (N_93,In_727,In_406);
nand U94 (N_94,In_221,In_73);
nor U95 (N_95,In_293,In_401);
nand U96 (N_96,In_564,In_596);
nor U97 (N_97,In_693,In_190);
nor U98 (N_98,In_219,In_107);
nand U99 (N_99,In_522,In_680);
or U100 (N_100,In_90,In_748);
nand U101 (N_101,In_112,In_538);
nor U102 (N_102,In_463,In_143);
nand U103 (N_103,In_525,In_617);
nand U104 (N_104,In_180,In_546);
xor U105 (N_105,In_524,In_586);
nor U106 (N_106,In_273,In_63);
nor U107 (N_107,In_597,In_99);
nand U108 (N_108,In_683,In_193);
nand U109 (N_109,In_223,In_382);
and U110 (N_110,In_682,In_640);
or U111 (N_111,In_58,In_18);
nor U112 (N_112,In_157,In_705);
nor U113 (N_113,In_630,In_144);
nand U114 (N_114,In_481,In_578);
and U115 (N_115,In_81,In_147);
nand U116 (N_116,In_696,In_11);
nand U117 (N_117,In_681,In_484);
and U118 (N_118,In_340,In_345);
nor U119 (N_119,In_84,In_474);
nor U120 (N_120,In_199,In_21);
nand U121 (N_121,In_365,In_451);
nor U122 (N_122,In_8,In_673);
or U123 (N_123,In_267,In_217);
and U124 (N_124,In_403,In_398);
or U125 (N_125,In_348,In_249);
or U126 (N_126,In_749,In_119);
and U127 (N_127,In_394,In_473);
and U128 (N_128,In_200,In_305);
nand U129 (N_129,In_129,In_10);
nand U130 (N_130,In_448,In_601);
nor U131 (N_131,In_386,In_381);
or U132 (N_132,In_312,In_580);
or U133 (N_133,In_307,In_457);
nand U134 (N_134,In_408,In_66);
nand U135 (N_135,In_719,In_412);
nor U136 (N_136,In_527,In_253);
and U137 (N_137,In_303,In_202);
nand U138 (N_138,In_295,In_227);
nor U139 (N_139,In_483,In_629);
nor U140 (N_140,In_171,In_329);
or U141 (N_141,In_516,In_424);
or U142 (N_142,In_493,In_709);
or U143 (N_143,In_68,In_279);
or U144 (N_144,In_77,In_501);
and U145 (N_145,In_363,In_332);
or U146 (N_146,In_612,In_468);
or U147 (N_147,In_226,In_743);
or U148 (N_148,In_645,In_111);
or U149 (N_149,In_428,In_698);
nand U150 (N_150,In_395,In_264);
nand U151 (N_151,In_337,In_519);
or U152 (N_152,In_211,In_545);
nor U153 (N_153,In_557,In_196);
and U154 (N_154,In_50,In_235);
nor U155 (N_155,In_360,In_498);
nand U156 (N_156,In_738,In_469);
or U157 (N_157,In_676,In_515);
nor U158 (N_158,In_666,In_526);
nand U159 (N_159,In_206,In_594);
nand U160 (N_160,In_9,In_414);
nand U161 (N_161,In_446,In_690);
or U162 (N_162,In_38,In_602);
or U163 (N_163,In_477,In_688);
nor U164 (N_164,In_3,In_742);
or U165 (N_165,In_49,In_358);
nor U166 (N_166,In_32,In_150);
nor U167 (N_167,In_435,In_355);
nor U168 (N_168,In_170,In_1);
and U169 (N_169,In_169,In_628);
or U170 (N_170,In_562,In_254);
or U171 (N_171,In_511,In_731);
and U172 (N_172,In_678,In_240);
nor U173 (N_173,In_101,In_416);
nor U174 (N_174,In_439,In_257);
nand U175 (N_175,In_214,In_216);
and U176 (N_176,In_93,In_261);
and U177 (N_177,In_338,In_142);
or U178 (N_178,In_179,In_145);
and U179 (N_179,In_5,In_400);
nand U180 (N_180,In_542,In_725);
and U181 (N_181,In_376,In_521);
nor U182 (N_182,In_582,In_464);
nor U183 (N_183,In_97,In_52);
or U184 (N_184,In_242,In_686);
or U185 (N_185,In_53,In_646);
nor U186 (N_186,In_317,In_116);
or U187 (N_187,In_614,In_128);
nor U188 (N_188,In_373,In_417);
nor U189 (N_189,In_74,In_368);
nor U190 (N_190,In_353,In_737);
nor U191 (N_191,In_318,In_34);
and U192 (N_192,In_173,In_491);
nand U193 (N_193,In_662,In_118);
nand U194 (N_194,In_637,In_689);
and U195 (N_195,In_503,In_387);
or U196 (N_196,In_393,In_215);
or U197 (N_197,In_44,In_547);
nand U198 (N_198,In_310,In_561);
nor U199 (N_199,In_278,In_258);
and U200 (N_200,In_591,In_238);
or U201 (N_201,In_620,In_533);
or U202 (N_202,In_194,In_42);
nor U203 (N_203,In_20,In_711);
nand U204 (N_204,In_156,In_404);
and U205 (N_205,In_283,In_76);
nand U206 (N_206,In_182,In_225);
nand U207 (N_207,In_198,In_425);
nor U208 (N_208,In_83,In_470);
nand U209 (N_209,In_195,In_671);
and U210 (N_210,In_415,In_418);
or U211 (N_211,In_618,In_536);
nor U212 (N_212,In_649,In_51);
nand U213 (N_213,In_313,In_569);
nand U214 (N_214,In_286,In_595);
and U215 (N_215,In_482,In_706);
and U216 (N_216,In_409,In_486);
or U217 (N_217,In_397,In_656);
nand U218 (N_218,In_647,In_367);
nor U219 (N_219,In_452,In_304);
or U220 (N_220,In_664,In_25);
nor U221 (N_221,In_230,In_655);
or U222 (N_222,In_454,In_733);
or U223 (N_223,In_652,In_247);
or U224 (N_224,In_496,In_328);
and U225 (N_225,In_276,In_108);
nand U226 (N_226,In_507,In_632);
and U227 (N_227,In_721,In_535);
nand U228 (N_228,In_739,In_336);
or U229 (N_229,In_191,In_389);
nor U230 (N_230,In_152,In_325);
or U231 (N_231,In_6,In_28);
nor U232 (N_232,In_285,In_532);
or U233 (N_233,In_256,In_281);
nand U234 (N_234,In_205,In_550);
nand U235 (N_235,In_378,In_565);
or U236 (N_236,In_131,In_104);
nand U237 (N_237,In_183,In_716);
and U238 (N_238,In_540,In_492);
nor U239 (N_239,In_56,In_100);
or U240 (N_240,In_531,In_236);
or U241 (N_241,In_91,In_55);
xnor U242 (N_242,In_23,In_222);
nor U243 (N_243,In_500,In_105);
and U244 (N_244,In_567,In_121);
or U245 (N_245,In_178,In_566);
nor U246 (N_246,In_603,In_36);
nor U247 (N_247,In_723,In_396);
or U248 (N_248,In_65,In_33);
and U249 (N_249,In_440,In_164);
and U250 (N_250,In_132,In_60);
nor U251 (N_251,In_499,In_349);
and U252 (N_252,In_443,In_520);
or U253 (N_253,In_54,In_554);
xnor U254 (N_254,In_490,In_271);
nand U255 (N_255,In_675,In_302);
nor U256 (N_256,In_246,In_626);
or U257 (N_257,In_445,In_207);
or U258 (N_258,In_4,In_37);
nor U259 (N_259,In_447,In_487);
or U260 (N_260,In_239,In_48);
or U261 (N_261,In_552,In_461);
or U262 (N_262,In_86,In_383);
nand U263 (N_263,In_208,In_89);
or U264 (N_264,In_366,In_702);
nor U265 (N_265,In_518,In_123);
or U266 (N_266,In_627,In_421);
and U267 (N_267,In_604,In_233);
or U268 (N_268,In_75,In_139);
and U269 (N_269,In_718,In_275);
nand U270 (N_270,In_466,In_229);
or U271 (N_271,In_291,In_300);
and U272 (N_272,In_674,In_621);
nand U273 (N_273,In_159,In_695);
nor U274 (N_274,In_177,In_176);
and U275 (N_275,In_350,In_347);
nor U276 (N_276,In_708,In_600);
and U277 (N_277,In_622,In_699);
nor U278 (N_278,In_650,In_642);
or U279 (N_279,In_504,In_430);
or U280 (N_280,In_192,In_45);
and U281 (N_281,In_115,In_185);
nor U282 (N_282,In_342,In_311);
nor U283 (N_283,In_479,In_138);
or U284 (N_284,In_529,In_472);
and U285 (N_285,In_22,In_266);
nand U286 (N_286,In_361,In_419);
nor U287 (N_287,In_125,In_67);
and U288 (N_288,In_234,In_658);
or U289 (N_289,In_320,In_534);
and U290 (N_290,In_64,In_606);
and U291 (N_291,In_583,In_346);
nand U292 (N_292,In_687,In_459);
or U293 (N_293,In_356,In_669);
nor U294 (N_294,In_140,In_453);
or U295 (N_295,In_636,In_523);
or U296 (N_296,In_585,In_588);
nand U297 (N_297,In_380,In_265);
nand U298 (N_298,In_16,In_29);
and U299 (N_299,In_335,In_712);
nor U300 (N_300,In_654,In_57);
or U301 (N_301,In_537,In_19);
or U302 (N_302,In_0,In_344);
and U303 (N_303,In_181,In_130);
nor U304 (N_304,In_141,In_551);
nand U305 (N_305,In_506,In_334);
nor U306 (N_306,In_710,In_726);
nand U307 (N_307,In_85,In_667);
nor U308 (N_308,In_243,In_270);
and U309 (N_309,In_377,In_441);
nor U310 (N_310,In_610,In_127);
nand U311 (N_311,In_309,In_660);
nor U312 (N_312,In_747,In_274);
xor U313 (N_313,In_162,In_109);
and U314 (N_314,In_290,In_541);
nand U315 (N_315,In_122,In_268);
nand U316 (N_316,In_135,In_590);
nand U317 (N_317,In_364,In_707);
and U318 (N_318,In_599,In_745);
and U319 (N_319,In_379,In_94);
or U320 (N_320,In_634,In_544);
nor U321 (N_321,In_13,In_92);
nand U322 (N_322,In_213,In_260);
nand U323 (N_323,In_231,In_241);
and U324 (N_324,In_694,In_252);
nor U325 (N_325,In_572,In_120);
or U326 (N_326,In_126,In_272);
nor U327 (N_327,In_576,In_581);
and U328 (N_328,In_251,In_280);
nand U329 (N_329,In_437,In_584);
nor U330 (N_330,In_72,In_82);
nand U331 (N_331,In_607,In_308);
nand U332 (N_332,In_255,In_568);
or U333 (N_333,In_729,In_319);
nand U334 (N_334,In_61,In_704);
and U335 (N_335,In_17,In_301);
or U336 (N_336,In_110,In_433);
nand U337 (N_337,In_476,In_728);
nand U338 (N_338,In_232,In_220);
or U339 (N_339,In_14,In_354);
nor U340 (N_340,In_245,In_384);
or U341 (N_341,In_420,In_555);
nand U342 (N_342,In_450,In_434);
nand U343 (N_343,In_619,In_41);
nand U344 (N_344,In_263,In_146);
nand U345 (N_345,In_70,In_613);
nor U346 (N_346,In_322,In_357);
and U347 (N_347,In_697,In_167);
and U348 (N_348,In_343,In_136);
nor U349 (N_349,In_700,In_549);
nor U350 (N_350,In_7,In_668);
and U351 (N_351,In_548,In_508);
and U352 (N_352,In_593,In_559);
and U353 (N_353,In_392,In_714);
nand U354 (N_354,In_692,In_316);
nand U355 (N_355,In_444,In_174);
nand U356 (N_356,In_323,In_352);
or U357 (N_357,In_639,In_31);
nor U358 (N_358,In_35,In_713);
nand U359 (N_359,In_282,In_616);
nand U360 (N_360,In_47,In_623);
nand U361 (N_361,In_341,In_321);
nor U362 (N_362,In_186,In_43);
nand U363 (N_363,In_269,In_289);
and U364 (N_364,In_12,In_432);
or U365 (N_365,In_458,In_362);
nor U366 (N_366,In_201,In_732);
nand U367 (N_367,In_410,In_587);
and U368 (N_368,In_371,In_505);
nor U369 (N_369,In_720,In_250);
and U370 (N_370,In_717,In_114);
or U371 (N_371,In_624,In_399);
nor U372 (N_372,In_703,In_339);
or U373 (N_373,In_98,In_741);
or U374 (N_374,In_411,In_615);
and U375 (N_375,In_452,In_158);
and U376 (N_376,In_60,In_401);
nor U377 (N_377,In_117,In_699);
nor U378 (N_378,In_33,In_247);
and U379 (N_379,In_593,In_663);
nand U380 (N_380,In_409,In_354);
or U381 (N_381,In_194,In_412);
and U382 (N_382,In_565,In_369);
nand U383 (N_383,In_288,In_259);
and U384 (N_384,In_47,In_40);
nor U385 (N_385,In_689,In_45);
nand U386 (N_386,In_607,In_511);
or U387 (N_387,In_614,In_162);
nand U388 (N_388,In_221,In_467);
nor U389 (N_389,In_11,In_485);
nand U390 (N_390,In_183,In_311);
and U391 (N_391,In_215,In_704);
or U392 (N_392,In_285,In_172);
or U393 (N_393,In_84,In_107);
nand U394 (N_394,In_282,In_195);
and U395 (N_395,In_78,In_584);
nor U396 (N_396,In_86,In_203);
and U397 (N_397,In_336,In_15);
nor U398 (N_398,In_415,In_41);
or U399 (N_399,In_63,In_681);
and U400 (N_400,In_248,In_1);
and U401 (N_401,In_212,In_410);
and U402 (N_402,In_624,In_120);
nor U403 (N_403,In_740,In_113);
nand U404 (N_404,In_546,In_595);
nand U405 (N_405,In_86,In_51);
nand U406 (N_406,In_253,In_338);
and U407 (N_407,In_329,In_250);
nand U408 (N_408,In_9,In_234);
and U409 (N_409,In_50,In_669);
nand U410 (N_410,In_226,In_668);
nand U411 (N_411,In_612,In_311);
nand U412 (N_412,In_475,In_432);
nand U413 (N_413,In_681,In_585);
nand U414 (N_414,In_214,In_40);
nor U415 (N_415,In_166,In_365);
and U416 (N_416,In_491,In_54);
nor U417 (N_417,In_275,In_625);
nor U418 (N_418,In_470,In_743);
nor U419 (N_419,In_646,In_160);
nor U420 (N_420,In_633,In_46);
nand U421 (N_421,In_127,In_69);
or U422 (N_422,In_416,In_155);
xnor U423 (N_423,In_509,In_108);
nand U424 (N_424,In_538,In_421);
and U425 (N_425,In_441,In_548);
nand U426 (N_426,In_26,In_746);
nor U427 (N_427,In_652,In_556);
nand U428 (N_428,In_530,In_384);
and U429 (N_429,In_169,In_328);
and U430 (N_430,In_592,In_340);
nand U431 (N_431,In_205,In_111);
nor U432 (N_432,In_229,In_313);
and U433 (N_433,In_45,In_229);
and U434 (N_434,In_252,In_334);
nand U435 (N_435,In_198,In_719);
nand U436 (N_436,In_163,In_537);
nor U437 (N_437,In_281,In_296);
and U438 (N_438,In_103,In_391);
or U439 (N_439,In_302,In_0);
and U440 (N_440,In_319,In_407);
or U441 (N_441,In_677,In_521);
nor U442 (N_442,In_209,In_167);
and U443 (N_443,In_124,In_74);
and U444 (N_444,In_543,In_339);
and U445 (N_445,In_42,In_137);
nor U446 (N_446,In_429,In_479);
and U447 (N_447,In_57,In_327);
nand U448 (N_448,In_692,In_657);
nand U449 (N_449,In_96,In_158);
nor U450 (N_450,In_465,In_621);
or U451 (N_451,In_347,In_338);
and U452 (N_452,In_281,In_623);
nor U453 (N_453,In_579,In_519);
nand U454 (N_454,In_523,In_493);
nand U455 (N_455,In_52,In_469);
or U456 (N_456,In_622,In_162);
nand U457 (N_457,In_176,In_135);
and U458 (N_458,In_682,In_45);
and U459 (N_459,In_207,In_174);
nand U460 (N_460,In_692,In_440);
nor U461 (N_461,In_0,In_22);
nand U462 (N_462,In_184,In_523);
or U463 (N_463,In_645,In_196);
nor U464 (N_464,In_273,In_123);
or U465 (N_465,In_353,In_691);
or U466 (N_466,In_199,In_134);
nand U467 (N_467,In_500,In_157);
and U468 (N_468,In_179,In_173);
nor U469 (N_469,In_561,In_35);
nor U470 (N_470,In_495,In_319);
or U471 (N_471,In_518,In_280);
nand U472 (N_472,In_485,In_602);
and U473 (N_473,In_417,In_205);
nand U474 (N_474,In_71,In_66);
nor U475 (N_475,In_175,In_31);
nand U476 (N_476,In_205,In_303);
nand U477 (N_477,In_152,In_707);
nand U478 (N_478,In_738,In_624);
nor U479 (N_479,In_544,In_398);
and U480 (N_480,In_163,In_353);
nor U481 (N_481,In_487,In_270);
or U482 (N_482,In_505,In_652);
or U483 (N_483,In_577,In_138);
and U484 (N_484,In_600,In_688);
nand U485 (N_485,In_223,In_74);
nand U486 (N_486,In_547,In_272);
nor U487 (N_487,In_726,In_294);
or U488 (N_488,In_141,In_707);
nor U489 (N_489,In_244,In_131);
nand U490 (N_490,In_62,In_326);
nor U491 (N_491,In_485,In_279);
or U492 (N_492,In_28,In_81);
and U493 (N_493,In_200,In_408);
and U494 (N_494,In_376,In_561);
nor U495 (N_495,In_706,In_284);
or U496 (N_496,In_593,In_190);
nor U497 (N_497,In_213,In_67);
nor U498 (N_498,In_600,In_490);
and U499 (N_499,In_320,In_462);
nand U500 (N_500,N_298,N_432);
or U501 (N_501,N_466,N_157);
and U502 (N_502,N_373,N_45);
nand U503 (N_503,N_226,N_104);
or U504 (N_504,N_50,N_346);
or U505 (N_505,N_303,N_124);
nor U506 (N_506,N_138,N_391);
nor U507 (N_507,N_61,N_151);
and U508 (N_508,N_195,N_60);
or U509 (N_509,N_110,N_116);
nand U510 (N_510,N_160,N_268);
nor U511 (N_511,N_206,N_299);
nand U512 (N_512,N_410,N_21);
and U513 (N_513,N_123,N_261);
or U514 (N_514,N_263,N_483);
nor U515 (N_515,N_314,N_360);
nand U516 (N_516,N_407,N_477);
or U517 (N_517,N_357,N_193);
and U518 (N_518,N_215,N_15);
and U519 (N_519,N_435,N_280);
nor U520 (N_520,N_384,N_205);
nand U521 (N_521,N_78,N_338);
nor U522 (N_522,N_284,N_118);
or U523 (N_523,N_81,N_198);
nor U524 (N_524,N_452,N_153);
nand U525 (N_525,N_34,N_207);
xnor U526 (N_526,N_492,N_159);
and U527 (N_527,N_386,N_352);
nor U528 (N_528,N_25,N_6);
nand U529 (N_529,N_276,N_250);
nor U530 (N_530,N_120,N_409);
nand U531 (N_531,N_289,N_12);
nand U532 (N_532,N_281,N_128);
nand U533 (N_533,N_443,N_48);
nand U534 (N_534,N_259,N_163);
nor U535 (N_535,N_145,N_8);
nor U536 (N_536,N_457,N_442);
nor U537 (N_537,N_449,N_376);
or U538 (N_538,N_393,N_112);
and U539 (N_539,N_392,N_271);
nand U540 (N_540,N_94,N_101);
nor U541 (N_541,N_139,N_349);
nor U542 (N_542,N_476,N_368);
and U543 (N_543,N_91,N_295);
or U544 (N_544,N_83,N_180);
and U545 (N_545,N_72,N_258);
or U546 (N_546,N_149,N_265);
nor U547 (N_547,N_321,N_305);
nor U548 (N_548,N_92,N_458);
nor U549 (N_549,N_194,N_228);
nor U550 (N_550,N_76,N_47);
and U551 (N_551,N_366,N_146);
nor U552 (N_552,N_319,N_428);
and U553 (N_553,N_309,N_42);
or U554 (N_554,N_64,N_465);
nand U555 (N_555,N_396,N_292);
or U556 (N_556,N_86,N_115);
and U557 (N_557,N_296,N_154);
and U558 (N_558,N_54,N_494);
or U559 (N_559,N_109,N_63);
or U560 (N_560,N_414,N_80);
nor U561 (N_561,N_317,N_274);
nand U562 (N_562,N_254,N_301);
nor U563 (N_563,N_406,N_106);
and U564 (N_564,N_41,N_275);
nor U565 (N_565,N_369,N_129);
or U566 (N_566,N_345,N_155);
nor U567 (N_567,N_479,N_491);
and U568 (N_568,N_221,N_127);
nor U569 (N_569,N_310,N_378);
nand U570 (N_570,N_256,N_37);
and U571 (N_571,N_260,N_171);
or U572 (N_572,N_196,N_168);
nand U573 (N_573,N_453,N_436);
nand U574 (N_574,N_133,N_282);
or U575 (N_575,N_200,N_411);
nand U576 (N_576,N_499,N_242);
nand U577 (N_577,N_342,N_401);
and U578 (N_578,N_403,N_188);
or U579 (N_579,N_247,N_29);
nor U580 (N_580,N_445,N_438);
nand U581 (N_581,N_4,N_39);
or U582 (N_582,N_277,N_167);
nand U583 (N_583,N_337,N_400);
and U584 (N_584,N_474,N_460);
and U585 (N_585,N_144,N_380);
and U586 (N_586,N_174,N_119);
and U587 (N_587,N_20,N_387);
nand U588 (N_588,N_66,N_439);
and U589 (N_589,N_99,N_287);
or U590 (N_590,N_251,N_44);
and U591 (N_591,N_297,N_100);
or U592 (N_592,N_448,N_70);
nor U593 (N_593,N_257,N_130);
nand U594 (N_594,N_31,N_362);
nor U595 (N_595,N_137,N_239);
or U596 (N_596,N_84,N_344);
nor U597 (N_597,N_397,N_473);
and U598 (N_598,N_192,N_253);
or U599 (N_599,N_135,N_184);
and U600 (N_600,N_96,N_212);
xnor U601 (N_601,N_7,N_33);
and U602 (N_602,N_481,N_142);
nand U603 (N_603,N_389,N_385);
and U604 (N_604,N_286,N_244);
nand U605 (N_605,N_418,N_482);
nor U606 (N_606,N_102,N_147);
or U607 (N_607,N_354,N_90);
or U608 (N_608,N_480,N_293);
or U609 (N_609,N_404,N_381);
nand U610 (N_610,N_177,N_5);
and U611 (N_611,N_93,N_113);
nand U612 (N_612,N_107,N_374);
nand U613 (N_613,N_176,N_136);
nor U614 (N_614,N_422,N_343);
nand U615 (N_615,N_464,N_427);
nor U616 (N_616,N_300,N_375);
or U617 (N_617,N_189,N_248);
nor U618 (N_618,N_313,N_450);
nor U619 (N_619,N_495,N_35);
and U620 (N_620,N_351,N_235);
or U621 (N_621,N_187,N_324);
nand U622 (N_622,N_365,N_150);
and U623 (N_623,N_463,N_53);
nor U624 (N_624,N_55,N_49);
or U625 (N_625,N_164,N_227);
xor U626 (N_626,N_423,N_370);
nand U627 (N_627,N_67,N_417);
nand U628 (N_628,N_493,N_203);
or U629 (N_629,N_348,N_197);
nand U630 (N_630,N_68,N_267);
nor U631 (N_631,N_191,N_325);
nand U632 (N_632,N_290,N_405);
and U633 (N_633,N_336,N_62);
or U634 (N_634,N_108,N_341);
and U635 (N_635,N_350,N_470);
and U636 (N_636,N_304,N_97);
and U637 (N_637,N_475,N_223);
nand U638 (N_638,N_140,N_339);
or U639 (N_639,N_111,N_364);
and U640 (N_640,N_199,N_307);
xor U641 (N_641,N_413,N_173);
nand U642 (N_642,N_59,N_455);
and U643 (N_643,N_231,N_272);
nor U644 (N_644,N_285,N_326);
nand U645 (N_645,N_132,N_18);
and U646 (N_646,N_148,N_323);
or U647 (N_647,N_426,N_51);
or U648 (N_648,N_121,N_316);
nor U649 (N_649,N_43,N_182);
and U650 (N_650,N_262,N_161);
and U651 (N_651,N_415,N_371);
nor U652 (N_652,N_447,N_273);
and U653 (N_653,N_213,N_1);
nand U654 (N_654,N_388,N_234);
nand U655 (N_655,N_255,N_82);
or U656 (N_656,N_216,N_98);
or U657 (N_657,N_114,N_421);
nor U658 (N_658,N_269,N_11);
or U659 (N_659,N_429,N_266);
or U660 (N_660,N_478,N_141);
or U661 (N_661,N_122,N_252);
or U662 (N_662,N_56,N_14);
and U663 (N_663,N_165,N_169);
nand U664 (N_664,N_420,N_416);
nand U665 (N_665,N_243,N_288);
nor U666 (N_666,N_158,N_65);
nor U667 (N_667,N_87,N_451);
nand U668 (N_668,N_322,N_156);
or U669 (N_669,N_125,N_430);
nand U670 (N_670,N_240,N_249);
nor U671 (N_671,N_408,N_166);
or U672 (N_672,N_390,N_85);
or U673 (N_673,N_238,N_209);
and U674 (N_674,N_472,N_383);
or U675 (N_675,N_245,N_334);
or U676 (N_676,N_16,N_327);
nand U677 (N_677,N_105,N_224);
nand U678 (N_678,N_237,N_73);
nor U679 (N_679,N_27,N_469);
or U680 (N_680,N_335,N_181);
nand U681 (N_681,N_441,N_359);
nand U682 (N_682,N_355,N_40);
or U683 (N_683,N_74,N_311);
nor U684 (N_684,N_270,N_279);
nor U685 (N_685,N_236,N_211);
nor U686 (N_686,N_318,N_17);
nand U687 (N_687,N_79,N_498);
nand U688 (N_688,N_103,N_331);
and U689 (N_689,N_328,N_382);
nor U690 (N_690,N_496,N_283);
nand U691 (N_691,N_294,N_13);
nor U692 (N_692,N_208,N_497);
or U693 (N_693,N_399,N_402);
or U694 (N_694,N_329,N_201);
or U695 (N_695,N_214,N_379);
and U696 (N_696,N_229,N_134);
nor U697 (N_697,N_488,N_3);
nand U698 (N_698,N_89,N_117);
or U699 (N_699,N_419,N_486);
nor U700 (N_700,N_433,N_372);
or U701 (N_701,N_461,N_179);
nand U702 (N_702,N_425,N_95);
or U703 (N_703,N_356,N_71);
and U704 (N_704,N_490,N_330);
nor U705 (N_705,N_77,N_126);
or U706 (N_706,N_456,N_52);
nor U707 (N_707,N_444,N_431);
nor U708 (N_708,N_22,N_315);
or U709 (N_709,N_398,N_485);
and U710 (N_710,N_202,N_19);
or U711 (N_711,N_222,N_36);
and U712 (N_712,N_264,N_424);
nand U713 (N_713,N_308,N_26);
and U714 (N_714,N_172,N_183);
nor U715 (N_715,N_0,N_467);
nor U716 (N_716,N_437,N_24);
and U717 (N_717,N_306,N_302);
and U718 (N_718,N_204,N_175);
or U719 (N_719,N_232,N_162);
nand U720 (N_720,N_312,N_218);
nand U721 (N_721,N_361,N_178);
and U722 (N_722,N_434,N_487);
or U723 (N_723,N_394,N_233);
nor U724 (N_724,N_332,N_333);
and U725 (N_725,N_210,N_454);
or U726 (N_726,N_57,N_412);
or U727 (N_727,N_69,N_9);
or U728 (N_728,N_489,N_75);
or U729 (N_729,N_10,N_358);
nand U730 (N_730,N_462,N_440);
nor U731 (N_731,N_186,N_471);
or U732 (N_732,N_246,N_468);
or U733 (N_733,N_38,N_32);
xnor U734 (N_734,N_353,N_446);
xnor U735 (N_735,N_152,N_230);
or U736 (N_736,N_278,N_28);
nand U737 (N_737,N_131,N_363);
and U738 (N_738,N_367,N_88);
and U739 (N_739,N_185,N_377);
and U740 (N_740,N_241,N_347);
or U741 (N_741,N_46,N_2);
or U742 (N_742,N_30,N_225);
or U743 (N_743,N_395,N_459);
and U744 (N_744,N_217,N_340);
or U745 (N_745,N_291,N_220);
nand U746 (N_746,N_320,N_190);
or U747 (N_747,N_143,N_219);
or U748 (N_748,N_58,N_170);
or U749 (N_749,N_484,N_23);
or U750 (N_750,N_296,N_379);
or U751 (N_751,N_390,N_402);
or U752 (N_752,N_350,N_498);
or U753 (N_753,N_26,N_42);
or U754 (N_754,N_347,N_322);
and U755 (N_755,N_71,N_443);
and U756 (N_756,N_141,N_196);
or U757 (N_757,N_336,N_125);
and U758 (N_758,N_283,N_121);
nand U759 (N_759,N_192,N_423);
nand U760 (N_760,N_338,N_439);
nand U761 (N_761,N_463,N_394);
and U762 (N_762,N_401,N_442);
or U763 (N_763,N_9,N_110);
or U764 (N_764,N_374,N_420);
nand U765 (N_765,N_8,N_282);
nand U766 (N_766,N_186,N_434);
nor U767 (N_767,N_11,N_128);
nor U768 (N_768,N_136,N_359);
and U769 (N_769,N_177,N_224);
nor U770 (N_770,N_105,N_334);
or U771 (N_771,N_216,N_63);
nor U772 (N_772,N_327,N_155);
nand U773 (N_773,N_350,N_495);
nand U774 (N_774,N_460,N_171);
or U775 (N_775,N_323,N_277);
and U776 (N_776,N_159,N_364);
and U777 (N_777,N_60,N_101);
nand U778 (N_778,N_33,N_422);
or U779 (N_779,N_210,N_29);
nor U780 (N_780,N_174,N_382);
nor U781 (N_781,N_169,N_6);
nand U782 (N_782,N_85,N_361);
and U783 (N_783,N_196,N_251);
nor U784 (N_784,N_233,N_101);
or U785 (N_785,N_91,N_40);
xnor U786 (N_786,N_101,N_152);
and U787 (N_787,N_356,N_240);
nor U788 (N_788,N_408,N_356);
nor U789 (N_789,N_99,N_375);
nand U790 (N_790,N_374,N_33);
or U791 (N_791,N_390,N_73);
and U792 (N_792,N_20,N_248);
and U793 (N_793,N_394,N_41);
and U794 (N_794,N_89,N_58);
nand U795 (N_795,N_495,N_164);
or U796 (N_796,N_54,N_388);
and U797 (N_797,N_303,N_129);
nand U798 (N_798,N_272,N_200);
or U799 (N_799,N_348,N_388);
or U800 (N_800,N_148,N_366);
nor U801 (N_801,N_417,N_410);
nand U802 (N_802,N_291,N_247);
and U803 (N_803,N_174,N_231);
or U804 (N_804,N_298,N_73);
nor U805 (N_805,N_428,N_480);
nand U806 (N_806,N_90,N_352);
nor U807 (N_807,N_420,N_18);
or U808 (N_808,N_274,N_112);
or U809 (N_809,N_106,N_330);
and U810 (N_810,N_308,N_326);
and U811 (N_811,N_12,N_227);
and U812 (N_812,N_334,N_192);
or U813 (N_813,N_432,N_451);
nor U814 (N_814,N_193,N_130);
nor U815 (N_815,N_170,N_98);
or U816 (N_816,N_467,N_432);
and U817 (N_817,N_12,N_15);
or U818 (N_818,N_3,N_404);
and U819 (N_819,N_254,N_53);
nor U820 (N_820,N_39,N_355);
nand U821 (N_821,N_335,N_260);
xor U822 (N_822,N_100,N_391);
or U823 (N_823,N_410,N_68);
or U824 (N_824,N_207,N_312);
nor U825 (N_825,N_355,N_114);
or U826 (N_826,N_426,N_148);
and U827 (N_827,N_226,N_166);
nor U828 (N_828,N_361,N_406);
nand U829 (N_829,N_496,N_179);
nor U830 (N_830,N_305,N_370);
and U831 (N_831,N_490,N_401);
nand U832 (N_832,N_258,N_140);
nor U833 (N_833,N_226,N_216);
and U834 (N_834,N_302,N_288);
or U835 (N_835,N_210,N_346);
or U836 (N_836,N_94,N_275);
nor U837 (N_837,N_312,N_28);
nor U838 (N_838,N_55,N_74);
and U839 (N_839,N_42,N_388);
nand U840 (N_840,N_76,N_105);
nand U841 (N_841,N_297,N_22);
nor U842 (N_842,N_65,N_59);
nor U843 (N_843,N_318,N_56);
and U844 (N_844,N_264,N_495);
nor U845 (N_845,N_15,N_124);
nand U846 (N_846,N_367,N_148);
nor U847 (N_847,N_231,N_499);
nor U848 (N_848,N_240,N_101);
nor U849 (N_849,N_192,N_453);
nand U850 (N_850,N_196,N_307);
or U851 (N_851,N_435,N_244);
nor U852 (N_852,N_268,N_27);
or U853 (N_853,N_311,N_90);
and U854 (N_854,N_466,N_24);
nor U855 (N_855,N_88,N_122);
nor U856 (N_856,N_299,N_3);
and U857 (N_857,N_403,N_87);
nand U858 (N_858,N_420,N_152);
nand U859 (N_859,N_105,N_399);
nand U860 (N_860,N_488,N_44);
nand U861 (N_861,N_0,N_114);
nor U862 (N_862,N_370,N_281);
nor U863 (N_863,N_291,N_184);
or U864 (N_864,N_33,N_322);
and U865 (N_865,N_386,N_50);
nor U866 (N_866,N_495,N_497);
nand U867 (N_867,N_158,N_300);
nor U868 (N_868,N_454,N_158);
nor U869 (N_869,N_444,N_384);
nand U870 (N_870,N_318,N_120);
and U871 (N_871,N_59,N_69);
and U872 (N_872,N_181,N_111);
and U873 (N_873,N_194,N_132);
and U874 (N_874,N_244,N_197);
nor U875 (N_875,N_410,N_142);
and U876 (N_876,N_382,N_262);
or U877 (N_877,N_55,N_352);
nor U878 (N_878,N_45,N_214);
and U879 (N_879,N_286,N_285);
nand U880 (N_880,N_163,N_47);
or U881 (N_881,N_266,N_417);
or U882 (N_882,N_234,N_233);
and U883 (N_883,N_302,N_459);
nand U884 (N_884,N_90,N_332);
nor U885 (N_885,N_47,N_321);
nor U886 (N_886,N_254,N_131);
and U887 (N_887,N_223,N_182);
nand U888 (N_888,N_10,N_284);
nor U889 (N_889,N_476,N_263);
nand U890 (N_890,N_165,N_467);
or U891 (N_891,N_169,N_140);
and U892 (N_892,N_215,N_166);
nor U893 (N_893,N_138,N_211);
nor U894 (N_894,N_3,N_464);
nor U895 (N_895,N_147,N_37);
nor U896 (N_896,N_397,N_102);
and U897 (N_897,N_197,N_81);
nor U898 (N_898,N_128,N_10);
and U899 (N_899,N_69,N_161);
nor U900 (N_900,N_263,N_55);
nor U901 (N_901,N_398,N_237);
and U902 (N_902,N_262,N_220);
and U903 (N_903,N_63,N_238);
nor U904 (N_904,N_130,N_414);
or U905 (N_905,N_439,N_21);
and U906 (N_906,N_293,N_405);
or U907 (N_907,N_85,N_412);
and U908 (N_908,N_119,N_19);
nand U909 (N_909,N_356,N_57);
nor U910 (N_910,N_57,N_295);
nor U911 (N_911,N_32,N_120);
and U912 (N_912,N_188,N_127);
or U913 (N_913,N_330,N_307);
or U914 (N_914,N_193,N_137);
and U915 (N_915,N_60,N_447);
nor U916 (N_916,N_151,N_86);
and U917 (N_917,N_52,N_279);
and U918 (N_918,N_286,N_75);
or U919 (N_919,N_90,N_249);
and U920 (N_920,N_418,N_456);
and U921 (N_921,N_162,N_0);
or U922 (N_922,N_423,N_39);
nor U923 (N_923,N_353,N_155);
and U924 (N_924,N_381,N_59);
and U925 (N_925,N_74,N_489);
and U926 (N_926,N_397,N_390);
nand U927 (N_927,N_304,N_359);
or U928 (N_928,N_228,N_358);
or U929 (N_929,N_414,N_92);
and U930 (N_930,N_188,N_175);
nand U931 (N_931,N_59,N_309);
or U932 (N_932,N_390,N_359);
nand U933 (N_933,N_328,N_454);
and U934 (N_934,N_372,N_90);
and U935 (N_935,N_320,N_14);
xor U936 (N_936,N_134,N_491);
or U937 (N_937,N_413,N_47);
and U938 (N_938,N_177,N_381);
nor U939 (N_939,N_36,N_488);
or U940 (N_940,N_236,N_451);
or U941 (N_941,N_351,N_468);
nor U942 (N_942,N_290,N_189);
nand U943 (N_943,N_301,N_54);
or U944 (N_944,N_133,N_121);
nor U945 (N_945,N_484,N_384);
nand U946 (N_946,N_456,N_450);
and U947 (N_947,N_154,N_388);
nor U948 (N_948,N_496,N_123);
nor U949 (N_949,N_478,N_102);
or U950 (N_950,N_441,N_137);
and U951 (N_951,N_45,N_249);
nand U952 (N_952,N_356,N_182);
or U953 (N_953,N_385,N_349);
xor U954 (N_954,N_259,N_235);
nand U955 (N_955,N_51,N_307);
and U956 (N_956,N_426,N_490);
or U957 (N_957,N_13,N_417);
or U958 (N_958,N_335,N_436);
nor U959 (N_959,N_226,N_136);
nand U960 (N_960,N_216,N_451);
xnor U961 (N_961,N_380,N_32);
and U962 (N_962,N_402,N_108);
nor U963 (N_963,N_391,N_74);
nor U964 (N_964,N_25,N_32);
or U965 (N_965,N_65,N_146);
nor U966 (N_966,N_355,N_489);
or U967 (N_967,N_227,N_13);
nand U968 (N_968,N_465,N_347);
nand U969 (N_969,N_17,N_175);
nand U970 (N_970,N_385,N_246);
and U971 (N_971,N_401,N_479);
nor U972 (N_972,N_402,N_453);
nand U973 (N_973,N_105,N_323);
nor U974 (N_974,N_413,N_299);
nand U975 (N_975,N_485,N_317);
or U976 (N_976,N_417,N_68);
nand U977 (N_977,N_472,N_491);
nand U978 (N_978,N_198,N_103);
nand U979 (N_979,N_363,N_347);
or U980 (N_980,N_113,N_251);
or U981 (N_981,N_144,N_242);
nor U982 (N_982,N_11,N_423);
nand U983 (N_983,N_102,N_110);
nor U984 (N_984,N_438,N_230);
nand U985 (N_985,N_104,N_361);
nand U986 (N_986,N_250,N_323);
or U987 (N_987,N_471,N_74);
or U988 (N_988,N_492,N_229);
or U989 (N_989,N_157,N_322);
nor U990 (N_990,N_169,N_282);
and U991 (N_991,N_321,N_110);
nand U992 (N_992,N_244,N_209);
nor U993 (N_993,N_394,N_12);
nand U994 (N_994,N_335,N_306);
nor U995 (N_995,N_141,N_431);
and U996 (N_996,N_303,N_76);
nand U997 (N_997,N_14,N_234);
nor U998 (N_998,N_198,N_445);
and U999 (N_999,N_411,N_205);
nor U1000 (N_1000,N_971,N_925);
nor U1001 (N_1001,N_822,N_812);
nand U1002 (N_1002,N_569,N_869);
nand U1003 (N_1003,N_969,N_556);
xnor U1004 (N_1004,N_661,N_967);
and U1005 (N_1005,N_761,N_974);
nand U1006 (N_1006,N_549,N_851);
or U1007 (N_1007,N_573,N_729);
nor U1008 (N_1008,N_558,N_766);
nand U1009 (N_1009,N_989,N_616);
or U1010 (N_1010,N_696,N_805);
or U1011 (N_1011,N_957,N_914);
nand U1012 (N_1012,N_928,N_600);
and U1013 (N_1013,N_744,N_735);
and U1014 (N_1014,N_560,N_620);
nor U1015 (N_1015,N_929,N_849);
and U1016 (N_1016,N_688,N_977);
xnor U1017 (N_1017,N_954,N_791);
or U1018 (N_1018,N_917,N_644);
nor U1019 (N_1019,N_763,N_997);
nor U1020 (N_1020,N_764,N_937);
nor U1021 (N_1021,N_955,N_528);
nand U1022 (N_1022,N_539,N_519);
nand U1023 (N_1023,N_594,N_523);
nand U1024 (N_1024,N_613,N_831);
nand U1025 (N_1025,N_837,N_704);
or U1026 (N_1026,N_727,N_730);
and U1027 (N_1027,N_570,N_793);
and U1028 (N_1028,N_529,N_920);
and U1029 (N_1029,N_625,N_733);
nor U1030 (N_1030,N_976,N_842);
and U1031 (N_1031,N_577,N_888);
and U1032 (N_1032,N_916,N_605);
and U1033 (N_1033,N_634,N_682);
nand U1034 (N_1034,N_774,N_742);
nand U1035 (N_1035,N_778,N_972);
and U1036 (N_1036,N_843,N_904);
and U1037 (N_1037,N_609,N_502);
nor U1038 (N_1038,N_617,N_859);
and U1039 (N_1039,N_676,N_825);
nor U1040 (N_1040,N_965,N_959);
nand U1041 (N_1041,N_692,N_941);
nand U1042 (N_1042,N_695,N_855);
nand U1043 (N_1043,N_503,N_884);
or U1044 (N_1044,N_902,N_897);
nor U1045 (N_1045,N_611,N_581);
or U1046 (N_1046,N_792,N_547);
and U1047 (N_1047,N_653,N_794);
or U1048 (N_1048,N_621,N_555);
and U1049 (N_1049,N_991,N_602);
nor U1050 (N_1050,N_639,N_557);
nor U1051 (N_1051,N_681,N_599);
and U1052 (N_1052,N_685,N_747);
and U1053 (N_1053,N_619,N_840);
nor U1054 (N_1054,N_996,N_584);
and U1055 (N_1055,N_736,N_618);
nand U1056 (N_1056,N_782,N_811);
nor U1057 (N_1057,N_820,N_576);
nor U1058 (N_1058,N_873,N_567);
and U1059 (N_1059,N_891,N_731);
nand U1060 (N_1060,N_658,N_823);
nor U1061 (N_1061,N_648,N_777);
and U1062 (N_1062,N_881,N_901);
nand U1063 (N_1063,N_948,N_745);
nand U1064 (N_1064,N_604,N_583);
and U1065 (N_1065,N_728,N_850);
nor U1066 (N_1066,N_958,N_741);
nor U1067 (N_1067,N_910,N_776);
nand U1068 (N_1068,N_527,N_511);
and U1069 (N_1069,N_746,N_799);
nor U1070 (N_1070,N_828,N_757);
and U1071 (N_1071,N_980,N_815);
or U1072 (N_1072,N_537,N_554);
nor U1073 (N_1073,N_934,N_927);
or U1074 (N_1074,N_988,N_614);
or U1075 (N_1075,N_877,N_943);
nand U1076 (N_1076,N_845,N_572);
nor U1077 (N_1077,N_932,N_838);
and U1078 (N_1078,N_771,N_802);
or U1079 (N_1079,N_908,N_933);
and U1080 (N_1080,N_804,N_713);
and U1081 (N_1081,N_912,N_669);
and U1082 (N_1082,N_952,N_524);
nand U1083 (N_1083,N_889,N_720);
and U1084 (N_1084,N_754,N_919);
and U1085 (N_1085,N_907,N_854);
and U1086 (N_1086,N_945,N_737);
nor U1087 (N_1087,N_672,N_807);
and U1088 (N_1088,N_551,N_751);
or U1089 (N_1089,N_610,N_668);
or U1090 (N_1090,N_832,N_652);
nor U1091 (N_1091,N_906,N_562);
and U1092 (N_1092,N_939,N_810);
nand U1093 (N_1093,N_702,N_998);
and U1094 (N_1094,N_630,N_699);
and U1095 (N_1095,N_515,N_824);
nor U1096 (N_1096,N_638,N_657);
nand U1097 (N_1097,N_856,N_615);
nor U1098 (N_1098,N_979,N_505);
or U1099 (N_1099,N_871,N_646);
and U1100 (N_1100,N_755,N_975);
and U1101 (N_1101,N_973,N_950);
nor U1102 (N_1102,N_852,N_809);
nor U1103 (N_1103,N_595,N_698);
nor U1104 (N_1104,N_743,N_675);
or U1105 (N_1105,N_775,N_946);
and U1106 (N_1106,N_585,N_773);
nand U1107 (N_1107,N_844,N_705);
nor U1108 (N_1108,N_506,N_772);
and U1109 (N_1109,N_701,N_748);
and U1110 (N_1110,N_936,N_833);
or U1111 (N_1111,N_964,N_947);
or U1112 (N_1112,N_753,N_689);
nor U1113 (N_1113,N_968,N_836);
nand U1114 (N_1114,N_752,N_848);
nand U1115 (N_1115,N_953,N_714);
and U1116 (N_1116,N_880,N_995);
or U1117 (N_1117,N_885,N_983);
and U1118 (N_1118,N_538,N_990);
or U1119 (N_1119,N_545,N_926);
nor U1120 (N_1120,N_588,N_740);
nand U1121 (N_1121,N_949,N_924);
nor U1122 (N_1122,N_978,N_870);
or U1123 (N_1123,N_544,N_798);
nor U1124 (N_1124,N_711,N_700);
nor U1125 (N_1125,N_826,N_874);
nor U1126 (N_1126,N_655,N_865);
nand U1127 (N_1127,N_803,N_708);
nand U1128 (N_1128,N_520,N_944);
nor U1129 (N_1129,N_568,N_629);
nor U1130 (N_1130,N_863,N_670);
and U1131 (N_1131,N_517,N_500);
and U1132 (N_1132,N_637,N_717);
nand U1133 (N_1133,N_666,N_656);
or U1134 (N_1134,N_636,N_531);
nor U1135 (N_1135,N_886,N_516);
and U1136 (N_1136,N_834,N_624);
nor U1137 (N_1137,N_598,N_726);
and U1138 (N_1138,N_808,N_786);
or U1139 (N_1139,N_862,N_680);
nand U1140 (N_1140,N_841,N_892);
nor U1141 (N_1141,N_795,N_574);
nand U1142 (N_1142,N_853,N_898);
nand U1143 (N_1143,N_739,N_984);
and U1144 (N_1144,N_543,N_864);
nor U1145 (N_1145,N_663,N_521);
nand U1146 (N_1146,N_903,N_597);
nor U1147 (N_1147,N_921,N_918);
nand U1148 (N_1148,N_501,N_632);
nand U1149 (N_1149,N_900,N_876);
or U1150 (N_1150,N_905,N_533);
and U1151 (N_1151,N_575,N_963);
nor U1152 (N_1152,N_565,N_915);
nor U1153 (N_1153,N_719,N_878);
nand U1154 (N_1154,N_942,N_541);
or U1155 (N_1155,N_857,N_797);
nor U1156 (N_1156,N_966,N_821);
or U1157 (N_1157,N_718,N_767);
nor U1158 (N_1158,N_591,N_830);
nand U1159 (N_1159,N_665,N_899);
nor U1160 (N_1160,N_522,N_703);
nor U1161 (N_1161,N_961,N_694);
nand U1162 (N_1162,N_813,N_985);
nand U1163 (N_1163,N_587,N_866);
and U1164 (N_1164,N_534,N_530);
and U1165 (N_1165,N_765,N_819);
and U1166 (N_1166,N_686,N_654);
nand U1167 (N_1167,N_986,N_643);
xor U1168 (N_1168,N_867,N_930);
and U1169 (N_1169,N_548,N_607);
nand U1170 (N_1170,N_879,N_514);
nor U1171 (N_1171,N_715,N_509);
nor U1172 (N_1172,N_860,N_635);
nor U1173 (N_1173,N_586,N_525);
nor U1174 (N_1174,N_536,N_893);
and U1175 (N_1175,N_691,N_542);
nor U1176 (N_1176,N_938,N_716);
nor U1177 (N_1177,N_706,N_962);
or U1178 (N_1178,N_895,N_999);
nor U1179 (N_1179,N_667,N_896);
nand U1180 (N_1180,N_783,N_582);
nor U1181 (N_1181,N_508,N_817);
and U1182 (N_1182,N_970,N_801);
nor U1183 (N_1183,N_606,N_951);
nor U1184 (N_1184,N_738,N_861);
nand U1185 (N_1185,N_993,N_762);
and U1186 (N_1186,N_535,N_553);
and U1187 (N_1187,N_806,N_758);
nand U1188 (N_1188,N_723,N_697);
nand U1189 (N_1189,N_872,N_818);
and U1190 (N_1190,N_931,N_829);
and U1191 (N_1191,N_725,N_790);
or U1192 (N_1192,N_566,N_677);
nor U1193 (N_1193,N_679,N_796);
or U1194 (N_1194,N_913,N_875);
and U1195 (N_1195,N_507,N_526);
or U1196 (N_1196,N_512,N_552);
and U1197 (N_1197,N_759,N_724);
and U1198 (N_1198,N_592,N_601);
and U1199 (N_1199,N_827,N_603);
and U1200 (N_1200,N_664,N_923);
xnor U1201 (N_1201,N_642,N_956);
or U1202 (N_1202,N_981,N_780);
nor U1203 (N_1203,N_847,N_684);
and U1204 (N_1204,N_641,N_589);
and U1205 (N_1205,N_504,N_707);
and U1206 (N_1206,N_712,N_649);
and U1207 (N_1207,N_540,N_868);
nand U1208 (N_1208,N_960,N_633);
and U1209 (N_1209,N_647,N_890);
nor U1210 (N_1210,N_561,N_883);
and U1211 (N_1211,N_580,N_563);
or U1212 (N_1212,N_922,N_769);
nand U1213 (N_1213,N_674,N_690);
or U1214 (N_1214,N_631,N_640);
nor U1215 (N_1215,N_816,N_660);
and U1216 (N_1216,N_887,N_628);
nand U1217 (N_1217,N_546,N_596);
nor U1218 (N_1218,N_846,N_659);
xnor U1219 (N_1219,N_785,N_709);
nand U1220 (N_1220,N_882,N_909);
nor U1221 (N_1221,N_651,N_518);
nand U1222 (N_1222,N_940,N_781);
or U1223 (N_1223,N_662,N_590);
and U1224 (N_1224,N_578,N_749);
nor U1225 (N_1225,N_510,N_835);
nor U1226 (N_1226,N_650,N_722);
or U1227 (N_1227,N_788,N_559);
nand U1228 (N_1228,N_721,N_992);
or U1229 (N_1229,N_678,N_612);
or U1230 (N_1230,N_693,N_645);
nor U1231 (N_1231,N_894,N_710);
or U1232 (N_1232,N_687,N_814);
nor U1233 (N_1233,N_779,N_787);
and U1234 (N_1234,N_671,N_839);
nor U1235 (N_1235,N_513,N_784);
nand U1236 (N_1236,N_550,N_626);
or U1237 (N_1237,N_579,N_732);
nand U1238 (N_1238,N_760,N_770);
and U1239 (N_1239,N_532,N_683);
nor U1240 (N_1240,N_564,N_750);
nor U1241 (N_1241,N_768,N_982);
and U1242 (N_1242,N_673,N_734);
nor U1243 (N_1243,N_935,N_994);
and U1244 (N_1244,N_756,N_800);
and U1245 (N_1245,N_593,N_608);
nor U1246 (N_1246,N_571,N_622);
or U1247 (N_1247,N_789,N_911);
or U1248 (N_1248,N_627,N_623);
nand U1249 (N_1249,N_858,N_987);
nand U1250 (N_1250,N_956,N_775);
nand U1251 (N_1251,N_511,N_552);
and U1252 (N_1252,N_585,N_750);
nor U1253 (N_1253,N_849,N_517);
nand U1254 (N_1254,N_750,N_921);
or U1255 (N_1255,N_901,N_821);
nor U1256 (N_1256,N_840,N_788);
xnor U1257 (N_1257,N_990,N_666);
and U1258 (N_1258,N_890,N_790);
and U1259 (N_1259,N_995,N_623);
nand U1260 (N_1260,N_811,N_871);
or U1261 (N_1261,N_693,N_809);
nand U1262 (N_1262,N_806,N_797);
nand U1263 (N_1263,N_916,N_889);
and U1264 (N_1264,N_727,N_863);
and U1265 (N_1265,N_838,N_752);
nor U1266 (N_1266,N_954,N_988);
and U1267 (N_1267,N_821,N_610);
or U1268 (N_1268,N_607,N_843);
nor U1269 (N_1269,N_663,N_849);
nand U1270 (N_1270,N_838,N_949);
and U1271 (N_1271,N_830,N_561);
nand U1272 (N_1272,N_873,N_886);
or U1273 (N_1273,N_596,N_531);
and U1274 (N_1274,N_587,N_697);
nand U1275 (N_1275,N_986,N_593);
nor U1276 (N_1276,N_705,N_500);
and U1277 (N_1277,N_779,N_903);
or U1278 (N_1278,N_884,N_804);
or U1279 (N_1279,N_944,N_905);
and U1280 (N_1280,N_913,N_818);
or U1281 (N_1281,N_707,N_703);
and U1282 (N_1282,N_669,N_854);
and U1283 (N_1283,N_616,N_599);
nand U1284 (N_1284,N_779,N_877);
and U1285 (N_1285,N_600,N_818);
nand U1286 (N_1286,N_807,N_787);
and U1287 (N_1287,N_615,N_764);
nand U1288 (N_1288,N_639,N_535);
nor U1289 (N_1289,N_822,N_756);
and U1290 (N_1290,N_967,N_766);
xor U1291 (N_1291,N_985,N_910);
nor U1292 (N_1292,N_738,N_668);
nor U1293 (N_1293,N_802,N_821);
or U1294 (N_1294,N_561,N_920);
nand U1295 (N_1295,N_720,N_780);
nand U1296 (N_1296,N_654,N_746);
nor U1297 (N_1297,N_507,N_912);
nor U1298 (N_1298,N_560,N_603);
and U1299 (N_1299,N_746,N_844);
nand U1300 (N_1300,N_889,N_896);
or U1301 (N_1301,N_578,N_558);
nand U1302 (N_1302,N_601,N_895);
and U1303 (N_1303,N_567,N_854);
or U1304 (N_1304,N_521,N_974);
or U1305 (N_1305,N_914,N_999);
nor U1306 (N_1306,N_502,N_887);
nand U1307 (N_1307,N_921,N_599);
or U1308 (N_1308,N_669,N_881);
or U1309 (N_1309,N_858,N_915);
or U1310 (N_1310,N_661,N_525);
nor U1311 (N_1311,N_566,N_731);
nor U1312 (N_1312,N_642,N_801);
nor U1313 (N_1313,N_820,N_727);
nor U1314 (N_1314,N_598,N_789);
or U1315 (N_1315,N_551,N_565);
nor U1316 (N_1316,N_524,N_836);
or U1317 (N_1317,N_797,N_755);
nor U1318 (N_1318,N_780,N_599);
nand U1319 (N_1319,N_859,N_637);
nand U1320 (N_1320,N_964,N_539);
nand U1321 (N_1321,N_861,N_626);
or U1322 (N_1322,N_694,N_887);
nor U1323 (N_1323,N_537,N_925);
and U1324 (N_1324,N_841,N_838);
and U1325 (N_1325,N_832,N_918);
nand U1326 (N_1326,N_563,N_927);
nor U1327 (N_1327,N_518,N_645);
and U1328 (N_1328,N_786,N_989);
nor U1329 (N_1329,N_539,N_861);
nor U1330 (N_1330,N_959,N_512);
and U1331 (N_1331,N_968,N_647);
nor U1332 (N_1332,N_873,N_993);
and U1333 (N_1333,N_840,N_870);
or U1334 (N_1334,N_785,N_988);
and U1335 (N_1335,N_745,N_650);
nand U1336 (N_1336,N_729,N_821);
nand U1337 (N_1337,N_513,N_562);
xnor U1338 (N_1338,N_594,N_650);
nor U1339 (N_1339,N_527,N_623);
and U1340 (N_1340,N_549,N_830);
nand U1341 (N_1341,N_861,N_844);
and U1342 (N_1342,N_514,N_530);
and U1343 (N_1343,N_512,N_606);
or U1344 (N_1344,N_739,N_691);
nand U1345 (N_1345,N_673,N_860);
and U1346 (N_1346,N_606,N_977);
nand U1347 (N_1347,N_796,N_706);
nand U1348 (N_1348,N_733,N_724);
nand U1349 (N_1349,N_525,N_734);
and U1350 (N_1350,N_805,N_543);
nor U1351 (N_1351,N_670,N_986);
nand U1352 (N_1352,N_758,N_750);
or U1353 (N_1353,N_908,N_723);
and U1354 (N_1354,N_807,N_837);
xnor U1355 (N_1355,N_711,N_548);
nand U1356 (N_1356,N_984,N_541);
nor U1357 (N_1357,N_604,N_508);
and U1358 (N_1358,N_770,N_545);
nand U1359 (N_1359,N_689,N_576);
nor U1360 (N_1360,N_983,N_946);
and U1361 (N_1361,N_786,N_986);
and U1362 (N_1362,N_793,N_770);
nand U1363 (N_1363,N_602,N_749);
nand U1364 (N_1364,N_992,N_887);
nor U1365 (N_1365,N_974,N_562);
and U1366 (N_1366,N_561,N_907);
or U1367 (N_1367,N_530,N_628);
nand U1368 (N_1368,N_920,N_904);
or U1369 (N_1369,N_993,N_820);
or U1370 (N_1370,N_750,N_711);
nand U1371 (N_1371,N_680,N_737);
nand U1372 (N_1372,N_935,N_688);
nand U1373 (N_1373,N_940,N_954);
nand U1374 (N_1374,N_698,N_934);
or U1375 (N_1375,N_575,N_854);
and U1376 (N_1376,N_617,N_993);
nand U1377 (N_1377,N_901,N_579);
and U1378 (N_1378,N_785,N_846);
nor U1379 (N_1379,N_833,N_736);
nor U1380 (N_1380,N_647,N_706);
or U1381 (N_1381,N_822,N_989);
or U1382 (N_1382,N_752,N_831);
or U1383 (N_1383,N_854,N_951);
or U1384 (N_1384,N_763,N_511);
nand U1385 (N_1385,N_844,N_837);
or U1386 (N_1386,N_533,N_808);
nor U1387 (N_1387,N_862,N_755);
or U1388 (N_1388,N_511,N_628);
nand U1389 (N_1389,N_912,N_536);
and U1390 (N_1390,N_908,N_525);
nor U1391 (N_1391,N_857,N_501);
nor U1392 (N_1392,N_904,N_592);
nor U1393 (N_1393,N_684,N_691);
nand U1394 (N_1394,N_870,N_652);
and U1395 (N_1395,N_565,N_917);
and U1396 (N_1396,N_750,N_924);
nor U1397 (N_1397,N_877,N_529);
nor U1398 (N_1398,N_570,N_711);
nand U1399 (N_1399,N_933,N_884);
nand U1400 (N_1400,N_973,N_731);
and U1401 (N_1401,N_512,N_542);
and U1402 (N_1402,N_563,N_834);
or U1403 (N_1403,N_953,N_709);
or U1404 (N_1404,N_667,N_990);
or U1405 (N_1405,N_875,N_667);
and U1406 (N_1406,N_536,N_866);
nand U1407 (N_1407,N_524,N_699);
and U1408 (N_1408,N_595,N_908);
nand U1409 (N_1409,N_647,N_884);
and U1410 (N_1410,N_705,N_850);
nand U1411 (N_1411,N_989,N_673);
nor U1412 (N_1412,N_509,N_982);
and U1413 (N_1413,N_588,N_930);
nor U1414 (N_1414,N_595,N_794);
nor U1415 (N_1415,N_993,N_975);
or U1416 (N_1416,N_572,N_785);
nor U1417 (N_1417,N_690,N_884);
and U1418 (N_1418,N_847,N_992);
and U1419 (N_1419,N_697,N_946);
or U1420 (N_1420,N_974,N_713);
or U1421 (N_1421,N_970,N_972);
and U1422 (N_1422,N_685,N_534);
and U1423 (N_1423,N_967,N_952);
or U1424 (N_1424,N_526,N_879);
nor U1425 (N_1425,N_906,N_502);
or U1426 (N_1426,N_701,N_836);
nor U1427 (N_1427,N_692,N_805);
nand U1428 (N_1428,N_704,N_962);
or U1429 (N_1429,N_921,N_875);
or U1430 (N_1430,N_626,N_879);
nand U1431 (N_1431,N_646,N_685);
nor U1432 (N_1432,N_874,N_617);
xnor U1433 (N_1433,N_840,N_881);
nor U1434 (N_1434,N_751,N_785);
and U1435 (N_1435,N_623,N_528);
nor U1436 (N_1436,N_559,N_905);
nand U1437 (N_1437,N_826,N_511);
nand U1438 (N_1438,N_507,N_892);
and U1439 (N_1439,N_744,N_687);
nand U1440 (N_1440,N_884,N_593);
nor U1441 (N_1441,N_625,N_958);
and U1442 (N_1442,N_700,N_802);
nand U1443 (N_1443,N_904,N_969);
or U1444 (N_1444,N_596,N_995);
and U1445 (N_1445,N_568,N_818);
and U1446 (N_1446,N_574,N_873);
nor U1447 (N_1447,N_799,N_932);
or U1448 (N_1448,N_837,N_630);
or U1449 (N_1449,N_597,N_602);
and U1450 (N_1450,N_520,N_719);
nor U1451 (N_1451,N_658,N_808);
nand U1452 (N_1452,N_875,N_570);
nor U1453 (N_1453,N_971,N_930);
or U1454 (N_1454,N_735,N_873);
and U1455 (N_1455,N_516,N_902);
nor U1456 (N_1456,N_739,N_697);
and U1457 (N_1457,N_510,N_696);
nand U1458 (N_1458,N_608,N_815);
or U1459 (N_1459,N_823,N_739);
nor U1460 (N_1460,N_524,N_962);
or U1461 (N_1461,N_727,N_978);
and U1462 (N_1462,N_988,N_726);
nand U1463 (N_1463,N_849,N_571);
nand U1464 (N_1464,N_702,N_842);
or U1465 (N_1465,N_958,N_815);
or U1466 (N_1466,N_517,N_701);
and U1467 (N_1467,N_711,N_777);
nor U1468 (N_1468,N_857,N_679);
nor U1469 (N_1469,N_596,N_967);
nand U1470 (N_1470,N_514,N_618);
and U1471 (N_1471,N_977,N_773);
or U1472 (N_1472,N_791,N_898);
and U1473 (N_1473,N_610,N_932);
and U1474 (N_1474,N_845,N_721);
nand U1475 (N_1475,N_714,N_924);
nand U1476 (N_1476,N_549,N_845);
nand U1477 (N_1477,N_840,N_662);
nor U1478 (N_1478,N_952,N_883);
nand U1479 (N_1479,N_913,N_844);
and U1480 (N_1480,N_759,N_749);
nor U1481 (N_1481,N_844,N_882);
nand U1482 (N_1482,N_858,N_761);
or U1483 (N_1483,N_900,N_938);
and U1484 (N_1484,N_983,N_884);
or U1485 (N_1485,N_838,N_818);
and U1486 (N_1486,N_807,N_968);
nor U1487 (N_1487,N_977,N_992);
nand U1488 (N_1488,N_671,N_655);
or U1489 (N_1489,N_730,N_565);
nand U1490 (N_1490,N_650,N_619);
or U1491 (N_1491,N_974,N_501);
and U1492 (N_1492,N_959,N_942);
or U1493 (N_1493,N_922,N_699);
nor U1494 (N_1494,N_919,N_739);
or U1495 (N_1495,N_944,N_893);
or U1496 (N_1496,N_547,N_738);
nor U1497 (N_1497,N_592,N_869);
nor U1498 (N_1498,N_787,N_788);
nor U1499 (N_1499,N_881,N_947);
and U1500 (N_1500,N_1116,N_1275);
and U1501 (N_1501,N_1355,N_1246);
and U1502 (N_1502,N_1405,N_1408);
nor U1503 (N_1503,N_1137,N_1264);
or U1504 (N_1504,N_1345,N_1253);
or U1505 (N_1505,N_1321,N_1184);
nor U1506 (N_1506,N_1258,N_1112);
and U1507 (N_1507,N_1295,N_1333);
or U1508 (N_1508,N_1243,N_1160);
and U1509 (N_1509,N_1127,N_1259);
or U1510 (N_1510,N_1149,N_1486);
nor U1511 (N_1511,N_1226,N_1467);
nand U1512 (N_1512,N_1483,N_1182);
nand U1513 (N_1513,N_1366,N_1435);
and U1514 (N_1514,N_1474,N_1393);
nand U1515 (N_1515,N_1102,N_1398);
or U1516 (N_1516,N_1278,N_1338);
or U1517 (N_1517,N_1005,N_1101);
xor U1518 (N_1518,N_1011,N_1097);
or U1519 (N_1519,N_1282,N_1456);
and U1520 (N_1520,N_1470,N_1285);
nand U1521 (N_1521,N_1340,N_1047);
nand U1522 (N_1522,N_1466,N_1414);
and U1523 (N_1523,N_1025,N_1214);
nor U1524 (N_1524,N_1030,N_1409);
or U1525 (N_1525,N_1225,N_1114);
and U1526 (N_1526,N_1041,N_1000);
nor U1527 (N_1527,N_1187,N_1056);
or U1528 (N_1528,N_1147,N_1174);
nand U1529 (N_1529,N_1216,N_1058);
nand U1530 (N_1530,N_1150,N_1080);
or U1531 (N_1531,N_1165,N_1015);
nor U1532 (N_1532,N_1337,N_1077);
or U1533 (N_1533,N_1177,N_1403);
nor U1534 (N_1534,N_1031,N_1069);
nor U1535 (N_1535,N_1319,N_1361);
and U1536 (N_1536,N_1176,N_1021);
or U1537 (N_1537,N_1094,N_1286);
nor U1538 (N_1538,N_1054,N_1356);
nand U1539 (N_1539,N_1382,N_1477);
and U1540 (N_1540,N_1059,N_1302);
or U1541 (N_1541,N_1301,N_1341);
and U1542 (N_1542,N_1084,N_1418);
and U1543 (N_1543,N_1252,N_1083);
nand U1544 (N_1544,N_1230,N_1202);
nor U1545 (N_1545,N_1063,N_1436);
nand U1546 (N_1546,N_1003,N_1429);
or U1547 (N_1547,N_1343,N_1401);
nor U1548 (N_1548,N_1048,N_1368);
nand U1549 (N_1549,N_1392,N_1499);
nor U1550 (N_1550,N_1210,N_1411);
nand U1551 (N_1551,N_1215,N_1413);
nor U1552 (N_1552,N_1068,N_1035);
nor U1553 (N_1553,N_1399,N_1380);
nand U1554 (N_1554,N_1189,N_1120);
or U1555 (N_1555,N_1344,N_1296);
or U1556 (N_1556,N_1490,N_1001);
nand U1557 (N_1557,N_1416,N_1424);
nor U1558 (N_1558,N_1024,N_1394);
or U1559 (N_1559,N_1208,N_1211);
or U1560 (N_1560,N_1240,N_1062);
and U1561 (N_1561,N_1316,N_1133);
nor U1562 (N_1562,N_1373,N_1004);
and U1563 (N_1563,N_1443,N_1363);
nor U1564 (N_1564,N_1110,N_1449);
or U1565 (N_1565,N_1379,N_1061);
nand U1566 (N_1566,N_1152,N_1014);
and U1567 (N_1567,N_1064,N_1100);
and U1568 (N_1568,N_1417,N_1346);
and U1569 (N_1569,N_1268,N_1447);
or U1570 (N_1570,N_1348,N_1074);
and U1571 (N_1571,N_1075,N_1153);
or U1572 (N_1572,N_1023,N_1205);
nor U1573 (N_1573,N_1495,N_1406);
nand U1574 (N_1574,N_1428,N_1473);
nor U1575 (N_1575,N_1260,N_1249);
nor U1576 (N_1576,N_1010,N_1318);
nor U1577 (N_1577,N_1197,N_1026);
and U1578 (N_1578,N_1376,N_1088);
nand U1579 (N_1579,N_1217,N_1493);
and U1580 (N_1580,N_1463,N_1172);
xor U1581 (N_1581,N_1335,N_1310);
and U1582 (N_1582,N_1410,N_1300);
or U1583 (N_1583,N_1146,N_1385);
nand U1584 (N_1584,N_1288,N_1272);
or U1585 (N_1585,N_1257,N_1207);
and U1586 (N_1586,N_1388,N_1081);
or U1587 (N_1587,N_1400,N_1314);
or U1588 (N_1588,N_1232,N_1455);
nand U1589 (N_1589,N_1175,N_1224);
nand U1590 (N_1590,N_1007,N_1038);
and U1591 (N_1591,N_1108,N_1183);
nor U1592 (N_1592,N_1421,N_1471);
or U1593 (N_1593,N_1046,N_1496);
nor U1594 (N_1594,N_1027,N_1076);
or U1595 (N_1595,N_1485,N_1367);
and U1596 (N_1596,N_1298,N_1129);
nand U1597 (N_1597,N_1223,N_1292);
nand U1598 (N_1598,N_1180,N_1441);
or U1599 (N_1599,N_1209,N_1434);
nand U1600 (N_1600,N_1099,N_1248);
nor U1601 (N_1601,N_1142,N_1353);
nor U1602 (N_1602,N_1154,N_1482);
nor U1603 (N_1603,N_1136,N_1008);
nor U1604 (N_1604,N_1096,N_1036);
or U1605 (N_1605,N_1322,N_1185);
nor U1606 (N_1606,N_1438,N_1148);
nand U1607 (N_1607,N_1073,N_1118);
and U1608 (N_1608,N_1238,N_1093);
and U1609 (N_1609,N_1186,N_1053);
and U1610 (N_1610,N_1378,N_1109);
and U1611 (N_1611,N_1254,N_1289);
nor U1612 (N_1612,N_1130,N_1022);
and U1613 (N_1613,N_1283,N_1122);
nand U1614 (N_1614,N_1263,N_1126);
or U1615 (N_1615,N_1281,N_1370);
and U1616 (N_1616,N_1028,N_1293);
and U1617 (N_1617,N_1279,N_1043);
nor U1618 (N_1618,N_1222,N_1395);
nor U1619 (N_1619,N_1018,N_1291);
nor U1620 (N_1620,N_1212,N_1372);
or U1621 (N_1621,N_1044,N_1389);
or U1622 (N_1622,N_1359,N_1419);
or U1623 (N_1623,N_1358,N_1488);
nand U1624 (N_1624,N_1432,N_1237);
or U1625 (N_1625,N_1362,N_1071);
nor U1626 (N_1626,N_1271,N_1190);
or U1627 (N_1627,N_1082,N_1095);
nor U1628 (N_1628,N_1227,N_1104);
nor U1629 (N_1629,N_1342,N_1002);
or U1630 (N_1630,N_1234,N_1369);
or U1631 (N_1631,N_1461,N_1164);
or U1632 (N_1632,N_1173,N_1312);
and U1633 (N_1633,N_1420,N_1480);
or U1634 (N_1634,N_1135,N_1060);
nor U1635 (N_1635,N_1475,N_1115);
nor U1636 (N_1636,N_1422,N_1006);
nor U1637 (N_1637,N_1103,N_1241);
or U1638 (N_1638,N_1009,N_1313);
and U1639 (N_1639,N_1427,N_1119);
or U1640 (N_1640,N_1171,N_1303);
and U1641 (N_1641,N_1269,N_1347);
nor U1642 (N_1642,N_1106,N_1016);
nand U1643 (N_1643,N_1323,N_1228);
and U1644 (N_1644,N_1045,N_1251);
or U1645 (N_1645,N_1280,N_1066);
or U1646 (N_1646,N_1140,N_1162);
and U1647 (N_1647,N_1229,N_1049);
nor U1648 (N_1648,N_1277,N_1247);
nand U1649 (N_1649,N_1448,N_1381);
nor U1650 (N_1650,N_1206,N_1360);
and U1651 (N_1651,N_1188,N_1377);
nor U1652 (N_1652,N_1452,N_1105);
and U1653 (N_1653,N_1270,N_1426);
nand U1654 (N_1654,N_1236,N_1297);
nor U1655 (N_1655,N_1339,N_1364);
nand U1656 (N_1656,N_1325,N_1161);
or U1657 (N_1657,N_1498,N_1351);
nand U1658 (N_1658,N_1086,N_1425);
nand U1659 (N_1659,N_1163,N_1334);
nor U1660 (N_1660,N_1092,N_1042);
or U1661 (N_1661,N_1065,N_1201);
and U1662 (N_1662,N_1191,N_1431);
nand U1663 (N_1663,N_1111,N_1087);
or U1664 (N_1664,N_1132,N_1446);
and U1665 (N_1665,N_1294,N_1052);
and U1666 (N_1666,N_1158,N_1039);
and U1667 (N_1667,N_1433,N_1194);
and U1668 (N_1668,N_1013,N_1218);
nand U1669 (N_1669,N_1117,N_1451);
nor U1670 (N_1670,N_1145,N_1315);
nor U1671 (N_1671,N_1469,N_1274);
or U1672 (N_1672,N_1309,N_1440);
nand U1673 (N_1673,N_1349,N_1311);
nand U1674 (N_1674,N_1179,N_1196);
or U1675 (N_1675,N_1078,N_1113);
nand U1676 (N_1676,N_1487,N_1267);
or U1677 (N_1677,N_1037,N_1131);
nand U1678 (N_1678,N_1442,N_1462);
nor U1679 (N_1679,N_1199,N_1465);
or U1680 (N_1680,N_1166,N_1144);
or U1681 (N_1681,N_1012,N_1139);
nor U1682 (N_1682,N_1261,N_1134);
nand U1683 (N_1683,N_1244,N_1407);
or U1684 (N_1684,N_1235,N_1329);
nor U1685 (N_1685,N_1181,N_1423);
or U1686 (N_1686,N_1159,N_1320);
and U1687 (N_1687,N_1157,N_1330);
and U1688 (N_1688,N_1479,N_1307);
or U1689 (N_1689,N_1284,N_1266);
or U1690 (N_1690,N_1265,N_1067);
or U1691 (N_1691,N_1029,N_1481);
nor U1692 (N_1692,N_1437,N_1085);
nor U1693 (N_1693,N_1444,N_1245);
and U1694 (N_1694,N_1231,N_1445);
nor U1695 (N_1695,N_1458,N_1387);
or U1696 (N_1696,N_1138,N_1170);
and U1697 (N_1697,N_1412,N_1352);
nand U1698 (N_1698,N_1220,N_1213);
or U1699 (N_1699,N_1178,N_1478);
xnor U1700 (N_1700,N_1365,N_1121);
nor U1701 (N_1701,N_1090,N_1386);
nand U1702 (N_1702,N_1169,N_1304);
and U1703 (N_1703,N_1439,N_1290);
nor U1704 (N_1704,N_1040,N_1256);
or U1705 (N_1705,N_1384,N_1453);
nor U1706 (N_1706,N_1255,N_1391);
and U1707 (N_1707,N_1331,N_1476);
nor U1708 (N_1708,N_1242,N_1089);
nor U1709 (N_1709,N_1489,N_1203);
xor U1710 (N_1710,N_1107,N_1468);
or U1711 (N_1711,N_1198,N_1193);
or U1712 (N_1712,N_1156,N_1155);
and U1713 (N_1713,N_1354,N_1195);
xor U1714 (N_1714,N_1276,N_1430);
and U1715 (N_1715,N_1192,N_1051);
nand U1716 (N_1716,N_1459,N_1200);
nor U1717 (N_1717,N_1327,N_1492);
or U1718 (N_1718,N_1057,N_1305);
or U1719 (N_1719,N_1221,N_1472);
nor U1720 (N_1720,N_1262,N_1494);
or U1721 (N_1721,N_1123,N_1141);
nor U1722 (N_1722,N_1460,N_1143);
nand U1723 (N_1723,N_1032,N_1404);
or U1724 (N_1724,N_1374,N_1306);
nor U1725 (N_1725,N_1033,N_1034);
nand U1726 (N_1726,N_1128,N_1125);
nor U1727 (N_1727,N_1019,N_1396);
and U1728 (N_1728,N_1020,N_1375);
nor U1729 (N_1729,N_1357,N_1390);
or U1730 (N_1730,N_1317,N_1239);
or U1731 (N_1731,N_1336,N_1332);
or U1732 (N_1732,N_1328,N_1457);
and U1733 (N_1733,N_1464,N_1072);
or U1734 (N_1734,N_1151,N_1050);
or U1735 (N_1735,N_1491,N_1350);
and U1736 (N_1736,N_1308,N_1287);
and U1737 (N_1737,N_1079,N_1415);
or U1738 (N_1738,N_1454,N_1402);
and U1739 (N_1739,N_1383,N_1299);
or U1740 (N_1740,N_1371,N_1098);
and U1741 (N_1741,N_1091,N_1250);
nor U1742 (N_1742,N_1204,N_1168);
nor U1743 (N_1743,N_1219,N_1484);
or U1744 (N_1744,N_1324,N_1450);
or U1745 (N_1745,N_1124,N_1497);
or U1746 (N_1746,N_1397,N_1017);
or U1747 (N_1747,N_1326,N_1273);
and U1748 (N_1748,N_1055,N_1070);
and U1749 (N_1749,N_1167,N_1233);
or U1750 (N_1750,N_1351,N_1370);
nor U1751 (N_1751,N_1040,N_1456);
or U1752 (N_1752,N_1456,N_1356);
nor U1753 (N_1753,N_1445,N_1199);
or U1754 (N_1754,N_1147,N_1425);
and U1755 (N_1755,N_1012,N_1471);
nand U1756 (N_1756,N_1363,N_1385);
and U1757 (N_1757,N_1011,N_1074);
nand U1758 (N_1758,N_1061,N_1269);
nor U1759 (N_1759,N_1057,N_1145);
nor U1760 (N_1760,N_1313,N_1166);
nor U1761 (N_1761,N_1297,N_1216);
nor U1762 (N_1762,N_1420,N_1033);
nand U1763 (N_1763,N_1161,N_1212);
and U1764 (N_1764,N_1049,N_1082);
nor U1765 (N_1765,N_1306,N_1381);
or U1766 (N_1766,N_1267,N_1174);
nand U1767 (N_1767,N_1494,N_1177);
or U1768 (N_1768,N_1332,N_1208);
or U1769 (N_1769,N_1022,N_1219);
and U1770 (N_1770,N_1463,N_1363);
and U1771 (N_1771,N_1250,N_1323);
or U1772 (N_1772,N_1200,N_1086);
nor U1773 (N_1773,N_1482,N_1163);
and U1774 (N_1774,N_1422,N_1499);
nor U1775 (N_1775,N_1062,N_1412);
nor U1776 (N_1776,N_1436,N_1026);
and U1777 (N_1777,N_1498,N_1499);
nor U1778 (N_1778,N_1140,N_1316);
nand U1779 (N_1779,N_1216,N_1343);
nand U1780 (N_1780,N_1027,N_1081);
nand U1781 (N_1781,N_1028,N_1400);
nor U1782 (N_1782,N_1200,N_1120);
nand U1783 (N_1783,N_1324,N_1328);
nor U1784 (N_1784,N_1186,N_1434);
nor U1785 (N_1785,N_1375,N_1062);
nand U1786 (N_1786,N_1420,N_1324);
and U1787 (N_1787,N_1378,N_1200);
or U1788 (N_1788,N_1324,N_1032);
nor U1789 (N_1789,N_1485,N_1326);
and U1790 (N_1790,N_1265,N_1132);
nand U1791 (N_1791,N_1298,N_1043);
xor U1792 (N_1792,N_1371,N_1177);
nand U1793 (N_1793,N_1207,N_1037);
nand U1794 (N_1794,N_1348,N_1477);
nand U1795 (N_1795,N_1170,N_1372);
and U1796 (N_1796,N_1351,N_1424);
and U1797 (N_1797,N_1256,N_1457);
nand U1798 (N_1798,N_1144,N_1456);
or U1799 (N_1799,N_1244,N_1099);
or U1800 (N_1800,N_1120,N_1180);
nand U1801 (N_1801,N_1175,N_1172);
and U1802 (N_1802,N_1354,N_1119);
or U1803 (N_1803,N_1209,N_1088);
or U1804 (N_1804,N_1138,N_1187);
nand U1805 (N_1805,N_1267,N_1433);
nand U1806 (N_1806,N_1039,N_1278);
and U1807 (N_1807,N_1058,N_1422);
or U1808 (N_1808,N_1017,N_1452);
or U1809 (N_1809,N_1476,N_1491);
or U1810 (N_1810,N_1383,N_1298);
nand U1811 (N_1811,N_1037,N_1306);
or U1812 (N_1812,N_1319,N_1393);
or U1813 (N_1813,N_1441,N_1177);
nand U1814 (N_1814,N_1293,N_1123);
and U1815 (N_1815,N_1102,N_1035);
and U1816 (N_1816,N_1222,N_1337);
and U1817 (N_1817,N_1287,N_1066);
and U1818 (N_1818,N_1158,N_1064);
and U1819 (N_1819,N_1147,N_1469);
or U1820 (N_1820,N_1449,N_1498);
nand U1821 (N_1821,N_1281,N_1082);
or U1822 (N_1822,N_1120,N_1338);
nor U1823 (N_1823,N_1119,N_1012);
or U1824 (N_1824,N_1329,N_1454);
or U1825 (N_1825,N_1148,N_1370);
nor U1826 (N_1826,N_1383,N_1468);
and U1827 (N_1827,N_1472,N_1001);
nor U1828 (N_1828,N_1001,N_1222);
nand U1829 (N_1829,N_1056,N_1109);
or U1830 (N_1830,N_1158,N_1117);
nor U1831 (N_1831,N_1317,N_1095);
nor U1832 (N_1832,N_1319,N_1173);
nor U1833 (N_1833,N_1261,N_1149);
and U1834 (N_1834,N_1343,N_1335);
nand U1835 (N_1835,N_1432,N_1062);
nand U1836 (N_1836,N_1142,N_1457);
nor U1837 (N_1837,N_1222,N_1235);
or U1838 (N_1838,N_1411,N_1372);
xor U1839 (N_1839,N_1492,N_1236);
and U1840 (N_1840,N_1277,N_1170);
or U1841 (N_1841,N_1383,N_1046);
or U1842 (N_1842,N_1190,N_1407);
and U1843 (N_1843,N_1254,N_1070);
nand U1844 (N_1844,N_1201,N_1164);
nand U1845 (N_1845,N_1282,N_1127);
nand U1846 (N_1846,N_1018,N_1150);
nand U1847 (N_1847,N_1465,N_1055);
and U1848 (N_1848,N_1389,N_1356);
nor U1849 (N_1849,N_1223,N_1387);
and U1850 (N_1850,N_1350,N_1450);
and U1851 (N_1851,N_1469,N_1240);
nor U1852 (N_1852,N_1453,N_1077);
nand U1853 (N_1853,N_1329,N_1497);
nand U1854 (N_1854,N_1101,N_1275);
nand U1855 (N_1855,N_1217,N_1334);
nand U1856 (N_1856,N_1216,N_1464);
or U1857 (N_1857,N_1482,N_1495);
nand U1858 (N_1858,N_1149,N_1331);
or U1859 (N_1859,N_1499,N_1154);
and U1860 (N_1860,N_1420,N_1000);
or U1861 (N_1861,N_1370,N_1139);
or U1862 (N_1862,N_1060,N_1139);
nor U1863 (N_1863,N_1466,N_1119);
or U1864 (N_1864,N_1483,N_1024);
or U1865 (N_1865,N_1166,N_1101);
nor U1866 (N_1866,N_1344,N_1397);
nor U1867 (N_1867,N_1374,N_1404);
nand U1868 (N_1868,N_1292,N_1062);
or U1869 (N_1869,N_1371,N_1235);
nor U1870 (N_1870,N_1106,N_1388);
xor U1871 (N_1871,N_1479,N_1346);
nor U1872 (N_1872,N_1207,N_1375);
and U1873 (N_1873,N_1287,N_1288);
nand U1874 (N_1874,N_1056,N_1104);
nand U1875 (N_1875,N_1117,N_1461);
nor U1876 (N_1876,N_1318,N_1017);
nor U1877 (N_1877,N_1436,N_1183);
and U1878 (N_1878,N_1041,N_1446);
and U1879 (N_1879,N_1485,N_1222);
or U1880 (N_1880,N_1226,N_1425);
nor U1881 (N_1881,N_1203,N_1137);
nor U1882 (N_1882,N_1380,N_1128);
or U1883 (N_1883,N_1233,N_1146);
nand U1884 (N_1884,N_1249,N_1497);
nor U1885 (N_1885,N_1117,N_1367);
or U1886 (N_1886,N_1315,N_1219);
nand U1887 (N_1887,N_1035,N_1257);
or U1888 (N_1888,N_1128,N_1041);
or U1889 (N_1889,N_1129,N_1447);
and U1890 (N_1890,N_1191,N_1334);
nand U1891 (N_1891,N_1481,N_1389);
nand U1892 (N_1892,N_1178,N_1001);
or U1893 (N_1893,N_1063,N_1308);
and U1894 (N_1894,N_1236,N_1497);
nor U1895 (N_1895,N_1207,N_1194);
nor U1896 (N_1896,N_1271,N_1294);
and U1897 (N_1897,N_1121,N_1327);
nor U1898 (N_1898,N_1411,N_1266);
nand U1899 (N_1899,N_1310,N_1309);
nand U1900 (N_1900,N_1030,N_1168);
or U1901 (N_1901,N_1079,N_1478);
nand U1902 (N_1902,N_1094,N_1428);
nor U1903 (N_1903,N_1408,N_1080);
and U1904 (N_1904,N_1148,N_1184);
nor U1905 (N_1905,N_1499,N_1236);
nor U1906 (N_1906,N_1102,N_1018);
nand U1907 (N_1907,N_1104,N_1218);
or U1908 (N_1908,N_1428,N_1409);
or U1909 (N_1909,N_1329,N_1472);
or U1910 (N_1910,N_1436,N_1355);
nor U1911 (N_1911,N_1091,N_1381);
and U1912 (N_1912,N_1339,N_1430);
xnor U1913 (N_1913,N_1054,N_1477);
or U1914 (N_1914,N_1157,N_1419);
and U1915 (N_1915,N_1370,N_1292);
or U1916 (N_1916,N_1245,N_1195);
or U1917 (N_1917,N_1321,N_1065);
or U1918 (N_1918,N_1448,N_1075);
nor U1919 (N_1919,N_1145,N_1033);
and U1920 (N_1920,N_1432,N_1225);
or U1921 (N_1921,N_1209,N_1454);
and U1922 (N_1922,N_1298,N_1253);
or U1923 (N_1923,N_1321,N_1325);
nor U1924 (N_1924,N_1055,N_1039);
or U1925 (N_1925,N_1225,N_1246);
nor U1926 (N_1926,N_1312,N_1299);
or U1927 (N_1927,N_1090,N_1493);
nand U1928 (N_1928,N_1288,N_1232);
and U1929 (N_1929,N_1216,N_1166);
and U1930 (N_1930,N_1408,N_1216);
or U1931 (N_1931,N_1182,N_1265);
nand U1932 (N_1932,N_1032,N_1084);
nor U1933 (N_1933,N_1469,N_1438);
and U1934 (N_1934,N_1491,N_1473);
nor U1935 (N_1935,N_1047,N_1235);
or U1936 (N_1936,N_1363,N_1402);
nand U1937 (N_1937,N_1226,N_1308);
nand U1938 (N_1938,N_1190,N_1376);
nand U1939 (N_1939,N_1295,N_1411);
and U1940 (N_1940,N_1054,N_1185);
and U1941 (N_1941,N_1088,N_1272);
and U1942 (N_1942,N_1090,N_1071);
and U1943 (N_1943,N_1090,N_1317);
nand U1944 (N_1944,N_1489,N_1447);
nand U1945 (N_1945,N_1123,N_1345);
and U1946 (N_1946,N_1360,N_1000);
and U1947 (N_1947,N_1005,N_1200);
nand U1948 (N_1948,N_1020,N_1349);
nor U1949 (N_1949,N_1053,N_1270);
and U1950 (N_1950,N_1137,N_1465);
or U1951 (N_1951,N_1176,N_1135);
nand U1952 (N_1952,N_1458,N_1261);
xor U1953 (N_1953,N_1362,N_1304);
nor U1954 (N_1954,N_1091,N_1143);
and U1955 (N_1955,N_1137,N_1334);
nor U1956 (N_1956,N_1393,N_1249);
and U1957 (N_1957,N_1197,N_1165);
nor U1958 (N_1958,N_1213,N_1429);
nor U1959 (N_1959,N_1159,N_1221);
and U1960 (N_1960,N_1248,N_1463);
nand U1961 (N_1961,N_1168,N_1072);
and U1962 (N_1962,N_1206,N_1173);
nand U1963 (N_1963,N_1362,N_1196);
nand U1964 (N_1964,N_1359,N_1271);
or U1965 (N_1965,N_1414,N_1448);
nand U1966 (N_1966,N_1277,N_1057);
nor U1967 (N_1967,N_1233,N_1222);
nor U1968 (N_1968,N_1340,N_1442);
nand U1969 (N_1969,N_1447,N_1177);
nor U1970 (N_1970,N_1024,N_1306);
or U1971 (N_1971,N_1281,N_1156);
xor U1972 (N_1972,N_1235,N_1415);
and U1973 (N_1973,N_1022,N_1238);
or U1974 (N_1974,N_1412,N_1277);
nand U1975 (N_1975,N_1254,N_1033);
nor U1976 (N_1976,N_1150,N_1158);
xor U1977 (N_1977,N_1407,N_1050);
and U1978 (N_1978,N_1328,N_1251);
or U1979 (N_1979,N_1276,N_1433);
or U1980 (N_1980,N_1031,N_1290);
and U1981 (N_1981,N_1028,N_1480);
or U1982 (N_1982,N_1114,N_1075);
and U1983 (N_1983,N_1177,N_1098);
or U1984 (N_1984,N_1227,N_1397);
nand U1985 (N_1985,N_1248,N_1487);
and U1986 (N_1986,N_1321,N_1233);
and U1987 (N_1987,N_1391,N_1178);
and U1988 (N_1988,N_1256,N_1264);
or U1989 (N_1989,N_1002,N_1149);
and U1990 (N_1990,N_1388,N_1004);
and U1991 (N_1991,N_1316,N_1131);
and U1992 (N_1992,N_1384,N_1235);
nand U1993 (N_1993,N_1110,N_1391);
nand U1994 (N_1994,N_1164,N_1363);
nand U1995 (N_1995,N_1214,N_1142);
or U1996 (N_1996,N_1040,N_1355);
or U1997 (N_1997,N_1174,N_1055);
nor U1998 (N_1998,N_1272,N_1265);
and U1999 (N_1999,N_1112,N_1016);
and U2000 (N_2000,N_1529,N_1650);
or U2001 (N_2001,N_1520,N_1987);
nand U2002 (N_2002,N_1672,N_1569);
or U2003 (N_2003,N_1622,N_1904);
or U2004 (N_2004,N_1628,N_1631);
or U2005 (N_2005,N_1821,N_1866);
or U2006 (N_2006,N_1928,N_1571);
or U2007 (N_2007,N_1759,N_1875);
or U2008 (N_2008,N_1990,N_1692);
nand U2009 (N_2009,N_1696,N_1828);
nor U2010 (N_2010,N_1547,N_1732);
nor U2011 (N_2011,N_1906,N_1666);
nand U2012 (N_2012,N_1534,N_1818);
nand U2013 (N_2013,N_1680,N_1761);
or U2014 (N_2014,N_1936,N_1537);
and U2015 (N_2015,N_1823,N_1768);
and U2016 (N_2016,N_1796,N_1709);
nor U2017 (N_2017,N_1740,N_1797);
and U2018 (N_2018,N_1954,N_1703);
nor U2019 (N_2019,N_1806,N_1746);
nor U2020 (N_2020,N_1671,N_1829);
nor U2021 (N_2021,N_1659,N_1813);
and U2022 (N_2022,N_1728,N_1771);
nor U2023 (N_2023,N_1785,N_1519);
nor U2024 (N_2024,N_1763,N_1981);
nor U2025 (N_2025,N_1688,N_1691);
nand U2026 (N_2026,N_1645,N_1675);
nor U2027 (N_2027,N_1798,N_1802);
nand U2028 (N_2028,N_1749,N_1634);
nor U2029 (N_2029,N_1915,N_1863);
nor U2030 (N_2030,N_1725,N_1794);
and U2031 (N_2031,N_1830,N_1572);
and U2032 (N_2032,N_1862,N_1879);
and U2033 (N_2033,N_1908,N_1530);
nand U2034 (N_2034,N_1847,N_1963);
and U2035 (N_2035,N_1930,N_1948);
or U2036 (N_2036,N_1809,N_1870);
nand U2037 (N_2037,N_1722,N_1550);
nor U2038 (N_2038,N_1651,N_1783);
or U2039 (N_2039,N_1535,N_1943);
and U2040 (N_2040,N_1678,N_1734);
nor U2041 (N_2041,N_1514,N_1881);
and U2042 (N_2042,N_1557,N_1882);
and U2043 (N_2043,N_1538,N_1938);
nand U2044 (N_2044,N_1695,N_1625);
and U2045 (N_2045,N_1949,N_1561);
or U2046 (N_2046,N_1834,N_1737);
and U2047 (N_2047,N_1873,N_1974);
or U2048 (N_2048,N_1849,N_1854);
or U2049 (N_2049,N_1629,N_1711);
and U2050 (N_2050,N_1694,N_1564);
nand U2051 (N_2051,N_1892,N_1690);
or U2052 (N_2052,N_1613,N_1764);
nor U2053 (N_2053,N_1693,N_1961);
and U2054 (N_2054,N_1889,N_1788);
nor U2055 (N_2055,N_1585,N_1618);
nor U2056 (N_2056,N_1986,N_1833);
xnor U2057 (N_2057,N_1756,N_1998);
and U2058 (N_2058,N_1903,N_1942);
nor U2059 (N_2059,N_1793,N_1861);
or U2060 (N_2060,N_1857,N_1616);
nand U2061 (N_2061,N_1744,N_1837);
nor U2062 (N_2062,N_1518,N_1922);
nand U2063 (N_2063,N_1855,N_1787);
nor U2064 (N_2064,N_1750,N_1820);
or U2065 (N_2065,N_1699,N_1812);
nand U2066 (N_2066,N_1856,N_1864);
or U2067 (N_2067,N_1673,N_1836);
nand U2068 (N_2068,N_1698,N_1975);
and U2069 (N_2069,N_1941,N_1905);
or U2070 (N_2070,N_1839,N_1636);
nor U2071 (N_2071,N_1758,N_1757);
nand U2072 (N_2072,N_1597,N_1884);
nand U2073 (N_2073,N_1517,N_1681);
nor U2074 (N_2074,N_1997,N_1956);
and U2075 (N_2075,N_1623,N_1966);
and U2076 (N_2076,N_1978,N_1951);
nor U2077 (N_2077,N_1633,N_1773);
and U2078 (N_2078,N_1995,N_1977);
or U2079 (N_2079,N_1581,N_1614);
or U2080 (N_2080,N_1924,N_1845);
nor U2081 (N_2081,N_1901,N_1610);
nor U2082 (N_2082,N_1502,N_1540);
or U2083 (N_2083,N_1962,N_1587);
nor U2084 (N_2084,N_1653,N_1742);
nand U2085 (N_2085,N_1810,N_1996);
or U2086 (N_2086,N_1982,N_1669);
nor U2087 (N_2087,N_1670,N_1957);
and U2088 (N_2088,N_1687,N_1710);
or U2089 (N_2089,N_1853,N_1655);
nand U2090 (N_2090,N_1880,N_1824);
and U2091 (N_2091,N_1874,N_1641);
nand U2092 (N_2092,N_1601,N_1707);
nand U2093 (N_2093,N_1804,N_1933);
nand U2094 (N_2094,N_1743,N_1767);
nor U2095 (N_2095,N_1584,N_1781);
and U2096 (N_2096,N_1894,N_1970);
nor U2097 (N_2097,N_1776,N_1549);
nand U2098 (N_2098,N_1638,N_1701);
nor U2099 (N_2099,N_1683,N_1664);
nand U2100 (N_2100,N_1819,N_1512);
nor U2101 (N_2101,N_1643,N_1532);
nand U2102 (N_2102,N_1603,N_1911);
and U2103 (N_2103,N_1567,N_1989);
or U2104 (N_2104,N_1544,N_1604);
nand U2105 (N_2105,N_1891,N_1826);
and U2106 (N_2106,N_1865,N_1927);
or U2107 (N_2107,N_1992,N_1570);
or U2108 (N_2108,N_1723,N_1593);
nor U2109 (N_2109,N_1800,N_1541);
nor U2110 (N_2110,N_1984,N_1971);
nand U2111 (N_2111,N_1575,N_1522);
or U2112 (N_2112,N_1558,N_1685);
nor U2113 (N_2113,N_1913,N_1718);
or U2114 (N_2114,N_1546,N_1775);
and U2115 (N_2115,N_1825,N_1503);
nand U2116 (N_2116,N_1999,N_1955);
nand U2117 (N_2117,N_1607,N_1579);
nand U2118 (N_2118,N_1814,N_1890);
nand U2119 (N_2119,N_1729,N_1686);
nor U2120 (N_2120,N_1751,N_1719);
and U2121 (N_2121,N_1553,N_1554);
nor U2122 (N_2122,N_1720,N_1578);
and U2123 (N_2123,N_1676,N_1510);
nand U2124 (N_2124,N_1566,N_1886);
and U2125 (N_2125,N_1663,N_1619);
and U2126 (N_2126,N_1598,N_1790);
nand U2127 (N_2127,N_1747,N_1586);
nand U2128 (N_2128,N_1795,N_1516);
nor U2129 (N_2129,N_1505,N_1662);
nor U2130 (N_2130,N_1786,N_1762);
nand U2131 (N_2131,N_1934,N_1574);
and U2132 (N_2132,N_1885,N_1868);
and U2133 (N_2133,N_1832,N_1926);
nand U2134 (N_2134,N_1754,N_1646);
nand U2135 (N_2135,N_1594,N_1736);
nand U2136 (N_2136,N_1612,N_1972);
or U2137 (N_2137,N_1748,N_1831);
nor U2138 (N_2138,N_1944,N_1765);
nor U2139 (N_2139,N_1952,N_1624);
and U2140 (N_2140,N_1649,N_1501);
nand U2141 (N_2141,N_1640,N_1967);
nand U2142 (N_2142,N_1543,N_1937);
or U2143 (N_2143,N_1697,N_1850);
or U2144 (N_2144,N_1777,N_1822);
nor U2145 (N_2145,N_1887,N_1876);
nand U2146 (N_2146,N_1991,N_1596);
and U2147 (N_2147,N_1896,N_1976);
and U2148 (N_2148,N_1583,N_1515);
nor U2149 (N_2149,N_1920,N_1621);
nor U2150 (N_2150,N_1968,N_1635);
or U2151 (N_2151,N_1760,N_1925);
or U2152 (N_2152,N_1888,N_1648);
or U2153 (N_2153,N_1741,N_1929);
nor U2154 (N_2154,N_1755,N_1509);
or U2155 (N_2155,N_1657,N_1682);
and U2156 (N_2156,N_1573,N_1595);
and U2157 (N_2157,N_1893,N_1877);
nor U2158 (N_2158,N_1859,N_1656);
or U2159 (N_2159,N_1835,N_1867);
or U2160 (N_2160,N_1801,N_1652);
or U2161 (N_2161,N_1782,N_1559);
nand U2162 (N_2162,N_1947,N_1808);
nand U2163 (N_2163,N_1907,N_1713);
nor U2164 (N_2164,N_1789,N_1735);
or U2165 (N_2165,N_1766,N_1731);
or U2166 (N_2166,N_1917,N_1769);
and U2167 (N_2167,N_1580,N_1939);
or U2168 (N_2168,N_1637,N_1871);
and U2169 (N_2169,N_1902,N_1807);
nor U2170 (N_2170,N_1708,N_1811);
and U2171 (N_2171,N_1883,N_1525);
and U2172 (N_2172,N_1858,N_1803);
nor U2173 (N_2173,N_1983,N_1899);
and U2174 (N_2174,N_1528,N_1668);
and U2175 (N_2175,N_1679,N_1665);
and U2176 (N_2176,N_1506,N_1551);
or U2177 (N_2177,N_1568,N_1960);
and U2178 (N_2178,N_1591,N_1533);
and U2179 (N_2179,N_1620,N_1843);
nand U2180 (N_2180,N_1730,N_1900);
nor U2181 (N_2181,N_1916,N_1545);
or U2182 (N_2182,N_1556,N_1630);
nor U2183 (N_2183,N_1923,N_1919);
nand U2184 (N_2184,N_1774,N_1869);
nand U2185 (N_2185,N_1577,N_1626);
nor U2186 (N_2186,N_1784,N_1935);
and U2187 (N_2187,N_1539,N_1644);
and U2188 (N_2188,N_1851,N_1617);
nand U2189 (N_2189,N_1548,N_1660);
and U2190 (N_2190,N_1827,N_1609);
nand U2191 (N_2191,N_1940,N_1745);
or U2192 (N_2192,N_1508,N_1931);
nand U2193 (N_2193,N_1959,N_1842);
and U2194 (N_2194,N_1689,N_1779);
or U2195 (N_2195,N_1565,N_1964);
and U2196 (N_2196,N_1946,N_1791);
and U2197 (N_2197,N_1932,N_1504);
or U2198 (N_2198,N_1817,N_1582);
or U2199 (N_2199,N_1526,N_1852);
and U2200 (N_2200,N_1969,N_1770);
and U2201 (N_2201,N_1500,N_1642);
nor U2202 (N_2202,N_1844,N_1706);
nor U2203 (N_2203,N_1897,N_1753);
xnor U2204 (N_2204,N_1872,N_1838);
or U2205 (N_2205,N_1552,N_1527);
or U2206 (N_2206,N_1727,N_1599);
or U2207 (N_2207,N_1945,N_1799);
nor U2208 (N_2208,N_1772,N_1684);
or U2209 (N_2209,N_1985,N_1605);
nor U2210 (N_2210,N_1523,N_1531);
nor U2211 (N_2211,N_1717,N_1521);
or U2212 (N_2212,N_1738,N_1592);
and U2213 (N_2213,N_1958,N_1667);
nand U2214 (N_2214,N_1511,N_1627);
nand U2215 (N_2215,N_1606,N_1953);
and U2216 (N_2216,N_1778,N_1815);
nand U2217 (N_2217,N_1705,N_1674);
nor U2218 (N_2218,N_1914,N_1840);
nor U2219 (N_2219,N_1576,N_1700);
nand U2220 (N_2220,N_1846,N_1542);
nand U2221 (N_2221,N_1600,N_1639);
nand U2222 (N_2222,N_1752,N_1715);
or U2223 (N_2223,N_1702,N_1965);
and U2224 (N_2224,N_1816,N_1909);
nand U2225 (N_2225,N_1910,N_1524);
nand U2226 (N_2226,N_1588,N_1860);
and U2227 (N_2227,N_1988,N_1973);
nand U2228 (N_2228,N_1739,N_1608);
nand U2229 (N_2229,N_1780,N_1792);
or U2230 (N_2230,N_1513,N_1980);
nor U2231 (N_2231,N_1805,N_1848);
or U2232 (N_2232,N_1898,N_1562);
or U2233 (N_2233,N_1921,N_1602);
and U2234 (N_2234,N_1979,N_1721);
nor U2235 (N_2235,N_1993,N_1507);
nor U2236 (N_2236,N_1555,N_1994);
nand U2237 (N_2237,N_1733,N_1918);
nor U2238 (N_2238,N_1661,N_1895);
or U2239 (N_2239,N_1912,N_1950);
nor U2240 (N_2240,N_1563,N_1536);
or U2241 (N_2241,N_1704,N_1658);
nand U2242 (N_2242,N_1726,N_1589);
nor U2243 (N_2243,N_1878,N_1714);
or U2244 (N_2244,N_1716,N_1724);
nor U2245 (N_2245,N_1590,N_1841);
nand U2246 (N_2246,N_1632,N_1677);
or U2247 (N_2247,N_1615,N_1712);
nand U2248 (N_2248,N_1611,N_1560);
nor U2249 (N_2249,N_1647,N_1654);
nor U2250 (N_2250,N_1888,N_1612);
or U2251 (N_2251,N_1811,N_1897);
nor U2252 (N_2252,N_1703,N_1834);
nor U2253 (N_2253,N_1735,N_1687);
or U2254 (N_2254,N_1633,N_1527);
or U2255 (N_2255,N_1887,N_1654);
and U2256 (N_2256,N_1610,N_1565);
nand U2257 (N_2257,N_1855,N_1975);
nand U2258 (N_2258,N_1798,N_1581);
nand U2259 (N_2259,N_1751,N_1972);
and U2260 (N_2260,N_1697,N_1756);
or U2261 (N_2261,N_1869,N_1832);
nand U2262 (N_2262,N_1692,N_1524);
nand U2263 (N_2263,N_1921,N_1976);
xnor U2264 (N_2264,N_1642,N_1775);
or U2265 (N_2265,N_1791,N_1664);
nand U2266 (N_2266,N_1819,N_1912);
nand U2267 (N_2267,N_1703,N_1971);
and U2268 (N_2268,N_1822,N_1573);
nand U2269 (N_2269,N_1665,N_1984);
nor U2270 (N_2270,N_1761,N_1623);
nand U2271 (N_2271,N_1578,N_1812);
and U2272 (N_2272,N_1719,N_1907);
or U2273 (N_2273,N_1833,N_1784);
nor U2274 (N_2274,N_1748,N_1506);
or U2275 (N_2275,N_1794,N_1736);
or U2276 (N_2276,N_1660,N_1730);
or U2277 (N_2277,N_1589,N_1837);
nor U2278 (N_2278,N_1956,N_1780);
or U2279 (N_2279,N_1989,N_1653);
nor U2280 (N_2280,N_1670,N_1522);
and U2281 (N_2281,N_1968,N_1971);
or U2282 (N_2282,N_1501,N_1676);
nand U2283 (N_2283,N_1652,N_1672);
nor U2284 (N_2284,N_1945,N_1505);
or U2285 (N_2285,N_1732,N_1600);
nor U2286 (N_2286,N_1623,N_1905);
or U2287 (N_2287,N_1975,N_1624);
or U2288 (N_2288,N_1805,N_1938);
and U2289 (N_2289,N_1808,N_1773);
and U2290 (N_2290,N_1794,N_1534);
nor U2291 (N_2291,N_1626,N_1994);
or U2292 (N_2292,N_1822,N_1501);
nand U2293 (N_2293,N_1528,N_1784);
nor U2294 (N_2294,N_1874,N_1720);
and U2295 (N_2295,N_1528,N_1536);
nor U2296 (N_2296,N_1562,N_1839);
nand U2297 (N_2297,N_1790,N_1621);
nand U2298 (N_2298,N_1851,N_1717);
and U2299 (N_2299,N_1930,N_1692);
nand U2300 (N_2300,N_1702,N_1704);
nor U2301 (N_2301,N_1670,N_1929);
or U2302 (N_2302,N_1871,N_1820);
nand U2303 (N_2303,N_1543,N_1631);
nand U2304 (N_2304,N_1926,N_1756);
nor U2305 (N_2305,N_1764,N_1921);
nand U2306 (N_2306,N_1908,N_1846);
or U2307 (N_2307,N_1812,N_1645);
nand U2308 (N_2308,N_1913,N_1885);
or U2309 (N_2309,N_1820,N_1999);
or U2310 (N_2310,N_1763,N_1839);
nor U2311 (N_2311,N_1741,N_1668);
nor U2312 (N_2312,N_1667,N_1720);
nor U2313 (N_2313,N_1962,N_1699);
nand U2314 (N_2314,N_1928,N_1500);
and U2315 (N_2315,N_1748,N_1719);
nor U2316 (N_2316,N_1827,N_1869);
and U2317 (N_2317,N_1534,N_1831);
nor U2318 (N_2318,N_1757,N_1548);
and U2319 (N_2319,N_1544,N_1869);
nand U2320 (N_2320,N_1778,N_1566);
or U2321 (N_2321,N_1611,N_1644);
nor U2322 (N_2322,N_1646,N_1514);
or U2323 (N_2323,N_1521,N_1921);
xnor U2324 (N_2324,N_1588,N_1796);
nand U2325 (N_2325,N_1518,N_1571);
or U2326 (N_2326,N_1805,N_1781);
or U2327 (N_2327,N_1774,N_1971);
and U2328 (N_2328,N_1681,N_1678);
or U2329 (N_2329,N_1910,N_1704);
and U2330 (N_2330,N_1885,N_1636);
nor U2331 (N_2331,N_1758,N_1510);
nand U2332 (N_2332,N_1833,N_1552);
and U2333 (N_2333,N_1833,N_1823);
or U2334 (N_2334,N_1691,N_1540);
or U2335 (N_2335,N_1532,N_1517);
nand U2336 (N_2336,N_1853,N_1580);
nor U2337 (N_2337,N_1751,N_1791);
nor U2338 (N_2338,N_1903,N_1779);
or U2339 (N_2339,N_1647,N_1540);
nor U2340 (N_2340,N_1762,N_1897);
or U2341 (N_2341,N_1732,N_1655);
and U2342 (N_2342,N_1809,N_1558);
nor U2343 (N_2343,N_1996,N_1578);
or U2344 (N_2344,N_1768,N_1539);
nand U2345 (N_2345,N_1904,N_1510);
or U2346 (N_2346,N_1686,N_1623);
or U2347 (N_2347,N_1985,N_1768);
nor U2348 (N_2348,N_1938,N_1916);
or U2349 (N_2349,N_1634,N_1843);
or U2350 (N_2350,N_1860,N_1899);
or U2351 (N_2351,N_1655,N_1810);
nor U2352 (N_2352,N_1899,N_1633);
and U2353 (N_2353,N_1745,N_1834);
nand U2354 (N_2354,N_1917,N_1896);
nor U2355 (N_2355,N_1569,N_1632);
xor U2356 (N_2356,N_1733,N_1845);
nor U2357 (N_2357,N_1746,N_1570);
nor U2358 (N_2358,N_1663,N_1625);
nor U2359 (N_2359,N_1771,N_1801);
nand U2360 (N_2360,N_1837,N_1894);
nand U2361 (N_2361,N_1966,N_1860);
or U2362 (N_2362,N_1568,N_1542);
and U2363 (N_2363,N_1538,N_1505);
nand U2364 (N_2364,N_1622,N_1556);
nand U2365 (N_2365,N_1715,N_1788);
or U2366 (N_2366,N_1999,N_1991);
nor U2367 (N_2367,N_1749,N_1764);
or U2368 (N_2368,N_1664,N_1514);
and U2369 (N_2369,N_1651,N_1906);
nand U2370 (N_2370,N_1867,N_1633);
or U2371 (N_2371,N_1917,N_1530);
nor U2372 (N_2372,N_1586,N_1555);
nor U2373 (N_2373,N_1632,N_1741);
and U2374 (N_2374,N_1943,N_1655);
nor U2375 (N_2375,N_1984,N_1556);
or U2376 (N_2376,N_1992,N_1743);
nor U2377 (N_2377,N_1519,N_1805);
nand U2378 (N_2378,N_1986,N_1992);
and U2379 (N_2379,N_1927,N_1619);
nor U2380 (N_2380,N_1659,N_1572);
nor U2381 (N_2381,N_1514,N_1773);
and U2382 (N_2382,N_1744,N_1715);
and U2383 (N_2383,N_1889,N_1969);
nand U2384 (N_2384,N_1911,N_1842);
nor U2385 (N_2385,N_1856,N_1936);
nor U2386 (N_2386,N_1614,N_1882);
nand U2387 (N_2387,N_1595,N_1525);
and U2388 (N_2388,N_1722,N_1671);
nor U2389 (N_2389,N_1575,N_1776);
nor U2390 (N_2390,N_1927,N_1630);
nor U2391 (N_2391,N_1859,N_1935);
and U2392 (N_2392,N_1995,N_1652);
nor U2393 (N_2393,N_1868,N_1717);
or U2394 (N_2394,N_1526,N_1798);
nor U2395 (N_2395,N_1641,N_1707);
and U2396 (N_2396,N_1682,N_1881);
or U2397 (N_2397,N_1717,N_1543);
nand U2398 (N_2398,N_1610,N_1622);
nor U2399 (N_2399,N_1955,N_1899);
or U2400 (N_2400,N_1529,N_1708);
and U2401 (N_2401,N_1540,N_1763);
or U2402 (N_2402,N_1519,N_1721);
or U2403 (N_2403,N_1529,N_1855);
nor U2404 (N_2404,N_1900,N_1627);
nor U2405 (N_2405,N_1608,N_1662);
and U2406 (N_2406,N_1608,N_1803);
and U2407 (N_2407,N_1894,N_1758);
nand U2408 (N_2408,N_1944,N_1908);
nor U2409 (N_2409,N_1870,N_1623);
and U2410 (N_2410,N_1656,N_1862);
nand U2411 (N_2411,N_1986,N_1748);
or U2412 (N_2412,N_1917,N_1762);
nand U2413 (N_2413,N_1953,N_1631);
xnor U2414 (N_2414,N_1666,N_1692);
or U2415 (N_2415,N_1730,N_1556);
or U2416 (N_2416,N_1517,N_1668);
and U2417 (N_2417,N_1572,N_1566);
nand U2418 (N_2418,N_1547,N_1786);
nand U2419 (N_2419,N_1568,N_1799);
nand U2420 (N_2420,N_1905,N_1638);
and U2421 (N_2421,N_1600,N_1961);
xor U2422 (N_2422,N_1519,N_1666);
nand U2423 (N_2423,N_1914,N_1598);
and U2424 (N_2424,N_1542,N_1582);
and U2425 (N_2425,N_1696,N_1728);
nor U2426 (N_2426,N_1831,N_1503);
and U2427 (N_2427,N_1911,N_1922);
nor U2428 (N_2428,N_1781,N_1915);
and U2429 (N_2429,N_1694,N_1589);
and U2430 (N_2430,N_1671,N_1677);
nand U2431 (N_2431,N_1672,N_1624);
or U2432 (N_2432,N_1586,N_1724);
and U2433 (N_2433,N_1651,N_1995);
or U2434 (N_2434,N_1781,N_1874);
and U2435 (N_2435,N_1805,N_1662);
nand U2436 (N_2436,N_1543,N_1984);
nor U2437 (N_2437,N_1695,N_1581);
or U2438 (N_2438,N_1682,N_1558);
and U2439 (N_2439,N_1874,N_1998);
xor U2440 (N_2440,N_1850,N_1880);
nor U2441 (N_2441,N_1618,N_1504);
nand U2442 (N_2442,N_1564,N_1908);
nor U2443 (N_2443,N_1668,N_1545);
or U2444 (N_2444,N_1603,N_1674);
or U2445 (N_2445,N_1923,N_1863);
nor U2446 (N_2446,N_1691,N_1907);
or U2447 (N_2447,N_1692,N_1700);
or U2448 (N_2448,N_1603,N_1783);
nand U2449 (N_2449,N_1916,N_1976);
nand U2450 (N_2450,N_1767,N_1835);
and U2451 (N_2451,N_1502,N_1914);
and U2452 (N_2452,N_1680,N_1543);
and U2453 (N_2453,N_1914,N_1543);
nand U2454 (N_2454,N_1896,N_1551);
nor U2455 (N_2455,N_1647,N_1795);
nor U2456 (N_2456,N_1788,N_1664);
nor U2457 (N_2457,N_1991,N_1644);
nand U2458 (N_2458,N_1711,N_1682);
nand U2459 (N_2459,N_1664,N_1779);
nor U2460 (N_2460,N_1838,N_1731);
or U2461 (N_2461,N_1880,N_1776);
and U2462 (N_2462,N_1975,N_1960);
or U2463 (N_2463,N_1997,N_1724);
nand U2464 (N_2464,N_1635,N_1691);
and U2465 (N_2465,N_1511,N_1951);
and U2466 (N_2466,N_1611,N_1528);
nor U2467 (N_2467,N_1756,N_1569);
nor U2468 (N_2468,N_1628,N_1690);
nand U2469 (N_2469,N_1698,N_1931);
nand U2470 (N_2470,N_1766,N_1593);
or U2471 (N_2471,N_1777,N_1721);
xor U2472 (N_2472,N_1627,N_1504);
and U2473 (N_2473,N_1506,N_1526);
nand U2474 (N_2474,N_1821,N_1988);
or U2475 (N_2475,N_1729,N_1897);
xor U2476 (N_2476,N_1918,N_1947);
or U2477 (N_2477,N_1561,N_1669);
and U2478 (N_2478,N_1613,N_1527);
nor U2479 (N_2479,N_1747,N_1569);
nand U2480 (N_2480,N_1556,N_1990);
or U2481 (N_2481,N_1944,N_1625);
nand U2482 (N_2482,N_1717,N_1830);
or U2483 (N_2483,N_1708,N_1795);
xor U2484 (N_2484,N_1726,N_1854);
nand U2485 (N_2485,N_1921,N_1837);
and U2486 (N_2486,N_1752,N_1831);
or U2487 (N_2487,N_1622,N_1712);
or U2488 (N_2488,N_1619,N_1502);
nor U2489 (N_2489,N_1788,N_1820);
nand U2490 (N_2490,N_1586,N_1503);
nand U2491 (N_2491,N_1736,N_1840);
nand U2492 (N_2492,N_1899,N_1697);
or U2493 (N_2493,N_1926,N_1578);
or U2494 (N_2494,N_1933,N_1880);
or U2495 (N_2495,N_1706,N_1700);
and U2496 (N_2496,N_1755,N_1783);
nor U2497 (N_2497,N_1607,N_1865);
nand U2498 (N_2498,N_1945,N_1528);
nand U2499 (N_2499,N_1906,N_1853);
nand U2500 (N_2500,N_2051,N_2141);
and U2501 (N_2501,N_2113,N_2292);
or U2502 (N_2502,N_2247,N_2120);
nand U2503 (N_2503,N_2361,N_2265);
or U2504 (N_2504,N_2284,N_2432);
nand U2505 (N_2505,N_2473,N_2032);
nor U2506 (N_2506,N_2167,N_2068);
nand U2507 (N_2507,N_2045,N_2468);
nor U2508 (N_2508,N_2023,N_2406);
nor U2509 (N_2509,N_2036,N_2460);
nor U2510 (N_2510,N_2208,N_2298);
nand U2511 (N_2511,N_2271,N_2211);
or U2512 (N_2512,N_2417,N_2127);
xor U2513 (N_2513,N_2356,N_2479);
nor U2514 (N_2514,N_2395,N_2379);
nand U2515 (N_2515,N_2267,N_2179);
nand U2516 (N_2516,N_2001,N_2454);
or U2517 (N_2517,N_2092,N_2290);
or U2518 (N_2518,N_2198,N_2436);
nor U2519 (N_2519,N_2178,N_2297);
nand U2520 (N_2520,N_2386,N_2106);
nor U2521 (N_2521,N_2035,N_2328);
nand U2522 (N_2522,N_2121,N_2004);
and U2523 (N_2523,N_2329,N_2472);
nand U2524 (N_2524,N_2133,N_2316);
nand U2525 (N_2525,N_2124,N_2230);
nor U2526 (N_2526,N_2273,N_2084);
and U2527 (N_2527,N_2170,N_2233);
and U2528 (N_2528,N_2214,N_2094);
nand U2529 (N_2529,N_2061,N_2163);
and U2530 (N_2530,N_2040,N_2189);
nand U2531 (N_2531,N_2197,N_2082);
or U2532 (N_2532,N_2222,N_2087);
and U2533 (N_2533,N_2209,N_2097);
nor U2534 (N_2534,N_2168,N_2025);
nand U2535 (N_2535,N_2042,N_2227);
nor U2536 (N_2536,N_2487,N_2365);
and U2537 (N_2537,N_2080,N_2058);
nor U2538 (N_2538,N_2412,N_2358);
nand U2539 (N_2539,N_2370,N_2494);
nand U2540 (N_2540,N_2264,N_2414);
nand U2541 (N_2541,N_2413,N_2394);
nand U2542 (N_2542,N_2321,N_2186);
and U2543 (N_2543,N_2334,N_2043);
or U2544 (N_2544,N_2218,N_2176);
and U2545 (N_2545,N_2044,N_2085);
and U2546 (N_2546,N_2174,N_2215);
and U2547 (N_2547,N_2266,N_2449);
or U2548 (N_2548,N_2399,N_2232);
or U2549 (N_2549,N_2072,N_2115);
nor U2550 (N_2550,N_2439,N_2246);
and U2551 (N_2551,N_2341,N_2461);
and U2552 (N_2552,N_2095,N_2389);
or U2553 (N_2553,N_2342,N_2303);
nand U2554 (N_2554,N_2162,N_2295);
or U2555 (N_2555,N_2305,N_2301);
and U2556 (N_2556,N_2136,N_2360);
and U2557 (N_2557,N_2482,N_2257);
nor U2558 (N_2558,N_2228,N_2005);
nand U2559 (N_2559,N_2003,N_2201);
or U2560 (N_2560,N_2135,N_2242);
nor U2561 (N_2561,N_2028,N_2492);
or U2562 (N_2562,N_2418,N_2076);
nand U2563 (N_2563,N_2021,N_2407);
nand U2564 (N_2564,N_2263,N_2485);
and U2565 (N_2565,N_2445,N_2156);
nor U2566 (N_2566,N_2011,N_2309);
nor U2567 (N_2567,N_2338,N_2054);
nor U2568 (N_2568,N_2333,N_2427);
nand U2569 (N_2569,N_2426,N_2304);
nor U2570 (N_2570,N_2364,N_2355);
nor U2571 (N_2571,N_2374,N_2375);
and U2572 (N_2572,N_2446,N_2307);
nor U2573 (N_2573,N_2107,N_2249);
or U2574 (N_2574,N_2421,N_2038);
and U2575 (N_2575,N_2433,N_2016);
nor U2576 (N_2576,N_2039,N_2311);
nor U2577 (N_2577,N_2289,N_2410);
and U2578 (N_2578,N_2172,N_2149);
nand U2579 (N_2579,N_2455,N_2363);
nor U2580 (N_2580,N_2238,N_2404);
or U2581 (N_2581,N_2254,N_2026);
or U2582 (N_2582,N_2420,N_2274);
nand U2583 (N_2583,N_2102,N_2148);
nor U2584 (N_2584,N_2474,N_2291);
xor U2585 (N_2585,N_2069,N_2437);
nand U2586 (N_2586,N_2348,N_2315);
nor U2587 (N_2587,N_2319,N_2392);
nor U2588 (N_2588,N_2422,N_2486);
nand U2589 (N_2589,N_2125,N_2020);
or U2590 (N_2590,N_2116,N_2447);
and U2591 (N_2591,N_2203,N_2337);
or U2592 (N_2592,N_2497,N_2223);
nand U2593 (N_2593,N_2184,N_2411);
nor U2594 (N_2594,N_2287,N_2047);
nor U2595 (N_2595,N_2111,N_2123);
or U2596 (N_2596,N_2405,N_2083);
nand U2597 (N_2597,N_2268,N_2217);
nand U2598 (N_2598,N_2464,N_2381);
and U2599 (N_2599,N_2450,N_2160);
or U2600 (N_2600,N_2213,N_2330);
nor U2601 (N_2601,N_2367,N_2430);
or U2602 (N_2602,N_2112,N_2452);
and U2603 (N_2603,N_2091,N_2165);
and U2604 (N_2604,N_2014,N_2368);
nor U2605 (N_2605,N_2402,N_2489);
xnor U2606 (N_2606,N_2182,N_2006);
and U2607 (N_2607,N_2324,N_2100);
or U2608 (N_2608,N_2296,N_2423);
nor U2609 (N_2609,N_2434,N_2164);
nor U2610 (N_2610,N_2057,N_2340);
nand U2611 (N_2611,N_2226,N_2105);
or U2612 (N_2612,N_2088,N_2109);
xnor U2613 (N_2613,N_2459,N_2477);
and U2614 (N_2614,N_2187,N_2012);
nor U2615 (N_2615,N_2188,N_2318);
or U2616 (N_2616,N_2033,N_2140);
or U2617 (N_2617,N_2219,N_2308);
nand U2618 (N_2618,N_2387,N_2017);
and U2619 (N_2619,N_2326,N_2131);
nor U2620 (N_2620,N_2431,N_2438);
or U2621 (N_2621,N_2099,N_2066);
xor U2622 (N_2622,N_2441,N_2101);
nand U2623 (N_2623,N_2074,N_2122);
nand U2624 (N_2624,N_2052,N_2031);
nand U2625 (N_2625,N_2384,N_2269);
or U2626 (N_2626,N_2442,N_2322);
nand U2627 (N_2627,N_2331,N_2185);
nor U2628 (N_2628,N_2344,N_2060);
nand U2629 (N_2629,N_2081,N_2484);
nand U2630 (N_2630,N_2142,N_2152);
or U2631 (N_2631,N_2067,N_2428);
or U2632 (N_2632,N_2171,N_2018);
nand U2633 (N_2633,N_2096,N_2471);
or U2634 (N_2634,N_2192,N_2312);
nor U2635 (N_2635,N_2408,N_2002);
nor U2636 (N_2636,N_2065,N_2498);
and U2637 (N_2637,N_2053,N_2138);
nor U2638 (N_2638,N_2030,N_2119);
and U2639 (N_2639,N_2396,N_2177);
or U2640 (N_2640,N_2098,N_2354);
and U2641 (N_2641,N_2481,N_2332);
or U2642 (N_2642,N_2229,N_2378);
nand U2643 (N_2643,N_2008,N_2104);
or U2644 (N_2644,N_2466,N_2173);
nor U2645 (N_2645,N_2346,N_2458);
or U2646 (N_2646,N_2078,N_2251);
or U2647 (N_2647,N_2118,N_2357);
nor U2648 (N_2648,N_2110,N_2415);
and U2649 (N_2649,N_2280,N_2161);
nor U2650 (N_2650,N_2306,N_2429);
nor U2651 (N_2651,N_2159,N_2241);
and U2652 (N_2652,N_2327,N_2493);
or U2653 (N_2653,N_2245,N_2248);
or U2654 (N_2654,N_2169,N_2335);
or U2655 (N_2655,N_2055,N_2224);
and U2656 (N_2656,N_2108,N_2050);
nand U2657 (N_2657,N_2270,N_2191);
or U2658 (N_2658,N_2231,N_2202);
or U2659 (N_2659,N_2444,N_2352);
nor U2660 (N_2660,N_2300,N_2345);
nand U2661 (N_2661,N_2279,N_2443);
nor U2662 (N_2662,N_2147,N_2313);
and U2663 (N_2663,N_2288,N_2259);
nand U2664 (N_2664,N_2491,N_2073);
nor U2665 (N_2665,N_2323,N_2480);
nor U2666 (N_2666,N_2193,N_2007);
xnor U2667 (N_2667,N_2180,N_2234);
and U2668 (N_2668,N_2139,N_2158);
nor U2669 (N_2669,N_2151,N_2393);
nor U2670 (N_2670,N_2293,N_2130);
nor U2671 (N_2671,N_2250,N_2390);
nand U2672 (N_2672,N_2022,N_2310);
and U2673 (N_2673,N_2143,N_2350);
nor U2674 (N_2674,N_2144,N_2062);
and U2675 (N_2675,N_2013,N_2325);
and U2676 (N_2676,N_2194,N_2093);
and U2677 (N_2677,N_2294,N_2244);
or U2678 (N_2678,N_2046,N_2283);
nor U2679 (N_2679,N_2478,N_2369);
nand U2680 (N_2680,N_2220,N_2451);
nand U2681 (N_2681,N_2200,N_2282);
and U2682 (N_2682,N_2440,N_2351);
nor U2683 (N_2683,N_2488,N_2196);
nand U2684 (N_2684,N_2373,N_2145);
and U2685 (N_2685,N_2153,N_2388);
or U2686 (N_2686,N_2475,N_2339);
nor U2687 (N_2687,N_2103,N_2225);
nand U2688 (N_2688,N_2400,N_2463);
and U2689 (N_2689,N_2070,N_2401);
and U2690 (N_2690,N_2314,N_2077);
nor U2691 (N_2691,N_2041,N_2383);
nor U2692 (N_2692,N_2009,N_2255);
and U2693 (N_2693,N_2336,N_2237);
or U2694 (N_2694,N_2372,N_2240);
or U2695 (N_2695,N_2207,N_2079);
nand U2696 (N_2696,N_2275,N_2272);
and U2697 (N_2697,N_2382,N_2114);
and U2698 (N_2698,N_2256,N_2126);
nand U2699 (N_2699,N_2490,N_2260);
nor U2700 (N_2700,N_2048,N_2376);
nor U2701 (N_2701,N_2470,N_2398);
nand U2702 (N_2702,N_2469,N_2128);
or U2703 (N_2703,N_2075,N_2166);
or U2704 (N_2704,N_2302,N_2276);
nand U2705 (N_2705,N_2063,N_2037);
nand U2706 (N_2706,N_2391,N_2448);
or U2707 (N_2707,N_2495,N_2216);
nor U2708 (N_2708,N_2086,N_2467);
or U2709 (N_2709,N_2132,N_2347);
nor U2710 (N_2710,N_2146,N_2258);
or U2711 (N_2711,N_2236,N_2221);
and U2712 (N_2712,N_2397,N_2155);
nand U2713 (N_2713,N_2317,N_2015);
and U2714 (N_2714,N_2137,N_2261);
or U2715 (N_2715,N_2253,N_2286);
nand U2716 (N_2716,N_2195,N_2034);
or U2717 (N_2717,N_2154,N_2206);
nor U2718 (N_2718,N_2496,N_2019);
or U2719 (N_2719,N_2134,N_2157);
and U2720 (N_2720,N_2349,N_2150);
nor U2721 (N_2721,N_2380,N_2205);
nor U2722 (N_2722,N_2252,N_2049);
and U2723 (N_2723,N_2385,N_2210);
nor U2724 (N_2724,N_2343,N_2281);
and U2725 (N_2725,N_2435,N_2320);
xnor U2726 (N_2726,N_2371,N_2059);
or U2727 (N_2727,N_2056,N_2064);
nand U2728 (N_2728,N_2262,N_2366);
and U2729 (N_2729,N_2359,N_2483);
nor U2730 (N_2730,N_2353,N_2000);
and U2731 (N_2731,N_2403,N_2377);
nor U2732 (N_2732,N_2476,N_2029);
nand U2733 (N_2733,N_2285,N_2277);
nand U2734 (N_2734,N_2278,N_2010);
nand U2735 (N_2735,N_2199,N_2419);
nand U2736 (N_2736,N_2425,N_2027);
or U2737 (N_2737,N_2462,N_2465);
nand U2738 (N_2738,N_2299,N_2457);
and U2739 (N_2739,N_2235,N_2090);
and U2740 (N_2740,N_2409,N_2499);
or U2741 (N_2741,N_2117,N_2212);
and U2742 (N_2742,N_2071,N_2181);
and U2743 (N_2743,N_2453,N_2456);
nor U2744 (N_2744,N_2024,N_2416);
or U2745 (N_2745,N_2183,N_2175);
and U2746 (N_2746,N_2362,N_2190);
or U2747 (N_2747,N_2129,N_2243);
and U2748 (N_2748,N_2089,N_2424);
nand U2749 (N_2749,N_2239,N_2204);
or U2750 (N_2750,N_2049,N_2145);
nor U2751 (N_2751,N_2158,N_2250);
or U2752 (N_2752,N_2158,N_2071);
and U2753 (N_2753,N_2058,N_2426);
nor U2754 (N_2754,N_2054,N_2378);
nand U2755 (N_2755,N_2175,N_2297);
and U2756 (N_2756,N_2327,N_2478);
nand U2757 (N_2757,N_2034,N_2340);
and U2758 (N_2758,N_2465,N_2377);
and U2759 (N_2759,N_2391,N_2437);
nand U2760 (N_2760,N_2083,N_2181);
or U2761 (N_2761,N_2344,N_2497);
nand U2762 (N_2762,N_2150,N_2388);
and U2763 (N_2763,N_2491,N_2093);
nand U2764 (N_2764,N_2335,N_2475);
or U2765 (N_2765,N_2074,N_2111);
or U2766 (N_2766,N_2346,N_2358);
or U2767 (N_2767,N_2222,N_2290);
or U2768 (N_2768,N_2355,N_2260);
nor U2769 (N_2769,N_2436,N_2199);
nor U2770 (N_2770,N_2030,N_2342);
or U2771 (N_2771,N_2258,N_2058);
and U2772 (N_2772,N_2388,N_2172);
nor U2773 (N_2773,N_2177,N_2085);
xnor U2774 (N_2774,N_2071,N_2210);
or U2775 (N_2775,N_2174,N_2447);
nand U2776 (N_2776,N_2499,N_2201);
nand U2777 (N_2777,N_2219,N_2314);
nand U2778 (N_2778,N_2028,N_2493);
and U2779 (N_2779,N_2010,N_2371);
or U2780 (N_2780,N_2073,N_2309);
nor U2781 (N_2781,N_2200,N_2141);
and U2782 (N_2782,N_2246,N_2278);
and U2783 (N_2783,N_2187,N_2019);
nor U2784 (N_2784,N_2228,N_2178);
nand U2785 (N_2785,N_2298,N_2318);
and U2786 (N_2786,N_2360,N_2003);
or U2787 (N_2787,N_2307,N_2414);
nor U2788 (N_2788,N_2121,N_2352);
or U2789 (N_2789,N_2320,N_2119);
nand U2790 (N_2790,N_2400,N_2107);
and U2791 (N_2791,N_2116,N_2203);
or U2792 (N_2792,N_2113,N_2373);
nand U2793 (N_2793,N_2421,N_2160);
or U2794 (N_2794,N_2240,N_2050);
nor U2795 (N_2795,N_2303,N_2318);
nor U2796 (N_2796,N_2349,N_2295);
and U2797 (N_2797,N_2332,N_2174);
nand U2798 (N_2798,N_2436,N_2274);
or U2799 (N_2799,N_2426,N_2344);
and U2800 (N_2800,N_2424,N_2061);
nand U2801 (N_2801,N_2164,N_2216);
or U2802 (N_2802,N_2009,N_2203);
or U2803 (N_2803,N_2186,N_2228);
nand U2804 (N_2804,N_2124,N_2028);
nor U2805 (N_2805,N_2082,N_2130);
and U2806 (N_2806,N_2205,N_2239);
nor U2807 (N_2807,N_2103,N_2230);
nand U2808 (N_2808,N_2015,N_2160);
and U2809 (N_2809,N_2343,N_2108);
nor U2810 (N_2810,N_2171,N_2236);
nor U2811 (N_2811,N_2251,N_2240);
nor U2812 (N_2812,N_2339,N_2471);
nand U2813 (N_2813,N_2043,N_2186);
or U2814 (N_2814,N_2178,N_2315);
and U2815 (N_2815,N_2284,N_2116);
nor U2816 (N_2816,N_2319,N_2089);
or U2817 (N_2817,N_2162,N_2170);
nand U2818 (N_2818,N_2031,N_2180);
and U2819 (N_2819,N_2451,N_2108);
nor U2820 (N_2820,N_2264,N_2228);
nand U2821 (N_2821,N_2220,N_2437);
and U2822 (N_2822,N_2077,N_2310);
xnor U2823 (N_2823,N_2096,N_2338);
nand U2824 (N_2824,N_2447,N_2056);
or U2825 (N_2825,N_2319,N_2149);
nand U2826 (N_2826,N_2105,N_2316);
and U2827 (N_2827,N_2080,N_2051);
and U2828 (N_2828,N_2151,N_2274);
nand U2829 (N_2829,N_2061,N_2181);
nand U2830 (N_2830,N_2405,N_2070);
nor U2831 (N_2831,N_2413,N_2223);
nor U2832 (N_2832,N_2321,N_2306);
or U2833 (N_2833,N_2305,N_2231);
nor U2834 (N_2834,N_2445,N_2292);
or U2835 (N_2835,N_2467,N_2354);
nand U2836 (N_2836,N_2336,N_2212);
or U2837 (N_2837,N_2323,N_2109);
nor U2838 (N_2838,N_2248,N_2077);
nand U2839 (N_2839,N_2271,N_2220);
and U2840 (N_2840,N_2011,N_2281);
or U2841 (N_2841,N_2401,N_2487);
or U2842 (N_2842,N_2221,N_2375);
nor U2843 (N_2843,N_2139,N_2330);
and U2844 (N_2844,N_2320,N_2052);
and U2845 (N_2845,N_2106,N_2148);
or U2846 (N_2846,N_2398,N_2433);
nand U2847 (N_2847,N_2106,N_2020);
and U2848 (N_2848,N_2297,N_2197);
nor U2849 (N_2849,N_2383,N_2038);
or U2850 (N_2850,N_2331,N_2377);
or U2851 (N_2851,N_2120,N_2056);
nor U2852 (N_2852,N_2235,N_2092);
and U2853 (N_2853,N_2494,N_2402);
or U2854 (N_2854,N_2415,N_2185);
nor U2855 (N_2855,N_2407,N_2113);
or U2856 (N_2856,N_2090,N_2468);
and U2857 (N_2857,N_2067,N_2025);
nor U2858 (N_2858,N_2280,N_2303);
nor U2859 (N_2859,N_2334,N_2154);
and U2860 (N_2860,N_2103,N_2070);
nor U2861 (N_2861,N_2102,N_2115);
and U2862 (N_2862,N_2313,N_2344);
and U2863 (N_2863,N_2384,N_2362);
or U2864 (N_2864,N_2170,N_2294);
nor U2865 (N_2865,N_2311,N_2397);
nand U2866 (N_2866,N_2115,N_2235);
or U2867 (N_2867,N_2330,N_2086);
nand U2868 (N_2868,N_2331,N_2188);
nand U2869 (N_2869,N_2340,N_2262);
nand U2870 (N_2870,N_2368,N_2180);
and U2871 (N_2871,N_2268,N_2123);
nor U2872 (N_2872,N_2408,N_2182);
nand U2873 (N_2873,N_2241,N_2383);
nand U2874 (N_2874,N_2179,N_2460);
nor U2875 (N_2875,N_2447,N_2439);
nor U2876 (N_2876,N_2050,N_2098);
and U2877 (N_2877,N_2154,N_2172);
nand U2878 (N_2878,N_2487,N_2097);
nand U2879 (N_2879,N_2431,N_2239);
nor U2880 (N_2880,N_2423,N_2164);
and U2881 (N_2881,N_2298,N_2034);
or U2882 (N_2882,N_2313,N_2436);
nand U2883 (N_2883,N_2354,N_2471);
and U2884 (N_2884,N_2474,N_2114);
nand U2885 (N_2885,N_2444,N_2057);
nor U2886 (N_2886,N_2470,N_2142);
and U2887 (N_2887,N_2376,N_2446);
or U2888 (N_2888,N_2262,N_2445);
nor U2889 (N_2889,N_2495,N_2092);
or U2890 (N_2890,N_2025,N_2343);
nand U2891 (N_2891,N_2325,N_2493);
nand U2892 (N_2892,N_2381,N_2451);
and U2893 (N_2893,N_2281,N_2120);
and U2894 (N_2894,N_2159,N_2398);
or U2895 (N_2895,N_2006,N_2453);
nor U2896 (N_2896,N_2272,N_2109);
or U2897 (N_2897,N_2416,N_2336);
and U2898 (N_2898,N_2058,N_2133);
nor U2899 (N_2899,N_2382,N_2375);
or U2900 (N_2900,N_2481,N_2354);
and U2901 (N_2901,N_2491,N_2191);
and U2902 (N_2902,N_2260,N_2414);
or U2903 (N_2903,N_2373,N_2166);
or U2904 (N_2904,N_2193,N_2403);
nand U2905 (N_2905,N_2114,N_2237);
nand U2906 (N_2906,N_2022,N_2441);
nor U2907 (N_2907,N_2320,N_2041);
nor U2908 (N_2908,N_2271,N_2053);
and U2909 (N_2909,N_2459,N_2398);
and U2910 (N_2910,N_2296,N_2257);
and U2911 (N_2911,N_2285,N_2299);
nand U2912 (N_2912,N_2081,N_2053);
nand U2913 (N_2913,N_2149,N_2211);
nand U2914 (N_2914,N_2453,N_2319);
nand U2915 (N_2915,N_2486,N_2400);
nor U2916 (N_2916,N_2242,N_2124);
nor U2917 (N_2917,N_2225,N_2167);
and U2918 (N_2918,N_2405,N_2343);
nand U2919 (N_2919,N_2340,N_2137);
nor U2920 (N_2920,N_2112,N_2039);
nor U2921 (N_2921,N_2073,N_2494);
nor U2922 (N_2922,N_2081,N_2283);
and U2923 (N_2923,N_2160,N_2385);
or U2924 (N_2924,N_2260,N_2020);
or U2925 (N_2925,N_2342,N_2212);
or U2926 (N_2926,N_2003,N_2446);
nor U2927 (N_2927,N_2465,N_2353);
nand U2928 (N_2928,N_2250,N_2097);
xor U2929 (N_2929,N_2327,N_2424);
and U2930 (N_2930,N_2155,N_2137);
nand U2931 (N_2931,N_2430,N_2145);
nand U2932 (N_2932,N_2227,N_2226);
and U2933 (N_2933,N_2477,N_2331);
nor U2934 (N_2934,N_2492,N_2171);
nand U2935 (N_2935,N_2095,N_2384);
nand U2936 (N_2936,N_2292,N_2092);
and U2937 (N_2937,N_2120,N_2302);
nor U2938 (N_2938,N_2066,N_2481);
or U2939 (N_2939,N_2261,N_2272);
nand U2940 (N_2940,N_2185,N_2269);
nor U2941 (N_2941,N_2456,N_2151);
nand U2942 (N_2942,N_2303,N_2284);
or U2943 (N_2943,N_2488,N_2132);
nor U2944 (N_2944,N_2333,N_2399);
nand U2945 (N_2945,N_2056,N_2274);
nor U2946 (N_2946,N_2246,N_2372);
or U2947 (N_2947,N_2158,N_2408);
or U2948 (N_2948,N_2159,N_2074);
nand U2949 (N_2949,N_2220,N_2174);
and U2950 (N_2950,N_2177,N_2033);
nand U2951 (N_2951,N_2254,N_2261);
nand U2952 (N_2952,N_2279,N_2055);
nand U2953 (N_2953,N_2483,N_2394);
nand U2954 (N_2954,N_2450,N_2308);
or U2955 (N_2955,N_2339,N_2057);
or U2956 (N_2956,N_2242,N_2136);
or U2957 (N_2957,N_2214,N_2228);
nand U2958 (N_2958,N_2095,N_2240);
nand U2959 (N_2959,N_2006,N_2069);
nand U2960 (N_2960,N_2495,N_2441);
xnor U2961 (N_2961,N_2207,N_2039);
nand U2962 (N_2962,N_2072,N_2288);
nor U2963 (N_2963,N_2045,N_2259);
and U2964 (N_2964,N_2142,N_2350);
and U2965 (N_2965,N_2450,N_2327);
and U2966 (N_2966,N_2086,N_2473);
nor U2967 (N_2967,N_2288,N_2457);
or U2968 (N_2968,N_2385,N_2353);
or U2969 (N_2969,N_2228,N_2472);
or U2970 (N_2970,N_2054,N_2301);
or U2971 (N_2971,N_2153,N_2451);
or U2972 (N_2972,N_2240,N_2309);
nor U2973 (N_2973,N_2444,N_2079);
and U2974 (N_2974,N_2466,N_2487);
nor U2975 (N_2975,N_2001,N_2400);
and U2976 (N_2976,N_2456,N_2489);
nand U2977 (N_2977,N_2022,N_2243);
nor U2978 (N_2978,N_2353,N_2424);
and U2979 (N_2979,N_2379,N_2274);
or U2980 (N_2980,N_2448,N_2103);
or U2981 (N_2981,N_2115,N_2030);
nand U2982 (N_2982,N_2207,N_2259);
and U2983 (N_2983,N_2295,N_2256);
nor U2984 (N_2984,N_2396,N_2337);
and U2985 (N_2985,N_2011,N_2411);
nand U2986 (N_2986,N_2156,N_2029);
and U2987 (N_2987,N_2179,N_2091);
nand U2988 (N_2988,N_2468,N_2145);
and U2989 (N_2989,N_2166,N_2396);
or U2990 (N_2990,N_2085,N_2126);
nand U2991 (N_2991,N_2341,N_2176);
nor U2992 (N_2992,N_2103,N_2013);
or U2993 (N_2993,N_2122,N_2131);
or U2994 (N_2994,N_2167,N_2276);
nand U2995 (N_2995,N_2451,N_2391);
nand U2996 (N_2996,N_2270,N_2396);
nand U2997 (N_2997,N_2320,N_2266);
nand U2998 (N_2998,N_2150,N_2325);
and U2999 (N_2999,N_2323,N_2219);
and U3000 (N_3000,N_2983,N_2849);
nand U3001 (N_3001,N_2953,N_2800);
or U3002 (N_3002,N_2592,N_2927);
nand U3003 (N_3003,N_2694,N_2510);
nor U3004 (N_3004,N_2935,N_2790);
or U3005 (N_3005,N_2956,N_2746);
or U3006 (N_3006,N_2518,N_2699);
or U3007 (N_3007,N_2507,N_2855);
nand U3008 (N_3008,N_2614,N_2812);
or U3009 (N_3009,N_2639,N_2880);
nor U3010 (N_3010,N_2512,N_2535);
and U3011 (N_3011,N_2958,N_2545);
or U3012 (N_3012,N_2587,N_2965);
nand U3013 (N_3013,N_2934,N_2649);
nand U3014 (N_3014,N_2827,N_2964);
and U3015 (N_3015,N_2750,N_2659);
nor U3016 (N_3016,N_2591,N_2967);
nand U3017 (N_3017,N_2796,N_2763);
nor U3018 (N_3018,N_2868,N_2735);
or U3019 (N_3019,N_2787,N_2807);
and U3020 (N_3020,N_2685,N_2679);
and U3021 (N_3021,N_2904,N_2543);
or U3022 (N_3022,N_2624,N_2665);
nand U3023 (N_3023,N_2526,N_2889);
or U3024 (N_3024,N_2742,N_2814);
and U3025 (N_3025,N_2896,N_2806);
or U3026 (N_3026,N_2505,N_2982);
or U3027 (N_3027,N_2860,N_2627);
or U3028 (N_3028,N_2762,N_2723);
and U3029 (N_3029,N_2539,N_2662);
nor U3030 (N_3030,N_2852,N_2745);
nor U3031 (N_3031,N_2758,N_2845);
nand U3032 (N_3032,N_2566,N_2701);
and U3033 (N_3033,N_2950,N_2754);
or U3034 (N_3034,N_2756,N_2932);
and U3035 (N_3035,N_2985,N_2791);
nor U3036 (N_3036,N_2987,N_2912);
and U3037 (N_3037,N_2644,N_2603);
nor U3038 (N_3038,N_2672,N_2997);
or U3039 (N_3039,N_2640,N_2653);
or U3040 (N_3040,N_2940,N_2892);
or U3041 (N_3041,N_2559,N_2586);
nor U3042 (N_3042,N_2669,N_2631);
nor U3043 (N_3043,N_2575,N_2552);
nand U3044 (N_3044,N_2719,N_2870);
nand U3045 (N_3045,N_2712,N_2817);
or U3046 (N_3046,N_2700,N_2891);
nor U3047 (N_3047,N_2897,N_2576);
or U3048 (N_3048,N_2560,N_2609);
or U3049 (N_3049,N_2504,N_2532);
nand U3050 (N_3050,N_2764,N_2687);
nand U3051 (N_3051,N_2972,N_2671);
or U3052 (N_3052,N_2689,N_2995);
nor U3053 (N_3053,N_2973,N_2678);
nand U3054 (N_3054,N_2563,N_2548);
or U3055 (N_3055,N_2819,N_2970);
nand U3056 (N_3056,N_2741,N_2946);
or U3057 (N_3057,N_2632,N_2770);
and U3058 (N_3058,N_2585,N_2838);
and U3059 (N_3059,N_2936,N_2625);
nand U3060 (N_3060,N_2966,N_2692);
and U3061 (N_3061,N_2590,N_2593);
nor U3062 (N_3062,N_2710,N_2668);
and U3063 (N_3063,N_2841,N_2979);
or U3064 (N_3064,N_2894,N_2840);
nand U3065 (N_3065,N_2984,N_2820);
nor U3066 (N_3066,N_2582,N_2988);
and U3067 (N_3067,N_2651,N_2833);
and U3068 (N_3068,N_2907,N_2724);
and U3069 (N_3069,N_2879,N_2867);
or U3070 (N_3070,N_2739,N_2551);
nor U3071 (N_3071,N_2768,N_2565);
nor U3072 (N_3072,N_2989,N_2620);
nand U3073 (N_3073,N_2813,N_2610);
nor U3074 (N_3074,N_2788,N_2866);
or U3075 (N_3075,N_2957,N_2853);
or U3076 (N_3076,N_2748,N_2971);
and U3077 (N_3077,N_2622,N_2772);
nor U3078 (N_3078,N_2513,N_2830);
or U3079 (N_3079,N_2882,N_2584);
nor U3080 (N_3080,N_2781,N_2914);
nand U3081 (N_3081,N_2617,N_2899);
and U3082 (N_3082,N_2562,N_2888);
or U3083 (N_3083,N_2643,N_2977);
nand U3084 (N_3084,N_2789,N_2976);
or U3085 (N_3085,N_2792,N_2616);
nor U3086 (N_3086,N_2637,N_2721);
nand U3087 (N_3087,N_2878,N_2893);
nand U3088 (N_3088,N_2810,N_2686);
nand U3089 (N_3089,N_2842,N_2900);
and U3090 (N_3090,N_2760,N_2567);
nand U3091 (N_3091,N_2655,N_2947);
nand U3092 (N_3092,N_2991,N_2994);
and U3093 (N_3093,N_2844,N_2980);
nand U3094 (N_3094,N_2529,N_2978);
or U3095 (N_3095,N_2629,N_2874);
nor U3096 (N_3096,N_2804,N_2647);
and U3097 (N_3097,N_2704,N_2909);
nor U3098 (N_3098,N_2732,N_2531);
or U3099 (N_3099,N_2933,N_2795);
and U3100 (N_3100,N_2917,N_2915);
or U3101 (N_3101,N_2524,N_2523);
or U3102 (N_3102,N_2646,N_2831);
or U3103 (N_3103,N_2717,N_2902);
and U3104 (N_3104,N_2501,N_2670);
and U3105 (N_3105,N_2581,N_2780);
and U3106 (N_3106,N_2821,N_2619);
nand U3107 (N_3107,N_2778,N_2805);
or U3108 (N_3108,N_2691,N_2534);
or U3109 (N_3109,N_2895,N_2937);
nand U3110 (N_3110,N_2736,N_2568);
and U3111 (N_3111,N_2744,N_2816);
nand U3112 (N_3112,N_2733,N_2919);
nand U3113 (N_3113,N_2588,N_2943);
nor U3114 (N_3114,N_2579,N_2537);
or U3115 (N_3115,N_2873,N_2863);
and U3116 (N_3116,N_2607,N_2515);
nand U3117 (N_3117,N_2839,N_2901);
nor U3118 (N_3118,N_2544,N_2595);
and U3119 (N_3119,N_2922,N_2598);
or U3120 (N_3120,N_2924,N_2986);
or U3121 (N_3121,N_2589,N_2858);
and U3122 (N_3122,N_2837,N_2695);
nand U3123 (N_3123,N_2635,N_2711);
and U3124 (N_3124,N_2561,N_2541);
or U3125 (N_3125,N_2641,N_2705);
nor U3126 (N_3126,N_2520,N_2801);
or U3127 (N_3127,N_2911,N_2884);
or U3128 (N_3128,N_2527,N_2533);
or U3129 (N_3129,N_2675,N_2749);
or U3130 (N_3130,N_2784,N_2573);
or U3131 (N_3131,N_2734,N_2621);
nand U3132 (N_3132,N_2612,N_2886);
nand U3133 (N_3133,N_2572,N_2877);
nand U3134 (N_3134,N_2753,N_2508);
nand U3135 (N_3135,N_2954,N_2913);
and U3136 (N_3136,N_2777,N_2664);
or U3137 (N_3137,N_2803,N_2769);
nor U3138 (N_3138,N_2557,N_2822);
nand U3139 (N_3139,N_2615,N_2570);
nor U3140 (N_3140,N_2611,N_2890);
nor U3141 (N_3141,N_2887,N_2826);
nor U3142 (N_3142,N_2981,N_2680);
or U3143 (N_3143,N_2514,N_2857);
nand U3144 (N_3144,N_2709,N_2864);
nor U3145 (N_3145,N_2843,N_2952);
nor U3146 (N_3146,N_2536,N_2525);
or U3147 (N_3147,N_2725,N_2799);
nand U3148 (N_3148,N_2761,N_2702);
nand U3149 (N_3149,N_2517,N_2809);
xor U3150 (N_3150,N_2785,N_2628);
nand U3151 (N_3151,N_2693,N_2715);
or U3152 (N_3152,N_2776,N_2553);
or U3153 (N_3153,N_2930,N_2941);
and U3154 (N_3154,N_2522,N_2728);
nand U3155 (N_3155,N_2706,N_2881);
nand U3156 (N_3156,N_2650,N_2757);
or U3157 (N_3157,N_2682,N_2818);
or U3158 (N_3158,N_2794,N_2920);
nand U3159 (N_3159,N_2564,N_2752);
nand U3160 (N_3160,N_2835,N_2856);
or U3161 (N_3161,N_2727,N_2638);
nand U3162 (N_3162,N_2908,N_2848);
nand U3163 (N_3163,N_2751,N_2718);
nand U3164 (N_3164,N_2993,N_2998);
nor U3165 (N_3165,N_2939,N_2519);
nor U3166 (N_3166,N_2729,N_2688);
nor U3167 (N_3167,N_2829,N_2600);
nand U3168 (N_3168,N_2931,N_2916);
and U3169 (N_3169,N_2854,N_2743);
and U3170 (N_3170,N_2633,N_2596);
and U3171 (N_3171,N_2949,N_2577);
or U3172 (N_3172,N_2793,N_2872);
or U3173 (N_3173,N_2846,N_2851);
nor U3174 (N_3174,N_2597,N_2948);
or U3175 (N_3175,N_2928,N_2996);
or U3176 (N_3176,N_2766,N_2569);
nand U3177 (N_3177,N_2716,N_2602);
or U3178 (N_3178,N_2975,N_2926);
nor U3179 (N_3179,N_2847,N_2773);
nor U3180 (N_3180,N_2869,N_2755);
or U3181 (N_3181,N_2663,N_2951);
or U3182 (N_3182,N_2580,N_2623);
nand U3183 (N_3183,N_2774,N_2673);
or U3184 (N_3184,N_2658,N_2731);
nor U3185 (N_3185,N_2759,N_2502);
nor U3186 (N_3186,N_2765,N_2938);
nor U3187 (N_3187,N_2963,N_2824);
nand U3188 (N_3188,N_2500,N_2815);
or U3189 (N_3189,N_2604,N_2549);
nor U3190 (N_3190,N_2506,N_2942);
nor U3191 (N_3191,N_2960,N_2516);
nor U3192 (N_3192,N_2962,N_2528);
nand U3193 (N_3193,N_2906,N_2720);
and U3194 (N_3194,N_2677,N_2836);
and U3195 (N_3195,N_2594,N_2546);
or U3196 (N_3196,N_2905,N_2811);
nand U3197 (N_3197,N_2921,N_2697);
or U3198 (N_3198,N_2636,N_2802);
nand U3199 (N_3199,N_2634,N_2608);
nor U3200 (N_3200,N_2558,N_2674);
or U3201 (N_3201,N_2511,N_2613);
or U3202 (N_3202,N_2554,N_2775);
and U3203 (N_3203,N_2992,N_2605);
or U3204 (N_3204,N_2503,N_2898);
nor U3205 (N_3205,N_2865,N_2601);
or U3206 (N_3206,N_2767,N_2681);
nor U3207 (N_3207,N_2656,N_2871);
and U3208 (N_3208,N_2999,N_2862);
and U3209 (N_3209,N_2797,N_2910);
and U3210 (N_3210,N_2944,N_2959);
or U3211 (N_3211,N_2630,N_2808);
or U3212 (N_3212,N_2666,N_2556);
or U3213 (N_3213,N_2786,N_2823);
and U3214 (N_3214,N_2509,N_2683);
or U3215 (N_3215,N_2885,N_2676);
nor U3216 (N_3216,N_2714,N_2883);
or U3217 (N_3217,N_2925,N_2645);
and U3218 (N_3218,N_2903,N_2707);
nand U3219 (N_3219,N_2555,N_2667);
and U3220 (N_3220,N_2990,N_2859);
nand U3221 (N_3221,N_2547,N_2779);
and U3222 (N_3222,N_2626,N_2726);
nor U3223 (N_3223,N_2832,N_2747);
nand U3224 (N_3224,N_2618,N_2969);
or U3225 (N_3225,N_2652,N_2530);
nand U3226 (N_3226,N_2713,N_2642);
or U3227 (N_3227,N_2825,N_2703);
nor U3228 (N_3228,N_2540,N_2738);
nor U3229 (N_3229,N_2834,N_2955);
nand U3230 (N_3230,N_2737,N_2661);
nor U3231 (N_3231,N_2875,N_2696);
nor U3232 (N_3232,N_2918,N_2783);
nand U3233 (N_3233,N_2876,N_2648);
or U3234 (N_3234,N_2571,N_2771);
or U3235 (N_3235,N_2740,N_2538);
or U3236 (N_3236,N_2782,N_2929);
xnor U3237 (N_3237,N_2542,N_2730);
or U3238 (N_3238,N_2861,N_2599);
or U3239 (N_3239,N_2684,N_2550);
or U3240 (N_3240,N_2657,N_2698);
nor U3241 (N_3241,N_2974,N_2660);
or U3242 (N_3242,N_2798,N_2945);
and U3243 (N_3243,N_2583,N_2578);
nor U3244 (N_3244,N_2574,N_2606);
and U3245 (N_3245,N_2923,N_2961);
or U3246 (N_3246,N_2828,N_2654);
nand U3247 (N_3247,N_2708,N_2722);
or U3248 (N_3248,N_2690,N_2968);
or U3249 (N_3249,N_2850,N_2521);
nand U3250 (N_3250,N_2564,N_2905);
or U3251 (N_3251,N_2870,N_2664);
nand U3252 (N_3252,N_2990,N_2665);
or U3253 (N_3253,N_2604,N_2889);
xnor U3254 (N_3254,N_2712,N_2645);
nand U3255 (N_3255,N_2745,N_2626);
nand U3256 (N_3256,N_2988,N_2917);
or U3257 (N_3257,N_2914,N_2813);
or U3258 (N_3258,N_2530,N_2808);
nand U3259 (N_3259,N_2748,N_2562);
nor U3260 (N_3260,N_2561,N_2659);
and U3261 (N_3261,N_2890,N_2801);
nand U3262 (N_3262,N_2694,N_2625);
nor U3263 (N_3263,N_2746,N_2965);
and U3264 (N_3264,N_2589,N_2957);
and U3265 (N_3265,N_2930,N_2807);
and U3266 (N_3266,N_2626,N_2662);
or U3267 (N_3267,N_2884,N_2793);
and U3268 (N_3268,N_2890,N_2994);
or U3269 (N_3269,N_2500,N_2799);
nand U3270 (N_3270,N_2957,N_2786);
or U3271 (N_3271,N_2822,N_2666);
or U3272 (N_3272,N_2835,N_2686);
and U3273 (N_3273,N_2516,N_2522);
nor U3274 (N_3274,N_2911,N_2976);
nor U3275 (N_3275,N_2838,N_2643);
xor U3276 (N_3276,N_2698,N_2601);
or U3277 (N_3277,N_2780,N_2834);
nor U3278 (N_3278,N_2626,N_2554);
nor U3279 (N_3279,N_2584,N_2687);
and U3280 (N_3280,N_2876,N_2762);
nand U3281 (N_3281,N_2602,N_2765);
nor U3282 (N_3282,N_2889,N_2895);
and U3283 (N_3283,N_2623,N_2620);
or U3284 (N_3284,N_2645,N_2577);
nand U3285 (N_3285,N_2677,N_2693);
nor U3286 (N_3286,N_2745,N_2664);
nand U3287 (N_3287,N_2811,N_2766);
and U3288 (N_3288,N_2607,N_2810);
or U3289 (N_3289,N_2675,N_2516);
nor U3290 (N_3290,N_2673,N_2681);
and U3291 (N_3291,N_2946,N_2876);
nand U3292 (N_3292,N_2665,N_2538);
or U3293 (N_3293,N_2728,N_2662);
nand U3294 (N_3294,N_2554,N_2933);
nor U3295 (N_3295,N_2536,N_2871);
and U3296 (N_3296,N_2612,N_2818);
nor U3297 (N_3297,N_2711,N_2956);
nand U3298 (N_3298,N_2846,N_2822);
nor U3299 (N_3299,N_2747,N_2901);
and U3300 (N_3300,N_2797,N_2819);
nand U3301 (N_3301,N_2898,N_2535);
nand U3302 (N_3302,N_2717,N_2751);
and U3303 (N_3303,N_2998,N_2725);
nand U3304 (N_3304,N_2571,N_2794);
nand U3305 (N_3305,N_2633,N_2676);
nand U3306 (N_3306,N_2877,N_2860);
nor U3307 (N_3307,N_2752,N_2793);
and U3308 (N_3308,N_2990,N_2612);
or U3309 (N_3309,N_2507,N_2506);
nand U3310 (N_3310,N_2977,N_2550);
nor U3311 (N_3311,N_2612,N_2580);
nor U3312 (N_3312,N_2836,N_2810);
nand U3313 (N_3313,N_2730,N_2558);
nand U3314 (N_3314,N_2851,N_2793);
or U3315 (N_3315,N_2900,N_2596);
or U3316 (N_3316,N_2642,N_2657);
and U3317 (N_3317,N_2957,N_2619);
and U3318 (N_3318,N_2882,N_2975);
nor U3319 (N_3319,N_2921,N_2608);
and U3320 (N_3320,N_2876,N_2738);
or U3321 (N_3321,N_2548,N_2875);
nand U3322 (N_3322,N_2967,N_2726);
or U3323 (N_3323,N_2843,N_2858);
or U3324 (N_3324,N_2704,N_2932);
and U3325 (N_3325,N_2744,N_2649);
nor U3326 (N_3326,N_2527,N_2713);
and U3327 (N_3327,N_2759,N_2873);
and U3328 (N_3328,N_2905,N_2699);
and U3329 (N_3329,N_2943,N_2595);
or U3330 (N_3330,N_2838,N_2603);
nand U3331 (N_3331,N_2801,N_2937);
or U3332 (N_3332,N_2890,N_2697);
nor U3333 (N_3333,N_2631,N_2613);
or U3334 (N_3334,N_2974,N_2648);
nor U3335 (N_3335,N_2731,N_2925);
or U3336 (N_3336,N_2840,N_2826);
nand U3337 (N_3337,N_2640,N_2896);
and U3338 (N_3338,N_2905,N_2896);
nor U3339 (N_3339,N_2724,N_2944);
or U3340 (N_3340,N_2938,N_2748);
and U3341 (N_3341,N_2783,N_2986);
nand U3342 (N_3342,N_2610,N_2900);
and U3343 (N_3343,N_2675,N_2594);
and U3344 (N_3344,N_2606,N_2842);
or U3345 (N_3345,N_2928,N_2886);
or U3346 (N_3346,N_2691,N_2872);
nor U3347 (N_3347,N_2966,N_2667);
or U3348 (N_3348,N_2946,N_2671);
nor U3349 (N_3349,N_2582,N_2984);
nand U3350 (N_3350,N_2689,N_2703);
nor U3351 (N_3351,N_2999,N_2705);
nand U3352 (N_3352,N_2974,N_2714);
or U3353 (N_3353,N_2551,N_2867);
nand U3354 (N_3354,N_2730,N_2601);
or U3355 (N_3355,N_2820,N_2979);
and U3356 (N_3356,N_2731,N_2578);
and U3357 (N_3357,N_2614,N_2559);
nand U3358 (N_3358,N_2552,N_2727);
nor U3359 (N_3359,N_2567,N_2512);
and U3360 (N_3360,N_2904,N_2578);
or U3361 (N_3361,N_2507,N_2646);
nor U3362 (N_3362,N_2905,N_2600);
or U3363 (N_3363,N_2683,N_2719);
nand U3364 (N_3364,N_2710,N_2771);
and U3365 (N_3365,N_2887,N_2856);
nor U3366 (N_3366,N_2546,N_2799);
and U3367 (N_3367,N_2704,N_2628);
and U3368 (N_3368,N_2661,N_2725);
or U3369 (N_3369,N_2558,N_2675);
nor U3370 (N_3370,N_2922,N_2904);
nand U3371 (N_3371,N_2674,N_2966);
or U3372 (N_3372,N_2773,N_2632);
and U3373 (N_3373,N_2512,N_2659);
nor U3374 (N_3374,N_2968,N_2752);
nor U3375 (N_3375,N_2855,N_2589);
nand U3376 (N_3376,N_2669,N_2723);
xor U3377 (N_3377,N_2947,N_2850);
nand U3378 (N_3378,N_2944,N_2826);
and U3379 (N_3379,N_2805,N_2530);
nor U3380 (N_3380,N_2797,N_2500);
and U3381 (N_3381,N_2677,N_2800);
nor U3382 (N_3382,N_2910,N_2733);
and U3383 (N_3383,N_2904,N_2703);
nand U3384 (N_3384,N_2522,N_2815);
nor U3385 (N_3385,N_2887,N_2906);
and U3386 (N_3386,N_2762,N_2825);
nor U3387 (N_3387,N_2638,N_2558);
and U3388 (N_3388,N_2515,N_2653);
nand U3389 (N_3389,N_2791,N_2732);
nand U3390 (N_3390,N_2865,N_2929);
nand U3391 (N_3391,N_2961,N_2548);
and U3392 (N_3392,N_2686,N_2560);
and U3393 (N_3393,N_2931,N_2613);
or U3394 (N_3394,N_2647,N_2803);
or U3395 (N_3395,N_2901,N_2637);
or U3396 (N_3396,N_2920,N_2691);
nor U3397 (N_3397,N_2782,N_2703);
and U3398 (N_3398,N_2700,N_2810);
nor U3399 (N_3399,N_2666,N_2617);
and U3400 (N_3400,N_2508,N_2864);
and U3401 (N_3401,N_2656,N_2615);
or U3402 (N_3402,N_2888,N_2647);
and U3403 (N_3403,N_2671,N_2689);
and U3404 (N_3404,N_2840,N_2651);
nand U3405 (N_3405,N_2829,N_2536);
nor U3406 (N_3406,N_2629,N_2883);
and U3407 (N_3407,N_2907,N_2900);
or U3408 (N_3408,N_2769,N_2707);
or U3409 (N_3409,N_2613,N_2604);
nor U3410 (N_3410,N_2816,N_2800);
nand U3411 (N_3411,N_2793,N_2719);
nor U3412 (N_3412,N_2832,N_2611);
or U3413 (N_3413,N_2932,N_2990);
nand U3414 (N_3414,N_2532,N_2743);
nor U3415 (N_3415,N_2692,N_2695);
nor U3416 (N_3416,N_2596,N_2652);
and U3417 (N_3417,N_2833,N_2986);
nor U3418 (N_3418,N_2974,N_2893);
nor U3419 (N_3419,N_2780,N_2517);
nor U3420 (N_3420,N_2776,N_2837);
and U3421 (N_3421,N_2632,N_2840);
and U3422 (N_3422,N_2700,N_2832);
nand U3423 (N_3423,N_2794,N_2560);
nor U3424 (N_3424,N_2868,N_2653);
nor U3425 (N_3425,N_2797,N_2958);
nor U3426 (N_3426,N_2679,N_2587);
or U3427 (N_3427,N_2752,N_2884);
or U3428 (N_3428,N_2953,N_2598);
or U3429 (N_3429,N_2644,N_2566);
nand U3430 (N_3430,N_2866,N_2528);
nor U3431 (N_3431,N_2545,N_2949);
nor U3432 (N_3432,N_2820,N_2510);
nand U3433 (N_3433,N_2711,N_2960);
nor U3434 (N_3434,N_2831,N_2999);
or U3435 (N_3435,N_2742,N_2641);
or U3436 (N_3436,N_2656,N_2824);
nor U3437 (N_3437,N_2678,N_2568);
nand U3438 (N_3438,N_2875,N_2925);
and U3439 (N_3439,N_2794,N_2562);
or U3440 (N_3440,N_2712,N_2564);
and U3441 (N_3441,N_2753,N_2899);
and U3442 (N_3442,N_2993,N_2658);
nor U3443 (N_3443,N_2923,N_2848);
or U3444 (N_3444,N_2729,N_2527);
and U3445 (N_3445,N_2978,N_2837);
nor U3446 (N_3446,N_2676,N_2626);
or U3447 (N_3447,N_2704,N_2648);
nand U3448 (N_3448,N_2631,N_2761);
or U3449 (N_3449,N_2879,N_2632);
nor U3450 (N_3450,N_2530,N_2842);
nor U3451 (N_3451,N_2804,N_2505);
nand U3452 (N_3452,N_2807,N_2977);
or U3453 (N_3453,N_2756,N_2737);
and U3454 (N_3454,N_2992,N_2997);
nand U3455 (N_3455,N_2919,N_2929);
nor U3456 (N_3456,N_2854,N_2603);
or U3457 (N_3457,N_2687,N_2941);
and U3458 (N_3458,N_2621,N_2526);
nand U3459 (N_3459,N_2852,N_2872);
or U3460 (N_3460,N_2802,N_2572);
and U3461 (N_3461,N_2870,N_2617);
nand U3462 (N_3462,N_2629,N_2723);
or U3463 (N_3463,N_2560,N_2612);
nor U3464 (N_3464,N_2736,N_2656);
or U3465 (N_3465,N_2626,N_2584);
or U3466 (N_3466,N_2645,N_2900);
and U3467 (N_3467,N_2950,N_2946);
or U3468 (N_3468,N_2710,N_2536);
nand U3469 (N_3469,N_2602,N_2701);
nand U3470 (N_3470,N_2928,N_2966);
or U3471 (N_3471,N_2632,N_2605);
nand U3472 (N_3472,N_2658,N_2593);
nand U3473 (N_3473,N_2675,N_2830);
nor U3474 (N_3474,N_2898,N_2855);
and U3475 (N_3475,N_2976,N_2592);
nand U3476 (N_3476,N_2744,N_2742);
nand U3477 (N_3477,N_2575,N_2768);
or U3478 (N_3478,N_2842,N_2754);
nand U3479 (N_3479,N_2967,N_2979);
and U3480 (N_3480,N_2851,N_2605);
nor U3481 (N_3481,N_2775,N_2637);
nand U3482 (N_3482,N_2572,N_2748);
and U3483 (N_3483,N_2753,N_2897);
and U3484 (N_3484,N_2958,N_2750);
nor U3485 (N_3485,N_2766,N_2955);
and U3486 (N_3486,N_2509,N_2836);
nor U3487 (N_3487,N_2914,N_2537);
and U3488 (N_3488,N_2620,N_2879);
and U3489 (N_3489,N_2755,N_2571);
and U3490 (N_3490,N_2610,N_2546);
nor U3491 (N_3491,N_2885,N_2639);
or U3492 (N_3492,N_2972,N_2828);
or U3493 (N_3493,N_2856,N_2980);
or U3494 (N_3494,N_2768,N_2853);
nor U3495 (N_3495,N_2512,N_2947);
nor U3496 (N_3496,N_2742,N_2540);
nor U3497 (N_3497,N_2925,N_2771);
nor U3498 (N_3498,N_2734,N_2571);
nor U3499 (N_3499,N_2816,N_2798);
nor U3500 (N_3500,N_3160,N_3477);
nor U3501 (N_3501,N_3004,N_3220);
nor U3502 (N_3502,N_3460,N_3494);
nor U3503 (N_3503,N_3044,N_3439);
and U3504 (N_3504,N_3257,N_3221);
nor U3505 (N_3505,N_3045,N_3374);
nand U3506 (N_3506,N_3147,N_3383);
nand U3507 (N_3507,N_3134,N_3133);
xor U3508 (N_3508,N_3096,N_3017);
or U3509 (N_3509,N_3399,N_3464);
nand U3510 (N_3510,N_3060,N_3027);
nor U3511 (N_3511,N_3358,N_3371);
and U3512 (N_3512,N_3061,N_3049);
nand U3513 (N_3513,N_3122,N_3127);
and U3514 (N_3514,N_3055,N_3236);
and U3515 (N_3515,N_3175,N_3142);
nor U3516 (N_3516,N_3245,N_3014);
or U3517 (N_3517,N_3080,N_3113);
or U3518 (N_3518,N_3377,N_3214);
and U3519 (N_3519,N_3025,N_3046);
nor U3520 (N_3520,N_3264,N_3429);
nor U3521 (N_3521,N_3106,N_3481);
nor U3522 (N_3522,N_3135,N_3485);
nand U3523 (N_3523,N_3354,N_3253);
and U3524 (N_3524,N_3433,N_3097);
nor U3525 (N_3525,N_3015,N_3416);
nor U3526 (N_3526,N_3476,N_3376);
nor U3527 (N_3527,N_3161,N_3471);
nand U3528 (N_3528,N_3090,N_3149);
or U3529 (N_3529,N_3265,N_3187);
nor U3530 (N_3530,N_3268,N_3283);
or U3531 (N_3531,N_3037,N_3168);
nor U3532 (N_3532,N_3478,N_3100);
and U3533 (N_3533,N_3165,N_3255);
nor U3534 (N_3534,N_3269,N_3229);
nand U3535 (N_3535,N_3170,N_3203);
nand U3536 (N_3536,N_3288,N_3086);
and U3537 (N_3537,N_3370,N_3167);
and U3538 (N_3538,N_3031,N_3355);
nand U3539 (N_3539,N_3330,N_3217);
or U3540 (N_3540,N_3453,N_3091);
and U3541 (N_3541,N_3077,N_3419);
nor U3542 (N_3542,N_3201,N_3137);
and U3543 (N_3543,N_3191,N_3144);
or U3544 (N_3544,N_3036,N_3448);
and U3545 (N_3545,N_3298,N_3223);
nand U3546 (N_3546,N_3193,N_3305);
or U3547 (N_3547,N_3226,N_3342);
nand U3548 (N_3548,N_3001,N_3428);
and U3549 (N_3549,N_3467,N_3402);
and U3550 (N_3550,N_3317,N_3480);
or U3551 (N_3551,N_3300,N_3483);
or U3552 (N_3552,N_3486,N_3256);
nor U3553 (N_3553,N_3387,N_3487);
or U3554 (N_3554,N_3436,N_3301);
or U3555 (N_3555,N_3224,N_3280);
or U3556 (N_3556,N_3492,N_3414);
nor U3557 (N_3557,N_3169,N_3457);
nor U3558 (N_3558,N_3115,N_3083);
nand U3559 (N_3559,N_3089,N_3472);
or U3560 (N_3560,N_3054,N_3219);
and U3561 (N_3561,N_3351,N_3064);
nor U3562 (N_3562,N_3328,N_3171);
or U3563 (N_3563,N_3456,N_3353);
or U3564 (N_3564,N_3408,N_3141);
nand U3565 (N_3565,N_3110,N_3199);
nor U3566 (N_3566,N_3067,N_3121);
nand U3567 (N_3567,N_3407,N_3378);
nand U3568 (N_3568,N_3120,N_3043);
and U3569 (N_3569,N_3241,N_3381);
and U3570 (N_3570,N_3275,N_3156);
xnor U3571 (N_3571,N_3286,N_3003);
nor U3572 (N_3572,N_3279,N_3430);
and U3573 (N_3573,N_3158,N_3357);
and U3574 (N_3574,N_3196,N_3272);
and U3575 (N_3575,N_3021,N_3173);
nand U3576 (N_3576,N_3291,N_3386);
or U3577 (N_3577,N_3350,N_3271);
or U3578 (N_3578,N_3002,N_3069);
and U3579 (N_3579,N_3406,N_3440);
or U3580 (N_3580,N_3493,N_3312);
nor U3581 (N_3581,N_3023,N_3356);
and U3582 (N_3582,N_3375,N_3028);
nor U3583 (N_3583,N_3461,N_3012);
nor U3584 (N_3584,N_3401,N_3324);
and U3585 (N_3585,N_3212,N_3185);
and U3586 (N_3586,N_3232,N_3125);
xnor U3587 (N_3587,N_3333,N_3108);
and U3588 (N_3588,N_3183,N_3336);
and U3589 (N_3589,N_3085,N_3029);
or U3590 (N_3590,N_3020,N_3435);
nand U3591 (N_3591,N_3200,N_3395);
or U3592 (N_3592,N_3344,N_3289);
nor U3593 (N_3593,N_3321,N_3058);
nand U3594 (N_3594,N_3182,N_3403);
or U3595 (N_3595,N_3041,N_3062);
and U3596 (N_3596,N_3458,N_3293);
nor U3597 (N_3597,N_3186,N_3410);
nor U3598 (N_3598,N_3263,N_3206);
nand U3599 (N_3599,N_3011,N_3065);
nor U3600 (N_3600,N_3415,N_3208);
nand U3601 (N_3601,N_3299,N_3207);
or U3602 (N_3602,N_3024,N_3442);
and U3603 (N_3603,N_3252,N_3192);
nor U3604 (N_3604,N_3095,N_3038);
and U3605 (N_3605,N_3155,N_3325);
nor U3606 (N_3606,N_3094,N_3396);
nor U3607 (N_3607,N_3444,N_3007);
nor U3608 (N_3608,N_3304,N_3088);
nand U3609 (N_3609,N_3222,N_3490);
and U3610 (N_3610,N_3303,N_3392);
nor U3611 (N_3611,N_3382,N_3384);
nand U3612 (N_3612,N_3451,N_3248);
and U3613 (N_3613,N_3260,N_3393);
and U3614 (N_3614,N_3176,N_3491);
nand U3615 (N_3615,N_3297,N_3425);
and U3616 (N_3616,N_3282,N_3322);
or U3617 (N_3617,N_3126,N_3261);
nand U3618 (N_3618,N_3215,N_3475);
nor U3619 (N_3619,N_3441,N_3231);
nand U3620 (N_3620,N_3163,N_3497);
nand U3621 (N_3621,N_3057,N_3109);
nand U3622 (N_3622,N_3296,N_3309);
nand U3623 (N_3623,N_3400,N_3104);
and U3624 (N_3624,N_3213,N_3019);
and U3625 (N_3625,N_3420,N_3434);
nor U3626 (N_3626,N_3499,N_3398);
or U3627 (N_3627,N_3107,N_3445);
nor U3628 (N_3628,N_3427,N_3285);
or U3629 (N_3629,N_3438,N_3459);
and U3630 (N_3630,N_3240,N_3372);
or U3631 (N_3631,N_3292,N_3337);
and U3632 (N_3632,N_3359,N_3202);
nand U3633 (N_3633,N_3323,N_3394);
and U3634 (N_3634,N_3413,N_3363);
or U3635 (N_3635,N_3112,N_3313);
nand U3636 (N_3636,N_3194,N_3295);
nand U3637 (N_3637,N_3010,N_3216);
or U3638 (N_3638,N_3385,N_3454);
nor U3639 (N_3639,N_3397,N_3235);
and U3640 (N_3640,N_3103,N_3138);
nand U3641 (N_3641,N_3152,N_3349);
and U3642 (N_3642,N_3123,N_3034);
nor U3643 (N_3643,N_3172,N_3076);
or U3644 (N_3644,N_3048,N_3056);
nand U3645 (N_3645,N_3450,N_3154);
nor U3646 (N_3646,N_3243,N_3273);
or U3647 (N_3647,N_3465,N_3379);
nor U3648 (N_3648,N_3190,N_3008);
and U3649 (N_3649,N_3059,N_3130);
and U3650 (N_3650,N_3022,N_3005);
or U3651 (N_3651,N_3405,N_3119);
and U3652 (N_3652,N_3489,N_3117);
and U3653 (N_3653,N_3033,N_3074);
and U3654 (N_3654,N_3227,N_3341);
nor U3655 (N_3655,N_3267,N_3150);
or U3656 (N_3656,N_3079,N_3431);
nand U3657 (N_3657,N_3035,N_3040);
and U3658 (N_3658,N_3073,N_3262);
and U3659 (N_3659,N_3075,N_3482);
nor U3660 (N_3660,N_3488,N_3391);
or U3661 (N_3661,N_3166,N_3159);
nand U3662 (N_3662,N_3345,N_3181);
or U3663 (N_3663,N_3140,N_3306);
nor U3664 (N_3664,N_3270,N_3237);
nor U3665 (N_3665,N_3361,N_3198);
nor U3666 (N_3666,N_3278,N_3225);
nor U3667 (N_3667,N_3098,N_3013);
or U3668 (N_3668,N_3368,N_3211);
nand U3669 (N_3669,N_3334,N_3039);
or U3670 (N_3670,N_3006,N_3143);
nor U3671 (N_3671,N_3189,N_3238);
and U3672 (N_3672,N_3145,N_3082);
or U3673 (N_3673,N_3174,N_3246);
nor U3674 (N_3674,N_3209,N_3327);
nand U3675 (N_3675,N_3116,N_3228);
or U3676 (N_3676,N_3131,N_3178);
nor U3677 (N_3677,N_3151,N_3360);
or U3678 (N_3678,N_3157,N_3281);
and U3679 (N_3679,N_3446,N_3409);
and U3680 (N_3680,N_3426,N_3466);
nor U3681 (N_3681,N_3188,N_3026);
nand U3682 (N_3682,N_3197,N_3093);
or U3683 (N_3683,N_3463,N_3329);
nor U3684 (N_3684,N_3072,N_3081);
nand U3685 (N_3685,N_3352,N_3332);
or U3686 (N_3686,N_3251,N_3422);
and U3687 (N_3687,N_3418,N_3244);
nand U3688 (N_3688,N_3318,N_3259);
or U3689 (N_3689,N_3099,N_3452);
and U3690 (N_3690,N_3469,N_3326);
and U3691 (N_3691,N_3230,N_3319);
or U3692 (N_3692,N_3473,N_3348);
and U3693 (N_3693,N_3102,N_3484);
nand U3694 (N_3694,N_3364,N_3071);
nand U3695 (N_3695,N_3447,N_3432);
nor U3696 (N_3696,N_3070,N_3016);
and U3697 (N_3697,N_3316,N_3314);
nand U3698 (N_3698,N_3114,N_3294);
nor U3699 (N_3699,N_3346,N_3132);
and U3700 (N_3700,N_3498,N_3195);
nand U3701 (N_3701,N_3366,N_3404);
and U3702 (N_3702,N_3302,N_3000);
or U3703 (N_3703,N_3277,N_3105);
nand U3704 (N_3704,N_3479,N_3320);
or U3705 (N_3705,N_3247,N_3210);
nor U3706 (N_3706,N_3412,N_3276);
and U3707 (N_3707,N_3335,N_3424);
nor U3708 (N_3708,N_3339,N_3290);
nand U3709 (N_3709,N_3331,N_3139);
nor U3710 (N_3710,N_3051,N_3032);
or U3711 (N_3711,N_3087,N_3084);
nor U3712 (N_3712,N_3343,N_3148);
or U3713 (N_3713,N_3030,N_3411);
or U3714 (N_3714,N_3249,N_3233);
nor U3715 (N_3715,N_3254,N_3179);
and U3716 (N_3716,N_3164,N_3052);
nor U3717 (N_3717,N_3242,N_3129);
nand U3718 (N_3718,N_3449,N_3218);
nand U3719 (N_3719,N_3496,N_3362);
nand U3720 (N_3720,N_3307,N_3340);
nor U3721 (N_3721,N_3347,N_3101);
nand U3722 (N_3722,N_3287,N_3423);
xnor U3723 (N_3723,N_3417,N_3205);
and U3724 (N_3724,N_3388,N_3068);
nor U3725 (N_3725,N_3443,N_3162);
nor U3726 (N_3726,N_3310,N_3470);
nand U3727 (N_3727,N_3308,N_3234);
or U3728 (N_3728,N_3258,N_3421);
and U3729 (N_3729,N_3380,N_3266);
nor U3730 (N_3730,N_3042,N_3136);
and U3731 (N_3731,N_3390,N_3250);
or U3732 (N_3732,N_3311,N_3365);
or U3733 (N_3733,N_3315,N_3177);
nand U3734 (N_3734,N_3389,N_3124);
nor U3735 (N_3735,N_3066,N_3128);
nor U3736 (N_3736,N_3437,N_3204);
nand U3737 (N_3737,N_3239,N_3468);
nor U3738 (N_3738,N_3050,N_3338);
nand U3739 (N_3739,N_3284,N_3092);
nor U3740 (N_3740,N_3367,N_3047);
nor U3741 (N_3741,N_3180,N_3495);
nand U3742 (N_3742,N_3153,N_3369);
nor U3743 (N_3743,N_3078,N_3009);
or U3744 (N_3744,N_3118,N_3063);
nand U3745 (N_3745,N_3455,N_3111);
nor U3746 (N_3746,N_3462,N_3274);
and U3747 (N_3747,N_3373,N_3184);
nor U3748 (N_3748,N_3146,N_3018);
nor U3749 (N_3749,N_3053,N_3474);
nand U3750 (N_3750,N_3416,N_3141);
or U3751 (N_3751,N_3318,N_3391);
or U3752 (N_3752,N_3379,N_3132);
or U3753 (N_3753,N_3370,N_3335);
nor U3754 (N_3754,N_3382,N_3348);
and U3755 (N_3755,N_3400,N_3410);
or U3756 (N_3756,N_3285,N_3018);
nor U3757 (N_3757,N_3339,N_3495);
or U3758 (N_3758,N_3333,N_3015);
and U3759 (N_3759,N_3310,N_3119);
or U3760 (N_3760,N_3209,N_3189);
nand U3761 (N_3761,N_3183,N_3169);
and U3762 (N_3762,N_3170,N_3063);
or U3763 (N_3763,N_3275,N_3377);
or U3764 (N_3764,N_3007,N_3256);
and U3765 (N_3765,N_3183,N_3290);
nand U3766 (N_3766,N_3299,N_3455);
nor U3767 (N_3767,N_3448,N_3160);
and U3768 (N_3768,N_3143,N_3414);
nand U3769 (N_3769,N_3129,N_3486);
nand U3770 (N_3770,N_3009,N_3353);
nor U3771 (N_3771,N_3027,N_3125);
and U3772 (N_3772,N_3346,N_3120);
nor U3773 (N_3773,N_3283,N_3008);
or U3774 (N_3774,N_3234,N_3486);
or U3775 (N_3775,N_3041,N_3087);
nor U3776 (N_3776,N_3186,N_3356);
nand U3777 (N_3777,N_3233,N_3096);
and U3778 (N_3778,N_3154,N_3260);
or U3779 (N_3779,N_3179,N_3004);
nand U3780 (N_3780,N_3066,N_3225);
or U3781 (N_3781,N_3440,N_3224);
and U3782 (N_3782,N_3111,N_3322);
nor U3783 (N_3783,N_3253,N_3475);
or U3784 (N_3784,N_3159,N_3181);
nor U3785 (N_3785,N_3237,N_3376);
and U3786 (N_3786,N_3001,N_3119);
nand U3787 (N_3787,N_3010,N_3095);
nand U3788 (N_3788,N_3442,N_3160);
and U3789 (N_3789,N_3381,N_3300);
nand U3790 (N_3790,N_3103,N_3365);
nand U3791 (N_3791,N_3291,N_3287);
nand U3792 (N_3792,N_3402,N_3499);
nand U3793 (N_3793,N_3479,N_3445);
or U3794 (N_3794,N_3463,N_3247);
nor U3795 (N_3795,N_3336,N_3089);
and U3796 (N_3796,N_3221,N_3311);
nand U3797 (N_3797,N_3337,N_3113);
or U3798 (N_3798,N_3346,N_3489);
nand U3799 (N_3799,N_3025,N_3261);
and U3800 (N_3800,N_3301,N_3077);
or U3801 (N_3801,N_3365,N_3440);
or U3802 (N_3802,N_3460,N_3229);
and U3803 (N_3803,N_3345,N_3395);
nand U3804 (N_3804,N_3084,N_3376);
nor U3805 (N_3805,N_3225,N_3121);
or U3806 (N_3806,N_3405,N_3107);
or U3807 (N_3807,N_3495,N_3257);
or U3808 (N_3808,N_3276,N_3025);
or U3809 (N_3809,N_3162,N_3333);
nor U3810 (N_3810,N_3321,N_3333);
nor U3811 (N_3811,N_3158,N_3459);
nand U3812 (N_3812,N_3270,N_3365);
nor U3813 (N_3813,N_3098,N_3195);
or U3814 (N_3814,N_3482,N_3166);
and U3815 (N_3815,N_3304,N_3305);
and U3816 (N_3816,N_3424,N_3451);
or U3817 (N_3817,N_3006,N_3493);
nand U3818 (N_3818,N_3018,N_3340);
or U3819 (N_3819,N_3375,N_3200);
nand U3820 (N_3820,N_3241,N_3214);
or U3821 (N_3821,N_3166,N_3314);
nand U3822 (N_3822,N_3385,N_3126);
and U3823 (N_3823,N_3432,N_3451);
nor U3824 (N_3824,N_3450,N_3389);
nand U3825 (N_3825,N_3195,N_3429);
nand U3826 (N_3826,N_3252,N_3012);
or U3827 (N_3827,N_3016,N_3294);
nand U3828 (N_3828,N_3312,N_3094);
nand U3829 (N_3829,N_3010,N_3299);
nor U3830 (N_3830,N_3247,N_3224);
xor U3831 (N_3831,N_3332,N_3273);
or U3832 (N_3832,N_3394,N_3322);
and U3833 (N_3833,N_3179,N_3309);
or U3834 (N_3834,N_3171,N_3381);
and U3835 (N_3835,N_3076,N_3337);
nand U3836 (N_3836,N_3159,N_3499);
or U3837 (N_3837,N_3102,N_3379);
nand U3838 (N_3838,N_3008,N_3002);
nor U3839 (N_3839,N_3109,N_3004);
xnor U3840 (N_3840,N_3016,N_3051);
or U3841 (N_3841,N_3410,N_3453);
xor U3842 (N_3842,N_3128,N_3479);
nand U3843 (N_3843,N_3473,N_3210);
nand U3844 (N_3844,N_3499,N_3467);
and U3845 (N_3845,N_3116,N_3104);
and U3846 (N_3846,N_3160,N_3289);
or U3847 (N_3847,N_3100,N_3329);
nand U3848 (N_3848,N_3161,N_3099);
and U3849 (N_3849,N_3439,N_3345);
and U3850 (N_3850,N_3390,N_3261);
and U3851 (N_3851,N_3173,N_3215);
nor U3852 (N_3852,N_3004,N_3120);
nor U3853 (N_3853,N_3292,N_3210);
and U3854 (N_3854,N_3475,N_3054);
and U3855 (N_3855,N_3347,N_3484);
and U3856 (N_3856,N_3272,N_3151);
nand U3857 (N_3857,N_3062,N_3111);
nand U3858 (N_3858,N_3281,N_3063);
nand U3859 (N_3859,N_3005,N_3183);
and U3860 (N_3860,N_3347,N_3346);
nand U3861 (N_3861,N_3137,N_3391);
and U3862 (N_3862,N_3224,N_3389);
nand U3863 (N_3863,N_3354,N_3192);
nor U3864 (N_3864,N_3260,N_3461);
or U3865 (N_3865,N_3063,N_3120);
or U3866 (N_3866,N_3497,N_3322);
or U3867 (N_3867,N_3421,N_3050);
nor U3868 (N_3868,N_3292,N_3401);
and U3869 (N_3869,N_3203,N_3208);
nor U3870 (N_3870,N_3217,N_3034);
or U3871 (N_3871,N_3099,N_3251);
and U3872 (N_3872,N_3081,N_3051);
or U3873 (N_3873,N_3150,N_3050);
and U3874 (N_3874,N_3255,N_3321);
or U3875 (N_3875,N_3154,N_3098);
and U3876 (N_3876,N_3078,N_3491);
or U3877 (N_3877,N_3094,N_3028);
nor U3878 (N_3878,N_3494,N_3358);
or U3879 (N_3879,N_3109,N_3434);
and U3880 (N_3880,N_3233,N_3143);
nand U3881 (N_3881,N_3325,N_3492);
nor U3882 (N_3882,N_3342,N_3314);
nand U3883 (N_3883,N_3258,N_3223);
nand U3884 (N_3884,N_3014,N_3313);
or U3885 (N_3885,N_3445,N_3222);
or U3886 (N_3886,N_3289,N_3128);
and U3887 (N_3887,N_3489,N_3119);
nand U3888 (N_3888,N_3460,N_3035);
or U3889 (N_3889,N_3362,N_3269);
nor U3890 (N_3890,N_3329,N_3295);
nand U3891 (N_3891,N_3327,N_3174);
nor U3892 (N_3892,N_3325,N_3331);
nor U3893 (N_3893,N_3343,N_3077);
nor U3894 (N_3894,N_3233,N_3473);
xor U3895 (N_3895,N_3463,N_3250);
xnor U3896 (N_3896,N_3450,N_3453);
nand U3897 (N_3897,N_3368,N_3228);
or U3898 (N_3898,N_3372,N_3451);
nor U3899 (N_3899,N_3216,N_3232);
nand U3900 (N_3900,N_3312,N_3084);
and U3901 (N_3901,N_3423,N_3249);
nor U3902 (N_3902,N_3065,N_3458);
nor U3903 (N_3903,N_3095,N_3241);
nand U3904 (N_3904,N_3394,N_3138);
nand U3905 (N_3905,N_3207,N_3469);
nand U3906 (N_3906,N_3022,N_3235);
and U3907 (N_3907,N_3054,N_3353);
and U3908 (N_3908,N_3136,N_3409);
nor U3909 (N_3909,N_3028,N_3308);
and U3910 (N_3910,N_3489,N_3466);
nor U3911 (N_3911,N_3349,N_3451);
nand U3912 (N_3912,N_3238,N_3350);
nand U3913 (N_3913,N_3306,N_3232);
nor U3914 (N_3914,N_3062,N_3245);
or U3915 (N_3915,N_3149,N_3257);
or U3916 (N_3916,N_3024,N_3065);
or U3917 (N_3917,N_3466,N_3087);
or U3918 (N_3918,N_3304,N_3290);
nand U3919 (N_3919,N_3452,N_3391);
nor U3920 (N_3920,N_3132,N_3415);
nor U3921 (N_3921,N_3183,N_3107);
nand U3922 (N_3922,N_3315,N_3354);
or U3923 (N_3923,N_3153,N_3363);
nor U3924 (N_3924,N_3162,N_3044);
nor U3925 (N_3925,N_3209,N_3414);
and U3926 (N_3926,N_3469,N_3037);
and U3927 (N_3927,N_3206,N_3339);
or U3928 (N_3928,N_3282,N_3465);
nor U3929 (N_3929,N_3340,N_3190);
or U3930 (N_3930,N_3192,N_3390);
nand U3931 (N_3931,N_3016,N_3388);
nor U3932 (N_3932,N_3043,N_3279);
or U3933 (N_3933,N_3131,N_3382);
or U3934 (N_3934,N_3024,N_3012);
and U3935 (N_3935,N_3046,N_3448);
or U3936 (N_3936,N_3380,N_3429);
and U3937 (N_3937,N_3234,N_3249);
nand U3938 (N_3938,N_3184,N_3403);
nand U3939 (N_3939,N_3356,N_3123);
or U3940 (N_3940,N_3110,N_3238);
or U3941 (N_3941,N_3115,N_3256);
nor U3942 (N_3942,N_3130,N_3218);
nand U3943 (N_3943,N_3355,N_3112);
and U3944 (N_3944,N_3284,N_3279);
or U3945 (N_3945,N_3218,N_3076);
or U3946 (N_3946,N_3361,N_3356);
nand U3947 (N_3947,N_3118,N_3078);
and U3948 (N_3948,N_3013,N_3452);
and U3949 (N_3949,N_3019,N_3245);
and U3950 (N_3950,N_3422,N_3095);
and U3951 (N_3951,N_3090,N_3020);
and U3952 (N_3952,N_3306,N_3187);
and U3953 (N_3953,N_3065,N_3397);
or U3954 (N_3954,N_3405,N_3301);
or U3955 (N_3955,N_3403,N_3130);
or U3956 (N_3956,N_3227,N_3131);
or U3957 (N_3957,N_3178,N_3139);
nor U3958 (N_3958,N_3397,N_3069);
and U3959 (N_3959,N_3217,N_3413);
nand U3960 (N_3960,N_3400,N_3129);
and U3961 (N_3961,N_3057,N_3457);
nand U3962 (N_3962,N_3092,N_3162);
and U3963 (N_3963,N_3131,N_3118);
and U3964 (N_3964,N_3343,N_3213);
or U3965 (N_3965,N_3043,N_3328);
nor U3966 (N_3966,N_3005,N_3167);
nand U3967 (N_3967,N_3445,N_3356);
nor U3968 (N_3968,N_3014,N_3124);
nor U3969 (N_3969,N_3269,N_3424);
nand U3970 (N_3970,N_3252,N_3160);
or U3971 (N_3971,N_3141,N_3200);
nor U3972 (N_3972,N_3432,N_3245);
nor U3973 (N_3973,N_3332,N_3244);
nand U3974 (N_3974,N_3378,N_3151);
and U3975 (N_3975,N_3279,N_3206);
or U3976 (N_3976,N_3483,N_3371);
nand U3977 (N_3977,N_3491,N_3223);
nand U3978 (N_3978,N_3130,N_3167);
nand U3979 (N_3979,N_3132,N_3152);
nand U3980 (N_3980,N_3112,N_3180);
and U3981 (N_3981,N_3112,N_3013);
nand U3982 (N_3982,N_3377,N_3248);
nor U3983 (N_3983,N_3123,N_3153);
nand U3984 (N_3984,N_3422,N_3461);
and U3985 (N_3985,N_3343,N_3426);
or U3986 (N_3986,N_3136,N_3494);
nand U3987 (N_3987,N_3119,N_3378);
and U3988 (N_3988,N_3024,N_3300);
or U3989 (N_3989,N_3358,N_3090);
nor U3990 (N_3990,N_3195,N_3108);
and U3991 (N_3991,N_3297,N_3149);
and U3992 (N_3992,N_3368,N_3005);
or U3993 (N_3993,N_3059,N_3282);
or U3994 (N_3994,N_3476,N_3119);
nor U3995 (N_3995,N_3496,N_3177);
nand U3996 (N_3996,N_3098,N_3407);
nand U3997 (N_3997,N_3378,N_3198);
nand U3998 (N_3998,N_3476,N_3039);
and U3999 (N_3999,N_3453,N_3226);
nand U4000 (N_4000,N_3805,N_3937);
or U4001 (N_4001,N_3702,N_3698);
or U4002 (N_4002,N_3783,N_3674);
and U4003 (N_4003,N_3505,N_3885);
and U4004 (N_4004,N_3917,N_3817);
nand U4005 (N_4005,N_3528,N_3942);
nand U4006 (N_4006,N_3566,N_3831);
nor U4007 (N_4007,N_3875,N_3830);
or U4008 (N_4008,N_3992,N_3598);
nand U4009 (N_4009,N_3696,N_3761);
nand U4010 (N_4010,N_3539,N_3624);
nand U4011 (N_4011,N_3789,N_3765);
nand U4012 (N_4012,N_3990,N_3754);
and U4013 (N_4013,N_3526,N_3959);
and U4014 (N_4014,N_3997,N_3685);
nand U4015 (N_4015,N_3623,N_3574);
or U4016 (N_4016,N_3671,N_3512);
nand U4017 (N_4017,N_3953,N_3824);
or U4018 (N_4018,N_3715,N_3753);
and U4019 (N_4019,N_3838,N_3889);
and U4020 (N_4020,N_3515,N_3676);
and U4021 (N_4021,N_3656,N_3866);
nor U4022 (N_4022,N_3617,N_3701);
nand U4023 (N_4023,N_3968,N_3863);
nor U4024 (N_4024,N_3669,N_3606);
nor U4025 (N_4025,N_3800,N_3864);
or U4026 (N_4026,N_3938,N_3544);
nand U4027 (N_4027,N_3768,N_3608);
and U4028 (N_4028,N_3548,N_3776);
and U4029 (N_4029,N_3913,N_3688);
or U4030 (N_4030,N_3999,N_3891);
and U4031 (N_4031,N_3711,N_3507);
and U4032 (N_4032,N_3991,N_3687);
or U4033 (N_4033,N_3995,N_3751);
and U4034 (N_4034,N_3612,N_3533);
and U4035 (N_4035,N_3731,N_3684);
or U4036 (N_4036,N_3925,N_3918);
and U4037 (N_4037,N_3758,N_3596);
and U4038 (N_4038,N_3663,N_3910);
or U4039 (N_4039,N_3589,N_3924);
nand U4040 (N_4040,N_3996,N_3895);
nand U4041 (N_4041,N_3736,N_3646);
nor U4042 (N_4042,N_3590,N_3974);
nand U4043 (N_4043,N_3607,N_3909);
or U4044 (N_4044,N_3841,N_3954);
nand U4045 (N_4045,N_3520,N_3662);
nand U4046 (N_4046,N_3767,N_3639);
or U4047 (N_4047,N_3522,N_3980);
nand U4048 (N_4048,N_3986,N_3989);
nand U4049 (N_4049,N_3724,N_3616);
nand U4050 (N_4050,N_3788,N_3772);
or U4051 (N_4051,N_3549,N_3967);
or U4052 (N_4052,N_3970,N_3689);
or U4053 (N_4053,N_3920,N_3745);
or U4054 (N_4054,N_3835,N_3700);
or U4055 (N_4055,N_3516,N_3706);
or U4056 (N_4056,N_3638,N_3538);
nand U4057 (N_4057,N_3903,N_3501);
nor U4058 (N_4058,N_3845,N_3525);
nand U4059 (N_4059,N_3908,N_3605);
xnor U4060 (N_4060,N_3813,N_3514);
and U4061 (N_4061,N_3553,N_3868);
nor U4062 (N_4062,N_3630,N_3641);
nor U4063 (N_4063,N_3665,N_3977);
nor U4064 (N_4064,N_3948,N_3531);
nor U4065 (N_4065,N_3880,N_3878);
nor U4066 (N_4066,N_3994,N_3527);
nand U4067 (N_4067,N_3626,N_3896);
nor U4068 (N_4068,N_3567,N_3771);
or U4069 (N_4069,N_3927,N_3888);
or U4070 (N_4070,N_3844,N_3584);
nor U4071 (N_4071,N_3945,N_3562);
nor U4072 (N_4072,N_3764,N_3691);
or U4073 (N_4073,N_3934,N_3818);
and U4074 (N_4074,N_3550,N_3826);
nand U4075 (N_4075,N_3756,N_3946);
nand U4076 (N_4076,N_3849,N_3710);
nor U4077 (N_4077,N_3618,N_3784);
xnor U4078 (N_4078,N_3673,N_3517);
and U4079 (N_4079,N_3931,N_3523);
or U4080 (N_4080,N_3703,N_3983);
nor U4081 (N_4081,N_3763,N_3949);
or U4082 (N_4082,N_3534,N_3922);
nor U4083 (N_4083,N_3914,N_3693);
xor U4084 (N_4084,N_3928,N_3935);
or U4085 (N_4085,N_3732,N_3654);
nand U4086 (N_4086,N_3781,N_3972);
and U4087 (N_4087,N_3836,N_3859);
and U4088 (N_4088,N_3879,N_3510);
and U4089 (N_4089,N_3647,N_3964);
nand U4090 (N_4090,N_3750,N_3657);
nand U4091 (N_4091,N_3681,N_3894);
nand U4092 (N_4092,N_3890,N_3797);
or U4093 (N_4093,N_3982,N_3856);
and U4094 (N_4094,N_3737,N_3837);
and U4095 (N_4095,N_3819,N_3719);
or U4096 (N_4096,N_3762,N_3943);
or U4097 (N_4097,N_3883,N_3573);
nand U4098 (N_4098,N_3851,N_3658);
nor U4099 (N_4099,N_3969,N_3786);
and U4100 (N_4100,N_3643,N_3503);
nor U4101 (N_4101,N_3855,N_3653);
and U4102 (N_4102,N_3560,N_3872);
or U4103 (N_4103,N_3815,N_3871);
nor U4104 (N_4104,N_3822,N_3563);
and U4105 (N_4105,N_3551,N_3811);
or U4106 (N_4106,N_3747,N_3536);
nor U4107 (N_4107,N_3916,N_3893);
or U4108 (N_4108,N_3509,N_3963);
nor U4109 (N_4109,N_3939,N_3508);
nand U4110 (N_4110,N_3981,N_3930);
nor U4111 (N_4111,N_3741,N_3632);
and U4112 (N_4112,N_3541,N_3808);
nand U4113 (N_4113,N_3947,N_3901);
and U4114 (N_4114,N_3840,N_3556);
and U4115 (N_4115,N_3609,N_3727);
or U4116 (N_4116,N_3791,N_3785);
or U4117 (N_4117,N_3827,N_3718);
nand U4118 (N_4118,N_3881,N_3611);
nor U4119 (N_4119,N_3592,N_3940);
nand U4120 (N_4120,N_3692,N_3686);
and U4121 (N_4121,N_3814,N_3746);
nor U4122 (N_4122,N_3904,N_3717);
or U4123 (N_4123,N_3559,N_3902);
and U4124 (N_4124,N_3952,N_3804);
nand U4125 (N_4125,N_3586,N_3571);
and U4126 (N_4126,N_3670,N_3979);
nor U4127 (N_4127,N_3518,N_3899);
or U4128 (N_4128,N_3846,N_3809);
or U4129 (N_4129,N_3985,N_3587);
nand U4130 (N_4130,N_3993,N_3690);
nor U4131 (N_4131,N_3782,N_3744);
nand U4132 (N_4132,N_3900,N_3604);
and U4133 (N_4133,N_3694,N_3680);
or U4134 (N_4134,N_3545,N_3739);
nor U4135 (N_4135,N_3798,N_3554);
nand U4136 (N_4136,N_3803,N_3529);
nand U4137 (N_4137,N_3912,N_3721);
or U4138 (N_4138,N_3860,N_3829);
nand U4139 (N_4139,N_3678,N_3629);
and U4140 (N_4140,N_3652,N_3622);
and U4141 (N_4141,N_3886,N_3599);
nand U4142 (N_4142,N_3722,N_3787);
nand U4143 (N_4143,N_3569,N_3796);
or U4144 (N_4144,N_3504,N_3759);
nand U4145 (N_4145,N_3540,N_3511);
or U4146 (N_4146,N_3749,N_3882);
nor U4147 (N_4147,N_3588,N_3779);
or U4148 (N_4148,N_3677,N_3820);
nand U4149 (N_4149,N_3790,N_3695);
nor U4150 (N_4150,N_3568,N_3561);
nand U4151 (N_4151,N_3595,N_3714);
nand U4152 (N_4152,N_3887,N_3513);
or U4153 (N_4153,N_3748,N_3780);
nand U4154 (N_4154,N_3839,N_3898);
or U4155 (N_4155,N_3848,N_3712);
nor U4156 (N_4156,N_3601,N_3971);
and U4157 (N_4157,N_3842,N_3960);
or U4158 (N_4158,N_3506,N_3857);
or U4159 (N_4159,N_3770,N_3884);
nor U4160 (N_4160,N_3966,N_3801);
and U4161 (N_4161,N_3582,N_3615);
nand U4162 (N_4162,N_3897,N_3524);
or U4163 (N_4163,N_3821,N_3730);
nor U4164 (N_4164,N_3650,N_3537);
or U4165 (N_4165,N_3597,N_3557);
and U4166 (N_4166,N_3600,N_3661);
nand U4167 (N_4167,N_3666,N_3728);
nand U4168 (N_4168,N_3577,N_3740);
nand U4169 (N_4169,N_3555,N_3905);
nand U4170 (N_4170,N_3799,N_3683);
nand U4171 (N_4171,N_3775,N_3532);
or U4172 (N_4172,N_3825,N_3644);
nor U4173 (N_4173,N_3955,N_3519);
nor U4174 (N_4174,N_3521,N_3944);
or U4175 (N_4175,N_3729,N_3757);
nor U4176 (N_4176,N_3535,N_3823);
and U4177 (N_4177,N_3627,N_3933);
nand U4178 (N_4178,N_3742,N_3929);
or U4179 (N_4179,N_3865,N_3734);
nor U4180 (N_4180,N_3564,N_3907);
and U4181 (N_4181,N_3932,N_3614);
nand U4182 (N_4182,N_3672,N_3649);
nor U4183 (N_4183,N_3707,N_3709);
nor U4184 (N_4184,N_3957,N_3645);
nor U4185 (N_4185,N_3572,N_3716);
or U4186 (N_4186,N_3580,N_3591);
and U4187 (N_4187,N_3558,N_3593);
or U4188 (N_4188,N_3941,N_3628);
nor U4189 (N_4189,N_3565,N_3755);
and U4190 (N_4190,N_3915,N_3723);
nor U4191 (N_4191,N_3631,N_3936);
or U4192 (N_4192,N_3832,N_3926);
or U4193 (N_4193,N_3834,N_3651);
nor U4194 (N_4194,N_3642,N_3570);
nor U4195 (N_4195,N_3610,N_3769);
nand U4196 (N_4196,N_3575,N_3733);
or U4197 (N_4197,N_3976,N_3726);
or U4198 (N_4198,N_3705,N_3738);
nand U4199 (N_4199,N_3984,N_3682);
or U4200 (N_4200,N_3870,N_3636);
nor U4201 (N_4201,N_3720,N_3911);
nand U4202 (N_4202,N_3667,N_3853);
nor U4203 (N_4203,N_3874,N_3978);
and U4204 (N_4204,N_3635,N_3828);
nor U4205 (N_4205,N_3648,N_3965);
nand U4206 (N_4206,N_3675,N_3552);
and U4207 (N_4207,N_3973,N_3578);
or U4208 (N_4208,N_3619,N_3699);
nand U4209 (N_4209,N_3655,N_3697);
and U4210 (N_4210,N_3810,N_3816);
or U4211 (N_4211,N_3958,N_3713);
nor U4212 (N_4212,N_3951,N_3542);
nor U4213 (N_4213,N_3843,N_3664);
and U4214 (N_4214,N_3660,N_3962);
or U4215 (N_4215,N_3576,N_3774);
or U4216 (N_4216,N_3766,N_3530);
nand U4217 (N_4217,N_3752,N_3975);
nand U4218 (N_4218,N_3850,N_3594);
or U4219 (N_4219,N_3725,N_3613);
nand U4220 (N_4220,N_3987,N_3988);
or U4221 (N_4221,N_3583,N_3950);
xor U4222 (N_4222,N_3877,N_3585);
or U4223 (N_4223,N_3633,N_3659);
and U4224 (N_4224,N_3602,N_3812);
and U4225 (N_4225,N_3640,N_3869);
and U4226 (N_4226,N_3858,N_3679);
or U4227 (N_4227,N_3906,N_3876);
or U4228 (N_4228,N_3704,N_3621);
nand U4229 (N_4229,N_3923,N_3802);
or U4230 (N_4230,N_3795,N_3777);
nor U4231 (N_4231,N_3892,N_3862);
or U4232 (N_4232,N_3637,N_3543);
or U4233 (N_4233,N_3998,N_3961);
and U4234 (N_4234,N_3854,N_3581);
nor U4235 (N_4235,N_3546,N_3735);
nor U4236 (N_4236,N_3861,N_3668);
or U4237 (N_4237,N_3603,N_3620);
nand U4238 (N_4238,N_3625,N_3502);
xnor U4239 (N_4239,N_3919,N_3793);
or U4240 (N_4240,N_3873,N_3743);
nor U4241 (N_4241,N_3807,N_3547);
nor U4242 (N_4242,N_3778,N_3773);
and U4243 (N_4243,N_3867,N_3921);
or U4244 (N_4244,N_3806,N_3579);
nor U4245 (N_4245,N_3760,N_3833);
or U4246 (N_4246,N_3708,N_3500);
or U4247 (N_4247,N_3634,N_3847);
nor U4248 (N_4248,N_3956,N_3794);
nor U4249 (N_4249,N_3852,N_3792);
nor U4250 (N_4250,N_3869,N_3601);
and U4251 (N_4251,N_3941,N_3725);
and U4252 (N_4252,N_3809,N_3830);
and U4253 (N_4253,N_3879,N_3673);
and U4254 (N_4254,N_3728,N_3752);
or U4255 (N_4255,N_3795,N_3733);
nand U4256 (N_4256,N_3901,N_3586);
nand U4257 (N_4257,N_3949,N_3910);
nor U4258 (N_4258,N_3578,N_3600);
or U4259 (N_4259,N_3533,N_3834);
nand U4260 (N_4260,N_3648,N_3876);
and U4261 (N_4261,N_3607,N_3843);
nor U4262 (N_4262,N_3700,N_3960);
and U4263 (N_4263,N_3539,N_3963);
nor U4264 (N_4264,N_3814,N_3834);
nor U4265 (N_4265,N_3691,N_3746);
or U4266 (N_4266,N_3697,N_3978);
and U4267 (N_4267,N_3933,N_3706);
or U4268 (N_4268,N_3804,N_3524);
nand U4269 (N_4269,N_3845,N_3770);
and U4270 (N_4270,N_3773,N_3830);
and U4271 (N_4271,N_3983,N_3871);
nand U4272 (N_4272,N_3925,N_3581);
and U4273 (N_4273,N_3579,N_3551);
nand U4274 (N_4274,N_3774,N_3523);
nor U4275 (N_4275,N_3745,N_3526);
or U4276 (N_4276,N_3582,N_3575);
nand U4277 (N_4277,N_3701,N_3595);
or U4278 (N_4278,N_3761,N_3908);
nand U4279 (N_4279,N_3573,N_3515);
nand U4280 (N_4280,N_3787,N_3538);
nand U4281 (N_4281,N_3995,N_3881);
nand U4282 (N_4282,N_3739,N_3679);
nor U4283 (N_4283,N_3596,N_3765);
nand U4284 (N_4284,N_3840,N_3938);
or U4285 (N_4285,N_3976,N_3931);
or U4286 (N_4286,N_3508,N_3592);
or U4287 (N_4287,N_3868,N_3550);
and U4288 (N_4288,N_3690,N_3620);
nor U4289 (N_4289,N_3716,N_3814);
or U4290 (N_4290,N_3964,N_3962);
nand U4291 (N_4291,N_3719,N_3611);
nand U4292 (N_4292,N_3690,N_3760);
nor U4293 (N_4293,N_3675,N_3742);
nor U4294 (N_4294,N_3816,N_3684);
or U4295 (N_4295,N_3626,N_3511);
nor U4296 (N_4296,N_3945,N_3542);
nand U4297 (N_4297,N_3997,N_3948);
or U4298 (N_4298,N_3915,N_3705);
nor U4299 (N_4299,N_3769,N_3683);
and U4300 (N_4300,N_3968,N_3975);
nor U4301 (N_4301,N_3666,N_3931);
or U4302 (N_4302,N_3897,N_3817);
or U4303 (N_4303,N_3783,N_3614);
xnor U4304 (N_4304,N_3808,N_3542);
nand U4305 (N_4305,N_3645,N_3863);
and U4306 (N_4306,N_3979,N_3742);
or U4307 (N_4307,N_3960,N_3566);
and U4308 (N_4308,N_3936,N_3829);
and U4309 (N_4309,N_3982,N_3984);
nand U4310 (N_4310,N_3728,N_3799);
and U4311 (N_4311,N_3696,N_3682);
nor U4312 (N_4312,N_3901,N_3687);
nor U4313 (N_4313,N_3801,N_3518);
or U4314 (N_4314,N_3530,N_3653);
and U4315 (N_4315,N_3831,N_3590);
nor U4316 (N_4316,N_3513,N_3959);
nand U4317 (N_4317,N_3749,N_3767);
nand U4318 (N_4318,N_3652,N_3913);
and U4319 (N_4319,N_3936,N_3861);
and U4320 (N_4320,N_3926,N_3961);
nor U4321 (N_4321,N_3744,N_3931);
nor U4322 (N_4322,N_3964,N_3897);
nand U4323 (N_4323,N_3917,N_3502);
or U4324 (N_4324,N_3718,N_3858);
or U4325 (N_4325,N_3773,N_3967);
and U4326 (N_4326,N_3864,N_3729);
nand U4327 (N_4327,N_3636,N_3547);
and U4328 (N_4328,N_3604,N_3903);
or U4329 (N_4329,N_3720,N_3590);
or U4330 (N_4330,N_3530,N_3966);
nand U4331 (N_4331,N_3631,N_3834);
nor U4332 (N_4332,N_3569,N_3507);
and U4333 (N_4333,N_3636,N_3765);
or U4334 (N_4334,N_3577,N_3890);
nand U4335 (N_4335,N_3581,N_3928);
or U4336 (N_4336,N_3655,N_3917);
nor U4337 (N_4337,N_3981,N_3911);
nor U4338 (N_4338,N_3620,N_3524);
and U4339 (N_4339,N_3715,N_3676);
nand U4340 (N_4340,N_3913,N_3695);
nand U4341 (N_4341,N_3654,N_3834);
or U4342 (N_4342,N_3567,N_3739);
nor U4343 (N_4343,N_3876,N_3758);
nand U4344 (N_4344,N_3942,N_3783);
nand U4345 (N_4345,N_3919,N_3605);
and U4346 (N_4346,N_3946,N_3578);
nor U4347 (N_4347,N_3522,N_3918);
or U4348 (N_4348,N_3789,N_3529);
or U4349 (N_4349,N_3617,N_3994);
or U4350 (N_4350,N_3742,N_3553);
nand U4351 (N_4351,N_3676,N_3716);
or U4352 (N_4352,N_3619,N_3680);
and U4353 (N_4353,N_3909,N_3990);
and U4354 (N_4354,N_3808,N_3859);
or U4355 (N_4355,N_3654,N_3749);
and U4356 (N_4356,N_3533,N_3580);
nor U4357 (N_4357,N_3666,N_3689);
or U4358 (N_4358,N_3744,N_3504);
nand U4359 (N_4359,N_3842,N_3764);
nand U4360 (N_4360,N_3558,N_3806);
nand U4361 (N_4361,N_3567,N_3638);
nand U4362 (N_4362,N_3510,N_3987);
nor U4363 (N_4363,N_3868,N_3960);
and U4364 (N_4364,N_3545,N_3852);
nor U4365 (N_4365,N_3779,N_3855);
or U4366 (N_4366,N_3535,N_3517);
and U4367 (N_4367,N_3983,N_3744);
and U4368 (N_4368,N_3987,N_3574);
or U4369 (N_4369,N_3890,N_3883);
or U4370 (N_4370,N_3680,N_3788);
or U4371 (N_4371,N_3879,N_3768);
nand U4372 (N_4372,N_3663,N_3965);
nor U4373 (N_4373,N_3630,N_3650);
nor U4374 (N_4374,N_3765,N_3505);
and U4375 (N_4375,N_3686,N_3516);
nor U4376 (N_4376,N_3897,N_3799);
and U4377 (N_4377,N_3828,N_3928);
or U4378 (N_4378,N_3827,N_3801);
nand U4379 (N_4379,N_3701,N_3764);
or U4380 (N_4380,N_3528,N_3547);
nor U4381 (N_4381,N_3846,N_3875);
and U4382 (N_4382,N_3586,N_3980);
or U4383 (N_4383,N_3877,N_3835);
nor U4384 (N_4384,N_3777,N_3759);
or U4385 (N_4385,N_3926,N_3688);
or U4386 (N_4386,N_3896,N_3630);
nand U4387 (N_4387,N_3709,N_3624);
and U4388 (N_4388,N_3703,N_3935);
nand U4389 (N_4389,N_3816,N_3799);
and U4390 (N_4390,N_3540,N_3689);
nand U4391 (N_4391,N_3756,N_3666);
nand U4392 (N_4392,N_3823,N_3605);
nor U4393 (N_4393,N_3687,N_3954);
nor U4394 (N_4394,N_3845,N_3846);
nand U4395 (N_4395,N_3968,N_3730);
nand U4396 (N_4396,N_3861,N_3808);
nor U4397 (N_4397,N_3638,N_3819);
nand U4398 (N_4398,N_3846,N_3933);
or U4399 (N_4399,N_3542,N_3717);
and U4400 (N_4400,N_3773,N_3719);
and U4401 (N_4401,N_3572,N_3956);
nand U4402 (N_4402,N_3851,N_3902);
and U4403 (N_4403,N_3567,N_3730);
nor U4404 (N_4404,N_3730,N_3880);
and U4405 (N_4405,N_3792,N_3975);
nor U4406 (N_4406,N_3941,N_3518);
nor U4407 (N_4407,N_3875,N_3548);
nand U4408 (N_4408,N_3577,N_3747);
nand U4409 (N_4409,N_3551,N_3882);
or U4410 (N_4410,N_3633,N_3868);
nor U4411 (N_4411,N_3631,N_3975);
nor U4412 (N_4412,N_3822,N_3858);
or U4413 (N_4413,N_3966,N_3678);
nor U4414 (N_4414,N_3590,N_3626);
or U4415 (N_4415,N_3789,N_3574);
or U4416 (N_4416,N_3630,N_3966);
nor U4417 (N_4417,N_3624,N_3980);
xnor U4418 (N_4418,N_3840,N_3557);
nor U4419 (N_4419,N_3878,N_3524);
nor U4420 (N_4420,N_3757,N_3740);
and U4421 (N_4421,N_3804,N_3886);
nand U4422 (N_4422,N_3629,N_3624);
nor U4423 (N_4423,N_3726,N_3623);
and U4424 (N_4424,N_3786,N_3986);
or U4425 (N_4425,N_3807,N_3754);
nor U4426 (N_4426,N_3834,N_3912);
or U4427 (N_4427,N_3998,N_3666);
and U4428 (N_4428,N_3593,N_3942);
nand U4429 (N_4429,N_3990,N_3502);
or U4430 (N_4430,N_3531,N_3783);
nand U4431 (N_4431,N_3703,N_3986);
or U4432 (N_4432,N_3943,N_3509);
nand U4433 (N_4433,N_3661,N_3659);
nor U4434 (N_4434,N_3608,N_3760);
nor U4435 (N_4435,N_3565,N_3616);
or U4436 (N_4436,N_3563,N_3550);
nand U4437 (N_4437,N_3547,N_3560);
and U4438 (N_4438,N_3859,N_3582);
and U4439 (N_4439,N_3627,N_3514);
nand U4440 (N_4440,N_3657,N_3641);
nor U4441 (N_4441,N_3729,N_3754);
or U4442 (N_4442,N_3558,N_3654);
or U4443 (N_4443,N_3772,N_3883);
and U4444 (N_4444,N_3895,N_3752);
or U4445 (N_4445,N_3964,N_3715);
or U4446 (N_4446,N_3948,N_3638);
or U4447 (N_4447,N_3533,N_3859);
or U4448 (N_4448,N_3791,N_3546);
nand U4449 (N_4449,N_3750,N_3920);
nand U4450 (N_4450,N_3813,N_3870);
and U4451 (N_4451,N_3633,N_3806);
and U4452 (N_4452,N_3857,N_3727);
or U4453 (N_4453,N_3818,N_3962);
or U4454 (N_4454,N_3890,N_3662);
nor U4455 (N_4455,N_3957,N_3890);
nor U4456 (N_4456,N_3813,N_3641);
or U4457 (N_4457,N_3808,N_3594);
and U4458 (N_4458,N_3636,N_3743);
and U4459 (N_4459,N_3520,N_3968);
nand U4460 (N_4460,N_3630,N_3691);
nand U4461 (N_4461,N_3955,N_3740);
and U4462 (N_4462,N_3871,N_3826);
nand U4463 (N_4463,N_3627,N_3573);
and U4464 (N_4464,N_3826,N_3672);
or U4465 (N_4465,N_3719,N_3943);
or U4466 (N_4466,N_3740,N_3693);
xnor U4467 (N_4467,N_3894,N_3825);
and U4468 (N_4468,N_3644,N_3792);
or U4469 (N_4469,N_3859,N_3815);
nand U4470 (N_4470,N_3554,N_3748);
nand U4471 (N_4471,N_3677,N_3982);
and U4472 (N_4472,N_3623,N_3614);
and U4473 (N_4473,N_3803,N_3888);
nand U4474 (N_4474,N_3567,N_3980);
and U4475 (N_4475,N_3666,N_3516);
and U4476 (N_4476,N_3984,N_3641);
nand U4477 (N_4477,N_3608,N_3611);
or U4478 (N_4478,N_3514,N_3940);
or U4479 (N_4479,N_3994,N_3615);
nor U4480 (N_4480,N_3813,N_3696);
or U4481 (N_4481,N_3938,N_3603);
and U4482 (N_4482,N_3817,N_3871);
nand U4483 (N_4483,N_3511,N_3759);
nand U4484 (N_4484,N_3855,N_3528);
nor U4485 (N_4485,N_3673,N_3786);
or U4486 (N_4486,N_3894,N_3511);
or U4487 (N_4487,N_3651,N_3539);
nor U4488 (N_4488,N_3664,N_3934);
and U4489 (N_4489,N_3976,N_3844);
nand U4490 (N_4490,N_3546,N_3894);
and U4491 (N_4491,N_3705,N_3846);
and U4492 (N_4492,N_3917,N_3718);
nand U4493 (N_4493,N_3701,N_3789);
and U4494 (N_4494,N_3855,N_3660);
nor U4495 (N_4495,N_3742,N_3810);
nor U4496 (N_4496,N_3897,N_3681);
nand U4497 (N_4497,N_3775,N_3675);
nand U4498 (N_4498,N_3526,N_3634);
nand U4499 (N_4499,N_3816,N_3692);
nor U4500 (N_4500,N_4135,N_4174);
nor U4501 (N_4501,N_4103,N_4257);
nor U4502 (N_4502,N_4260,N_4142);
nand U4503 (N_4503,N_4352,N_4277);
and U4504 (N_4504,N_4356,N_4252);
nand U4505 (N_4505,N_4053,N_4253);
and U4506 (N_4506,N_4312,N_4293);
nand U4507 (N_4507,N_4242,N_4096);
or U4508 (N_4508,N_4362,N_4485);
nor U4509 (N_4509,N_4049,N_4063);
and U4510 (N_4510,N_4351,N_4000);
nand U4511 (N_4511,N_4061,N_4069);
nand U4512 (N_4512,N_4421,N_4296);
nor U4513 (N_4513,N_4249,N_4457);
nor U4514 (N_4514,N_4133,N_4112);
and U4515 (N_4515,N_4340,N_4004);
or U4516 (N_4516,N_4186,N_4466);
nand U4517 (N_4517,N_4192,N_4413);
and U4518 (N_4518,N_4393,N_4348);
and U4519 (N_4519,N_4084,N_4342);
and U4520 (N_4520,N_4355,N_4411);
and U4521 (N_4521,N_4073,N_4254);
nor U4522 (N_4522,N_4276,N_4006);
nor U4523 (N_4523,N_4415,N_4064);
nor U4524 (N_4524,N_4136,N_4450);
or U4525 (N_4525,N_4204,N_4095);
or U4526 (N_4526,N_4027,N_4202);
nand U4527 (N_4527,N_4106,N_4494);
and U4528 (N_4528,N_4427,N_4265);
or U4529 (N_4529,N_4247,N_4471);
nand U4530 (N_4530,N_4020,N_4057);
or U4531 (N_4531,N_4123,N_4217);
nor U4532 (N_4532,N_4469,N_4042);
and U4533 (N_4533,N_4041,N_4168);
and U4534 (N_4534,N_4177,N_4323);
and U4535 (N_4535,N_4270,N_4200);
and U4536 (N_4536,N_4250,N_4470);
or U4537 (N_4537,N_4132,N_4304);
nor U4538 (N_4538,N_4187,N_4325);
nor U4539 (N_4539,N_4286,N_4137);
or U4540 (N_4540,N_4279,N_4234);
nor U4541 (N_4541,N_4126,N_4374);
and U4542 (N_4542,N_4288,N_4266);
nand U4543 (N_4543,N_4213,N_4284);
or U4544 (N_4544,N_4237,N_4281);
nor U4545 (N_4545,N_4306,N_4321);
nor U4546 (N_4546,N_4206,N_4464);
or U4547 (N_4547,N_4332,N_4179);
nor U4548 (N_4548,N_4230,N_4129);
nand U4549 (N_4549,N_4045,N_4317);
or U4550 (N_4550,N_4181,N_4228);
nor U4551 (N_4551,N_4403,N_4369);
and U4552 (N_4552,N_4319,N_4259);
nor U4553 (N_4553,N_4046,N_4175);
nand U4554 (N_4554,N_4074,N_4017);
or U4555 (N_4555,N_4238,N_4387);
nor U4556 (N_4556,N_4327,N_4170);
xor U4557 (N_4557,N_4068,N_4191);
nand U4558 (N_4558,N_4113,N_4219);
xor U4559 (N_4559,N_4141,N_4377);
or U4560 (N_4560,N_4108,N_4039);
or U4561 (N_4561,N_4445,N_4368);
nor U4562 (N_4562,N_4493,N_4161);
or U4563 (N_4563,N_4302,N_4070);
or U4564 (N_4564,N_4489,N_4062);
and U4565 (N_4565,N_4067,N_4299);
nand U4566 (N_4566,N_4227,N_4184);
and U4567 (N_4567,N_4090,N_4468);
nor U4568 (N_4568,N_4243,N_4056);
or U4569 (N_4569,N_4373,N_4154);
nor U4570 (N_4570,N_4490,N_4205);
nor U4571 (N_4571,N_4498,N_4140);
or U4572 (N_4572,N_4122,N_4147);
or U4573 (N_4573,N_4367,N_4152);
nor U4574 (N_4574,N_4479,N_4245);
nand U4575 (N_4575,N_4310,N_4059);
nand U4576 (N_4576,N_4159,N_4436);
or U4577 (N_4577,N_4282,N_4400);
or U4578 (N_4578,N_4314,N_4207);
and U4579 (N_4579,N_4343,N_4385);
nand U4580 (N_4580,N_4478,N_4440);
nor U4581 (N_4581,N_4289,N_4088);
and U4582 (N_4582,N_4497,N_4496);
or U4583 (N_4583,N_4318,N_4405);
nand U4584 (N_4584,N_4475,N_4029);
nand U4585 (N_4585,N_4486,N_4109);
or U4586 (N_4586,N_4298,N_4320);
nand U4587 (N_4587,N_4264,N_4155);
and U4588 (N_4588,N_4392,N_4231);
nand U4589 (N_4589,N_4458,N_4297);
nand U4590 (N_4590,N_4402,N_4158);
nand U4591 (N_4591,N_4114,N_4051);
or U4592 (N_4592,N_4434,N_4290);
or U4593 (N_4593,N_4328,N_4417);
and U4594 (N_4594,N_4212,N_4223);
nand U4595 (N_4595,N_4262,N_4148);
nand U4596 (N_4596,N_4229,N_4087);
and U4597 (N_4597,N_4075,N_4216);
nand U4598 (N_4598,N_4308,N_4003);
or U4599 (N_4599,N_4214,N_4009);
or U4600 (N_4600,N_4366,N_4078);
or U4601 (N_4601,N_4337,N_4153);
nand U4602 (N_4602,N_4481,N_4345);
nand U4603 (N_4603,N_4022,N_4483);
or U4604 (N_4604,N_4050,N_4360);
nand U4605 (N_4605,N_4484,N_4097);
nor U4606 (N_4606,N_4072,N_4339);
nand U4607 (N_4607,N_4165,N_4433);
or U4608 (N_4608,N_4294,N_4083);
or U4609 (N_4609,N_4156,N_4431);
nand U4610 (N_4610,N_4472,N_4295);
nand U4611 (N_4611,N_4491,N_4305);
nand U4612 (N_4612,N_4026,N_4447);
nand U4613 (N_4613,N_4086,N_4363);
nor U4614 (N_4614,N_4410,N_4397);
nand U4615 (N_4615,N_4409,N_4394);
nand U4616 (N_4616,N_4380,N_4128);
and U4617 (N_4617,N_4467,N_4338);
nor U4618 (N_4618,N_4210,N_4438);
nand U4619 (N_4619,N_4169,N_4364);
nand U4620 (N_4620,N_4199,N_4024);
and U4621 (N_4621,N_4261,N_4221);
and U4622 (N_4622,N_4193,N_4019);
nor U4623 (N_4623,N_4442,N_4031);
or U4624 (N_4624,N_4033,N_4335);
or U4625 (N_4625,N_4111,N_4058);
and U4626 (N_4626,N_4150,N_4025);
and U4627 (N_4627,N_4182,N_4085);
or U4628 (N_4628,N_4383,N_4256);
and U4629 (N_4629,N_4370,N_4435);
or U4630 (N_4630,N_4418,N_4273);
nand U4631 (N_4631,N_4016,N_4118);
and U4632 (N_4632,N_4007,N_4315);
or U4633 (N_4633,N_4336,N_4313);
nand U4634 (N_4634,N_4190,N_4149);
or U4635 (N_4635,N_4124,N_4303);
nand U4636 (N_4636,N_4071,N_4121);
nand U4637 (N_4637,N_4399,N_4038);
nor U4638 (N_4638,N_4350,N_4251);
and U4639 (N_4639,N_4263,N_4396);
nand U4640 (N_4640,N_4301,N_4198);
and U4641 (N_4641,N_4218,N_4384);
or U4642 (N_4642,N_4163,N_4185);
nor U4643 (N_4643,N_4349,N_4480);
and U4644 (N_4644,N_4171,N_4089);
nand U4645 (N_4645,N_4180,N_4422);
nor U4646 (N_4646,N_4102,N_4167);
nor U4647 (N_4647,N_4116,N_4379);
or U4648 (N_4648,N_4201,N_4376);
and U4649 (N_4649,N_4462,N_4011);
nand U4650 (N_4650,N_4215,N_4131);
and U4651 (N_4651,N_4292,N_4082);
nand U4652 (N_4652,N_4188,N_4178);
or U4653 (N_4653,N_4398,N_4424);
nand U4654 (N_4654,N_4115,N_4439);
nand U4655 (N_4655,N_4454,N_4287);
or U4656 (N_4656,N_4414,N_4101);
nand U4657 (N_4657,N_4010,N_4117);
or U4658 (N_4658,N_4425,N_4423);
nor U4659 (N_4659,N_4081,N_4119);
nand U4660 (N_4660,N_4048,N_4334);
nor U4661 (N_4661,N_4278,N_4382);
nand U4662 (N_4662,N_4280,N_4331);
nor U4663 (N_4663,N_4066,N_4144);
nor U4664 (N_4664,N_4477,N_4138);
nand U4665 (N_4665,N_4034,N_4455);
and U4666 (N_4666,N_4134,N_4104);
and U4667 (N_4667,N_4499,N_4333);
nor U4668 (N_4668,N_4463,N_4021);
nor U4669 (N_4669,N_4151,N_4437);
and U4670 (N_4670,N_4145,N_4269);
or U4671 (N_4671,N_4065,N_4488);
or U4672 (N_4672,N_4209,N_4419);
nor U4673 (N_4673,N_4143,N_4446);
and U4674 (N_4674,N_4372,N_4125);
and U4675 (N_4675,N_4358,N_4459);
nor U4676 (N_4676,N_4222,N_4271);
or U4677 (N_4677,N_4040,N_4401);
nor U4678 (N_4678,N_4473,N_4487);
nand U4679 (N_4679,N_4015,N_4449);
xnor U4680 (N_4680,N_4316,N_4091);
or U4681 (N_4681,N_4157,N_4420);
or U4682 (N_4682,N_4324,N_4211);
nand U4683 (N_4683,N_4375,N_4311);
nand U4684 (N_4684,N_4404,N_4241);
nor U4685 (N_4685,N_4030,N_4307);
nor U4686 (N_4686,N_4052,N_4233);
nand U4687 (N_4687,N_4274,N_4285);
nor U4688 (N_4688,N_4098,N_4130);
nand U4689 (N_4689,N_4093,N_4407);
and U4690 (N_4690,N_4291,N_4002);
nor U4691 (N_4691,N_4461,N_4441);
and U4692 (N_4692,N_4060,N_4054);
or U4693 (N_4693,N_4023,N_4267);
or U4694 (N_4694,N_4452,N_4244);
and U4695 (N_4695,N_4428,N_4354);
and U4696 (N_4696,N_4197,N_4208);
nand U4697 (N_4697,N_4395,N_4239);
and U4698 (N_4698,N_4357,N_4035);
or U4699 (N_4699,N_4482,N_4196);
nor U4700 (N_4700,N_4176,N_4326);
nor U4701 (N_4701,N_4235,N_4258);
nor U4702 (N_4702,N_4094,N_4347);
and U4703 (N_4703,N_4160,N_4460);
nand U4704 (N_4704,N_4353,N_4139);
nand U4705 (N_4705,N_4448,N_4172);
xor U4706 (N_4706,N_4224,N_4028);
nand U4707 (N_4707,N_4162,N_4389);
or U4708 (N_4708,N_4300,N_4365);
nor U4709 (N_4709,N_4476,N_4344);
or U4710 (N_4710,N_4341,N_4120);
and U4711 (N_4711,N_4391,N_4001);
or U4712 (N_4712,N_4195,N_4189);
xor U4713 (N_4713,N_4248,N_4465);
nand U4714 (N_4714,N_4164,N_4426);
nor U4715 (N_4715,N_4107,N_4008);
or U4716 (N_4716,N_4005,N_4386);
nor U4717 (N_4717,N_4080,N_4443);
or U4718 (N_4718,N_4329,N_4432);
nor U4719 (N_4719,N_4127,N_4346);
or U4720 (N_4720,N_4225,N_4076);
nand U4721 (N_4721,N_4378,N_4236);
nand U4722 (N_4722,N_4272,N_4203);
or U4723 (N_4723,N_4013,N_4246);
or U4724 (N_4724,N_4330,N_4444);
and U4725 (N_4725,N_4412,N_4408);
or U4726 (N_4726,N_4268,N_4220);
nand U4727 (N_4727,N_4453,N_4240);
and U4728 (N_4728,N_4429,N_4043);
nor U4729 (N_4729,N_4255,N_4381);
and U4730 (N_4730,N_4146,N_4012);
nand U4731 (N_4731,N_4416,N_4232);
nand U4732 (N_4732,N_4044,N_4014);
or U4733 (N_4733,N_4055,N_4166);
nor U4734 (N_4734,N_4037,N_4079);
nor U4735 (N_4735,N_4105,N_4099);
and U4736 (N_4736,N_4100,N_4018);
and U4737 (N_4737,N_4283,N_4092);
and U4738 (N_4738,N_4036,N_4275);
and U4739 (N_4739,N_4032,N_4309);
and U4740 (N_4740,N_4110,N_4047);
and U4741 (N_4741,N_4430,N_4361);
nand U4742 (N_4742,N_4173,N_4388);
nor U4743 (N_4743,N_4474,N_4183);
or U4744 (N_4744,N_4456,N_4322);
nand U4745 (N_4745,N_4194,N_4492);
or U4746 (N_4746,N_4359,N_4406);
nor U4747 (N_4747,N_4226,N_4390);
nand U4748 (N_4748,N_4371,N_4451);
nor U4749 (N_4749,N_4077,N_4495);
nor U4750 (N_4750,N_4372,N_4342);
nand U4751 (N_4751,N_4284,N_4348);
xor U4752 (N_4752,N_4380,N_4284);
nor U4753 (N_4753,N_4050,N_4263);
nand U4754 (N_4754,N_4476,N_4211);
nor U4755 (N_4755,N_4049,N_4148);
and U4756 (N_4756,N_4486,N_4343);
nor U4757 (N_4757,N_4184,N_4249);
or U4758 (N_4758,N_4005,N_4248);
nand U4759 (N_4759,N_4424,N_4466);
nand U4760 (N_4760,N_4419,N_4439);
or U4761 (N_4761,N_4450,N_4182);
nand U4762 (N_4762,N_4012,N_4477);
and U4763 (N_4763,N_4301,N_4333);
nor U4764 (N_4764,N_4044,N_4155);
and U4765 (N_4765,N_4156,N_4288);
nor U4766 (N_4766,N_4438,N_4081);
nand U4767 (N_4767,N_4321,N_4465);
nor U4768 (N_4768,N_4120,N_4000);
nor U4769 (N_4769,N_4336,N_4181);
nand U4770 (N_4770,N_4379,N_4000);
nand U4771 (N_4771,N_4259,N_4088);
nor U4772 (N_4772,N_4254,N_4386);
nand U4773 (N_4773,N_4157,N_4106);
nand U4774 (N_4774,N_4205,N_4086);
nor U4775 (N_4775,N_4470,N_4091);
nand U4776 (N_4776,N_4106,N_4199);
nand U4777 (N_4777,N_4198,N_4327);
nand U4778 (N_4778,N_4315,N_4070);
nand U4779 (N_4779,N_4205,N_4030);
nand U4780 (N_4780,N_4303,N_4335);
and U4781 (N_4781,N_4023,N_4108);
or U4782 (N_4782,N_4161,N_4184);
xnor U4783 (N_4783,N_4092,N_4091);
and U4784 (N_4784,N_4374,N_4192);
and U4785 (N_4785,N_4346,N_4066);
and U4786 (N_4786,N_4057,N_4310);
nor U4787 (N_4787,N_4057,N_4427);
nor U4788 (N_4788,N_4461,N_4373);
and U4789 (N_4789,N_4089,N_4485);
and U4790 (N_4790,N_4161,N_4373);
nor U4791 (N_4791,N_4208,N_4493);
and U4792 (N_4792,N_4047,N_4337);
and U4793 (N_4793,N_4399,N_4339);
and U4794 (N_4794,N_4216,N_4107);
nand U4795 (N_4795,N_4072,N_4203);
nor U4796 (N_4796,N_4068,N_4460);
nor U4797 (N_4797,N_4016,N_4193);
nand U4798 (N_4798,N_4474,N_4043);
nand U4799 (N_4799,N_4460,N_4021);
nor U4800 (N_4800,N_4314,N_4218);
nor U4801 (N_4801,N_4444,N_4185);
nor U4802 (N_4802,N_4399,N_4079);
or U4803 (N_4803,N_4121,N_4208);
or U4804 (N_4804,N_4454,N_4034);
nand U4805 (N_4805,N_4167,N_4191);
and U4806 (N_4806,N_4036,N_4028);
and U4807 (N_4807,N_4444,N_4280);
or U4808 (N_4808,N_4143,N_4322);
and U4809 (N_4809,N_4177,N_4115);
nand U4810 (N_4810,N_4020,N_4216);
or U4811 (N_4811,N_4405,N_4378);
and U4812 (N_4812,N_4084,N_4074);
and U4813 (N_4813,N_4405,N_4074);
nor U4814 (N_4814,N_4080,N_4314);
and U4815 (N_4815,N_4111,N_4381);
and U4816 (N_4816,N_4348,N_4447);
nor U4817 (N_4817,N_4240,N_4335);
or U4818 (N_4818,N_4056,N_4329);
nor U4819 (N_4819,N_4014,N_4045);
and U4820 (N_4820,N_4040,N_4086);
nor U4821 (N_4821,N_4095,N_4217);
nor U4822 (N_4822,N_4411,N_4292);
nand U4823 (N_4823,N_4138,N_4113);
nor U4824 (N_4824,N_4251,N_4492);
nor U4825 (N_4825,N_4433,N_4077);
nand U4826 (N_4826,N_4088,N_4439);
nand U4827 (N_4827,N_4107,N_4039);
nand U4828 (N_4828,N_4337,N_4144);
nand U4829 (N_4829,N_4089,N_4024);
and U4830 (N_4830,N_4332,N_4162);
or U4831 (N_4831,N_4051,N_4071);
and U4832 (N_4832,N_4301,N_4428);
or U4833 (N_4833,N_4350,N_4484);
nand U4834 (N_4834,N_4130,N_4024);
nand U4835 (N_4835,N_4021,N_4496);
nor U4836 (N_4836,N_4100,N_4050);
or U4837 (N_4837,N_4138,N_4191);
and U4838 (N_4838,N_4197,N_4353);
or U4839 (N_4839,N_4312,N_4078);
or U4840 (N_4840,N_4257,N_4297);
or U4841 (N_4841,N_4247,N_4478);
nand U4842 (N_4842,N_4351,N_4027);
or U4843 (N_4843,N_4184,N_4304);
or U4844 (N_4844,N_4116,N_4272);
and U4845 (N_4845,N_4189,N_4421);
nor U4846 (N_4846,N_4156,N_4202);
nand U4847 (N_4847,N_4236,N_4465);
or U4848 (N_4848,N_4274,N_4464);
and U4849 (N_4849,N_4349,N_4385);
nand U4850 (N_4850,N_4031,N_4291);
nor U4851 (N_4851,N_4025,N_4015);
nand U4852 (N_4852,N_4437,N_4451);
and U4853 (N_4853,N_4421,N_4346);
and U4854 (N_4854,N_4363,N_4160);
nor U4855 (N_4855,N_4366,N_4370);
and U4856 (N_4856,N_4445,N_4493);
nand U4857 (N_4857,N_4172,N_4496);
nor U4858 (N_4858,N_4006,N_4281);
and U4859 (N_4859,N_4218,N_4251);
or U4860 (N_4860,N_4237,N_4498);
and U4861 (N_4861,N_4017,N_4483);
and U4862 (N_4862,N_4040,N_4426);
or U4863 (N_4863,N_4422,N_4306);
or U4864 (N_4864,N_4250,N_4308);
or U4865 (N_4865,N_4200,N_4185);
or U4866 (N_4866,N_4046,N_4319);
and U4867 (N_4867,N_4215,N_4030);
or U4868 (N_4868,N_4387,N_4233);
nand U4869 (N_4869,N_4231,N_4009);
and U4870 (N_4870,N_4258,N_4114);
nand U4871 (N_4871,N_4074,N_4338);
nor U4872 (N_4872,N_4206,N_4312);
nor U4873 (N_4873,N_4290,N_4343);
nor U4874 (N_4874,N_4461,N_4128);
and U4875 (N_4875,N_4076,N_4025);
or U4876 (N_4876,N_4024,N_4316);
or U4877 (N_4877,N_4476,N_4373);
nand U4878 (N_4878,N_4412,N_4402);
and U4879 (N_4879,N_4357,N_4260);
nor U4880 (N_4880,N_4031,N_4262);
nor U4881 (N_4881,N_4429,N_4036);
nand U4882 (N_4882,N_4426,N_4467);
or U4883 (N_4883,N_4370,N_4401);
and U4884 (N_4884,N_4169,N_4193);
and U4885 (N_4885,N_4252,N_4342);
nor U4886 (N_4886,N_4465,N_4117);
xnor U4887 (N_4887,N_4006,N_4185);
and U4888 (N_4888,N_4074,N_4174);
nor U4889 (N_4889,N_4018,N_4218);
and U4890 (N_4890,N_4127,N_4147);
nor U4891 (N_4891,N_4045,N_4398);
nor U4892 (N_4892,N_4475,N_4336);
nor U4893 (N_4893,N_4482,N_4027);
or U4894 (N_4894,N_4106,N_4335);
nor U4895 (N_4895,N_4376,N_4332);
or U4896 (N_4896,N_4356,N_4317);
xor U4897 (N_4897,N_4312,N_4162);
or U4898 (N_4898,N_4062,N_4119);
nor U4899 (N_4899,N_4087,N_4481);
xnor U4900 (N_4900,N_4072,N_4307);
xnor U4901 (N_4901,N_4458,N_4419);
or U4902 (N_4902,N_4339,N_4168);
and U4903 (N_4903,N_4446,N_4433);
and U4904 (N_4904,N_4133,N_4371);
and U4905 (N_4905,N_4335,N_4242);
or U4906 (N_4906,N_4310,N_4017);
nand U4907 (N_4907,N_4095,N_4198);
nor U4908 (N_4908,N_4293,N_4135);
and U4909 (N_4909,N_4147,N_4457);
nand U4910 (N_4910,N_4355,N_4020);
nand U4911 (N_4911,N_4367,N_4160);
nor U4912 (N_4912,N_4158,N_4456);
nand U4913 (N_4913,N_4308,N_4083);
nand U4914 (N_4914,N_4477,N_4107);
and U4915 (N_4915,N_4003,N_4076);
and U4916 (N_4916,N_4060,N_4281);
nand U4917 (N_4917,N_4102,N_4393);
nor U4918 (N_4918,N_4198,N_4377);
or U4919 (N_4919,N_4298,N_4015);
or U4920 (N_4920,N_4182,N_4173);
and U4921 (N_4921,N_4065,N_4120);
or U4922 (N_4922,N_4211,N_4399);
and U4923 (N_4923,N_4402,N_4049);
or U4924 (N_4924,N_4136,N_4251);
and U4925 (N_4925,N_4347,N_4114);
nor U4926 (N_4926,N_4136,N_4342);
nand U4927 (N_4927,N_4334,N_4188);
nor U4928 (N_4928,N_4363,N_4217);
or U4929 (N_4929,N_4436,N_4209);
and U4930 (N_4930,N_4305,N_4347);
and U4931 (N_4931,N_4477,N_4446);
nor U4932 (N_4932,N_4175,N_4406);
nand U4933 (N_4933,N_4493,N_4463);
or U4934 (N_4934,N_4248,N_4112);
and U4935 (N_4935,N_4417,N_4062);
nor U4936 (N_4936,N_4090,N_4079);
nand U4937 (N_4937,N_4285,N_4381);
nor U4938 (N_4938,N_4143,N_4157);
nand U4939 (N_4939,N_4059,N_4144);
nor U4940 (N_4940,N_4490,N_4459);
nand U4941 (N_4941,N_4190,N_4198);
and U4942 (N_4942,N_4167,N_4377);
or U4943 (N_4943,N_4218,N_4169);
and U4944 (N_4944,N_4444,N_4089);
and U4945 (N_4945,N_4273,N_4434);
and U4946 (N_4946,N_4008,N_4458);
nor U4947 (N_4947,N_4284,N_4095);
nand U4948 (N_4948,N_4254,N_4420);
xnor U4949 (N_4949,N_4368,N_4096);
or U4950 (N_4950,N_4480,N_4301);
and U4951 (N_4951,N_4314,N_4266);
or U4952 (N_4952,N_4120,N_4133);
nand U4953 (N_4953,N_4184,N_4136);
and U4954 (N_4954,N_4369,N_4161);
or U4955 (N_4955,N_4275,N_4474);
and U4956 (N_4956,N_4057,N_4180);
or U4957 (N_4957,N_4317,N_4459);
nand U4958 (N_4958,N_4259,N_4478);
nand U4959 (N_4959,N_4196,N_4218);
nor U4960 (N_4960,N_4157,N_4232);
or U4961 (N_4961,N_4353,N_4096);
nor U4962 (N_4962,N_4034,N_4021);
or U4963 (N_4963,N_4436,N_4257);
and U4964 (N_4964,N_4297,N_4324);
nor U4965 (N_4965,N_4413,N_4440);
and U4966 (N_4966,N_4363,N_4423);
and U4967 (N_4967,N_4298,N_4042);
nand U4968 (N_4968,N_4406,N_4418);
or U4969 (N_4969,N_4213,N_4343);
or U4970 (N_4970,N_4157,N_4293);
nor U4971 (N_4971,N_4168,N_4394);
nand U4972 (N_4972,N_4125,N_4263);
or U4973 (N_4973,N_4292,N_4440);
and U4974 (N_4974,N_4287,N_4137);
nor U4975 (N_4975,N_4090,N_4199);
nand U4976 (N_4976,N_4105,N_4165);
nand U4977 (N_4977,N_4207,N_4437);
or U4978 (N_4978,N_4432,N_4164);
nand U4979 (N_4979,N_4466,N_4372);
or U4980 (N_4980,N_4360,N_4113);
nand U4981 (N_4981,N_4113,N_4422);
nor U4982 (N_4982,N_4019,N_4138);
nand U4983 (N_4983,N_4312,N_4445);
nor U4984 (N_4984,N_4311,N_4129);
or U4985 (N_4985,N_4136,N_4446);
nor U4986 (N_4986,N_4030,N_4044);
and U4987 (N_4987,N_4432,N_4298);
nor U4988 (N_4988,N_4381,N_4196);
nor U4989 (N_4989,N_4235,N_4403);
nor U4990 (N_4990,N_4281,N_4249);
and U4991 (N_4991,N_4352,N_4279);
and U4992 (N_4992,N_4094,N_4424);
and U4993 (N_4993,N_4369,N_4126);
nor U4994 (N_4994,N_4018,N_4457);
and U4995 (N_4995,N_4463,N_4006);
nor U4996 (N_4996,N_4488,N_4052);
nor U4997 (N_4997,N_4354,N_4102);
nand U4998 (N_4998,N_4188,N_4019);
nand U4999 (N_4999,N_4342,N_4002);
or UO_0 (O_0,N_4704,N_4862);
nand UO_1 (O_1,N_4569,N_4831);
or UO_2 (O_2,N_4891,N_4906);
nor UO_3 (O_3,N_4757,N_4624);
nand UO_4 (O_4,N_4746,N_4881);
or UO_5 (O_5,N_4965,N_4604);
nor UO_6 (O_6,N_4567,N_4660);
or UO_7 (O_7,N_4824,N_4713);
nand UO_8 (O_8,N_4783,N_4555);
or UO_9 (O_9,N_4806,N_4989);
and UO_10 (O_10,N_4932,N_4759);
or UO_11 (O_11,N_4724,N_4728);
nor UO_12 (O_12,N_4751,N_4793);
and UO_13 (O_13,N_4636,N_4692);
and UO_14 (O_14,N_4639,N_4694);
or UO_15 (O_15,N_4651,N_4707);
or UO_16 (O_16,N_4761,N_4556);
nand UO_17 (O_17,N_4633,N_4655);
nor UO_18 (O_18,N_4517,N_4538);
nand UO_19 (O_19,N_4928,N_4672);
nor UO_20 (O_20,N_4661,N_4869);
nor UO_21 (O_21,N_4777,N_4947);
nor UO_22 (O_22,N_4948,N_4966);
and UO_23 (O_23,N_4668,N_4587);
or UO_24 (O_24,N_4962,N_4852);
nor UO_25 (O_25,N_4986,N_4585);
nand UO_26 (O_26,N_4836,N_4542);
nand UO_27 (O_27,N_4853,N_4586);
or UO_28 (O_28,N_4877,N_4580);
nand UO_29 (O_29,N_4848,N_4764);
or UO_30 (O_30,N_4969,N_4863);
and UO_31 (O_31,N_4916,N_4794);
nand UO_32 (O_32,N_4894,N_4755);
nand UO_33 (O_33,N_4768,N_4611);
or UO_34 (O_34,N_4758,N_4994);
nand UO_35 (O_35,N_4914,N_4696);
nor UO_36 (O_36,N_4892,N_4533);
nand UO_37 (O_37,N_4987,N_4921);
xor UO_38 (O_38,N_4695,N_4875);
nor UO_39 (O_39,N_4900,N_4539);
nor UO_40 (O_40,N_4945,N_4572);
or UO_41 (O_41,N_4792,N_4804);
nor UO_42 (O_42,N_4521,N_4674);
nor UO_43 (O_43,N_4664,N_4647);
or UO_44 (O_44,N_4573,N_4646);
and UO_45 (O_45,N_4977,N_4609);
and UO_46 (O_46,N_4529,N_4748);
or UO_47 (O_47,N_4690,N_4844);
and UO_48 (O_48,N_4870,N_4558);
nand UO_49 (O_49,N_4920,N_4599);
or UO_50 (O_50,N_4548,N_4910);
and UO_51 (O_51,N_4665,N_4918);
nor UO_52 (O_52,N_4867,N_4562);
nor UO_53 (O_53,N_4929,N_4712);
or UO_54 (O_54,N_4574,N_4973);
or UO_55 (O_55,N_4709,N_4710);
xor UO_56 (O_56,N_4503,N_4830);
and UO_57 (O_57,N_4559,N_4508);
nor UO_58 (O_58,N_4524,N_4765);
and UO_59 (O_59,N_4640,N_4941);
or UO_60 (O_60,N_4922,N_4782);
or UO_61 (O_61,N_4780,N_4882);
nand UO_62 (O_62,N_4718,N_4700);
nand UO_63 (O_63,N_4752,N_4741);
nand UO_64 (O_64,N_4807,N_4545);
or UO_65 (O_65,N_4818,N_4543);
and UO_66 (O_66,N_4846,N_4607);
nand UO_67 (O_67,N_4630,N_4974);
or UO_68 (O_68,N_4978,N_4519);
and UO_69 (O_69,N_4618,N_4887);
nor UO_70 (O_70,N_4589,N_4554);
and UO_71 (O_71,N_4591,N_4971);
and UO_72 (O_72,N_4808,N_4682);
or UO_73 (O_73,N_4801,N_4854);
nor UO_74 (O_74,N_4512,N_4522);
or UO_75 (O_75,N_4619,N_4934);
or UO_76 (O_76,N_4841,N_4845);
nor UO_77 (O_77,N_4731,N_4735);
nor UO_78 (O_78,N_4851,N_4739);
or UO_79 (O_79,N_4884,N_4866);
and UO_80 (O_80,N_4504,N_4871);
nand UO_81 (O_81,N_4507,N_4738);
and UO_82 (O_82,N_4627,N_4924);
or UO_83 (O_83,N_4581,N_4776);
or UO_84 (O_84,N_4600,N_4826);
nand UO_85 (O_85,N_4528,N_4642);
and UO_86 (O_86,N_4859,N_4822);
or UO_87 (O_87,N_4530,N_4925);
nand UO_88 (O_88,N_4985,N_4702);
and UO_89 (O_89,N_4850,N_4975);
or UO_90 (O_90,N_4769,N_4720);
nor UO_91 (O_91,N_4886,N_4608);
nor UO_92 (O_92,N_4904,N_4502);
nor UO_93 (O_93,N_4798,N_4963);
and UO_94 (O_94,N_4744,N_4896);
or UO_95 (O_95,N_4880,N_4876);
nor UO_96 (O_96,N_4775,N_4899);
and UO_97 (O_97,N_4706,N_4595);
nor UO_98 (O_98,N_4737,N_4897);
and UO_99 (O_99,N_4520,N_4957);
and UO_100 (O_100,N_4961,N_4726);
nor UO_101 (O_101,N_4908,N_4756);
nand UO_102 (O_102,N_4685,N_4536);
or UO_103 (O_103,N_4983,N_4729);
and UO_104 (O_104,N_4805,N_4617);
nand UO_105 (O_105,N_4641,N_4500);
nand UO_106 (O_106,N_4570,N_4864);
and UO_107 (O_107,N_4679,N_4677);
and UO_108 (O_108,N_4721,N_4571);
nor UO_109 (O_109,N_4960,N_4635);
nand UO_110 (O_110,N_4861,N_4733);
and UO_111 (O_111,N_4820,N_4849);
nand UO_112 (O_112,N_4628,N_4631);
nand UO_113 (O_113,N_4763,N_4708);
or UO_114 (O_114,N_4936,N_4791);
nand UO_115 (O_115,N_4509,N_4950);
and UO_116 (O_116,N_4693,N_4614);
or UO_117 (O_117,N_4858,N_4909);
nand UO_118 (O_118,N_4691,N_4515);
nand UO_119 (O_119,N_4550,N_4847);
or UO_120 (O_120,N_4903,N_4905);
nand UO_121 (O_121,N_4557,N_4680);
nor UO_122 (O_122,N_4937,N_4547);
nand UO_123 (O_123,N_4955,N_4993);
nand UO_124 (O_124,N_4531,N_4800);
and UO_125 (O_125,N_4514,N_4988);
nand UO_126 (O_126,N_4964,N_4926);
nor UO_127 (O_127,N_4781,N_4927);
nor UO_128 (O_128,N_4666,N_4774);
and UO_129 (O_129,N_4566,N_4885);
nor UO_130 (O_130,N_4770,N_4879);
nand UO_131 (O_131,N_4659,N_4883);
nor UO_132 (O_132,N_4865,N_4564);
nand UO_133 (O_133,N_4546,N_4812);
nor UO_134 (O_134,N_4603,N_4827);
nor UO_135 (O_135,N_4513,N_4995);
and UO_136 (O_136,N_4938,N_4687);
nand UO_137 (O_137,N_4943,N_4578);
or UO_138 (O_138,N_4576,N_4760);
nand UO_139 (O_139,N_4742,N_4874);
nand UO_140 (O_140,N_4681,N_4915);
or UO_141 (O_141,N_4772,N_4953);
nor UO_142 (O_142,N_4951,N_4992);
nor UO_143 (O_143,N_4670,N_4810);
nor UO_144 (O_144,N_4590,N_4982);
or UO_145 (O_145,N_4518,N_4942);
nand UO_146 (O_146,N_4823,N_4549);
nor UO_147 (O_147,N_4623,N_4819);
and UO_148 (O_148,N_4563,N_4779);
nand UO_149 (O_149,N_4786,N_4778);
and UO_150 (O_150,N_4996,N_4855);
or UO_151 (O_151,N_4568,N_4825);
nand UO_152 (O_152,N_4584,N_4582);
and UO_153 (O_153,N_4832,N_4967);
and UO_154 (O_154,N_4727,N_4814);
nand UO_155 (O_155,N_4809,N_4597);
nor UO_156 (O_156,N_4663,N_4997);
and UO_157 (O_157,N_4911,N_4616);
nand UO_158 (O_158,N_4979,N_4923);
nor UO_159 (O_159,N_4534,N_4613);
and UO_160 (O_160,N_4753,N_4560);
nand UO_161 (O_161,N_4817,N_4610);
and UO_162 (O_162,N_4723,N_4544);
and UO_163 (O_163,N_4771,N_4889);
nand UO_164 (O_164,N_4671,N_4821);
nand UO_165 (O_165,N_4816,N_4552);
or UO_166 (O_166,N_4537,N_4698);
and UO_167 (O_167,N_4583,N_4784);
nor UO_168 (O_168,N_4526,N_4605);
nor UO_169 (O_169,N_4675,N_4888);
or UO_170 (O_170,N_4743,N_4991);
and UO_171 (O_171,N_4593,N_4648);
or UO_172 (O_172,N_4541,N_4510);
or UO_173 (O_173,N_4873,N_4754);
nor UO_174 (O_174,N_4952,N_4703);
and UO_175 (O_175,N_4717,N_4787);
and UO_176 (O_176,N_4652,N_4990);
nor UO_177 (O_177,N_4634,N_4688);
or UO_178 (O_178,N_4622,N_4829);
or UO_179 (O_179,N_4676,N_4621);
and UO_180 (O_180,N_4868,N_4740);
and UO_181 (O_181,N_4762,N_4656);
or UO_182 (O_182,N_4615,N_4683);
and UO_183 (O_183,N_4797,N_4940);
nand UO_184 (O_184,N_4535,N_4697);
nor UO_185 (O_185,N_4767,N_4840);
nand UO_186 (O_186,N_4523,N_4669);
nor UO_187 (O_187,N_4912,N_4984);
nor UO_188 (O_188,N_4980,N_4790);
nand UO_189 (O_189,N_4629,N_4872);
nand UO_190 (O_190,N_4745,N_4959);
and UO_191 (O_191,N_4860,N_4540);
or UO_192 (O_192,N_4917,N_4699);
and UO_193 (O_193,N_4701,N_4588);
nand UO_194 (O_194,N_4838,N_4898);
nand UO_195 (O_195,N_4785,N_4795);
or UO_196 (O_196,N_4750,N_4525);
or UO_197 (O_197,N_4946,N_4653);
and UO_198 (O_198,N_4592,N_4833);
nand UO_199 (O_199,N_4725,N_4913);
or UO_200 (O_200,N_4714,N_4901);
and UO_201 (O_201,N_4893,N_4976);
or UO_202 (O_202,N_4902,N_4970);
nand UO_203 (O_203,N_4705,N_4662);
nor UO_204 (O_204,N_4788,N_4715);
nor UO_205 (O_205,N_4645,N_4527);
nor UO_206 (O_206,N_4650,N_4749);
nand UO_207 (O_207,N_4575,N_4842);
nor UO_208 (O_208,N_4594,N_4620);
and UO_209 (O_209,N_4632,N_4501);
and UO_210 (O_210,N_4722,N_4684);
nor UO_211 (O_211,N_4828,N_4834);
or UO_212 (O_212,N_4766,N_4730);
nand UO_213 (O_213,N_4532,N_4657);
nand UO_214 (O_214,N_4689,N_4907);
and UO_215 (O_215,N_4856,N_4837);
nand UO_216 (O_216,N_4747,N_4505);
or UO_217 (O_217,N_4658,N_4796);
and UO_218 (O_218,N_4673,N_4506);
nand UO_219 (O_219,N_4956,N_4895);
nand UO_220 (O_220,N_4843,N_4561);
nand UO_221 (O_221,N_4930,N_4637);
nor UO_222 (O_222,N_4579,N_4813);
or UO_223 (O_223,N_4649,N_4711);
nand UO_224 (O_224,N_4565,N_4516);
or UO_225 (O_225,N_4716,N_4933);
nor UO_226 (O_226,N_4954,N_4602);
nand UO_227 (O_227,N_4686,N_4654);
nand UO_228 (O_228,N_4643,N_4644);
and UO_229 (O_229,N_4839,N_4734);
and UO_230 (O_230,N_4811,N_4835);
and UO_231 (O_231,N_4625,N_4719);
or UO_232 (O_232,N_4968,N_4972);
nor UO_233 (O_233,N_4981,N_4612);
and UO_234 (O_234,N_4999,N_4598);
or UO_235 (O_235,N_4551,N_4803);
or UO_236 (O_236,N_4736,N_4890);
nor UO_237 (O_237,N_4802,N_4773);
nor UO_238 (O_238,N_4626,N_4667);
and UO_239 (O_239,N_4553,N_4878);
nand UO_240 (O_240,N_4577,N_4935);
and UO_241 (O_241,N_4732,N_4919);
or UO_242 (O_242,N_4857,N_4601);
or UO_243 (O_243,N_4511,N_4799);
and UO_244 (O_244,N_4638,N_4596);
nor UO_245 (O_245,N_4944,N_4998);
nand UO_246 (O_246,N_4958,N_4931);
and UO_247 (O_247,N_4815,N_4678);
or UO_248 (O_248,N_4606,N_4789);
or UO_249 (O_249,N_4949,N_4939);
and UO_250 (O_250,N_4522,N_4642);
nand UO_251 (O_251,N_4953,N_4708);
xor UO_252 (O_252,N_4769,N_4786);
nand UO_253 (O_253,N_4534,N_4829);
or UO_254 (O_254,N_4725,N_4742);
and UO_255 (O_255,N_4954,N_4678);
and UO_256 (O_256,N_4819,N_4998);
and UO_257 (O_257,N_4762,N_4952);
nand UO_258 (O_258,N_4929,N_4610);
or UO_259 (O_259,N_4538,N_4925);
or UO_260 (O_260,N_4542,N_4994);
nor UO_261 (O_261,N_4717,N_4815);
or UO_262 (O_262,N_4873,N_4746);
or UO_263 (O_263,N_4650,N_4776);
and UO_264 (O_264,N_4761,N_4691);
or UO_265 (O_265,N_4710,N_4776);
nor UO_266 (O_266,N_4556,N_4880);
nand UO_267 (O_267,N_4783,N_4713);
or UO_268 (O_268,N_4559,N_4714);
nor UO_269 (O_269,N_4648,N_4694);
nor UO_270 (O_270,N_4960,N_4837);
nand UO_271 (O_271,N_4691,N_4696);
and UO_272 (O_272,N_4604,N_4913);
and UO_273 (O_273,N_4977,N_4526);
nor UO_274 (O_274,N_4546,N_4558);
and UO_275 (O_275,N_4806,N_4951);
nor UO_276 (O_276,N_4910,N_4757);
nand UO_277 (O_277,N_4805,N_4716);
or UO_278 (O_278,N_4821,N_4529);
and UO_279 (O_279,N_4724,N_4877);
nor UO_280 (O_280,N_4959,N_4704);
and UO_281 (O_281,N_4802,N_4581);
or UO_282 (O_282,N_4914,N_4607);
or UO_283 (O_283,N_4997,N_4895);
nor UO_284 (O_284,N_4728,N_4975);
nor UO_285 (O_285,N_4569,N_4561);
or UO_286 (O_286,N_4860,N_4834);
nor UO_287 (O_287,N_4847,N_4986);
nor UO_288 (O_288,N_4981,N_4726);
nor UO_289 (O_289,N_4535,N_4992);
nor UO_290 (O_290,N_4569,N_4917);
and UO_291 (O_291,N_4884,N_4887);
and UO_292 (O_292,N_4609,N_4891);
or UO_293 (O_293,N_4507,N_4704);
nor UO_294 (O_294,N_4880,N_4564);
nand UO_295 (O_295,N_4540,N_4857);
or UO_296 (O_296,N_4952,N_4550);
and UO_297 (O_297,N_4552,N_4959);
or UO_298 (O_298,N_4931,N_4969);
nand UO_299 (O_299,N_4702,N_4648);
and UO_300 (O_300,N_4836,N_4918);
nor UO_301 (O_301,N_4784,N_4560);
nor UO_302 (O_302,N_4786,N_4761);
or UO_303 (O_303,N_4867,N_4981);
nand UO_304 (O_304,N_4589,N_4637);
and UO_305 (O_305,N_4584,N_4624);
or UO_306 (O_306,N_4776,N_4518);
and UO_307 (O_307,N_4514,N_4955);
and UO_308 (O_308,N_4943,N_4589);
or UO_309 (O_309,N_4620,N_4520);
or UO_310 (O_310,N_4967,N_4970);
nor UO_311 (O_311,N_4781,N_4638);
or UO_312 (O_312,N_4554,N_4550);
and UO_313 (O_313,N_4856,N_4886);
or UO_314 (O_314,N_4595,N_4796);
nor UO_315 (O_315,N_4942,N_4997);
nand UO_316 (O_316,N_4957,N_4512);
and UO_317 (O_317,N_4720,N_4887);
or UO_318 (O_318,N_4594,N_4512);
and UO_319 (O_319,N_4945,N_4509);
nand UO_320 (O_320,N_4917,N_4739);
or UO_321 (O_321,N_4875,N_4984);
nand UO_322 (O_322,N_4753,N_4660);
and UO_323 (O_323,N_4858,N_4709);
or UO_324 (O_324,N_4836,N_4594);
and UO_325 (O_325,N_4881,N_4772);
nand UO_326 (O_326,N_4776,N_4784);
xor UO_327 (O_327,N_4668,N_4725);
or UO_328 (O_328,N_4922,N_4928);
or UO_329 (O_329,N_4681,N_4568);
nor UO_330 (O_330,N_4923,N_4726);
nor UO_331 (O_331,N_4930,N_4733);
and UO_332 (O_332,N_4519,N_4997);
nor UO_333 (O_333,N_4856,N_4652);
and UO_334 (O_334,N_4837,N_4655);
or UO_335 (O_335,N_4980,N_4688);
nand UO_336 (O_336,N_4628,N_4758);
and UO_337 (O_337,N_4828,N_4902);
nor UO_338 (O_338,N_4566,N_4764);
nand UO_339 (O_339,N_4885,N_4585);
nor UO_340 (O_340,N_4577,N_4880);
nor UO_341 (O_341,N_4987,N_4758);
nor UO_342 (O_342,N_4865,N_4645);
nor UO_343 (O_343,N_4722,N_4575);
nand UO_344 (O_344,N_4669,N_4531);
nor UO_345 (O_345,N_4581,N_4991);
or UO_346 (O_346,N_4623,N_4956);
nor UO_347 (O_347,N_4709,N_4990);
or UO_348 (O_348,N_4675,N_4812);
nand UO_349 (O_349,N_4627,N_4802);
or UO_350 (O_350,N_4872,N_4846);
and UO_351 (O_351,N_4965,N_4903);
nand UO_352 (O_352,N_4783,N_4942);
nand UO_353 (O_353,N_4849,N_4969);
nor UO_354 (O_354,N_4562,N_4951);
and UO_355 (O_355,N_4843,N_4886);
nor UO_356 (O_356,N_4666,N_4696);
nor UO_357 (O_357,N_4509,N_4605);
or UO_358 (O_358,N_4841,N_4593);
or UO_359 (O_359,N_4512,N_4755);
or UO_360 (O_360,N_4835,N_4704);
or UO_361 (O_361,N_4787,N_4838);
nor UO_362 (O_362,N_4786,N_4767);
nor UO_363 (O_363,N_4971,N_4601);
nand UO_364 (O_364,N_4931,N_4771);
nand UO_365 (O_365,N_4716,N_4741);
and UO_366 (O_366,N_4648,N_4655);
and UO_367 (O_367,N_4729,N_4693);
or UO_368 (O_368,N_4557,N_4951);
and UO_369 (O_369,N_4642,N_4900);
nor UO_370 (O_370,N_4886,N_4747);
and UO_371 (O_371,N_4686,N_4919);
or UO_372 (O_372,N_4743,N_4570);
or UO_373 (O_373,N_4968,N_4762);
nand UO_374 (O_374,N_4770,N_4565);
and UO_375 (O_375,N_4993,N_4885);
or UO_376 (O_376,N_4664,N_4646);
nor UO_377 (O_377,N_4533,N_4601);
nand UO_378 (O_378,N_4695,N_4708);
nor UO_379 (O_379,N_4543,N_4977);
nand UO_380 (O_380,N_4532,N_4950);
nand UO_381 (O_381,N_4708,N_4535);
nor UO_382 (O_382,N_4731,N_4722);
nand UO_383 (O_383,N_4871,N_4968);
or UO_384 (O_384,N_4516,N_4761);
and UO_385 (O_385,N_4634,N_4773);
or UO_386 (O_386,N_4899,N_4963);
nor UO_387 (O_387,N_4937,N_4619);
and UO_388 (O_388,N_4569,N_4992);
and UO_389 (O_389,N_4708,N_4653);
nor UO_390 (O_390,N_4871,N_4928);
nor UO_391 (O_391,N_4587,N_4939);
and UO_392 (O_392,N_4516,N_4692);
or UO_393 (O_393,N_4949,N_4771);
and UO_394 (O_394,N_4983,N_4747);
nor UO_395 (O_395,N_4775,N_4519);
or UO_396 (O_396,N_4515,N_4857);
nand UO_397 (O_397,N_4824,N_4698);
nand UO_398 (O_398,N_4907,N_4628);
nand UO_399 (O_399,N_4848,N_4917);
or UO_400 (O_400,N_4622,N_4995);
nor UO_401 (O_401,N_4558,N_4835);
nor UO_402 (O_402,N_4870,N_4973);
nand UO_403 (O_403,N_4643,N_4816);
or UO_404 (O_404,N_4639,N_4978);
nor UO_405 (O_405,N_4762,N_4606);
nand UO_406 (O_406,N_4828,N_4969);
nand UO_407 (O_407,N_4648,N_4893);
nand UO_408 (O_408,N_4817,N_4835);
nor UO_409 (O_409,N_4883,N_4750);
and UO_410 (O_410,N_4862,N_4673);
or UO_411 (O_411,N_4696,N_4742);
nand UO_412 (O_412,N_4789,N_4807);
nor UO_413 (O_413,N_4996,N_4938);
nand UO_414 (O_414,N_4677,N_4766);
nor UO_415 (O_415,N_4919,N_4817);
nand UO_416 (O_416,N_4505,N_4873);
and UO_417 (O_417,N_4858,N_4550);
nor UO_418 (O_418,N_4566,N_4838);
nand UO_419 (O_419,N_4950,N_4556);
nand UO_420 (O_420,N_4612,N_4701);
xnor UO_421 (O_421,N_4604,N_4933);
and UO_422 (O_422,N_4947,N_4825);
or UO_423 (O_423,N_4604,N_4889);
and UO_424 (O_424,N_4657,N_4566);
or UO_425 (O_425,N_4642,N_4941);
or UO_426 (O_426,N_4838,N_4724);
and UO_427 (O_427,N_4880,N_4643);
and UO_428 (O_428,N_4674,N_4970);
or UO_429 (O_429,N_4796,N_4757);
or UO_430 (O_430,N_4868,N_4534);
or UO_431 (O_431,N_4811,N_4599);
and UO_432 (O_432,N_4836,N_4823);
nor UO_433 (O_433,N_4618,N_4926);
and UO_434 (O_434,N_4732,N_4908);
nor UO_435 (O_435,N_4802,N_4934);
and UO_436 (O_436,N_4820,N_4610);
nand UO_437 (O_437,N_4717,N_4664);
nand UO_438 (O_438,N_4712,N_4963);
nor UO_439 (O_439,N_4953,N_4578);
and UO_440 (O_440,N_4880,N_4686);
nand UO_441 (O_441,N_4798,N_4665);
nand UO_442 (O_442,N_4865,N_4732);
and UO_443 (O_443,N_4884,N_4717);
and UO_444 (O_444,N_4840,N_4520);
and UO_445 (O_445,N_4648,N_4801);
or UO_446 (O_446,N_4597,N_4821);
and UO_447 (O_447,N_4782,N_4891);
nor UO_448 (O_448,N_4904,N_4810);
or UO_449 (O_449,N_4512,N_4570);
nand UO_450 (O_450,N_4820,N_4785);
or UO_451 (O_451,N_4781,N_4696);
nand UO_452 (O_452,N_4730,N_4741);
or UO_453 (O_453,N_4804,N_4565);
nand UO_454 (O_454,N_4793,N_4737);
nand UO_455 (O_455,N_4873,N_4694);
or UO_456 (O_456,N_4879,N_4687);
nor UO_457 (O_457,N_4801,N_4813);
or UO_458 (O_458,N_4730,N_4715);
and UO_459 (O_459,N_4547,N_4863);
nand UO_460 (O_460,N_4792,N_4753);
or UO_461 (O_461,N_4506,N_4586);
xor UO_462 (O_462,N_4856,N_4748);
or UO_463 (O_463,N_4503,N_4770);
and UO_464 (O_464,N_4819,N_4713);
nor UO_465 (O_465,N_4699,N_4738);
and UO_466 (O_466,N_4542,N_4913);
nand UO_467 (O_467,N_4882,N_4909);
nor UO_468 (O_468,N_4594,N_4821);
nand UO_469 (O_469,N_4770,N_4866);
and UO_470 (O_470,N_4604,N_4908);
or UO_471 (O_471,N_4835,N_4954);
or UO_472 (O_472,N_4871,N_4750);
nand UO_473 (O_473,N_4576,N_4867);
and UO_474 (O_474,N_4832,N_4968);
nand UO_475 (O_475,N_4995,N_4859);
nand UO_476 (O_476,N_4883,N_4621);
nor UO_477 (O_477,N_4685,N_4540);
nand UO_478 (O_478,N_4574,N_4612);
nand UO_479 (O_479,N_4799,N_4820);
or UO_480 (O_480,N_4714,N_4763);
nor UO_481 (O_481,N_4537,N_4735);
nor UO_482 (O_482,N_4892,N_4776);
or UO_483 (O_483,N_4856,N_4924);
nor UO_484 (O_484,N_4828,N_4602);
nor UO_485 (O_485,N_4890,N_4613);
nand UO_486 (O_486,N_4859,N_4752);
nand UO_487 (O_487,N_4943,N_4937);
xor UO_488 (O_488,N_4681,N_4585);
or UO_489 (O_489,N_4939,N_4650);
nand UO_490 (O_490,N_4764,N_4556);
nor UO_491 (O_491,N_4911,N_4606);
and UO_492 (O_492,N_4972,N_4819);
or UO_493 (O_493,N_4607,N_4965);
nor UO_494 (O_494,N_4822,N_4816);
or UO_495 (O_495,N_4815,N_4754);
nand UO_496 (O_496,N_4770,N_4900);
and UO_497 (O_497,N_4976,N_4727);
nor UO_498 (O_498,N_4731,N_4581);
nor UO_499 (O_499,N_4532,N_4986);
nand UO_500 (O_500,N_4645,N_4711);
and UO_501 (O_501,N_4697,N_4647);
nor UO_502 (O_502,N_4670,N_4961);
nor UO_503 (O_503,N_4761,N_4716);
or UO_504 (O_504,N_4762,N_4613);
or UO_505 (O_505,N_4753,N_4856);
nor UO_506 (O_506,N_4818,N_4969);
or UO_507 (O_507,N_4667,N_4884);
and UO_508 (O_508,N_4747,N_4677);
nor UO_509 (O_509,N_4688,N_4869);
or UO_510 (O_510,N_4740,N_4534);
nand UO_511 (O_511,N_4745,N_4945);
nor UO_512 (O_512,N_4724,N_4682);
or UO_513 (O_513,N_4929,N_4676);
nand UO_514 (O_514,N_4555,N_4867);
and UO_515 (O_515,N_4951,N_4961);
and UO_516 (O_516,N_4657,N_4703);
or UO_517 (O_517,N_4890,N_4638);
nor UO_518 (O_518,N_4770,N_4600);
nand UO_519 (O_519,N_4981,N_4679);
nand UO_520 (O_520,N_4727,N_4536);
nand UO_521 (O_521,N_4792,N_4741);
and UO_522 (O_522,N_4783,N_4554);
or UO_523 (O_523,N_4515,N_4598);
or UO_524 (O_524,N_4538,N_4784);
and UO_525 (O_525,N_4869,N_4707);
nand UO_526 (O_526,N_4866,N_4826);
or UO_527 (O_527,N_4901,N_4860);
nand UO_528 (O_528,N_4794,N_4550);
nand UO_529 (O_529,N_4593,N_4670);
nor UO_530 (O_530,N_4723,N_4982);
nand UO_531 (O_531,N_4810,N_4875);
and UO_532 (O_532,N_4912,N_4648);
and UO_533 (O_533,N_4826,N_4569);
nor UO_534 (O_534,N_4534,N_4903);
or UO_535 (O_535,N_4945,N_4763);
or UO_536 (O_536,N_4563,N_4608);
nor UO_537 (O_537,N_4671,N_4554);
and UO_538 (O_538,N_4510,N_4586);
nor UO_539 (O_539,N_4722,N_4868);
and UO_540 (O_540,N_4893,N_4653);
nor UO_541 (O_541,N_4510,N_4582);
nand UO_542 (O_542,N_4542,N_4594);
and UO_543 (O_543,N_4559,N_4865);
and UO_544 (O_544,N_4661,N_4566);
nor UO_545 (O_545,N_4815,N_4876);
nor UO_546 (O_546,N_4664,N_4883);
nand UO_547 (O_547,N_4766,N_4579);
and UO_548 (O_548,N_4790,N_4956);
nand UO_549 (O_549,N_4955,N_4628);
or UO_550 (O_550,N_4697,N_4644);
nand UO_551 (O_551,N_4770,N_4859);
or UO_552 (O_552,N_4550,N_4664);
nor UO_553 (O_553,N_4881,N_4984);
and UO_554 (O_554,N_4999,N_4550);
and UO_555 (O_555,N_4636,N_4698);
nor UO_556 (O_556,N_4845,N_4626);
or UO_557 (O_557,N_4794,N_4636);
nand UO_558 (O_558,N_4885,N_4633);
or UO_559 (O_559,N_4821,N_4796);
xor UO_560 (O_560,N_4901,N_4581);
or UO_561 (O_561,N_4536,N_4763);
or UO_562 (O_562,N_4764,N_4585);
nand UO_563 (O_563,N_4623,N_4760);
nand UO_564 (O_564,N_4819,N_4709);
and UO_565 (O_565,N_4780,N_4808);
nor UO_566 (O_566,N_4839,N_4544);
nand UO_567 (O_567,N_4886,N_4842);
nand UO_568 (O_568,N_4929,N_4591);
nor UO_569 (O_569,N_4786,N_4832);
and UO_570 (O_570,N_4601,N_4671);
nand UO_571 (O_571,N_4806,N_4860);
nor UO_572 (O_572,N_4987,N_4995);
nor UO_573 (O_573,N_4601,N_4885);
or UO_574 (O_574,N_4771,N_4822);
or UO_575 (O_575,N_4969,N_4700);
nand UO_576 (O_576,N_4517,N_4805);
or UO_577 (O_577,N_4759,N_4986);
or UO_578 (O_578,N_4775,N_4611);
and UO_579 (O_579,N_4847,N_4787);
nor UO_580 (O_580,N_4997,N_4709);
nor UO_581 (O_581,N_4542,N_4993);
nor UO_582 (O_582,N_4677,N_4988);
nor UO_583 (O_583,N_4968,N_4964);
and UO_584 (O_584,N_4873,N_4595);
nor UO_585 (O_585,N_4901,N_4951);
or UO_586 (O_586,N_4501,N_4956);
nor UO_587 (O_587,N_4634,N_4934);
and UO_588 (O_588,N_4779,N_4622);
or UO_589 (O_589,N_4837,N_4710);
nand UO_590 (O_590,N_4782,N_4671);
nor UO_591 (O_591,N_4504,N_4515);
and UO_592 (O_592,N_4589,N_4571);
or UO_593 (O_593,N_4778,N_4892);
nor UO_594 (O_594,N_4652,N_4580);
nor UO_595 (O_595,N_4669,N_4708);
or UO_596 (O_596,N_4610,N_4592);
nand UO_597 (O_597,N_4511,N_4930);
nand UO_598 (O_598,N_4503,N_4938);
and UO_599 (O_599,N_4725,N_4502);
or UO_600 (O_600,N_4727,N_4722);
nor UO_601 (O_601,N_4966,N_4665);
nand UO_602 (O_602,N_4884,N_4640);
nand UO_603 (O_603,N_4546,N_4994);
and UO_604 (O_604,N_4563,N_4889);
or UO_605 (O_605,N_4800,N_4822);
nor UO_606 (O_606,N_4515,N_4620);
nand UO_607 (O_607,N_4889,N_4630);
nand UO_608 (O_608,N_4954,N_4748);
nor UO_609 (O_609,N_4503,N_4917);
or UO_610 (O_610,N_4814,N_4881);
xor UO_611 (O_611,N_4625,N_4643);
or UO_612 (O_612,N_4720,N_4774);
or UO_613 (O_613,N_4772,N_4802);
or UO_614 (O_614,N_4865,N_4990);
and UO_615 (O_615,N_4578,N_4545);
or UO_616 (O_616,N_4618,N_4542);
and UO_617 (O_617,N_4798,N_4852);
or UO_618 (O_618,N_4643,N_4907);
nor UO_619 (O_619,N_4940,N_4969);
or UO_620 (O_620,N_4996,N_4920);
and UO_621 (O_621,N_4743,N_4613);
nor UO_622 (O_622,N_4733,N_4534);
and UO_623 (O_623,N_4753,N_4935);
or UO_624 (O_624,N_4558,N_4508);
nor UO_625 (O_625,N_4652,N_4785);
and UO_626 (O_626,N_4625,N_4772);
nand UO_627 (O_627,N_4793,N_4951);
nand UO_628 (O_628,N_4668,N_4859);
nand UO_629 (O_629,N_4554,N_4927);
nor UO_630 (O_630,N_4688,N_4661);
and UO_631 (O_631,N_4844,N_4514);
nor UO_632 (O_632,N_4899,N_4592);
and UO_633 (O_633,N_4752,N_4842);
nand UO_634 (O_634,N_4995,N_4816);
or UO_635 (O_635,N_4749,N_4776);
nand UO_636 (O_636,N_4893,N_4505);
nand UO_637 (O_637,N_4771,N_4667);
nor UO_638 (O_638,N_4592,N_4593);
and UO_639 (O_639,N_4683,N_4662);
xnor UO_640 (O_640,N_4543,N_4744);
and UO_641 (O_641,N_4884,N_4537);
nand UO_642 (O_642,N_4725,N_4854);
nand UO_643 (O_643,N_4864,N_4584);
nand UO_644 (O_644,N_4518,N_4999);
nand UO_645 (O_645,N_4864,N_4979);
or UO_646 (O_646,N_4945,N_4969);
nor UO_647 (O_647,N_4675,N_4956);
nor UO_648 (O_648,N_4543,N_4819);
and UO_649 (O_649,N_4880,N_4841);
nor UO_650 (O_650,N_4821,N_4945);
nor UO_651 (O_651,N_4675,N_4559);
or UO_652 (O_652,N_4865,N_4840);
nor UO_653 (O_653,N_4821,N_4921);
and UO_654 (O_654,N_4855,N_4660);
nand UO_655 (O_655,N_4727,N_4649);
and UO_656 (O_656,N_4956,N_4850);
nor UO_657 (O_657,N_4969,N_4894);
nand UO_658 (O_658,N_4976,N_4642);
or UO_659 (O_659,N_4839,N_4551);
or UO_660 (O_660,N_4797,N_4617);
and UO_661 (O_661,N_4952,N_4616);
and UO_662 (O_662,N_4907,N_4516);
and UO_663 (O_663,N_4931,N_4697);
or UO_664 (O_664,N_4723,N_4621);
or UO_665 (O_665,N_4783,N_4539);
nand UO_666 (O_666,N_4746,N_4672);
or UO_667 (O_667,N_4780,N_4903);
and UO_668 (O_668,N_4848,N_4993);
nor UO_669 (O_669,N_4743,N_4631);
nor UO_670 (O_670,N_4806,N_4821);
nand UO_671 (O_671,N_4513,N_4941);
and UO_672 (O_672,N_4900,N_4664);
nand UO_673 (O_673,N_4710,N_4852);
nand UO_674 (O_674,N_4509,N_4684);
nor UO_675 (O_675,N_4596,N_4625);
nor UO_676 (O_676,N_4746,N_4822);
and UO_677 (O_677,N_4500,N_4949);
or UO_678 (O_678,N_4912,N_4533);
nor UO_679 (O_679,N_4931,N_4888);
nand UO_680 (O_680,N_4907,N_4992);
nor UO_681 (O_681,N_4945,N_4867);
or UO_682 (O_682,N_4878,N_4858);
and UO_683 (O_683,N_4535,N_4893);
and UO_684 (O_684,N_4807,N_4544);
nand UO_685 (O_685,N_4570,N_4694);
or UO_686 (O_686,N_4680,N_4588);
nand UO_687 (O_687,N_4517,N_4972);
nand UO_688 (O_688,N_4664,N_4527);
or UO_689 (O_689,N_4641,N_4816);
and UO_690 (O_690,N_4735,N_4997);
nor UO_691 (O_691,N_4843,N_4700);
nand UO_692 (O_692,N_4917,N_4579);
nand UO_693 (O_693,N_4595,N_4533);
nor UO_694 (O_694,N_4909,N_4672);
and UO_695 (O_695,N_4915,N_4838);
nor UO_696 (O_696,N_4611,N_4560);
and UO_697 (O_697,N_4633,N_4960);
or UO_698 (O_698,N_4976,N_4842);
and UO_699 (O_699,N_4896,N_4748);
or UO_700 (O_700,N_4919,N_4846);
nor UO_701 (O_701,N_4500,N_4548);
or UO_702 (O_702,N_4782,N_4947);
nand UO_703 (O_703,N_4730,N_4989);
nand UO_704 (O_704,N_4940,N_4875);
or UO_705 (O_705,N_4682,N_4679);
or UO_706 (O_706,N_4659,N_4538);
and UO_707 (O_707,N_4946,N_4664);
nand UO_708 (O_708,N_4811,N_4577);
or UO_709 (O_709,N_4813,N_4715);
or UO_710 (O_710,N_4939,N_4796);
and UO_711 (O_711,N_4908,N_4643);
xor UO_712 (O_712,N_4871,N_4733);
nand UO_713 (O_713,N_4820,N_4842);
and UO_714 (O_714,N_4631,N_4637);
and UO_715 (O_715,N_4754,N_4524);
and UO_716 (O_716,N_4539,N_4860);
and UO_717 (O_717,N_4838,N_4803);
nand UO_718 (O_718,N_4649,N_4824);
nor UO_719 (O_719,N_4874,N_4812);
nand UO_720 (O_720,N_4809,N_4540);
or UO_721 (O_721,N_4694,N_4724);
or UO_722 (O_722,N_4921,N_4614);
or UO_723 (O_723,N_4665,N_4614);
and UO_724 (O_724,N_4955,N_4954);
nor UO_725 (O_725,N_4980,N_4804);
nor UO_726 (O_726,N_4750,N_4574);
or UO_727 (O_727,N_4885,N_4921);
nand UO_728 (O_728,N_4903,N_4573);
nand UO_729 (O_729,N_4887,N_4885);
nand UO_730 (O_730,N_4619,N_4947);
or UO_731 (O_731,N_4838,N_4624);
nand UO_732 (O_732,N_4935,N_4556);
or UO_733 (O_733,N_4649,N_4633);
or UO_734 (O_734,N_4505,N_4923);
or UO_735 (O_735,N_4939,N_4831);
and UO_736 (O_736,N_4901,N_4942);
or UO_737 (O_737,N_4786,N_4803);
and UO_738 (O_738,N_4919,N_4663);
nor UO_739 (O_739,N_4747,N_4518);
or UO_740 (O_740,N_4586,N_4527);
nor UO_741 (O_741,N_4961,N_4962);
or UO_742 (O_742,N_4797,N_4500);
nor UO_743 (O_743,N_4623,N_4639);
or UO_744 (O_744,N_4524,N_4788);
nor UO_745 (O_745,N_4577,N_4714);
and UO_746 (O_746,N_4682,N_4614);
nor UO_747 (O_747,N_4590,N_4751);
nor UO_748 (O_748,N_4677,N_4711);
or UO_749 (O_749,N_4869,N_4951);
nand UO_750 (O_750,N_4536,N_4575);
and UO_751 (O_751,N_4805,N_4829);
and UO_752 (O_752,N_4842,N_4534);
nand UO_753 (O_753,N_4650,N_4826);
and UO_754 (O_754,N_4570,N_4954);
or UO_755 (O_755,N_4694,N_4998);
and UO_756 (O_756,N_4987,N_4555);
nor UO_757 (O_757,N_4651,N_4701);
and UO_758 (O_758,N_4744,N_4653);
and UO_759 (O_759,N_4895,N_4524);
or UO_760 (O_760,N_4800,N_4750);
or UO_761 (O_761,N_4985,N_4813);
nand UO_762 (O_762,N_4879,N_4699);
nor UO_763 (O_763,N_4939,N_4564);
or UO_764 (O_764,N_4963,N_4538);
xnor UO_765 (O_765,N_4961,N_4821);
xnor UO_766 (O_766,N_4571,N_4649);
nor UO_767 (O_767,N_4771,N_4938);
or UO_768 (O_768,N_4794,N_4736);
nor UO_769 (O_769,N_4584,N_4988);
nand UO_770 (O_770,N_4871,N_4858);
and UO_771 (O_771,N_4660,N_4830);
and UO_772 (O_772,N_4603,N_4846);
or UO_773 (O_773,N_4669,N_4988);
and UO_774 (O_774,N_4794,N_4782);
nand UO_775 (O_775,N_4669,N_4878);
nand UO_776 (O_776,N_4591,N_4754);
nand UO_777 (O_777,N_4528,N_4644);
or UO_778 (O_778,N_4720,N_4697);
or UO_779 (O_779,N_4907,N_4911);
and UO_780 (O_780,N_4526,N_4863);
or UO_781 (O_781,N_4791,N_4899);
nor UO_782 (O_782,N_4725,N_4734);
nor UO_783 (O_783,N_4731,N_4857);
or UO_784 (O_784,N_4719,N_4933);
nand UO_785 (O_785,N_4927,N_4695);
and UO_786 (O_786,N_4758,N_4681);
or UO_787 (O_787,N_4644,N_4598);
or UO_788 (O_788,N_4614,N_4958);
or UO_789 (O_789,N_4594,N_4841);
nor UO_790 (O_790,N_4607,N_4830);
and UO_791 (O_791,N_4969,N_4733);
nand UO_792 (O_792,N_4778,N_4675);
or UO_793 (O_793,N_4600,N_4904);
nand UO_794 (O_794,N_4558,N_4534);
nand UO_795 (O_795,N_4608,N_4547);
and UO_796 (O_796,N_4831,N_4997);
nor UO_797 (O_797,N_4829,N_4678);
or UO_798 (O_798,N_4729,N_4735);
or UO_799 (O_799,N_4635,N_4615);
nor UO_800 (O_800,N_4835,N_4922);
nor UO_801 (O_801,N_4576,N_4566);
nor UO_802 (O_802,N_4690,N_4641);
or UO_803 (O_803,N_4807,N_4553);
and UO_804 (O_804,N_4620,N_4737);
and UO_805 (O_805,N_4748,N_4701);
or UO_806 (O_806,N_4630,N_4897);
or UO_807 (O_807,N_4657,N_4928);
nand UO_808 (O_808,N_4683,N_4674);
nor UO_809 (O_809,N_4538,N_4610);
or UO_810 (O_810,N_4724,N_4847);
and UO_811 (O_811,N_4957,N_4600);
or UO_812 (O_812,N_4558,N_4660);
nor UO_813 (O_813,N_4753,N_4766);
nor UO_814 (O_814,N_4979,N_4723);
nand UO_815 (O_815,N_4618,N_4982);
nand UO_816 (O_816,N_4532,N_4881);
nand UO_817 (O_817,N_4804,N_4874);
nor UO_818 (O_818,N_4508,N_4797);
nor UO_819 (O_819,N_4561,N_4824);
nand UO_820 (O_820,N_4805,N_4705);
nand UO_821 (O_821,N_4812,N_4906);
nand UO_822 (O_822,N_4912,N_4501);
nand UO_823 (O_823,N_4917,N_4796);
and UO_824 (O_824,N_4539,N_4959);
or UO_825 (O_825,N_4557,N_4515);
nor UO_826 (O_826,N_4617,N_4843);
nand UO_827 (O_827,N_4920,N_4787);
nor UO_828 (O_828,N_4672,N_4563);
and UO_829 (O_829,N_4765,N_4939);
nand UO_830 (O_830,N_4980,N_4825);
or UO_831 (O_831,N_4692,N_4989);
nand UO_832 (O_832,N_4653,N_4584);
nor UO_833 (O_833,N_4975,N_4936);
nand UO_834 (O_834,N_4982,N_4945);
nor UO_835 (O_835,N_4889,N_4928);
xnor UO_836 (O_836,N_4807,N_4571);
or UO_837 (O_837,N_4921,N_4564);
nor UO_838 (O_838,N_4855,N_4833);
nor UO_839 (O_839,N_4752,N_4541);
nand UO_840 (O_840,N_4954,N_4561);
and UO_841 (O_841,N_4853,N_4659);
nor UO_842 (O_842,N_4626,N_4708);
nand UO_843 (O_843,N_4960,N_4702);
or UO_844 (O_844,N_4543,N_4565);
or UO_845 (O_845,N_4911,N_4774);
nor UO_846 (O_846,N_4542,N_4755);
or UO_847 (O_847,N_4657,N_4847);
nor UO_848 (O_848,N_4607,N_4672);
nand UO_849 (O_849,N_4741,N_4842);
xor UO_850 (O_850,N_4638,N_4926);
and UO_851 (O_851,N_4782,N_4814);
nand UO_852 (O_852,N_4727,N_4706);
and UO_853 (O_853,N_4745,N_4723);
or UO_854 (O_854,N_4501,N_4899);
or UO_855 (O_855,N_4786,N_4737);
or UO_856 (O_856,N_4742,N_4749);
nor UO_857 (O_857,N_4597,N_4706);
nand UO_858 (O_858,N_4828,N_4847);
nand UO_859 (O_859,N_4999,N_4589);
nor UO_860 (O_860,N_4564,N_4929);
nand UO_861 (O_861,N_4781,N_4742);
and UO_862 (O_862,N_4511,N_4593);
or UO_863 (O_863,N_4674,N_4807);
nor UO_864 (O_864,N_4762,N_4600);
and UO_865 (O_865,N_4657,N_4874);
nor UO_866 (O_866,N_4729,N_4570);
and UO_867 (O_867,N_4592,N_4671);
and UO_868 (O_868,N_4658,N_4694);
and UO_869 (O_869,N_4667,N_4598);
or UO_870 (O_870,N_4701,N_4875);
and UO_871 (O_871,N_4759,N_4900);
or UO_872 (O_872,N_4964,N_4708);
and UO_873 (O_873,N_4985,N_4525);
nand UO_874 (O_874,N_4906,N_4951);
nand UO_875 (O_875,N_4950,N_4550);
nand UO_876 (O_876,N_4647,N_4823);
and UO_877 (O_877,N_4704,N_4568);
nor UO_878 (O_878,N_4884,N_4830);
nand UO_879 (O_879,N_4799,N_4653);
nand UO_880 (O_880,N_4518,N_4579);
nand UO_881 (O_881,N_4763,N_4659);
or UO_882 (O_882,N_4835,N_4532);
and UO_883 (O_883,N_4501,N_4542);
nand UO_884 (O_884,N_4938,N_4691);
nand UO_885 (O_885,N_4945,N_4528);
nor UO_886 (O_886,N_4655,N_4783);
nand UO_887 (O_887,N_4752,N_4872);
or UO_888 (O_888,N_4840,N_4597);
nor UO_889 (O_889,N_4723,N_4532);
nand UO_890 (O_890,N_4706,N_4866);
and UO_891 (O_891,N_4757,N_4742);
or UO_892 (O_892,N_4916,N_4948);
or UO_893 (O_893,N_4840,N_4957);
or UO_894 (O_894,N_4701,N_4510);
or UO_895 (O_895,N_4547,N_4969);
nor UO_896 (O_896,N_4809,N_4838);
and UO_897 (O_897,N_4671,N_4626);
nand UO_898 (O_898,N_4562,N_4791);
nor UO_899 (O_899,N_4878,N_4747);
nor UO_900 (O_900,N_4993,N_4878);
nor UO_901 (O_901,N_4977,N_4932);
or UO_902 (O_902,N_4922,N_4721);
nand UO_903 (O_903,N_4635,N_4862);
xor UO_904 (O_904,N_4634,N_4788);
nand UO_905 (O_905,N_4691,N_4931);
or UO_906 (O_906,N_4792,N_4900);
nor UO_907 (O_907,N_4773,N_4932);
nor UO_908 (O_908,N_4958,N_4774);
and UO_909 (O_909,N_4509,N_4859);
nand UO_910 (O_910,N_4879,N_4753);
nand UO_911 (O_911,N_4858,N_4886);
nor UO_912 (O_912,N_4546,N_4603);
or UO_913 (O_913,N_4501,N_4898);
or UO_914 (O_914,N_4586,N_4533);
or UO_915 (O_915,N_4512,N_4989);
and UO_916 (O_916,N_4646,N_4609);
nor UO_917 (O_917,N_4577,N_4877);
and UO_918 (O_918,N_4697,N_4914);
and UO_919 (O_919,N_4676,N_4733);
or UO_920 (O_920,N_4549,N_4984);
or UO_921 (O_921,N_4614,N_4660);
and UO_922 (O_922,N_4631,N_4998);
and UO_923 (O_923,N_4777,N_4812);
nor UO_924 (O_924,N_4628,N_4887);
nor UO_925 (O_925,N_4944,N_4636);
and UO_926 (O_926,N_4790,N_4804);
nor UO_927 (O_927,N_4968,N_4685);
or UO_928 (O_928,N_4935,N_4679);
nor UO_929 (O_929,N_4636,N_4946);
nor UO_930 (O_930,N_4513,N_4934);
or UO_931 (O_931,N_4905,N_4507);
nand UO_932 (O_932,N_4986,N_4648);
nor UO_933 (O_933,N_4897,N_4627);
or UO_934 (O_934,N_4660,N_4835);
or UO_935 (O_935,N_4877,N_4682);
and UO_936 (O_936,N_4558,N_4841);
nor UO_937 (O_937,N_4655,N_4626);
nand UO_938 (O_938,N_4691,N_4690);
and UO_939 (O_939,N_4909,N_4872);
and UO_940 (O_940,N_4919,N_4810);
or UO_941 (O_941,N_4897,N_4612);
and UO_942 (O_942,N_4676,N_4610);
or UO_943 (O_943,N_4920,N_4925);
and UO_944 (O_944,N_4780,N_4863);
nor UO_945 (O_945,N_4688,N_4520);
nor UO_946 (O_946,N_4920,N_4731);
nand UO_947 (O_947,N_4842,N_4986);
nor UO_948 (O_948,N_4601,N_4611);
nand UO_949 (O_949,N_4936,N_4797);
or UO_950 (O_950,N_4807,N_4896);
nor UO_951 (O_951,N_4579,N_4967);
nor UO_952 (O_952,N_4782,N_4756);
or UO_953 (O_953,N_4900,N_4943);
nor UO_954 (O_954,N_4945,N_4782);
nor UO_955 (O_955,N_4824,N_4715);
nand UO_956 (O_956,N_4620,N_4847);
nor UO_957 (O_957,N_4918,N_4637);
nor UO_958 (O_958,N_4807,N_4893);
nand UO_959 (O_959,N_4624,N_4569);
nor UO_960 (O_960,N_4540,N_4614);
nand UO_961 (O_961,N_4806,N_4935);
nor UO_962 (O_962,N_4525,N_4863);
or UO_963 (O_963,N_4634,N_4768);
or UO_964 (O_964,N_4956,N_4715);
nor UO_965 (O_965,N_4713,N_4895);
nand UO_966 (O_966,N_4683,N_4671);
nand UO_967 (O_967,N_4562,N_4826);
nor UO_968 (O_968,N_4573,N_4751);
or UO_969 (O_969,N_4573,N_4539);
or UO_970 (O_970,N_4693,N_4570);
or UO_971 (O_971,N_4900,N_4797);
nor UO_972 (O_972,N_4935,N_4672);
or UO_973 (O_973,N_4783,N_4600);
nor UO_974 (O_974,N_4623,N_4851);
nand UO_975 (O_975,N_4953,N_4646);
and UO_976 (O_976,N_4907,N_4983);
nand UO_977 (O_977,N_4853,N_4937);
nand UO_978 (O_978,N_4623,N_4820);
nor UO_979 (O_979,N_4885,N_4527);
nand UO_980 (O_980,N_4674,N_4981);
nand UO_981 (O_981,N_4928,N_4958);
nand UO_982 (O_982,N_4665,N_4716);
xor UO_983 (O_983,N_4606,N_4853);
and UO_984 (O_984,N_4580,N_4931);
or UO_985 (O_985,N_4810,N_4627);
and UO_986 (O_986,N_4653,N_4936);
or UO_987 (O_987,N_4939,N_4719);
nor UO_988 (O_988,N_4891,N_4904);
nand UO_989 (O_989,N_4834,N_4916);
nor UO_990 (O_990,N_4815,N_4660);
and UO_991 (O_991,N_4913,N_4941);
nand UO_992 (O_992,N_4572,N_4843);
nand UO_993 (O_993,N_4568,N_4586);
and UO_994 (O_994,N_4902,N_4609);
or UO_995 (O_995,N_4761,N_4679);
nor UO_996 (O_996,N_4683,N_4987);
nor UO_997 (O_997,N_4998,N_4502);
or UO_998 (O_998,N_4935,N_4846);
nand UO_999 (O_999,N_4705,N_4550);
endmodule