module basic_750_5000_1000_5_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_3,In_322);
and U1 (N_1,In_375,In_669);
and U2 (N_2,In_419,In_355);
or U3 (N_3,In_657,In_523);
and U4 (N_4,In_721,In_134);
nand U5 (N_5,In_553,In_439);
nor U6 (N_6,In_8,In_241);
and U7 (N_7,In_118,In_86);
or U8 (N_8,In_547,In_283);
nor U9 (N_9,In_369,In_569);
and U10 (N_10,In_452,In_313);
nor U11 (N_11,In_487,In_195);
or U12 (N_12,In_179,In_645);
xnor U13 (N_13,In_738,In_160);
and U14 (N_14,In_142,In_665);
nand U15 (N_15,In_646,In_559);
nor U16 (N_16,In_692,In_295);
nand U17 (N_17,In_704,In_232);
and U18 (N_18,In_649,In_708);
and U19 (N_19,In_183,In_586);
nor U20 (N_20,In_576,In_144);
or U21 (N_21,In_475,In_397);
xnor U22 (N_22,In_82,In_521);
xor U23 (N_23,In_428,In_100);
nor U24 (N_24,In_388,In_543);
nand U25 (N_25,In_61,In_145);
and U26 (N_26,In_595,In_59);
and U27 (N_27,In_701,In_433);
and U28 (N_28,In_39,In_719);
and U29 (N_29,In_174,In_19);
nor U30 (N_30,In_450,In_529);
and U31 (N_31,In_262,In_583);
and U32 (N_32,In_16,In_231);
nand U33 (N_33,In_371,In_703);
or U34 (N_34,In_45,In_598);
and U35 (N_35,In_527,In_123);
and U36 (N_36,In_97,In_289);
or U37 (N_37,In_87,In_648);
nor U38 (N_38,In_479,In_349);
xnor U39 (N_39,In_666,In_55);
nand U40 (N_40,In_619,In_182);
nor U41 (N_41,In_417,In_334);
nand U42 (N_42,In_474,In_101);
nor U43 (N_43,In_415,In_281);
nand U44 (N_44,In_406,In_278);
nor U45 (N_45,In_320,In_66);
or U46 (N_46,In_718,In_266);
and U47 (N_47,In_98,In_374);
or U48 (N_48,In_85,In_264);
nor U49 (N_49,In_36,In_272);
and U50 (N_50,In_137,In_331);
nand U51 (N_51,In_270,In_133);
nor U52 (N_52,In_386,In_378);
and U53 (N_53,In_490,In_291);
xnor U54 (N_54,In_336,In_443);
xnor U55 (N_55,In_421,In_494);
or U56 (N_56,In_637,In_298);
nor U57 (N_57,In_573,In_725);
or U58 (N_58,In_372,In_502);
xnor U59 (N_59,In_720,In_238);
nand U60 (N_60,In_459,In_636);
xor U61 (N_61,In_260,In_267);
and U62 (N_62,In_207,In_467);
and U63 (N_63,In_317,In_726);
or U64 (N_64,In_41,In_357);
nand U65 (N_65,In_37,In_444);
or U66 (N_66,In_611,In_481);
and U67 (N_67,In_668,In_729);
or U68 (N_68,In_642,In_618);
xnor U69 (N_69,In_578,In_199);
and U70 (N_70,In_736,In_18);
or U71 (N_71,In_147,In_628);
or U72 (N_72,In_461,In_276);
xnor U73 (N_73,In_456,In_634);
nand U74 (N_74,In_186,In_548);
and U75 (N_75,In_505,In_293);
xnor U76 (N_76,In_518,In_339);
nand U77 (N_77,In_333,In_414);
or U78 (N_78,In_128,In_542);
nand U79 (N_79,In_215,In_663);
nor U80 (N_80,In_237,In_165);
nor U81 (N_81,In_508,In_211);
xnor U82 (N_82,In_497,In_525);
or U83 (N_83,In_710,In_344);
nand U84 (N_84,In_492,In_437);
nand U85 (N_85,In_728,In_79);
xor U86 (N_86,In_201,In_617);
and U87 (N_87,In_105,In_124);
or U88 (N_88,In_149,In_687);
and U89 (N_89,In_288,In_341);
nor U90 (N_90,In_612,In_498);
nand U91 (N_91,In_310,In_602);
nor U92 (N_92,In_706,In_482);
nand U93 (N_93,In_562,In_458);
and U94 (N_94,In_307,In_185);
nor U95 (N_95,In_608,In_256);
and U96 (N_96,In_65,In_28);
and U97 (N_97,In_680,In_566);
nand U98 (N_98,In_248,In_399);
xnor U99 (N_99,In_172,In_99);
nor U100 (N_100,In_507,In_208);
and U101 (N_101,In_323,In_156);
and U102 (N_102,In_640,In_202);
nor U103 (N_103,In_17,In_486);
xnor U104 (N_104,In_345,In_153);
nor U105 (N_105,In_33,In_359);
nand U106 (N_106,In_579,In_113);
or U107 (N_107,In_632,In_620);
or U108 (N_108,In_730,In_330);
or U109 (N_109,In_629,In_429);
nor U110 (N_110,In_252,In_589);
or U111 (N_111,In_12,In_213);
nand U112 (N_112,In_679,In_613);
or U113 (N_113,In_173,In_681);
xnor U114 (N_114,In_551,In_549);
nand U115 (N_115,In_300,In_277);
xnor U116 (N_116,In_392,In_658);
nand U117 (N_117,In_122,In_70);
and U118 (N_118,In_240,In_84);
nor U119 (N_119,In_223,In_520);
or U120 (N_120,In_102,In_540);
or U121 (N_121,In_396,In_319);
and U122 (N_122,In_23,In_29);
or U123 (N_123,In_387,In_327);
or U124 (N_124,In_664,In_591);
and U125 (N_125,In_109,In_190);
and U126 (N_126,In_683,In_220);
or U127 (N_127,In_711,In_138);
or U128 (N_128,In_600,In_279);
nor U129 (N_129,In_219,In_626);
nand U130 (N_130,In_214,In_77);
nor U131 (N_131,In_38,In_390);
nor U132 (N_132,In_453,In_111);
nand U133 (N_133,In_188,In_503);
and U134 (N_134,In_709,In_115);
and U135 (N_135,In_381,In_321);
nor U136 (N_136,In_175,In_13);
nor U137 (N_137,In_483,In_303);
xor U138 (N_138,In_6,In_373);
nor U139 (N_139,In_739,In_366);
nor U140 (N_140,In_221,In_218);
and U141 (N_141,In_247,In_21);
or U142 (N_142,In_255,In_574);
and U143 (N_143,In_564,In_233);
and U144 (N_144,In_440,In_741);
nor U145 (N_145,In_103,In_325);
and U146 (N_146,In_744,In_141);
nand U147 (N_147,In_148,In_367);
nand U148 (N_148,In_460,In_676);
or U149 (N_149,In_376,In_187);
nand U150 (N_150,In_592,In_210);
nor U151 (N_151,In_60,In_723);
or U152 (N_152,In_157,In_621);
and U153 (N_153,In_674,In_88);
nor U154 (N_154,In_643,In_423);
nand U155 (N_155,In_614,In_362);
or U156 (N_156,In_418,In_596);
xnor U157 (N_157,In_538,In_478);
or U158 (N_158,In_318,In_58);
nor U159 (N_159,In_32,In_107);
nor U160 (N_160,In_116,In_383);
and U161 (N_161,In_567,In_447);
and U162 (N_162,In_470,In_168);
and U163 (N_163,In_68,In_501);
and U164 (N_164,In_560,In_351);
and U165 (N_165,In_308,In_693);
or U166 (N_166,In_571,In_197);
or U167 (N_167,In_382,In_302);
nor U168 (N_168,In_469,In_724);
and U169 (N_169,In_599,In_44);
or U170 (N_170,In_40,In_426);
nor U171 (N_171,In_352,In_697);
or U172 (N_172,In_517,In_408);
or U173 (N_173,In_412,In_347);
xor U174 (N_174,In_696,In_164);
or U175 (N_175,In_265,In_607);
nand U176 (N_176,In_268,In_212);
and U177 (N_177,In_454,In_413);
and U178 (N_178,In_76,In_631);
or U179 (N_179,In_274,In_269);
or U180 (N_180,In_416,In_531);
and U181 (N_181,In_594,In_656);
and U182 (N_182,In_226,In_53);
and U183 (N_183,In_635,In_14);
nand U184 (N_184,In_71,In_504);
xnor U185 (N_185,In_633,In_332);
or U186 (N_186,In_609,In_555);
nand U187 (N_187,In_306,In_316);
xnor U188 (N_188,In_151,In_89);
and U189 (N_189,In_203,In_11);
xnor U190 (N_190,In_575,In_191);
and U191 (N_191,In_511,In_250);
and U192 (N_192,In_280,In_652);
nand U193 (N_193,In_228,In_743);
or U194 (N_194,In_615,In_209);
nor U195 (N_195,In_493,In_732);
nor U196 (N_196,In_678,In_159);
nor U197 (N_197,In_401,In_353);
nor U198 (N_198,In_242,In_370);
and U199 (N_199,In_749,In_604);
or U200 (N_200,In_556,In_427);
nand U201 (N_201,In_731,In_328);
or U202 (N_202,In_557,In_499);
and U203 (N_203,In_129,In_305);
nand U204 (N_204,In_713,In_360);
nor U205 (N_205,In_534,In_154);
xnor U206 (N_206,In_180,In_488);
xnor U207 (N_207,In_660,In_442);
nand U208 (N_208,In_4,In_5);
nor U209 (N_209,In_584,In_410);
nand U210 (N_210,In_445,In_177);
xor U211 (N_211,In_27,In_398);
nor U212 (N_212,In_290,In_296);
or U213 (N_213,In_435,In_380);
and U214 (N_214,In_106,In_181);
or U215 (N_215,In_509,In_715);
xor U216 (N_216,In_403,In_193);
or U217 (N_217,In_249,In_130);
xor U218 (N_218,In_93,In_434);
nand U219 (N_219,In_235,In_155);
nor U220 (N_220,In_422,In_385);
nand U221 (N_221,In_343,In_489);
or U222 (N_222,In_405,In_10);
or U223 (N_223,In_52,In_47);
nor U224 (N_224,In_284,In_26);
nor U225 (N_225,In_143,In_158);
nand U226 (N_226,In_354,In_257);
nor U227 (N_227,In_108,In_312);
nor U228 (N_228,In_748,In_25);
nand U229 (N_229,In_473,In_364);
nand U230 (N_230,In_20,In_64);
and U231 (N_231,In_468,In_171);
nor U232 (N_232,In_389,In_733);
xnor U233 (N_233,In_72,In_451);
xnor U234 (N_234,In_593,In_229);
xnor U235 (N_235,In_50,In_261);
nor U236 (N_236,In_379,In_496);
and U237 (N_237,In_425,In_409);
nor U238 (N_238,In_348,In_301);
xnor U239 (N_239,In_342,In_515);
and U240 (N_240,In_234,In_178);
nor U241 (N_241,In_524,In_254);
or U242 (N_242,In_377,In_476);
and U243 (N_243,In_563,In_150);
nor U244 (N_244,In_324,In_304);
xor U245 (N_245,In_384,In_647);
or U246 (N_246,In_700,In_449);
xor U247 (N_247,In_688,In_69);
or U248 (N_248,In_169,In_682);
or U249 (N_249,In_712,In_35);
nor U250 (N_250,In_537,In_57);
nand U251 (N_251,In_63,In_56);
xnor U252 (N_252,In_641,In_484);
xnor U253 (N_253,In_73,In_438);
and U254 (N_254,In_539,In_239);
and U255 (N_255,In_590,In_691);
and U256 (N_256,In_734,In_400);
nor U257 (N_257,In_630,In_136);
or U258 (N_258,In_587,In_535);
and U259 (N_259,In_745,In_22);
nand U260 (N_260,In_135,In_554);
and U261 (N_261,In_217,In_495);
nand U262 (N_262,In_455,In_684);
xnor U263 (N_263,In_485,In_465);
and U264 (N_264,In_194,In_117);
nand U265 (N_265,In_140,In_127);
and U266 (N_266,In_287,In_533);
and U267 (N_267,In_477,In_163);
nor U268 (N_268,In_558,In_448);
and U269 (N_269,In_659,In_514);
nand U270 (N_270,In_605,In_603);
nor U271 (N_271,In_81,In_9);
nand U272 (N_272,In_532,In_189);
nand U273 (N_273,In_200,In_746);
or U274 (N_274,In_480,In_404);
xnor U275 (N_275,In_472,In_661);
nor U276 (N_276,In_622,In_356);
nand U277 (N_277,In_243,In_110);
nor U278 (N_278,In_338,In_638);
or U279 (N_279,In_653,In_541);
nor U280 (N_280,In_670,In_299);
or U281 (N_281,In_530,In_258);
nor U282 (N_282,In_580,In_132);
or U283 (N_283,In_120,In_430);
nor U284 (N_284,In_702,In_565);
and U285 (N_285,In_536,In_431);
nor U286 (N_286,In_62,In_275);
or U287 (N_287,In_528,In_735);
nor U288 (N_288,In_466,In_104);
and U289 (N_289,In_119,In_78);
nor U290 (N_290,In_623,In_315);
nor U291 (N_291,In_245,In_463);
nand U292 (N_292,In_314,In_716);
or U293 (N_293,In_273,In_146);
and U294 (N_294,In_92,In_606);
nor U295 (N_295,In_176,In_699);
nand U296 (N_296,In_694,In_162);
and U297 (N_297,In_125,In_131);
or U298 (N_298,In_685,In_94);
or U299 (N_299,In_625,In_184);
or U300 (N_300,In_246,In_552);
or U301 (N_301,In_206,In_747);
nand U302 (N_302,In_462,In_671);
nor U303 (N_303,In_727,In_624);
nand U304 (N_304,In_407,In_282);
nand U305 (N_305,In_610,In_457);
nand U306 (N_306,In_51,In_204);
nand U307 (N_307,In_506,In_491);
xor U308 (N_308,In_74,In_227);
or U309 (N_309,In_361,In_420);
and U310 (N_310,In_292,In_597);
or U311 (N_311,In_285,In_42);
and U312 (N_312,In_627,In_67);
nand U313 (N_313,In_54,In_644);
or U314 (N_314,In_395,In_675);
nor U315 (N_315,In_510,In_95);
or U316 (N_316,In_43,In_91);
nand U317 (N_317,In_49,In_550);
and U318 (N_318,In_311,In_286);
or U319 (N_319,In_263,In_695);
nor U320 (N_320,In_394,In_662);
xor U321 (N_321,In_441,In_253);
or U322 (N_322,In_698,In_737);
nor U323 (N_323,In_309,In_192);
or U324 (N_324,In_585,In_34);
nand U325 (N_325,In_740,In_650);
and U326 (N_326,In_561,In_714);
nand U327 (N_327,In_686,In_112);
and U328 (N_328,In_601,In_337);
nor U329 (N_329,In_424,In_7);
or U330 (N_330,In_546,In_513);
and U331 (N_331,In_329,In_225);
nand U332 (N_332,In_294,In_46);
nor U333 (N_333,In_0,In_1);
and U334 (N_334,In_655,In_335);
nand U335 (N_335,In_436,In_271);
xnor U336 (N_336,In_570,In_526);
nor U337 (N_337,In_616,In_639);
and U338 (N_338,In_161,In_30);
or U339 (N_339,In_368,In_689);
or U340 (N_340,In_2,In_167);
xnor U341 (N_341,In_500,In_690);
nand U342 (N_342,In_83,In_350);
nand U343 (N_343,In_402,In_90);
or U344 (N_344,In_654,In_577);
nand U345 (N_345,In_519,In_297);
xnor U346 (N_346,In_205,In_545);
and U347 (N_347,In_707,In_673);
nand U348 (N_348,In_121,In_464);
nor U349 (N_349,In_512,In_126);
nor U350 (N_350,In_651,In_236);
nand U351 (N_351,In_544,In_667);
or U352 (N_352,In_365,In_244);
nor U353 (N_353,In_588,In_224);
nand U354 (N_354,In_572,In_326);
and U355 (N_355,In_24,In_516);
and U356 (N_356,In_48,In_222);
or U357 (N_357,In_340,In_722);
nor U358 (N_358,In_251,In_522);
nand U359 (N_359,In_581,In_31);
nand U360 (N_360,In_196,In_80);
or U361 (N_361,In_432,In_717);
nor U362 (N_362,In_672,In_391);
and U363 (N_363,In_568,In_705);
nor U364 (N_364,In_15,In_170);
nand U365 (N_365,In_346,In_152);
nand U366 (N_366,In_198,In_259);
and U367 (N_367,In_96,In_411);
nor U368 (N_368,In_114,In_139);
nor U369 (N_369,In_471,In_393);
xor U370 (N_370,In_677,In_582);
or U371 (N_371,In_446,In_230);
and U372 (N_372,In_166,In_363);
or U373 (N_373,In_216,In_75);
or U374 (N_374,In_358,In_742);
and U375 (N_375,In_166,In_158);
nand U376 (N_376,In_387,In_479);
nand U377 (N_377,In_749,In_543);
and U378 (N_378,In_2,In_497);
nand U379 (N_379,In_343,In_702);
and U380 (N_380,In_494,In_460);
or U381 (N_381,In_119,In_511);
nand U382 (N_382,In_515,In_278);
or U383 (N_383,In_457,In_480);
or U384 (N_384,In_98,In_57);
xnor U385 (N_385,In_476,In_139);
or U386 (N_386,In_657,In_579);
nand U387 (N_387,In_245,In_695);
nand U388 (N_388,In_335,In_611);
and U389 (N_389,In_288,In_463);
nor U390 (N_390,In_279,In_535);
and U391 (N_391,In_348,In_528);
nor U392 (N_392,In_749,In_421);
xor U393 (N_393,In_746,In_89);
and U394 (N_394,In_655,In_330);
and U395 (N_395,In_265,In_198);
nand U396 (N_396,In_318,In_147);
nor U397 (N_397,In_272,In_486);
nand U398 (N_398,In_712,In_20);
and U399 (N_399,In_477,In_57);
xor U400 (N_400,In_58,In_112);
nand U401 (N_401,In_351,In_13);
or U402 (N_402,In_565,In_271);
and U403 (N_403,In_633,In_439);
nand U404 (N_404,In_98,In_592);
and U405 (N_405,In_702,In_149);
nand U406 (N_406,In_439,In_36);
and U407 (N_407,In_291,In_727);
nor U408 (N_408,In_181,In_703);
nand U409 (N_409,In_380,In_567);
nand U410 (N_410,In_633,In_229);
xnor U411 (N_411,In_397,In_148);
and U412 (N_412,In_678,In_558);
nor U413 (N_413,In_437,In_421);
nor U414 (N_414,In_565,In_666);
or U415 (N_415,In_529,In_230);
nand U416 (N_416,In_94,In_414);
nand U417 (N_417,In_163,In_716);
nand U418 (N_418,In_311,In_410);
nand U419 (N_419,In_93,In_506);
xor U420 (N_420,In_399,In_745);
and U421 (N_421,In_475,In_165);
xor U422 (N_422,In_260,In_626);
nor U423 (N_423,In_177,In_535);
or U424 (N_424,In_336,In_294);
and U425 (N_425,In_596,In_250);
nor U426 (N_426,In_581,In_377);
xnor U427 (N_427,In_186,In_513);
nor U428 (N_428,In_281,In_646);
xnor U429 (N_429,In_191,In_724);
and U430 (N_430,In_298,In_326);
and U431 (N_431,In_233,In_116);
xor U432 (N_432,In_608,In_44);
and U433 (N_433,In_598,In_18);
nand U434 (N_434,In_511,In_206);
nand U435 (N_435,In_626,In_223);
nand U436 (N_436,In_554,In_346);
or U437 (N_437,In_404,In_432);
or U438 (N_438,In_741,In_156);
nor U439 (N_439,In_738,In_526);
nor U440 (N_440,In_365,In_371);
nor U441 (N_441,In_251,In_587);
nand U442 (N_442,In_580,In_221);
nand U443 (N_443,In_75,In_647);
or U444 (N_444,In_48,In_203);
nand U445 (N_445,In_595,In_473);
nor U446 (N_446,In_5,In_601);
nand U447 (N_447,In_560,In_35);
or U448 (N_448,In_564,In_649);
and U449 (N_449,In_359,In_519);
and U450 (N_450,In_226,In_479);
nand U451 (N_451,In_96,In_589);
nand U452 (N_452,In_490,In_272);
or U453 (N_453,In_457,In_119);
nand U454 (N_454,In_398,In_697);
nand U455 (N_455,In_304,In_493);
nand U456 (N_456,In_228,In_541);
nand U457 (N_457,In_581,In_121);
or U458 (N_458,In_340,In_335);
nand U459 (N_459,In_149,In_415);
nor U460 (N_460,In_649,In_736);
or U461 (N_461,In_415,In_12);
nand U462 (N_462,In_301,In_634);
and U463 (N_463,In_90,In_558);
or U464 (N_464,In_547,In_387);
xnor U465 (N_465,In_198,In_504);
xnor U466 (N_466,In_6,In_414);
nor U467 (N_467,In_656,In_93);
or U468 (N_468,In_545,In_607);
nand U469 (N_469,In_110,In_156);
nor U470 (N_470,In_644,In_630);
or U471 (N_471,In_433,In_424);
nor U472 (N_472,In_660,In_587);
and U473 (N_473,In_213,In_358);
nor U474 (N_474,In_641,In_377);
or U475 (N_475,In_394,In_106);
nor U476 (N_476,In_697,In_93);
nor U477 (N_477,In_45,In_597);
nor U478 (N_478,In_149,In_524);
nand U479 (N_479,In_476,In_535);
nand U480 (N_480,In_536,In_166);
or U481 (N_481,In_315,In_399);
nand U482 (N_482,In_260,In_516);
or U483 (N_483,In_446,In_417);
nor U484 (N_484,In_234,In_26);
or U485 (N_485,In_364,In_281);
or U486 (N_486,In_400,In_559);
or U487 (N_487,In_319,In_391);
nor U488 (N_488,In_46,In_272);
nand U489 (N_489,In_260,In_181);
nand U490 (N_490,In_437,In_673);
nor U491 (N_491,In_549,In_595);
nand U492 (N_492,In_227,In_46);
nand U493 (N_493,In_174,In_514);
or U494 (N_494,In_433,In_320);
xor U495 (N_495,In_307,In_429);
nand U496 (N_496,In_203,In_526);
nand U497 (N_497,In_496,In_119);
nor U498 (N_498,In_701,In_331);
nand U499 (N_499,In_559,In_136);
nor U500 (N_500,In_703,In_670);
or U501 (N_501,In_591,In_144);
nor U502 (N_502,In_451,In_290);
xor U503 (N_503,In_106,In_101);
and U504 (N_504,In_350,In_496);
or U505 (N_505,In_286,In_366);
xnor U506 (N_506,In_58,In_30);
nor U507 (N_507,In_640,In_306);
and U508 (N_508,In_276,In_304);
nand U509 (N_509,In_128,In_312);
nand U510 (N_510,In_36,In_320);
nand U511 (N_511,In_747,In_120);
nor U512 (N_512,In_10,In_171);
nor U513 (N_513,In_68,In_71);
nor U514 (N_514,In_660,In_369);
and U515 (N_515,In_692,In_507);
nor U516 (N_516,In_726,In_18);
nor U517 (N_517,In_653,In_693);
nand U518 (N_518,In_727,In_425);
nor U519 (N_519,In_583,In_439);
nand U520 (N_520,In_543,In_568);
and U521 (N_521,In_568,In_337);
or U522 (N_522,In_677,In_498);
or U523 (N_523,In_664,In_197);
xnor U524 (N_524,In_720,In_128);
and U525 (N_525,In_306,In_26);
nand U526 (N_526,In_17,In_441);
nor U527 (N_527,In_330,In_70);
or U528 (N_528,In_169,In_295);
and U529 (N_529,In_577,In_488);
or U530 (N_530,In_285,In_211);
and U531 (N_531,In_641,In_243);
xor U532 (N_532,In_578,In_526);
nor U533 (N_533,In_690,In_71);
nand U534 (N_534,In_12,In_163);
and U535 (N_535,In_200,In_440);
nand U536 (N_536,In_547,In_612);
and U537 (N_537,In_226,In_669);
nor U538 (N_538,In_744,In_465);
nor U539 (N_539,In_22,In_32);
xnor U540 (N_540,In_605,In_38);
nand U541 (N_541,In_536,In_111);
xnor U542 (N_542,In_450,In_721);
and U543 (N_543,In_326,In_185);
and U544 (N_544,In_294,In_598);
nand U545 (N_545,In_269,In_74);
or U546 (N_546,In_304,In_194);
nor U547 (N_547,In_27,In_672);
xnor U548 (N_548,In_87,In_684);
or U549 (N_549,In_548,In_103);
nand U550 (N_550,In_440,In_729);
and U551 (N_551,In_39,In_20);
nand U552 (N_552,In_485,In_78);
or U553 (N_553,In_3,In_340);
nor U554 (N_554,In_97,In_118);
nand U555 (N_555,In_193,In_68);
or U556 (N_556,In_339,In_163);
or U557 (N_557,In_100,In_84);
or U558 (N_558,In_254,In_216);
xor U559 (N_559,In_639,In_315);
nor U560 (N_560,In_140,In_633);
and U561 (N_561,In_135,In_208);
nor U562 (N_562,In_422,In_541);
or U563 (N_563,In_199,In_22);
or U564 (N_564,In_31,In_155);
nand U565 (N_565,In_53,In_524);
and U566 (N_566,In_654,In_162);
nor U567 (N_567,In_365,In_250);
nor U568 (N_568,In_223,In_83);
or U569 (N_569,In_503,In_586);
or U570 (N_570,In_207,In_361);
xor U571 (N_571,In_424,In_518);
nor U572 (N_572,In_444,In_425);
nor U573 (N_573,In_705,In_486);
nor U574 (N_574,In_408,In_260);
nor U575 (N_575,In_143,In_120);
nand U576 (N_576,In_429,In_562);
nand U577 (N_577,In_233,In_566);
or U578 (N_578,In_675,In_714);
nand U579 (N_579,In_419,In_33);
nor U580 (N_580,In_406,In_606);
and U581 (N_581,In_382,In_284);
and U582 (N_582,In_291,In_256);
nor U583 (N_583,In_302,In_436);
and U584 (N_584,In_734,In_310);
nand U585 (N_585,In_743,In_620);
xnor U586 (N_586,In_599,In_149);
and U587 (N_587,In_126,In_572);
nor U588 (N_588,In_113,In_332);
or U589 (N_589,In_648,In_43);
or U590 (N_590,In_237,In_117);
or U591 (N_591,In_704,In_441);
nand U592 (N_592,In_78,In_333);
or U593 (N_593,In_254,In_407);
nand U594 (N_594,In_718,In_301);
and U595 (N_595,In_432,In_538);
and U596 (N_596,In_240,In_222);
nor U597 (N_597,In_531,In_63);
or U598 (N_598,In_719,In_141);
or U599 (N_599,In_405,In_217);
or U600 (N_600,In_23,In_409);
nand U601 (N_601,In_79,In_6);
nor U602 (N_602,In_357,In_625);
nor U603 (N_603,In_641,In_176);
or U604 (N_604,In_607,In_188);
nand U605 (N_605,In_614,In_523);
nand U606 (N_606,In_445,In_681);
or U607 (N_607,In_72,In_515);
nand U608 (N_608,In_349,In_609);
nor U609 (N_609,In_277,In_113);
nand U610 (N_610,In_181,In_397);
and U611 (N_611,In_575,In_708);
and U612 (N_612,In_366,In_64);
nor U613 (N_613,In_423,In_736);
xor U614 (N_614,In_433,In_79);
or U615 (N_615,In_746,In_385);
nor U616 (N_616,In_291,In_651);
or U617 (N_617,In_712,In_402);
nand U618 (N_618,In_241,In_42);
nand U619 (N_619,In_320,In_401);
nand U620 (N_620,In_634,In_413);
nor U621 (N_621,In_340,In_527);
nor U622 (N_622,In_598,In_460);
or U623 (N_623,In_245,In_265);
or U624 (N_624,In_123,In_721);
nor U625 (N_625,In_407,In_258);
nor U626 (N_626,In_147,In_270);
nand U627 (N_627,In_181,In_549);
nor U628 (N_628,In_183,In_476);
or U629 (N_629,In_130,In_572);
nand U630 (N_630,In_104,In_632);
nand U631 (N_631,In_635,In_94);
xor U632 (N_632,In_107,In_632);
nand U633 (N_633,In_648,In_190);
or U634 (N_634,In_111,In_235);
and U635 (N_635,In_652,In_357);
nor U636 (N_636,In_250,In_614);
nand U637 (N_637,In_367,In_201);
and U638 (N_638,In_587,In_227);
and U639 (N_639,In_99,In_676);
nor U640 (N_640,In_405,In_714);
nor U641 (N_641,In_173,In_591);
or U642 (N_642,In_447,In_632);
nand U643 (N_643,In_745,In_521);
and U644 (N_644,In_242,In_444);
xor U645 (N_645,In_663,In_311);
and U646 (N_646,In_286,In_171);
nand U647 (N_647,In_393,In_702);
and U648 (N_648,In_652,In_444);
and U649 (N_649,In_153,In_665);
and U650 (N_650,In_385,In_112);
and U651 (N_651,In_270,In_390);
nor U652 (N_652,In_8,In_305);
or U653 (N_653,In_485,In_724);
nor U654 (N_654,In_227,In_346);
or U655 (N_655,In_192,In_665);
xor U656 (N_656,In_367,In_177);
xor U657 (N_657,In_453,In_558);
xor U658 (N_658,In_66,In_154);
or U659 (N_659,In_318,In_378);
and U660 (N_660,In_155,In_426);
nand U661 (N_661,In_515,In_192);
nor U662 (N_662,In_416,In_51);
nand U663 (N_663,In_33,In_601);
nor U664 (N_664,In_107,In_156);
nor U665 (N_665,In_537,In_296);
or U666 (N_666,In_125,In_177);
nor U667 (N_667,In_312,In_302);
or U668 (N_668,In_552,In_243);
xnor U669 (N_669,In_573,In_564);
nor U670 (N_670,In_518,In_587);
or U671 (N_671,In_687,In_294);
or U672 (N_672,In_133,In_290);
nor U673 (N_673,In_494,In_67);
or U674 (N_674,In_28,In_415);
xor U675 (N_675,In_97,In_27);
and U676 (N_676,In_445,In_749);
and U677 (N_677,In_335,In_495);
and U678 (N_678,In_11,In_121);
nand U679 (N_679,In_627,In_508);
or U680 (N_680,In_35,In_332);
and U681 (N_681,In_173,In_514);
and U682 (N_682,In_549,In_643);
nand U683 (N_683,In_633,In_211);
or U684 (N_684,In_189,In_101);
nand U685 (N_685,In_474,In_673);
and U686 (N_686,In_589,In_674);
nor U687 (N_687,In_596,In_352);
nand U688 (N_688,In_222,In_735);
nor U689 (N_689,In_341,In_85);
nand U690 (N_690,In_520,In_373);
nand U691 (N_691,In_502,In_334);
nor U692 (N_692,In_744,In_523);
xor U693 (N_693,In_370,In_374);
or U694 (N_694,In_740,In_138);
nor U695 (N_695,In_259,In_465);
nor U696 (N_696,In_181,In_412);
and U697 (N_697,In_222,In_172);
xnor U698 (N_698,In_683,In_49);
and U699 (N_699,In_79,In_416);
or U700 (N_700,In_413,In_49);
and U701 (N_701,In_412,In_497);
or U702 (N_702,In_641,In_608);
or U703 (N_703,In_387,In_148);
and U704 (N_704,In_519,In_15);
nor U705 (N_705,In_210,In_295);
xor U706 (N_706,In_38,In_308);
nand U707 (N_707,In_560,In_371);
nor U708 (N_708,In_631,In_732);
nand U709 (N_709,In_79,In_467);
nor U710 (N_710,In_27,In_318);
nor U711 (N_711,In_733,In_266);
and U712 (N_712,In_455,In_434);
nor U713 (N_713,In_601,In_516);
and U714 (N_714,In_673,In_623);
and U715 (N_715,In_105,In_441);
or U716 (N_716,In_597,In_330);
nand U717 (N_717,In_342,In_130);
or U718 (N_718,In_93,In_407);
xor U719 (N_719,In_176,In_565);
and U720 (N_720,In_404,In_177);
and U721 (N_721,In_197,In_18);
and U722 (N_722,In_385,In_414);
or U723 (N_723,In_538,In_463);
xnor U724 (N_724,In_428,In_10);
nor U725 (N_725,In_602,In_86);
and U726 (N_726,In_107,In_184);
nor U727 (N_727,In_718,In_442);
and U728 (N_728,In_57,In_425);
nand U729 (N_729,In_38,In_134);
or U730 (N_730,In_312,In_437);
nor U731 (N_731,In_467,In_167);
and U732 (N_732,In_112,In_306);
and U733 (N_733,In_132,In_537);
nor U734 (N_734,In_499,In_713);
and U735 (N_735,In_401,In_555);
nor U736 (N_736,In_242,In_576);
or U737 (N_737,In_723,In_282);
nand U738 (N_738,In_580,In_507);
nor U739 (N_739,In_104,In_472);
or U740 (N_740,In_225,In_23);
nand U741 (N_741,In_464,In_534);
nand U742 (N_742,In_580,In_445);
nand U743 (N_743,In_273,In_602);
nor U744 (N_744,In_574,In_561);
nor U745 (N_745,In_637,In_353);
and U746 (N_746,In_297,In_178);
and U747 (N_747,In_600,In_651);
and U748 (N_748,In_638,In_246);
nand U749 (N_749,In_284,In_510);
nand U750 (N_750,In_429,In_366);
or U751 (N_751,In_7,In_740);
nor U752 (N_752,In_526,In_216);
or U753 (N_753,In_375,In_502);
and U754 (N_754,In_705,In_269);
nor U755 (N_755,In_442,In_261);
and U756 (N_756,In_56,In_341);
nand U757 (N_757,In_566,In_667);
and U758 (N_758,In_577,In_58);
nand U759 (N_759,In_293,In_151);
and U760 (N_760,In_137,In_249);
or U761 (N_761,In_668,In_243);
nand U762 (N_762,In_644,In_262);
nor U763 (N_763,In_31,In_393);
and U764 (N_764,In_199,In_738);
nand U765 (N_765,In_582,In_48);
xor U766 (N_766,In_662,In_34);
or U767 (N_767,In_111,In_481);
or U768 (N_768,In_650,In_581);
nor U769 (N_769,In_65,In_193);
or U770 (N_770,In_489,In_253);
nor U771 (N_771,In_468,In_304);
and U772 (N_772,In_416,In_126);
nand U773 (N_773,In_304,In_249);
nand U774 (N_774,In_734,In_550);
nand U775 (N_775,In_192,In_0);
nand U776 (N_776,In_18,In_488);
or U777 (N_777,In_390,In_52);
or U778 (N_778,In_234,In_256);
and U779 (N_779,In_375,In_531);
xor U780 (N_780,In_651,In_44);
xor U781 (N_781,In_424,In_511);
nand U782 (N_782,In_628,In_694);
nand U783 (N_783,In_250,In_90);
and U784 (N_784,In_620,In_47);
nand U785 (N_785,In_150,In_105);
nand U786 (N_786,In_364,In_645);
nand U787 (N_787,In_704,In_244);
nand U788 (N_788,In_599,In_523);
and U789 (N_789,In_258,In_515);
or U790 (N_790,In_416,In_252);
nand U791 (N_791,In_58,In_39);
nand U792 (N_792,In_404,In_135);
nor U793 (N_793,In_209,In_60);
and U794 (N_794,In_20,In_517);
nand U795 (N_795,In_438,In_380);
nor U796 (N_796,In_719,In_380);
and U797 (N_797,In_430,In_722);
or U798 (N_798,In_196,In_729);
xnor U799 (N_799,In_264,In_97);
or U800 (N_800,In_738,In_372);
and U801 (N_801,In_724,In_222);
nand U802 (N_802,In_404,In_304);
or U803 (N_803,In_470,In_711);
nand U804 (N_804,In_447,In_240);
nand U805 (N_805,In_408,In_693);
nor U806 (N_806,In_688,In_731);
nand U807 (N_807,In_486,In_745);
nor U808 (N_808,In_437,In_386);
or U809 (N_809,In_206,In_5);
or U810 (N_810,In_253,In_504);
nor U811 (N_811,In_31,In_451);
nor U812 (N_812,In_77,In_371);
nand U813 (N_813,In_610,In_620);
and U814 (N_814,In_517,In_651);
nor U815 (N_815,In_528,In_315);
xnor U816 (N_816,In_471,In_517);
xnor U817 (N_817,In_639,In_481);
nand U818 (N_818,In_623,In_261);
or U819 (N_819,In_192,In_481);
nand U820 (N_820,In_320,In_740);
and U821 (N_821,In_720,In_348);
or U822 (N_822,In_576,In_516);
or U823 (N_823,In_564,In_478);
nand U824 (N_824,In_675,In_560);
or U825 (N_825,In_583,In_392);
nor U826 (N_826,In_581,In_571);
nor U827 (N_827,In_495,In_246);
nor U828 (N_828,In_147,In_582);
and U829 (N_829,In_492,In_715);
nor U830 (N_830,In_235,In_218);
and U831 (N_831,In_20,In_131);
or U832 (N_832,In_240,In_519);
or U833 (N_833,In_584,In_44);
and U834 (N_834,In_28,In_194);
nor U835 (N_835,In_563,In_7);
xor U836 (N_836,In_6,In_311);
nor U837 (N_837,In_300,In_92);
xor U838 (N_838,In_112,In_120);
and U839 (N_839,In_208,In_407);
nand U840 (N_840,In_681,In_344);
and U841 (N_841,In_279,In_620);
nand U842 (N_842,In_736,In_644);
and U843 (N_843,In_662,In_713);
or U844 (N_844,In_220,In_194);
xnor U845 (N_845,In_530,In_499);
or U846 (N_846,In_510,In_493);
and U847 (N_847,In_245,In_78);
nor U848 (N_848,In_300,In_22);
xor U849 (N_849,In_651,In_196);
nand U850 (N_850,In_269,In_691);
and U851 (N_851,In_600,In_501);
and U852 (N_852,In_11,In_4);
nand U853 (N_853,In_143,In_567);
nor U854 (N_854,In_2,In_363);
nor U855 (N_855,In_198,In_297);
and U856 (N_856,In_206,In_717);
or U857 (N_857,In_461,In_618);
nand U858 (N_858,In_180,In_634);
nand U859 (N_859,In_716,In_97);
and U860 (N_860,In_379,In_198);
nor U861 (N_861,In_40,In_22);
nor U862 (N_862,In_443,In_34);
xor U863 (N_863,In_523,In_190);
xor U864 (N_864,In_0,In_514);
and U865 (N_865,In_282,In_179);
nand U866 (N_866,In_476,In_111);
xnor U867 (N_867,In_352,In_452);
and U868 (N_868,In_9,In_463);
nor U869 (N_869,In_112,In_491);
nand U870 (N_870,In_508,In_701);
nand U871 (N_871,In_14,In_715);
or U872 (N_872,In_552,In_346);
nor U873 (N_873,In_508,In_438);
xnor U874 (N_874,In_551,In_396);
xor U875 (N_875,In_543,In_625);
xnor U876 (N_876,In_219,In_186);
nand U877 (N_877,In_82,In_34);
or U878 (N_878,In_457,In_689);
and U879 (N_879,In_463,In_183);
or U880 (N_880,In_444,In_25);
nor U881 (N_881,In_594,In_610);
nor U882 (N_882,In_698,In_402);
and U883 (N_883,In_747,In_110);
xor U884 (N_884,In_69,In_351);
nor U885 (N_885,In_114,In_307);
nand U886 (N_886,In_158,In_542);
nand U887 (N_887,In_279,In_579);
nand U888 (N_888,In_154,In_83);
nand U889 (N_889,In_350,In_633);
nand U890 (N_890,In_600,In_499);
xnor U891 (N_891,In_531,In_208);
and U892 (N_892,In_505,In_167);
nand U893 (N_893,In_531,In_739);
and U894 (N_894,In_69,In_412);
nor U895 (N_895,In_618,In_84);
nand U896 (N_896,In_206,In_342);
nand U897 (N_897,In_432,In_255);
and U898 (N_898,In_730,In_14);
nand U899 (N_899,In_498,In_193);
nand U900 (N_900,In_600,In_74);
or U901 (N_901,In_680,In_135);
xnor U902 (N_902,In_702,In_362);
nand U903 (N_903,In_679,In_674);
nand U904 (N_904,In_641,In_328);
and U905 (N_905,In_78,In_516);
nor U906 (N_906,In_193,In_482);
nor U907 (N_907,In_657,In_235);
or U908 (N_908,In_100,In_602);
and U909 (N_909,In_589,In_130);
and U910 (N_910,In_87,In_178);
nand U911 (N_911,In_450,In_381);
nand U912 (N_912,In_538,In_200);
and U913 (N_913,In_86,In_735);
or U914 (N_914,In_130,In_631);
nand U915 (N_915,In_710,In_237);
or U916 (N_916,In_659,In_99);
nand U917 (N_917,In_346,In_658);
or U918 (N_918,In_53,In_282);
and U919 (N_919,In_666,In_396);
and U920 (N_920,In_579,In_513);
and U921 (N_921,In_659,In_651);
nand U922 (N_922,In_237,In_187);
nand U923 (N_923,In_528,In_644);
or U924 (N_924,In_412,In_740);
nand U925 (N_925,In_182,In_280);
nand U926 (N_926,In_124,In_474);
and U927 (N_927,In_576,In_96);
or U928 (N_928,In_566,In_82);
nor U929 (N_929,In_373,In_122);
nor U930 (N_930,In_596,In_636);
nor U931 (N_931,In_39,In_498);
nand U932 (N_932,In_330,In_376);
nand U933 (N_933,In_727,In_679);
or U934 (N_934,In_522,In_736);
nor U935 (N_935,In_460,In_501);
and U936 (N_936,In_275,In_90);
nand U937 (N_937,In_638,In_110);
nand U938 (N_938,In_301,In_745);
nor U939 (N_939,In_287,In_70);
nand U940 (N_940,In_107,In_702);
nor U941 (N_941,In_520,In_713);
and U942 (N_942,In_445,In_90);
and U943 (N_943,In_326,In_500);
nand U944 (N_944,In_333,In_605);
nor U945 (N_945,In_41,In_139);
nand U946 (N_946,In_251,In_322);
or U947 (N_947,In_395,In_377);
xnor U948 (N_948,In_301,In_451);
and U949 (N_949,In_650,In_276);
nand U950 (N_950,In_65,In_12);
or U951 (N_951,In_171,In_624);
and U952 (N_952,In_345,In_87);
nor U953 (N_953,In_445,In_380);
xnor U954 (N_954,In_239,In_554);
nand U955 (N_955,In_737,In_387);
nand U956 (N_956,In_546,In_718);
nor U957 (N_957,In_320,In_340);
or U958 (N_958,In_132,In_240);
and U959 (N_959,In_605,In_620);
nor U960 (N_960,In_83,In_288);
or U961 (N_961,In_196,In_252);
nor U962 (N_962,In_99,In_478);
nand U963 (N_963,In_602,In_360);
nor U964 (N_964,In_498,In_627);
xor U965 (N_965,In_290,In_682);
and U966 (N_966,In_335,In_275);
nand U967 (N_967,In_357,In_286);
nand U968 (N_968,In_510,In_274);
or U969 (N_969,In_731,In_608);
or U970 (N_970,In_384,In_2);
nand U971 (N_971,In_683,In_276);
nor U972 (N_972,In_259,In_610);
or U973 (N_973,In_699,In_547);
nor U974 (N_974,In_97,In_738);
xor U975 (N_975,In_82,In_309);
nor U976 (N_976,In_717,In_652);
xnor U977 (N_977,In_641,In_178);
xnor U978 (N_978,In_680,In_140);
nor U979 (N_979,In_468,In_631);
nor U980 (N_980,In_608,In_671);
or U981 (N_981,In_154,In_259);
xor U982 (N_982,In_181,In_518);
nand U983 (N_983,In_735,In_404);
nor U984 (N_984,In_470,In_708);
nor U985 (N_985,In_78,In_584);
or U986 (N_986,In_28,In_370);
nand U987 (N_987,In_248,In_208);
nand U988 (N_988,In_431,In_717);
and U989 (N_989,In_340,In_108);
nor U990 (N_990,In_398,In_714);
and U991 (N_991,In_533,In_324);
and U992 (N_992,In_4,In_417);
xor U993 (N_993,In_216,In_736);
nand U994 (N_994,In_552,In_678);
or U995 (N_995,In_673,In_62);
and U996 (N_996,In_457,In_31);
and U997 (N_997,In_682,In_614);
or U998 (N_998,In_81,In_349);
or U999 (N_999,In_517,In_75);
and U1000 (N_1000,N_53,N_167);
nand U1001 (N_1001,N_65,N_413);
or U1002 (N_1002,N_49,N_741);
and U1003 (N_1003,N_536,N_238);
or U1004 (N_1004,N_254,N_856);
or U1005 (N_1005,N_232,N_542);
or U1006 (N_1006,N_988,N_250);
xnor U1007 (N_1007,N_756,N_316);
and U1008 (N_1008,N_554,N_278);
or U1009 (N_1009,N_269,N_469);
nor U1010 (N_1010,N_858,N_173);
or U1011 (N_1011,N_146,N_932);
or U1012 (N_1012,N_15,N_527);
or U1013 (N_1013,N_255,N_959);
and U1014 (N_1014,N_490,N_234);
xnor U1015 (N_1015,N_514,N_508);
or U1016 (N_1016,N_279,N_248);
or U1017 (N_1017,N_775,N_732);
nand U1018 (N_1018,N_23,N_135);
nand U1019 (N_1019,N_894,N_540);
nor U1020 (N_1020,N_347,N_320);
nand U1021 (N_1021,N_130,N_193);
nand U1022 (N_1022,N_131,N_307);
nor U1023 (N_1023,N_369,N_571);
or U1024 (N_1024,N_640,N_925);
xor U1025 (N_1025,N_312,N_844);
or U1026 (N_1026,N_346,N_681);
or U1027 (N_1027,N_659,N_872);
nor U1028 (N_1028,N_475,N_372);
nor U1029 (N_1029,N_874,N_902);
or U1030 (N_1030,N_522,N_870);
or U1031 (N_1031,N_612,N_147);
nor U1032 (N_1032,N_271,N_914);
and U1033 (N_1033,N_938,N_877);
and U1034 (N_1034,N_976,N_333);
and U1035 (N_1035,N_133,N_543);
nor U1036 (N_1036,N_412,N_208);
and U1037 (N_1037,N_648,N_662);
nand U1038 (N_1038,N_275,N_785);
and U1039 (N_1039,N_991,N_348);
or U1040 (N_1040,N_229,N_647);
or U1041 (N_1041,N_887,N_898);
or U1042 (N_1042,N_521,N_551);
nor U1043 (N_1043,N_467,N_471);
or U1044 (N_1044,N_761,N_128);
and U1045 (N_1045,N_152,N_780);
nor U1046 (N_1046,N_450,N_159);
or U1047 (N_1047,N_60,N_441);
nor U1048 (N_1048,N_240,N_18);
and U1049 (N_1049,N_396,N_701);
and U1050 (N_1050,N_237,N_893);
and U1051 (N_1051,N_678,N_896);
and U1052 (N_1052,N_337,N_544);
or U1053 (N_1053,N_686,N_883);
nand U1054 (N_1054,N_206,N_903);
nand U1055 (N_1055,N_710,N_968);
nand U1056 (N_1056,N_7,N_297);
and U1057 (N_1057,N_364,N_804);
nand U1058 (N_1058,N_38,N_14);
nor U1059 (N_1059,N_688,N_504);
or U1060 (N_1060,N_430,N_443);
xnor U1061 (N_1061,N_773,N_358);
or U1062 (N_1062,N_731,N_470);
nand U1063 (N_1063,N_538,N_917);
and U1064 (N_1064,N_292,N_267);
nand U1065 (N_1065,N_264,N_162);
and U1066 (N_1066,N_194,N_165);
or U1067 (N_1067,N_454,N_217);
nor U1068 (N_1068,N_112,N_918);
nor U1069 (N_1069,N_17,N_27);
and U1070 (N_1070,N_599,N_825);
and U1071 (N_1071,N_954,N_286);
nor U1072 (N_1072,N_367,N_707);
or U1073 (N_1073,N_318,N_740);
or U1074 (N_1074,N_998,N_24);
or U1075 (N_1075,N_357,N_709);
nand U1076 (N_1076,N_848,N_510);
xnor U1077 (N_1077,N_853,N_805);
and U1078 (N_1078,N_936,N_205);
and U1079 (N_1079,N_990,N_826);
nor U1080 (N_1080,N_663,N_399);
nor U1081 (N_1081,N_45,N_493);
or U1082 (N_1082,N_488,N_572);
or U1083 (N_1083,N_892,N_733);
nor U1084 (N_1084,N_134,N_594);
nor U1085 (N_1085,N_174,N_287);
nand U1086 (N_1086,N_905,N_272);
and U1087 (N_1087,N_718,N_483);
nor U1088 (N_1088,N_180,N_717);
nand U1089 (N_1089,N_886,N_719);
nand U1090 (N_1090,N_751,N_580);
and U1091 (N_1091,N_379,N_632);
nor U1092 (N_1092,N_880,N_288);
nor U1093 (N_1093,N_639,N_523);
or U1094 (N_1094,N_949,N_285);
and U1095 (N_1095,N_728,N_608);
and U1096 (N_1096,N_373,N_378);
and U1097 (N_1097,N_142,N_314);
nor U1098 (N_1098,N_702,N_830);
nand U1099 (N_1099,N_303,N_416);
or U1100 (N_1100,N_43,N_214);
and U1101 (N_1101,N_813,N_164);
nor U1102 (N_1102,N_985,N_342);
nor U1103 (N_1103,N_793,N_634);
or U1104 (N_1104,N_111,N_439);
nor U1105 (N_1105,N_509,N_68);
and U1106 (N_1106,N_924,N_744);
nand U1107 (N_1107,N_74,N_6);
and U1108 (N_1108,N_435,N_777);
and U1109 (N_1109,N_228,N_85);
xor U1110 (N_1110,N_970,N_419);
xnor U1111 (N_1111,N_852,N_136);
nor U1112 (N_1112,N_245,N_930);
and U1113 (N_1113,N_166,N_101);
nand U1114 (N_1114,N_485,N_115);
and U1115 (N_1115,N_800,N_106);
and U1116 (N_1116,N_444,N_670);
and U1117 (N_1117,N_125,N_195);
and U1118 (N_1118,N_891,N_54);
or U1119 (N_1119,N_80,N_789);
xnor U1120 (N_1120,N_315,N_81);
or U1121 (N_1121,N_993,N_96);
nand U1122 (N_1122,N_846,N_550);
nand U1123 (N_1123,N_616,N_218);
nor U1124 (N_1124,N_646,N_332);
or U1125 (N_1125,N_463,N_713);
and U1126 (N_1126,N_834,N_452);
and U1127 (N_1127,N_477,N_197);
nand U1128 (N_1128,N_899,N_325);
xnor U1129 (N_1129,N_618,N_298);
or U1130 (N_1130,N_704,N_570);
or U1131 (N_1131,N_941,N_840);
nor U1132 (N_1132,N_155,N_847);
xnor U1133 (N_1133,N_273,N_423);
and U1134 (N_1134,N_869,N_171);
xnor U1135 (N_1135,N_620,N_839);
and U1136 (N_1136,N_952,N_829);
and U1137 (N_1137,N_909,N_482);
and U1138 (N_1138,N_185,N_446);
or U1139 (N_1139,N_35,N_625);
or U1140 (N_1140,N_613,N_922);
and U1141 (N_1141,N_951,N_345);
nand U1142 (N_1142,N_820,N_651);
and U1143 (N_1143,N_407,N_790);
nand U1144 (N_1144,N_355,N_884);
or U1145 (N_1145,N_833,N_803);
or U1146 (N_1146,N_807,N_335);
nor U1147 (N_1147,N_457,N_486);
or U1148 (N_1148,N_923,N_52);
or U1149 (N_1149,N_188,N_994);
and U1150 (N_1150,N_986,N_974);
nor U1151 (N_1151,N_199,N_593);
nor U1152 (N_1152,N_432,N_311);
nand U1153 (N_1153,N_811,N_461);
nor U1154 (N_1154,N_698,N_867);
or U1155 (N_1155,N_939,N_817);
nor U1156 (N_1156,N_151,N_411);
and U1157 (N_1157,N_402,N_445);
and U1158 (N_1158,N_908,N_674);
and U1159 (N_1159,N_759,N_97);
or U1160 (N_1160,N_32,N_462);
nor U1161 (N_1161,N_82,N_643);
nand U1162 (N_1162,N_502,N_601);
nand U1163 (N_1163,N_243,N_211);
and U1164 (N_1164,N_397,N_582);
nand U1165 (N_1165,N_221,N_108);
or U1166 (N_1166,N_61,N_263);
or U1167 (N_1167,N_177,N_530);
nor U1168 (N_1168,N_531,N_661);
nand U1169 (N_1169,N_276,N_414);
nor U1170 (N_1170,N_353,N_849);
xor U1171 (N_1171,N_799,N_226);
nand U1172 (N_1172,N_553,N_109);
nand U1173 (N_1173,N_683,N_447);
and U1174 (N_1174,N_972,N_11);
and U1175 (N_1175,N_695,N_390);
and U1176 (N_1176,N_202,N_566);
nand U1177 (N_1177,N_119,N_779);
xnor U1178 (N_1178,N_699,N_845);
or U1179 (N_1179,N_516,N_809);
or U1180 (N_1180,N_89,N_274);
or U1181 (N_1181,N_890,N_381);
or U1182 (N_1182,N_319,N_982);
nand U1183 (N_1183,N_50,N_642);
and U1184 (N_1184,N_64,N_772);
nand U1185 (N_1185,N_437,N_755);
nand U1186 (N_1186,N_587,N_495);
nand U1187 (N_1187,N_368,N_284);
nand U1188 (N_1188,N_393,N_818);
nor U1189 (N_1189,N_535,N_247);
and U1190 (N_1190,N_656,N_259);
and U1191 (N_1191,N_500,N_126);
or U1192 (N_1192,N_981,N_770);
nor U1193 (N_1193,N_657,N_231);
nand U1194 (N_1194,N_31,N_953);
nand U1195 (N_1195,N_676,N_121);
xnor U1196 (N_1196,N_838,N_889);
nand U1197 (N_1197,N_295,N_584);
nor U1198 (N_1198,N_305,N_351);
or U1199 (N_1199,N_564,N_113);
nand U1200 (N_1200,N_842,N_148);
or U1201 (N_1201,N_242,N_384);
nor U1202 (N_1202,N_746,N_673);
and U1203 (N_1203,N_734,N_900);
nand U1204 (N_1204,N_827,N_10);
xnor U1205 (N_1205,N_721,N_977);
xor U1206 (N_1206,N_754,N_230);
nand U1207 (N_1207,N_750,N_794);
nor U1208 (N_1208,N_862,N_340);
and U1209 (N_1209,N_532,N_545);
nor U1210 (N_1210,N_139,N_405);
nand U1211 (N_1211,N_588,N_198);
nand U1212 (N_1212,N_94,N_422);
and U1213 (N_1213,N_48,N_942);
or U1214 (N_1214,N_706,N_660);
and U1215 (N_1215,N_107,N_201);
or U1216 (N_1216,N_51,N_753);
nand U1217 (N_1217,N_603,N_802);
nor U1218 (N_1218,N_567,N_666);
and U1219 (N_1219,N_30,N_310);
and U1220 (N_1220,N_66,N_116);
and U1221 (N_1221,N_496,N_776);
and U1222 (N_1222,N_406,N_927);
or U1223 (N_1223,N_687,N_225);
or U1224 (N_1224,N_168,N_926);
nor U1225 (N_1225,N_768,N_836);
xor U1226 (N_1226,N_26,N_715);
and U1227 (N_1227,N_270,N_965);
and U1228 (N_1228,N_739,N_655);
and U1229 (N_1229,N_175,N_317);
nor U1230 (N_1230,N_784,N_868);
or U1231 (N_1231,N_955,N_336);
or U1232 (N_1232,N_19,N_921);
nand U1233 (N_1233,N_366,N_762);
nand U1234 (N_1234,N_421,N_29);
nand U1235 (N_1235,N_434,N_967);
nor U1236 (N_1236,N_418,N_34);
nor U1237 (N_1237,N_966,N_487);
or U1238 (N_1238,N_459,N_749);
xnor U1239 (N_1239,N_763,N_428);
or U1240 (N_1240,N_277,N_617);
nand U1241 (N_1241,N_971,N_598);
xor U1242 (N_1242,N_313,N_515);
nor U1243 (N_1243,N_863,N_28);
nor U1244 (N_1244,N_169,N_394);
nand U1245 (N_1245,N_77,N_433);
nor U1246 (N_1246,N_129,N_47);
or U1247 (N_1247,N_929,N_933);
nand U1248 (N_1248,N_525,N_283);
nand U1249 (N_1249,N_42,N_438);
or U1250 (N_1250,N_343,N_40);
and U1251 (N_1251,N_712,N_36);
and U1252 (N_1252,N_548,N_895);
xnor U1253 (N_1253,N_689,N_724);
xor U1254 (N_1254,N_947,N_363);
xnor U1255 (N_1255,N_92,N_677);
nand U1256 (N_1256,N_973,N_210);
nand U1257 (N_1257,N_987,N_296);
nor U1258 (N_1258,N_455,N_624);
or U1259 (N_1259,N_360,N_614);
nand U1260 (N_1260,N_999,N_653);
nor U1261 (N_1261,N_84,N_669);
or U1262 (N_1262,N_114,N_575);
and U1263 (N_1263,N_344,N_460);
and U1264 (N_1264,N_465,N_814);
xor U1265 (N_1265,N_480,N_391);
and U1266 (N_1266,N_958,N_980);
and U1267 (N_1267,N_67,N_760);
and U1268 (N_1268,N_200,N_160);
nand U1269 (N_1269,N_158,N_481);
and U1270 (N_1270,N_425,N_479);
xnor U1271 (N_1271,N_606,N_408);
nor U1272 (N_1272,N_427,N_86);
or U1273 (N_1273,N_291,N_220);
and U1274 (N_1274,N_581,N_127);
or U1275 (N_1275,N_641,N_507);
nor U1276 (N_1276,N_87,N_132);
and U1277 (N_1277,N_223,N_219);
nor U1278 (N_1278,N_843,N_574);
nor U1279 (N_1279,N_675,N_380);
nand U1280 (N_1280,N_453,N_309);
and U1281 (N_1281,N_871,N_705);
or U1282 (N_1282,N_140,N_714);
or U1283 (N_1283,N_104,N_63);
nor U1284 (N_1284,N_150,N_992);
and U1285 (N_1285,N_822,N_442);
or U1286 (N_1286,N_178,N_537);
and U1287 (N_1287,N_449,N_934);
nor U1288 (N_1288,N_781,N_484);
xnor U1289 (N_1289,N_806,N_984);
nor U1290 (N_1290,N_300,N_356);
nor U1291 (N_1291,N_837,N_638);
and U1292 (N_1292,N_769,N_143);
nor U1293 (N_1293,N_265,N_969);
nand U1294 (N_1294,N_576,N_742);
nor U1295 (N_1295,N_745,N_996);
and U1296 (N_1296,N_79,N_563);
and U1297 (N_1297,N_252,N_103);
nor U1298 (N_1298,N_352,N_39);
xnor U1299 (N_1299,N_771,N_534);
nor U1300 (N_1300,N_511,N_93);
nand U1301 (N_1301,N_21,N_385);
nor U1302 (N_1302,N_685,N_633);
or U1303 (N_1303,N_726,N_573);
nor U1304 (N_1304,N_748,N_610);
or U1305 (N_1305,N_565,N_915);
nor U1306 (N_1306,N_22,N_329);
nand U1307 (N_1307,N_370,N_943);
and U1308 (N_1308,N_680,N_561);
nor U1309 (N_1309,N_602,N_956);
nor U1310 (N_1310,N_362,N_398);
nor U1311 (N_1311,N_3,N_334);
and U1312 (N_1312,N_124,N_928);
nand U1313 (N_1313,N_190,N_528);
nand U1314 (N_1314,N_181,N_73);
nor U1315 (N_1315,N_268,N_556);
or U1316 (N_1316,N_56,N_4);
nor U1317 (N_1317,N_426,N_823);
nand U1318 (N_1318,N_585,N_559);
or U1319 (N_1319,N_489,N_722);
nor U1320 (N_1320,N_851,N_626);
nor U1321 (N_1321,N_747,N_163);
nor U1322 (N_1322,N_607,N_176);
nor U1323 (N_1323,N_725,N_239);
nand U1324 (N_1324,N_684,N_506);
xnor U1325 (N_1325,N_604,N_492);
and U1326 (N_1326,N_810,N_711);
and U1327 (N_1327,N_141,N_120);
and U1328 (N_1328,N_885,N_901);
and U1329 (N_1329,N_720,N_860);
or U1330 (N_1330,N_622,N_796);
nor U1331 (N_1331,N_730,N_964);
and U1332 (N_1332,N_907,N_186);
and U1333 (N_1333,N_583,N_474);
nor U1334 (N_1334,N_832,N_388);
nor U1335 (N_1335,N_875,N_667);
or U1336 (N_1336,N_946,N_555);
or U1337 (N_1337,N_321,N_57);
or U1338 (N_1338,N_505,N_855);
nand U1339 (N_1339,N_494,N_215);
nor U1340 (N_1340,N_558,N_302);
and U1341 (N_1341,N_299,N_615);
and U1342 (N_1342,N_560,N_361);
or U1343 (N_1343,N_919,N_191);
nand U1344 (N_1344,N_224,N_547);
xnor U1345 (N_1345,N_944,N_708);
nand U1346 (N_1346,N_801,N_664);
or U1347 (N_1347,N_161,N_5);
or U1348 (N_1348,N_940,N_882);
xor U1349 (N_1349,N_605,N_209);
nor U1350 (N_1350,N_382,N_812);
and U1351 (N_1351,N_78,N_137);
or U1352 (N_1352,N_149,N_13);
and U1353 (N_1353,N_100,N_931);
or U1354 (N_1354,N_1,N_904);
and U1355 (N_1355,N_696,N_693);
or U1356 (N_1356,N_568,N_935);
nand U1357 (N_1357,N_960,N_529);
xor U1358 (N_1358,N_184,N_339);
nor U1359 (N_1359,N_878,N_436);
nor U1360 (N_1360,N_637,N_609);
and U1361 (N_1361,N_415,N_472);
xor U1362 (N_1362,N_468,N_948);
nor U1363 (N_1363,N_526,N_577);
nor U1364 (N_1364,N_451,N_144);
or U1365 (N_1365,N_627,N_792);
nor U1366 (N_1366,N_513,N_349);
nand U1367 (N_1367,N_281,N_873);
nand U1368 (N_1368,N_682,N_650);
or U1369 (N_1369,N_758,N_404);
nand U1370 (N_1370,N_729,N_170);
or U1371 (N_1371,N_738,N_323);
nand U1372 (N_1372,N_401,N_520);
and U1373 (N_1373,N_517,N_304);
nor U1374 (N_1374,N_854,N_635);
nand U1375 (N_1375,N_253,N_403);
nand U1376 (N_1376,N_596,N_630);
nor U1377 (N_1377,N_409,N_154);
xnor U1378 (N_1378,N_757,N_306);
or U1379 (N_1379,N_90,N_961);
and U1380 (N_1380,N_0,N_541);
or U1381 (N_1381,N_597,N_458);
nand U1382 (N_1382,N_694,N_916);
and U1383 (N_1383,N_46,N_658);
nor U1384 (N_1384,N_595,N_983);
xor U1385 (N_1385,N_25,N_389);
xnor U1386 (N_1386,N_75,N_690);
nand U1387 (N_1387,N_798,N_881);
nor U1388 (N_1388,N_330,N_866);
or U1389 (N_1389,N_12,N_824);
nor U1390 (N_1390,N_280,N_497);
or U1391 (N_1391,N_499,N_350);
and U1392 (N_1392,N_979,N_957);
and U1393 (N_1393,N_2,N_569);
nand U1394 (N_1394,N_737,N_371);
and U1395 (N_1395,N_692,N_145);
and U1396 (N_1396,N_723,N_600);
nand U1397 (N_1397,N_241,N_290);
nor U1398 (N_1398,N_897,N_539);
or U1399 (N_1399,N_783,N_212);
xnor U1400 (N_1400,N_72,N_8);
and U1401 (N_1401,N_249,N_365);
and U1402 (N_1402,N_668,N_795);
xnor U1403 (N_1403,N_743,N_203);
nand U1404 (N_1404,N_294,N_512);
nand U1405 (N_1405,N_153,N_331);
nand U1406 (N_1406,N_328,N_579);
or U1407 (N_1407,N_417,N_697);
nand U1408 (N_1408,N_138,N_182);
or U1409 (N_1409,N_945,N_623);
nand U1410 (N_1410,N_105,N_359);
nor U1411 (N_1411,N_400,N_552);
and U1412 (N_1412,N_478,N_652);
and U1413 (N_1413,N_76,N_341);
and U1414 (N_1414,N_592,N_518);
nor U1415 (N_1415,N_631,N_448);
nor U1416 (N_1416,N_524,N_791);
and U1417 (N_1417,N_533,N_187);
or U1418 (N_1418,N_876,N_383);
and U1419 (N_1419,N_308,N_375);
nand U1420 (N_1420,N_671,N_557);
nand U1421 (N_1421,N_374,N_222);
nand U1422 (N_1422,N_102,N_69);
nand U1423 (N_1423,N_157,N_628);
and U1424 (N_1424,N_376,N_691);
xor U1425 (N_1425,N_110,N_207);
xnor U1426 (N_1426,N_491,N_59);
or U1427 (N_1427,N_562,N_227);
nor U1428 (N_1428,N_476,N_88);
nand U1429 (N_1429,N_118,N_621);
nor U1430 (N_1430,N_913,N_589);
xor U1431 (N_1431,N_619,N_727);
nand U1432 (N_1432,N_236,N_424);
nor U1433 (N_1433,N_466,N_420);
nor U1434 (N_1434,N_787,N_324);
nor U1435 (N_1435,N_258,N_864);
nand U1436 (N_1436,N_703,N_99);
and U1437 (N_1437,N_266,N_911);
or U1438 (N_1438,N_888,N_995);
nand U1439 (N_1439,N_192,N_962);
nand U1440 (N_1440,N_861,N_649);
nand U1441 (N_1441,N_821,N_122);
nand U1442 (N_1442,N_387,N_736);
or U1443 (N_1443,N_251,N_233);
nand U1444 (N_1444,N_44,N_71);
and U1445 (N_1445,N_354,N_473);
xnor U1446 (N_1446,N_9,N_256);
nand U1447 (N_1447,N_764,N_91);
and U1448 (N_1448,N_636,N_767);
nand U1449 (N_1449,N_189,N_246);
nand U1450 (N_1450,N_912,N_786);
nor U1451 (N_1451,N_440,N_33);
nor U1452 (N_1452,N_963,N_322);
xnor U1453 (N_1453,N_765,N_196);
and U1454 (N_1454,N_293,N_808);
xnor U1455 (N_1455,N_216,N_815);
xor U1456 (N_1456,N_503,N_865);
nor U1457 (N_1457,N_456,N_879);
and U1458 (N_1458,N_83,N_586);
nor U1459 (N_1459,N_766,N_778);
and U1460 (N_1460,N_857,N_282);
or U1461 (N_1461,N_20,N_395);
or U1462 (N_1462,N_498,N_117);
and U1463 (N_1463,N_546,N_327);
and U1464 (N_1464,N_590,N_204);
nor U1465 (N_1465,N_788,N_213);
nor U1466 (N_1466,N_549,N_519);
nand U1467 (N_1467,N_782,N_464);
or U1468 (N_1468,N_62,N_937);
and U1469 (N_1469,N_70,N_95);
and U1470 (N_1470,N_679,N_654);
and U1471 (N_1471,N_261,N_975);
nor U1472 (N_1472,N_797,N_716);
nor U1473 (N_1473,N_611,N_257);
nand U1474 (N_1474,N_429,N_672);
nand U1475 (N_1475,N_644,N_16);
nor U1476 (N_1476,N_997,N_338);
and U1477 (N_1477,N_123,N_816);
and U1478 (N_1478,N_301,N_235);
and U1479 (N_1479,N_629,N_156);
or U1480 (N_1480,N_98,N_501);
nand U1481 (N_1481,N_326,N_55);
nand U1482 (N_1482,N_774,N_37);
and U1483 (N_1483,N_645,N_578);
nor U1484 (N_1484,N_392,N_828);
nand U1485 (N_1485,N_386,N_920);
nand U1486 (N_1486,N_289,N_752);
or U1487 (N_1487,N_978,N_262);
nand U1488 (N_1488,N_700,N_244);
nor U1489 (N_1489,N_859,N_179);
xnor U1490 (N_1490,N_831,N_989);
and U1491 (N_1491,N_410,N_735);
xnor U1492 (N_1492,N_172,N_841);
or U1493 (N_1493,N_591,N_819);
nand U1494 (N_1494,N_950,N_183);
nor U1495 (N_1495,N_850,N_835);
and U1496 (N_1496,N_58,N_910);
nand U1497 (N_1497,N_260,N_377);
nor U1498 (N_1498,N_41,N_431);
nand U1499 (N_1499,N_665,N_906);
nand U1500 (N_1500,N_480,N_801);
or U1501 (N_1501,N_222,N_927);
xor U1502 (N_1502,N_618,N_225);
and U1503 (N_1503,N_720,N_801);
and U1504 (N_1504,N_398,N_168);
and U1505 (N_1505,N_596,N_821);
nor U1506 (N_1506,N_565,N_108);
or U1507 (N_1507,N_370,N_812);
or U1508 (N_1508,N_366,N_382);
and U1509 (N_1509,N_131,N_575);
or U1510 (N_1510,N_210,N_83);
nor U1511 (N_1511,N_468,N_690);
nand U1512 (N_1512,N_454,N_902);
or U1513 (N_1513,N_34,N_573);
and U1514 (N_1514,N_466,N_110);
and U1515 (N_1515,N_598,N_260);
and U1516 (N_1516,N_676,N_467);
xor U1517 (N_1517,N_851,N_779);
or U1518 (N_1518,N_105,N_292);
and U1519 (N_1519,N_285,N_733);
nand U1520 (N_1520,N_342,N_769);
and U1521 (N_1521,N_64,N_203);
nand U1522 (N_1522,N_950,N_427);
nand U1523 (N_1523,N_595,N_760);
and U1524 (N_1524,N_785,N_910);
or U1525 (N_1525,N_943,N_734);
and U1526 (N_1526,N_880,N_741);
or U1527 (N_1527,N_41,N_213);
or U1528 (N_1528,N_108,N_170);
and U1529 (N_1529,N_49,N_352);
nand U1530 (N_1530,N_641,N_679);
and U1531 (N_1531,N_904,N_560);
nor U1532 (N_1532,N_828,N_489);
nor U1533 (N_1533,N_851,N_143);
nand U1534 (N_1534,N_773,N_941);
and U1535 (N_1535,N_264,N_212);
and U1536 (N_1536,N_284,N_915);
nor U1537 (N_1537,N_272,N_955);
nand U1538 (N_1538,N_985,N_933);
nand U1539 (N_1539,N_30,N_953);
or U1540 (N_1540,N_769,N_362);
or U1541 (N_1541,N_654,N_985);
or U1542 (N_1542,N_627,N_993);
xnor U1543 (N_1543,N_14,N_312);
and U1544 (N_1544,N_807,N_611);
and U1545 (N_1545,N_680,N_72);
nor U1546 (N_1546,N_183,N_371);
nor U1547 (N_1547,N_278,N_987);
and U1548 (N_1548,N_702,N_620);
and U1549 (N_1549,N_674,N_880);
nor U1550 (N_1550,N_29,N_595);
and U1551 (N_1551,N_971,N_46);
and U1552 (N_1552,N_879,N_429);
nand U1553 (N_1553,N_80,N_460);
nor U1554 (N_1554,N_411,N_998);
nand U1555 (N_1555,N_928,N_984);
and U1556 (N_1556,N_118,N_447);
and U1557 (N_1557,N_602,N_609);
nor U1558 (N_1558,N_249,N_791);
nor U1559 (N_1559,N_998,N_247);
nor U1560 (N_1560,N_849,N_709);
and U1561 (N_1561,N_983,N_60);
nor U1562 (N_1562,N_948,N_530);
nor U1563 (N_1563,N_438,N_143);
xnor U1564 (N_1564,N_160,N_440);
or U1565 (N_1565,N_340,N_63);
nand U1566 (N_1566,N_564,N_415);
and U1567 (N_1567,N_564,N_301);
and U1568 (N_1568,N_821,N_51);
or U1569 (N_1569,N_36,N_399);
nor U1570 (N_1570,N_757,N_509);
nand U1571 (N_1571,N_255,N_120);
xor U1572 (N_1572,N_318,N_925);
nor U1573 (N_1573,N_104,N_131);
xor U1574 (N_1574,N_871,N_969);
or U1575 (N_1575,N_215,N_187);
xor U1576 (N_1576,N_729,N_297);
nor U1577 (N_1577,N_226,N_970);
or U1578 (N_1578,N_515,N_676);
nand U1579 (N_1579,N_510,N_601);
or U1580 (N_1580,N_279,N_656);
and U1581 (N_1581,N_334,N_278);
and U1582 (N_1582,N_48,N_343);
and U1583 (N_1583,N_757,N_384);
or U1584 (N_1584,N_401,N_565);
xnor U1585 (N_1585,N_441,N_937);
or U1586 (N_1586,N_562,N_710);
and U1587 (N_1587,N_540,N_979);
and U1588 (N_1588,N_23,N_150);
nand U1589 (N_1589,N_262,N_628);
and U1590 (N_1590,N_70,N_393);
nand U1591 (N_1591,N_966,N_787);
and U1592 (N_1592,N_758,N_308);
nand U1593 (N_1593,N_302,N_83);
nor U1594 (N_1594,N_20,N_15);
or U1595 (N_1595,N_197,N_657);
xor U1596 (N_1596,N_48,N_784);
nand U1597 (N_1597,N_212,N_106);
and U1598 (N_1598,N_190,N_362);
nor U1599 (N_1599,N_129,N_670);
nand U1600 (N_1600,N_216,N_546);
and U1601 (N_1601,N_629,N_931);
nand U1602 (N_1602,N_88,N_905);
xor U1603 (N_1603,N_659,N_944);
nor U1604 (N_1604,N_291,N_262);
xnor U1605 (N_1605,N_528,N_384);
xor U1606 (N_1606,N_616,N_805);
and U1607 (N_1607,N_650,N_329);
xnor U1608 (N_1608,N_653,N_382);
or U1609 (N_1609,N_429,N_533);
and U1610 (N_1610,N_888,N_615);
and U1611 (N_1611,N_256,N_866);
or U1612 (N_1612,N_245,N_493);
or U1613 (N_1613,N_458,N_106);
and U1614 (N_1614,N_879,N_110);
xnor U1615 (N_1615,N_34,N_610);
and U1616 (N_1616,N_850,N_874);
nand U1617 (N_1617,N_550,N_301);
or U1618 (N_1618,N_128,N_372);
and U1619 (N_1619,N_40,N_707);
xor U1620 (N_1620,N_924,N_215);
and U1621 (N_1621,N_535,N_420);
nor U1622 (N_1622,N_420,N_290);
nand U1623 (N_1623,N_459,N_624);
or U1624 (N_1624,N_234,N_734);
and U1625 (N_1625,N_626,N_301);
xor U1626 (N_1626,N_777,N_206);
or U1627 (N_1627,N_321,N_99);
xor U1628 (N_1628,N_761,N_309);
and U1629 (N_1629,N_867,N_873);
or U1630 (N_1630,N_508,N_80);
nand U1631 (N_1631,N_528,N_593);
or U1632 (N_1632,N_911,N_780);
or U1633 (N_1633,N_252,N_321);
nor U1634 (N_1634,N_63,N_750);
and U1635 (N_1635,N_722,N_966);
or U1636 (N_1636,N_285,N_317);
xnor U1637 (N_1637,N_206,N_576);
or U1638 (N_1638,N_207,N_580);
nor U1639 (N_1639,N_589,N_724);
and U1640 (N_1640,N_454,N_609);
nor U1641 (N_1641,N_105,N_12);
and U1642 (N_1642,N_744,N_459);
nand U1643 (N_1643,N_781,N_601);
or U1644 (N_1644,N_390,N_139);
or U1645 (N_1645,N_573,N_363);
nand U1646 (N_1646,N_420,N_760);
or U1647 (N_1647,N_641,N_78);
nor U1648 (N_1648,N_55,N_316);
and U1649 (N_1649,N_413,N_593);
or U1650 (N_1650,N_51,N_183);
or U1651 (N_1651,N_245,N_606);
nand U1652 (N_1652,N_512,N_485);
nand U1653 (N_1653,N_987,N_633);
and U1654 (N_1654,N_794,N_88);
and U1655 (N_1655,N_419,N_101);
and U1656 (N_1656,N_548,N_526);
and U1657 (N_1657,N_745,N_136);
xnor U1658 (N_1658,N_38,N_174);
nor U1659 (N_1659,N_39,N_356);
nor U1660 (N_1660,N_830,N_944);
and U1661 (N_1661,N_783,N_270);
or U1662 (N_1662,N_120,N_184);
or U1663 (N_1663,N_139,N_633);
nand U1664 (N_1664,N_354,N_874);
nor U1665 (N_1665,N_995,N_44);
nand U1666 (N_1666,N_672,N_149);
or U1667 (N_1667,N_13,N_717);
nand U1668 (N_1668,N_418,N_562);
and U1669 (N_1669,N_229,N_713);
and U1670 (N_1670,N_145,N_696);
nand U1671 (N_1671,N_564,N_920);
or U1672 (N_1672,N_600,N_663);
nand U1673 (N_1673,N_430,N_935);
and U1674 (N_1674,N_166,N_205);
nor U1675 (N_1675,N_560,N_819);
or U1676 (N_1676,N_136,N_187);
nor U1677 (N_1677,N_905,N_414);
or U1678 (N_1678,N_190,N_230);
or U1679 (N_1679,N_96,N_229);
nand U1680 (N_1680,N_286,N_168);
or U1681 (N_1681,N_348,N_997);
nand U1682 (N_1682,N_129,N_990);
or U1683 (N_1683,N_588,N_90);
and U1684 (N_1684,N_118,N_70);
nor U1685 (N_1685,N_757,N_618);
nor U1686 (N_1686,N_990,N_26);
nand U1687 (N_1687,N_193,N_83);
and U1688 (N_1688,N_457,N_605);
nand U1689 (N_1689,N_969,N_674);
or U1690 (N_1690,N_237,N_40);
and U1691 (N_1691,N_145,N_707);
and U1692 (N_1692,N_180,N_890);
xor U1693 (N_1693,N_828,N_79);
nand U1694 (N_1694,N_897,N_513);
nand U1695 (N_1695,N_637,N_621);
xnor U1696 (N_1696,N_821,N_331);
and U1697 (N_1697,N_495,N_868);
nor U1698 (N_1698,N_607,N_747);
or U1699 (N_1699,N_292,N_162);
nand U1700 (N_1700,N_107,N_401);
and U1701 (N_1701,N_878,N_363);
and U1702 (N_1702,N_252,N_971);
xor U1703 (N_1703,N_430,N_892);
nand U1704 (N_1704,N_396,N_165);
xnor U1705 (N_1705,N_929,N_962);
nor U1706 (N_1706,N_442,N_238);
nor U1707 (N_1707,N_371,N_102);
or U1708 (N_1708,N_395,N_89);
nand U1709 (N_1709,N_519,N_546);
or U1710 (N_1710,N_892,N_391);
nand U1711 (N_1711,N_603,N_107);
nand U1712 (N_1712,N_826,N_638);
and U1713 (N_1713,N_899,N_572);
nand U1714 (N_1714,N_168,N_527);
or U1715 (N_1715,N_315,N_761);
and U1716 (N_1716,N_972,N_329);
nor U1717 (N_1717,N_756,N_84);
and U1718 (N_1718,N_153,N_181);
or U1719 (N_1719,N_259,N_622);
or U1720 (N_1720,N_867,N_507);
nor U1721 (N_1721,N_255,N_616);
or U1722 (N_1722,N_881,N_323);
nor U1723 (N_1723,N_143,N_686);
nor U1724 (N_1724,N_655,N_875);
or U1725 (N_1725,N_67,N_991);
or U1726 (N_1726,N_433,N_359);
nor U1727 (N_1727,N_716,N_811);
nand U1728 (N_1728,N_912,N_858);
and U1729 (N_1729,N_317,N_714);
nand U1730 (N_1730,N_859,N_902);
and U1731 (N_1731,N_848,N_590);
nor U1732 (N_1732,N_417,N_908);
or U1733 (N_1733,N_9,N_757);
xnor U1734 (N_1734,N_164,N_433);
or U1735 (N_1735,N_309,N_949);
or U1736 (N_1736,N_461,N_745);
nor U1737 (N_1737,N_406,N_29);
or U1738 (N_1738,N_62,N_33);
nand U1739 (N_1739,N_808,N_314);
nor U1740 (N_1740,N_9,N_75);
nand U1741 (N_1741,N_824,N_723);
xor U1742 (N_1742,N_22,N_434);
and U1743 (N_1743,N_237,N_444);
nor U1744 (N_1744,N_189,N_243);
nor U1745 (N_1745,N_814,N_514);
or U1746 (N_1746,N_120,N_121);
nand U1747 (N_1747,N_306,N_157);
nor U1748 (N_1748,N_655,N_794);
and U1749 (N_1749,N_239,N_7);
or U1750 (N_1750,N_139,N_468);
xor U1751 (N_1751,N_755,N_412);
and U1752 (N_1752,N_186,N_847);
and U1753 (N_1753,N_287,N_693);
nand U1754 (N_1754,N_304,N_959);
and U1755 (N_1755,N_752,N_358);
and U1756 (N_1756,N_869,N_887);
or U1757 (N_1757,N_842,N_873);
nand U1758 (N_1758,N_270,N_126);
or U1759 (N_1759,N_524,N_464);
nor U1760 (N_1760,N_266,N_564);
xor U1761 (N_1761,N_661,N_145);
nor U1762 (N_1762,N_254,N_475);
nand U1763 (N_1763,N_112,N_784);
and U1764 (N_1764,N_666,N_571);
and U1765 (N_1765,N_491,N_519);
or U1766 (N_1766,N_363,N_563);
nand U1767 (N_1767,N_751,N_503);
nand U1768 (N_1768,N_799,N_99);
nand U1769 (N_1769,N_596,N_324);
nand U1770 (N_1770,N_394,N_968);
nor U1771 (N_1771,N_487,N_466);
and U1772 (N_1772,N_183,N_53);
nand U1773 (N_1773,N_344,N_847);
and U1774 (N_1774,N_410,N_575);
and U1775 (N_1775,N_252,N_71);
or U1776 (N_1776,N_845,N_317);
xor U1777 (N_1777,N_820,N_538);
or U1778 (N_1778,N_948,N_252);
or U1779 (N_1779,N_490,N_654);
or U1780 (N_1780,N_313,N_95);
nand U1781 (N_1781,N_677,N_660);
nor U1782 (N_1782,N_8,N_791);
and U1783 (N_1783,N_175,N_822);
nand U1784 (N_1784,N_701,N_574);
nor U1785 (N_1785,N_533,N_749);
and U1786 (N_1786,N_664,N_553);
xnor U1787 (N_1787,N_477,N_166);
nand U1788 (N_1788,N_523,N_968);
nand U1789 (N_1789,N_176,N_251);
nand U1790 (N_1790,N_793,N_391);
and U1791 (N_1791,N_226,N_746);
nand U1792 (N_1792,N_839,N_913);
nor U1793 (N_1793,N_610,N_816);
or U1794 (N_1794,N_964,N_542);
nand U1795 (N_1795,N_154,N_841);
nor U1796 (N_1796,N_797,N_437);
and U1797 (N_1797,N_815,N_412);
or U1798 (N_1798,N_801,N_786);
nor U1799 (N_1799,N_507,N_590);
xor U1800 (N_1800,N_6,N_881);
and U1801 (N_1801,N_63,N_699);
nand U1802 (N_1802,N_744,N_561);
nand U1803 (N_1803,N_576,N_355);
and U1804 (N_1804,N_651,N_94);
xnor U1805 (N_1805,N_566,N_44);
and U1806 (N_1806,N_804,N_480);
and U1807 (N_1807,N_424,N_674);
nor U1808 (N_1808,N_186,N_928);
xnor U1809 (N_1809,N_918,N_110);
nor U1810 (N_1810,N_791,N_927);
nor U1811 (N_1811,N_685,N_774);
nand U1812 (N_1812,N_138,N_822);
nor U1813 (N_1813,N_545,N_846);
and U1814 (N_1814,N_550,N_688);
nor U1815 (N_1815,N_855,N_674);
and U1816 (N_1816,N_264,N_311);
or U1817 (N_1817,N_217,N_45);
nor U1818 (N_1818,N_757,N_469);
nor U1819 (N_1819,N_868,N_754);
and U1820 (N_1820,N_316,N_89);
xor U1821 (N_1821,N_528,N_189);
nor U1822 (N_1822,N_977,N_912);
nor U1823 (N_1823,N_912,N_469);
and U1824 (N_1824,N_342,N_727);
nand U1825 (N_1825,N_577,N_200);
and U1826 (N_1826,N_163,N_254);
nor U1827 (N_1827,N_359,N_721);
nor U1828 (N_1828,N_125,N_915);
and U1829 (N_1829,N_600,N_399);
and U1830 (N_1830,N_180,N_217);
or U1831 (N_1831,N_283,N_468);
nor U1832 (N_1832,N_406,N_443);
or U1833 (N_1833,N_736,N_245);
nor U1834 (N_1834,N_130,N_330);
nor U1835 (N_1835,N_671,N_502);
nor U1836 (N_1836,N_928,N_107);
xnor U1837 (N_1837,N_843,N_77);
or U1838 (N_1838,N_918,N_777);
or U1839 (N_1839,N_647,N_302);
nor U1840 (N_1840,N_636,N_727);
nand U1841 (N_1841,N_212,N_564);
and U1842 (N_1842,N_515,N_411);
nand U1843 (N_1843,N_553,N_667);
nand U1844 (N_1844,N_320,N_977);
nor U1845 (N_1845,N_649,N_503);
or U1846 (N_1846,N_354,N_635);
nand U1847 (N_1847,N_854,N_279);
nand U1848 (N_1848,N_579,N_296);
or U1849 (N_1849,N_945,N_7);
or U1850 (N_1850,N_130,N_42);
nand U1851 (N_1851,N_968,N_166);
nand U1852 (N_1852,N_707,N_828);
or U1853 (N_1853,N_461,N_783);
xor U1854 (N_1854,N_337,N_972);
nand U1855 (N_1855,N_32,N_29);
nor U1856 (N_1856,N_605,N_596);
or U1857 (N_1857,N_869,N_659);
nand U1858 (N_1858,N_186,N_434);
nand U1859 (N_1859,N_519,N_482);
or U1860 (N_1860,N_875,N_207);
or U1861 (N_1861,N_485,N_450);
nand U1862 (N_1862,N_839,N_873);
nor U1863 (N_1863,N_213,N_628);
and U1864 (N_1864,N_741,N_42);
and U1865 (N_1865,N_594,N_95);
nand U1866 (N_1866,N_120,N_10);
and U1867 (N_1867,N_757,N_299);
and U1868 (N_1868,N_436,N_205);
nor U1869 (N_1869,N_386,N_149);
nand U1870 (N_1870,N_64,N_864);
nor U1871 (N_1871,N_682,N_476);
nand U1872 (N_1872,N_909,N_88);
and U1873 (N_1873,N_627,N_97);
nor U1874 (N_1874,N_306,N_779);
nand U1875 (N_1875,N_970,N_374);
nor U1876 (N_1876,N_757,N_480);
nor U1877 (N_1877,N_325,N_701);
or U1878 (N_1878,N_990,N_938);
nor U1879 (N_1879,N_312,N_556);
or U1880 (N_1880,N_682,N_314);
xor U1881 (N_1881,N_794,N_599);
or U1882 (N_1882,N_654,N_788);
or U1883 (N_1883,N_182,N_757);
nand U1884 (N_1884,N_373,N_246);
and U1885 (N_1885,N_819,N_988);
nand U1886 (N_1886,N_696,N_220);
xnor U1887 (N_1887,N_120,N_520);
or U1888 (N_1888,N_335,N_228);
xnor U1889 (N_1889,N_459,N_779);
nand U1890 (N_1890,N_715,N_180);
and U1891 (N_1891,N_882,N_588);
or U1892 (N_1892,N_263,N_249);
nand U1893 (N_1893,N_878,N_73);
or U1894 (N_1894,N_958,N_984);
or U1895 (N_1895,N_500,N_932);
nor U1896 (N_1896,N_314,N_456);
nor U1897 (N_1897,N_541,N_484);
nand U1898 (N_1898,N_331,N_695);
nor U1899 (N_1899,N_153,N_414);
and U1900 (N_1900,N_566,N_599);
nand U1901 (N_1901,N_443,N_449);
and U1902 (N_1902,N_151,N_777);
nand U1903 (N_1903,N_886,N_823);
or U1904 (N_1904,N_685,N_471);
nand U1905 (N_1905,N_84,N_419);
nand U1906 (N_1906,N_885,N_309);
nand U1907 (N_1907,N_901,N_181);
xnor U1908 (N_1908,N_59,N_77);
nand U1909 (N_1909,N_360,N_819);
nand U1910 (N_1910,N_226,N_172);
nor U1911 (N_1911,N_772,N_960);
nand U1912 (N_1912,N_898,N_294);
xnor U1913 (N_1913,N_891,N_38);
or U1914 (N_1914,N_65,N_837);
and U1915 (N_1915,N_439,N_112);
nand U1916 (N_1916,N_988,N_993);
or U1917 (N_1917,N_202,N_347);
nor U1918 (N_1918,N_963,N_273);
nor U1919 (N_1919,N_428,N_890);
nor U1920 (N_1920,N_238,N_712);
or U1921 (N_1921,N_490,N_335);
nand U1922 (N_1922,N_684,N_750);
or U1923 (N_1923,N_54,N_20);
xor U1924 (N_1924,N_460,N_331);
nand U1925 (N_1925,N_786,N_307);
nor U1926 (N_1926,N_282,N_718);
nor U1927 (N_1927,N_459,N_505);
nand U1928 (N_1928,N_176,N_299);
or U1929 (N_1929,N_526,N_259);
or U1930 (N_1930,N_149,N_562);
nand U1931 (N_1931,N_785,N_341);
nor U1932 (N_1932,N_467,N_964);
or U1933 (N_1933,N_44,N_275);
or U1934 (N_1934,N_384,N_490);
or U1935 (N_1935,N_862,N_554);
nand U1936 (N_1936,N_416,N_603);
or U1937 (N_1937,N_65,N_347);
and U1938 (N_1938,N_619,N_267);
or U1939 (N_1939,N_238,N_607);
nand U1940 (N_1940,N_759,N_753);
nand U1941 (N_1941,N_474,N_715);
and U1942 (N_1942,N_938,N_609);
nor U1943 (N_1943,N_695,N_586);
nor U1944 (N_1944,N_832,N_282);
nor U1945 (N_1945,N_203,N_121);
and U1946 (N_1946,N_352,N_24);
and U1947 (N_1947,N_111,N_714);
nor U1948 (N_1948,N_177,N_891);
or U1949 (N_1949,N_196,N_969);
or U1950 (N_1950,N_453,N_931);
nand U1951 (N_1951,N_248,N_390);
and U1952 (N_1952,N_100,N_333);
xor U1953 (N_1953,N_672,N_454);
and U1954 (N_1954,N_96,N_550);
xor U1955 (N_1955,N_906,N_163);
nor U1956 (N_1956,N_378,N_78);
nor U1957 (N_1957,N_883,N_93);
or U1958 (N_1958,N_244,N_340);
or U1959 (N_1959,N_720,N_444);
nand U1960 (N_1960,N_321,N_866);
and U1961 (N_1961,N_811,N_146);
or U1962 (N_1962,N_42,N_896);
and U1963 (N_1963,N_415,N_773);
or U1964 (N_1964,N_705,N_765);
nand U1965 (N_1965,N_920,N_218);
and U1966 (N_1966,N_178,N_503);
nor U1967 (N_1967,N_865,N_385);
nor U1968 (N_1968,N_774,N_392);
nand U1969 (N_1969,N_426,N_380);
nand U1970 (N_1970,N_553,N_290);
nand U1971 (N_1971,N_350,N_345);
nor U1972 (N_1972,N_212,N_463);
nor U1973 (N_1973,N_392,N_410);
nand U1974 (N_1974,N_371,N_187);
or U1975 (N_1975,N_414,N_430);
or U1976 (N_1976,N_937,N_210);
and U1977 (N_1977,N_379,N_905);
or U1978 (N_1978,N_579,N_956);
nor U1979 (N_1979,N_399,N_193);
or U1980 (N_1980,N_392,N_326);
or U1981 (N_1981,N_288,N_731);
nand U1982 (N_1982,N_80,N_283);
nand U1983 (N_1983,N_379,N_136);
nor U1984 (N_1984,N_821,N_446);
and U1985 (N_1985,N_635,N_558);
and U1986 (N_1986,N_319,N_99);
nand U1987 (N_1987,N_18,N_176);
nor U1988 (N_1988,N_509,N_129);
and U1989 (N_1989,N_809,N_845);
and U1990 (N_1990,N_520,N_857);
or U1991 (N_1991,N_45,N_165);
xor U1992 (N_1992,N_102,N_450);
or U1993 (N_1993,N_261,N_5);
and U1994 (N_1994,N_13,N_170);
and U1995 (N_1995,N_145,N_591);
and U1996 (N_1996,N_570,N_66);
xnor U1997 (N_1997,N_146,N_619);
nand U1998 (N_1998,N_988,N_232);
nor U1999 (N_1999,N_91,N_204);
and U2000 (N_2000,N_1337,N_1748);
nand U2001 (N_2001,N_1688,N_1473);
or U2002 (N_2002,N_1593,N_1757);
and U2003 (N_2003,N_1938,N_1316);
and U2004 (N_2004,N_1936,N_1461);
xor U2005 (N_2005,N_1297,N_1282);
nand U2006 (N_2006,N_1385,N_1235);
xnor U2007 (N_2007,N_1851,N_1369);
nand U2008 (N_2008,N_1345,N_1110);
nand U2009 (N_2009,N_1958,N_1326);
or U2010 (N_2010,N_1614,N_1608);
nand U2011 (N_2011,N_1454,N_1310);
and U2012 (N_2012,N_1531,N_1479);
xnor U2013 (N_2013,N_1018,N_1581);
nand U2014 (N_2014,N_1277,N_1508);
or U2015 (N_2015,N_1700,N_1962);
nor U2016 (N_2016,N_1585,N_1642);
nor U2017 (N_2017,N_1666,N_1114);
nor U2018 (N_2018,N_1848,N_1170);
nand U2019 (N_2019,N_1205,N_1653);
and U2020 (N_2020,N_1550,N_1339);
xnor U2021 (N_2021,N_1094,N_1861);
or U2022 (N_2022,N_1291,N_1472);
and U2023 (N_2023,N_1024,N_1828);
or U2024 (N_2024,N_1306,N_1395);
xor U2025 (N_2025,N_1836,N_1724);
nand U2026 (N_2026,N_1145,N_1838);
xnor U2027 (N_2027,N_1774,N_1554);
or U2028 (N_2028,N_1992,N_1049);
nor U2029 (N_2029,N_1712,N_1380);
nand U2030 (N_2030,N_1603,N_1545);
nand U2031 (N_2031,N_1892,N_1398);
or U2032 (N_2032,N_1661,N_1986);
nand U2033 (N_2033,N_1429,N_1328);
and U2034 (N_2034,N_1191,N_1257);
nand U2035 (N_2035,N_1839,N_1678);
nand U2036 (N_2036,N_1286,N_1227);
nand U2037 (N_2037,N_1807,N_1621);
xor U2038 (N_2038,N_1532,N_1402);
and U2039 (N_2039,N_1223,N_1054);
and U2040 (N_2040,N_1070,N_1565);
nor U2041 (N_2041,N_1616,N_1033);
and U2042 (N_2042,N_1761,N_1327);
nand U2043 (N_2043,N_1965,N_1733);
nor U2044 (N_2044,N_1460,N_1100);
and U2045 (N_2045,N_1721,N_1207);
and U2046 (N_2046,N_1014,N_1204);
nor U2047 (N_2047,N_1843,N_1841);
nor U2048 (N_2048,N_1809,N_1190);
nand U2049 (N_2049,N_1635,N_1879);
xor U2050 (N_2050,N_1760,N_1737);
nor U2051 (N_2051,N_1726,N_1899);
nor U2052 (N_2052,N_1939,N_1477);
or U2053 (N_2053,N_1978,N_1789);
nor U2054 (N_2054,N_1015,N_1209);
and U2055 (N_2055,N_1115,N_1269);
nor U2056 (N_2056,N_1423,N_1085);
nand U2057 (N_2057,N_1800,N_1592);
and U2058 (N_2058,N_1742,N_1975);
and U2059 (N_2059,N_1266,N_1336);
and U2060 (N_2060,N_1347,N_1571);
or U2061 (N_2061,N_1799,N_1776);
nand U2062 (N_2062,N_1989,N_1136);
nor U2063 (N_2063,N_1199,N_1882);
xnor U2064 (N_2064,N_1053,N_1759);
or U2065 (N_2065,N_1138,N_1216);
or U2066 (N_2066,N_1278,N_1427);
nor U2067 (N_2067,N_1459,N_1817);
nand U2068 (N_2068,N_1364,N_1262);
or U2069 (N_2069,N_1078,N_1343);
nor U2070 (N_2070,N_1378,N_1980);
or U2071 (N_2071,N_1436,N_1677);
or U2072 (N_2072,N_1811,N_1476);
nor U2073 (N_2073,N_1360,N_1627);
or U2074 (N_2074,N_1357,N_1599);
nand U2075 (N_2075,N_1243,N_1954);
and U2076 (N_2076,N_1417,N_1027);
or U2077 (N_2077,N_1346,N_1862);
xnor U2078 (N_2078,N_1596,N_1432);
or U2079 (N_2079,N_1098,N_1539);
nor U2080 (N_2080,N_1521,N_1864);
nor U2081 (N_2081,N_1034,N_1180);
nand U2082 (N_2082,N_1239,N_1323);
and U2083 (N_2083,N_1203,N_1820);
nand U2084 (N_2084,N_1998,N_1388);
or U2085 (N_2085,N_1729,N_1470);
nand U2086 (N_2086,N_1615,N_1969);
and U2087 (N_2087,N_1896,N_1823);
nor U2088 (N_2088,N_1156,N_1768);
or U2089 (N_2089,N_1943,N_1217);
nand U2090 (N_2090,N_1179,N_1650);
xnor U2091 (N_2091,N_1743,N_1013);
nand U2092 (N_2092,N_1077,N_1687);
or U2093 (N_2093,N_1988,N_1993);
nand U2094 (N_2094,N_1431,N_1569);
and U2095 (N_2095,N_1496,N_1734);
nor U2096 (N_2096,N_1693,N_1405);
nor U2097 (N_2097,N_1654,N_1104);
xnor U2098 (N_2098,N_1246,N_1029);
nand U2099 (N_2099,N_1884,N_1031);
and U2100 (N_2100,N_1491,N_1238);
nand U2101 (N_2101,N_1690,N_1983);
or U2102 (N_2102,N_1547,N_1544);
and U2103 (N_2103,N_1135,N_1872);
and U2104 (N_2104,N_1684,N_1072);
nand U2105 (N_2105,N_1795,N_1131);
nor U2106 (N_2106,N_1281,N_1708);
and U2107 (N_2107,N_1079,N_1801);
nor U2108 (N_2108,N_1723,N_1927);
xnor U2109 (N_2109,N_1169,N_1215);
or U2110 (N_2110,N_1572,N_1679);
and U2111 (N_2111,N_1959,N_1683);
nand U2112 (N_2112,N_1334,N_1852);
or U2113 (N_2113,N_1375,N_1964);
nand U2114 (N_2114,N_1561,N_1229);
or U2115 (N_2115,N_1793,N_1740);
nand U2116 (N_2116,N_1010,N_1917);
nor U2117 (N_2117,N_1154,N_1289);
nor U2118 (N_2118,N_1271,N_1102);
or U2119 (N_2119,N_1805,N_1058);
and U2120 (N_2120,N_1143,N_1503);
and U2121 (N_2121,N_1052,N_1391);
or U2122 (N_2122,N_1438,N_1556);
nand U2123 (N_2123,N_1363,N_1549);
and U2124 (N_2124,N_1171,N_1664);
xnor U2125 (N_2125,N_1329,N_1250);
and U2126 (N_2126,N_1971,N_1351);
nand U2127 (N_2127,N_1876,N_1855);
and U2128 (N_2128,N_1731,N_1221);
nand U2129 (N_2129,N_1292,N_1122);
and U2130 (N_2130,N_1060,N_1562);
nor U2131 (N_2131,N_1868,N_1057);
or U2132 (N_2132,N_1344,N_1056);
nor U2133 (N_2133,N_1301,N_1397);
or U2134 (N_2134,N_1232,N_1225);
xnor U2135 (N_2135,N_1727,N_1617);
nor U2136 (N_2136,N_1484,N_1538);
or U2137 (N_2137,N_1368,N_1824);
and U2138 (N_2138,N_1003,N_1008);
nand U2139 (N_2139,N_1691,N_1469);
or U2140 (N_2140,N_1042,N_1674);
nor U2141 (N_2141,N_1919,N_1973);
nand U2142 (N_2142,N_1059,N_1177);
and U2143 (N_2143,N_1092,N_1632);
nor U2144 (N_2144,N_1312,N_1744);
nand U2145 (N_2145,N_1443,N_1118);
nor U2146 (N_2146,N_1140,N_1730);
nand U2147 (N_2147,N_1619,N_1313);
and U2148 (N_2148,N_1854,N_1451);
or U2149 (N_2149,N_1831,N_1778);
nand U2150 (N_2150,N_1821,N_1739);
nor U2151 (N_2151,N_1133,N_1447);
or U2152 (N_2152,N_1910,N_1275);
nor U2153 (N_2153,N_1797,N_1338);
or U2154 (N_2154,N_1948,N_1520);
nor U2155 (N_2155,N_1048,N_1090);
and U2156 (N_2156,N_1967,N_1210);
nand U2157 (N_2157,N_1780,N_1694);
xor U2158 (N_2158,N_1643,N_1717);
or U2159 (N_2159,N_1941,N_1612);
or U2160 (N_2160,N_1833,N_1088);
nor U2161 (N_2161,N_1409,N_1152);
or U2162 (N_2162,N_1139,N_1883);
nand U2163 (N_2163,N_1907,N_1189);
nand U2164 (N_2164,N_1294,N_1400);
nand U2165 (N_2165,N_1132,N_1584);
nor U2166 (N_2166,N_1440,N_1428);
xor U2167 (N_2167,N_1555,N_1891);
and U2168 (N_2168,N_1652,N_1952);
or U2169 (N_2169,N_1366,N_1582);
and U2170 (N_2170,N_1228,N_1002);
nand U2171 (N_2171,N_1183,N_1559);
and U2172 (N_2172,N_1526,N_1722);
nand U2173 (N_2173,N_1951,N_1367);
and U2174 (N_2174,N_1163,N_1591);
or U2175 (N_2175,N_1548,N_1990);
nand U2176 (N_2176,N_1787,N_1030);
nor U2177 (N_2177,N_1038,N_1198);
nand U2178 (N_2178,N_1074,N_1573);
nor U2179 (N_2179,N_1705,N_1942);
nand U2180 (N_2180,N_1084,N_1706);
nand U2181 (N_2181,N_1127,N_1745);
or U2182 (N_2182,N_1396,N_1121);
nor U2183 (N_2183,N_1506,N_1937);
and U2184 (N_2184,N_1251,N_1898);
nor U2185 (N_2185,N_1285,N_1877);
and U2186 (N_2186,N_1697,N_1494);
or U2187 (N_2187,N_1445,N_1644);
nand U2188 (N_2188,N_1258,N_1835);
or U2189 (N_2189,N_1812,N_1467);
or U2190 (N_2190,N_1510,N_1887);
or U2191 (N_2191,N_1062,N_1816);
nor U2192 (N_2192,N_1782,N_1829);
nor U2193 (N_2193,N_1912,N_1097);
and U2194 (N_2194,N_1302,N_1441);
xor U2195 (N_2195,N_1178,N_1982);
nand U2196 (N_2196,N_1618,N_1752);
nor U2197 (N_2197,N_1840,N_1055);
nand U2198 (N_2198,N_1350,N_1685);
nand U2199 (N_2199,N_1325,N_1908);
or U2200 (N_2200,N_1558,N_1792);
nor U2201 (N_2201,N_1832,N_1750);
nand U2202 (N_2202,N_1767,N_1117);
nand U2203 (N_2203,N_1361,N_1699);
or U2204 (N_2204,N_1028,N_1321);
or U2205 (N_2205,N_1420,N_1991);
and U2206 (N_2206,N_1613,N_1270);
nand U2207 (N_2207,N_1267,N_1419);
or U2208 (N_2208,N_1846,N_1356);
and U2209 (N_2209,N_1575,N_1012);
and U2210 (N_2210,N_1148,N_1176);
nor U2211 (N_2211,N_1924,N_1537);
nor U2212 (N_2212,N_1576,N_1977);
nand U2213 (N_2213,N_1474,N_1637);
and U2214 (N_2214,N_1631,N_1211);
nand U2215 (N_2215,N_1994,N_1017);
or U2216 (N_2216,N_1482,N_1174);
nor U2217 (N_2217,N_1044,N_1925);
nand U2218 (N_2218,N_1681,N_1736);
or U2219 (N_2219,N_1112,N_1598);
xor U2220 (N_2220,N_1111,N_1830);
and U2221 (N_2221,N_1091,N_1206);
and U2222 (N_2222,N_1248,N_1659);
nand U2223 (N_2223,N_1252,N_1224);
or U2224 (N_2224,N_1777,N_1629);
and U2225 (N_2225,N_1318,N_1172);
nand U2226 (N_2226,N_1009,N_1738);
nor U2227 (N_2227,N_1847,N_1219);
or U2228 (N_2228,N_1624,N_1299);
or U2229 (N_2229,N_1231,N_1611);
nor U2230 (N_2230,N_1966,N_1963);
xor U2231 (N_2231,N_1089,N_1126);
nand U2232 (N_2232,N_1035,N_1513);
and U2233 (N_2233,N_1071,N_1481);
nor U2234 (N_2234,N_1947,N_1762);
nand U2235 (N_2235,N_1137,N_1061);
nor U2236 (N_2236,N_1023,N_1413);
nand U2237 (N_2237,N_1471,N_1715);
or U2238 (N_2238,N_1620,N_1920);
and U2239 (N_2239,N_1376,N_1628);
or U2240 (N_2240,N_1507,N_1151);
and U2241 (N_2241,N_1853,N_1452);
nand U2242 (N_2242,N_1895,N_1553);
nor U2243 (N_2243,N_1741,N_1185);
nand U2244 (N_2244,N_1610,N_1241);
nand U2245 (N_2245,N_1946,N_1645);
and U2246 (N_2246,N_1501,N_1930);
and U2247 (N_2247,N_1863,N_1214);
nor U2248 (N_2248,N_1844,N_1253);
or U2249 (N_2249,N_1113,N_1444);
nor U2250 (N_2250,N_1453,N_1746);
or U2251 (N_2251,N_1497,N_1913);
nor U2252 (N_2252,N_1213,N_1570);
nor U2253 (N_2253,N_1886,N_1311);
nand U2254 (N_2254,N_1640,N_1487);
nand U2255 (N_2255,N_1082,N_1716);
xnor U2256 (N_2256,N_1751,N_1803);
nand U2257 (N_2257,N_1871,N_1093);
or U2258 (N_2258,N_1196,N_1160);
or U2259 (N_2259,N_1530,N_1704);
nor U2260 (N_2260,N_1230,N_1625);
nand U2261 (N_2261,N_1928,N_1201);
and U2262 (N_2262,N_1394,N_1725);
or U2263 (N_2263,N_1668,N_1333);
or U2264 (N_2264,N_1902,N_1945);
or U2265 (N_2265,N_1511,N_1911);
nor U2266 (N_2266,N_1815,N_1290);
or U2267 (N_2267,N_1182,N_1656);
or U2268 (N_2268,N_1222,N_1081);
nand U2269 (N_2269,N_1401,N_1353);
nor U2270 (N_2270,N_1025,N_1466);
nor U2271 (N_2271,N_1646,N_1065);
or U2272 (N_2272,N_1961,N_1542);
and U2273 (N_2273,N_1247,N_1399);
nand U2274 (N_2274,N_1202,N_1516);
and U2275 (N_2275,N_1707,N_1387);
nand U2276 (N_2276,N_1826,N_1672);
nor U2277 (N_2277,N_1095,N_1181);
and U2278 (N_2278,N_1410,N_1845);
and U2279 (N_2279,N_1414,N_1173);
and U2280 (N_2280,N_1953,N_1875);
nand U2281 (N_2281,N_1775,N_1698);
or U2282 (N_2282,N_1192,N_1150);
or U2283 (N_2283,N_1280,N_1421);
and U2284 (N_2284,N_1448,N_1641);
nand U2285 (N_2285,N_1046,N_1566);
nor U2286 (N_2286,N_1430,N_1518);
nand U2287 (N_2287,N_1633,N_1208);
nor U2288 (N_2288,N_1063,N_1157);
and U2289 (N_2289,N_1418,N_1764);
nand U2290 (N_2290,N_1904,N_1987);
xor U2291 (N_2291,N_1673,N_1162);
and U2292 (N_2292,N_1985,N_1167);
nand U2293 (N_2293,N_1609,N_1878);
nor U2294 (N_2294,N_1341,N_1193);
nand U2295 (N_2295,N_1568,N_1352);
nor U2296 (N_2296,N_1424,N_1386);
nor U2297 (N_2297,N_1906,N_1116);
or U2298 (N_2298,N_1517,N_1279);
and U2299 (N_2299,N_1101,N_1567);
and U2300 (N_2300,N_1790,N_1703);
and U2301 (N_2301,N_1260,N_1307);
nand U2302 (N_2302,N_1944,N_1922);
nand U2303 (N_2303,N_1359,N_1660);
and U2304 (N_2304,N_1103,N_1859);
nor U2305 (N_2305,N_1293,N_1534);
xor U2306 (N_2306,N_1268,N_1076);
nand U2307 (N_2307,N_1422,N_1022);
and U2308 (N_2308,N_1415,N_1218);
and U2309 (N_2309,N_1036,N_1541);
nand U2310 (N_2310,N_1144,N_1766);
nor U2311 (N_2311,N_1814,N_1713);
and U2312 (N_2312,N_1272,N_1524);
or U2313 (N_2313,N_1769,N_1319);
nor U2314 (N_2314,N_1630,N_1686);
and U2315 (N_2315,N_1283,N_1869);
or U2316 (N_2316,N_1486,N_1589);
nor U2317 (N_2317,N_1075,N_1383);
xnor U2318 (N_2318,N_1256,N_1371);
nand U2319 (N_2319,N_1515,N_1043);
or U2320 (N_2320,N_1068,N_1340);
or U2321 (N_2321,N_1349,N_1918);
or U2322 (N_2322,N_1806,N_1128);
nand U2323 (N_2323,N_1265,N_1551);
nor U2324 (N_2324,N_1670,N_1066);
and U2325 (N_2325,N_1648,N_1155);
nor U2326 (N_2326,N_1184,N_1261);
or U2327 (N_2327,N_1514,N_1200);
nor U2328 (N_2328,N_1480,N_1425);
and U2329 (N_2329,N_1039,N_1634);
or U2330 (N_2330,N_1658,N_1695);
nand U2331 (N_2331,N_1949,N_1236);
nor U2332 (N_2332,N_1639,N_1956);
xor U2333 (N_2333,N_1234,N_1940);
nor U2334 (N_2334,N_1080,N_1273);
and U2335 (N_2335,N_1087,N_1332);
or U2336 (N_2336,N_1600,N_1696);
nor U2337 (N_2337,N_1682,N_1976);
and U2338 (N_2338,N_1525,N_1412);
nor U2339 (N_2339,N_1779,N_1314);
or U2340 (N_2340,N_1040,N_1096);
or U2341 (N_2341,N_1749,N_1365);
and U2342 (N_2342,N_1125,N_1502);
and U2343 (N_2343,N_1881,N_1588);
or U2344 (N_2344,N_1563,N_1086);
and U2345 (N_2345,N_1485,N_1373);
nor U2346 (N_2346,N_1870,N_1149);
and U2347 (N_2347,N_1099,N_1500);
and U2348 (N_2348,N_1680,N_1586);
or U2349 (N_2349,N_1298,N_1984);
nor U2350 (N_2350,N_1450,N_1000);
or U2351 (N_2351,N_1426,N_1934);
nor U2352 (N_2352,N_1860,N_1007);
or U2353 (N_2353,N_1651,N_1932);
and U2354 (N_2354,N_1249,N_1041);
or U2355 (N_2355,N_1276,N_1406);
and U2356 (N_2356,N_1305,N_1602);
and U2357 (N_2357,N_1923,N_1107);
or U2358 (N_2358,N_1390,N_1866);
nor U2359 (N_2359,N_1786,N_1164);
nor U2360 (N_2360,N_1073,N_1119);
nand U2361 (N_2361,N_1021,N_1888);
and U2362 (N_2362,N_1124,N_1106);
xnor U2363 (N_2363,N_1540,N_1929);
nor U2364 (N_2364,N_1755,N_1893);
or U2365 (N_2365,N_1161,N_1842);
or U2366 (N_2366,N_1926,N_1237);
nor U2367 (N_2367,N_1692,N_1153);
and U2368 (N_2368,N_1372,N_1979);
and U2369 (N_2369,N_1732,N_1449);
or U2370 (N_2370,N_1623,N_1168);
xnor U2371 (N_2371,N_1069,N_1259);
nor U2372 (N_2372,N_1462,N_1130);
or U2373 (N_2373,N_1788,N_1330);
nor U2374 (N_2374,N_1509,N_1579);
or U2375 (N_2375,N_1158,N_1972);
nor U2376 (N_2376,N_1950,N_1689);
xnor U2377 (N_2377,N_1523,N_1527);
nand U2378 (N_2378,N_1747,N_1032);
and U2379 (N_2379,N_1783,N_1295);
nor U2380 (N_2380,N_1499,N_1233);
or U2381 (N_2381,N_1622,N_1528);
and U2382 (N_2382,N_1770,N_1594);
and U2383 (N_2383,N_1287,N_1446);
or U2384 (N_2384,N_1226,N_1220);
and U2385 (N_2385,N_1504,N_1407);
and U2386 (N_2386,N_1194,N_1796);
nand U2387 (N_2387,N_1890,N_1605);
or U2388 (N_2388,N_1885,N_1141);
nor U2389 (N_2389,N_1362,N_1827);
or U2390 (N_2390,N_1996,N_1195);
or U2391 (N_2391,N_1304,N_1597);
and U2392 (N_2392,N_1331,N_1240);
xnor U2393 (N_2393,N_1120,N_1498);
and U2394 (N_2394,N_1564,N_1317);
nand U2395 (N_2395,N_1626,N_1047);
and U2396 (N_2396,N_1701,N_1519);
or U2397 (N_2397,N_1590,N_1456);
and U2398 (N_2398,N_1728,N_1358);
or U2399 (N_2399,N_1671,N_1475);
or U2400 (N_2400,N_1560,N_1051);
nor U2401 (N_2401,N_1765,N_1108);
and U2402 (N_2402,N_1416,N_1850);
or U2403 (N_2403,N_1134,N_1669);
nand U2404 (N_2404,N_1050,N_1300);
and U2405 (N_2405,N_1382,N_1490);
nor U2406 (N_2406,N_1675,N_1604);
nor U2407 (N_2407,N_1529,N_1802);
nand U2408 (N_2408,N_1756,N_1771);
or U2409 (N_2409,N_1935,N_1819);
and U2410 (N_2410,N_1245,N_1915);
xor U2411 (N_2411,N_1468,N_1636);
or U2412 (N_2412,N_1315,N_1997);
or U2413 (N_2413,N_1995,N_1595);
nand U2414 (N_2414,N_1109,N_1709);
and U2415 (N_2415,N_1370,N_1535);
nand U2416 (N_2416,N_1458,N_1914);
nand U2417 (N_2417,N_1026,N_1463);
nand U2418 (N_2418,N_1493,N_1492);
nor U2419 (N_2419,N_1004,N_1557);
and U2420 (N_2420,N_1244,N_1960);
or U2421 (N_2421,N_1808,N_1478);
nand U2422 (N_2422,N_1781,N_1186);
nand U2423 (N_2423,N_1791,N_1335);
and U2424 (N_2424,N_1483,N_1045);
nor U2425 (N_2425,N_1187,N_1166);
nand U2426 (N_2426,N_1857,N_1308);
or U2427 (N_2427,N_1754,N_1512);
nand U2428 (N_2428,N_1720,N_1255);
or U2429 (N_2429,N_1753,N_1019);
xnor U2430 (N_2430,N_1348,N_1900);
nand U2431 (N_2431,N_1322,N_1212);
and U2432 (N_2432,N_1505,N_1288);
nor U2433 (N_2433,N_1543,N_1536);
nand U2434 (N_2434,N_1874,N_1894);
nand U2435 (N_2435,N_1142,N_1354);
or U2436 (N_2436,N_1129,N_1083);
and U2437 (N_2437,N_1825,N_1433);
nand U2438 (N_2438,N_1442,N_1849);
or U2439 (N_2439,N_1710,N_1404);
nor U2440 (N_2440,N_1197,N_1324);
or U2441 (N_2441,N_1016,N_1758);
nand U2442 (N_2442,N_1037,N_1905);
nor U2443 (N_2443,N_1858,N_1665);
or U2444 (N_2444,N_1379,N_1403);
nor U2445 (N_2445,N_1655,N_1159);
and U2446 (N_2446,N_1455,N_1981);
nor U2447 (N_2447,N_1837,N_1264);
nand U2448 (N_2448,N_1242,N_1583);
nand U2449 (N_2449,N_1320,N_1916);
nor U2450 (N_2450,N_1901,N_1574);
nor U2451 (N_2451,N_1735,N_1384);
xor U2452 (N_2452,N_1105,N_1393);
nand U2453 (N_2453,N_1647,N_1020);
nand U2454 (N_2454,N_1810,N_1165);
nand U2455 (N_2455,N_1880,N_1968);
or U2456 (N_2456,N_1389,N_1957);
nor U2457 (N_2457,N_1649,N_1667);
nor U2458 (N_2458,N_1067,N_1522);
and U2459 (N_2459,N_1702,N_1970);
and U2460 (N_2460,N_1577,N_1607);
xnor U2461 (N_2461,N_1005,N_1785);
xor U2462 (N_2462,N_1711,N_1465);
nand U2463 (N_2463,N_1794,N_1818);
or U2464 (N_2464,N_1495,N_1773);
and U2465 (N_2465,N_1714,N_1552);
xnor U2466 (N_2466,N_1772,N_1488);
xor U2467 (N_2467,N_1903,N_1638);
nor U2468 (N_2468,N_1439,N_1889);
nand U2469 (N_2469,N_1657,N_1955);
nand U2470 (N_2470,N_1909,N_1263);
nor U2471 (N_2471,N_1408,N_1834);
nand U2472 (N_2472,N_1309,N_1254);
and U2473 (N_2473,N_1897,N_1011);
and U2474 (N_2474,N_1489,N_1974);
and U2475 (N_2475,N_1274,N_1784);
and U2476 (N_2476,N_1763,N_1296);
nor U2477 (N_2477,N_1437,N_1175);
and U2478 (N_2478,N_1411,N_1931);
nand U2479 (N_2479,N_1804,N_1676);
nand U2480 (N_2480,N_1303,N_1342);
nand U2481 (N_2481,N_1188,N_1146);
nor U2482 (N_2482,N_1377,N_1374);
nor U2483 (N_2483,N_1999,N_1064);
and U2484 (N_2484,N_1606,N_1578);
or U2485 (N_2485,N_1601,N_1434);
and U2486 (N_2486,N_1856,N_1933);
and U2487 (N_2487,N_1435,N_1123);
nand U2488 (N_2488,N_1663,N_1546);
or U2489 (N_2489,N_1873,N_1798);
and U2490 (N_2490,N_1580,N_1822);
and U2491 (N_2491,N_1381,N_1813);
nand U2492 (N_2492,N_1718,N_1006);
nor U2493 (N_2493,N_1719,N_1587);
nor U2494 (N_2494,N_1392,N_1284);
nor U2495 (N_2495,N_1867,N_1921);
and U2496 (N_2496,N_1355,N_1533);
or U2497 (N_2497,N_1865,N_1001);
nand U2498 (N_2498,N_1464,N_1662);
nand U2499 (N_2499,N_1457,N_1147);
xnor U2500 (N_2500,N_1100,N_1021);
and U2501 (N_2501,N_1275,N_1389);
nand U2502 (N_2502,N_1399,N_1471);
nand U2503 (N_2503,N_1707,N_1334);
nor U2504 (N_2504,N_1953,N_1599);
nand U2505 (N_2505,N_1170,N_1146);
nand U2506 (N_2506,N_1060,N_1302);
nor U2507 (N_2507,N_1917,N_1786);
xor U2508 (N_2508,N_1827,N_1005);
and U2509 (N_2509,N_1762,N_1051);
xnor U2510 (N_2510,N_1536,N_1403);
nor U2511 (N_2511,N_1912,N_1269);
or U2512 (N_2512,N_1733,N_1555);
or U2513 (N_2513,N_1379,N_1226);
and U2514 (N_2514,N_1506,N_1222);
nand U2515 (N_2515,N_1762,N_1439);
and U2516 (N_2516,N_1645,N_1568);
and U2517 (N_2517,N_1080,N_1678);
nand U2518 (N_2518,N_1638,N_1223);
nor U2519 (N_2519,N_1258,N_1506);
or U2520 (N_2520,N_1324,N_1533);
nand U2521 (N_2521,N_1044,N_1020);
nor U2522 (N_2522,N_1894,N_1674);
nor U2523 (N_2523,N_1990,N_1339);
xnor U2524 (N_2524,N_1157,N_1445);
or U2525 (N_2525,N_1011,N_1338);
nor U2526 (N_2526,N_1670,N_1057);
nor U2527 (N_2527,N_1690,N_1510);
nor U2528 (N_2528,N_1426,N_1677);
xnor U2529 (N_2529,N_1836,N_1906);
nor U2530 (N_2530,N_1783,N_1246);
or U2531 (N_2531,N_1875,N_1823);
nand U2532 (N_2532,N_1357,N_1897);
nand U2533 (N_2533,N_1209,N_1863);
nand U2534 (N_2534,N_1698,N_1472);
and U2535 (N_2535,N_1317,N_1741);
nor U2536 (N_2536,N_1917,N_1249);
nand U2537 (N_2537,N_1879,N_1368);
nand U2538 (N_2538,N_1592,N_1435);
nand U2539 (N_2539,N_1913,N_1542);
nor U2540 (N_2540,N_1588,N_1734);
nand U2541 (N_2541,N_1987,N_1440);
and U2542 (N_2542,N_1832,N_1346);
nand U2543 (N_2543,N_1924,N_1907);
nor U2544 (N_2544,N_1584,N_1157);
or U2545 (N_2545,N_1345,N_1861);
and U2546 (N_2546,N_1598,N_1993);
and U2547 (N_2547,N_1777,N_1489);
nor U2548 (N_2548,N_1443,N_1687);
nor U2549 (N_2549,N_1507,N_1369);
or U2550 (N_2550,N_1166,N_1672);
nand U2551 (N_2551,N_1167,N_1410);
nand U2552 (N_2552,N_1464,N_1025);
or U2553 (N_2553,N_1523,N_1349);
nand U2554 (N_2554,N_1037,N_1702);
xnor U2555 (N_2555,N_1534,N_1887);
nor U2556 (N_2556,N_1584,N_1062);
nor U2557 (N_2557,N_1449,N_1279);
nor U2558 (N_2558,N_1726,N_1059);
nand U2559 (N_2559,N_1173,N_1892);
and U2560 (N_2560,N_1995,N_1394);
nor U2561 (N_2561,N_1249,N_1798);
or U2562 (N_2562,N_1181,N_1520);
nand U2563 (N_2563,N_1844,N_1450);
or U2564 (N_2564,N_1142,N_1691);
nor U2565 (N_2565,N_1907,N_1989);
nand U2566 (N_2566,N_1343,N_1009);
nor U2567 (N_2567,N_1544,N_1284);
and U2568 (N_2568,N_1613,N_1119);
and U2569 (N_2569,N_1201,N_1256);
or U2570 (N_2570,N_1965,N_1148);
nand U2571 (N_2571,N_1790,N_1943);
nand U2572 (N_2572,N_1817,N_1154);
nor U2573 (N_2573,N_1666,N_1470);
nor U2574 (N_2574,N_1775,N_1737);
and U2575 (N_2575,N_1695,N_1140);
and U2576 (N_2576,N_1640,N_1454);
or U2577 (N_2577,N_1097,N_1146);
xnor U2578 (N_2578,N_1368,N_1355);
nand U2579 (N_2579,N_1949,N_1852);
or U2580 (N_2580,N_1268,N_1701);
xnor U2581 (N_2581,N_1121,N_1252);
xnor U2582 (N_2582,N_1378,N_1337);
and U2583 (N_2583,N_1364,N_1785);
and U2584 (N_2584,N_1402,N_1835);
and U2585 (N_2585,N_1920,N_1567);
nand U2586 (N_2586,N_1697,N_1210);
xor U2587 (N_2587,N_1263,N_1521);
nor U2588 (N_2588,N_1813,N_1785);
or U2589 (N_2589,N_1904,N_1823);
nor U2590 (N_2590,N_1273,N_1235);
or U2591 (N_2591,N_1952,N_1338);
or U2592 (N_2592,N_1122,N_1284);
and U2593 (N_2593,N_1588,N_1870);
nor U2594 (N_2594,N_1964,N_1444);
and U2595 (N_2595,N_1351,N_1651);
and U2596 (N_2596,N_1973,N_1513);
or U2597 (N_2597,N_1961,N_1392);
nor U2598 (N_2598,N_1847,N_1674);
nor U2599 (N_2599,N_1494,N_1958);
or U2600 (N_2600,N_1771,N_1427);
or U2601 (N_2601,N_1845,N_1317);
nor U2602 (N_2602,N_1409,N_1334);
and U2603 (N_2603,N_1612,N_1776);
or U2604 (N_2604,N_1310,N_1228);
and U2605 (N_2605,N_1890,N_1802);
or U2606 (N_2606,N_1971,N_1767);
and U2607 (N_2607,N_1577,N_1429);
nor U2608 (N_2608,N_1863,N_1119);
nand U2609 (N_2609,N_1939,N_1275);
or U2610 (N_2610,N_1186,N_1990);
nor U2611 (N_2611,N_1105,N_1315);
or U2612 (N_2612,N_1870,N_1404);
nand U2613 (N_2613,N_1951,N_1712);
xor U2614 (N_2614,N_1881,N_1147);
nand U2615 (N_2615,N_1434,N_1917);
or U2616 (N_2616,N_1685,N_1973);
xnor U2617 (N_2617,N_1459,N_1761);
nor U2618 (N_2618,N_1385,N_1133);
or U2619 (N_2619,N_1144,N_1111);
xor U2620 (N_2620,N_1241,N_1947);
and U2621 (N_2621,N_1250,N_1776);
nand U2622 (N_2622,N_1945,N_1632);
nand U2623 (N_2623,N_1924,N_1194);
and U2624 (N_2624,N_1818,N_1510);
and U2625 (N_2625,N_1961,N_1233);
nand U2626 (N_2626,N_1774,N_1414);
and U2627 (N_2627,N_1108,N_1106);
nor U2628 (N_2628,N_1777,N_1194);
or U2629 (N_2629,N_1058,N_1044);
nand U2630 (N_2630,N_1707,N_1374);
xor U2631 (N_2631,N_1422,N_1239);
nor U2632 (N_2632,N_1283,N_1246);
nand U2633 (N_2633,N_1742,N_1702);
or U2634 (N_2634,N_1442,N_1529);
and U2635 (N_2635,N_1393,N_1565);
and U2636 (N_2636,N_1375,N_1702);
nand U2637 (N_2637,N_1679,N_1346);
nand U2638 (N_2638,N_1340,N_1850);
nor U2639 (N_2639,N_1896,N_1075);
and U2640 (N_2640,N_1100,N_1121);
and U2641 (N_2641,N_1639,N_1077);
nand U2642 (N_2642,N_1613,N_1154);
or U2643 (N_2643,N_1432,N_1076);
nand U2644 (N_2644,N_1292,N_1284);
nand U2645 (N_2645,N_1204,N_1831);
nand U2646 (N_2646,N_1898,N_1951);
nor U2647 (N_2647,N_1063,N_1282);
and U2648 (N_2648,N_1157,N_1969);
nor U2649 (N_2649,N_1221,N_1172);
nand U2650 (N_2650,N_1452,N_1408);
and U2651 (N_2651,N_1613,N_1834);
or U2652 (N_2652,N_1912,N_1135);
and U2653 (N_2653,N_1857,N_1934);
and U2654 (N_2654,N_1876,N_1323);
xor U2655 (N_2655,N_1918,N_1107);
nand U2656 (N_2656,N_1757,N_1624);
nand U2657 (N_2657,N_1082,N_1423);
and U2658 (N_2658,N_1587,N_1471);
xor U2659 (N_2659,N_1424,N_1697);
nor U2660 (N_2660,N_1565,N_1138);
and U2661 (N_2661,N_1319,N_1234);
nor U2662 (N_2662,N_1893,N_1436);
nand U2663 (N_2663,N_1532,N_1517);
or U2664 (N_2664,N_1460,N_1983);
nand U2665 (N_2665,N_1162,N_1768);
nand U2666 (N_2666,N_1859,N_1382);
nand U2667 (N_2667,N_1756,N_1237);
nand U2668 (N_2668,N_1545,N_1626);
nand U2669 (N_2669,N_1271,N_1020);
nor U2670 (N_2670,N_1845,N_1334);
nor U2671 (N_2671,N_1864,N_1534);
and U2672 (N_2672,N_1360,N_1236);
nand U2673 (N_2673,N_1765,N_1484);
nor U2674 (N_2674,N_1143,N_1125);
nor U2675 (N_2675,N_1817,N_1132);
and U2676 (N_2676,N_1816,N_1753);
and U2677 (N_2677,N_1940,N_1859);
or U2678 (N_2678,N_1708,N_1831);
or U2679 (N_2679,N_1456,N_1337);
and U2680 (N_2680,N_1777,N_1918);
and U2681 (N_2681,N_1941,N_1042);
nand U2682 (N_2682,N_1737,N_1425);
or U2683 (N_2683,N_1436,N_1969);
and U2684 (N_2684,N_1995,N_1926);
nand U2685 (N_2685,N_1643,N_1670);
nand U2686 (N_2686,N_1289,N_1077);
or U2687 (N_2687,N_1664,N_1747);
nor U2688 (N_2688,N_1039,N_1231);
xor U2689 (N_2689,N_1502,N_1169);
xnor U2690 (N_2690,N_1677,N_1496);
nand U2691 (N_2691,N_1428,N_1194);
nor U2692 (N_2692,N_1749,N_1896);
or U2693 (N_2693,N_1260,N_1229);
nand U2694 (N_2694,N_1879,N_1022);
nor U2695 (N_2695,N_1663,N_1449);
nor U2696 (N_2696,N_1981,N_1600);
or U2697 (N_2697,N_1577,N_1421);
or U2698 (N_2698,N_1578,N_1840);
nor U2699 (N_2699,N_1907,N_1077);
xor U2700 (N_2700,N_1585,N_1064);
nand U2701 (N_2701,N_1460,N_1212);
or U2702 (N_2702,N_1196,N_1933);
nand U2703 (N_2703,N_1199,N_1468);
and U2704 (N_2704,N_1251,N_1072);
or U2705 (N_2705,N_1437,N_1999);
nand U2706 (N_2706,N_1091,N_1033);
and U2707 (N_2707,N_1151,N_1907);
nand U2708 (N_2708,N_1589,N_1796);
nor U2709 (N_2709,N_1392,N_1651);
nand U2710 (N_2710,N_1641,N_1655);
and U2711 (N_2711,N_1989,N_1870);
and U2712 (N_2712,N_1234,N_1211);
or U2713 (N_2713,N_1547,N_1734);
or U2714 (N_2714,N_1857,N_1433);
nor U2715 (N_2715,N_1591,N_1794);
and U2716 (N_2716,N_1265,N_1146);
and U2717 (N_2717,N_1520,N_1879);
and U2718 (N_2718,N_1625,N_1598);
and U2719 (N_2719,N_1349,N_1699);
and U2720 (N_2720,N_1679,N_1010);
xor U2721 (N_2721,N_1686,N_1152);
and U2722 (N_2722,N_1231,N_1446);
xor U2723 (N_2723,N_1205,N_1031);
or U2724 (N_2724,N_1164,N_1601);
nand U2725 (N_2725,N_1080,N_1730);
or U2726 (N_2726,N_1113,N_1971);
xnor U2727 (N_2727,N_1517,N_1670);
nor U2728 (N_2728,N_1935,N_1597);
nand U2729 (N_2729,N_1807,N_1289);
nand U2730 (N_2730,N_1359,N_1691);
nor U2731 (N_2731,N_1550,N_1736);
or U2732 (N_2732,N_1448,N_1513);
and U2733 (N_2733,N_1543,N_1524);
nand U2734 (N_2734,N_1314,N_1067);
and U2735 (N_2735,N_1101,N_1315);
xnor U2736 (N_2736,N_1264,N_1405);
and U2737 (N_2737,N_1799,N_1257);
or U2738 (N_2738,N_1171,N_1955);
nor U2739 (N_2739,N_1744,N_1933);
nand U2740 (N_2740,N_1538,N_1503);
nand U2741 (N_2741,N_1383,N_1015);
nand U2742 (N_2742,N_1090,N_1449);
and U2743 (N_2743,N_1670,N_1156);
or U2744 (N_2744,N_1814,N_1989);
or U2745 (N_2745,N_1939,N_1485);
or U2746 (N_2746,N_1272,N_1387);
nand U2747 (N_2747,N_1097,N_1647);
or U2748 (N_2748,N_1868,N_1988);
nand U2749 (N_2749,N_1341,N_1454);
nor U2750 (N_2750,N_1710,N_1891);
nand U2751 (N_2751,N_1453,N_1276);
nor U2752 (N_2752,N_1184,N_1136);
nor U2753 (N_2753,N_1659,N_1102);
nor U2754 (N_2754,N_1975,N_1424);
nor U2755 (N_2755,N_1172,N_1720);
nand U2756 (N_2756,N_1495,N_1981);
nor U2757 (N_2757,N_1476,N_1657);
nor U2758 (N_2758,N_1215,N_1949);
and U2759 (N_2759,N_1791,N_1177);
or U2760 (N_2760,N_1637,N_1804);
nand U2761 (N_2761,N_1843,N_1502);
nor U2762 (N_2762,N_1562,N_1406);
nor U2763 (N_2763,N_1764,N_1440);
and U2764 (N_2764,N_1574,N_1509);
or U2765 (N_2765,N_1481,N_1734);
nor U2766 (N_2766,N_1273,N_1361);
nand U2767 (N_2767,N_1903,N_1628);
nor U2768 (N_2768,N_1998,N_1185);
and U2769 (N_2769,N_1401,N_1847);
or U2770 (N_2770,N_1591,N_1428);
and U2771 (N_2771,N_1730,N_1553);
and U2772 (N_2772,N_1795,N_1769);
or U2773 (N_2773,N_1496,N_1709);
nand U2774 (N_2774,N_1683,N_1020);
xor U2775 (N_2775,N_1421,N_1469);
nor U2776 (N_2776,N_1861,N_1724);
or U2777 (N_2777,N_1573,N_1103);
or U2778 (N_2778,N_1829,N_1551);
and U2779 (N_2779,N_1930,N_1149);
nor U2780 (N_2780,N_1460,N_1481);
and U2781 (N_2781,N_1071,N_1543);
xor U2782 (N_2782,N_1447,N_1159);
nand U2783 (N_2783,N_1562,N_1251);
nand U2784 (N_2784,N_1154,N_1019);
and U2785 (N_2785,N_1145,N_1288);
and U2786 (N_2786,N_1341,N_1429);
nand U2787 (N_2787,N_1530,N_1964);
and U2788 (N_2788,N_1962,N_1890);
nor U2789 (N_2789,N_1113,N_1471);
nor U2790 (N_2790,N_1145,N_1507);
nor U2791 (N_2791,N_1027,N_1198);
or U2792 (N_2792,N_1636,N_1408);
and U2793 (N_2793,N_1689,N_1387);
or U2794 (N_2794,N_1485,N_1658);
nand U2795 (N_2795,N_1463,N_1090);
nand U2796 (N_2796,N_1585,N_1834);
nand U2797 (N_2797,N_1716,N_1525);
nor U2798 (N_2798,N_1246,N_1748);
nand U2799 (N_2799,N_1828,N_1007);
and U2800 (N_2800,N_1989,N_1917);
nor U2801 (N_2801,N_1526,N_1868);
and U2802 (N_2802,N_1780,N_1729);
and U2803 (N_2803,N_1279,N_1382);
nand U2804 (N_2804,N_1718,N_1763);
or U2805 (N_2805,N_1217,N_1657);
nor U2806 (N_2806,N_1678,N_1818);
nor U2807 (N_2807,N_1328,N_1698);
nand U2808 (N_2808,N_1423,N_1670);
nand U2809 (N_2809,N_1234,N_1664);
nor U2810 (N_2810,N_1157,N_1447);
nand U2811 (N_2811,N_1197,N_1034);
xnor U2812 (N_2812,N_1881,N_1175);
and U2813 (N_2813,N_1711,N_1520);
and U2814 (N_2814,N_1448,N_1521);
nor U2815 (N_2815,N_1442,N_1890);
nand U2816 (N_2816,N_1139,N_1584);
nand U2817 (N_2817,N_1605,N_1196);
nor U2818 (N_2818,N_1876,N_1209);
nand U2819 (N_2819,N_1314,N_1328);
nor U2820 (N_2820,N_1591,N_1300);
or U2821 (N_2821,N_1968,N_1704);
nand U2822 (N_2822,N_1819,N_1794);
nand U2823 (N_2823,N_1723,N_1189);
nand U2824 (N_2824,N_1561,N_1865);
xnor U2825 (N_2825,N_1807,N_1882);
or U2826 (N_2826,N_1944,N_1469);
nand U2827 (N_2827,N_1849,N_1465);
nand U2828 (N_2828,N_1433,N_1582);
and U2829 (N_2829,N_1800,N_1356);
xnor U2830 (N_2830,N_1980,N_1484);
nand U2831 (N_2831,N_1226,N_1742);
nand U2832 (N_2832,N_1694,N_1156);
nand U2833 (N_2833,N_1576,N_1533);
nor U2834 (N_2834,N_1563,N_1553);
and U2835 (N_2835,N_1296,N_1917);
and U2836 (N_2836,N_1314,N_1028);
nor U2837 (N_2837,N_1717,N_1951);
and U2838 (N_2838,N_1502,N_1058);
nor U2839 (N_2839,N_1042,N_1533);
and U2840 (N_2840,N_1849,N_1928);
xnor U2841 (N_2841,N_1588,N_1216);
xnor U2842 (N_2842,N_1291,N_1365);
nand U2843 (N_2843,N_1113,N_1492);
or U2844 (N_2844,N_1496,N_1746);
nor U2845 (N_2845,N_1945,N_1542);
nor U2846 (N_2846,N_1894,N_1062);
nand U2847 (N_2847,N_1066,N_1355);
or U2848 (N_2848,N_1424,N_1858);
nand U2849 (N_2849,N_1215,N_1088);
nor U2850 (N_2850,N_1306,N_1480);
or U2851 (N_2851,N_1635,N_1673);
nand U2852 (N_2852,N_1218,N_1947);
or U2853 (N_2853,N_1693,N_1503);
nor U2854 (N_2854,N_1972,N_1192);
nor U2855 (N_2855,N_1279,N_1831);
xnor U2856 (N_2856,N_1402,N_1423);
and U2857 (N_2857,N_1289,N_1339);
nor U2858 (N_2858,N_1829,N_1863);
xor U2859 (N_2859,N_1921,N_1842);
or U2860 (N_2860,N_1358,N_1831);
nor U2861 (N_2861,N_1724,N_1121);
nand U2862 (N_2862,N_1151,N_1768);
or U2863 (N_2863,N_1550,N_1000);
xor U2864 (N_2864,N_1753,N_1324);
nor U2865 (N_2865,N_1341,N_1959);
or U2866 (N_2866,N_1463,N_1180);
nand U2867 (N_2867,N_1671,N_1207);
nor U2868 (N_2868,N_1611,N_1937);
xor U2869 (N_2869,N_1005,N_1043);
nor U2870 (N_2870,N_1611,N_1307);
or U2871 (N_2871,N_1394,N_1670);
or U2872 (N_2872,N_1008,N_1948);
and U2873 (N_2873,N_1329,N_1753);
nor U2874 (N_2874,N_1788,N_1048);
and U2875 (N_2875,N_1474,N_1498);
nor U2876 (N_2876,N_1163,N_1181);
or U2877 (N_2877,N_1029,N_1650);
nand U2878 (N_2878,N_1772,N_1320);
and U2879 (N_2879,N_1237,N_1851);
nor U2880 (N_2880,N_1702,N_1938);
and U2881 (N_2881,N_1185,N_1649);
and U2882 (N_2882,N_1365,N_1021);
nand U2883 (N_2883,N_1563,N_1471);
nor U2884 (N_2884,N_1979,N_1613);
nand U2885 (N_2885,N_1881,N_1113);
nor U2886 (N_2886,N_1320,N_1969);
nor U2887 (N_2887,N_1993,N_1537);
or U2888 (N_2888,N_1870,N_1846);
and U2889 (N_2889,N_1862,N_1544);
and U2890 (N_2890,N_1980,N_1582);
or U2891 (N_2891,N_1224,N_1075);
nand U2892 (N_2892,N_1485,N_1606);
nor U2893 (N_2893,N_1813,N_1424);
or U2894 (N_2894,N_1016,N_1468);
nor U2895 (N_2895,N_1726,N_1426);
and U2896 (N_2896,N_1072,N_1746);
xor U2897 (N_2897,N_1340,N_1344);
nor U2898 (N_2898,N_1722,N_1745);
and U2899 (N_2899,N_1769,N_1086);
or U2900 (N_2900,N_1440,N_1759);
and U2901 (N_2901,N_1928,N_1500);
and U2902 (N_2902,N_1265,N_1702);
nand U2903 (N_2903,N_1529,N_1895);
nand U2904 (N_2904,N_1379,N_1446);
nor U2905 (N_2905,N_1137,N_1505);
or U2906 (N_2906,N_1685,N_1785);
and U2907 (N_2907,N_1741,N_1180);
and U2908 (N_2908,N_1838,N_1565);
nand U2909 (N_2909,N_1352,N_1855);
xor U2910 (N_2910,N_1837,N_1906);
and U2911 (N_2911,N_1973,N_1884);
nand U2912 (N_2912,N_1066,N_1151);
nor U2913 (N_2913,N_1977,N_1194);
nor U2914 (N_2914,N_1947,N_1970);
or U2915 (N_2915,N_1962,N_1689);
and U2916 (N_2916,N_1581,N_1057);
or U2917 (N_2917,N_1849,N_1487);
nand U2918 (N_2918,N_1233,N_1740);
xnor U2919 (N_2919,N_1255,N_1010);
and U2920 (N_2920,N_1844,N_1315);
and U2921 (N_2921,N_1050,N_1990);
nand U2922 (N_2922,N_1799,N_1041);
or U2923 (N_2923,N_1232,N_1404);
nor U2924 (N_2924,N_1319,N_1757);
nor U2925 (N_2925,N_1237,N_1717);
or U2926 (N_2926,N_1735,N_1843);
or U2927 (N_2927,N_1677,N_1650);
xnor U2928 (N_2928,N_1580,N_1102);
or U2929 (N_2929,N_1853,N_1255);
or U2930 (N_2930,N_1654,N_1903);
xor U2931 (N_2931,N_1788,N_1030);
nand U2932 (N_2932,N_1533,N_1263);
nand U2933 (N_2933,N_1719,N_1617);
and U2934 (N_2934,N_1172,N_1710);
nand U2935 (N_2935,N_1104,N_1268);
and U2936 (N_2936,N_1945,N_1730);
nor U2937 (N_2937,N_1983,N_1295);
nor U2938 (N_2938,N_1647,N_1189);
and U2939 (N_2939,N_1346,N_1245);
or U2940 (N_2940,N_1315,N_1669);
or U2941 (N_2941,N_1197,N_1487);
or U2942 (N_2942,N_1263,N_1810);
nor U2943 (N_2943,N_1764,N_1638);
nor U2944 (N_2944,N_1877,N_1425);
nand U2945 (N_2945,N_1662,N_1944);
or U2946 (N_2946,N_1983,N_1464);
and U2947 (N_2947,N_1221,N_1870);
nor U2948 (N_2948,N_1474,N_1683);
or U2949 (N_2949,N_1955,N_1402);
and U2950 (N_2950,N_1605,N_1389);
or U2951 (N_2951,N_1023,N_1769);
and U2952 (N_2952,N_1133,N_1869);
and U2953 (N_2953,N_1873,N_1430);
nor U2954 (N_2954,N_1042,N_1097);
or U2955 (N_2955,N_1690,N_1167);
nor U2956 (N_2956,N_1190,N_1769);
or U2957 (N_2957,N_1479,N_1853);
or U2958 (N_2958,N_1798,N_1687);
nor U2959 (N_2959,N_1008,N_1294);
and U2960 (N_2960,N_1013,N_1891);
or U2961 (N_2961,N_1632,N_1792);
and U2962 (N_2962,N_1251,N_1749);
or U2963 (N_2963,N_1018,N_1025);
or U2964 (N_2964,N_1445,N_1198);
nor U2965 (N_2965,N_1193,N_1399);
nor U2966 (N_2966,N_1065,N_1530);
and U2967 (N_2967,N_1879,N_1620);
or U2968 (N_2968,N_1469,N_1251);
xor U2969 (N_2969,N_1356,N_1766);
nand U2970 (N_2970,N_1374,N_1492);
nor U2971 (N_2971,N_1653,N_1890);
or U2972 (N_2972,N_1382,N_1483);
xor U2973 (N_2973,N_1468,N_1212);
nand U2974 (N_2974,N_1658,N_1241);
nor U2975 (N_2975,N_1848,N_1223);
and U2976 (N_2976,N_1722,N_1433);
or U2977 (N_2977,N_1576,N_1484);
nand U2978 (N_2978,N_1427,N_1118);
or U2979 (N_2979,N_1938,N_1061);
and U2980 (N_2980,N_1169,N_1534);
or U2981 (N_2981,N_1444,N_1245);
and U2982 (N_2982,N_1495,N_1768);
nor U2983 (N_2983,N_1267,N_1434);
xor U2984 (N_2984,N_1694,N_1031);
nor U2985 (N_2985,N_1735,N_1861);
nor U2986 (N_2986,N_1869,N_1284);
nand U2987 (N_2987,N_1415,N_1537);
nor U2988 (N_2988,N_1688,N_1921);
nor U2989 (N_2989,N_1367,N_1028);
or U2990 (N_2990,N_1289,N_1827);
nand U2991 (N_2991,N_1633,N_1672);
nand U2992 (N_2992,N_1040,N_1949);
or U2993 (N_2993,N_1929,N_1827);
and U2994 (N_2994,N_1376,N_1665);
nand U2995 (N_2995,N_1669,N_1550);
nand U2996 (N_2996,N_1498,N_1042);
nand U2997 (N_2997,N_1788,N_1618);
and U2998 (N_2998,N_1992,N_1175);
or U2999 (N_2999,N_1988,N_1901);
nor U3000 (N_3000,N_2179,N_2303);
nor U3001 (N_3001,N_2231,N_2013);
and U3002 (N_3002,N_2030,N_2415);
nor U3003 (N_3003,N_2291,N_2808);
or U3004 (N_3004,N_2929,N_2933);
or U3005 (N_3005,N_2942,N_2698);
xor U3006 (N_3006,N_2785,N_2901);
xor U3007 (N_3007,N_2598,N_2490);
and U3008 (N_3008,N_2920,N_2296);
nand U3009 (N_3009,N_2566,N_2500);
nor U3010 (N_3010,N_2791,N_2936);
or U3011 (N_3011,N_2648,N_2713);
nand U3012 (N_3012,N_2406,N_2905);
nor U3013 (N_3013,N_2056,N_2043);
or U3014 (N_3014,N_2225,N_2565);
nor U3015 (N_3015,N_2268,N_2844);
nor U3016 (N_3016,N_2839,N_2865);
nor U3017 (N_3017,N_2671,N_2174);
nor U3018 (N_3018,N_2053,N_2709);
nand U3019 (N_3019,N_2797,N_2629);
nand U3020 (N_3020,N_2503,N_2887);
nor U3021 (N_3021,N_2343,N_2677);
and U3022 (N_3022,N_2298,N_2872);
or U3023 (N_3023,N_2736,N_2351);
nand U3024 (N_3024,N_2441,N_2201);
xnor U3025 (N_3025,N_2474,N_2224);
and U3026 (N_3026,N_2293,N_2803);
and U3027 (N_3027,N_2238,N_2780);
nor U3028 (N_3028,N_2662,N_2970);
xor U3029 (N_3029,N_2276,N_2232);
nand U3030 (N_3030,N_2955,N_2753);
or U3031 (N_3031,N_2410,N_2317);
nor U3032 (N_3032,N_2842,N_2009);
nand U3033 (N_3033,N_2732,N_2895);
and U3034 (N_3034,N_2524,N_2748);
xnor U3035 (N_3035,N_2483,N_2636);
nand U3036 (N_3036,N_2012,N_2479);
nor U3037 (N_3037,N_2379,N_2337);
or U3038 (N_3038,N_2372,N_2959);
and U3039 (N_3039,N_2658,N_2985);
or U3040 (N_3040,N_2587,N_2850);
xnor U3041 (N_3041,N_2062,N_2127);
and U3042 (N_3042,N_2422,N_2830);
nand U3043 (N_3043,N_2618,N_2237);
nor U3044 (N_3044,N_2586,N_2359);
nand U3045 (N_3045,N_2761,N_2891);
nor U3046 (N_3046,N_2909,N_2172);
and U3047 (N_3047,N_2339,N_2494);
and U3048 (N_3048,N_2064,N_2057);
nand U3049 (N_3049,N_2082,N_2786);
nand U3050 (N_3050,N_2800,N_2570);
and U3051 (N_3051,N_2245,N_2347);
or U3052 (N_3052,N_2621,N_2171);
xor U3053 (N_3053,N_2571,N_2543);
nand U3054 (N_3054,N_2914,N_2605);
nand U3055 (N_3055,N_2390,N_2585);
or U3056 (N_3056,N_2362,N_2038);
and U3057 (N_3057,N_2488,N_2222);
or U3058 (N_3058,N_2823,N_2975);
or U3059 (N_3059,N_2870,N_2793);
nor U3060 (N_3060,N_2555,N_2625);
xnor U3061 (N_3061,N_2788,N_2664);
or U3062 (N_3062,N_2282,N_2158);
xnor U3063 (N_3063,N_2628,N_2663);
xor U3064 (N_3064,N_2350,N_2795);
nor U3065 (N_3065,N_2278,N_2965);
nand U3066 (N_3066,N_2110,N_2463);
nand U3067 (N_3067,N_2416,N_2783);
and U3068 (N_3068,N_2336,N_2502);
xnor U3069 (N_3069,N_2424,N_2049);
or U3070 (N_3070,N_2971,N_2136);
and U3071 (N_3071,N_2655,N_2029);
or U3072 (N_3072,N_2241,N_2468);
nor U3073 (N_3073,N_2335,N_2880);
nand U3074 (N_3074,N_2305,N_2690);
nor U3075 (N_3075,N_2515,N_2094);
xnor U3076 (N_3076,N_2000,N_2608);
or U3077 (N_3077,N_2884,N_2922);
and U3078 (N_3078,N_2024,N_2978);
nand U3079 (N_3079,N_2391,N_2779);
nor U3080 (N_3080,N_2322,N_2584);
nand U3081 (N_3081,N_2097,N_2411);
xor U3082 (N_3082,N_2506,N_2026);
or U3083 (N_3083,N_2686,N_2747);
or U3084 (N_3084,N_2235,N_2845);
nand U3085 (N_3085,N_2363,N_2849);
or U3086 (N_3086,N_2417,N_2617);
nor U3087 (N_3087,N_2561,N_2969);
or U3088 (N_3088,N_2544,N_2752);
and U3089 (N_3089,N_2126,N_2264);
xnor U3090 (N_3090,N_2145,N_2081);
nand U3091 (N_3091,N_2430,N_2270);
nand U3092 (N_3092,N_2011,N_2724);
and U3093 (N_3093,N_2115,N_2934);
nand U3094 (N_3094,N_2284,N_2730);
nand U3095 (N_3095,N_2819,N_2882);
or U3096 (N_3096,N_2279,N_2578);
and U3097 (N_3097,N_2841,N_2691);
nand U3098 (N_3098,N_2679,N_2318);
or U3099 (N_3099,N_2675,N_2700);
xnor U3100 (N_3100,N_2572,N_2715);
xnor U3101 (N_3101,N_2314,N_2722);
nor U3102 (N_3102,N_2414,N_2583);
nand U3103 (N_3103,N_2644,N_2501);
nor U3104 (N_3104,N_2874,N_2159);
xnor U3105 (N_3105,N_2961,N_2400);
or U3106 (N_3106,N_2864,N_2567);
nand U3107 (N_3107,N_2289,N_2701);
and U3108 (N_3108,N_2949,N_2230);
and U3109 (N_3109,N_2308,N_2492);
nand U3110 (N_3110,N_2717,N_2249);
nor U3111 (N_3111,N_2071,N_2067);
xor U3112 (N_3112,N_2092,N_2398);
nand U3113 (N_3113,N_2966,N_2560);
xor U3114 (N_3114,N_2862,N_2848);
or U3115 (N_3115,N_2728,N_2513);
and U3116 (N_3116,N_2354,N_2804);
xor U3117 (N_3117,N_2944,N_2353);
nand U3118 (N_3118,N_2453,N_2272);
nor U3119 (N_3119,N_2777,N_2749);
xor U3120 (N_3120,N_2462,N_2534);
nor U3121 (N_3121,N_2609,N_2801);
nand U3122 (N_3122,N_2155,N_2904);
nor U3123 (N_3123,N_2812,N_2497);
nand U3124 (N_3124,N_2200,N_2032);
or U3125 (N_3125,N_2196,N_2482);
nand U3126 (N_3126,N_2193,N_2247);
nor U3127 (N_3127,N_2370,N_2255);
xnor U3128 (N_3128,N_2729,N_2388);
or U3129 (N_3129,N_2073,N_2851);
or U3130 (N_3130,N_2437,N_2956);
nand U3131 (N_3131,N_2931,N_2499);
nor U3132 (N_3132,N_2569,N_2743);
and U3133 (N_3133,N_2214,N_2527);
nor U3134 (N_3134,N_2457,N_2537);
nand U3135 (N_3135,N_2757,N_2509);
nor U3136 (N_3136,N_2325,N_2526);
and U3137 (N_3137,N_2191,N_2602);
nand U3138 (N_3138,N_2460,N_2041);
or U3139 (N_3139,N_2871,N_2923);
or U3140 (N_3140,N_2769,N_2580);
and U3141 (N_3141,N_2295,N_2798);
xor U3142 (N_3142,N_2745,N_2858);
or U3143 (N_3143,N_2822,N_2723);
xnor U3144 (N_3144,N_2047,N_2084);
nand U3145 (N_3145,N_2764,N_2831);
nor U3146 (N_3146,N_2620,N_2215);
or U3147 (N_3147,N_2576,N_2987);
or U3148 (N_3148,N_2202,N_2055);
xor U3149 (N_3149,N_2896,N_2838);
nand U3150 (N_3150,N_2078,N_2974);
and U3151 (N_3151,N_2528,N_2883);
or U3152 (N_3152,N_2052,N_2563);
nand U3153 (N_3153,N_2031,N_2472);
nand U3154 (N_3154,N_2185,N_2926);
xnor U3155 (N_3155,N_2465,N_2135);
nor U3156 (N_3156,N_2319,N_2708);
and U3157 (N_3157,N_2133,N_2881);
and U3158 (N_3158,N_2297,N_2106);
or U3159 (N_3159,N_2643,N_2429);
nand U3160 (N_3160,N_2597,N_2045);
nor U3161 (N_3161,N_2138,N_2044);
or U3162 (N_3162,N_2143,N_2113);
or U3163 (N_3163,N_2328,N_2184);
nor U3164 (N_3164,N_2394,N_2893);
and U3165 (N_3165,N_2373,N_2682);
or U3166 (N_3166,N_2674,N_2892);
nand U3167 (N_3167,N_2688,N_2324);
nor U3168 (N_3168,N_2814,N_2401);
nand U3169 (N_3169,N_2491,N_2173);
xor U3170 (N_3170,N_2973,N_2562);
nand U3171 (N_3171,N_2330,N_2810);
nor U3172 (N_3172,N_2877,N_2635);
or U3173 (N_3173,N_2194,N_2456);
xor U3174 (N_3174,N_2913,N_2186);
nor U3175 (N_3175,N_2641,N_2271);
or U3176 (N_3176,N_2590,N_2523);
and U3177 (N_3177,N_2090,N_2349);
xnor U3178 (N_3178,N_2257,N_2639);
xnor U3179 (N_3179,N_2699,N_2767);
and U3180 (N_3180,N_2262,N_2710);
and U3181 (N_3181,N_2162,N_2156);
or U3182 (N_3182,N_2946,N_2873);
nand U3183 (N_3183,N_2380,N_2132);
nor U3184 (N_3184,N_2254,N_2903);
and U3185 (N_3185,N_2142,N_2852);
nor U3186 (N_3186,N_2593,N_2754);
nor U3187 (N_3187,N_2035,N_2573);
or U3188 (N_3188,N_2420,N_2089);
or U3189 (N_3189,N_2107,N_2004);
or U3190 (N_3190,N_2784,N_2863);
nor U3191 (N_3191,N_2403,N_2612);
and U3192 (N_3192,N_2988,N_2781);
and U3193 (N_3193,N_2725,N_2454);
nor U3194 (N_3194,N_2564,N_2079);
or U3195 (N_3195,N_2461,N_2939);
nand U3196 (N_3196,N_2742,N_2650);
and U3197 (N_3197,N_2080,N_2549);
nand U3198 (N_3198,N_2875,N_2274);
nand U3199 (N_3199,N_2310,N_2821);
nor U3200 (N_3200,N_2521,N_2997);
nor U3201 (N_3201,N_2344,N_2950);
and U3202 (N_3202,N_2258,N_2458);
or U3203 (N_3203,N_2672,N_2619);
nand U3204 (N_3204,N_2357,N_2157);
or U3205 (N_3205,N_2086,N_2015);
nor U3206 (N_3206,N_2227,N_2763);
and U3207 (N_3207,N_2361,N_2007);
nand U3208 (N_3208,N_2516,N_2554);
nor U3209 (N_3209,N_2886,N_2150);
nor U3210 (N_3210,N_2799,N_2427);
nor U3211 (N_3211,N_2796,N_2405);
nand U3212 (N_3212,N_2195,N_2510);
or U3213 (N_3213,N_2835,N_2475);
or U3214 (N_3214,N_2568,N_2464);
or U3215 (N_3215,N_2843,N_2476);
or U3216 (N_3216,N_2626,N_2466);
nand U3217 (N_3217,N_2065,N_2938);
and U3218 (N_3218,N_2436,N_2498);
or U3219 (N_3219,N_2037,N_2489);
or U3220 (N_3220,N_2299,N_2187);
nand U3221 (N_3221,N_2937,N_2811);
nand U3222 (N_3222,N_2229,N_2243);
or U3223 (N_3223,N_2286,N_2889);
and U3224 (N_3224,N_2911,N_2496);
nor U3225 (N_3225,N_2446,N_2396);
and U3226 (N_3226,N_2140,N_2263);
nor U3227 (N_3227,N_2377,N_2208);
or U3228 (N_3228,N_2166,N_2141);
nand U3229 (N_3229,N_2218,N_2867);
and U3230 (N_3230,N_2604,N_2669);
nor U3231 (N_3231,N_2902,N_2321);
or U3232 (N_3232,N_2930,N_2188);
nand U3233 (N_3233,N_2085,N_2681);
and U3234 (N_3234,N_2820,N_2768);
or U3235 (N_3235,N_2118,N_2802);
nor U3236 (N_3236,N_2642,N_2175);
nand U3237 (N_3237,N_2139,N_2021);
or U3238 (N_3238,N_2833,N_2450);
or U3239 (N_3239,N_2137,N_2213);
nand U3240 (N_3240,N_2477,N_2292);
xor U3241 (N_3241,N_2652,N_2792);
xnor U3242 (N_3242,N_2093,N_2773);
xnor U3243 (N_3243,N_2712,N_2306);
xor U3244 (N_3244,N_2759,N_2019);
or U3245 (N_3245,N_2269,N_2376);
and U3246 (N_3246,N_2209,N_2265);
nand U3247 (N_3247,N_2755,N_2687);
nand U3248 (N_3248,N_2806,N_2183);
and U3249 (N_3249,N_2693,N_2288);
nor U3250 (N_3250,N_2947,N_2083);
and U3251 (N_3251,N_2248,N_2253);
nor U3252 (N_3252,N_2582,N_2036);
or U3253 (N_3253,N_2025,N_2958);
or U3254 (N_3254,N_2001,N_2900);
and U3255 (N_3255,N_2720,N_2898);
nor U3256 (N_3256,N_2678,N_2577);
nor U3257 (N_3257,N_2112,N_2739);
and U3258 (N_3258,N_2522,N_2661);
and U3259 (N_3259,N_2480,N_2705);
xor U3260 (N_3260,N_2023,N_2756);
nand U3261 (N_3261,N_2550,N_2177);
nand U3262 (N_3262,N_2212,N_2766);
nand U3263 (N_3263,N_2878,N_2100);
or U3264 (N_3264,N_2868,N_2002);
nand U3265 (N_3265,N_2935,N_2242);
or U3266 (N_3266,N_2063,N_2256);
nand U3267 (N_3267,N_2431,N_2392);
nand U3268 (N_3268,N_2121,N_2369);
nor U3269 (N_3269,N_2342,N_2925);
or U3270 (N_3270,N_2828,N_2654);
nand U3271 (N_3271,N_2432,N_2114);
and U3272 (N_3272,N_2481,N_2711);
nand U3273 (N_3273,N_2345,N_2668);
nor U3274 (N_3274,N_2832,N_2540);
or U3275 (N_3275,N_2979,N_2125);
or U3276 (N_3276,N_2505,N_2435);
and U3277 (N_3277,N_2646,N_2575);
nor U3278 (N_3278,N_2060,N_2365);
xnor U3279 (N_3279,N_2951,N_2116);
or U3280 (N_3280,N_2408,N_2653);
xor U3281 (N_3281,N_2058,N_2630);
nor U3282 (N_3282,N_2824,N_2444);
xnor U3283 (N_3283,N_2706,N_2309);
nor U3284 (N_3284,N_2252,N_2447);
or U3285 (N_3285,N_2134,N_2632);
xnor U3286 (N_3286,N_2105,N_2221);
and U3287 (N_3287,N_2360,N_2834);
nand U3288 (N_3288,N_2197,N_2216);
and U3289 (N_3289,N_2300,N_2771);
nand U3290 (N_3290,N_2542,N_2574);
nand U3291 (N_3291,N_2579,N_2916);
or U3292 (N_3292,N_2374,N_2751);
nor U3293 (N_3293,N_2733,N_2130);
nand U3294 (N_3294,N_2856,N_2685);
or U3295 (N_3295,N_2010,N_2167);
and U3296 (N_3296,N_2980,N_2259);
nor U3297 (N_3297,N_2484,N_2765);
xor U3298 (N_3298,N_2393,N_2428);
or U3299 (N_3299,N_2233,N_2556);
xor U3300 (N_3300,N_2240,N_2774);
or U3301 (N_3301,N_2595,N_2531);
nand U3302 (N_3302,N_2530,N_2992);
and U3303 (N_3303,N_2277,N_2866);
nand U3304 (N_3304,N_2355,N_2707);
or U3305 (N_3305,N_2737,N_2689);
or U3306 (N_3306,N_2989,N_2680);
nor U3307 (N_3307,N_2017,N_2119);
nor U3308 (N_3308,N_2634,N_2807);
xnor U3309 (N_3309,N_2888,N_2847);
nand U3310 (N_3310,N_2968,N_2627);
nor U3311 (N_3311,N_2455,N_2818);
nor U3312 (N_3312,N_2948,N_2976);
and U3313 (N_3313,N_2986,N_2599);
xor U3314 (N_3314,N_2236,N_2860);
nand U3315 (N_3315,N_2122,N_2164);
and U3316 (N_3316,N_2525,N_2356);
nor U3317 (N_3317,N_2149,N_2199);
nand U3318 (N_3318,N_2512,N_2181);
xnor U3319 (N_3319,N_2311,N_2776);
and U3320 (N_3320,N_2389,N_2518);
nor U3321 (N_3321,N_2205,N_2897);
and U3322 (N_3322,N_2161,N_2760);
nand U3323 (N_3323,N_2696,N_2547);
nor U3324 (N_3324,N_2601,N_2998);
nor U3325 (N_3325,N_2616,N_2869);
or U3326 (N_3326,N_2294,N_2964);
or U3327 (N_3327,N_2407,N_2304);
nand U3328 (N_3328,N_2117,N_2261);
or U3329 (N_3329,N_2656,N_2719);
nor U3330 (N_3330,N_2470,N_2631);
nor U3331 (N_3331,N_2876,N_2419);
nand U3332 (N_3332,N_2469,N_2536);
and U3333 (N_3333,N_2421,N_2673);
or U3334 (N_3334,N_2640,N_2425);
or U3335 (N_3335,N_2283,N_2734);
nand U3336 (N_3336,N_2770,N_2695);
and U3337 (N_3337,N_2368,N_2022);
or U3338 (N_3338,N_2266,N_2124);
nand U3339 (N_3339,N_2163,N_2638);
nand U3340 (N_3340,N_2762,N_2659);
and U3341 (N_3341,N_2329,N_2147);
nand U3342 (N_3342,N_2327,N_2731);
nand U3343 (N_3343,N_2219,N_2211);
and U3344 (N_3344,N_2535,N_2596);
and U3345 (N_3345,N_2908,N_2637);
nor U3346 (N_3346,N_2782,N_2657);
nand U3347 (N_3347,N_2861,N_2120);
xor U3348 (N_3348,N_2532,N_2857);
nand U3349 (N_3349,N_2703,N_2813);
nor U3350 (N_3350,N_2854,N_2910);
nand U3351 (N_3351,N_2290,N_2945);
nand U3352 (N_3352,N_2932,N_2189);
nor U3353 (N_3353,N_2381,N_2907);
nor U3354 (N_3354,N_2846,N_2478);
xnor U3355 (N_3355,N_2840,N_2251);
xor U3356 (N_3356,N_2459,N_2072);
or U3357 (N_3357,N_2244,N_2624);
and U3358 (N_3358,N_2203,N_2412);
nor U3359 (N_3359,N_2787,N_2352);
or U3360 (N_3360,N_2042,N_2409);
or U3361 (N_3361,N_2750,N_2051);
nand U3362 (N_3362,N_2028,N_2103);
nand U3363 (N_3363,N_2285,N_2003);
nor U3364 (N_3364,N_2087,N_2967);
nor U3365 (N_3365,N_2921,N_2246);
and U3366 (N_3366,N_2899,N_2207);
or U3367 (N_3367,N_2538,N_2493);
or U3368 (N_3368,N_2735,N_2829);
nand U3369 (N_3369,N_2006,N_2551);
and U3370 (N_3370,N_2508,N_2367);
nor U3371 (N_3371,N_2364,N_2471);
nor U3372 (N_3372,N_2111,N_2467);
and U3373 (N_3373,N_2607,N_2316);
or U3374 (N_3374,N_2332,N_2452);
and U3375 (N_3375,N_2993,N_2890);
and U3376 (N_3376,N_2533,N_2495);
and U3377 (N_3377,N_2740,N_2995);
nand U3378 (N_3378,N_2287,N_2982);
and U3379 (N_3379,N_2387,N_2486);
or U3380 (N_3380,N_2553,N_2109);
nor U3381 (N_3381,N_2442,N_2439);
and U3382 (N_3382,N_2176,N_2014);
or U3383 (N_3383,N_2614,N_2894);
nand U3384 (N_3384,N_2331,N_2790);
nor U3385 (N_3385,N_2991,N_2273);
nand U3386 (N_3386,N_2267,N_2104);
xor U3387 (N_3387,N_2054,N_2504);
xor U3388 (N_3388,N_2836,N_2069);
nand U3389 (N_3389,N_2451,N_2676);
nand U3390 (N_3390,N_2144,N_2600);
or U3391 (N_3391,N_2076,N_2692);
or U3392 (N_3392,N_2558,N_2108);
nor U3393 (N_3393,N_2340,N_2741);
nand U3394 (N_3394,N_2772,N_2445);
xnor U3395 (N_3395,N_2928,N_2074);
and U3396 (N_3396,N_2101,N_2667);
nand U3397 (N_3397,N_2552,N_2927);
nor U3398 (N_3398,N_2018,N_2917);
nand U3399 (N_3399,N_2206,N_2048);
or U3400 (N_3400,N_2426,N_2423);
xor U3401 (N_3401,N_2716,N_2348);
nor U3402 (N_3402,N_2983,N_2260);
and U3403 (N_3403,N_2334,N_2095);
and U3404 (N_3404,N_2088,N_2039);
and U3405 (N_3405,N_2307,N_2603);
or U3406 (N_3406,N_2020,N_2622);
nand U3407 (N_3407,N_2154,N_2915);
nand U3408 (N_3408,N_2160,N_2529);
or U3409 (N_3409,N_2589,N_2281);
and U3410 (N_3410,N_2789,N_2302);
or U3411 (N_3411,N_2912,N_2228);
and U3412 (N_3412,N_2226,N_2702);
or U3413 (N_3413,N_2326,N_2885);
or U3414 (N_3414,N_2358,N_2981);
nand U3415 (N_3415,N_2404,N_2957);
nor U3416 (N_3416,N_2313,N_2962);
nand U3417 (N_3417,N_2744,N_2386);
xnor U3418 (N_3418,N_2613,N_2169);
xnor U3419 (N_3419,N_2418,N_2746);
and U3420 (N_3420,N_2953,N_2837);
or U3421 (N_3421,N_2507,N_2794);
or U3422 (N_3422,N_2046,N_2520);
xor U3423 (N_3423,N_2999,N_2485);
xnor U3424 (N_3424,N_2443,N_2610);
and U3425 (N_3425,N_2077,N_2952);
nand U3426 (N_3426,N_2972,N_2954);
nand U3427 (N_3427,N_2615,N_2098);
or U3428 (N_3428,N_2919,N_2148);
and U3429 (N_3429,N_2704,N_2034);
nor U3430 (N_3430,N_2977,N_2192);
nand U3431 (N_3431,N_2153,N_2384);
and U3432 (N_3432,N_2146,N_2996);
nor U3433 (N_3433,N_2817,N_2815);
nor U3434 (N_3434,N_2665,N_2606);
and U3435 (N_3435,N_2250,N_2190);
or U3436 (N_3436,N_2940,N_2438);
nor U3437 (N_3437,N_2320,N_2301);
nor U3438 (N_3438,N_2280,N_2514);
or U3439 (N_3439,N_2033,N_2559);
xnor U3440 (N_3440,N_2666,N_2341);
nand U3441 (N_3441,N_2721,N_2859);
nor U3442 (N_3442,N_2960,N_2855);
or U3443 (N_3443,N_2588,N_2963);
and U3444 (N_3444,N_2371,N_2546);
or U3445 (N_3445,N_2990,N_2448);
nand U3446 (N_3446,N_2726,N_2758);
xor U3447 (N_3447,N_2557,N_2548);
nand U3448 (N_3448,N_2397,N_2385);
or U3449 (N_3449,N_2008,N_2378);
or U3450 (N_3450,N_2694,N_2027);
nand U3451 (N_3451,N_2102,N_2519);
and U3452 (N_3452,N_2346,N_2449);
and U3453 (N_3453,N_2683,N_2738);
nand U3454 (N_3454,N_2775,N_2633);
nor U3455 (N_3455,N_2059,N_2220);
nor U3456 (N_3456,N_2096,N_2592);
nor U3457 (N_3457,N_2924,N_2918);
nand U3458 (N_3458,N_2210,N_2545);
and U3459 (N_3459,N_2198,N_2382);
and U3460 (N_3460,N_2315,N_2517);
nor U3461 (N_3461,N_2275,N_2234);
xnor U3462 (N_3462,N_2366,N_2223);
or U3463 (N_3463,N_2168,N_2239);
and U3464 (N_3464,N_2323,N_2050);
and U3465 (N_3465,N_2943,N_2152);
nand U3466 (N_3466,N_2217,N_2684);
or U3467 (N_3467,N_2016,N_2727);
nand U3468 (N_3468,N_2131,N_2816);
xnor U3469 (N_3469,N_2129,N_2151);
nor U3470 (N_3470,N_2809,N_2941);
and U3471 (N_3471,N_2853,N_2178);
nor U3472 (N_3472,N_2649,N_2825);
or U3473 (N_3473,N_2375,N_2165);
and U3474 (N_3474,N_2070,N_2651);
nand U3475 (N_3475,N_2906,N_2511);
and U3476 (N_3476,N_2123,N_2827);
nand U3477 (N_3477,N_2170,N_2075);
nor U3478 (N_3478,N_2204,N_2984);
nand U3479 (N_3479,N_2182,N_2099);
nor U3480 (N_3480,N_2434,N_2180);
nor U3481 (N_3481,N_2718,N_2312);
and U3482 (N_3482,N_2714,N_2338);
nor U3483 (N_3483,N_2066,N_2040);
nor U3484 (N_3484,N_2399,N_2826);
or U3485 (N_3485,N_2128,N_2879);
and U3486 (N_3486,N_2778,N_2660);
nand U3487 (N_3487,N_2068,N_2611);
and U3488 (N_3488,N_2697,N_2402);
or U3489 (N_3489,N_2383,N_2061);
or U3490 (N_3490,N_2645,N_2591);
or U3491 (N_3491,N_2091,N_2805);
nand U3492 (N_3492,N_2539,N_2581);
nor U3493 (N_3493,N_2433,N_2623);
nand U3494 (N_3494,N_2594,N_2487);
nor U3495 (N_3495,N_2413,N_2670);
nor U3496 (N_3496,N_2473,N_2440);
nand U3497 (N_3497,N_2541,N_2333);
nand U3498 (N_3498,N_2647,N_2005);
nor U3499 (N_3499,N_2395,N_2994);
xnor U3500 (N_3500,N_2296,N_2885);
nor U3501 (N_3501,N_2992,N_2002);
and U3502 (N_3502,N_2744,N_2190);
nand U3503 (N_3503,N_2979,N_2444);
nor U3504 (N_3504,N_2840,N_2669);
and U3505 (N_3505,N_2159,N_2528);
and U3506 (N_3506,N_2001,N_2953);
and U3507 (N_3507,N_2773,N_2535);
or U3508 (N_3508,N_2577,N_2995);
and U3509 (N_3509,N_2529,N_2337);
nor U3510 (N_3510,N_2971,N_2443);
or U3511 (N_3511,N_2545,N_2421);
and U3512 (N_3512,N_2448,N_2243);
nor U3513 (N_3513,N_2483,N_2015);
and U3514 (N_3514,N_2794,N_2431);
nor U3515 (N_3515,N_2677,N_2068);
or U3516 (N_3516,N_2923,N_2383);
nand U3517 (N_3517,N_2950,N_2049);
or U3518 (N_3518,N_2796,N_2113);
nand U3519 (N_3519,N_2966,N_2910);
xor U3520 (N_3520,N_2820,N_2040);
or U3521 (N_3521,N_2612,N_2175);
or U3522 (N_3522,N_2749,N_2696);
or U3523 (N_3523,N_2367,N_2739);
and U3524 (N_3524,N_2112,N_2717);
or U3525 (N_3525,N_2419,N_2637);
nand U3526 (N_3526,N_2885,N_2759);
nand U3527 (N_3527,N_2753,N_2500);
xor U3528 (N_3528,N_2550,N_2996);
or U3529 (N_3529,N_2289,N_2601);
nand U3530 (N_3530,N_2465,N_2576);
and U3531 (N_3531,N_2765,N_2820);
nand U3532 (N_3532,N_2052,N_2311);
xnor U3533 (N_3533,N_2758,N_2544);
nor U3534 (N_3534,N_2236,N_2064);
nor U3535 (N_3535,N_2594,N_2641);
and U3536 (N_3536,N_2366,N_2750);
and U3537 (N_3537,N_2233,N_2473);
xnor U3538 (N_3538,N_2583,N_2517);
nor U3539 (N_3539,N_2318,N_2028);
or U3540 (N_3540,N_2608,N_2856);
nand U3541 (N_3541,N_2898,N_2439);
nand U3542 (N_3542,N_2704,N_2422);
nand U3543 (N_3543,N_2588,N_2219);
nor U3544 (N_3544,N_2983,N_2862);
nand U3545 (N_3545,N_2142,N_2002);
nor U3546 (N_3546,N_2948,N_2496);
nor U3547 (N_3547,N_2664,N_2337);
nor U3548 (N_3548,N_2831,N_2203);
nor U3549 (N_3549,N_2054,N_2753);
xor U3550 (N_3550,N_2090,N_2763);
nor U3551 (N_3551,N_2889,N_2181);
nor U3552 (N_3552,N_2908,N_2811);
xor U3553 (N_3553,N_2985,N_2634);
or U3554 (N_3554,N_2252,N_2653);
or U3555 (N_3555,N_2154,N_2202);
xnor U3556 (N_3556,N_2454,N_2697);
nor U3557 (N_3557,N_2282,N_2192);
nand U3558 (N_3558,N_2066,N_2195);
nand U3559 (N_3559,N_2534,N_2153);
or U3560 (N_3560,N_2937,N_2026);
and U3561 (N_3561,N_2177,N_2555);
nor U3562 (N_3562,N_2817,N_2630);
nand U3563 (N_3563,N_2418,N_2554);
or U3564 (N_3564,N_2929,N_2983);
nand U3565 (N_3565,N_2459,N_2431);
nor U3566 (N_3566,N_2788,N_2748);
nor U3567 (N_3567,N_2687,N_2603);
nor U3568 (N_3568,N_2467,N_2633);
nor U3569 (N_3569,N_2668,N_2238);
and U3570 (N_3570,N_2782,N_2358);
nor U3571 (N_3571,N_2130,N_2272);
and U3572 (N_3572,N_2105,N_2592);
nor U3573 (N_3573,N_2140,N_2104);
and U3574 (N_3574,N_2085,N_2239);
nor U3575 (N_3575,N_2289,N_2641);
nor U3576 (N_3576,N_2992,N_2142);
nor U3577 (N_3577,N_2316,N_2541);
and U3578 (N_3578,N_2935,N_2772);
nand U3579 (N_3579,N_2792,N_2137);
or U3580 (N_3580,N_2865,N_2550);
nor U3581 (N_3581,N_2267,N_2439);
nor U3582 (N_3582,N_2298,N_2156);
nand U3583 (N_3583,N_2098,N_2304);
or U3584 (N_3584,N_2327,N_2567);
nor U3585 (N_3585,N_2885,N_2365);
xor U3586 (N_3586,N_2174,N_2995);
or U3587 (N_3587,N_2927,N_2829);
nand U3588 (N_3588,N_2126,N_2198);
xnor U3589 (N_3589,N_2259,N_2093);
nand U3590 (N_3590,N_2783,N_2159);
nor U3591 (N_3591,N_2271,N_2686);
nand U3592 (N_3592,N_2060,N_2711);
nand U3593 (N_3593,N_2682,N_2203);
nand U3594 (N_3594,N_2758,N_2872);
or U3595 (N_3595,N_2906,N_2093);
nand U3596 (N_3596,N_2568,N_2093);
xnor U3597 (N_3597,N_2547,N_2458);
xnor U3598 (N_3598,N_2945,N_2889);
nand U3599 (N_3599,N_2399,N_2014);
nor U3600 (N_3600,N_2763,N_2253);
or U3601 (N_3601,N_2125,N_2623);
nand U3602 (N_3602,N_2743,N_2813);
nand U3603 (N_3603,N_2912,N_2352);
and U3604 (N_3604,N_2329,N_2093);
nand U3605 (N_3605,N_2289,N_2580);
or U3606 (N_3606,N_2375,N_2700);
or U3607 (N_3607,N_2949,N_2601);
and U3608 (N_3608,N_2471,N_2745);
or U3609 (N_3609,N_2953,N_2636);
nor U3610 (N_3610,N_2549,N_2708);
and U3611 (N_3611,N_2655,N_2862);
or U3612 (N_3612,N_2668,N_2078);
nor U3613 (N_3613,N_2331,N_2586);
nand U3614 (N_3614,N_2630,N_2903);
or U3615 (N_3615,N_2258,N_2372);
and U3616 (N_3616,N_2307,N_2873);
and U3617 (N_3617,N_2831,N_2955);
or U3618 (N_3618,N_2169,N_2358);
or U3619 (N_3619,N_2569,N_2963);
or U3620 (N_3620,N_2920,N_2278);
xor U3621 (N_3621,N_2511,N_2503);
nand U3622 (N_3622,N_2868,N_2048);
nor U3623 (N_3623,N_2552,N_2939);
xor U3624 (N_3624,N_2831,N_2972);
or U3625 (N_3625,N_2593,N_2690);
nor U3626 (N_3626,N_2524,N_2850);
nor U3627 (N_3627,N_2416,N_2869);
and U3628 (N_3628,N_2010,N_2309);
nor U3629 (N_3629,N_2631,N_2578);
xnor U3630 (N_3630,N_2698,N_2929);
and U3631 (N_3631,N_2513,N_2626);
nand U3632 (N_3632,N_2834,N_2638);
or U3633 (N_3633,N_2247,N_2291);
and U3634 (N_3634,N_2537,N_2439);
or U3635 (N_3635,N_2368,N_2505);
nand U3636 (N_3636,N_2672,N_2282);
nand U3637 (N_3637,N_2350,N_2155);
nand U3638 (N_3638,N_2057,N_2059);
or U3639 (N_3639,N_2030,N_2757);
nor U3640 (N_3640,N_2013,N_2894);
nand U3641 (N_3641,N_2686,N_2937);
nand U3642 (N_3642,N_2165,N_2547);
nand U3643 (N_3643,N_2400,N_2740);
nand U3644 (N_3644,N_2629,N_2783);
or U3645 (N_3645,N_2721,N_2436);
nor U3646 (N_3646,N_2292,N_2834);
nor U3647 (N_3647,N_2554,N_2527);
nand U3648 (N_3648,N_2947,N_2817);
nor U3649 (N_3649,N_2567,N_2694);
or U3650 (N_3650,N_2637,N_2399);
nand U3651 (N_3651,N_2614,N_2170);
nand U3652 (N_3652,N_2732,N_2485);
xor U3653 (N_3653,N_2980,N_2856);
or U3654 (N_3654,N_2129,N_2810);
or U3655 (N_3655,N_2229,N_2320);
and U3656 (N_3656,N_2667,N_2954);
nand U3657 (N_3657,N_2109,N_2718);
or U3658 (N_3658,N_2643,N_2418);
and U3659 (N_3659,N_2853,N_2418);
nor U3660 (N_3660,N_2414,N_2945);
nor U3661 (N_3661,N_2341,N_2927);
xnor U3662 (N_3662,N_2391,N_2669);
xor U3663 (N_3663,N_2791,N_2782);
or U3664 (N_3664,N_2016,N_2160);
nand U3665 (N_3665,N_2814,N_2558);
nor U3666 (N_3666,N_2222,N_2959);
and U3667 (N_3667,N_2194,N_2563);
and U3668 (N_3668,N_2837,N_2133);
or U3669 (N_3669,N_2588,N_2477);
or U3670 (N_3670,N_2637,N_2901);
or U3671 (N_3671,N_2149,N_2890);
nand U3672 (N_3672,N_2010,N_2477);
nor U3673 (N_3673,N_2424,N_2707);
xnor U3674 (N_3674,N_2342,N_2417);
or U3675 (N_3675,N_2324,N_2050);
and U3676 (N_3676,N_2983,N_2028);
and U3677 (N_3677,N_2165,N_2426);
nand U3678 (N_3678,N_2087,N_2486);
or U3679 (N_3679,N_2523,N_2053);
and U3680 (N_3680,N_2898,N_2209);
and U3681 (N_3681,N_2411,N_2195);
and U3682 (N_3682,N_2437,N_2568);
nor U3683 (N_3683,N_2230,N_2929);
and U3684 (N_3684,N_2474,N_2006);
or U3685 (N_3685,N_2974,N_2060);
nand U3686 (N_3686,N_2273,N_2206);
xor U3687 (N_3687,N_2517,N_2680);
nor U3688 (N_3688,N_2516,N_2482);
nor U3689 (N_3689,N_2959,N_2954);
nand U3690 (N_3690,N_2711,N_2367);
nor U3691 (N_3691,N_2958,N_2614);
nand U3692 (N_3692,N_2794,N_2818);
nand U3693 (N_3693,N_2694,N_2713);
nor U3694 (N_3694,N_2703,N_2721);
nor U3695 (N_3695,N_2520,N_2925);
and U3696 (N_3696,N_2107,N_2846);
nor U3697 (N_3697,N_2762,N_2252);
or U3698 (N_3698,N_2169,N_2579);
or U3699 (N_3699,N_2025,N_2691);
or U3700 (N_3700,N_2073,N_2695);
nor U3701 (N_3701,N_2031,N_2102);
and U3702 (N_3702,N_2352,N_2817);
nor U3703 (N_3703,N_2487,N_2079);
or U3704 (N_3704,N_2028,N_2991);
nor U3705 (N_3705,N_2389,N_2790);
nand U3706 (N_3706,N_2575,N_2532);
nor U3707 (N_3707,N_2883,N_2155);
or U3708 (N_3708,N_2491,N_2920);
or U3709 (N_3709,N_2241,N_2368);
nor U3710 (N_3710,N_2078,N_2175);
or U3711 (N_3711,N_2529,N_2714);
and U3712 (N_3712,N_2958,N_2070);
nand U3713 (N_3713,N_2843,N_2401);
or U3714 (N_3714,N_2054,N_2849);
or U3715 (N_3715,N_2204,N_2221);
or U3716 (N_3716,N_2467,N_2203);
or U3717 (N_3717,N_2588,N_2364);
or U3718 (N_3718,N_2723,N_2909);
xor U3719 (N_3719,N_2913,N_2826);
and U3720 (N_3720,N_2944,N_2780);
nor U3721 (N_3721,N_2788,N_2842);
nor U3722 (N_3722,N_2635,N_2227);
or U3723 (N_3723,N_2689,N_2630);
and U3724 (N_3724,N_2648,N_2404);
nand U3725 (N_3725,N_2343,N_2846);
nor U3726 (N_3726,N_2757,N_2500);
or U3727 (N_3727,N_2516,N_2021);
nor U3728 (N_3728,N_2586,N_2637);
nor U3729 (N_3729,N_2258,N_2414);
and U3730 (N_3730,N_2488,N_2104);
or U3731 (N_3731,N_2862,N_2354);
or U3732 (N_3732,N_2152,N_2600);
nand U3733 (N_3733,N_2076,N_2633);
nand U3734 (N_3734,N_2740,N_2847);
or U3735 (N_3735,N_2765,N_2016);
xnor U3736 (N_3736,N_2974,N_2977);
or U3737 (N_3737,N_2251,N_2254);
or U3738 (N_3738,N_2333,N_2059);
and U3739 (N_3739,N_2422,N_2674);
and U3740 (N_3740,N_2252,N_2164);
and U3741 (N_3741,N_2255,N_2307);
nor U3742 (N_3742,N_2947,N_2427);
and U3743 (N_3743,N_2388,N_2980);
or U3744 (N_3744,N_2617,N_2636);
nor U3745 (N_3745,N_2038,N_2042);
and U3746 (N_3746,N_2874,N_2542);
and U3747 (N_3747,N_2872,N_2975);
nand U3748 (N_3748,N_2568,N_2551);
and U3749 (N_3749,N_2439,N_2355);
or U3750 (N_3750,N_2219,N_2428);
and U3751 (N_3751,N_2070,N_2110);
and U3752 (N_3752,N_2805,N_2034);
or U3753 (N_3753,N_2878,N_2371);
xor U3754 (N_3754,N_2668,N_2913);
or U3755 (N_3755,N_2888,N_2504);
or U3756 (N_3756,N_2277,N_2126);
or U3757 (N_3757,N_2070,N_2229);
or U3758 (N_3758,N_2943,N_2742);
or U3759 (N_3759,N_2858,N_2097);
nand U3760 (N_3760,N_2291,N_2127);
and U3761 (N_3761,N_2594,N_2178);
or U3762 (N_3762,N_2903,N_2045);
or U3763 (N_3763,N_2516,N_2594);
nor U3764 (N_3764,N_2022,N_2475);
or U3765 (N_3765,N_2840,N_2458);
nand U3766 (N_3766,N_2695,N_2653);
and U3767 (N_3767,N_2139,N_2286);
or U3768 (N_3768,N_2494,N_2806);
or U3769 (N_3769,N_2582,N_2880);
nand U3770 (N_3770,N_2819,N_2160);
or U3771 (N_3771,N_2477,N_2830);
or U3772 (N_3772,N_2310,N_2127);
nor U3773 (N_3773,N_2328,N_2074);
or U3774 (N_3774,N_2618,N_2684);
or U3775 (N_3775,N_2884,N_2075);
nor U3776 (N_3776,N_2188,N_2550);
nand U3777 (N_3777,N_2184,N_2537);
or U3778 (N_3778,N_2893,N_2261);
and U3779 (N_3779,N_2375,N_2763);
and U3780 (N_3780,N_2567,N_2449);
and U3781 (N_3781,N_2364,N_2425);
xnor U3782 (N_3782,N_2706,N_2525);
or U3783 (N_3783,N_2480,N_2291);
nand U3784 (N_3784,N_2783,N_2582);
nor U3785 (N_3785,N_2179,N_2149);
and U3786 (N_3786,N_2570,N_2449);
nand U3787 (N_3787,N_2699,N_2163);
and U3788 (N_3788,N_2138,N_2039);
nand U3789 (N_3789,N_2141,N_2535);
xor U3790 (N_3790,N_2568,N_2972);
nor U3791 (N_3791,N_2594,N_2441);
nand U3792 (N_3792,N_2465,N_2261);
or U3793 (N_3793,N_2023,N_2982);
xor U3794 (N_3794,N_2040,N_2705);
and U3795 (N_3795,N_2659,N_2105);
nand U3796 (N_3796,N_2248,N_2271);
or U3797 (N_3797,N_2357,N_2949);
nand U3798 (N_3798,N_2520,N_2780);
and U3799 (N_3799,N_2031,N_2022);
and U3800 (N_3800,N_2024,N_2663);
nand U3801 (N_3801,N_2558,N_2977);
and U3802 (N_3802,N_2183,N_2926);
nor U3803 (N_3803,N_2754,N_2356);
nor U3804 (N_3804,N_2295,N_2589);
nor U3805 (N_3805,N_2953,N_2593);
nand U3806 (N_3806,N_2255,N_2144);
or U3807 (N_3807,N_2779,N_2285);
nand U3808 (N_3808,N_2796,N_2523);
xor U3809 (N_3809,N_2054,N_2023);
or U3810 (N_3810,N_2070,N_2930);
nor U3811 (N_3811,N_2593,N_2583);
nor U3812 (N_3812,N_2050,N_2722);
nand U3813 (N_3813,N_2107,N_2461);
nor U3814 (N_3814,N_2792,N_2072);
and U3815 (N_3815,N_2327,N_2103);
nor U3816 (N_3816,N_2030,N_2801);
and U3817 (N_3817,N_2453,N_2422);
and U3818 (N_3818,N_2452,N_2241);
or U3819 (N_3819,N_2122,N_2894);
or U3820 (N_3820,N_2675,N_2423);
nand U3821 (N_3821,N_2334,N_2518);
nor U3822 (N_3822,N_2170,N_2508);
nor U3823 (N_3823,N_2969,N_2333);
and U3824 (N_3824,N_2764,N_2862);
or U3825 (N_3825,N_2604,N_2639);
and U3826 (N_3826,N_2226,N_2280);
nand U3827 (N_3827,N_2834,N_2058);
nor U3828 (N_3828,N_2300,N_2374);
xor U3829 (N_3829,N_2339,N_2699);
xor U3830 (N_3830,N_2006,N_2069);
xnor U3831 (N_3831,N_2681,N_2295);
and U3832 (N_3832,N_2821,N_2121);
or U3833 (N_3833,N_2155,N_2191);
and U3834 (N_3834,N_2244,N_2701);
or U3835 (N_3835,N_2245,N_2561);
nor U3836 (N_3836,N_2006,N_2550);
nand U3837 (N_3837,N_2835,N_2576);
or U3838 (N_3838,N_2350,N_2952);
and U3839 (N_3839,N_2742,N_2809);
nand U3840 (N_3840,N_2728,N_2262);
nor U3841 (N_3841,N_2913,N_2614);
and U3842 (N_3842,N_2423,N_2966);
or U3843 (N_3843,N_2791,N_2559);
and U3844 (N_3844,N_2115,N_2635);
nand U3845 (N_3845,N_2330,N_2319);
and U3846 (N_3846,N_2778,N_2084);
nand U3847 (N_3847,N_2889,N_2763);
nand U3848 (N_3848,N_2157,N_2817);
nand U3849 (N_3849,N_2292,N_2379);
and U3850 (N_3850,N_2986,N_2501);
nand U3851 (N_3851,N_2035,N_2013);
or U3852 (N_3852,N_2138,N_2868);
nor U3853 (N_3853,N_2189,N_2084);
nand U3854 (N_3854,N_2223,N_2433);
and U3855 (N_3855,N_2994,N_2747);
nor U3856 (N_3856,N_2635,N_2302);
and U3857 (N_3857,N_2747,N_2119);
nand U3858 (N_3858,N_2088,N_2473);
or U3859 (N_3859,N_2565,N_2826);
and U3860 (N_3860,N_2687,N_2214);
or U3861 (N_3861,N_2748,N_2506);
nand U3862 (N_3862,N_2922,N_2834);
nand U3863 (N_3863,N_2884,N_2649);
xnor U3864 (N_3864,N_2953,N_2150);
or U3865 (N_3865,N_2691,N_2288);
or U3866 (N_3866,N_2804,N_2556);
nand U3867 (N_3867,N_2212,N_2788);
nand U3868 (N_3868,N_2607,N_2651);
and U3869 (N_3869,N_2353,N_2589);
nand U3870 (N_3870,N_2504,N_2093);
xor U3871 (N_3871,N_2402,N_2061);
nand U3872 (N_3872,N_2298,N_2536);
nand U3873 (N_3873,N_2476,N_2977);
and U3874 (N_3874,N_2346,N_2556);
nor U3875 (N_3875,N_2521,N_2045);
or U3876 (N_3876,N_2639,N_2415);
nor U3877 (N_3877,N_2592,N_2495);
nand U3878 (N_3878,N_2600,N_2374);
or U3879 (N_3879,N_2243,N_2954);
nand U3880 (N_3880,N_2401,N_2658);
nand U3881 (N_3881,N_2299,N_2981);
nor U3882 (N_3882,N_2792,N_2533);
or U3883 (N_3883,N_2212,N_2871);
or U3884 (N_3884,N_2427,N_2591);
or U3885 (N_3885,N_2869,N_2176);
or U3886 (N_3886,N_2249,N_2369);
nor U3887 (N_3887,N_2504,N_2995);
nand U3888 (N_3888,N_2330,N_2301);
nor U3889 (N_3889,N_2690,N_2054);
xnor U3890 (N_3890,N_2158,N_2688);
or U3891 (N_3891,N_2937,N_2050);
xnor U3892 (N_3892,N_2373,N_2760);
or U3893 (N_3893,N_2659,N_2327);
and U3894 (N_3894,N_2925,N_2109);
or U3895 (N_3895,N_2867,N_2632);
nand U3896 (N_3896,N_2488,N_2610);
nor U3897 (N_3897,N_2634,N_2393);
nor U3898 (N_3898,N_2614,N_2598);
or U3899 (N_3899,N_2480,N_2698);
nand U3900 (N_3900,N_2210,N_2387);
nand U3901 (N_3901,N_2975,N_2706);
and U3902 (N_3902,N_2716,N_2811);
nand U3903 (N_3903,N_2987,N_2147);
and U3904 (N_3904,N_2837,N_2582);
nor U3905 (N_3905,N_2191,N_2340);
and U3906 (N_3906,N_2371,N_2574);
nor U3907 (N_3907,N_2656,N_2709);
or U3908 (N_3908,N_2015,N_2295);
nor U3909 (N_3909,N_2656,N_2078);
xnor U3910 (N_3910,N_2352,N_2348);
nand U3911 (N_3911,N_2794,N_2714);
nor U3912 (N_3912,N_2466,N_2160);
nand U3913 (N_3913,N_2436,N_2101);
xnor U3914 (N_3914,N_2720,N_2712);
nand U3915 (N_3915,N_2082,N_2066);
nand U3916 (N_3916,N_2153,N_2566);
and U3917 (N_3917,N_2931,N_2956);
and U3918 (N_3918,N_2592,N_2987);
nand U3919 (N_3919,N_2794,N_2370);
and U3920 (N_3920,N_2772,N_2807);
and U3921 (N_3921,N_2125,N_2736);
nor U3922 (N_3922,N_2313,N_2343);
nor U3923 (N_3923,N_2222,N_2472);
nor U3924 (N_3924,N_2169,N_2173);
nand U3925 (N_3925,N_2326,N_2353);
nand U3926 (N_3926,N_2821,N_2896);
and U3927 (N_3927,N_2884,N_2549);
xnor U3928 (N_3928,N_2906,N_2439);
xor U3929 (N_3929,N_2026,N_2199);
or U3930 (N_3930,N_2196,N_2057);
xor U3931 (N_3931,N_2344,N_2787);
and U3932 (N_3932,N_2795,N_2562);
nand U3933 (N_3933,N_2278,N_2519);
and U3934 (N_3934,N_2238,N_2747);
and U3935 (N_3935,N_2558,N_2969);
xnor U3936 (N_3936,N_2588,N_2570);
or U3937 (N_3937,N_2623,N_2732);
nor U3938 (N_3938,N_2583,N_2666);
and U3939 (N_3939,N_2625,N_2932);
and U3940 (N_3940,N_2510,N_2820);
and U3941 (N_3941,N_2933,N_2817);
or U3942 (N_3942,N_2486,N_2470);
and U3943 (N_3943,N_2602,N_2021);
nand U3944 (N_3944,N_2681,N_2955);
nand U3945 (N_3945,N_2737,N_2936);
nand U3946 (N_3946,N_2254,N_2195);
or U3947 (N_3947,N_2146,N_2302);
nand U3948 (N_3948,N_2557,N_2753);
or U3949 (N_3949,N_2920,N_2147);
nand U3950 (N_3950,N_2404,N_2289);
or U3951 (N_3951,N_2039,N_2056);
nor U3952 (N_3952,N_2699,N_2635);
nor U3953 (N_3953,N_2475,N_2458);
nor U3954 (N_3954,N_2595,N_2855);
nand U3955 (N_3955,N_2312,N_2058);
xor U3956 (N_3956,N_2264,N_2930);
xnor U3957 (N_3957,N_2050,N_2198);
nor U3958 (N_3958,N_2843,N_2180);
nor U3959 (N_3959,N_2677,N_2327);
or U3960 (N_3960,N_2302,N_2958);
nor U3961 (N_3961,N_2879,N_2860);
and U3962 (N_3962,N_2534,N_2592);
xnor U3963 (N_3963,N_2276,N_2256);
nor U3964 (N_3964,N_2021,N_2647);
nor U3965 (N_3965,N_2708,N_2031);
or U3966 (N_3966,N_2278,N_2477);
nor U3967 (N_3967,N_2035,N_2505);
nand U3968 (N_3968,N_2501,N_2131);
or U3969 (N_3969,N_2864,N_2108);
or U3970 (N_3970,N_2627,N_2644);
nand U3971 (N_3971,N_2727,N_2463);
xnor U3972 (N_3972,N_2336,N_2284);
nor U3973 (N_3973,N_2759,N_2527);
nor U3974 (N_3974,N_2998,N_2789);
or U3975 (N_3975,N_2423,N_2121);
or U3976 (N_3976,N_2652,N_2504);
and U3977 (N_3977,N_2774,N_2970);
xnor U3978 (N_3978,N_2581,N_2309);
or U3979 (N_3979,N_2643,N_2754);
nand U3980 (N_3980,N_2469,N_2453);
xor U3981 (N_3981,N_2822,N_2864);
xnor U3982 (N_3982,N_2132,N_2416);
or U3983 (N_3983,N_2549,N_2105);
xnor U3984 (N_3984,N_2158,N_2183);
nor U3985 (N_3985,N_2908,N_2456);
nand U3986 (N_3986,N_2947,N_2994);
nand U3987 (N_3987,N_2901,N_2432);
xor U3988 (N_3988,N_2548,N_2332);
nand U3989 (N_3989,N_2620,N_2427);
nand U3990 (N_3990,N_2677,N_2169);
and U3991 (N_3991,N_2397,N_2187);
and U3992 (N_3992,N_2498,N_2635);
and U3993 (N_3993,N_2552,N_2185);
and U3994 (N_3994,N_2601,N_2389);
and U3995 (N_3995,N_2146,N_2637);
nor U3996 (N_3996,N_2563,N_2839);
nor U3997 (N_3997,N_2445,N_2966);
and U3998 (N_3998,N_2311,N_2081);
nor U3999 (N_3999,N_2610,N_2663);
xnor U4000 (N_4000,N_3870,N_3448);
nor U4001 (N_4001,N_3468,N_3917);
nor U4002 (N_4002,N_3280,N_3384);
and U4003 (N_4003,N_3197,N_3725);
or U4004 (N_4004,N_3054,N_3415);
nor U4005 (N_4005,N_3406,N_3854);
nand U4006 (N_4006,N_3596,N_3571);
xor U4007 (N_4007,N_3199,N_3402);
nor U4008 (N_4008,N_3196,N_3212);
nand U4009 (N_4009,N_3033,N_3648);
or U4010 (N_4010,N_3646,N_3497);
nand U4011 (N_4011,N_3600,N_3387);
nand U4012 (N_4012,N_3179,N_3128);
nor U4013 (N_4013,N_3061,N_3136);
or U4014 (N_4014,N_3954,N_3473);
nor U4015 (N_4015,N_3877,N_3352);
nor U4016 (N_4016,N_3987,N_3676);
and U4017 (N_4017,N_3368,N_3325);
and U4018 (N_4018,N_3577,N_3157);
or U4019 (N_4019,N_3747,N_3006);
and U4020 (N_4020,N_3193,N_3720);
or U4021 (N_4021,N_3728,N_3811);
and U4022 (N_4022,N_3994,N_3546);
nor U4023 (N_4023,N_3618,N_3267);
or U4024 (N_4024,N_3372,N_3268);
nor U4025 (N_4025,N_3550,N_3132);
nand U4026 (N_4026,N_3135,N_3871);
and U4027 (N_4027,N_3866,N_3506);
nand U4028 (N_4028,N_3974,N_3669);
and U4029 (N_4029,N_3141,N_3575);
nor U4030 (N_4030,N_3278,N_3553);
or U4031 (N_4031,N_3013,N_3951);
nand U4032 (N_4032,N_3508,N_3859);
and U4033 (N_4033,N_3805,N_3122);
nand U4034 (N_4034,N_3181,N_3828);
nand U4035 (N_4035,N_3922,N_3228);
or U4036 (N_4036,N_3538,N_3541);
nor U4037 (N_4037,N_3925,N_3860);
nand U4038 (N_4038,N_3029,N_3028);
or U4039 (N_4039,N_3200,N_3785);
nor U4040 (N_4040,N_3602,N_3024);
and U4041 (N_4041,N_3915,N_3856);
and U4042 (N_4042,N_3957,N_3800);
nand U4043 (N_4043,N_3053,N_3313);
or U4044 (N_4044,N_3680,N_3023);
nor U4045 (N_4045,N_3751,N_3099);
or U4046 (N_4046,N_3074,N_3520);
xor U4047 (N_4047,N_3684,N_3430);
or U4048 (N_4048,N_3231,N_3766);
and U4049 (N_4049,N_3270,N_3153);
and U4050 (N_4050,N_3757,N_3797);
nor U4051 (N_4051,N_3302,N_3044);
and U4052 (N_4052,N_3039,N_3235);
xor U4053 (N_4053,N_3381,N_3007);
nand U4054 (N_4054,N_3320,N_3882);
or U4055 (N_4055,N_3396,N_3894);
nand U4056 (N_4056,N_3752,N_3753);
and U4057 (N_4057,N_3000,N_3607);
nand U4058 (N_4058,N_3830,N_3485);
nor U4059 (N_4059,N_3932,N_3590);
nand U4060 (N_4060,N_3187,N_3282);
nor U4061 (N_4061,N_3813,N_3218);
or U4062 (N_4062,N_3317,N_3453);
nor U4063 (N_4063,N_3512,N_3429);
and U4064 (N_4064,N_3247,N_3134);
nand U4065 (N_4065,N_3662,N_3846);
or U4066 (N_4066,N_3471,N_3149);
nand U4067 (N_4067,N_3502,N_3695);
or U4068 (N_4068,N_3616,N_3563);
nor U4069 (N_4069,N_3927,N_3089);
or U4070 (N_4070,N_3166,N_3850);
nand U4071 (N_4071,N_3963,N_3524);
and U4072 (N_4072,N_3182,N_3449);
nor U4073 (N_4073,N_3867,N_3126);
nor U4074 (N_4074,N_3582,N_3992);
and U4075 (N_4075,N_3975,N_3514);
nor U4076 (N_4076,N_3085,N_3838);
xor U4077 (N_4077,N_3970,N_3729);
and U4078 (N_4078,N_3673,N_3110);
and U4079 (N_4079,N_3581,N_3643);
and U4080 (N_4080,N_3385,N_3878);
nand U4081 (N_4081,N_3005,N_3879);
or U4082 (N_4082,N_3848,N_3906);
nand U4083 (N_4083,N_3272,N_3437);
or U4084 (N_4084,N_3542,N_3857);
or U4085 (N_4085,N_3714,N_3455);
and U4086 (N_4086,N_3319,N_3652);
nand U4087 (N_4087,N_3779,N_3470);
or U4088 (N_4088,N_3158,N_3048);
nand U4089 (N_4089,N_3480,N_3892);
nor U4090 (N_4090,N_3331,N_3275);
and U4091 (N_4091,N_3745,N_3641);
or U4092 (N_4092,N_3088,N_3463);
nor U4093 (N_4093,N_3472,N_3672);
and U4094 (N_4094,N_3020,N_3904);
nor U4095 (N_4095,N_3003,N_3809);
and U4096 (N_4096,N_3622,N_3012);
or U4097 (N_4097,N_3359,N_3941);
nor U4098 (N_4098,N_3503,N_3988);
and U4099 (N_4099,N_3035,N_3215);
nand U4100 (N_4100,N_3043,N_3305);
or U4101 (N_4101,N_3469,N_3420);
or U4102 (N_4102,N_3694,N_3880);
or U4103 (N_4103,N_3277,N_3221);
and U4104 (N_4104,N_3298,N_3883);
or U4105 (N_4105,N_3789,N_3203);
nor U4106 (N_4106,N_3810,N_3321);
and U4107 (N_4107,N_3307,N_3464);
nand U4108 (N_4108,N_3504,N_3601);
or U4109 (N_4109,N_3640,N_3572);
or U4110 (N_4110,N_3711,N_3527);
xor U4111 (N_4111,N_3682,N_3719);
or U4112 (N_4112,N_3667,N_3744);
or U4113 (N_4113,N_3253,N_3511);
nand U4114 (N_4114,N_3353,N_3299);
or U4115 (N_4115,N_3380,N_3565);
and U4116 (N_4116,N_3056,N_3069);
or U4117 (N_4117,N_3525,N_3544);
or U4118 (N_4118,N_3981,N_3400);
nor U4119 (N_4119,N_3706,N_3351);
and U4120 (N_4120,N_3580,N_3423);
and U4121 (N_4121,N_3083,N_3814);
nand U4122 (N_4122,N_3358,N_3130);
nand U4123 (N_4123,N_3881,N_3274);
or U4124 (N_4124,N_3658,N_3617);
xnor U4125 (N_4125,N_3865,N_3096);
xor U4126 (N_4126,N_3258,N_3775);
nand U4127 (N_4127,N_3047,N_3248);
and U4128 (N_4128,N_3819,N_3914);
and U4129 (N_4129,N_3487,N_3995);
and U4130 (N_4130,N_3038,N_3833);
or U4131 (N_4131,N_3446,N_3063);
nor U4132 (N_4132,N_3761,N_3588);
or U4133 (N_4133,N_3561,N_3960);
and U4134 (N_4134,N_3839,N_3606);
and U4135 (N_4135,N_3366,N_3997);
and U4136 (N_4136,N_3486,N_3064);
and U4137 (N_4137,N_3004,N_3303);
nor U4138 (N_4138,N_3481,N_3836);
nand U4139 (N_4139,N_3240,N_3345);
xor U4140 (N_4140,N_3650,N_3117);
or U4141 (N_4141,N_3555,N_3427);
xnor U4142 (N_4142,N_3796,N_3623);
or U4143 (N_4143,N_3885,N_3092);
and U4144 (N_4144,N_3102,N_3383);
or U4145 (N_4145,N_3727,N_3644);
and U4146 (N_4146,N_3259,N_3018);
nor U4147 (N_4147,N_3146,N_3972);
and U4148 (N_4148,N_3505,N_3993);
nor U4149 (N_4149,N_3645,N_3151);
xnor U4150 (N_4150,N_3619,N_3046);
or U4151 (N_4151,N_3614,N_3287);
or U4152 (N_4152,N_3490,N_3492);
nand U4153 (N_4153,N_3842,N_3549);
nor U4154 (N_4154,N_3116,N_3440);
nand U4155 (N_4155,N_3685,N_3863);
or U4156 (N_4156,N_3337,N_3334);
or U4157 (N_4157,N_3315,N_3653);
xnor U4158 (N_4158,N_3447,N_3767);
nand U4159 (N_4159,N_3891,N_3501);
and U4160 (N_4160,N_3771,N_3160);
nor U4161 (N_4161,N_3924,N_3256);
xor U4162 (N_4162,N_3573,N_3935);
or U4163 (N_4163,N_3584,N_3300);
nand U4164 (N_4164,N_3609,N_3521);
and U4165 (N_4165,N_3647,N_3100);
nor U4166 (N_4166,N_3593,N_3586);
nand U4167 (N_4167,N_3079,N_3740);
xor U4168 (N_4168,N_3008,N_3297);
nor U4169 (N_4169,N_3246,N_3482);
nand U4170 (N_4170,N_3245,N_3495);
nand U4171 (N_4171,N_3161,N_3786);
or U4172 (N_4172,N_3214,N_3407);
nand U4173 (N_4173,N_3795,N_3206);
xnor U4174 (N_4174,N_3635,N_3462);
nor U4175 (N_4175,N_3379,N_3296);
or U4176 (N_4176,N_3147,N_3283);
nand U4177 (N_4177,N_3808,N_3661);
and U4178 (N_4178,N_3792,N_3874);
nand U4179 (N_4179,N_3216,N_3333);
or U4180 (N_4180,N_3564,N_3363);
and U4181 (N_4181,N_3843,N_3207);
xor U4182 (N_4182,N_3944,N_3458);
nand U4183 (N_4183,N_3718,N_3756);
nand U4184 (N_4184,N_3519,N_3841);
or U4185 (N_4185,N_3513,N_3651);
nor U4186 (N_4186,N_3224,N_3286);
nand U4187 (N_4187,N_3289,N_3243);
xor U4188 (N_4188,N_3461,N_3738);
nor U4189 (N_4189,N_3721,N_3201);
or U4190 (N_4190,N_3824,N_3691);
nor U4191 (N_4191,N_3120,N_3236);
nor U4192 (N_4192,N_3734,N_3080);
nor U4193 (N_4193,N_3949,N_3075);
and U4194 (N_4194,N_3763,N_3143);
nand U4195 (N_4195,N_3377,N_3965);
nor U4196 (N_4196,N_3531,N_3888);
or U4197 (N_4197,N_3019,N_3290);
nand U4198 (N_4198,N_3239,N_3457);
nor U4199 (N_4199,N_3750,N_3923);
nor U4200 (N_4200,N_3444,N_3101);
and U4201 (N_4201,N_3194,N_3421);
nor U4202 (N_4202,N_3165,N_3176);
xnor U4203 (N_4203,N_3847,N_3627);
nor U4204 (N_4204,N_3826,N_3391);
nand U4205 (N_4205,N_3356,N_3148);
and U4206 (N_4206,N_3093,N_3168);
nand U4207 (N_4207,N_3189,N_3760);
or U4208 (N_4208,N_3350,N_3405);
or U4209 (N_4209,N_3835,N_3125);
and U4210 (N_4210,N_3144,N_3741);
nor U4211 (N_4211,N_3518,N_3633);
and U4212 (N_4212,N_3570,N_3712);
nand U4213 (N_4213,N_3953,N_3178);
and U4214 (N_4214,N_3362,N_3827);
or U4215 (N_4215,N_3790,N_3227);
and U4216 (N_4216,N_3416,N_3678);
or U4217 (N_4217,N_3604,N_3802);
nand U4218 (N_4218,N_3288,N_3670);
or U4219 (N_4219,N_3220,N_3493);
nor U4220 (N_4220,N_3817,N_3939);
or U4221 (N_4221,N_3475,N_3984);
nor U4222 (N_4222,N_3884,N_3109);
or U4223 (N_4223,N_3636,N_3783);
nor U4224 (N_4224,N_3155,N_3360);
xor U4225 (N_4225,N_3709,N_3365);
nor U4226 (N_4226,N_3361,N_3295);
nand U4227 (N_4227,N_3737,N_3509);
xnor U4228 (N_4228,N_3169,N_3392);
or U4229 (N_4229,N_3742,N_3174);
or U4230 (N_4230,N_3081,N_3566);
and U4231 (N_4231,N_3731,N_3699);
nand U4232 (N_4232,N_3530,N_3578);
nor U4233 (N_4233,N_3620,N_3467);
nand U4234 (N_4234,N_3666,N_3431);
nand U4235 (N_4235,N_3326,N_3608);
nor U4236 (N_4236,N_3060,N_3373);
nand U4237 (N_4237,N_3409,N_3386);
or U4238 (N_4238,N_3942,N_3094);
and U4239 (N_4239,N_3034,N_3098);
nand U4240 (N_4240,N_3341,N_3129);
xor U4241 (N_4241,N_3930,N_3724);
and U4242 (N_4242,N_3554,N_3660);
nor U4243 (N_4243,N_3323,N_3599);
or U4244 (N_4244,N_3823,N_3820);
nand U4245 (N_4245,N_3688,N_3017);
or U4246 (N_4246,N_3042,N_3086);
and U4247 (N_4247,N_3723,N_3929);
nor U4248 (N_4248,N_3276,N_3626);
nor U4249 (N_4249,N_3324,N_3774);
nor U4250 (N_4250,N_3702,N_3118);
or U4251 (N_4251,N_3336,N_3142);
xnor U4252 (N_4252,N_3574,N_3908);
and U4253 (N_4253,N_3829,N_3818);
nand U4254 (N_4254,N_3696,N_3252);
nand U4255 (N_4255,N_3106,N_3339);
nor U4256 (N_4256,N_3713,N_3560);
or U4257 (N_4257,N_3022,N_3170);
nor U4258 (N_4258,N_3213,N_3764);
or U4259 (N_4259,N_3119,N_3355);
nor U4260 (N_4260,N_3968,N_3983);
and U4261 (N_4261,N_3112,N_3587);
or U4262 (N_4262,N_3912,N_3517);
and U4263 (N_4263,N_3016,N_3612);
nor U4264 (N_4264,N_3435,N_3853);
or U4265 (N_4265,N_3145,N_3733);
or U4266 (N_4266,N_3346,N_3537);
nor U4267 (N_4267,N_3998,N_3154);
nand U4268 (N_4268,N_3639,N_3484);
or U4269 (N_4269,N_3002,N_3410);
nand U4270 (N_4270,N_3759,N_3269);
and U4271 (N_4271,N_3011,N_3015);
nor U4272 (N_4272,N_3690,N_3748);
and U4273 (N_4273,N_3067,N_3831);
nor U4274 (N_4274,N_3318,N_3255);
or U4275 (N_4275,N_3439,N_3115);
nand U4276 (N_4276,N_3969,N_3322);
nor U4277 (N_4277,N_3801,N_3664);
or U4278 (N_4278,N_3338,N_3671);
and U4279 (N_4279,N_3412,N_3466);
and U4280 (N_4280,N_3111,N_3180);
and U4281 (N_4281,N_3798,N_3279);
nor U4282 (N_4282,N_3913,N_3589);
xnor U4283 (N_4283,N_3657,N_3855);
or U4284 (N_4284,N_3233,N_3933);
or U4285 (N_4285,N_3059,N_3401);
or U4286 (N_4286,N_3476,N_3991);
and U4287 (N_4287,N_3556,N_3743);
xnor U4288 (N_4288,N_3097,N_3496);
and U4289 (N_4289,N_3971,N_3611);
nand U4290 (N_4290,N_3167,N_3585);
or U4291 (N_4291,N_3301,N_3522);
and U4292 (N_4292,N_3294,N_3442);
nor U4293 (N_4293,N_3202,N_3821);
and U4294 (N_4294,N_3683,N_3794);
nand U4295 (N_4295,N_3436,N_3162);
or U4296 (N_4296,N_3438,N_3876);
nor U4297 (N_4297,N_3844,N_3597);
and U4298 (N_4298,N_3896,N_3979);
xnor U4299 (N_4299,N_3621,N_3077);
xnor U4300 (N_4300,N_3705,N_3432);
and U4301 (N_4301,N_3958,N_3121);
nand U4302 (N_4302,N_3411,N_3171);
nor U4303 (N_4303,N_3583,N_3625);
and U4304 (N_4304,N_3834,N_3045);
nand U4305 (N_4305,N_3769,N_3569);
or U4306 (N_4306,N_3659,N_3348);
nor U4307 (N_4307,N_3579,N_3443);
xnor U4308 (N_4308,N_3137,N_3488);
nor U4309 (N_4309,N_3413,N_3945);
nor U4310 (N_4310,N_3113,N_3311);
nor U4311 (N_4311,N_3675,N_3225);
nor U4312 (N_4312,N_3708,N_3902);
or U4313 (N_4313,N_3428,N_3799);
and U4314 (N_4314,N_3404,N_3940);
and U4315 (N_4315,N_3887,N_3124);
nor U4316 (N_4316,N_3539,N_3852);
nor U4317 (N_4317,N_3175,N_3610);
nor U4318 (N_4318,N_3191,N_3397);
nor U4319 (N_4319,N_3285,N_3104);
nor U4320 (N_4320,N_3700,N_3232);
xor U4321 (N_4321,N_3367,N_3898);
and U4322 (N_4322,N_3825,N_3768);
or U4323 (N_4323,N_3291,N_3784);
nand U4324 (N_4324,N_3192,N_3424);
nand U4325 (N_4325,N_3864,N_3076);
nor U4326 (N_4326,N_3631,N_3780);
xor U4327 (N_4327,N_3687,N_3188);
and U4328 (N_4328,N_3393,N_3982);
nand U4329 (N_4329,N_3812,N_3494);
nor U4330 (N_4330,N_3138,N_3370);
nand U4331 (N_4331,N_3445,N_3907);
nand U4332 (N_4332,N_3547,N_3755);
xor U4333 (N_4333,N_3920,N_3164);
xor U4334 (N_4334,N_3332,N_3237);
nor U4335 (N_4335,N_3679,N_3273);
nor U4336 (N_4336,N_3663,N_3217);
xor U4337 (N_4337,N_3782,N_3306);
or U4338 (N_4338,N_3919,N_3489);
and U4339 (N_4339,N_3027,N_3454);
nand U4340 (N_4340,N_3535,N_3426);
or U4341 (N_4341,N_3634,N_3330);
or U4342 (N_4342,N_3703,N_3545);
or U4343 (N_4343,N_3058,N_3689);
nand U4344 (N_4344,N_3183,N_3050);
nand U4345 (N_4345,N_3918,N_3875);
nor U4346 (N_4346,N_3964,N_3375);
or U4347 (N_4347,N_3459,N_3281);
nor U4348 (N_4348,N_3230,N_3551);
nor U4349 (N_4349,N_3715,N_3414);
xnor U4350 (N_4350,N_3500,N_3567);
nand U4351 (N_4351,N_3936,N_3591);
and U4352 (N_4352,N_3009,N_3343);
nor U4353 (N_4353,N_3816,N_3603);
or U4354 (N_4354,N_3967,N_3868);
or U4355 (N_4355,N_3873,N_3140);
nor U4356 (N_4356,N_3133,N_3533);
nor U4357 (N_4357,N_3976,N_3931);
nand U4358 (N_4358,N_3395,N_3265);
and U4359 (N_4359,N_3893,N_3342);
nor U4360 (N_4360,N_3382,N_3219);
nor U4361 (N_4361,N_3707,N_3491);
xnor U4362 (N_4362,N_3722,N_3765);
nand U4363 (N_4363,N_3791,N_3736);
or U4364 (N_4364,N_3562,N_3777);
and U4365 (N_4365,N_3642,N_3516);
nor U4366 (N_4366,N_3686,N_3605);
nor U4367 (N_4367,N_3677,N_3251);
and U4368 (N_4368,N_3090,N_3450);
nor U4369 (N_4369,N_3204,N_3895);
and U4370 (N_4370,N_3398,N_3250);
nor U4371 (N_4371,N_3376,N_3190);
and U4372 (N_4372,N_3532,N_3107);
and U4373 (N_4373,N_3014,N_3793);
nand U4374 (N_4374,N_3576,N_3041);
or U4375 (N_4375,N_3840,N_3293);
and U4376 (N_4376,N_3477,N_3364);
and U4377 (N_4377,N_3095,N_3901);
nand U4378 (N_4378,N_3973,N_3049);
xnor U4379 (N_4379,N_3889,N_3552);
and U4380 (N_4380,N_3886,N_3507);
and U4381 (N_4381,N_3483,N_3928);
or U4382 (N_4382,N_3210,N_3529);
and U4383 (N_4383,N_3335,N_3152);
xnor U4384 (N_4384,N_3292,N_3613);
or U4385 (N_4385,N_3946,N_3776);
nor U4386 (N_4386,N_3804,N_3630);
and U4387 (N_4387,N_3899,N_3754);
or U4388 (N_4388,N_3072,N_3349);
nor U4389 (N_4389,N_3615,N_3284);
and U4390 (N_4390,N_3717,N_3177);
or U4391 (N_4391,N_3226,N_3628);
xor U4392 (N_4392,N_3985,N_3937);
nand U4393 (N_4393,N_3948,N_3238);
nor U4394 (N_4394,N_3378,N_3716);
nand U4395 (N_4395,N_3952,N_3434);
nand U4396 (N_4396,N_3934,N_3425);
or U4397 (N_4397,N_3926,N_3528);
xor U4398 (N_4398,N_3950,N_3354);
xnor U4399 (N_4399,N_3961,N_3257);
xor U4400 (N_4400,N_3592,N_3955);
nand U4401 (N_4401,N_3103,N_3244);
or U4402 (N_4402,N_3770,N_3959);
xor U4403 (N_4403,N_3832,N_3543);
or U4404 (N_4404,N_3131,N_3123);
and U4405 (N_4405,N_3499,N_3869);
and U4406 (N_4406,N_3082,N_3465);
nand U4407 (N_4407,N_3845,N_3858);
and U4408 (N_4408,N_3418,N_3989);
or U4409 (N_4409,N_3655,N_3114);
and U4410 (N_4410,N_3862,N_3730);
or U4411 (N_4411,N_3388,N_3693);
nor U4412 (N_4412,N_3523,N_3911);
or U4413 (N_4413,N_3105,N_3222);
nor U4414 (N_4414,N_3403,N_3595);
and U4415 (N_4415,N_3638,N_3897);
nor U4416 (N_4416,N_3903,N_3851);
and U4417 (N_4417,N_3229,N_3422);
nand U4418 (N_4418,N_3025,N_3456);
or U4419 (N_4419,N_3515,N_3371);
nand U4420 (N_4420,N_3656,N_3781);
or U4421 (N_4421,N_3732,N_3815);
or U4422 (N_4422,N_3921,N_3778);
nor U4423 (N_4423,N_3962,N_3762);
and U4424 (N_4424,N_3697,N_3668);
xnor U4425 (N_4425,N_3108,N_3394);
nand U4426 (N_4426,N_3540,N_3156);
and U4427 (N_4427,N_3710,N_3254);
and U4428 (N_4428,N_3417,N_3329);
or U4429 (N_4429,N_3195,N_3433);
nor U4430 (N_4430,N_3701,N_3308);
or U4431 (N_4431,N_3788,N_3890);
or U4432 (N_4432,N_3309,N_3787);
or U4433 (N_4433,N_3807,N_3205);
xor U4434 (N_4434,N_3441,N_3637);
or U4435 (N_4435,N_3073,N_3938);
and U4436 (N_4436,N_3150,N_3037);
and U4437 (N_4437,N_3026,N_3068);
nor U4438 (N_4438,N_3837,N_3328);
or U4439 (N_4439,N_3030,N_3084);
nor U4440 (N_4440,N_3674,N_3966);
nor U4441 (N_4441,N_3057,N_3310);
nor U4442 (N_4442,N_3806,N_3389);
nand U4443 (N_4443,N_3548,N_3772);
nor U4444 (N_4444,N_3186,N_3594);
nand U4445 (N_4445,N_3452,N_3803);
nand U4446 (N_4446,N_3263,N_3460);
or U4447 (N_4447,N_3249,N_3172);
and U4448 (N_4448,N_3905,N_3261);
nand U4449 (N_4449,N_3849,N_3173);
nor U4450 (N_4450,N_3980,N_3065);
xor U4451 (N_4451,N_3304,N_3598);
xor U4452 (N_4452,N_3052,N_3316);
and U4453 (N_4453,N_3340,N_3051);
nand U4454 (N_4454,N_3978,N_3001);
nand U4455 (N_4455,N_3749,N_3451);
nor U4456 (N_4456,N_3314,N_3369);
or U4457 (N_4457,N_3559,N_3070);
or U4458 (N_4458,N_3419,N_3735);
xnor U4459 (N_4459,N_3986,N_3271);
or U4460 (N_4460,N_3260,N_3698);
xor U4461 (N_4461,N_3184,N_3947);
nand U4462 (N_4462,N_3223,N_3536);
and U4463 (N_4463,N_3557,N_3266);
and U4464 (N_4464,N_3040,N_3479);
xnor U4465 (N_4465,N_3498,N_3900);
nor U4466 (N_4466,N_3861,N_3632);
and U4467 (N_4467,N_3078,N_3665);
nor U4468 (N_4468,N_3159,N_3909);
and U4469 (N_4469,N_3185,N_3071);
nor U4470 (N_4470,N_3624,N_3066);
xnor U4471 (N_4471,N_3055,N_3534);
nand U4472 (N_4472,N_3127,N_3357);
nand U4473 (N_4473,N_3010,N_3726);
nor U4474 (N_4474,N_3264,N_3822);
and U4475 (N_4475,N_3568,N_3021);
nor U4476 (N_4476,N_3347,N_3091);
nor U4477 (N_4477,N_3739,N_3374);
or U4478 (N_4478,N_3241,N_3526);
or U4479 (N_4479,N_3692,N_3087);
xor U4480 (N_4480,N_3209,N_3242);
nor U4481 (N_4481,N_3327,N_3996);
nand U4482 (N_4482,N_3943,N_3408);
or U4483 (N_4483,N_3478,N_3916);
and U4484 (N_4484,N_3390,N_3399);
nor U4485 (N_4485,N_3558,N_3746);
and U4486 (N_4486,N_3139,N_3681);
xor U4487 (N_4487,N_3198,N_3344);
nand U4488 (N_4488,N_3910,N_3977);
or U4489 (N_4489,N_3510,N_3163);
xnor U4490 (N_4490,N_3234,N_3031);
nand U4491 (N_4491,N_3474,N_3208);
or U4492 (N_4492,N_3654,N_3032);
or U4493 (N_4493,N_3211,N_3990);
and U4494 (N_4494,N_3773,N_3629);
or U4495 (N_4495,N_3062,N_3872);
or U4496 (N_4496,N_3704,N_3999);
nand U4497 (N_4497,N_3262,N_3956);
nor U4498 (N_4498,N_3312,N_3758);
nor U4499 (N_4499,N_3649,N_3036);
and U4500 (N_4500,N_3839,N_3752);
or U4501 (N_4501,N_3085,N_3364);
nor U4502 (N_4502,N_3142,N_3026);
nor U4503 (N_4503,N_3352,N_3727);
xnor U4504 (N_4504,N_3532,N_3895);
and U4505 (N_4505,N_3405,N_3762);
or U4506 (N_4506,N_3840,N_3826);
xor U4507 (N_4507,N_3154,N_3132);
nor U4508 (N_4508,N_3699,N_3257);
or U4509 (N_4509,N_3164,N_3329);
or U4510 (N_4510,N_3542,N_3131);
xnor U4511 (N_4511,N_3604,N_3418);
or U4512 (N_4512,N_3824,N_3389);
or U4513 (N_4513,N_3362,N_3168);
nor U4514 (N_4514,N_3548,N_3276);
and U4515 (N_4515,N_3713,N_3561);
nor U4516 (N_4516,N_3432,N_3022);
or U4517 (N_4517,N_3130,N_3987);
nor U4518 (N_4518,N_3718,N_3370);
nand U4519 (N_4519,N_3222,N_3503);
or U4520 (N_4520,N_3213,N_3890);
xor U4521 (N_4521,N_3947,N_3143);
and U4522 (N_4522,N_3550,N_3764);
and U4523 (N_4523,N_3609,N_3292);
xnor U4524 (N_4524,N_3475,N_3429);
nor U4525 (N_4525,N_3605,N_3749);
and U4526 (N_4526,N_3895,N_3527);
or U4527 (N_4527,N_3188,N_3753);
and U4528 (N_4528,N_3017,N_3396);
nor U4529 (N_4529,N_3694,N_3720);
nor U4530 (N_4530,N_3632,N_3327);
nor U4531 (N_4531,N_3885,N_3318);
nand U4532 (N_4532,N_3988,N_3579);
nor U4533 (N_4533,N_3070,N_3063);
or U4534 (N_4534,N_3325,N_3970);
nor U4535 (N_4535,N_3281,N_3009);
and U4536 (N_4536,N_3808,N_3144);
nand U4537 (N_4537,N_3731,N_3282);
nand U4538 (N_4538,N_3384,N_3262);
and U4539 (N_4539,N_3587,N_3135);
and U4540 (N_4540,N_3579,N_3213);
nor U4541 (N_4541,N_3627,N_3814);
or U4542 (N_4542,N_3813,N_3115);
nor U4543 (N_4543,N_3817,N_3731);
or U4544 (N_4544,N_3643,N_3904);
and U4545 (N_4545,N_3844,N_3836);
and U4546 (N_4546,N_3458,N_3192);
nand U4547 (N_4547,N_3931,N_3996);
nand U4548 (N_4548,N_3764,N_3640);
nand U4549 (N_4549,N_3398,N_3110);
nor U4550 (N_4550,N_3580,N_3460);
and U4551 (N_4551,N_3032,N_3166);
or U4552 (N_4552,N_3885,N_3304);
nand U4553 (N_4553,N_3796,N_3554);
nand U4554 (N_4554,N_3080,N_3962);
xnor U4555 (N_4555,N_3339,N_3082);
nor U4556 (N_4556,N_3760,N_3814);
nor U4557 (N_4557,N_3669,N_3892);
nor U4558 (N_4558,N_3107,N_3701);
and U4559 (N_4559,N_3313,N_3996);
nand U4560 (N_4560,N_3827,N_3087);
nor U4561 (N_4561,N_3060,N_3123);
and U4562 (N_4562,N_3804,N_3657);
nand U4563 (N_4563,N_3617,N_3059);
and U4564 (N_4564,N_3427,N_3853);
or U4565 (N_4565,N_3587,N_3425);
or U4566 (N_4566,N_3181,N_3633);
nor U4567 (N_4567,N_3443,N_3441);
xor U4568 (N_4568,N_3232,N_3272);
nand U4569 (N_4569,N_3200,N_3058);
nand U4570 (N_4570,N_3182,N_3159);
nand U4571 (N_4571,N_3280,N_3162);
or U4572 (N_4572,N_3803,N_3345);
nor U4573 (N_4573,N_3255,N_3894);
nor U4574 (N_4574,N_3796,N_3466);
or U4575 (N_4575,N_3237,N_3428);
and U4576 (N_4576,N_3798,N_3619);
or U4577 (N_4577,N_3934,N_3255);
and U4578 (N_4578,N_3893,N_3455);
or U4579 (N_4579,N_3576,N_3995);
nor U4580 (N_4580,N_3155,N_3326);
nor U4581 (N_4581,N_3699,N_3458);
nor U4582 (N_4582,N_3971,N_3140);
nor U4583 (N_4583,N_3038,N_3352);
xnor U4584 (N_4584,N_3585,N_3415);
nor U4585 (N_4585,N_3544,N_3788);
or U4586 (N_4586,N_3200,N_3239);
nand U4587 (N_4587,N_3650,N_3480);
nor U4588 (N_4588,N_3507,N_3973);
and U4589 (N_4589,N_3048,N_3987);
and U4590 (N_4590,N_3409,N_3362);
or U4591 (N_4591,N_3012,N_3944);
xor U4592 (N_4592,N_3874,N_3091);
nor U4593 (N_4593,N_3039,N_3741);
nand U4594 (N_4594,N_3808,N_3577);
or U4595 (N_4595,N_3528,N_3511);
xnor U4596 (N_4596,N_3226,N_3473);
and U4597 (N_4597,N_3285,N_3689);
or U4598 (N_4598,N_3404,N_3843);
xor U4599 (N_4599,N_3048,N_3271);
and U4600 (N_4600,N_3224,N_3592);
nor U4601 (N_4601,N_3688,N_3661);
nand U4602 (N_4602,N_3439,N_3856);
nand U4603 (N_4603,N_3839,N_3450);
nand U4604 (N_4604,N_3299,N_3803);
nor U4605 (N_4605,N_3400,N_3048);
nand U4606 (N_4606,N_3898,N_3687);
nand U4607 (N_4607,N_3239,N_3983);
or U4608 (N_4608,N_3348,N_3240);
or U4609 (N_4609,N_3749,N_3745);
or U4610 (N_4610,N_3199,N_3073);
or U4611 (N_4611,N_3750,N_3536);
or U4612 (N_4612,N_3664,N_3098);
nor U4613 (N_4613,N_3130,N_3477);
and U4614 (N_4614,N_3851,N_3535);
xnor U4615 (N_4615,N_3147,N_3626);
and U4616 (N_4616,N_3851,N_3261);
and U4617 (N_4617,N_3241,N_3788);
and U4618 (N_4618,N_3472,N_3235);
or U4619 (N_4619,N_3212,N_3039);
and U4620 (N_4620,N_3229,N_3102);
nand U4621 (N_4621,N_3232,N_3524);
nor U4622 (N_4622,N_3949,N_3748);
and U4623 (N_4623,N_3048,N_3344);
nand U4624 (N_4624,N_3429,N_3082);
nor U4625 (N_4625,N_3509,N_3284);
nor U4626 (N_4626,N_3878,N_3359);
xor U4627 (N_4627,N_3743,N_3609);
and U4628 (N_4628,N_3490,N_3980);
or U4629 (N_4629,N_3361,N_3922);
and U4630 (N_4630,N_3084,N_3877);
xnor U4631 (N_4631,N_3600,N_3632);
and U4632 (N_4632,N_3148,N_3085);
nand U4633 (N_4633,N_3019,N_3727);
and U4634 (N_4634,N_3775,N_3321);
nor U4635 (N_4635,N_3450,N_3557);
or U4636 (N_4636,N_3722,N_3532);
or U4637 (N_4637,N_3430,N_3110);
nor U4638 (N_4638,N_3477,N_3026);
or U4639 (N_4639,N_3501,N_3357);
nor U4640 (N_4640,N_3592,N_3074);
or U4641 (N_4641,N_3522,N_3316);
nor U4642 (N_4642,N_3094,N_3729);
or U4643 (N_4643,N_3053,N_3805);
xnor U4644 (N_4644,N_3284,N_3211);
and U4645 (N_4645,N_3326,N_3437);
xnor U4646 (N_4646,N_3371,N_3293);
and U4647 (N_4647,N_3155,N_3276);
or U4648 (N_4648,N_3523,N_3108);
or U4649 (N_4649,N_3895,N_3826);
or U4650 (N_4650,N_3566,N_3626);
nand U4651 (N_4651,N_3717,N_3866);
or U4652 (N_4652,N_3043,N_3705);
and U4653 (N_4653,N_3931,N_3914);
nand U4654 (N_4654,N_3032,N_3795);
or U4655 (N_4655,N_3451,N_3196);
and U4656 (N_4656,N_3939,N_3186);
or U4657 (N_4657,N_3915,N_3369);
or U4658 (N_4658,N_3412,N_3489);
nand U4659 (N_4659,N_3474,N_3524);
xor U4660 (N_4660,N_3770,N_3663);
or U4661 (N_4661,N_3584,N_3107);
or U4662 (N_4662,N_3116,N_3565);
nor U4663 (N_4663,N_3979,N_3079);
nand U4664 (N_4664,N_3222,N_3542);
xnor U4665 (N_4665,N_3511,N_3965);
nor U4666 (N_4666,N_3662,N_3337);
nor U4667 (N_4667,N_3110,N_3819);
and U4668 (N_4668,N_3833,N_3926);
and U4669 (N_4669,N_3949,N_3253);
and U4670 (N_4670,N_3517,N_3317);
nor U4671 (N_4671,N_3185,N_3848);
nor U4672 (N_4672,N_3823,N_3728);
and U4673 (N_4673,N_3485,N_3026);
xor U4674 (N_4674,N_3655,N_3782);
nor U4675 (N_4675,N_3742,N_3810);
nand U4676 (N_4676,N_3948,N_3689);
nor U4677 (N_4677,N_3100,N_3739);
and U4678 (N_4678,N_3762,N_3497);
nor U4679 (N_4679,N_3856,N_3999);
and U4680 (N_4680,N_3314,N_3800);
or U4681 (N_4681,N_3653,N_3115);
nand U4682 (N_4682,N_3152,N_3101);
or U4683 (N_4683,N_3247,N_3451);
xnor U4684 (N_4684,N_3553,N_3452);
or U4685 (N_4685,N_3564,N_3210);
nand U4686 (N_4686,N_3601,N_3645);
or U4687 (N_4687,N_3237,N_3660);
nor U4688 (N_4688,N_3748,N_3023);
xor U4689 (N_4689,N_3455,N_3675);
nand U4690 (N_4690,N_3858,N_3563);
or U4691 (N_4691,N_3647,N_3608);
nand U4692 (N_4692,N_3029,N_3882);
nand U4693 (N_4693,N_3929,N_3604);
or U4694 (N_4694,N_3371,N_3047);
and U4695 (N_4695,N_3017,N_3049);
or U4696 (N_4696,N_3878,N_3649);
and U4697 (N_4697,N_3930,N_3719);
nand U4698 (N_4698,N_3842,N_3764);
nor U4699 (N_4699,N_3249,N_3983);
nand U4700 (N_4700,N_3635,N_3773);
nor U4701 (N_4701,N_3360,N_3125);
or U4702 (N_4702,N_3445,N_3935);
and U4703 (N_4703,N_3148,N_3719);
or U4704 (N_4704,N_3527,N_3765);
nor U4705 (N_4705,N_3018,N_3293);
or U4706 (N_4706,N_3432,N_3234);
nor U4707 (N_4707,N_3576,N_3186);
nand U4708 (N_4708,N_3830,N_3400);
xnor U4709 (N_4709,N_3228,N_3993);
nor U4710 (N_4710,N_3590,N_3983);
and U4711 (N_4711,N_3827,N_3981);
xor U4712 (N_4712,N_3859,N_3690);
nor U4713 (N_4713,N_3403,N_3482);
nand U4714 (N_4714,N_3095,N_3277);
or U4715 (N_4715,N_3966,N_3244);
or U4716 (N_4716,N_3175,N_3691);
nand U4717 (N_4717,N_3096,N_3899);
or U4718 (N_4718,N_3290,N_3017);
nor U4719 (N_4719,N_3335,N_3984);
nor U4720 (N_4720,N_3726,N_3705);
nand U4721 (N_4721,N_3658,N_3665);
nor U4722 (N_4722,N_3869,N_3570);
or U4723 (N_4723,N_3011,N_3732);
nor U4724 (N_4724,N_3018,N_3747);
nor U4725 (N_4725,N_3462,N_3397);
nor U4726 (N_4726,N_3090,N_3696);
nand U4727 (N_4727,N_3719,N_3458);
or U4728 (N_4728,N_3351,N_3450);
nor U4729 (N_4729,N_3387,N_3796);
nand U4730 (N_4730,N_3334,N_3661);
or U4731 (N_4731,N_3775,N_3070);
xor U4732 (N_4732,N_3150,N_3159);
or U4733 (N_4733,N_3153,N_3088);
or U4734 (N_4734,N_3006,N_3088);
nor U4735 (N_4735,N_3365,N_3647);
and U4736 (N_4736,N_3062,N_3812);
nor U4737 (N_4737,N_3812,N_3155);
or U4738 (N_4738,N_3808,N_3294);
and U4739 (N_4739,N_3869,N_3575);
and U4740 (N_4740,N_3228,N_3365);
or U4741 (N_4741,N_3139,N_3095);
nand U4742 (N_4742,N_3777,N_3184);
or U4743 (N_4743,N_3671,N_3002);
nor U4744 (N_4744,N_3884,N_3394);
and U4745 (N_4745,N_3298,N_3712);
nand U4746 (N_4746,N_3477,N_3707);
or U4747 (N_4747,N_3853,N_3897);
and U4748 (N_4748,N_3190,N_3356);
and U4749 (N_4749,N_3906,N_3841);
or U4750 (N_4750,N_3367,N_3957);
nor U4751 (N_4751,N_3735,N_3311);
nand U4752 (N_4752,N_3183,N_3069);
or U4753 (N_4753,N_3989,N_3388);
and U4754 (N_4754,N_3193,N_3729);
or U4755 (N_4755,N_3435,N_3469);
and U4756 (N_4756,N_3109,N_3107);
and U4757 (N_4757,N_3470,N_3207);
and U4758 (N_4758,N_3452,N_3878);
nand U4759 (N_4759,N_3713,N_3063);
nand U4760 (N_4760,N_3099,N_3594);
nand U4761 (N_4761,N_3508,N_3369);
nor U4762 (N_4762,N_3543,N_3260);
and U4763 (N_4763,N_3064,N_3491);
or U4764 (N_4764,N_3531,N_3535);
nand U4765 (N_4765,N_3774,N_3558);
xor U4766 (N_4766,N_3073,N_3998);
nor U4767 (N_4767,N_3774,N_3772);
nand U4768 (N_4768,N_3721,N_3956);
xor U4769 (N_4769,N_3116,N_3107);
nand U4770 (N_4770,N_3232,N_3993);
nor U4771 (N_4771,N_3322,N_3015);
and U4772 (N_4772,N_3638,N_3989);
and U4773 (N_4773,N_3058,N_3822);
or U4774 (N_4774,N_3125,N_3769);
or U4775 (N_4775,N_3578,N_3193);
nand U4776 (N_4776,N_3814,N_3612);
xnor U4777 (N_4777,N_3408,N_3768);
or U4778 (N_4778,N_3769,N_3424);
nand U4779 (N_4779,N_3583,N_3024);
and U4780 (N_4780,N_3752,N_3597);
xor U4781 (N_4781,N_3557,N_3668);
nand U4782 (N_4782,N_3721,N_3811);
and U4783 (N_4783,N_3578,N_3459);
nor U4784 (N_4784,N_3051,N_3843);
xnor U4785 (N_4785,N_3244,N_3461);
and U4786 (N_4786,N_3767,N_3327);
nor U4787 (N_4787,N_3727,N_3852);
or U4788 (N_4788,N_3324,N_3597);
and U4789 (N_4789,N_3931,N_3906);
nor U4790 (N_4790,N_3254,N_3961);
or U4791 (N_4791,N_3153,N_3004);
nand U4792 (N_4792,N_3195,N_3637);
nand U4793 (N_4793,N_3635,N_3639);
nand U4794 (N_4794,N_3005,N_3483);
and U4795 (N_4795,N_3805,N_3474);
nand U4796 (N_4796,N_3103,N_3092);
or U4797 (N_4797,N_3507,N_3188);
or U4798 (N_4798,N_3977,N_3172);
xor U4799 (N_4799,N_3518,N_3179);
nand U4800 (N_4800,N_3736,N_3001);
nor U4801 (N_4801,N_3133,N_3782);
and U4802 (N_4802,N_3291,N_3743);
nor U4803 (N_4803,N_3665,N_3111);
or U4804 (N_4804,N_3247,N_3911);
or U4805 (N_4805,N_3381,N_3598);
or U4806 (N_4806,N_3683,N_3080);
xor U4807 (N_4807,N_3566,N_3538);
nand U4808 (N_4808,N_3437,N_3868);
or U4809 (N_4809,N_3081,N_3860);
and U4810 (N_4810,N_3127,N_3630);
xor U4811 (N_4811,N_3846,N_3920);
and U4812 (N_4812,N_3809,N_3197);
nor U4813 (N_4813,N_3963,N_3105);
and U4814 (N_4814,N_3804,N_3038);
nand U4815 (N_4815,N_3995,N_3859);
nand U4816 (N_4816,N_3005,N_3575);
nand U4817 (N_4817,N_3670,N_3311);
or U4818 (N_4818,N_3554,N_3297);
nor U4819 (N_4819,N_3887,N_3377);
or U4820 (N_4820,N_3347,N_3606);
nand U4821 (N_4821,N_3650,N_3460);
nor U4822 (N_4822,N_3953,N_3048);
or U4823 (N_4823,N_3268,N_3915);
nor U4824 (N_4824,N_3628,N_3466);
nand U4825 (N_4825,N_3942,N_3296);
or U4826 (N_4826,N_3963,N_3254);
and U4827 (N_4827,N_3693,N_3877);
nor U4828 (N_4828,N_3087,N_3182);
and U4829 (N_4829,N_3079,N_3512);
and U4830 (N_4830,N_3916,N_3302);
or U4831 (N_4831,N_3865,N_3123);
nand U4832 (N_4832,N_3669,N_3250);
nand U4833 (N_4833,N_3090,N_3405);
or U4834 (N_4834,N_3148,N_3975);
nand U4835 (N_4835,N_3379,N_3426);
xnor U4836 (N_4836,N_3479,N_3697);
nor U4837 (N_4837,N_3351,N_3092);
xor U4838 (N_4838,N_3547,N_3226);
nand U4839 (N_4839,N_3042,N_3263);
or U4840 (N_4840,N_3483,N_3590);
nor U4841 (N_4841,N_3085,N_3791);
or U4842 (N_4842,N_3544,N_3230);
and U4843 (N_4843,N_3554,N_3990);
or U4844 (N_4844,N_3579,N_3057);
and U4845 (N_4845,N_3731,N_3956);
or U4846 (N_4846,N_3429,N_3897);
or U4847 (N_4847,N_3710,N_3547);
nand U4848 (N_4848,N_3597,N_3526);
or U4849 (N_4849,N_3042,N_3490);
nor U4850 (N_4850,N_3751,N_3874);
and U4851 (N_4851,N_3946,N_3869);
and U4852 (N_4852,N_3850,N_3732);
or U4853 (N_4853,N_3825,N_3704);
nor U4854 (N_4854,N_3632,N_3576);
nand U4855 (N_4855,N_3410,N_3097);
nor U4856 (N_4856,N_3544,N_3906);
nand U4857 (N_4857,N_3928,N_3705);
or U4858 (N_4858,N_3810,N_3376);
xnor U4859 (N_4859,N_3205,N_3785);
nand U4860 (N_4860,N_3323,N_3735);
nor U4861 (N_4861,N_3694,N_3811);
nor U4862 (N_4862,N_3841,N_3309);
nand U4863 (N_4863,N_3427,N_3183);
and U4864 (N_4864,N_3507,N_3278);
and U4865 (N_4865,N_3625,N_3049);
or U4866 (N_4866,N_3315,N_3285);
or U4867 (N_4867,N_3415,N_3952);
nand U4868 (N_4868,N_3552,N_3814);
nand U4869 (N_4869,N_3301,N_3960);
and U4870 (N_4870,N_3646,N_3408);
nand U4871 (N_4871,N_3779,N_3948);
or U4872 (N_4872,N_3080,N_3599);
nand U4873 (N_4873,N_3040,N_3616);
and U4874 (N_4874,N_3538,N_3940);
nor U4875 (N_4875,N_3866,N_3122);
and U4876 (N_4876,N_3790,N_3946);
nor U4877 (N_4877,N_3797,N_3658);
or U4878 (N_4878,N_3363,N_3669);
nand U4879 (N_4879,N_3666,N_3952);
or U4880 (N_4880,N_3380,N_3538);
nor U4881 (N_4881,N_3465,N_3592);
or U4882 (N_4882,N_3164,N_3695);
or U4883 (N_4883,N_3184,N_3622);
or U4884 (N_4884,N_3419,N_3707);
nand U4885 (N_4885,N_3129,N_3405);
nor U4886 (N_4886,N_3049,N_3065);
and U4887 (N_4887,N_3639,N_3173);
and U4888 (N_4888,N_3752,N_3587);
or U4889 (N_4889,N_3290,N_3215);
or U4890 (N_4890,N_3191,N_3178);
or U4891 (N_4891,N_3173,N_3122);
xnor U4892 (N_4892,N_3848,N_3382);
and U4893 (N_4893,N_3587,N_3945);
and U4894 (N_4894,N_3786,N_3341);
nand U4895 (N_4895,N_3187,N_3879);
nand U4896 (N_4896,N_3421,N_3208);
xnor U4897 (N_4897,N_3332,N_3384);
xor U4898 (N_4898,N_3243,N_3111);
and U4899 (N_4899,N_3110,N_3151);
and U4900 (N_4900,N_3347,N_3966);
and U4901 (N_4901,N_3865,N_3044);
and U4902 (N_4902,N_3463,N_3813);
and U4903 (N_4903,N_3664,N_3694);
nand U4904 (N_4904,N_3420,N_3128);
and U4905 (N_4905,N_3749,N_3172);
nor U4906 (N_4906,N_3063,N_3002);
and U4907 (N_4907,N_3094,N_3230);
nor U4908 (N_4908,N_3802,N_3469);
or U4909 (N_4909,N_3987,N_3531);
xor U4910 (N_4910,N_3557,N_3127);
nand U4911 (N_4911,N_3539,N_3470);
or U4912 (N_4912,N_3547,N_3694);
nand U4913 (N_4913,N_3838,N_3880);
or U4914 (N_4914,N_3692,N_3842);
xnor U4915 (N_4915,N_3306,N_3419);
nand U4916 (N_4916,N_3276,N_3772);
nor U4917 (N_4917,N_3773,N_3591);
xnor U4918 (N_4918,N_3812,N_3529);
nand U4919 (N_4919,N_3869,N_3198);
nand U4920 (N_4920,N_3622,N_3950);
nand U4921 (N_4921,N_3429,N_3842);
nand U4922 (N_4922,N_3582,N_3697);
or U4923 (N_4923,N_3242,N_3736);
and U4924 (N_4924,N_3802,N_3246);
nand U4925 (N_4925,N_3709,N_3344);
and U4926 (N_4926,N_3231,N_3721);
xnor U4927 (N_4927,N_3589,N_3357);
nand U4928 (N_4928,N_3926,N_3647);
and U4929 (N_4929,N_3946,N_3071);
nand U4930 (N_4930,N_3192,N_3433);
or U4931 (N_4931,N_3683,N_3696);
and U4932 (N_4932,N_3563,N_3627);
nor U4933 (N_4933,N_3780,N_3131);
xor U4934 (N_4934,N_3411,N_3661);
nand U4935 (N_4935,N_3466,N_3940);
xnor U4936 (N_4936,N_3067,N_3759);
nand U4937 (N_4937,N_3489,N_3777);
or U4938 (N_4938,N_3686,N_3714);
nor U4939 (N_4939,N_3047,N_3459);
nor U4940 (N_4940,N_3042,N_3305);
xnor U4941 (N_4941,N_3816,N_3398);
nor U4942 (N_4942,N_3177,N_3251);
and U4943 (N_4943,N_3532,N_3718);
or U4944 (N_4944,N_3918,N_3798);
and U4945 (N_4945,N_3447,N_3598);
xor U4946 (N_4946,N_3352,N_3403);
xnor U4947 (N_4947,N_3844,N_3811);
nor U4948 (N_4948,N_3437,N_3015);
and U4949 (N_4949,N_3037,N_3177);
or U4950 (N_4950,N_3976,N_3836);
nor U4951 (N_4951,N_3920,N_3522);
nand U4952 (N_4952,N_3484,N_3937);
and U4953 (N_4953,N_3781,N_3594);
and U4954 (N_4954,N_3163,N_3388);
and U4955 (N_4955,N_3582,N_3366);
or U4956 (N_4956,N_3769,N_3103);
and U4957 (N_4957,N_3203,N_3278);
nand U4958 (N_4958,N_3473,N_3242);
nor U4959 (N_4959,N_3230,N_3318);
nor U4960 (N_4960,N_3873,N_3636);
nor U4961 (N_4961,N_3311,N_3488);
or U4962 (N_4962,N_3491,N_3840);
and U4963 (N_4963,N_3810,N_3737);
nand U4964 (N_4964,N_3856,N_3298);
nand U4965 (N_4965,N_3982,N_3818);
xnor U4966 (N_4966,N_3398,N_3863);
or U4967 (N_4967,N_3007,N_3860);
or U4968 (N_4968,N_3209,N_3935);
and U4969 (N_4969,N_3748,N_3729);
and U4970 (N_4970,N_3661,N_3337);
and U4971 (N_4971,N_3175,N_3718);
or U4972 (N_4972,N_3331,N_3268);
nor U4973 (N_4973,N_3089,N_3963);
nand U4974 (N_4974,N_3569,N_3191);
nor U4975 (N_4975,N_3217,N_3631);
xor U4976 (N_4976,N_3176,N_3280);
nand U4977 (N_4977,N_3495,N_3573);
nor U4978 (N_4978,N_3895,N_3902);
and U4979 (N_4979,N_3630,N_3932);
nor U4980 (N_4980,N_3847,N_3117);
xnor U4981 (N_4981,N_3827,N_3305);
and U4982 (N_4982,N_3782,N_3662);
nor U4983 (N_4983,N_3123,N_3626);
nor U4984 (N_4984,N_3104,N_3452);
nor U4985 (N_4985,N_3675,N_3606);
and U4986 (N_4986,N_3336,N_3208);
and U4987 (N_4987,N_3657,N_3619);
xor U4988 (N_4988,N_3255,N_3613);
nand U4989 (N_4989,N_3932,N_3378);
and U4990 (N_4990,N_3236,N_3217);
nor U4991 (N_4991,N_3707,N_3845);
and U4992 (N_4992,N_3937,N_3619);
or U4993 (N_4993,N_3219,N_3135);
and U4994 (N_4994,N_3396,N_3462);
nand U4995 (N_4995,N_3175,N_3271);
or U4996 (N_4996,N_3905,N_3287);
or U4997 (N_4997,N_3213,N_3544);
and U4998 (N_4998,N_3949,N_3865);
nor U4999 (N_4999,N_3692,N_3097);
or UO_0 (O_0,N_4116,N_4166);
xor UO_1 (O_1,N_4551,N_4845);
xor UO_2 (O_2,N_4142,N_4029);
xor UO_3 (O_3,N_4396,N_4727);
and UO_4 (O_4,N_4780,N_4145);
and UO_5 (O_5,N_4947,N_4352);
nor UO_6 (O_6,N_4858,N_4067);
nor UO_7 (O_7,N_4597,N_4457);
nand UO_8 (O_8,N_4185,N_4903);
or UO_9 (O_9,N_4991,N_4507);
nand UO_10 (O_10,N_4515,N_4082);
and UO_11 (O_11,N_4728,N_4688);
or UO_12 (O_12,N_4062,N_4025);
nand UO_13 (O_13,N_4641,N_4754);
nor UO_14 (O_14,N_4246,N_4004);
nand UO_15 (O_15,N_4623,N_4872);
or UO_16 (O_16,N_4472,N_4381);
nand UO_17 (O_17,N_4708,N_4810);
or UO_18 (O_18,N_4096,N_4178);
nor UO_19 (O_19,N_4588,N_4385);
nand UO_20 (O_20,N_4379,N_4630);
nor UO_21 (O_21,N_4408,N_4935);
nand UO_22 (O_22,N_4198,N_4536);
nand UO_23 (O_23,N_4672,N_4291);
xor UO_24 (O_24,N_4686,N_4595);
and UO_25 (O_25,N_4348,N_4835);
nand UO_26 (O_26,N_4525,N_4661);
nand UO_27 (O_27,N_4806,N_4224);
and UO_28 (O_28,N_4059,N_4443);
and UO_29 (O_29,N_4932,N_4325);
and UO_30 (O_30,N_4288,N_4502);
nand UO_31 (O_31,N_4962,N_4985);
nand UO_32 (O_32,N_4775,N_4337);
nand UO_33 (O_33,N_4570,N_4216);
nor UO_34 (O_34,N_4383,N_4697);
and UO_35 (O_35,N_4434,N_4862);
nand UO_36 (O_36,N_4659,N_4492);
and UO_37 (O_37,N_4812,N_4479);
and UO_38 (O_38,N_4131,N_4821);
or UO_39 (O_39,N_4008,N_4531);
nor UO_40 (O_40,N_4388,N_4290);
nor UO_41 (O_41,N_4248,N_4762);
and UO_42 (O_42,N_4350,N_4374);
and UO_43 (O_43,N_4704,N_4868);
nor UO_44 (O_44,N_4860,N_4552);
nand UO_45 (O_45,N_4016,N_4820);
or UO_46 (O_46,N_4665,N_4929);
nand UO_47 (O_47,N_4347,N_4009);
nand UO_48 (O_48,N_4486,N_4683);
and UO_49 (O_49,N_4524,N_4395);
nor UO_50 (O_50,N_4458,N_4709);
nor UO_51 (O_51,N_4756,N_4996);
and UO_52 (O_52,N_4787,N_4968);
xor UO_53 (O_53,N_4323,N_4258);
nor UO_54 (O_54,N_4900,N_4828);
or UO_55 (O_55,N_4153,N_4508);
or UO_56 (O_56,N_4199,N_4169);
nand UO_57 (O_57,N_4529,N_4975);
and UO_58 (O_58,N_4275,N_4423);
nor UO_59 (O_59,N_4808,N_4783);
and UO_60 (O_60,N_4670,N_4411);
nand UO_61 (O_61,N_4882,N_4401);
or UO_62 (O_62,N_4539,N_4889);
nand UO_63 (O_63,N_4130,N_4738);
or UO_64 (O_64,N_4654,N_4462);
and UO_65 (O_65,N_4279,N_4612);
nand UO_66 (O_66,N_4941,N_4818);
and UO_67 (O_67,N_4015,N_4768);
nand UO_68 (O_68,N_4723,N_4600);
nand UO_69 (O_69,N_4755,N_4629);
and UO_70 (O_70,N_4563,N_4773);
nor UO_71 (O_71,N_4950,N_4518);
and UO_72 (O_72,N_4856,N_4281);
or UO_73 (O_73,N_4483,N_4249);
or UO_74 (O_74,N_4446,N_4440);
nand UO_75 (O_75,N_4316,N_4834);
nor UO_76 (O_76,N_4376,N_4003);
and UO_77 (O_77,N_4372,N_4952);
nor UO_78 (O_78,N_4102,N_4286);
nand UO_79 (O_79,N_4439,N_4310);
and UO_80 (O_80,N_4548,N_4874);
nor UO_81 (O_81,N_4026,N_4849);
nor UO_82 (O_82,N_4922,N_4657);
and UO_83 (O_83,N_4705,N_4645);
and UO_84 (O_84,N_4888,N_4099);
xor UO_85 (O_85,N_4306,N_4092);
and UO_86 (O_86,N_4087,N_4118);
nand UO_87 (O_87,N_4468,N_4135);
and UO_88 (O_88,N_4075,N_4829);
xor UO_89 (O_89,N_4471,N_4558);
nand UO_90 (O_90,N_4326,N_4115);
nor UO_91 (O_91,N_4898,N_4210);
nor UO_92 (O_92,N_4123,N_4170);
nor UO_93 (O_93,N_4542,N_4986);
nand UO_94 (O_94,N_4419,N_4865);
and UO_95 (O_95,N_4431,N_4490);
nor UO_96 (O_96,N_4073,N_4174);
nand UO_97 (O_97,N_4477,N_4740);
nor UO_98 (O_98,N_4220,N_4318);
or UO_99 (O_99,N_4392,N_4349);
and UO_100 (O_100,N_4072,N_4267);
and UO_101 (O_101,N_4724,N_4988);
nand UO_102 (O_102,N_4070,N_4071);
nor UO_103 (O_103,N_4041,N_4666);
nand UO_104 (O_104,N_4734,N_4211);
and UO_105 (O_105,N_4736,N_4180);
nand UO_106 (O_106,N_4273,N_4790);
and UO_107 (O_107,N_4944,N_4295);
or UO_108 (O_108,N_4864,N_4580);
or UO_109 (O_109,N_4535,N_4713);
nand UO_110 (O_110,N_4532,N_4887);
and UO_111 (O_111,N_4816,N_4857);
xnor UO_112 (O_112,N_4658,N_4896);
nand UO_113 (O_113,N_4157,N_4877);
or UO_114 (O_114,N_4549,N_4173);
nor UO_115 (O_115,N_4924,N_4160);
nor UO_116 (O_116,N_4863,N_4520);
xor UO_117 (O_117,N_4753,N_4319);
or UO_118 (O_118,N_4565,N_4582);
xnor UO_119 (O_119,N_4236,N_4353);
nand UO_120 (O_120,N_4989,N_4876);
nor UO_121 (O_121,N_4936,N_4403);
and UO_122 (O_122,N_4745,N_4107);
xnor UO_123 (O_123,N_4938,N_4052);
or UO_124 (O_124,N_4796,N_4801);
and UO_125 (O_125,N_4089,N_4496);
nand UO_126 (O_126,N_4470,N_4878);
and UO_127 (O_127,N_4636,N_4345);
nand UO_128 (O_128,N_4282,N_4194);
and UO_129 (O_129,N_4788,N_4843);
nor UO_130 (O_130,N_4296,N_4497);
nor UO_131 (O_131,N_4533,N_4589);
or UO_132 (O_132,N_4177,N_4425);
or UO_133 (O_133,N_4449,N_4424);
or UO_134 (O_134,N_4831,N_4807);
xnor UO_135 (O_135,N_4870,N_4769);
and UO_136 (O_136,N_4106,N_4933);
and UO_137 (O_137,N_4779,N_4967);
or UO_138 (O_138,N_4233,N_4585);
nor UO_139 (O_139,N_4019,N_4668);
and UO_140 (O_140,N_4368,N_4786);
xor UO_141 (O_141,N_4854,N_4561);
nand UO_142 (O_142,N_4676,N_4259);
nand UO_143 (O_143,N_4303,N_4250);
nand UO_144 (O_144,N_4873,N_4977);
or UO_145 (O_145,N_4133,N_4207);
and UO_146 (O_146,N_4719,N_4333);
nor UO_147 (O_147,N_4732,N_4189);
and UO_148 (O_148,N_4715,N_4839);
and UO_149 (O_149,N_4455,N_4038);
xor UO_150 (O_150,N_4778,N_4583);
or UO_151 (O_151,N_4712,N_4545);
and UO_152 (O_152,N_4761,N_4223);
or UO_153 (O_153,N_4114,N_4027);
nand UO_154 (O_154,N_4091,N_4201);
or UO_155 (O_155,N_4833,N_4797);
nand UO_156 (O_156,N_4921,N_4265);
or UO_157 (O_157,N_4257,N_4369);
or UO_158 (O_158,N_4167,N_4001);
nor UO_159 (O_159,N_4855,N_4940);
and UO_160 (O_160,N_4799,N_4138);
or UO_161 (O_161,N_4386,N_4244);
nand UO_162 (O_162,N_4811,N_4726);
nand UO_163 (O_163,N_4871,N_4809);
nor UO_164 (O_164,N_4897,N_4886);
or UO_165 (O_165,N_4108,N_4042);
nor UO_166 (O_166,N_4414,N_4866);
or UO_167 (O_167,N_4971,N_4074);
or UO_168 (O_168,N_4928,N_4032);
nor UO_169 (O_169,N_4599,N_4667);
and UO_170 (O_170,N_4113,N_4905);
or UO_171 (O_171,N_4766,N_4841);
nor UO_172 (O_172,N_4651,N_4315);
nor UO_173 (O_173,N_4733,N_4673);
and UO_174 (O_174,N_4716,N_4393);
nand UO_175 (O_175,N_4634,N_4321);
xnor UO_176 (O_176,N_4172,N_4689);
or UO_177 (O_177,N_4627,N_4010);
nand UO_178 (O_178,N_4238,N_4404);
and UO_179 (O_179,N_4503,N_4669);
and UO_180 (O_180,N_4023,N_4622);
xnor UO_181 (O_181,N_4421,N_4840);
nand UO_182 (O_182,N_4390,N_4464);
xor UO_183 (O_183,N_4541,N_4293);
or UO_184 (O_184,N_4292,N_4847);
xor UO_185 (O_185,N_4498,N_4024);
or UO_186 (O_186,N_4789,N_4491);
or UO_187 (O_187,N_4149,N_4322);
and UO_188 (O_188,N_4884,N_4328);
nor UO_189 (O_189,N_4137,N_4729);
nand UO_190 (O_190,N_4992,N_4313);
and UO_191 (O_191,N_4056,N_4330);
nor UO_192 (O_192,N_4798,N_4528);
and UO_193 (O_193,N_4191,N_4263);
or UO_194 (O_194,N_4981,N_4557);
xor UO_195 (O_195,N_4466,N_4662);
and UO_196 (O_196,N_4268,N_4362);
nand UO_197 (O_197,N_4150,N_4144);
or UO_198 (O_198,N_4183,N_4159);
xnor UO_199 (O_199,N_4710,N_4117);
or UO_200 (O_200,N_4367,N_4785);
and UO_201 (O_201,N_4516,N_4976);
or UO_202 (O_202,N_4299,N_4413);
and UO_203 (O_203,N_4744,N_4039);
xor UO_204 (O_204,N_4523,N_4053);
and UO_205 (O_205,N_4894,N_4500);
or UO_206 (O_206,N_4499,N_4221);
nor UO_207 (O_207,N_4982,N_4909);
nand UO_208 (O_208,N_4463,N_4815);
nor UO_209 (O_209,N_4495,N_4482);
and UO_210 (O_210,N_4690,N_4954);
xor UO_211 (O_211,N_4493,N_4359);
nor UO_212 (O_212,N_4742,N_4603);
and UO_213 (O_213,N_4791,N_4964);
nor UO_214 (O_214,N_4692,N_4842);
or UO_215 (O_215,N_4782,N_4602);
or UO_216 (O_216,N_4080,N_4002);
or UO_217 (O_217,N_4021,N_4478);
and UO_218 (O_218,N_4823,N_4202);
nand UO_219 (O_219,N_4934,N_4187);
nand UO_220 (O_220,N_4794,N_4994);
xor UO_221 (O_221,N_4747,N_4143);
nor UO_222 (O_222,N_4384,N_4848);
xor UO_223 (O_223,N_4714,N_4200);
or UO_224 (O_224,N_4939,N_4687);
nor UO_225 (O_225,N_4895,N_4550);
and UO_226 (O_226,N_4346,N_4800);
xnor UO_227 (O_227,N_4427,N_4453);
or UO_228 (O_228,N_4663,N_4925);
nor UO_229 (O_229,N_4718,N_4433);
and UO_230 (O_230,N_4355,N_4125);
nor UO_231 (O_231,N_4022,N_4320);
and UO_232 (O_232,N_4045,N_4360);
and UO_233 (O_233,N_4227,N_4832);
nand UO_234 (O_234,N_4767,N_4608);
or UO_235 (O_235,N_4266,N_4481);
or UO_236 (O_236,N_4949,N_4154);
nor UO_237 (O_237,N_4633,N_4112);
nand UO_238 (O_238,N_4624,N_4556);
nand UO_239 (O_239,N_4051,N_4494);
or UO_240 (O_240,N_4615,N_4540);
nor UO_241 (O_241,N_4474,N_4030);
nand UO_242 (O_242,N_4046,N_4721);
nor UO_243 (O_243,N_4122,N_4324);
nand UO_244 (O_244,N_4792,N_4918);
and UO_245 (O_245,N_4604,N_4093);
nand UO_246 (O_246,N_4095,N_4068);
nor UO_247 (O_247,N_4339,N_4429);
or UO_248 (O_248,N_4394,N_4011);
or UO_249 (O_249,N_4356,N_4906);
or UO_250 (O_250,N_4061,N_4338);
or UO_251 (O_251,N_4576,N_4640);
or UO_252 (O_252,N_4014,N_4642);
or UO_253 (O_253,N_4653,N_4127);
or UO_254 (O_254,N_4711,N_4892);
nor UO_255 (O_255,N_4880,N_4245);
and UO_256 (O_256,N_4475,N_4917);
and UO_257 (O_257,N_4579,N_4416);
or UO_258 (O_258,N_4047,N_4340);
nand UO_259 (O_259,N_4572,N_4526);
nand UO_260 (O_260,N_4217,N_4243);
nand UO_261 (O_261,N_4241,N_4262);
nor UO_262 (O_262,N_4336,N_4289);
and UO_263 (O_263,N_4237,N_4972);
nor UO_264 (O_264,N_4311,N_4447);
nor UO_265 (O_265,N_4239,N_4420);
nand UO_266 (O_266,N_4555,N_4229);
and UO_267 (O_267,N_4077,N_4625);
or UO_268 (O_268,N_4442,N_4639);
or UO_269 (O_269,N_4450,N_4737);
nor UO_270 (O_270,N_4487,N_4955);
nor UO_271 (O_271,N_4158,N_4119);
nand UO_272 (O_272,N_4136,N_4278);
nor UO_273 (O_273,N_4469,N_4456);
nor UO_274 (O_274,N_4152,N_4534);
and UO_275 (O_275,N_4054,N_4912);
and UO_276 (O_276,N_4701,N_4100);
and UO_277 (O_277,N_4104,N_4771);
or UO_278 (O_278,N_4448,N_4830);
nor UO_279 (O_279,N_4717,N_4838);
nor UO_280 (O_280,N_4410,N_4260);
or UO_281 (O_281,N_4691,N_4171);
and UO_282 (O_282,N_4121,N_4269);
or UO_283 (O_283,N_4436,N_4759);
nand UO_284 (O_284,N_4638,N_4997);
xor UO_285 (O_285,N_4521,N_4405);
nor UO_286 (O_286,N_4824,N_4007);
xnor UO_287 (O_287,N_4990,N_4276);
nor UO_288 (O_288,N_4943,N_4650);
nand UO_289 (O_289,N_4695,N_4389);
nand UO_290 (O_290,N_4930,N_4036);
or UO_291 (O_291,N_4937,N_4948);
and UO_292 (O_292,N_4357,N_4438);
or UO_293 (O_293,N_4140,N_4378);
or UO_294 (O_294,N_4147,N_4611);
nand UO_295 (O_295,N_4358,N_4432);
nand UO_296 (O_296,N_4048,N_4309);
or UO_297 (O_297,N_4272,N_4510);
and UO_298 (O_298,N_4722,N_4974);
nand UO_299 (O_299,N_4213,N_4097);
and UO_300 (O_300,N_4261,N_4228);
nor UO_301 (O_301,N_4538,N_4514);
or UO_302 (O_302,N_4527,N_4225);
xor UO_303 (O_303,N_4020,N_4836);
nor UO_304 (O_304,N_4752,N_4908);
xnor UO_305 (O_305,N_4837,N_4043);
nor UO_306 (O_306,N_4057,N_4120);
and UO_307 (O_307,N_4594,N_4033);
or UO_308 (O_308,N_4684,N_4215);
nor UO_309 (O_309,N_4957,N_4085);
and UO_310 (O_310,N_4825,N_4980);
nand UO_311 (O_311,N_4226,N_4146);
nand UO_312 (O_312,N_4387,N_4031);
nand UO_313 (O_313,N_4373,N_4567);
and UO_314 (O_314,N_4028,N_4979);
and UO_315 (O_315,N_4195,N_4664);
and UO_316 (O_316,N_4467,N_4298);
nand UO_317 (O_317,N_4465,N_4605);
nand UO_318 (O_318,N_4793,N_4370);
nor UO_319 (O_319,N_4619,N_4182);
nand UO_320 (O_320,N_4511,N_4546);
nand UO_321 (O_321,N_4277,N_4256);
or UO_322 (O_322,N_4418,N_4614);
nand UO_323 (O_323,N_4307,N_4560);
nand UO_324 (O_324,N_4616,N_4564);
or UO_325 (O_325,N_4763,N_4966);
nor UO_326 (O_326,N_4190,N_4040);
nand UO_327 (O_327,N_4537,N_4105);
and UO_328 (O_328,N_4331,N_4126);
or UO_329 (O_329,N_4601,N_4214);
nor UO_330 (O_330,N_4018,N_4205);
or UO_331 (O_331,N_4700,N_4817);
and UO_332 (O_332,N_4509,N_4079);
nor UO_333 (O_333,N_4720,N_4212);
nor UO_334 (O_334,N_4441,N_4451);
nor UO_335 (O_335,N_4592,N_4590);
or UO_336 (O_336,N_4678,N_4480);
nand UO_337 (O_337,N_4607,N_4251);
xnor UO_338 (O_338,N_4402,N_4308);
nand UO_339 (O_339,N_4682,N_4219);
nor UO_340 (O_340,N_4218,N_4757);
or UO_341 (O_341,N_4343,N_4013);
nor UO_342 (O_342,N_4517,N_4132);
xnor UO_343 (O_343,N_4805,N_4294);
nand UO_344 (O_344,N_4460,N_4513);
xnor UO_345 (O_345,N_4772,N_4885);
or UO_346 (O_346,N_4090,N_4553);
nor UO_347 (O_347,N_4803,N_4973);
and UO_348 (O_348,N_4861,N_4562);
nor UO_349 (O_349,N_4083,N_4312);
xnor UO_350 (O_350,N_4428,N_4883);
nand UO_351 (O_351,N_4066,N_4301);
nand UO_352 (O_352,N_4911,N_4270);
nor UO_353 (O_353,N_4240,N_4999);
xor UO_354 (O_354,N_4559,N_4648);
and UO_355 (O_355,N_4609,N_4910);
and UO_356 (O_356,N_4730,N_4060);
nand UO_357 (O_357,N_4875,N_4649);
xor UO_358 (O_358,N_4109,N_4504);
nand UO_359 (O_359,N_4179,N_4577);
nand UO_360 (O_360,N_4005,N_4501);
nand UO_361 (O_361,N_4231,N_4963);
nand UO_362 (O_362,N_4165,N_4366);
nand UO_363 (O_363,N_4965,N_4852);
nor UO_364 (O_364,N_4554,N_4488);
nand UO_365 (O_365,N_4680,N_4774);
or UO_366 (O_366,N_4012,N_4208);
nand UO_367 (O_367,N_4222,N_4591);
nand UO_368 (O_368,N_4620,N_4255);
nand UO_369 (O_369,N_4035,N_4445);
nand UO_370 (O_370,N_4902,N_4637);
nand UO_371 (O_371,N_4371,N_4881);
and UO_372 (O_372,N_4660,N_4430);
or UO_373 (O_373,N_4867,N_4086);
nand UO_374 (O_374,N_4000,N_4391);
nand UO_375 (O_375,N_4098,N_4890);
and UO_376 (O_376,N_4593,N_4959);
nand UO_377 (O_377,N_4969,N_4399);
and UO_378 (O_378,N_4646,N_4252);
nand UO_379 (O_379,N_4181,N_4891);
nor UO_380 (O_380,N_4505,N_4739);
and UO_381 (O_381,N_4081,N_4058);
or UO_382 (O_382,N_4644,N_4951);
or UO_383 (O_383,N_4613,N_4186);
xnor UO_384 (O_384,N_4899,N_4703);
or UO_385 (O_385,N_4827,N_4743);
and UO_386 (O_386,N_4017,N_4044);
nand UO_387 (O_387,N_4361,N_4784);
or UO_388 (O_388,N_4751,N_4846);
nand UO_389 (O_389,N_4234,N_4412);
and UO_390 (O_390,N_4363,N_4643);
nor UO_391 (O_391,N_4377,N_4101);
xnor UO_392 (O_392,N_4452,N_4437);
nand UO_393 (O_393,N_4063,N_4764);
or UO_394 (O_394,N_4034,N_4314);
nand UO_395 (O_395,N_4305,N_4163);
or UO_396 (O_396,N_4489,N_4656);
and UO_397 (O_397,N_4571,N_4317);
or UO_398 (O_398,N_4380,N_4998);
xnor UO_399 (O_399,N_4110,N_4506);
or UO_400 (O_400,N_4164,N_4354);
nor UO_401 (O_401,N_4204,N_4161);
xnor UO_402 (O_402,N_4581,N_4084);
nor UO_403 (O_403,N_4335,N_4055);
nor UO_404 (O_404,N_4904,N_4444);
nand UO_405 (O_405,N_4334,N_4970);
or UO_406 (O_406,N_4748,N_4573);
and UO_407 (O_407,N_4400,N_4919);
or UO_408 (O_408,N_4409,N_4731);
xor UO_409 (O_409,N_4770,N_4078);
nor UO_410 (O_410,N_4626,N_4916);
or UO_411 (O_411,N_4587,N_4674);
nand UO_412 (O_412,N_4679,N_4203);
and UO_413 (O_413,N_4632,N_4958);
nor UO_414 (O_414,N_4776,N_4826);
or UO_415 (O_415,N_4351,N_4926);
nand UO_416 (O_416,N_4332,N_4280);
nor UO_417 (O_417,N_4365,N_4702);
nand UO_418 (O_418,N_4129,N_4397);
nand UO_419 (O_419,N_4417,N_4574);
and UO_420 (O_420,N_4302,N_4610);
and UO_421 (O_421,N_4813,N_4196);
nor UO_422 (O_422,N_4543,N_4156);
or UO_423 (O_423,N_4706,N_4635);
xnor UO_424 (O_424,N_4920,N_4765);
nand UO_425 (O_425,N_4426,N_4235);
and UO_426 (O_426,N_4923,N_4942);
nand UO_427 (O_427,N_4735,N_4422);
nand UO_428 (O_428,N_4327,N_4901);
nand UO_429 (O_429,N_4076,N_4148);
nand UO_430 (O_430,N_4192,N_4584);
or UO_431 (O_431,N_4993,N_4382);
or UO_432 (O_432,N_4741,N_4344);
nor UO_433 (O_433,N_4802,N_4284);
and UO_434 (O_434,N_4287,N_4264);
nor UO_435 (O_435,N_4795,N_4655);
nor UO_436 (O_436,N_4193,N_4777);
nand UO_437 (O_437,N_4155,N_4859);
nand UO_438 (O_438,N_4415,N_4978);
nand UO_439 (O_439,N_4168,N_4869);
nor UO_440 (O_440,N_4064,N_4915);
and UO_441 (O_441,N_4652,N_4484);
or UO_442 (O_442,N_4230,N_4522);
nand UO_443 (O_443,N_4253,N_4454);
or UO_444 (O_444,N_4151,N_4247);
or UO_445 (O_445,N_4677,N_4931);
and UO_446 (O_446,N_4621,N_4341);
nor UO_447 (O_447,N_4398,N_4175);
and UO_448 (O_448,N_4647,N_4134);
nand UO_449 (O_449,N_4300,N_4530);
and UO_450 (O_450,N_4435,N_4283);
and UO_451 (O_451,N_4271,N_4519);
or UO_452 (O_452,N_4822,N_4725);
nand UO_453 (O_453,N_4512,N_4907);
nand UO_454 (O_454,N_4197,N_4707);
nor UO_455 (O_455,N_4049,N_4342);
nand UO_456 (O_456,N_4699,N_4631);
nand UO_457 (O_457,N_4065,N_4914);
or UO_458 (O_458,N_4547,N_4606);
nand UO_459 (O_459,N_4750,N_4139);
or UO_460 (O_460,N_4566,N_4111);
and UO_461 (O_461,N_4050,N_4578);
nor UO_462 (O_462,N_4209,N_4184);
and UO_463 (O_463,N_4274,N_4617);
nor UO_464 (O_464,N_4006,N_4618);
and UO_465 (O_465,N_4814,N_4176);
nor UO_466 (O_466,N_4987,N_4232);
and UO_467 (O_467,N_4844,N_4094);
nand UO_468 (O_468,N_4853,N_4961);
or UO_469 (O_469,N_4983,N_4407);
or UO_470 (O_470,N_4671,N_4128);
nand UO_471 (O_471,N_4953,N_4285);
or UO_472 (O_472,N_4746,N_4696);
and UO_473 (O_473,N_4596,N_4485);
or UO_474 (O_474,N_4141,N_4375);
nor UO_475 (O_475,N_4188,N_4984);
nor UO_476 (O_476,N_4037,N_4694);
nor UO_477 (O_477,N_4758,N_4995);
nand UO_478 (O_478,N_4893,N_4781);
nor UO_479 (O_479,N_4819,N_4946);
and UO_480 (O_480,N_4598,N_4254);
xor UO_481 (O_481,N_4851,N_4459);
or UO_482 (O_482,N_4088,N_4304);
and UO_483 (O_483,N_4956,N_4103);
and UO_484 (O_484,N_4242,N_4162);
nand UO_485 (O_485,N_4124,N_4206);
nor UO_486 (O_486,N_4568,N_4850);
nand UO_487 (O_487,N_4685,N_4913);
nor UO_488 (O_488,N_4681,N_4749);
nor UO_489 (O_489,N_4569,N_4544);
or UO_490 (O_490,N_4575,N_4476);
and UO_491 (O_491,N_4461,N_4804);
xnor UO_492 (O_492,N_4675,N_4760);
nor UO_493 (O_493,N_4927,N_4473);
or UO_494 (O_494,N_4879,N_4364);
and UO_495 (O_495,N_4693,N_4586);
and UO_496 (O_496,N_4945,N_4698);
xnor UO_497 (O_497,N_4069,N_4960);
or UO_498 (O_498,N_4329,N_4406);
nand UO_499 (O_499,N_4297,N_4628);
and UO_500 (O_500,N_4027,N_4833);
and UO_501 (O_501,N_4370,N_4263);
and UO_502 (O_502,N_4679,N_4528);
or UO_503 (O_503,N_4204,N_4073);
xnor UO_504 (O_504,N_4124,N_4824);
and UO_505 (O_505,N_4481,N_4711);
or UO_506 (O_506,N_4414,N_4315);
or UO_507 (O_507,N_4515,N_4985);
and UO_508 (O_508,N_4156,N_4232);
or UO_509 (O_509,N_4618,N_4297);
nand UO_510 (O_510,N_4651,N_4609);
and UO_511 (O_511,N_4204,N_4841);
or UO_512 (O_512,N_4972,N_4770);
and UO_513 (O_513,N_4832,N_4620);
nor UO_514 (O_514,N_4846,N_4473);
nor UO_515 (O_515,N_4580,N_4744);
or UO_516 (O_516,N_4804,N_4205);
and UO_517 (O_517,N_4008,N_4499);
nor UO_518 (O_518,N_4529,N_4931);
and UO_519 (O_519,N_4063,N_4214);
nand UO_520 (O_520,N_4114,N_4799);
nand UO_521 (O_521,N_4274,N_4290);
nand UO_522 (O_522,N_4893,N_4310);
xnor UO_523 (O_523,N_4882,N_4438);
or UO_524 (O_524,N_4778,N_4874);
or UO_525 (O_525,N_4126,N_4779);
nor UO_526 (O_526,N_4653,N_4000);
nand UO_527 (O_527,N_4876,N_4495);
or UO_528 (O_528,N_4005,N_4565);
nor UO_529 (O_529,N_4756,N_4072);
and UO_530 (O_530,N_4062,N_4696);
and UO_531 (O_531,N_4984,N_4094);
and UO_532 (O_532,N_4235,N_4928);
nand UO_533 (O_533,N_4418,N_4582);
and UO_534 (O_534,N_4468,N_4655);
or UO_535 (O_535,N_4122,N_4308);
and UO_536 (O_536,N_4302,N_4931);
and UO_537 (O_537,N_4970,N_4732);
xnor UO_538 (O_538,N_4210,N_4290);
or UO_539 (O_539,N_4319,N_4371);
or UO_540 (O_540,N_4425,N_4200);
and UO_541 (O_541,N_4944,N_4306);
or UO_542 (O_542,N_4473,N_4877);
or UO_543 (O_543,N_4936,N_4242);
nand UO_544 (O_544,N_4752,N_4767);
xor UO_545 (O_545,N_4154,N_4757);
or UO_546 (O_546,N_4808,N_4218);
nand UO_547 (O_547,N_4548,N_4846);
nor UO_548 (O_548,N_4033,N_4693);
nor UO_549 (O_549,N_4357,N_4119);
nand UO_550 (O_550,N_4586,N_4363);
nor UO_551 (O_551,N_4538,N_4065);
nand UO_552 (O_552,N_4403,N_4427);
and UO_553 (O_553,N_4019,N_4269);
or UO_554 (O_554,N_4850,N_4555);
xor UO_555 (O_555,N_4209,N_4067);
nand UO_556 (O_556,N_4471,N_4531);
and UO_557 (O_557,N_4662,N_4429);
nand UO_558 (O_558,N_4153,N_4675);
nand UO_559 (O_559,N_4287,N_4885);
or UO_560 (O_560,N_4298,N_4431);
or UO_561 (O_561,N_4561,N_4514);
nand UO_562 (O_562,N_4417,N_4081);
nor UO_563 (O_563,N_4224,N_4145);
and UO_564 (O_564,N_4523,N_4081);
or UO_565 (O_565,N_4394,N_4762);
or UO_566 (O_566,N_4076,N_4949);
nor UO_567 (O_567,N_4909,N_4633);
and UO_568 (O_568,N_4281,N_4267);
nor UO_569 (O_569,N_4770,N_4354);
nor UO_570 (O_570,N_4735,N_4193);
and UO_571 (O_571,N_4580,N_4929);
nand UO_572 (O_572,N_4983,N_4676);
and UO_573 (O_573,N_4100,N_4700);
and UO_574 (O_574,N_4824,N_4492);
and UO_575 (O_575,N_4589,N_4367);
or UO_576 (O_576,N_4245,N_4904);
nand UO_577 (O_577,N_4667,N_4593);
nand UO_578 (O_578,N_4962,N_4527);
or UO_579 (O_579,N_4822,N_4973);
nand UO_580 (O_580,N_4114,N_4189);
or UO_581 (O_581,N_4631,N_4799);
nand UO_582 (O_582,N_4939,N_4925);
or UO_583 (O_583,N_4700,N_4169);
or UO_584 (O_584,N_4121,N_4034);
and UO_585 (O_585,N_4236,N_4743);
nor UO_586 (O_586,N_4993,N_4386);
and UO_587 (O_587,N_4644,N_4881);
or UO_588 (O_588,N_4430,N_4235);
nand UO_589 (O_589,N_4558,N_4004);
nor UO_590 (O_590,N_4287,N_4488);
and UO_591 (O_591,N_4844,N_4346);
or UO_592 (O_592,N_4745,N_4247);
and UO_593 (O_593,N_4668,N_4136);
nor UO_594 (O_594,N_4555,N_4164);
nand UO_595 (O_595,N_4700,N_4553);
and UO_596 (O_596,N_4155,N_4667);
xor UO_597 (O_597,N_4425,N_4290);
and UO_598 (O_598,N_4937,N_4529);
nor UO_599 (O_599,N_4066,N_4118);
nor UO_600 (O_600,N_4765,N_4299);
or UO_601 (O_601,N_4602,N_4047);
or UO_602 (O_602,N_4393,N_4442);
and UO_603 (O_603,N_4166,N_4314);
xor UO_604 (O_604,N_4365,N_4382);
nand UO_605 (O_605,N_4667,N_4035);
nor UO_606 (O_606,N_4798,N_4319);
nor UO_607 (O_607,N_4420,N_4370);
nand UO_608 (O_608,N_4767,N_4349);
and UO_609 (O_609,N_4229,N_4121);
nand UO_610 (O_610,N_4940,N_4546);
nand UO_611 (O_611,N_4489,N_4814);
nor UO_612 (O_612,N_4631,N_4864);
xor UO_613 (O_613,N_4263,N_4398);
nor UO_614 (O_614,N_4992,N_4125);
nand UO_615 (O_615,N_4314,N_4810);
nor UO_616 (O_616,N_4994,N_4772);
and UO_617 (O_617,N_4287,N_4074);
or UO_618 (O_618,N_4981,N_4761);
and UO_619 (O_619,N_4367,N_4722);
and UO_620 (O_620,N_4048,N_4336);
and UO_621 (O_621,N_4878,N_4299);
nor UO_622 (O_622,N_4769,N_4448);
nand UO_623 (O_623,N_4415,N_4563);
or UO_624 (O_624,N_4491,N_4042);
and UO_625 (O_625,N_4935,N_4599);
nor UO_626 (O_626,N_4007,N_4235);
or UO_627 (O_627,N_4961,N_4951);
nand UO_628 (O_628,N_4639,N_4285);
nor UO_629 (O_629,N_4117,N_4854);
nor UO_630 (O_630,N_4583,N_4995);
or UO_631 (O_631,N_4569,N_4433);
nand UO_632 (O_632,N_4693,N_4849);
and UO_633 (O_633,N_4873,N_4013);
nor UO_634 (O_634,N_4861,N_4815);
nand UO_635 (O_635,N_4895,N_4216);
or UO_636 (O_636,N_4579,N_4100);
nor UO_637 (O_637,N_4217,N_4640);
nand UO_638 (O_638,N_4779,N_4574);
xnor UO_639 (O_639,N_4879,N_4977);
nor UO_640 (O_640,N_4239,N_4685);
nand UO_641 (O_641,N_4071,N_4850);
nand UO_642 (O_642,N_4486,N_4881);
nor UO_643 (O_643,N_4014,N_4830);
nand UO_644 (O_644,N_4128,N_4156);
and UO_645 (O_645,N_4512,N_4028);
and UO_646 (O_646,N_4827,N_4395);
nand UO_647 (O_647,N_4556,N_4635);
xor UO_648 (O_648,N_4256,N_4173);
nor UO_649 (O_649,N_4933,N_4530);
nor UO_650 (O_650,N_4721,N_4363);
xor UO_651 (O_651,N_4019,N_4744);
and UO_652 (O_652,N_4389,N_4720);
nor UO_653 (O_653,N_4176,N_4179);
nand UO_654 (O_654,N_4921,N_4712);
or UO_655 (O_655,N_4939,N_4214);
or UO_656 (O_656,N_4514,N_4101);
or UO_657 (O_657,N_4900,N_4257);
or UO_658 (O_658,N_4197,N_4290);
nand UO_659 (O_659,N_4276,N_4202);
and UO_660 (O_660,N_4392,N_4854);
and UO_661 (O_661,N_4483,N_4560);
and UO_662 (O_662,N_4423,N_4152);
nand UO_663 (O_663,N_4556,N_4463);
or UO_664 (O_664,N_4695,N_4778);
nor UO_665 (O_665,N_4825,N_4773);
nor UO_666 (O_666,N_4577,N_4491);
nor UO_667 (O_667,N_4004,N_4401);
nor UO_668 (O_668,N_4393,N_4429);
or UO_669 (O_669,N_4046,N_4661);
nand UO_670 (O_670,N_4432,N_4790);
and UO_671 (O_671,N_4634,N_4748);
or UO_672 (O_672,N_4636,N_4534);
and UO_673 (O_673,N_4764,N_4880);
and UO_674 (O_674,N_4266,N_4005);
and UO_675 (O_675,N_4877,N_4308);
nor UO_676 (O_676,N_4288,N_4120);
and UO_677 (O_677,N_4711,N_4568);
nor UO_678 (O_678,N_4024,N_4601);
or UO_679 (O_679,N_4782,N_4922);
or UO_680 (O_680,N_4630,N_4699);
nor UO_681 (O_681,N_4603,N_4940);
nand UO_682 (O_682,N_4258,N_4915);
or UO_683 (O_683,N_4910,N_4570);
nor UO_684 (O_684,N_4936,N_4261);
nor UO_685 (O_685,N_4619,N_4910);
nand UO_686 (O_686,N_4857,N_4007);
or UO_687 (O_687,N_4962,N_4511);
and UO_688 (O_688,N_4675,N_4058);
and UO_689 (O_689,N_4414,N_4148);
or UO_690 (O_690,N_4001,N_4472);
or UO_691 (O_691,N_4444,N_4288);
or UO_692 (O_692,N_4125,N_4421);
nor UO_693 (O_693,N_4192,N_4466);
nand UO_694 (O_694,N_4644,N_4535);
nor UO_695 (O_695,N_4040,N_4441);
and UO_696 (O_696,N_4635,N_4337);
xor UO_697 (O_697,N_4555,N_4861);
nor UO_698 (O_698,N_4510,N_4564);
nor UO_699 (O_699,N_4148,N_4809);
and UO_700 (O_700,N_4442,N_4710);
nand UO_701 (O_701,N_4839,N_4959);
nand UO_702 (O_702,N_4392,N_4730);
xnor UO_703 (O_703,N_4745,N_4495);
nor UO_704 (O_704,N_4262,N_4531);
nand UO_705 (O_705,N_4725,N_4391);
and UO_706 (O_706,N_4381,N_4867);
and UO_707 (O_707,N_4432,N_4169);
nand UO_708 (O_708,N_4899,N_4035);
nand UO_709 (O_709,N_4221,N_4805);
and UO_710 (O_710,N_4476,N_4707);
nor UO_711 (O_711,N_4891,N_4085);
or UO_712 (O_712,N_4383,N_4220);
nand UO_713 (O_713,N_4289,N_4287);
and UO_714 (O_714,N_4868,N_4969);
or UO_715 (O_715,N_4550,N_4903);
nor UO_716 (O_716,N_4313,N_4687);
or UO_717 (O_717,N_4491,N_4966);
nand UO_718 (O_718,N_4876,N_4507);
nor UO_719 (O_719,N_4528,N_4223);
xnor UO_720 (O_720,N_4845,N_4271);
and UO_721 (O_721,N_4818,N_4200);
nand UO_722 (O_722,N_4539,N_4581);
nor UO_723 (O_723,N_4534,N_4482);
nor UO_724 (O_724,N_4525,N_4599);
or UO_725 (O_725,N_4783,N_4814);
nand UO_726 (O_726,N_4871,N_4366);
nor UO_727 (O_727,N_4787,N_4690);
nand UO_728 (O_728,N_4100,N_4977);
or UO_729 (O_729,N_4211,N_4536);
and UO_730 (O_730,N_4654,N_4653);
nand UO_731 (O_731,N_4822,N_4645);
xor UO_732 (O_732,N_4833,N_4103);
xor UO_733 (O_733,N_4480,N_4519);
nor UO_734 (O_734,N_4673,N_4312);
xor UO_735 (O_735,N_4535,N_4742);
nand UO_736 (O_736,N_4762,N_4178);
nor UO_737 (O_737,N_4363,N_4613);
or UO_738 (O_738,N_4561,N_4610);
nor UO_739 (O_739,N_4188,N_4885);
or UO_740 (O_740,N_4900,N_4738);
and UO_741 (O_741,N_4103,N_4230);
nand UO_742 (O_742,N_4374,N_4569);
and UO_743 (O_743,N_4530,N_4435);
nor UO_744 (O_744,N_4538,N_4273);
xor UO_745 (O_745,N_4454,N_4245);
or UO_746 (O_746,N_4166,N_4427);
nor UO_747 (O_747,N_4721,N_4119);
or UO_748 (O_748,N_4775,N_4652);
nand UO_749 (O_749,N_4695,N_4077);
nor UO_750 (O_750,N_4278,N_4484);
and UO_751 (O_751,N_4220,N_4015);
or UO_752 (O_752,N_4201,N_4339);
or UO_753 (O_753,N_4750,N_4722);
xnor UO_754 (O_754,N_4100,N_4265);
and UO_755 (O_755,N_4254,N_4524);
and UO_756 (O_756,N_4546,N_4684);
nor UO_757 (O_757,N_4709,N_4969);
nand UO_758 (O_758,N_4666,N_4979);
and UO_759 (O_759,N_4244,N_4096);
or UO_760 (O_760,N_4333,N_4557);
nand UO_761 (O_761,N_4582,N_4932);
nand UO_762 (O_762,N_4588,N_4126);
or UO_763 (O_763,N_4555,N_4688);
or UO_764 (O_764,N_4168,N_4860);
nor UO_765 (O_765,N_4053,N_4817);
nand UO_766 (O_766,N_4156,N_4428);
nor UO_767 (O_767,N_4436,N_4555);
and UO_768 (O_768,N_4808,N_4416);
and UO_769 (O_769,N_4246,N_4860);
or UO_770 (O_770,N_4271,N_4539);
or UO_771 (O_771,N_4506,N_4024);
or UO_772 (O_772,N_4799,N_4632);
nand UO_773 (O_773,N_4866,N_4091);
nand UO_774 (O_774,N_4067,N_4221);
xnor UO_775 (O_775,N_4691,N_4661);
nor UO_776 (O_776,N_4465,N_4947);
or UO_777 (O_777,N_4308,N_4186);
nor UO_778 (O_778,N_4180,N_4182);
nor UO_779 (O_779,N_4979,N_4944);
xnor UO_780 (O_780,N_4695,N_4880);
and UO_781 (O_781,N_4515,N_4632);
nand UO_782 (O_782,N_4265,N_4315);
nand UO_783 (O_783,N_4633,N_4773);
and UO_784 (O_784,N_4655,N_4037);
nand UO_785 (O_785,N_4876,N_4312);
or UO_786 (O_786,N_4615,N_4076);
or UO_787 (O_787,N_4854,N_4678);
or UO_788 (O_788,N_4605,N_4199);
xor UO_789 (O_789,N_4753,N_4307);
or UO_790 (O_790,N_4721,N_4768);
or UO_791 (O_791,N_4247,N_4236);
nand UO_792 (O_792,N_4490,N_4089);
and UO_793 (O_793,N_4154,N_4897);
nand UO_794 (O_794,N_4729,N_4798);
and UO_795 (O_795,N_4043,N_4815);
xnor UO_796 (O_796,N_4711,N_4082);
or UO_797 (O_797,N_4526,N_4059);
and UO_798 (O_798,N_4363,N_4063);
or UO_799 (O_799,N_4883,N_4510);
nor UO_800 (O_800,N_4333,N_4284);
nand UO_801 (O_801,N_4202,N_4688);
xnor UO_802 (O_802,N_4258,N_4968);
nor UO_803 (O_803,N_4133,N_4961);
or UO_804 (O_804,N_4879,N_4904);
or UO_805 (O_805,N_4026,N_4317);
or UO_806 (O_806,N_4213,N_4190);
nor UO_807 (O_807,N_4785,N_4953);
and UO_808 (O_808,N_4709,N_4175);
nor UO_809 (O_809,N_4830,N_4553);
or UO_810 (O_810,N_4538,N_4680);
nand UO_811 (O_811,N_4575,N_4734);
or UO_812 (O_812,N_4856,N_4678);
nand UO_813 (O_813,N_4921,N_4517);
nand UO_814 (O_814,N_4283,N_4469);
nor UO_815 (O_815,N_4626,N_4864);
nor UO_816 (O_816,N_4599,N_4868);
and UO_817 (O_817,N_4652,N_4361);
and UO_818 (O_818,N_4189,N_4641);
nand UO_819 (O_819,N_4247,N_4685);
nor UO_820 (O_820,N_4728,N_4779);
nor UO_821 (O_821,N_4863,N_4208);
and UO_822 (O_822,N_4247,N_4754);
nand UO_823 (O_823,N_4571,N_4879);
and UO_824 (O_824,N_4832,N_4223);
nand UO_825 (O_825,N_4541,N_4306);
xor UO_826 (O_826,N_4517,N_4277);
nand UO_827 (O_827,N_4275,N_4429);
and UO_828 (O_828,N_4075,N_4747);
nor UO_829 (O_829,N_4016,N_4391);
xnor UO_830 (O_830,N_4182,N_4676);
and UO_831 (O_831,N_4445,N_4637);
and UO_832 (O_832,N_4064,N_4196);
and UO_833 (O_833,N_4667,N_4774);
nand UO_834 (O_834,N_4295,N_4129);
nor UO_835 (O_835,N_4669,N_4696);
or UO_836 (O_836,N_4616,N_4590);
xor UO_837 (O_837,N_4908,N_4664);
or UO_838 (O_838,N_4287,N_4111);
nand UO_839 (O_839,N_4834,N_4144);
nor UO_840 (O_840,N_4500,N_4293);
nand UO_841 (O_841,N_4316,N_4957);
nor UO_842 (O_842,N_4265,N_4483);
nand UO_843 (O_843,N_4504,N_4818);
nor UO_844 (O_844,N_4342,N_4362);
nor UO_845 (O_845,N_4692,N_4726);
and UO_846 (O_846,N_4629,N_4438);
or UO_847 (O_847,N_4265,N_4749);
or UO_848 (O_848,N_4690,N_4181);
nor UO_849 (O_849,N_4885,N_4800);
xnor UO_850 (O_850,N_4834,N_4431);
or UO_851 (O_851,N_4147,N_4940);
and UO_852 (O_852,N_4462,N_4717);
and UO_853 (O_853,N_4750,N_4938);
nor UO_854 (O_854,N_4857,N_4668);
and UO_855 (O_855,N_4319,N_4629);
and UO_856 (O_856,N_4096,N_4499);
nor UO_857 (O_857,N_4078,N_4874);
nand UO_858 (O_858,N_4934,N_4936);
xor UO_859 (O_859,N_4262,N_4514);
or UO_860 (O_860,N_4512,N_4429);
xor UO_861 (O_861,N_4697,N_4448);
nand UO_862 (O_862,N_4427,N_4970);
nand UO_863 (O_863,N_4711,N_4616);
xor UO_864 (O_864,N_4399,N_4780);
or UO_865 (O_865,N_4330,N_4602);
xnor UO_866 (O_866,N_4244,N_4402);
or UO_867 (O_867,N_4194,N_4905);
nor UO_868 (O_868,N_4964,N_4457);
or UO_869 (O_869,N_4668,N_4557);
nor UO_870 (O_870,N_4171,N_4085);
or UO_871 (O_871,N_4295,N_4628);
or UO_872 (O_872,N_4595,N_4025);
nor UO_873 (O_873,N_4623,N_4970);
or UO_874 (O_874,N_4332,N_4317);
or UO_875 (O_875,N_4277,N_4903);
and UO_876 (O_876,N_4665,N_4128);
and UO_877 (O_877,N_4632,N_4866);
or UO_878 (O_878,N_4977,N_4923);
nor UO_879 (O_879,N_4284,N_4421);
xnor UO_880 (O_880,N_4847,N_4995);
xor UO_881 (O_881,N_4301,N_4493);
nor UO_882 (O_882,N_4070,N_4625);
and UO_883 (O_883,N_4940,N_4264);
or UO_884 (O_884,N_4385,N_4043);
nor UO_885 (O_885,N_4308,N_4234);
or UO_886 (O_886,N_4667,N_4341);
nor UO_887 (O_887,N_4541,N_4328);
nand UO_888 (O_888,N_4487,N_4385);
nand UO_889 (O_889,N_4010,N_4139);
nand UO_890 (O_890,N_4250,N_4736);
nand UO_891 (O_891,N_4183,N_4298);
nor UO_892 (O_892,N_4823,N_4320);
nand UO_893 (O_893,N_4720,N_4376);
nand UO_894 (O_894,N_4300,N_4987);
or UO_895 (O_895,N_4957,N_4094);
and UO_896 (O_896,N_4965,N_4361);
nand UO_897 (O_897,N_4415,N_4299);
nor UO_898 (O_898,N_4941,N_4912);
nor UO_899 (O_899,N_4850,N_4139);
and UO_900 (O_900,N_4555,N_4103);
nand UO_901 (O_901,N_4799,N_4028);
xor UO_902 (O_902,N_4854,N_4725);
nor UO_903 (O_903,N_4660,N_4269);
nor UO_904 (O_904,N_4939,N_4935);
nor UO_905 (O_905,N_4774,N_4095);
and UO_906 (O_906,N_4067,N_4358);
or UO_907 (O_907,N_4669,N_4338);
nand UO_908 (O_908,N_4772,N_4781);
or UO_909 (O_909,N_4419,N_4189);
nor UO_910 (O_910,N_4484,N_4926);
and UO_911 (O_911,N_4741,N_4573);
nand UO_912 (O_912,N_4564,N_4482);
nor UO_913 (O_913,N_4382,N_4360);
and UO_914 (O_914,N_4542,N_4904);
nand UO_915 (O_915,N_4854,N_4363);
and UO_916 (O_916,N_4448,N_4904);
or UO_917 (O_917,N_4311,N_4818);
nand UO_918 (O_918,N_4676,N_4587);
nand UO_919 (O_919,N_4828,N_4728);
or UO_920 (O_920,N_4199,N_4087);
nand UO_921 (O_921,N_4385,N_4980);
nand UO_922 (O_922,N_4584,N_4351);
nor UO_923 (O_923,N_4540,N_4960);
xnor UO_924 (O_924,N_4593,N_4836);
nor UO_925 (O_925,N_4534,N_4279);
and UO_926 (O_926,N_4616,N_4815);
nor UO_927 (O_927,N_4732,N_4628);
nor UO_928 (O_928,N_4540,N_4403);
nand UO_929 (O_929,N_4448,N_4763);
or UO_930 (O_930,N_4119,N_4062);
nand UO_931 (O_931,N_4332,N_4021);
nor UO_932 (O_932,N_4897,N_4583);
nor UO_933 (O_933,N_4370,N_4379);
nand UO_934 (O_934,N_4883,N_4294);
nor UO_935 (O_935,N_4516,N_4714);
nand UO_936 (O_936,N_4922,N_4870);
and UO_937 (O_937,N_4306,N_4333);
nand UO_938 (O_938,N_4261,N_4959);
and UO_939 (O_939,N_4304,N_4560);
nor UO_940 (O_940,N_4154,N_4506);
nor UO_941 (O_941,N_4940,N_4306);
or UO_942 (O_942,N_4259,N_4263);
nand UO_943 (O_943,N_4550,N_4198);
nand UO_944 (O_944,N_4184,N_4927);
or UO_945 (O_945,N_4311,N_4145);
or UO_946 (O_946,N_4703,N_4249);
and UO_947 (O_947,N_4172,N_4096);
or UO_948 (O_948,N_4032,N_4281);
or UO_949 (O_949,N_4575,N_4389);
or UO_950 (O_950,N_4747,N_4570);
and UO_951 (O_951,N_4624,N_4772);
or UO_952 (O_952,N_4225,N_4550);
nor UO_953 (O_953,N_4336,N_4639);
xnor UO_954 (O_954,N_4135,N_4415);
nor UO_955 (O_955,N_4660,N_4373);
nor UO_956 (O_956,N_4223,N_4964);
nor UO_957 (O_957,N_4503,N_4480);
nor UO_958 (O_958,N_4742,N_4694);
or UO_959 (O_959,N_4764,N_4756);
and UO_960 (O_960,N_4876,N_4340);
nor UO_961 (O_961,N_4621,N_4052);
nor UO_962 (O_962,N_4834,N_4961);
or UO_963 (O_963,N_4025,N_4265);
xnor UO_964 (O_964,N_4944,N_4326);
and UO_965 (O_965,N_4426,N_4106);
or UO_966 (O_966,N_4654,N_4951);
and UO_967 (O_967,N_4599,N_4351);
nor UO_968 (O_968,N_4503,N_4627);
or UO_969 (O_969,N_4119,N_4938);
or UO_970 (O_970,N_4945,N_4673);
nand UO_971 (O_971,N_4270,N_4246);
nand UO_972 (O_972,N_4492,N_4929);
nand UO_973 (O_973,N_4274,N_4492);
nand UO_974 (O_974,N_4533,N_4682);
and UO_975 (O_975,N_4872,N_4413);
nor UO_976 (O_976,N_4449,N_4345);
nor UO_977 (O_977,N_4980,N_4229);
nor UO_978 (O_978,N_4348,N_4399);
and UO_979 (O_979,N_4586,N_4010);
nor UO_980 (O_980,N_4926,N_4501);
and UO_981 (O_981,N_4049,N_4073);
xnor UO_982 (O_982,N_4328,N_4527);
and UO_983 (O_983,N_4430,N_4323);
nand UO_984 (O_984,N_4910,N_4025);
nor UO_985 (O_985,N_4568,N_4116);
nand UO_986 (O_986,N_4665,N_4000);
nor UO_987 (O_987,N_4226,N_4959);
and UO_988 (O_988,N_4107,N_4564);
nor UO_989 (O_989,N_4550,N_4713);
and UO_990 (O_990,N_4287,N_4255);
or UO_991 (O_991,N_4922,N_4757);
nor UO_992 (O_992,N_4647,N_4445);
or UO_993 (O_993,N_4091,N_4369);
or UO_994 (O_994,N_4777,N_4394);
nand UO_995 (O_995,N_4212,N_4641);
nand UO_996 (O_996,N_4752,N_4051);
and UO_997 (O_997,N_4834,N_4225);
nor UO_998 (O_998,N_4162,N_4581);
or UO_999 (O_999,N_4699,N_4887);
endmodule