module basic_500_3000_500_5_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_232,In_429);
nor U1 (N_1,In_128,In_185);
nor U2 (N_2,In_245,In_34);
or U3 (N_3,In_399,In_310);
or U4 (N_4,In_2,In_167);
nor U5 (N_5,In_218,In_290);
nand U6 (N_6,In_78,In_363);
nand U7 (N_7,In_331,In_272);
nand U8 (N_8,In_327,In_396);
nor U9 (N_9,In_208,In_186);
and U10 (N_10,In_155,In_161);
nand U11 (N_11,In_472,In_19);
nand U12 (N_12,In_392,In_428);
nor U13 (N_13,In_465,In_442);
nand U14 (N_14,In_118,In_201);
xor U15 (N_15,In_261,In_190);
and U16 (N_16,In_371,In_9);
and U17 (N_17,In_26,In_336);
nand U18 (N_18,In_418,In_348);
nand U19 (N_19,In_318,In_131);
xor U20 (N_20,In_152,In_397);
nand U21 (N_21,In_460,In_87);
nand U22 (N_22,In_91,In_69);
nand U23 (N_23,In_115,In_247);
nor U24 (N_24,In_335,In_226);
or U25 (N_25,In_70,In_33);
nand U26 (N_26,In_277,In_296);
and U27 (N_27,In_469,In_352);
nand U28 (N_28,In_367,In_256);
nor U29 (N_29,In_94,In_284);
and U30 (N_30,In_306,In_324);
or U31 (N_31,In_294,In_23);
or U32 (N_32,In_433,In_426);
nand U33 (N_33,In_75,In_17);
or U34 (N_34,In_386,In_89);
nand U35 (N_35,In_188,In_171);
nor U36 (N_36,In_302,In_270);
nand U37 (N_37,In_441,In_478);
and U38 (N_38,In_140,In_410);
nand U39 (N_39,In_436,In_391);
nor U40 (N_40,In_79,In_273);
nand U41 (N_41,In_210,In_252);
xnor U42 (N_42,In_305,In_317);
or U43 (N_43,In_71,In_353);
xor U44 (N_44,In_340,In_38);
xnor U45 (N_45,In_108,In_51);
and U46 (N_46,In_445,In_46);
and U47 (N_47,In_477,In_434);
nand U48 (N_48,In_269,In_438);
nand U49 (N_49,In_159,In_239);
nand U50 (N_50,In_286,In_345);
nand U51 (N_51,In_11,In_142);
nand U52 (N_52,In_328,In_212);
nor U53 (N_53,In_405,In_113);
nand U54 (N_54,In_129,In_96);
or U55 (N_55,In_448,In_378);
or U56 (N_56,In_278,In_422);
and U57 (N_57,In_41,In_57);
xnor U58 (N_58,In_487,In_62);
and U59 (N_59,In_497,In_390);
and U60 (N_60,In_132,In_29);
or U61 (N_61,In_202,In_380);
xor U62 (N_62,In_330,In_114);
nand U63 (N_63,In_203,In_425);
nor U64 (N_64,In_287,In_65);
nand U65 (N_65,In_80,In_319);
nand U66 (N_66,In_249,In_77);
and U67 (N_67,In_309,In_407);
or U68 (N_68,In_480,In_414);
xor U69 (N_69,In_308,In_106);
nor U70 (N_70,In_147,In_137);
nand U71 (N_71,In_216,In_412);
nand U72 (N_72,In_343,In_355);
and U73 (N_73,In_104,In_116);
nand U74 (N_74,In_432,In_37);
xor U75 (N_75,In_409,In_381);
nand U76 (N_76,In_25,In_234);
nor U77 (N_77,In_431,In_35);
nor U78 (N_78,In_440,In_398);
nor U79 (N_79,In_358,In_122);
or U80 (N_80,In_344,In_27);
and U81 (N_81,In_450,In_219);
nand U82 (N_82,In_362,In_361);
or U83 (N_83,In_120,In_488);
nor U84 (N_84,In_15,In_192);
nor U85 (N_85,In_285,In_356);
or U86 (N_86,In_149,In_183);
and U87 (N_87,In_209,In_125);
and U88 (N_88,In_498,In_21);
xnor U89 (N_89,In_156,In_264);
xnor U90 (N_90,In_134,In_283);
or U91 (N_91,In_30,In_300);
nand U92 (N_92,In_6,In_389);
and U93 (N_93,In_334,In_90);
or U94 (N_94,In_45,In_101);
or U95 (N_95,In_98,In_377);
and U96 (N_96,In_292,In_10);
and U97 (N_97,In_313,In_350);
nand U98 (N_98,In_401,In_5);
or U99 (N_99,In_173,In_311);
and U100 (N_100,In_259,In_177);
and U101 (N_101,In_168,In_325);
nor U102 (N_102,In_246,In_326);
or U103 (N_103,In_424,In_233);
or U104 (N_104,In_315,In_13);
and U105 (N_105,In_242,In_262);
and U106 (N_106,In_48,In_102);
nand U107 (N_107,In_107,In_144);
nand U108 (N_108,In_402,In_342);
nor U109 (N_109,In_241,In_56);
xor U110 (N_110,In_320,In_126);
and U111 (N_111,In_307,In_314);
nand U112 (N_112,In_194,In_179);
nand U113 (N_113,In_473,In_332);
nor U114 (N_114,In_254,In_109);
nand U115 (N_115,In_105,In_265);
nand U116 (N_116,In_281,In_206);
nor U117 (N_117,In_298,In_421);
or U118 (N_118,In_54,In_258);
or U119 (N_119,In_240,In_267);
and U120 (N_120,In_112,In_133);
or U121 (N_121,In_160,In_427);
nor U122 (N_122,In_395,In_484);
or U123 (N_123,In_150,In_63);
or U124 (N_124,In_76,In_388);
or U125 (N_125,In_141,In_375);
or U126 (N_126,In_467,In_251);
or U127 (N_127,In_64,In_490);
nor U128 (N_128,In_153,In_175);
and U129 (N_129,In_151,In_165);
nor U130 (N_130,In_82,In_146);
nor U131 (N_131,In_213,In_143);
nand U132 (N_132,In_374,In_387);
nor U133 (N_133,In_458,In_333);
nor U134 (N_134,In_135,In_403);
xor U135 (N_135,In_238,In_36);
nor U136 (N_136,In_73,In_124);
or U137 (N_137,In_176,In_408);
nor U138 (N_138,In_92,In_139);
nor U139 (N_139,In_288,In_215);
nor U140 (N_140,In_385,In_172);
nand U141 (N_141,In_279,In_293);
xor U142 (N_142,In_338,In_466);
and U143 (N_143,In_457,In_379);
and U144 (N_144,In_86,In_468);
or U145 (N_145,In_282,In_66);
or U146 (N_146,In_485,In_14);
nor U147 (N_147,In_164,In_236);
or U148 (N_148,In_220,In_1);
nor U149 (N_149,In_280,In_406);
and U150 (N_150,In_44,In_103);
or U151 (N_151,In_68,In_205);
xor U152 (N_152,In_244,In_456);
or U153 (N_153,In_323,In_299);
or U154 (N_154,In_470,In_148);
nand U155 (N_155,In_83,In_174);
nand U156 (N_156,In_276,In_42);
or U157 (N_157,In_483,In_154);
nor U158 (N_158,In_214,In_28);
or U159 (N_159,In_235,In_72);
and U160 (N_160,In_437,In_453);
nor U161 (N_161,In_260,In_291);
or U162 (N_162,In_455,In_257);
and U163 (N_163,In_464,In_184);
nor U164 (N_164,In_304,In_158);
nor U165 (N_165,In_346,In_354);
and U166 (N_166,In_170,In_357);
nand U167 (N_167,In_95,In_400);
nand U168 (N_168,In_50,In_61);
or U169 (N_169,In_474,In_372);
or U170 (N_170,In_84,In_248);
nand U171 (N_171,In_3,In_180);
or U172 (N_172,In_60,In_222);
or U173 (N_173,In_223,In_74);
and U174 (N_174,In_32,In_47);
nor U175 (N_175,In_169,In_16);
and U176 (N_176,In_369,In_221);
nand U177 (N_177,In_393,In_435);
or U178 (N_178,In_494,In_49);
nor U179 (N_179,In_446,In_138);
nand U180 (N_180,In_163,In_0);
nand U181 (N_181,In_253,In_471);
nor U182 (N_182,In_198,In_491);
xor U183 (N_183,In_419,In_119);
nor U184 (N_184,In_199,In_12);
nor U185 (N_185,In_187,In_20);
or U186 (N_186,In_443,In_200);
nor U187 (N_187,In_423,In_97);
and U188 (N_188,In_364,In_341);
nor U189 (N_189,In_211,In_394);
nor U190 (N_190,In_376,In_439);
and U191 (N_191,In_263,In_452);
and U192 (N_192,In_495,In_136);
nand U193 (N_193,In_237,In_365);
xor U194 (N_194,In_373,In_40);
nand U195 (N_195,In_266,In_420);
and U196 (N_196,In_415,In_181);
and U197 (N_197,In_382,In_271);
and U198 (N_198,In_417,In_322);
nand U199 (N_199,In_444,In_43);
or U200 (N_200,In_339,In_289);
nor U201 (N_201,In_255,In_8);
nor U202 (N_202,In_110,In_227);
and U203 (N_203,In_197,In_100);
nor U204 (N_204,In_461,In_88);
and U205 (N_205,In_231,In_349);
or U206 (N_206,In_360,In_193);
nor U207 (N_207,In_430,In_59);
nand U208 (N_208,In_479,In_204);
or U209 (N_209,In_111,In_250);
and U210 (N_210,In_321,In_81);
nand U211 (N_211,In_195,In_225);
nor U212 (N_212,In_24,In_22);
nor U213 (N_213,In_4,In_127);
xnor U214 (N_214,In_295,In_99);
nor U215 (N_215,In_217,In_53);
nor U216 (N_216,In_85,In_123);
and U217 (N_217,In_493,In_145);
nor U218 (N_218,In_454,In_275);
or U219 (N_219,In_476,In_301);
xor U220 (N_220,In_351,In_475);
or U221 (N_221,In_93,In_462);
nor U222 (N_222,In_368,In_481);
or U223 (N_223,In_359,In_383);
nor U224 (N_224,In_224,In_18);
and U225 (N_225,In_182,In_312);
nand U226 (N_226,In_121,In_189);
nor U227 (N_227,In_39,In_303);
or U228 (N_228,In_347,In_130);
and U229 (N_229,In_447,In_411);
or U230 (N_230,In_463,In_162);
nor U231 (N_231,In_230,In_166);
and U232 (N_232,In_117,In_370);
or U233 (N_233,In_7,In_496);
nand U234 (N_234,In_191,In_486);
nand U235 (N_235,In_52,In_297);
nand U236 (N_236,In_413,In_499);
and U237 (N_237,In_196,In_451);
nand U238 (N_238,In_243,In_268);
nand U239 (N_239,In_157,In_274);
and U240 (N_240,In_489,In_329);
nor U241 (N_241,In_67,In_55);
nand U242 (N_242,In_178,In_384);
or U243 (N_243,In_207,In_31);
nor U244 (N_244,In_449,In_58);
xnor U245 (N_245,In_228,In_316);
xor U246 (N_246,In_416,In_366);
nand U247 (N_247,In_492,In_337);
nor U248 (N_248,In_229,In_459);
xnor U249 (N_249,In_404,In_482);
nand U250 (N_250,In_406,In_39);
nor U251 (N_251,In_83,In_59);
and U252 (N_252,In_71,In_474);
xnor U253 (N_253,In_360,In_380);
and U254 (N_254,In_342,In_275);
and U255 (N_255,In_146,In_325);
or U256 (N_256,In_39,In_399);
nor U257 (N_257,In_80,In_71);
or U258 (N_258,In_493,In_393);
nor U259 (N_259,In_280,In_135);
nand U260 (N_260,In_98,In_225);
or U261 (N_261,In_474,In_287);
or U262 (N_262,In_117,In_417);
and U263 (N_263,In_367,In_182);
nand U264 (N_264,In_11,In_460);
nor U265 (N_265,In_349,In_392);
and U266 (N_266,In_303,In_376);
nor U267 (N_267,In_313,In_302);
xnor U268 (N_268,In_240,In_442);
and U269 (N_269,In_137,In_410);
and U270 (N_270,In_474,In_377);
nand U271 (N_271,In_68,In_493);
nand U272 (N_272,In_154,In_418);
nand U273 (N_273,In_415,In_98);
and U274 (N_274,In_56,In_369);
xor U275 (N_275,In_79,In_378);
and U276 (N_276,In_429,In_417);
nand U277 (N_277,In_137,In_308);
nand U278 (N_278,In_293,In_274);
and U279 (N_279,In_149,In_405);
nand U280 (N_280,In_43,In_462);
and U281 (N_281,In_290,In_73);
nand U282 (N_282,In_495,In_272);
or U283 (N_283,In_90,In_402);
nand U284 (N_284,In_85,In_335);
xor U285 (N_285,In_311,In_47);
nor U286 (N_286,In_124,In_18);
nand U287 (N_287,In_447,In_261);
and U288 (N_288,In_162,In_267);
and U289 (N_289,In_491,In_273);
or U290 (N_290,In_393,In_53);
nor U291 (N_291,In_251,In_248);
nor U292 (N_292,In_124,In_250);
or U293 (N_293,In_353,In_160);
nor U294 (N_294,In_415,In_174);
nor U295 (N_295,In_464,In_254);
or U296 (N_296,In_344,In_53);
nand U297 (N_297,In_28,In_232);
and U298 (N_298,In_121,In_147);
nor U299 (N_299,In_31,In_223);
nand U300 (N_300,In_224,In_252);
or U301 (N_301,In_189,In_226);
nor U302 (N_302,In_166,In_201);
nor U303 (N_303,In_241,In_103);
or U304 (N_304,In_170,In_280);
nand U305 (N_305,In_437,In_487);
xnor U306 (N_306,In_37,In_308);
nor U307 (N_307,In_396,In_74);
xnor U308 (N_308,In_265,In_453);
xnor U309 (N_309,In_195,In_162);
nor U310 (N_310,In_400,In_485);
xnor U311 (N_311,In_350,In_118);
or U312 (N_312,In_202,In_420);
and U313 (N_313,In_83,In_380);
and U314 (N_314,In_426,In_400);
nand U315 (N_315,In_308,In_267);
nand U316 (N_316,In_108,In_68);
and U317 (N_317,In_49,In_343);
and U318 (N_318,In_375,In_41);
xor U319 (N_319,In_113,In_218);
nand U320 (N_320,In_446,In_401);
nor U321 (N_321,In_360,In_226);
and U322 (N_322,In_452,In_364);
nand U323 (N_323,In_147,In_397);
nand U324 (N_324,In_321,In_450);
xnor U325 (N_325,In_272,In_424);
xor U326 (N_326,In_254,In_244);
nand U327 (N_327,In_73,In_422);
or U328 (N_328,In_444,In_393);
and U329 (N_329,In_499,In_86);
nor U330 (N_330,In_243,In_203);
nand U331 (N_331,In_62,In_472);
xor U332 (N_332,In_433,In_20);
and U333 (N_333,In_134,In_392);
xnor U334 (N_334,In_156,In_254);
or U335 (N_335,In_360,In_278);
and U336 (N_336,In_150,In_316);
and U337 (N_337,In_131,In_345);
xnor U338 (N_338,In_492,In_192);
and U339 (N_339,In_480,In_39);
or U340 (N_340,In_377,In_470);
and U341 (N_341,In_251,In_196);
nor U342 (N_342,In_353,In_95);
and U343 (N_343,In_32,In_327);
nand U344 (N_344,In_44,In_166);
or U345 (N_345,In_307,In_265);
nand U346 (N_346,In_297,In_293);
nor U347 (N_347,In_465,In_284);
nand U348 (N_348,In_312,In_219);
or U349 (N_349,In_364,In_406);
and U350 (N_350,In_243,In_301);
or U351 (N_351,In_148,In_262);
and U352 (N_352,In_47,In_400);
xnor U353 (N_353,In_120,In_231);
nor U354 (N_354,In_115,In_111);
nor U355 (N_355,In_82,In_78);
or U356 (N_356,In_474,In_97);
and U357 (N_357,In_239,In_227);
and U358 (N_358,In_408,In_221);
nand U359 (N_359,In_290,In_350);
or U360 (N_360,In_421,In_92);
or U361 (N_361,In_254,In_286);
nand U362 (N_362,In_438,In_335);
nor U363 (N_363,In_162,In_202);
nand U364 (N_364,In_62,In_280);
nand U365 (N_365,In_236,In_205);
xnor U366 (N_366,In_212,In_109);
nor U367 (N_367,In_66,In_369);
or U368 (N_368,In_224,In_223);
or U369 (N_369,In_88,In_31);
or U370 (N_370,In_92,In_164);
and U371 (N_371,In_489,In_31);
nand U372 (N_372,In_329,In_246);
and U373 (N_373,In_228,In_272);
nand U374 (N_374,In_429,In_139);
and U375 (N_375,In_160,In_87);
nand U376 (N_376,In_185,In_307);
and U377 (N_377,In_21,In_422);
and U378 (N_378,In_469,In_199);
nor U379 (N_379,In_421,In_112);
or U380 (N_380,In_196,In_248);
nand U381 (N_381,In_29,In_36);
nand U382 (N_382,In_83,In_283);
or U383 (N_383,In_8,In_80);
nand U384 (N_384,In_323,In_194);
nor U385 (N_385,In_110,In_121);
nor U386 (N_386,In_116,In_496);
xor U387 (N_387,In_394,In_152);
or U388 (N_388,In_180,In_161);
nand U389 (N_389,In_17,In_66);
nor U390 (N_390,In_91,In_264);
nor U391 (N_391,In_332,In_137);
nand U392 (N_392,In_53,In_159);
or U393 (N_393,In_39,In_144);
nand U394 (N_394,In_226,In_451);
xnor U395 (N_395,In_281,In_395);
xnor U396 (N_396,In_99,In_439);
and U397 (N_397,In_485,In_214);
and U398 (N_398,In_478,In_310);
nor U399 (N_399,In_129,In_0);
and U400 (N_400,In_334,In_22);
nor U401 (N_401,In_42,In_252);
or U402 (N_402,In_12,In_167);
or U403 (N_403,In_211,In_255);
nand U404 (N_404,In_448,In_164);
or U405 (N_405,In_5,In_194);
or U406 (N_406,In_411,In_118);
nor U407 (N_407,In_179,In_293);
and U408 (N_408,In_187,In_403);
nand U409 (N_409,In_375,In_346);
nor U410 (N_410,In_390,In_391);
or U411 (N_411,In_150,In_460);
or U412 (N_412,In_293,In_191);
nand U413 (N_413,In_98,In_134);
or U414 (N_414,In_221,In_4);
or U415 (N_415,In_444,In_2);
or U416 (N_416,In_309,In_466);
xnor U417 (N_417,In_208,In_46);
or U418 (N_418,In_466,In_139);
nor U419 (N_419,In_359,In_68);
xnor U420 (N_420,In_76,In_410);
or U421 (N_421,In_161,In_154);
nor U422 (N_422,In_2,In_355);
nand U423 (N_423,In_188,In_182);
nand U424 (N_424,In_492,In_417);
or U425 (N_425,In_134,In_470);
nor U426 (N_426,In_0,In_393);
nor U427 (N_427,In_279,In_222);
and U428 (N_428,In_243,In_131);
nor U429 (N_429,In_297,In_389);
and U430 (N_430,In_455,In_26);
nor U431 (N_431,In_266,In_301);
and U432 (N_432,In_157,In_56);
nor U433 (N_433,In_387,In_444);
and U434 (N_434,In_14,In_72);
and U435 (N_435,In_289,In_124);
or U436 (N_436,In_23,In_462);
nor U437 (N_437,In_324,In_124);
nor U438 (N_438,In_75,In_135);
or U439 (N_439,In_212,In_486);
xor U440 (N_440,In_223,In_436);
xor U441 (N_441,In_372,In_266);
and U442 (N_442,In_395,In_198);
nand U443 (N_443,In_83,In_480);
nand U444 (N_444,In_159,In_413);
nor U445 (N_445,In_497,In_163);
nor U446 (N_446,In_117,In_404);
nand U447 (N_447,In_166,In_9);
xnor U448 (N_448,In_426,In_476);
and U449 (N_449,In_431,In_495);
xnor U450 (N_450,In_36,In_335);
or U451 (N_451,In_112,In_288);
nand U452 (N_452,In_389,In_31);
nor U453 (N_453,In_416,In_106);
or U454 (N_454,In_215,In_65);
xnor U455 (N_455,In_99,In_286);
or U456 (N_456,In_27,In_339);
or U457 (N_457,In_263,In_443);
nor U458 (N_458,In_394,In_492);
nor U459 (N_459,In_373,In_374);
or U460 (N_460,In_301,In_252);
nand U461 (N_461,In_279,In_35);
nand U462 (N_462,In_138,In_121);
and U463 (N_463,In_430,In_73);
nand U464 (N_464,In_294,In_65);
and U465 (N_465,In_150,In_184);
nor U466 (N_466,In_399,In_298);
nand U467 (N_467,In_227,In_89);
or U468 (N_468,In_86,In_124);
or U469 (N_469,In_202,In_41);
nor U470 (N_470,In_427,In_492);
or U471 (N_471,In_155,In_257);
or U472 (N_472,In_437,In_327);
or U473 (N_473,In_421,In_427);
or U474 (N_474,In_111,In_316);
or U475 (N_475,In_215,In_99);
nor U476 (N_476,In_25,In_463);
nor U477 (N_477,In_469,In_306);
nor U478 (N_478,In_11,In_108);
nand U479 (N_479,In_475,In_444);
and U480 (N_480,In_386,In_334);
nand U481 (N_481,In_168,In_140);
and U482 (N_482,In_85,In_168);
nor U483 (N_483,In_84,In_443);
or U484 (N_484,In_172,In_87);
and U485 (N_485,In_358,In_468);
nor U486 (N_486,In_205,In_93);
nand U487 (N_487,In_447,In_74);
nand U488 (N_488,In_42,In_281);
and U489 (N_489,In_1,In_118);
nand U490 (N_490,In_109,In_87);
nor U491 (N_491,In_27,In_278);
or U492 (N_492,In_145,In_284);
nor U493 (N_493,In_180,In_150);
nand U494 (N_494,In_414,In_206);
and U495 (N_495,In_297,In_151);
nor U496 (N_496,In_465,In_128);
nand U497 (N_497,In_281,In_228);
and U498 (N_498,In_326,In_378);
nand U499 (N_499,In_193,In_283);
and U500 (N_500,In_444,In_472);
or U501 (N_501,In_314,In_285);
or U502 (N_502,In_112,In_458);
nor U503 (N_503,In_240,In_200);
and U504 (N_504,In_19,In_388);
nor U505 (N_505,In_218,In_141);
or U506 (N_506,In_382,In_355);
or U507 (N_507,In_113,In_497);
xor U508 (N_508,In_115,In_55);
and U509 (N_509,In_243,In_2);
or U510 (N_510,In_14,In_404);
or U511 (N_511,In_386,In_470);
and U512 (N_512,In_106,In_45);
or U513 (N_513,In_218,In_447);
and U514 (N_514,In_435,In_316);
and U515 (N_515,In_498,In_220);
nand U516 (N_516,In_126,In_400);
or U517 (N_517,In_451,In_271);
nor U518 (N_518,In_194,In_338);
or U519 (N_519,In_177,In_499);
nand U520 (N_520,In_308,In_401);
or U521 (N_521,In_272,In_432);
nand U522 (N_522,In_392,In_378);
and U523 (N_523,In_117,In_218);
nor U524 (N_524,In_221,In_479);
and U525 (N_525,In_23,In_126);
or U526 (N_526,In_250,In_229);
and U527 (N_527,In_20,In_176);
xor U528 (N_528,In_274,In_379);
nand U529 (N_529,In_39,In_325);
and U530 (N_530,In_448,In_288);
and U531 (N_531,In_198,In_458);
and U532 (N_532,In_294,In_431);
nor U533 (N_533,In_170,In_239);
or U534 (N_534,In_108,In_111);
and U535 (N_535,In_391,In_185);
or U536 (N_536,In_115,In_324);
nor U537 (N_537,In_261,In_198);
nor U538 (N_538,In_342,In_400);
or U539 (N_539,In_95,In_375);
and U540 (N_540,In_375,In_203);
and U541 (N_541,In_86,In_402);
nand U542 (N_542,In_0,In_338);
or U543 (N_543,In_309,In_449);
and U544 (N_544,In_242,In_16);
or U545 (N_545,In_279,In_0);
and U546 (N_546,In_249,In_30);
nand U547 (N_547,In_482,In_288);
or U548 (N_548,In_358,In_370);
nor U549 (N_549,In_24,In_458);
nor U550 (N_550,In_75,In_386);
nand U551 (N_551,In_453,In_358);
xnor U552 (N_552,In_75,In_421);
and U553 (N_553,In_451,In_37);
or U554 (N_554,In_458,In_295);
or U555 (N_555,In_378,In_204);
nor U556 (N_556,In_431,In_430);
nor U557 (N_557,In_39,In_17);
nor U558 (N_558,In_331,In_273);
nand U559 (N_559,In_204,In_321);
nor U560 (N_560,In_172,In_320);
nor U561 (N_561,In_202,In_363);
nand U562 (N_562,In_286,In_491);
or U563 (N_563,In_286,In_93);
nand U564 (N_564,In_230,In_194);
nand U565 (N_565,In_411,In_351);
or U566 (N_566,In_265,In_74);
nand U567 (N_567,In_403,In_218);
nand U568 (N_568,In_366,In_40);
and U569 (N_569,In_142,In_389);
and U570 (N_570,In_205,In_91);
nor U571 (N_571,In_484,In_266);
and U572 (N_572,In_14,In_314);
nor U573 (N_573,In_353,In_328);
and U574 (N_574,In_458,In_401);
or U575 (N_575,In_492,In_203);
nor U576 (N_576,In_71,In_340);
nor U577 (N_577,In_83,In_163);
and U578 (N_578,In_249,In_225);
or U579 (N_579,In_492,In_404);
and U580 (N_580,In_484,In_32);
and U581 (N_581,In_241,In_226);
nor U582 (N_582,In_166,In_274);
or U583 (N_583,In_26,In_64);
nand U584 (N_584,In_352,In_175);
nor U585 (N_585,In_189,In_225);
nand U586 (N_586,In_494,In_405);
and U587 (N_587,In_419,In_225);
or U588 (N_588,In_124,In_83);
or U589 (N_589,In_405,In_150);
nand U590 (N_590,In_20,In_247);
and U591 (N_591,In_24,In_58);
nand U592 (N_592,In_96,In_212);
xnor U593 (N_593,In_241,In_335);
nor U594 (N_594,In_101,In_499);
or U595 (N_595,In_92,In_425);
nand U596 (N_596,In_336,In_34);
nor U597 (N_597,In_94,In_101);
and U598 (N_598,In_26,In_252);
nand U599 (N_599,In_11,In_127);
and U600 (N_600,N_0,N_125);
or U601 (N_601,N_288,N_88);
nand U602 (N_602,N_514,N_593);
nand U603 (N_603,N_369,N_383);
or U604 (N_604,N_447,N_375);
and U605 (N_605,N_431,N_192);
nand U606 (N_606,N_417,N_235);
nand U607 (N_607,N_79,N_212);
nand U608 (N_608,N_435,N_409);
nor U609 (N_609,N_584,N_84);
nand U610 (N_610,N_489,N_199);
nor U611 (N_611,N_393,N_534);
nand U612 (N_612,N_130,N_58);
nor U613 (N_613,N_213,N_239);
nand U614 (N_614,N_585,N_226);
xor U615 (N_615,N_492,N_7);
and U616 (N_616,N_330,N_372);
nand U617 (N_617,N_452,N_547);
nor U618 (N_618,N_538,N_385);
nor U619 (N_619,N_15,N_362);
nand U620 (N_620,N_578,N_19);
nand U621 (N_621,N_497,N_532);
or U622 (N_622,N_165,N_371);
or U623 (N_623,N_341,N_530);
and U624 (N_624,N_1,N_563);
nand U625 (N_625,N_451,N_574);
and U626 (N_626,N_386,N_461);
nand U627 (N_627,N_21,N_243);
and U628 (N_628,N_307,N_579);
xnor U629 (N_629,N_303,N_396);
or U630 (N_630,N_129,N_367);
and U631 (N_631,N_16,N_140);
and U632 (N_632,N_536,N_250);
and U633 (N_633,N_528,N_517);
nor U634 (N_634,N_123,N_177);
and U635 (N_635,N_121,N_221);
nand U636 (N_636,N_304,N_397);
xor U637 (N_637,N_413,N_315);
nor U638 (N_638,N_388,N_107);
xor U639 (N_639,N_214,N_160);
nand U640 (N_640,N_496,N_73);
nand U641 (N_641,N_117,N_311);
or U642 (N_642,N_436,N_398);
or U643 (N_643,N_201,N_249);
and U644 (N_644,N_460,N_470);
nor U645 (N_645,N_483,N_169);
nor U646 (N_646,N_599,N_93);
or U647 (N_647,N_18,N_64);
nand U648 (N_648,N_523,N_332);
or U649 (N_649,N_429,N_335);
or U650 (N_650,N_159,N_96);
and U651 (N_651,N_309,N_175);
nor U652 (N_652,N_289,N_402);
nand U653 (N_653,N_72,N_317);
and U654 (N_654,N_180,N_487);
nand U655 (N_655,N_109,N_52);
nor U656 (N_656,N_83,N_441);
xnor U657 (N_657,N_531,N_268);
xnor U658 (N_658,N_66,N_455);
or U659 (N_659,N_522,N_32);
and U660 (N_660,N_596,N_568);
nand U661 (N_661,N_331,N_529);
or U662 (N_662,N_459,N_89);
or U663 (N_663,N_105,N_551);
nand U664 (N_664,N_525,N_555);
xnor U665 (N_665,N_406,N_296);
or U666 (N_666,N_27,N_422);
and U667 (N_667,N_493,N_294);
nand U668 (N_668,N_61,N_333);
or U669 (N_669,N_374,N_527);
xnor U670 (N_670,N_395,N_265);
nand U671 (N_671,N_301,N_427);
nor U672 (N_672,N_586,N_518);
nand U673 (N_673,N_370,N_182);
nor U674 (N_674,N_572,N_118);
nor U675 (N_675,N_245,N_173);
nor U676 (N_676,N_548,N_486);
or U677 (N_677,N_399,N_44);
and U678 (N_678,N_465,N_34);
and U679 (N_679,N_69,N_188);
nand U680 (N_680,N_229,N_195);
or U681 (N_681,N_325,N_98);
and U682 (N_682,N_198,N_426);
xor U683 (N_683,N_379,N_102);
or U684 (N_684,N_25,N_51);
nand U685 (N_685,N_446,N_276);
or U686 (N_686,N_485,N_170);
and U687 (N_687,N_113,N_368);
nand U688 (N_688,N_4,N_166);
nor U689 (N_689,N_209,N_9);
nand U690 (N_690,N_473,N_207);
and U691 (N_691,N_230,N_78);
and U692 (N_692,N_206,N_3);
nor U693 (N_693,N_122,N_306);
or U694 (N_694,N_280,N_457);
or U695 (N_695,N_478,N_127);
nor U696 (N_696,N_222,N_266);
nor U697 (N_697,N_236,N_167);
nand U698 (N_698,N_546,N_231);
or U699 (N_699,N_591,N_91);
or U700 (N_700,N_274,N_410);
xor U701 (N_701,N_87,N_225);
nand U702 (N_702,N_381,N_139);
or U703 (N_703,N_420,N_277);
nor U704 (N_704,N_310,N_285);
and U705 (N_705,N_543,N_100);
nor U706 (N_706,N_53,N_158);
nand U707 (N_707,N_128,N_11);
nor U708 (N_708,N_503,N_146);
or U709 (N_709,N_434,N_554);
nor U710 (N_710,N_124,N_344);
nand U711 (N_711,N_187,N_71);
nand U712 (N_712,N_394,N_35);
nand U713 (N_713,N_141,N_445);
nand U714 (N_714,N_498,N_358);
or U715 (N_715,N_200,N_500);
nand U716 (N_716,N_81,N_38);
nor U717 (N_717,N_558,N_55);
nand U718 (N_718,N_537,N_544);
and U719 (N_719,N_570,N_24);
nor U720 (N_720,N_90,N_161);
nor U721 (N_721,N_490,N_321);
nand U722 (N_722,N_194,N_580);
nor U723 (N_723,N_407,N_36);
and U724 (N_724,N_464,N_346);
or U725 (N_725,N_111,N_261);
and U726 (N_726,N_556,N_152);
nand U727 (N_727,N_168,N_360);
nor U728 (N_728,N_26,N_495);
and U729 (N_729,N_10,N_504);
nor U730 (N_730,N_244,N_132);
xor U731 (N_731,N_308,N_373);
xnor U732 (N_732,N_219,N_519);
and U733 (N_733,N_502,N_279);
or U734 (N_734,N_463,N_562);
or U735 (N_735,N_2,N_106);
nor U736 (N_736,N_415,N_475);
nand U737 (N_737,N_252,N_193);
xor U738 (N_738,N_582,N_184);
nor U739 (N_739,N_322,N_233);
xnor U740 (N_740,N_454,N_238);
nor U741 (N_741,N_75,N_5);
and U742 (N_742,N_509,N_271);
nor U743 (N_743,N_510,N_550);
nand U744 (N_744,N_458,N_23);
nand U745 (N_745,N_20,N_217);
and U746 (N_746,N_218,N_86);
and U747 (N_747,N_43,N_95);
xnor U748 (N_748,N_355,N_576);
nand U749 (N_749,N_380,N_376);
xor U750 (N_750,N_389,N_92);
nand U751 (N_751,N_466,N_46);
nand U752 (N_752,N_6,N_133);
and U753 (N_753,N_232,N_126);
and U754 (N_754,N_506,N_357);
nand U755 (N_755,N_253,N_392);
xnor U756 (N_756,N_312,N_539);
nand U757 (N_757,N_101,N_540);
or U758 (N_758,N_324,N_31);
or U759 (N_759,N_505,N_155);
nor U760 (N_760,N_45,N_248);
nand U761 (N_761,N_97,N_571);
and U762 (N_762,N_224,N_40);
or U763 (N_763,N_197,N_143);
xor U764 (N_764,N_208,N_488);
or U765 (N_765,N_284,N_247);
or U766 (N_766,N_8,N_33);
nand U767 (N_767,N_14,N_80);
nor U768 (N_768,N_354,N_255);
nand U769 (N_769,N_329,N_147);
nor U770 (N_770,N_264,N_144);
nor U771 (N_771,N_428,N_150);
xor U772 (N_772,N_202,N_120);
nor U773 (N_773,N_366,N_211);
and U774 (N_774,N_104,N_468);
and U775 (N_775,N_577,N_382);
or U776 (N_776,N_82,N_553);
nand U777 (N_777,N_293,N_482);
nor U778 (N_778,N_450,N_178);
and U779 (N_779,N_291,N_153);
or U780 (N_780,N_587,N_67);
nor U781 (N_781,N_569,N_328);
nand U782 (N_782,N_340,N_237);
and U783 (N_783,N_94,N_12);
or U784 (N_784,N_275,N_37);
and U785 (N_785,N_416,N_444);
and U786 (N_786,N_13,N_583);
or U787 (N_787,N_251,N_305);
nor U788 (N_788,N_56,N_60);
nor U789 (N_789,N_48,N_323);
nor U790 (N_790,N_287,N_292);
nand U791 (N_791,N_575,N_240);
nand U792 (N_792,N_403,N_592);
nor U793 (N_793,N_316,N_598);
and U794 (N_794,N_430,N_353);
nor U795 (N_795,N_507,N_438);
nand U796 (N_796,N_347,N_561);
or U797 (N_797,N_295,N_419);
nand U798 (N_798,N_350,N_270);
or U799 (N_799,N_414,N_99);
and U800 (N_800,N_164,N_50);
or U801 (N_801,N_28,N_516);
nor U802 (N_802,N_565,N_110);
nand U803 (N_803,N_131,N_390);
nor U804 (N_804,N_508,N_318);
and U805 (N_805,N_471,N_391);
nand U806 (N_806,N_480,N_216);
and U807 (N_807,N_400,N_595);
nand U808 (N_808,N_282,N_228);
nor U809 (N_809,N_183,N_137);
and U810 (N_810,N_511,N_343);
nor U811 (N_811,N_545,N_520);
nor U812 (N_812,N_549,N_559);
and U813 (N_813,N_361,N_203);
nand U814 (N_814,N_521,N_149);
nand U815 (N_815,N_112,N_186);
or U816 (N_816,N_437,N_63);
nand U817 (N_817,N_448,N_242);
and U818 (N_818,N_567,N_334);
and U819 (N_819,N_439,N_42);
and U820 (N_820,N_283,N_77);
nor U821 (N_821,N_472,N_210);
and U822 (N_822,N_338,N_138);
and U823 (N_823,N_566,N_57);
or U824 (N_824,N_220,N_345);
xor U825 (N_825,N_462,N_474);
nor U826 (N_826,N_281,N_134);
or U827 (N_827,N_467,N_154);
or U828 (N_828,N_30,N_533);
and U829 (N_829,N_246,N_352);
or U830 (N_830,N_425,N_541);
nand U831 (N_831,N_589,N_564);
nor U832 (N_832,N_313,N_257);
or U833 (N_833,N_223,N_39);
or U834 (N_834,N_476,N_481);
and U835 (N_835,N_515,N_234);
xor U836 (N_836,N_171,N_442);
xnor U837 (N_837,N_254,N_359);
or U838 (N_838,N_114,N_387);
nand U839 (N_839,N_349,N_456);
and U840 (N_840,N_286,N_542);
nor U841 (N_841,N_267,N_174);
nor U842 (N_842,N_378,N_479);
or U843 (N_843,N_588,N_262);
nor U844 (N_844,N_557,N_17);
and U845 (N_845,N_172,N_260);
xor U846 (N_846,N_119,N_302);
or U847 (N_847,N_115,N_421);
and U848 (N_848,N_342,N_594);
nand U849 (N_849,N_408,N_103);
nor U850 (N_850,N_157,N_298);
nand U851 (N_851,N_484,N_142);
nand U852 (N_852,N_499,N_401);
and U853 (N_853,N_189,N_65);
and U854 (N_854,N_405,N_29);
nor U855 (N_855,N_526,N_59);
nand U856 (N_856,N_162,N_560);
nand U857 (N_857,N_22,N_336);
nor U858 (N_858,N_449,N_116);
or U859 (N_859,N_70,N_524);
xor U860 (N_860,N_76,N_258);
nor U861 (N_861,N_319,N_440);
or U862 (N_862,N_227,N_299);
or U863 (N_863,N_573,N_263);
nand U864 (N_864,N_54,N_156);
and U865 (N_865,N_552,N_163);
or U866 (N_866,N_513,N_41);
or U867 (N_867,N_535,N_337);
or U868 (N_868,N_185,N_49);
nor U869 (N_869,N_85,N_364);
or U870 (N_870,N_151,N_453);
nand U871 (N_871,N_377,N_365);
xor U872 (N_872,N_590,N_196);
xor U873 (N_873,N_269,N_581);
xor U874 (N_874,N_363,N_314);
xnor U875 (N_875,N_300,N_181);
and U876 (N_876,N_204,N_418);
xor U877 (N_877,N_491,N_327);
nor U878 (N_878,N_411,N_494);
and U879 (N_879,N_272,N_443);
nor U880 (N_880,N_297,N_433);
nand U881 (N_881,N_74,N_62);
xnor U882 (N_882,N_290,N_256);
nand U883 (N_883,N_477,N_47);
or U884 (N_884,N_469,N_136);
nor U885 (N_885,N_404,N_351);
or U886 (N_886,N_501,N_326);
or U887 (N_887,N_412,N_191);
nor U888 (N_888,N_215,N_356);
nand U889 (N_889,N_384,N_148);
or U890 (N_890,N_278,N_179);
nand U891 (N_891,N_424,N_145);
xor U892 (N_892,N_68,N_423);
nor U893 (N_893,N_512,N_190);
and U894 (N_894,N_176,N_135);
or U895 (N_895,N_205,N_241);
nand U896 (N_896,N_597,N_320);
nand U897 (N_897,N_339,N_273);
or U898 (N_898,N_108,N_432);
and U899 (N_899,N_259,N_348);
and U900 (N_900,N_270,N_431);
nand U901 (N_901,N_300,N_441);
and U902 (N_902,N_48,N_51);
nor U903 (N_903,N_403,N_15);
or U904 (N_904,N_170,N_536);
and U905 (N_905,N_84,N_417);
xor U906 (N_906,N_47,N_179);
and U907 (N_907,N_527,N_46);
nor U908 (N_908,N_269,N_61);
nor U909 (N_909,N_322,N_396);
nor U910 (N_910,N_67,N_503);
or U911 (N_911,N_445,N_232);
and U912 (N_912,N_149,N_77);
nor U913 (N_913,N_40,N_165);
xnor U914 (N_914,N_282,N_279);
nor U915 (N_915,N_555,N_51);
nor U916 (N_916,N_460,N_570);
or U917 (N_917,N_162,N_420);
nand U918 (N_918,N_511,N_49);
and U919 (N_919,N_492,N_222);
nor U920 (N_920,N_487,N_376);
and U921 (N_921,N_87,N_187);
and U922 (N_922,N_304,N_486);
nor U923 (N_923,N_131,N_512);
or U924 (N_924,N_444,N_572);
and U925 (N_925,N_294,N_63);
nand U926 (N_926,N_104,N_342);
and U927 (N_927,N_22,N_18);
nor U928 (N_928,N_175,N_288);
nor U929 (N_929,N_374,N_395);
nand U930 (N_930,N_541,N_23);
xor U931 (N_931,N_508,N_286);
and U932 (N_932,N_586,N_151);
or U933 (N_933,N_431,N_277);
nor U934 (N_934,N_538,N_311);
xor U935 (N_935,N_524,N_288);
and U936 (N_936,N_501,N_441);
nor U937 (N_937,N_199,N_83);
or U938 (N_938,N_46,N_274);
or U939 (N_939,N_372,N_51);
nand U940 (N_940,N_227,N_567);
and U941 (N_941,N_3,N_179);
and U942 (N_942,N_347,N_298);
nor U943 (N_943,N_429,N_326);
nor U944 (N_944,N_438,N_548);
nand U945 (N_945,N_110,N_180);
nand U946 (N_946,N_534,N_343);
and U947 (N_947,N_441,N_477);
nor U948 (N_948,N_500,N_401);
xnor U949 (N_949,N_45,N_423);
nor U950 (N_950,N_108,N_187);
or U951 (N_951,N_189,N_54);
or U952 (N_952,N_428,N_268);
nand U953 (N_953,N_252,N_312);
nand U954 (N_954,N_402,N_111);
xnor U955 (N_955,N_220,N_167);
and U956 (N_956,N_253,N_543);
nand U957 (N_957,N_114,N_334);
nand U958 (N_958,N_358,N_416);
nor U959 (N_959,N_142,N_583);
nor U960 (N_960,N_261,N_367);
nand U961 (N_961,N_409,N_56);
and U962 (N_962,N_357,N_492);
nand U963 (N_963,N_417,N_489);
nor U964 (N_964,N_54,N_355);
xor U965 (N_965,N_76,N_555);
nor U966 (N_966,N_507,N_281);
nand U967 (N_967,N_288,N_276);
or U968 (N_968,N_594,N_555);
nand U969 (N_969,N_363,N_90);
and U970 (N_970,N_265,N_317);
and U971 (N_971,N_434,N_281);
and U972 (N_972,N_297,N_469);
nor U973 (N_973,N_5,N_390);
nor U974 (N_974,N_132,N_299);
or U975 (N_975,N_465,N_90);
or U976 (N_976,N_310,N_471);
or U977 (N_977,N_290,N_254);
nand U978 (N_978,N_307,N_454);
nand U979 (N_979,N_377,N_96);
or U980 (N_980,N_447,N_86);
and U981 (N_981,N_168,N_208);
xnor U982 (N_982,N_487,N_61);
xor U983 (N_983,N_55,N_340);
nand U984 (N_984,N_437,N_71);
nand U985 (N_985,N_238,N_92);
and U986 (N_986,N_70,N_592);
nand U987 (N_987,N_107,N_427);
and U988 (N_988,N_553,N_284);
or U989 (N_989,N_307,N_123);
or U990 (N_990,N_540,N_585);
nor U991 (N_991,N_333,N_351);
nor U992 (N_992,N_161,N_336);
xor U993 (N_993,N_160,N_368);
or U994 (N_994,N_535,N_345);
nand U995 (N_995,N_515,N_400);
and U996 (N_996,N_562,N_341);
nand U997 (N_997,N_77,N_503);
nor U998 (N_998,N_450,N_477);
or U999 (N_999,N_548,N_33);
nand U1000 (N_1000,N_574,N_359);
or U1001 (N_1001,N_331,N_226);
nor U1002 (N_1002,N_309,N_370);
and U1003 (N_1003,N_225,N_494);
xor U1004 (N_1004,N_598,N_231);
or U1005 (N_1005,N_545,N_120);
nand U1006 (N_1006,N_383,N_26);
nor U1007 (N_1007,N_167,N_141);
nand U1008 (N_1008,N_121,N_257);
nor U1009 (N_1009,N_67,N_457);
nor U1010 (N_1010,N_257,N_89);
nand U1011 (N_1011,N_442,N_17);
nand U1012 (N_1012,N_466,N_554);
or U1013 (N_1013,N_126,N_382);
nor U1014 (N_1014,N_313,N_382);
or U1015 (N_1015,N_396,N_239);
nor U1016 (N_1016,N_184,N_26);
nand U1017 (N_1017,N_432,N_426);
nand U1018 (N_1018,N_127,N_485);
nor U1019 (N_1019,N_111,N_256);
nor U1020 (N_1020,N_135,N_16);
or U1021 (N_1021,N_393,N_106);
xnor U1022 (N_1022,N_458,N_490);
nor U1023 (N_1023,N_545,N_97);
xnor U1024 (N_1024,N_453,N_280);
or U1025 (N_1025,N_107,N_366);
or U1026 (N_1026,N_364,N_387);
xor U1027 (N_1027,N_195,N_588);
and U1028 (N_1028,N_374,N_467);
nand U1029 (N_1029,N_448,N_126);
nor U1030 (N_1030,N_392,N_363);
nor U1031 (N_1031,N_95,N_251);
nor U1032 (N_1032,N_452,N_491);
or U1033 (N_1033,N_575,N_315);
nand U1034 (N_1034,N_298,N_582);
nor U1035 (N_1035,N_110,N_91);
nor U1036 (N_1036,N_197,N_328);
nor U1037 (N_1037,N_273,N_62);
or U1038 (N_1038,N_472,N_60);
and U1039 (N_1039,N_391,N_326);
nor U1040 (N_1040,N_590,N_84);
nor U1041 (N_1041,N_242,N_588);
nand U1042 (N_1042,N_229,N_26);
or U1043 (N_1043,N_52,N_164);
and U1044 (N_1044,N_309,N_119);
nor U1045 (N_1045,N_195,N_238);
or U1046 (N_1046,N_428,N_246);
nor U1047 (N_1047,N_403,N_80);
nor U1048 (N_1048,N_512,N_218);
nor U1049 (N_1049,N_494,N_387);
nand U1050 (N_1050,N_259,N_576);
or U1051 (N_1051,N_426,N_324);
nor U1052 (N_1052,N_373,N_424);
or U1053 (N_1053,N_402,N_108);
and U1054 (N_1054,N_368,N_530);
or U1055 (N_1055,N_318,N_78);
and U1056 (N_1056,N_324,N_377);
nand U1057 (N_1057,N_170,N_443);
nor U1058 (N_1058,N_528,N_161);
xor U1059 (N_1059,N_309,N_576);
nand U1060 (N_1060,N_236,N_533);
nor U1061 (N_1061,N_557,N_35);
or U1062 (N_1062,N_210,N_233);
nor U1063 (N_1063,N_36,N_127);
and U1064 (N_1064,N_353,N_164);
xor U1065 (N_1065,N_583,N_196);
nor U1066 (N_1066,N_409,N_536);
and U1067 (N_1067,N_485,N_240);
xor U1068 (N_1068,N_531,N_228);
nor U1069 (N_1069,N_147,N_85);
and U1070 (N_1070,N_571,N_267);
nand U1071 (N_1071,N_597,N_308);
or U1072 (N_1072,N_79,N_308);
xnor U1073 (N_1073,N_209,N_81);
nor U1074 (N_1074,N_556,N_514);
or U1075 (N_1075,N_49,N_100);
nand U1076 (N_1076,N_6,N_251);
nand U1077 (N_1077,N_277,N_80);
xnor U1078 (N_1078,N_55,N_573);
nor U1079 (N_1079,N_14,N_450);
or U1080 (N_1080,N_296,N_43);
nand U1081 (N_1081,N_400,N_265);
and U1082 (N_1082,N_25,N_119);
nor U1083 (N_1083,N_362,N_27);
nor U1084 (N_1084,N_52,N_436);
or U1085 (N_1085,N_404,N_504);
and U1086 (N_1086,N_187,N_469);
xnor U1087 (N_1087,N_570,N_542);
nor U1088 (N_1088,N_142,N_505);
nand U1089 (N_1089,N_92,N_437);
nand U1090 (N_1090,N_306,N_534);
or U1091 (N_1091,N_583,N_541);
or U1092 (N_1092,N_246,N_94);
or U1093 (N_1093,N_174,N_269);
nor U1094 (N_1094,N_378,N_428);
and U1095 (N_1095,N_126,N_416);
xnor U1096 (N_1096,N_351,N_573);
nand U1097 (N_1097,N_307,N_512);
nand U1098 (N_1098,N_312,N_14);
or U1099 (N_1099,N_493,N_197);
or U1100 (N_1100,N_216,N_524);
nand U1101 (N_1101,N_312,N_377);
nand U1102 (N_1102,N_558,N_132);
nor U1103 (N_1103,N_553,N_425);
and U1104 (N_1104,N_489,N_415);
nor U1105 (N_1105,N_20,N_323);
xor U1106 (N_1106,N_335,N_38);
and U1107 (N_1107,N_4,N_149);
and U1108 (N_1108,N_404,N_574);
and U1109 (N_1109,N_97,N_420);
nor U1110 (N_1110,N_75,N_181);
and U1111 (N_1111,N_151,N_217);
nand U1112 (N_1112,N_183,N_300);
and U1113 (N_1113,N_374,N_236);
and U1114 (N_1114,N_287,N_1);
nor U1115 (N_1115,N_414,N_93);
and U1116 (N_1116,N_498,N_563);
nand U1117 (N_1117,N_278,N_508);
or U1118 (N_1118,N_35,N_156);
or U1119 (N_1119,N_570,N_3);
nor U1120 (N_1120,N_363,N_218);
or U1121 (N_1121,N_137,N_252);
and U1122 (N_1122,N_520,N_561);
and U1123 (N_1123,N_510,N_33);
or U1124 (N_1124,N_10,N_104);
nor U1125 (N_1125,N_376,N_97);
and U1126 (N_1126,N_96,N_25);
nand U1127 (N_1127,N_275,N_448);
and U1128 (N_1128,N_405,N_418);
or U1129 (N_1129,N_278,N_384);
and U1130 (N_1130,N_83,N_127);
and U1131 (N_1131,N_561,N_240);
nor U1132 (N_1132,N_50,N_184);
nor U1133 (N_1133,N_396,N_383);
or U1134 (N_1134,N_1,N_254);
or U1135 (N_1135,N_346,N_18);
and U1136 (N_1136,N_435,N_563);
or U1137 (N_1137,N_487,N_455);
or U1138 (N_1138,N_560,N_543);
xnor U1139 (N_1139,N_378,N_433);
nand U1140 (N_1140,N_386,N_476);
nand U1141 (N_1141,N_432,N_449);
and U1142 (N_1142,N_447,N_243);
nand U1143 (N_1143,N_198,N_535);
or U1144 (N_1144,N_261,N_293);
xor U1145 (N_1145,N_560,N_305);
nand U1146 (N_1146,N_333,N_156);
or U1147 (N_1147,N_491,N_477);
or U1148 (N_1148,N_272,N_279);
nand U1149 (N_1149,N_216,N_130);
nand U1150 (N_1150,N_455,N_167);
nand U1151 (N_1151,N_464,N_237);
nor U1152 (N_1152,N_298,N_120);
and U1153 (N_1153,N_592,N_28);
xnor U1154 (N_1154,N_506,N_427);
or U1155 (N_1155,N_478,N_542);
nor U1156 (N_1156,N_89,N_369);
and U1157 (N_1157,N_347,N_510);
nor U1158 (N_1158,N_56,N_192);
and U1159 (N_1159,N_356,N_412);
and U1160 (N_1160,N_393,N_501);
nor U1161 (N_1161,N_575,N_553);
nand U1162 (N_1162,N_492,N_302);
nor U1163 (N_1163,N_220,N_500);
nor U1164 (N_1164,N_116,N_387);
nand U1165 (N_1165,N_88,N_523);
nor U1166 (N_1166,N_542,N_329);
nand U1167 (N_1167,N_415,N_37);
xnor U1168 (N_1168,N_99,N_51);
nand U1169 (N_1169,N_420,N_197);
or U1170 (N_1170,N_460,N_245);
nor U1171 (N_1171,N_480,N_341);
or U1172 (N_1172,N_188,N_417);
or U1173 (N_1173,N_87,N_445);
and U1174 (N_1174,N_304,N_382);
nand U1175 (N_1175,N_168,N_285);
or U1176 (N_1176,N_240,N_234);
nor U1177 (N_1177,N_350,N_382);
nor U1178 (N_1178,N_468,N_147);
or U1179 (N_1179,N_55,N_30);
nor U1180 (N_1180,N_61,N_221);
nand U1181 (N_1181,N_11,N_268);
xnor U1182 (N_1182,N_232,N_487);
or U1183 (N_1183,N_162,N_513);
nor U1184 (N_1184,N_502,N_296);
nor U1185 (N_1185,N_404,N_433);
xnor U1186 (N_1186,N_506,N_174);
and U1187 (N_1187,N_51,N_84);
or U1188 (N_1188,N_230,N_545);
and U1189 (N_1189,N_371,N_123);
and U1190 (N_1190,N_219,N_478);
xnor U1191 (N_1191,N_351,N_174);
nor U1192 (N_1192,N_313,N_232);
nor U1193 (N_1193,N_278,N_245);
nand U1194 (N_1194,N_260,N_412);
or U1195 (N_1195,N_154,N_141);
and U1196 (N_1196,N_322,N_346);
nor U1197 (N_1197,N_93,N_367);
or U1198 (N_1198,N_147,N_499);
nand U1199 (N_1199,N_301,N_426);
or U1200 (N_1200,N_803,N_696);
and U1201 (N_1201,N_765,N_871);
or U1202 (N_1202,N_918,N_978);
or U1203 (N_1203,N_866,N_1189);
nand U1204 (N_1204,N_669,N_772);
or U1205 (N_1205,N_1029,N_694);
nor U1206 (N_1206,N_603,N_848);
or U1207 (N_1207,N_835,N_974);
nand U1208 (N_1208,N_882,N_644);
or U1209 (N_1209,N_760,N_1197);
and U1210 (N_1210,N_650,N_1105);
and U1211 (N_1211,N_635,N_612);
or U1212 (N_1212,N_770,N_1153);
nor U1213 (N_1213,N_954,N_683);
or U1214 (N_1214,N_963,N_1099);
and U1215 (N_1215,N_1007,N_867);
or U1216 (N_1216,N_1194,N_890);
and U1217 (N_1217,N_641,N_657);
nor U1218 (N_1218,N_606,N_673);
nor U1219 (N_1219,N_927,N_802);
and U1220 (N_1220,N_864,N_762);
or U1221 (N_1221,N_1097,N_884);
or U1222 (N_1222,N_821,N_638);
and U1223 (N_1223,N_862,N_759);
or U1224 (N_1224,N_861,N_713);
nor U1225 (N_1225,N_892,N_659);
or U1226 (N_1226,N_677,N_928);
and U1227 (N_1227,N_1134,N_744);
and U1228 (N_1228,N_850,N_739);
xor U1229 (N_1229,N_1191,N_908);
nand U1230 (N_1230,N_779,N_932);
xor U1231 (N_1231,N_629,N_647);
and U1232 (N_1232,N_1090,N_665);
and U1233 (N_1233,N_1091,N_632);
nor U1234 (N_1234,N_895,N_930);
nand U1235 (N_1235,N_922,N_1149);
nor U1236 (N_1236,N_1107,N_883);
nor U1237 (N_1237,N_1047,N_952);
and U1238 (N_1238,N_986,N_875);
or U1239 (N_1239,N_1161,N_799);
nand U1240 (N_1240,N_728,N_977);
or U1241 (N_1241,N_1108,N_661);
and U1242 (N_1242,N_1019,N_705);
or U1243 (N_1243,N_839,N_783);
nand U1244 (N_1244,N_847,N_1138);
and U1245 (N_1245,N_637,N_923);
and U1246 (N_1246,N_944,N_732);
nor U1247 (N_1247,N_849,N_703);
nand U1248 (N_1248,N_995,N_1068);
or U1249 (N_1249,N_1013,N_1085);
nand U1250 (N_1250,N_698,N_1142);
and U1251 (N_1251,N_721,N_961);
nand U1252 (N_1252,N_1115,N_1146);
xor U1253 (N_1253,N_725,N_1185);
nor U1254 (N_1254,N_999,N_1167);
and U1255 (N_1255,N_1101,N_768);
nand U1256 (N_1256,N_766,N_1177);
nand U1257 (N_1257,N_1032,N_1192);
xor U1258 (N_1258,N_860,N_1152);
nand U1259 (N_1259,N_623,N_748);
nor U1260 (N_1260,N_1089,N_877);
xor U1261 (N_1261,N_1122,N_1008);
nand U1262 (N_1262,N_962,N_1096);
nand U1263 (N_1263,N_610,N_617);
nand U1264 (N_1264,N_758,N_820);
and U1265 (N_1265,N_642,N_989);
and U1266 (N_1266,N_1158,N_790);
xnor U1267 (N_1267,N_807,N_789);
xnor U1268 (N_1268,N_894,N_852);
and U1269 (N_1269,N_1184,N_602);
or U1270 (N_1270,N_897,N_828);
or U1271 (N_1271,N_1103,N_806);
nor U1272 (N_1272,N_1009,N_1088);
nand U1273 (N_1273,N_858,N_798);
or U1274 (N_1274,N_787,N_733);
nand U1275 (N_1275,N_992,N_745);
nand U1276 (N_1276,N_656,N_1056);
or U1277 (N_1277,N_1140,N_1175);
or U1278 (N_1278,N_1049,N_1126);
nor U1279 (N_1279,N_797,N_788);
nand U1280 (N_1280,N_822,N_662);
or U1281 (N_1281,N_845,N_697);
and U1282 (N_1282,N_856,N_826);
nand U1283 (N_1283,N_940,N_920);
or U1284 (N_1284,N_785,N_953);
nand U1285 (N_1285,N_921,N_1015);
or U1286 (N_1286,N_619,N_1163);
nor U1287 (N_1287,N_924,N_775);
and U1288 (N_1288,N_959,N_1120);
nand U1289 (N_1289,N_899,N_915);
or U1290 (N_1290,N_838,N_675);
and U1291 (N_1291,N_936,N_605);
or U1292 (N_1292,N_1081,N_1058);
xnor U1293 (N_1293,N_947,N_1180);
and U1294 (N_1294,N_960,N_722);
or U1295 (N_1295,N_670,N_625);
nor U1296 (N_1296,N_782,N_1154);
nor U1297 (N_1297,N_1166,N_925);
nor U1298 (N_1298,N_907,N_1135);
nor U1299 (N_1299,N_633,N_950);
or U1300 (N_1300,N_709,N_701);
and U1301 (N_1301,N_1075,N_649);
nand U1302 (N_1302,N_1044,N_851);
nand U1303 (N_1303,N_715,N_1035);
nor U1304 (N_1304,N_1109,N_906);
or U1305 (N_1305,N_780,N_613);
nor U1306 (N_1306,N_1181,N_793);
nand U1307 (N_1307,N_640,N_695);
and U1308 (N_1308,N_1036,N_916);
and U1309 (N_1309,N_655,N_704);
and U1310 (N_1310,N_621,N_898);
or U1311 (N_1311,N_742,N_691);
and U1312 (N_1312,N_809,N_935);
xor U1313 (N_1313,N_651,N_912);
nand U1314 (N_1314,N_1136,N_919);
nor U1315 (N_1315,N_729,N_943);
nand U1316 (N_1316,N_1017,N_1102);
nand U1317 (N_1317,N_972,N_749);
and U1318 (N_1318,N_873,N_1073);
nand U1319 (N_1319,N_1114,N_700);
nor U1320 (N_1320,N_1055,N_991);
nand U1321 (N_1321,N_681,N_841);
nand U1322 (N_1322,N_1119,N_1030);
or U1323 (N_1323,N_1160,N_1024);
or U1324 (N_1324,N_904,N_1168);
nand U1325 (N_1325,N_1034,N_805);
nand U1326 (N_1326,N_979,N_840);
xnor U1327 (N_1327,N_639,N_668);
nor U1328 (N_1328,N_689,N_1172);
or U1329 (N_1329,N_938,N_753);
and U1330 (N_1330,N_1054,N_718);
nor U1331 (N_1331,N_1023,N_1143);
nand U1332 (N_1332,N_827,N_769);
and U1333 (N_1333,N_636,N_844);
nand U1334 (N_1334,N_1069,N_1179);
xor U1335 (N_1335,N_1072,N_857);
nand U1336 (N_1336,N_843,N_816);
xnor U1337 (N_1337,N_1018,N_1004);
or U1338 (N_1338,N_981,N_717);
nor U1339 (N_1339,N_755,N_1020);
or U1340 (N_1340,N_975,N_740);
or U1341 (N_1341,N_654,N_716);
xnor U1342 (N_1342,N_955,N_653);
or U1343 (N_1343,N_600,N_863);
or U1344 (N_1344,N_1026,N_1157);
and U1345 (N_1345,N_970,N_939);
nor U1346 (N_1346,N_660,N_988);
nor U1347 (N_1347,N_869,N_674);
nand U1348 (N_1348,N_887,N_664);
nor U1349 (N_1349,N_968,N_814);
or U1350 (N_1350,N_846,N_946);
or U1351 (N_1351,N_627,N_804);
or U1352 (N_1352,N_648,N_687);
nand U1353 (N_1353,N_751,N_1150);
and U1354 (N_1354,N_1042,N_1043);
and U1355 (N_1355,N_1074,N_1076);
and U1356 (N_1356,N_795,N_1104);
nor U1357 (N_1357,N_824,N_1063);
and U1358 (N_1358,N_726,N_889);
and U1359 (N_1359,N_646,N_692);
and U1360 (N_1360,N_735,N_1174);
or U1361 (N_1361,N_1038,N_604);
or U1362 (N_1362,N_1005,N_1012);
or U1363 (N_1363,N_791,N_690);
nor U1364 (N_1364,N_830,N_1128);
and U1365 (N_1365,N_792,N_615);
xor U1366 (N_1366,N_818,N_1070);
nand U1367 (N_1367,N_1125,N_1195);
xnor U1368 (N_1368,N_1051,N_982);
nand U1369 (N_1369,N_917,N_933);
and U1370 (N_1370,N_730,N_984);
or U1371 (N_1371,N_881,N_750);
and U1372 (N_1372,N_736,N_987);
nand U1373 (N_1373,N_1010,N_1027);
nand U1374 (N_1374,N_994,N_872);
or U1375 (N_1375,N_1118,N_1022);
nand U1376 (N_1376,N_1129,N_680);
and U1377 (N_1377,N_1000,N_1165);
nand U1378 (N_1378,N_693,N_737);
or U1379 (N_1379,N_741,N_1188);
nand U1380 (N_1380,N_1060,N_608);
xor U1381 (N_1381,N_1186,N_1100);
or U1382 (N_1382,N_719,N_1199);
or U1383 (N_1383,N_1137,N_1077);
nand U1384 (N_1384,N_1046,N_879);
nor U1385 (N_1385,N_786,N_1130);
or U1386 (N_1386,N_1132,N_859);
nor U1387 (N_1387,N_909,N_980);
nand U1388 (N_1388,N_1078,N_951);
nand U1389 (N_1389,N_1173,N_958);
nand U1390 (N_1390,N_1011,N_1169);
nor U1391 (N_1391,N_1062,N_634);
nor U1392 (N_1392,N_1061,N_626);
or U1393 (N_1393,N_1052,N_672);
nor U1394 (N_1394,N_712,N_624);
or U1395 (N_1395,N_874,N_1139);
nor U1396 (N_1396,N_1082,N_1123);
nand U1397 (N_1397,N_1147,N_817);
and U1398 (N_1398,N_893,N_973);
nor U1399 (N_1399,N_834,N_937);
nand U1400 (N_1400,N_880,N_965);
or U1401 (N_1401,N_800,N_902);
nor U1402 (N_1402,N_1021,N_1196);
nand U1403 (N_1403,N_1039,N_724);
or U1404 (N_1404,N_1040,N_773);
and U1405 (N_1405,N_996,N_1193);
nand U1406 (N_1406,N_891,N_688);
nand U1407 (N_1407,N_1066,N_784);
and U1408 (N_1408,N_756,N_1031);
and U1409 (N_1409,N_1124,N_810);
nand U1410 (N_1410,N_900,N_855);
or U1411 (N_1411,N_1144,N_607);
nand U1412 (N_1412,N_752,N_990);
and U1413 (N_1413,N_993,N_1176);
and U1414 (N_1414,N_1190,N_777);
nand U1415 (N_1415,N_914,N_774);
xor U1416 (N_1416,N_618,N_1113);
xnor U1417 (N_1417,N_983,N_1162);
nor U1418 (N_1418,N_949,N_868);
nand U1419 (N_1419,N_738,N_1071);
nor U1420 (N_1420,N_676,N_1145);
xor U1421 (N_1421,N_1116,N_1014);
or U1422 (N_1422,N_763,N_708);
nor U1423 (N_1423,N_1164,N_747);
nor U1424 (N_1424,N_616,N_1131);
nor U1425 (N_1425,N_1065,N_658);
nand U1426 (N_1426,N_1053,N_1084);
xor U1427 (N_1427,N_948,N_1045);
or U1428 (N_1428,N_966,N_667);
and U1429 (N_1429,N_1106,N_630);
and U1430 (N_1430,N_903,N_885);
nand U1431 (N_1431,N_1178,N_1133);
or U1432 (N_1432,N_710,N_812);
xnor U1433 (N_1433,N_825,N_876);
nor U1434 (N_1434,N_1003,N_778);
nand U1435 (N_1435,N_1087,N_967);
and U1436 (N_1436,N_1092,N_643);
xnor U1437 (N_1437,N_842,N_706);
nand U1438 (N_1438,N_1083,N_985);
nor U1439 (N_1439,N_1057,N_813);
xnor U1440 (N_1440,N_685,N_666);
and U1441 (N_1441,N_1080,N_1098);
nand U1442 (N_1442,N_1086,N_1064);
and U1443 (N_1443,N_714,N_905);
nor U1444 (N_1444,N_611,N_878);
and U1445 (N_1445,N_865,N_1059);
or U1446 (N_1446,N_957,N_886);
and U1447 (N_1447,N_836,N_1006);
nand U1448 (N_1448,N_645,N_671);
and U1449 (N_1449,N_601,N_767);
xor U1450 (N_1450,N_942,N_1002);
nor U1451 (N_1451,N_734,N_911);
and U1452 (N_1452,N_853,N_901);
nor U1453 (N_1453,N_757,N_997);
nand U1454 (N_1454,N_746,N_1028);
nor U1455 (N_1455,N_831,N_754);
nand U1456 (N_1456,N_1187,N_854);
or U1457 (N_1457,N_829,N_1155);
and U1458 (N_1458,N_945,N_609);
nand U1459 (N_1459,N_620,N_819);
and U1460 (N_1460,N_1183,N_870);
nand U1461 (N_1461,N_663,N_964);
nor U1462 (N_1462,N_1121,N_815);
or U1463 (N_1463,N_1148,N_956);
nand U1464 (N_1464,N_837,N_743);
and U1465 (N_1465,N_678,N_808);
and U1466 (N_1466,N_1110,N_1111);
nand U1467 (N_1467,N_1117,N_781);
or U1468 (N_1468,N_1171,N_1050);
nand U1469 (N_1469,N_699,N_1037);
or U1470 (N_1470,N_1001,N_1079);
nor U1471 (N_1471,N_811,N_888);
nor U1472 (N_1472,N_833,N_652);
and U1473 (N_1473,N_764,N_1198);
or U1474 (N_1474,N_702,N_969);
or U1475 (N_1475,N_801,N_941);
nor U1476 (N_1476,N_1041,N_686);
nor U1477 (N_1477,N_679,N_684);
nor U1478 (N_1478,N_1127,N_1094);
and U1479 (N_1479,N_934,N_1033);
nor U1480 (N_1480,N_910,N_707);
nor U1481 (N_1481,N_976,N_628);
and U1482 (N_1482,N_711,N_929);
and U1483 (N_1483,N_926,N_1016);
xnor U1484 (N_1484,N_631,N_1112);
nand U1485 (N_1485,N_1025,N_1151);
nor U1486 (N_1486,N_832,N_1170);
nand U1487 (N_1487,N_1093,N_796);
or U1488 (N_1488,N_1156,N_776);
or U1489 (N_1489,N_913,N_720);
nand U1490 (N_1490,N_896,N_614);
and U1491 (N_1491,N_1159,N_931);
nand U1492 (N_1492,N_1095,N_1048);
or U1493 (N_1493,N_998,N_682);
nand U1494 (N_1494,N_761,N_823);
and U1495 (N_1495,N_1067,N_622);
xnor U1496 (N_1496,N_971,N_723);
nor U1497 (N_1497,N_794,N_1141);
nor U1498 (N_1498,N_727,N_1182);
nor U1499 (N_1499,N_771,N_731);
or U1500 (N_1500,N_618,N_675);
or U1501 (N_1501,N_1000,N_607);
nand U1502 (N_1502,N_1089,N_956);
or U1503 (N_1503,N_1095,N_618);
and U1504 (N_1504,N_1026,N_957);
xor U1505 (N_1505,N_710,N_1046);
or U1506 (N_1506,N_940,N_833);
nand U1507 (N_1507,N_630,N_742);
nand U1508 (N_1508,N_917,N_705);
and U1509 (N_1509,N_1133,N_619);
and U1510 (N_1510,N_1054,N_927);
and U1511 (N_1511,N_1184,N_1028);
and U1512 (N_1512,N_903,N_928);
nor U1513 (N_1513,N_856,N_816);
and U1514 (N_1514,N_1186,N_971);
nor U1515 (N_1515,N_616,N_759);
xor U1516 (N_1516,N_1198,N_1155);
xnor U1517 (N_1517,N_986,N_711);
nand U1518 (N_1518,N_978,N_837);
nor U1519 (N_1519,N_1147,N_1144);
nand U1520 (N_1520,N_1114,N_1015);
or U1521 (N_1521,N_1161,N_1011);
and U1522 (N_1522,N_636,N_1003);
nand U1523 (N_1523,N_925,N_1054);
xor U1524 (N_1524,N_797,N_1061);
or U1525 (N_1525,N_1191,N_617);
nand U1526 (N_1526,N_1194,N_889);
nor U1527 (N_1527,N_668,N_848);
xnor U1528 (N_1528,N_877,N_773);
nor U1529 (N_1529,N_889,N_969);
and U1530 (N_1530,N_614,N_783);
nor U1531 (N_1531,N_699,N_860);
or U1532 (N_1532,N_811,N_1090);
nand U1533 (N_1533,N_1174,N_667);
and U1534 (N_1534,N_1034,N_1118);
or U1535 (N_1535,N_953,N_772);
xnor U1536 (N_1536,N_793,N_1011);
or U1537 (N_1537,N_1173,N_675);
nand U1538 (N_1538,N_761,N_1178);
nand U1539 (N_1539,N_814,N_1165);
nor U1540 (N_1540,N_716,N_1011);
nand U1541 (N_1541,N_645,N_767);
nand U1542 (N_1542,N_850,N_758);
and U1543 (N_1543,N_875,N_866);
nor U1544 (N_1544,N_1024,N_678);
nand U1545 (N_1545,N_626,N_867);
or U1546 (N_1546,N_1130,N_878);
nand U1547 (N_1547,N_617,N_969);
or U1548 (N_1548,N_787,N_629);
nand U1549 (N_1549,N_1153,N_1011);
or U1550 (N_1550,N_1088,N_966);
nor U1551 (N_1551,N_718,N_720);
nand U1552 (N_1552,N_657,N_796);
nor U1553 (N_1553,N_1040,N_1042);
or U1554 (N_1554,N_816,N_985);
xor U1555 (N_1555,N_913,N_660);
or U1556 (N_1556,N_659,N_1014);
xor U1557 (N_1557,N_1143,N_885);
xor U1558 (N_1558,N_804,N_1062);
nor U1559 (N_1559,N_761,N_659);
nor U1560 (N_1560,N_902,N_1073);
nor U1561 (N_1561,N_802,N_809);
or U1562 (N_1562,N_1161,N_834);
xor U1563 (N_1563,N_872,N_881);
or U1564 (N_1564,N_1095,N_641);
or U1565 (N_1565,N_945,N_1032);
and U1566 (N_1566,N_942,N_776);
nor U1567 (N_1567,N_618,N_614);
and U1568 (N_1568,N_811,N_951);
or U1569 (N_1569,N_1081,N_1078);
and U1570 (N_1570,N_750,N_827);
nand U1571 (N_1571,N_632,N_825);
nor U1572 (N_1572,N_804,N_790);
and U1573 (N_1573,N_943,N_1013);
nand U1574 (N_1574,N_634,N_622);
or U1575 (N_1575,N_862,N_626);
nand U1576 (N_1576,N_722,N_614);
nand U1577 (N_1577,N_799,N_882);
nor U1578 (N_1578,N_851,N_660);
and U1579 (N_1579,N_650,N_816);
and U1580 (N_1580,N_851,N_1112);
nor U1581 (N_1581,N_968,N_707);
nor U1582 (N_1582,N_1094,N_736);
nand U1583 (N_1583,N_608,N_1198);
xnor U1584 (N_1584,N_627,N_638);
nor U1585 (N_1585,N_1023,N_1076);
and U1586 (N_1586,N_1007,N_710);
and U1587 (N_1587,N_1027,N_651);
nand U1588 (N_1588,N_1105,N_859);
or U1589 (N_1589,N_769,N_958);
or U1590 (N_1590,N_740,N_965);
and U1591 (N_1591,N_831,N_922);
and U1592 (N_1592,N_611,N_960);
nor U1593 (N_1593,N_706,N_1153);
or U1594 (N_1594,N_722,N_1059);
nor U1595 (N_1595,N_1129,N_883);
nor U1596 (N_1596,N_1148,N_642);
nor U1597 (N_1597,N_1006,N_952);
or U1598 (N_1598,N_949,N_1009);
nand U1599 (N_1599,N_666,N_868);
or U1600 (N_1600,N_1092,N_704);
nand U1601 (N_1601,N_1149,N_866);
nand U1602 (N_1602,N_731,N_669);
or U1603 (N_1603,N_1037,N_1099);
nor U1604 (N_1604,N_856,N_785);
and U1605 (N_1605,N_1095,N_1195);
nand U1606 (N_1606,N_1117,N_1031);
or U1607 (N_1607,N_768,N_785);
nand U1608 (N_1608,N_1086,N_974);
xnor U1609 (N_1609,N_802,N_1080);
or U1610 (N_1610,N_943,N_1043);
or U1611 (N_1611,N_755,N_676);
xnor U1612 (N_1612,N_749,N_781);
nand U1613 (N_1613,N_641,N_638);
xor U1614 (N_1614,N_630,N_862);
or U1615 (N_1615,N_813,N_1098);
nor U1616 (N_1616,N_929,N_1062);
xnor U1617 (N_1617,N_918,N_664);
or U1618 (N_1618,N_1169,N_1135);
nor U1619 (N_1619,N_654,N_673);
xor U1620 (N_1620,N_742,N_938);
xor U1621 (N_1621,N_677,N_1171);
nand U1622 (N_1622,N_1145,N_703);
and U1623 (N_1623,N_743,N_1091);
and U1624 (N_1624,N_932,N_840);
and U1625 (N_1625,N_686,N_1102);
nand U1626 (N_1626,N_1030,N_619);
xor U1627 (N_1627,N_1004,N_632);
and U1628 (N_1628,N_1020,N_893);
xor U1629 (N_1629,N_723,N_671);
nand U1630 (N_1630,N_1006,N_1066);
nor U1631 (N_1631,N_1199,N_912);
or U1632 (N_1632,N_1020,N_1087);
xor U1633 (N_1633,N_780,N_928);
nor U1634 (N_1634,N_1162,N_604);
or U1635 (N_1635,N_785,N_825);
nor U1636 (N_1636,N_826,N_1192);
and U1637 (N_1637,N_1020,N_1184);
xnor U1638 (N_1638,N_707,N_999);
nor U1639 (N_1639,N_1042,N_1100);
and U1640 (N_1640,N_729,N_719);
xnor U1641 (N_1641,N_728,N_853);
or U1642 (N_1642,N_1158,N_788);
nand U1643 (N_1643,N_733,N_901);
nand U1644 (N_1644,N_809,N_1141);
or U1645 (N_1645,N_904,N_667);
and U1646 (N_1646,N_1125,N_686);
nand U1647 (N_1647,N_922,N_881);
nor U1648 (N_1648,N_738,N_1112);
nand U1649 (N_1649,N_1135,N_732);
nor U1650 (N_1650,N_971,N_645);
nand U1651 (N_1651,N_930,N_1025);
and U1652 (N_1652,N_848,N_928);
nand U1653 (N_1653,N_1110,N_808);
or U1654 (N_1654,N_967,N_878);
or U1655 (N_1655,N_968,N_650);
nand U1656 (N_1656,N_1050,N_1124);
nand U1657 (N_1657,N_687,N_837);
and U1658 (N_1658,N_806,N_1173);
or U1659 (N_1659,N_938,N_615);
and U1660 (N_1660,N_955,N_603);
nand U1661 (N_1661,N_1174,N_732);
nand U1662 (N_1662,N_904,N_777);
or U1663 (N_1663,N_871,N_1172);
nor U1664 (N_1664,N_648,N_1084);
or U1665 (N_1665,N_762,N_994);
nor U1666 (N_1666,N_649,N_1150);
and U1667 (N_1667,N_1184,N_933);
nor U1668 (N_1668,N_696,N_634);
nand U1669 (N_1669,N_1190,N_678);
or U1670 (N_1670,N_706,N_1071);
nand U1671 (N_1671,N_1097,N_822);
and U1672 (N_1672,N_877,N_905);
nand U1673 (N_1673,N_1030,N_648);
xnor U1674 (N_1674,N_744,N_757);
or U1675 (N_1675,N_799,N_1058);
or U1676 (N_1676,N_1061,N_1103);
and U1677 (N_1677,N_1138,N_825);
nor U1678 (N_1678,N_1044,N_889);
and U1679 (N_1679,N_1040,N_1179);
nor U1680 (N_1680,N_649,N_908);
nor U1681 (N_1681,N_885,N_937);
or U1682 (N_1682,N_1150,N_909);
nand U1683 (N_1683,N_1122,N_981);
nand U1684 (N_1684,N_939,N_895);
nor U1685 (N_1685,N_929,N_666);
nand U1686 (N_1686,N_1184,N_1061);
xnor U1687 (N_1687,N_1169,N_785);
nor U1688 (N_1688,N_818,N_817);
nand U1689 (N_1689,N_923,N_1040);
nand U1690 (N_1690,N_641,N_659);
nor U1691 (N_1691,N_997,N_953);
nand U1692 (N_1692,N_1182,N_802);
nand U1693 (N_1693,N_982,N_1027);
or U1694 (N_1694,N_882,N_1073);
nand U1695 (N_1695,N_918,N_1194);
or U1696 (N_1696,N_646,N_687);
or U1697 (N_1697,N_942,N_748);
nand U1698 (N_1698,N_840,N_1195);
nand U1699 (N_1699,N_711,N_632);
nor U1700 (N_1700,N_669,N_919);
or U1701 (N_1701,N_1049,N_1153);
nor U1702 (N_1702,N_1102,N_964);
nor U1703 (N_1703,N_1042,N_1120);
xor U1704 (N_1704,N_1104,N_1140);
and U1705 (N_1705,N_720,N_706);
nand U1706 (N_1706,N_702,N_938);
and U1707 (N_1707,N_1156,N_619);
nand U1708 (N_1708,N_960,N_962);
or U1709 (N_1709,N_1124,N_904);
nand U1710 (N_1710,N_875,N_1175);
nand U1711 (N_1711,N_1180,N_1095);
nand U1712 (N_1712,N_832,N_818);
nand U1713 (N_1713,N_1087,N_991);
and U1714 (N_1714,N_1027,N_967);
and U1715 (N_1715,N_631,N_782);
nor U1716 (N_1716,N_1112,N_694);
nand U1717 (N_1717,N_1163,N_1199);
or U1718 (N_1718,N_977,N_1000);
xor U1719 (N_1719,N_813,N_922);
and U1720 (N_1720,N_1137,N_815);
xnor U1721 (N_1721,N_1086,N_659);
and U1722 (N_1722,N_1072,N_1000);
and U1723 (N_1723,N_1074,N_692);
nor U1724 (N_1724,N_648,N_869);
nand U1725 (N_1725,N_1013,N_634);
nor U1726 (N_1726,N_1102,N_957);
and U1727 (N_1727,N_702,N_831);
nand U1728 (N_1728,N_1197,N_1055);
nor U1729 (N_1729,N_1009,N_998);
nand U1730 (N_1730,N_621,N_673);
nand U1731 (N_1731,N_927,N_1131);
or U1732 (N_1732,N_1029,N_767);
nor U1733 (N_1733,N_874,N_939);
nand U1734 (N_1734,N_1033,N_605);
and U1735 (N_1735,N_1014,N_670);
and U1736 (N_1736,N_881,N_1155);
nand U1737 (N_1737,N_687,N_1137);
and U1738 (N_1738,N_815,N_836);
nor U1739 (N_1739,N_819,N_1044);
or U1740 (N_1740,N_738,N_769);
nor U1741 (N_1741,N_891,N_1066);
nor U1742 (N_1742,N_892,N_933);
and U1743 (N_1743,N_871,N_1091);
nand U1744 (N_1744,N_940,N_937);
or U1745 (N_1745,N_703,N_1052);
and U1746 (N_1746,N_987,N_877);
or U1747 (N_1747,N_903,N_1013);
nor U1748 (N_1748,N_946,N_941);
and U1749 (N_1749,N_897,N_1078);
or U1750 (N_1750,N_1158,N_1160);
and U1751 (N_1751,N_1004,N_836);
nor U1752 (N_1752,N_1151,N_895);
nand U1753 (N_1753,N_936,N_1035);
nand U1754 (N_1754,N_1148,N_904);
or U1755 (N_1755,N_983,N_693);
and U1756 (N_1756,N_868,N_1089);
nor U1757 (N_1757,N_660,N_828);
nor U1758 (N_1758,N_657,N_906);
nor U1759 (N_1759,N_945,N_688);
nor U1760 (N_1760,N_1018,N_1172);
and U1761 (N_1761,N_824,N_1077);
xnor U1762 (N_1762,N_1085,N_802);
nor U1763 (N_1763,N_1026,N_661);
nand U1764 (N_1764,N_641,N_667);
nand U1765 (N_1765,N_980,N_911);
or U1766 (N_1766,N_966,N_733);
and U1767 (N_1767,N_1054,N_1090);
nand U1768 (N_1768,N_749,N_682);
or U1769 (N_1769,N_901,N_987);
nand U1770 (N_1770,N_800,N_1051);
xor U1771 (N_1771,N_678,N_610);
and U1772 (N_1772,N_1192,N_630);
nand U1773 (N_1773,N_760,N_793);
or U1774 (N_1774,N_912,N_829);
xor U1775 (N_1775,N_664,N_967);
and U1776 (N_1776,N_1122,N_989);
nand U1777 (N_1777,N_833,N_703);
or U1778 (N_1778,N_757,N_769);
and U1779 (N_1779,N_1155,N_830);
and U1780 (N_1780,N_899,N_1158);
nand U1781 (N_1781,N_1047,N_826);
nand U1782 (N_1782,N_1016,N_1107);
and U1783 (N_1783,N_1088,N_1039);
nand U1784 (N_1784,N_1012,N_737);
nor U1785 (N_1785,N_1162,N_682);
or U1786 (N_1786,N_872,N_815);
and U1787 (N_1787,N_779,N_948);
nor U1788 (N_1788,N_1008,N_865);
xnor U1789 (N_1789,N_616,N_777);
and U1790 (N_1790,N_762,N_917);
nor U1791 (N_1791,N_1067,N_827);
nand U1792 (N_1792,N_632,N_963);
xor U1793 (N_1793,N_1002,N_943);
nand U1794 (N_1794,N_732,N_1170);
or U1795 (N_1795,N_897,N_762);
or U1796 (N_1796,N_777,N_955);
and U1797 (N_1797,N_1084,N_1130);
nor U1798 (N_1798,N_724,N_1191);
xor U1799 (N_1799,N_1149,N_1138);
or U1800 (N_1800,N_1426,N_1799);
or U1801 (N_1801,N_1330,N_1327);
nor U1802 (N_1802,N_1266,N_1739);
nor U1803 (N_1803,N_1428,N_1316);
xor U1804 (N_1804,N_1408,N_1645);
nor U1805 (N_1805,N_1405,N_1675);
nor U1806 (N_1806,N_1781,N_1219);
or U1807 (N_1807,N_1478,N_1716);
and U1808 (N_1808,N_1289,N_1696);
and U1809 (N_1809,N_1424,N_1782);
or U1810 (N_1810,N_1208,N_1298);
xor U1811 (N_1811,N_1394,N_1772);
nand U1812 (N_1812,N_1701,N_1381);
or U1813 (N_1813,N_1679,N_1248);
and U1814 (N_1814,N_1361,N_1324);
or U1815 (N_1815,N_1542,N_1616);
xnor U1816 (N_1816,N_1486,N_1367);
xor U1817 (N_1817,N_1618,N_1301);
xnor U1818 (N_1818,N_1547,N_1212);
xnor U1819 (N_1819,N_1791,N_1431);
or U1820 (N_1820,N_1328,N_1797);
xor U1821 (N_1821,N_1231,N_1583);
nor U1822 (N_1822,N_1278,N_1430);
or U1823 (N_1823,N_1629,N_1352);
or U1824 (N_1824,N_1242,N_1648);
xor U1825 (N_1825,N_1545,N_1685);
nand U1826 (N_1826,N_1306,N_1731);
and U1827 (N_1827,N_1245,N_1738);
and U1828 (N_1828,N_1377,N_1207);
xnor U1829 (N_1829,N_1234,N_1259);
or U1830 (N_1830,N_1502,N_1365);
and U1831 (N_1831,N_1356,N_1669);
and U1832 (N_1832,N_1476,N_1753);
and U1833 (N_1833,N_1413,N_1334);
or U1834 (N_1834,N_1787,N_1758);
xnor U1835 (N_1835,N_1415,N_1261);
and U1836 (N_1836,N_1490,N_1247);
and U1837 (N_1837,N_1639,N_1390);
nand U1838 (N_1838,N_1273,N_1578);
nor U1839 (N_1839,N_1748,N_1354);
or U1840 (N_1840,N_1751,N_1315);
xnor U1841 (N_1841,N_1345,N_1517);
nand U1842 (N_1842,N_1469,N_1760);
or U1843 (N_1843,N_1655,N_1628);
xnor U1844 (N_1844,N_1224,N_1551);
nor U1845 (N_1845,N_1577,N_1603);
nand U1846 (N_1846,N_1684,N_1205);
or U1847 (N_1847,N_1200,N_1590);
nor U1848 (N_1848,N_1601,N_1719);
or U1849 (N_1849,N_1682,N_1470);
nor U1850 (N_1850,N_1265,N_1371);
or U1851 (N_1851,N_1796,N_1454);
or U1852 (N_1852,N_1249,N_1457);
and U1853 (N_1853,N_1699,N_1398);
xor U1854 (N_1854,N_1269,N_1262);
nand U1855 (N_1855,N_1712,N_1335);
and U1856 (N_1856,N_1794,N_1724);
or U1857 (N_1857,N_1539,N_1664);
nor U1858 (N_1858,N_1680,N_1586);
nor U1859 (N_1859,N_1492,N_1533);
nand U1860 (N_1860,N_1402,N_1216);
and U1861 (N_1861,N_1323,N_1624);
nand U1862 (N_1862,N_1757,N_1737);
nand U1863 (N_1863,N_1686,N_1666);
and U1864 (N_1864,N_1777,N_1244);
nor U1865 (N_1865,N_1725,N_1310);
nand U1866 (N_1866,N_1728,N_1373);
xnor U1867 (N_1867,N_1581,N_1732);
and U1868 (N_1868,N_1561,N_1213);
and U1869 (N_1869,N_1348,N_1764);
nand U1870 (N_1870,N_1425,N_1589);
or U1871 (N_1871,N_1564,N_1579);
nor U1872 (N_1872,N_1297,N_1511);
nor U1873 (N_1873,N_1246,N_1752);
nor U1874 (N_1874,N_1597,N_1339);
and U1875 (N_1875,N_1455,N_1754);
nor U1876 (N_1876,N_1575,N_1562);
xor U1877 (N_1877,N_1366,N_1556);
or U1878 (N_1878,N_1745,N_1295);
nor U1879 (N_1879,N_1694,N_1636);
xor U1880 (N_1880,N_1223,N_1474);
and U1881 (N_1881,N_1678,N_1277);
nor U1882 (N_1882,N_1765,N_1567);
or U1883 (N_1883,N_1203,N_1483);
nand U1884 (N_1884,N_1710,N_1656);
or U1885 (N_1885,N_1341,N_1633);
nor U1886 (N_1886,N_1617,N_1351);
nand U1887 (N_1887,N_1689,N_1419);
or U1888 (N_1888,N_1433,N_1228);
and U1889 (N_1889,N_1784,N_1641);
nand U1890 (N_1890,N_1608,N_1282);
nand U1891 (N_1891,N_1414,N_1549);
and U1892 (N_1892,N_1347,N_1535);
nand U1893 (N_1893,N_1604,N_1225);
xnor U1894 (N_1894,N_1622,N_1485);
and U1895 (N_1895,N_1400,N_1467);
and U1896 (N_1896,N_1344,N_1670);
nor U1897 (N_1897,N_1741,N_1210);
or U1898 (N_1898,N_1538,N_1683);
or U1899 (N_1899,N_1333,N_1250);
nor U1900 (N_1900,N_1294,N_1593);
nand U1901 (N_1901,N_1755,N_1598);
nor U1902 (N_1902,N_1226,N_1704);
and U1903 (N_1903,N_1392,N_1720);
and U1904 (N_1904,N_1441,N_1771);
and U1905 (N_1905,N_1709,N_1506);
nor U1906 (N_1906,N_1337,N_1342);
or U1907 (N_1907,N_1667,N_1461);
or U1908 (N_1908,N_1388,N_1369);
and U1909 (N_1909,N_1509,N_1449);
or U1910 (N_1910,N_1375,N_1465);
and U1911 (N_1911,N_1254,N_1240);
nor U1912 (N_1912,N_1293,N_1411);
and U1913 (N_1913,N_1463,N_1627);
nand U1914 (N_1914,N_1436,N_1255);
and U1915 (N_1915,N_1421,N_1632);
or U1916 (N_1916,N_1279,N_1512);
nand U1917 (N_1917,N_1498,N_1767);
and U1918 (N_1918,N_1355,N_1391);
and U1919 (N_1919,N_1364,N_1493);
or U1920 (N_1920,N_1500,N_1582);
or U1921 (N_1921,N_1241,N_1239);
and U1922 (N_1922,N_1514,N_1299);
xnor U1923 (N_1923,N_1396,N_1770);
xnor U1924 (N_1924,N_1734,N_1705);
nand U1925 (N_1925,N_1527,N_1427);
and U1926 (N_1926,N_1762,N_1360);
and U1927 (N_1927,N_1651,N_1251);
or U1928 (N_1928,N_1769,N_1256);
nor U1929 (N_1929,N_1437,N_1275);
nand U1930 (N_1930,N_1588,N_1574);
and U1931 (N_1931,N_1473,N_1580);
and U1932 (N_1932,N_1599,N_1384);
nand U1933 (N_1933,N_1718,N_1422);
and U1934 (N_1934,N_1510,N_1326);
and U1935 (N_1935,N_1280,N_1729);
nand U1936 (N_1936,N_1218,N_1291);
nor U1937 (N_1937,N_1494,N_1495);
nor U1938 (N_1938,N_1565,N_1663);
nor U1939 (N_1939,N_1635,N_1215);
xnor U1940 (N_1940,N_1443,N_1585);
and U1941 (N_1941,N_1503,N_1550);
and U1942 (N_1942,N_1343,N_1202);
nor U1943 (N_1943,N_1573,N_1222);
nand U1944 (N_1944,N_1448,N_1372);
nor U1945 (N_1945,N_1672,N_1761);
or U1946 (N_1946,N_1359,N_1605);
xor U1947 (N_1947,N_1558,N_1401);
nor U1948 (N_1948,N_1692,N_1717);
xnor U1949 (N_1949,N_1206,N_1385);
nand U1950 (N_1950,N_1479,N_1320);
nand U1951 (N_1951,N_1412,N_1795);
nand U1952 (N_1952,N_1743,N_1650);
nand U1953 (N_1953,N_1687,N_1319);
nor U1954 (N_1954,N_1541,N_1393);
or U1955 (N_1955,N_1453,N_1395);
nor U1956 (N_1956,N_1721,N_1768);
nand U1957 (N_1957,N_1735,N_1270);
nor U1958 (N_1958,N_1505,N_1304);
nor U1959 (N_1959,N_1303,N_1418);
and U1960 (N_1960,N_1288,N_1480);
nand U1961 (N_1961,N_1285,N_1524);
or U1962 (N_1962,N_1518,N_1232);
nand U1963 (N_1963,N_1563,N_1370);
and U1964 (N_1964,N_1477,N_1526);
nor U1965 (N_1965,N_1349,N_1708);
and U1966 (N_1966,N_1296,N_1357);
nand U1967 (N_1967,N_1338,N_1475);
xnor U1968 (N_1968,N_1759,N_1271);
and U1969 (N_1969,N_1286,N_1706);
or U1970 (N_1970,N_1445,N_1253);
or U1971 (N_1971,N_1774,N_1410);
nand U1972 (N_1972,N_1610,N_1466);
nand U1973 (N_1973,N_1432,N_1733);
nand U1974 (N_1974,N_1657,N_1625);
nand U1975 (N_1975,N_1233,N_1267);
and U1976 (N_1976,N_1688,N_1642);
and U1977 (N_1977,N_1560,N_1317);
xor U1978 (N_1978,N_1727,N_1438);
nor U1979 (N_1979,N_1464,N_1281);
xnor U1980 (N_1980,N_1647,N_1658);
or U1981 (N_1981,N_1715,N_1525);
nor U1982 (N_1982,N_1340,N_1272);
xor U1983 (N_1983,N_1609,N_1460);
nor U1984 (N_1984,N_1504,N_1350);
or U1985 (N_1985,N_1792,N_1543);
or U1986 (N_1986,N_1363,N_1209);
xor U1987 (N_1987,N_1798,N_1450);
and U1988 (N_1988,N_1302,N_1287);
nand U1989 (N_1989,N_1536,N_1446);
nor U1990 (N_1990,N_1435,N_1481);
nor U1991 (N_1991,N_1230,N_1429);
and U1992 (N_1992,N_1615,N_1379);
nand U1993 (N_1993,N_1530,N_1440);
nor U1994 (N_1994,N_1221,N_1386);
nor U1995 (N_1995,N_1331,N_1723);
nor U1996 (N_1996,N_1631,N_1746);
nand U1997 (N_1997,N_1491,N_1204);
nor U1998 (N_1998,N_1730,N_1529);
and U1999 (N_1999,N_1559,N_1776);
nor U2000 (N_2000,N_1644,N_1660);
nor U2001 (N_2001,N_1569,N_1546);
or U2002 (N_2002,N_1659,N_1703);
nand U2003 (N_2003,N_1522,N_1638);
nand U2004 (N_2004,N_1621,N_1566);
or U2005 (N_2005,N_1607,N_1691);
nand U2006 (N_2006,N_1534,N_1778);
nor U2007 (N_2007,N_1264,N_1308);
or U2008 (N_2008,N_1693,N_1309);
and U2009 (N_2009,N_1406,N_1346);
and U2010 (N_2010,N_1300,N_1380);
nor U2011 (N_2011,N_1654,N_1596);
nand U2012 (N_2012,N_1362,N_1358);
and U2013 (N_2013,N_1389,N_1668);
and U2014 (N_2014,N_1726,N_1488);
nand U2015 (N_2015,N_1750,N_1417);
nand U2016 (N_2016,N_1788,N_1217);
xor U2017 (N_2017,N_1677,N_1439);
or U2018 (N_2018,N_1520,N_1637);
nor U2019 (N_2019,N_1742,N_1416);
and U2020 (N_2020,N_1653,N_1555);
or U2021 (N_2021,N_1507,N_1674);
nand U2022 (N_2022,N_1652,N_1258);
nand U2023 (N_2023,N_1749,N_1387);
or U2024 (N_2024,N_1274,N_1284);
and U2025 (N_2025,N_1252,N_1489);
or U2026 (N_2026,N_1236,N_1201);
nand U2027 (N_2027,N_1766,N_1235);
xor U2028 (N_2028,N_1785,N_1790);
nand U2029 (N_2029,N_1591,N_1747);
nand U2030 (N_2030,N_1508,N_1404);
nor U2031 (N_2031,N_1576,N_1472);
nor U2032 (N_2032,N_1214,N_1515);
or U2033 (N_2033,N_1698,N_1403);
nand U2034 (N_2034,N_1459,N_1643);
and U2035 (N_2035,N_1501,N_1697);
and U2036 (N_2036,N_1312,N_1553);
nand U2037 (N_2037,N_1711,N_1613);
or U2038 (N_2038,N_1513,N_1786);
nor U2039 (N_2039,N_1484,N_1531);
nand U2040 (N_2040,N_1487,N_1673);
nor U2041 (N_2041,N_1521,N_1447);
nor U2042 (N_2042,N_1313,N_1211);
or U2043 (N_2043,N_1557,N_1707);
xor U2044 (N_2044,N_1740,N_1584);
and U2045 (N_2045,N_1257,N_1736);
or U2046 (N_2046,N_1260,N_1744);
nor U2047 (N_2047,N_1763,N_1516);
and U2048 (N_2048,N_1540,N_1671);
nor U2049 (N_2049,N_1458,N_1681);
nor U2050 (N_2050,N_1544,N_1452);
and U2051 (N_2051,N_1793,N_1570);
nor U2052 (N_2052,N_1321,N_1614);
and U2053 (N_2053,N_1773,N_1383);
xor U2054 (N_2054,N_1661,N_1568);
nand U2055 (N_2055,N_1376,N_1528);
nor U2056 (N_2056,N_1420,N_1519);
and U2057 (N_2057,N_1789,N_1662);
or U2058 (N_2058,N_1409,N_1263);
nand U2059 (N_2059,N_1423,N_1756);
or U2060 (N_2060,N_1592,N_1336);
or U2061 (N_2061,N_1399,N_1537);
nand U2062 (N_2062,N_1451,N_1602);
and U2063 (N_2063,N_1322,N_1595);
nand U2064 (N_2064,N_1276,N_1665);
nor U2065 (N_2065,N_1397,N_1571);
or U2066 (N_2066,N_1314,N_1318);
or U2067 (N_2067,N_1290,N_1623);
and U2068 (N_2068,N_1649,N_1552);
or U2069 (N_2069,N_1779,N_1434);
or U2070 (N_2070,N_1307,N_1594);
nor U2071 (N_2071,N_1587,N_1626);
or U2072 (N_2072,N_1243,N_1620);
or U2073 (N_2073,N_1311,N_1482);
nor U2074 (N_2074,N_1332,N_1700);
nand U2075 (N_2075,N_1325,N_1283);
and U2076 (N_2076,N_1378,N_1600);
nand U2077 (N_2077,N_1634,N_1227);
nor U2078 (N_2078,N_1523,N_1329);
and U2079 (N_2079,N_1238,N_1676);
xnor U2080 (N_2080,N_1442,N_1690);
nor U2081 (N_2081,N_1237,N_1532);
nor U2082 (N_2082,N_1468,N_1353);
nand U2083 (N_2083,N_1268,N_1407);
xnor U2084 (N_2084,N_1619,N_1646);
nor U2085 (N_2085,N_1496,N_1640);
and U2086 (N_2086,N_1229,N_1780);
xnor U2087 (N_2087,N_1702,N_1499);
and U2088 (N_2088,N_1374,N_1382);
or U2089 (N_2089,N_1714,N_1713);
nand U2090 (N_2090,N_1292,N_1368);
and U2091 (N_2091,N_1606,N_1630);
and U2092 (N_2092,N_1305,N_1471);
nor U2093 (N_2093,N_1722,N_1554);
and U2094 (N_2094,N_1572,N_1695);
and U2095 (N_2095,N_1548,N_1497);
or U2096 (N_2096,N_1462,N_1775);
nand U2097 (N_2097,N_1612,N_1611);
nand U2098 (N_2098,N_1783,N_1456);
and U2099 (N_2099,N_1220,N_1444);
xnor U2100 (N_2100,N_1777,N_1529);
and U2101 (N_2101,N_1408,N_1486);
nand U2102 (N_2102,N_1721,N_1670);
nand U2103 (N_2103,N_1611,N_1411);
nor U2104 (N_2104,N_1760,N_1529);
nand U2105 (N_2105,N_1258,N_1361);
xor U2106 (N_2106,N_1287,N_1616);
nand U2107 (N_2107,N_1675,N_1605);
and U2108 (N_2108,N_1617,N_1779);
nor U2109 (N_2109,N_1211,N_1661);
or U2110 (N_2110,N_1401,N_1734);
and U2111 (N_2111,N_1717,N_1446);
nand U2112 (N_2112,N_1291,N_1420);
nor U2113 (N_2113,N_1617,N_1732);
and U2114 (N_2114,N_1640,N_1395);
nand U2115 (N_2115,N_1526,N_1395);
or U2116 (N_2116,N_1401,N_1762);
nand U2117 (N_2117,N_1320,N_1604);
xnor U2118 (N_2118,N_1415,N_1695);
nor U2119 (N_2119,N_1691,N_1743);
nor U2120 (N_2120,N_1355,N_1319);
xnor U2121 (N_2121,N_1594,N_1451);
nand U2122 (N_2122,N_1766,N_1293);
nand U2123 (N_2123,N_1399,N_1267);
nor U2124 (N_2124,N_1724,N_1755);
nand U2125 (N_2125,N_1641,N_1376);
nor U2126 (N_2126,N_1492,N_1553);
or U2127 (N_2127,N_1487,N_1798);
or U2128 (N_2128,N_1752,N_1661);
or U2129 (N_2129,N_1407,N_1469);
nand U2130 (N_2130,N_1628,N_1328);
and U2131 (N_2131,N_1661,N_1475);
and U2132 (N_2132,N_1700,N_1625);
and U2133 (N_2133,N_1577,N_1334);
or U2134 (N_2134,N_1511,N_1304);
xnor U2135 (N_2135,N_1717,N_1203);
nand U2136 (N_2136,N_1571,N_1458);
or U2137 (N_2137,N_1555,N_1217);
nand U2138 (N_2138,N_1325,N_1348);
or U2139 (N_2139,N_1330,N_1239);
and U2140 (N_2140,N_1732,N_1399);
and U2141 (N_2141,N_1662,N_1538);
nand U2142 (N_2142,N_1209,N_1607);
nor U2143 (N_2143,N_1492,N_1585);
nor U2144 (N_2144,N_1288,N_1349);
or U2145 (N_2145,N_1508,N_1708);
nor U2146 (N_2146,N_1711,N_1688);
or U2147 (N_2147,N_1562,N_1492);
or U2148 (N_2148,N_1716,N_1709);
and U2149 (N_2149,N_1589,N_1279);
or U2150 (N_2150,N_1778,N_1630);
nand U2151 (N_2151,N_1779,N_1713);
nand U2152 (N_2152,N_1510,N_1703);
nor U2153 (N_2153,N_1511,N_1435);
nor U2154 (N_2154,N_1743,N_1304);
nand U2155 (N_2155,N_1745,N_1214);
nor U2156 (N_2156,N_1724,N_1595);
and U2157 (N_2157,N_1265,N_1215);
xor U2158 (N_2158,N_1434,N_1432);
xnor U2159 (N_2159,N_1469,N_1384);
or U2160 (N_2160,N_1215,N_1347);
nand U2161 (N_2161,N_1669,N_1608);
and U2162 (N_2162,N_1765,N_1242);
nor U2163 (N_2163,N_1641,N_1589);
nor U2164 (N_2164,N_1748,N_1236);
or U2165 (N_2165,N_1411,N_1758);
or U2166 (N_2166,N_1374,N_1543);
nand U2167 (N_2167,N_1334,N_1478);
or U2168 (N_2168,N_1510,N_1799);
nor U2169 (N_2169,N_1520,N_1676);
or U2170 (N_2170,N_1246,N_1483);
xnor U2171 (N_2171,N_1256,N_1729);
xor U2172 (N_2172,N_1727,N_1545);
nand U2173 (N_2173,N_1459,N_1240);
and U2174 (N_2174,N_1518,N_1771);
or U2175 (N_2175,N_1466,N_1278);
nor U2176 (N_2176,N_1520,N_1678);
and U2177 (N_2177,N_1321,N_1580);
and U2178 (N_2178,N_1316,N_1532);
nand U2179 (N_2179,N_1219,N_1569);
nand U2180 (N_2180,N_1656,N_1441);
xor U2181 (N_2181,N_1643,N_1509);
nand U2182 (N_2182,N_1449,N_1448);
xnor U2183 (N_2183,N_1606,N_1223);
or U2184 (N_2184,N_1451,N_1591);
xnor U2185 (N_2185,N_1609,N_1620);
and U2186 (N_2186,N_1346,N_1267);
nor U2187 (N_2187,N_1454,N_1586);
nor U2188 (N_2188,N_1515,N_1597);
nor U2189 (N_2189,N_1458,N_1560);
nor U2190 (N_2190,N_1689,N_1209);
nand U2191 (N_2191,N_1512,N_1351);
xnor U2192 (N_2192,N_1388,N_1352);
nand U2193 (N_2193,N_1573,N_1520);
nand U2194 (N_2194,N_1578,N_1535);
nor U2195 (N_2195,N_1631,N_1506);
or U2196 (N_2196,N_1454,N_1455);
or U2197 (N_2197,N_1727,N_1771);
and U2198 (N_2198,N_1728,N_1221);
nand U2199 (N_2199,N_1389,N_1795);
xnor U2200 (N_2200,N_1646,N_1256);
nand U2201 (N_2201,N_1432,N_1618);
nand U2202 (N_2202,N_1753,N_1294);
nor U2203 (N_2203,N_1728,N_1734);
nand U2204 (N_2204,N_1666,N_1783);
and U2205 (N_2205,N_1769,N_1220);
and U2206 (N_2206,N_1618,N_1575);
nand U2207 (N_2207,N_1776,N_1659);
and U2208 (N_2208,N_1667,N_1659);
nor U2209 (N_2209,N_1433,N_1777);
nand U2210 (N_2210,N_1500,N_1597);
or U2211 (N_2211,N_1712,N_1387);
and U2212 (N_2212,N_1443,N_1656);
and U2213 (N_2213,N_1416,N_1773);
nand U2214 (N_2214,N_1454,N_1529);
nand U2215 (N_2215,N_1278,N_1666);
or U2216 (N_2216,N_1281,N_1462);
and U2217 (N_2217,N_1525,N_1612);
and U2218 (N_2218,N_1739,N_1600);
or U2219 (N_2219,N_1750,N_1435);
and U2220 (N_2220,N_1491,N_1315);
nand U2221 (N_2221,N_1200,N_1690);
nand U2222 (N_2222,N_1642,N_1470);
or U2223 (N_2223,N_1628,N_1411);
and U2224 (N_2224,N_1782,N_1592);
nor U2225 (N_2225,N_1595,N_1630);
xor U2226 (N_2226,N_1635,N_1734);
and U2227 (N_2227,N_1682,N_1485);
nand U2228 (N_2228,N_1782,N_1714);
xnor U2229 (N_2229,N_1724,N_1511);
xnor U2230 (N_2230,N_1248,N_1781);
nand U2231 (N_2231,N_1563,N_1312);
and U2232 (N_2232,N_1618,N_1719);
and U2233 (N_2233,N_1299,N_1795);
and U2234 (N_2234,N_1361,N_1580);
and U2235 (N_2235,N_1789,N_1524);
nand U2236 (N_2236,N_1657,N_1663);
nand U2237 (N_2237,N_1289,N_1584);
nand U2238 (N_2238,N_1747,N_1755);
or U2239 (N_2239,N_1275,N_1456);
xor U2240 (N_2240,N_1561,N_1635);
nand U2241 (N_2241,N_1549,N_1574);
xor U2242 (N_2242,N_1615,N_1402);
nand U2243 (N_2243,N_1723,N_1470);
or U2244 (N_2244,N_1434,N_1382);
or U2245 (N_2245,N_1410,N_1595);
or U2246 (N_2246,N_1458,N_1616);
and U2247 (N_2247,N_1387,N_1349);
and U2248 (N_2248,N_1625,N_1470);
nand U2249 (N_2249,N_1405,N_1282);
and U2250 (N_2250,N_1577,N_1600);
nor U2251 (N_2251,N_1533,N_1707);
or U2252 (N_2252,N_1281,N_1316);
nand U2253 (N_2253,N_1212,N_1460);
nor U2254 (N_2254,N_1431,N_1708);
and U2255 (N_2255,N_1357,N_1556);
and U2256 (N_2256,N_1763,N_1260);
xor U2257 (N_2257,N_1717,N_1704);
nand U2258 (N_2258,N_1705,N_1447);
nand U2259 (N_2259,N_1514,N_1235);
nor U2260 (N_2260,N_1411,N_1765);
or U2261 (N_2261,N_1614,N_1292);
or U2262 (N_2262,N_1700,N_1638);
and U2263 (N_2263,N_1446,N_1398);
nand U2264 (N_2264,N_1360,N_1271);
nand U2265 (N_2265,N_1483,N_1540);
or U2266 (N_2266,N_1729,N_1429);
nor U2267 (N_2267,N_1739,N_1520);
nand U2268 (N_2268,N_1234,N_1734);
or U2269 (N_2269,N_1694,N_1441);
nand U2270 (N_2270,N_1478,N_1651);
nor U2271 (N_2271,N_1313,N_1517);
or U2272 (N_2272,N_1335,N_1333);
and U2273 (N_2273,N_1676,N_1270);
or U2274 (N_2274,N_1258,N_1376);
nand U2275 (N_2275,N_1666,N_1461);
nor U2276 (N_2276,N_1483,N_1423);
and U2277 (N_2277,N_1479,N_1708);
or U2278 (N_2278,N_1617,N_1381);
nor U2279 (N_2279,N_1691,N_1732);
nand U2280 (N_2280,N_1285,N_1744);
and U2281 (N_2281,N_1232,N_1343);
nand U2282 (N_2282,N_1692,N_1645);
nand U2283 (N_2283,N_1764,N_1666);
nand U2284 (N_2284,N_1755,N_1568);
and U2285 (N_2285,N_1608,N_1656);
or U2286 (N_2286,N_1379,N_1306);
nand U2287 (N_2287,N_1724,N_1532);
and U2288 (N_2288,N_1398,N_1762);
or U2289 (N_2289,N_1472,N_1281);
nor U2290 (N_2290,N_1390,N_1223);
and U2291 (N_2291,N_1283,N_1267);
and U2292 (N_2292,N_1799,N_1708);
nand U2293 (N_2293,N_1731,N_1552);
or U2294 (N_2294,N_1253,N_1511);
nand U2295 (N_2295,N_1743,N_1267);
nor U2296 (N_2296,N_1574,N_1652);
nor U2297 (N_2297,N_1738,N_1201);
nand U2298 (N_2298,N_1572,N_1293);
nand U2299 (N_2299,N_1281,N_1618);
xnor U2300 (N_2300,N_1658,N_1670);
nor U2301 (N_2301,N_1565,N_1479);
or U2302 (N_2302,N_1446,N_1649);
nand U2303 (N_2303,N_1714,N_1500);
nor U2304 (N_2304,N_1304,N_1485);
nand U2305 (N_2305,N_1200,N_1396);
nor U2306 (N_2306,N_1784,N_1518);
or U2307 (N_2307,N_1223,N_1412);
and U2308 (N_2308,N_1517,N_1296);
or U2309 (N_2309,N_1561,N_1671);
nand U2310 (N_2310,N_1676,N_1667);
nand U2311 (N_2311,N_1409,N_1243);
and U2312 (N_2312,N_1495,N_1260);
or U2313 (N_2313,N_1784,N_1324);
nor U2314 (N_2314,N_1642,N_1266);
nand U2315 (N_2315,N_1335,N_1483);
nand U2316 (N_2316,N_1708,N_1615);
nand U2317 (N_2317,N_1206,N_1339);
nand U2318 (N_2318,N_1608,N_1277);
nor U2319 (N_2319,N_1208,N_1726);
or U2320 (N_2320,N_1226,N_1387);
xor U2321 (N_2321,N_1794,N_1722);
xnor U2322 (N_2322,N_1443,N_1276);
or U2323 (N_2323,N_1653,N_1634);
nand U2324 (N_2324,N_1798,N_1329);
nor U2325 (N_2325,N_1592,N_1653);
nand U2326 (N_2326,N_1639,N_1764);
nand U2327 (N_2327,N_1382,N_1384);
and U2328 (N_2328,N_1200,N_1731);
and U2329 (N_2329,N_1244,N_1606);
xnor U2330 (N_2330,N_1402,N_1435);
nor U2331 (N_2331,N_1538,N_1686);
nor U2332 (N_2332,N_1273,N_1442);
nand U2333 (N_2333,N_1462,N_1280);
nand U2334 (N_2334,N_1716,N_1769);
xnor U2335 (N_2335,N_1638,N_1352);
nor U2336 (N_2336,N_1239,N_1755);
or U2337 (N_2337,N_1749,N_1722);
nor U2338 (N_2338,N_1789,N_1390);
nand U2339 (N_2339,N_1625,N_1638);
nand U2340 (N_2340,N_1519,N_1540);
nor U2341 (N_2341,N_1623,N_1216);
and U2342 (N_2342,N_1725,N_1645);
and U2343 (N_2343,N_1396,N_1295);
or U2344 (N_2344,N_1327,N_1343);
nand U2345 (N_2345,N_1293,N_1556);
nand U2346 (N_2346,N_1386,N_1545);
xor U2347 (N_2347,N_1652,N_1522);
xnor U2348 (N_2348,N_1419,N_1213);
and U2349 (N_2349,N_1478,N_1453);
xor U2350 (N_2350,N_1234,N_1717);
and U2351 (N_2351,N_1278,N_1617);
and U2352 (N_2352,N_1596,N_1650);
or U2353 (N_2353,N_1275,N_1377);
and U2354 (N_2354,N_1783,N_1214);
nand U2355 (N_2355,N_1760,N_1713);
nor U2356 (N_2356,N_1313,N_1372);
nor U2357 (N_2357,N_1446,N_1421);
and U2358 (N_2358,N_1740,N_1764);
nor U2359 (N_2359,N_1794,N_1454);
and U2360 (N_2360,N_1266,N_1281);
nand U2361 (N_2361,N_1242,N_1787);
xor U2362 (N_2362,N_1560,N_1224);
and U2363 (N_2363,N_1654,N_1256);
nand U2364 (N_2364,N_1512,N_1292);
and U2365 (N_2365,N_1679,N_1615);
or U2366 (N_2366,N_1626,N_1296);
and U2367 (N_2367,N_1634,N_1689);
nand U2368 (N_2368,N_1788,N_1522);
and U2369 (N_2369,N_1571,N_1319);
or U2370 (N_2370,N_1764,N_1571);
nor U2371 (N_2371,N_1778,N_1459);
or U2372 (N_2372,N_1599,N_1488);
and U2373 (N_2373,N_1594,N_1663);
and U2374 (N_2374,N_1513,N_1725);
nor U2375 (N_2375,N_1425,N_1711);
or U2376 (N_2376,N_1620,N_1618);
nor U2377 (N_2377,N_1225,N_1592);
nand U2378 (N_2378,N_1582,N_1435);
nor U2379 (N_2379,N_1281,N_1641);
nor U2380 (N_2380,N_1246,N_1758);
xnor U2381 (N_2381,N_1621,N_1582);
nor U2382 (N_2382,N_1765,N_1649);
or U2383 (N_2383,N_1648,N_1614);
nand U2384 (N_2384,N_1507,N_1349);
xnor U2385 (N_2385,N_1431,N_1481);
xor U2386 (N_2386,N_1223,N_1538);
nor U2387 (N_2387,N_1395,N_1333);
or U2388 (N_2388,N_1329,N_1435);
and U2389 (N_2389,N_1439,N_1698);
or U2390 (N_2390,N_1322,N_1386);
nor U2391 (N_2391,N_1475,N_1479);
xor U2392 (N_2392,N_1635,N_1639);
nor U2393 (N_2393,N_1580,N_1271);
or U2394 (N_2394,N_1646,N_1225);
or U2395 (N_2395,N_1687,N_1606);
or U2396 (N_2396,N_1625,N_1771);
and U2397 (N_2397,N_1646,N_1677);
nand U2398 (N_2398,N_1654,N_1466);
nand U2399 (N_2399,N_1762,N_1295);
and U2400 (N_2400,N_1808,N_1893);
nor U2401 (N_2401,N_2243,N_1887);
nor U2402 (N_2402,N_2013,N_2119);
nand U2403 (N_2403,N_1918,N_2066);
or U2404 (N_2404,N_2394,N_1870);
nor U2405 (N_2405,N_2020,N_2374);
nand U2406 (N_2406,N_2065,N_2152);
nand U2407 (N_2407,N_2171,N_2354);
and U2408 (N_2408,N_1980,N_2241);
and U2409 (N_2409,N_2036,N_2068);
xnor U2410 (N_2410,N_1902,N_1979);
nor U2411 (N_2411,N_2052,N_2247);
or U2412 (N_2412,N_1842,N_2115);
nor U2413 (N_2413,N_2064,N_2028);
or U2414 (N_2414,N_1818,N_1996);
xor U2415 (N_2415,N_2378,N_2251);
nand U2416 (N_2416,N_2387,N_1803);
nor U2417 (N_2417,N_2209,N_2039);
or U2418 (N_2418,N_1827,N_2325);
xor U2419 (N_2419,N_2099,N_1913);
nand U2420 (N_2420,N_1961,N_2193);
nand U2421 (N_2421,N_1800,N_2238);
or U2422 (N_2422,N_1978,N_2163);
nand U2423 (N_2423,N_2026,N_2205);
or U2424 (N_2424,N_2058,N_2141);
nand U2425 (N_2425,N_2321,N_2237);
or U2426 (N_2426,N_2273,N_2051);
and U2427 (N_2427,N_2023,N_2083);
and U2428 (N_2428,N_2173,N_2148);
or U2429 (N_2429,N_2264,N_2153);
and U2430 (N_2430,N_2085,N_2226);
nand U2431 (N_2431,N_2197,N_2343);
and U2432 (N_2432,N_2130,N_1891);
and U2433 (N_2433,N_1998,N_2244);
or U2434 (N_2434,N_2118,N_1817);
or U2435 (N_2435,N_2363,N_2348);
nor U2436 (N_2436,N_1855,N_2090);
and U2437 (N_2437,N_2249,N_2033);
xnor U2438 (N_2438,N_1850,N_1879);
or U2439 (N_2439,N_2042,N_2071);
nor U2440 (N_2440,N_2196,N_1819);
and U2441 (N_2441,N_1853,N_2109);
or U2442 (N_2442,N_1858,N_2259);
nand U2443 (N_2443,N_2011,N_2035);
nor U2444 (N_2444,N_2157,N_2313);
nand U2445 (N_2445,N_1851,N_2038);
nor U2446 (N_2446,N_2124,N_2345);
or U2447 (N_2447,N_2088,N_2166);
and U2448 (N_2448,N_1824,N_1992);
xor U2449 (N_2449,N_2175,N_2139);
and U2450 (N_2450,N_2395,N_1954);
nand U2451 (N_2451,N_2017,N_2281);
nand U2452 (N_2452,N_2122,N_1971);
xor U2453 (N_2453,N_2257,N_2303);
nand U2454 (N_2454,N_1991,N_2311);
xor U2455 (N_2455,N_2194,N_2106);
nand U2456 (N_2456,N_2270,N_2239);
or U2457 (N_2457,N_2199,N_1906);
xnor U2458 (N_2458,N_1890,N_2108);
or U2459 (N_2459,N_2304,N_1936);
nand U2460 (N_2460,N_2168,N_2097);
nor U2461 (N_2461,N_1865,N_1986);
and U2462 (N_2462,N_2004,N_1934);
and U2463 (N_2463,N_1895,N_2302);
xor U2464 (N_2464,N_2120,N_1888);
and U2465 (N_2465,N_2265,N_1812);
or U2466 (N_2466,N_2396,N_2006);
and U2467 (N_2467,N_2263,N_1944);
nand U2468 (N_2468,N_2008,N_2382);
nor U2469 (N_2469,N_2350,N_1881);
and U2470 (N_2470,N_1814,N_2138);
nand U2471 (N_2471,N_2339,N_2332);
nand U2472 (N_2472,N_1901,N_1805);
nor U2473 (N_2473,N_2142,N_2292);
or U2474 (N_2474,N_2346,N_1951);
xor U2475 (N_2475,N_2319,N_2369);
or U2476 (N_2476,N_1833,N_2105);
nor U2477 (N_2477,N_2001,N_1928);
or U2478 (N_2478,N_1802,N_2094);
nand U2479 (N_2479,N_2208,N_1903);
or U2480 (N_2480,N_2131,N_1924);
nor U2481 (N_2481,N_2132,N_2082);
and U2482 (N_2482,N_2310,N_2164);
or U2483 (N_2483,N_2268,N_1969);
nand U2484 (N_2484,N_2383,N_1874);
xor U2485 (N_2485,N_2136,N_2341);
nor U2486 (N_2486,N_1860,N_2025);
nand U2487 (N_2487,N_2254,N_2252);
and U2488 (N_2488,N_1941,N_2024);
nor U2489 (N_2489,N_2046,N_2112);
or U2490 (N_2490,N_1958,N_1880);
nand U2491 (N_2491,N_2328,N_2358);
and U2492 (N_2492,N_1939,N_2117);
or U2493 (N_2493,N_1873,N_1857);
or U2494 (N_2494,N_1830,N_2338);
nor U2495 (N_2495,N_1810,N_1862);
nand U2496 (N_2496,N_2312,N_1963);
nand U2497 (N_2497,N_1999,N_2127);
nand U2498 (N_2498,N_1977,N_2022);
xor U2499 (N_2499,N_2393,N_1844);
or U2500 (N_2500,N_2352,N_2256);
or U2501 (N_2501,N_2329,N_2289);
or U2502 (N_2502,N_1972,N_2018);
nor U2503 (N_2503,N_2231,N_1975);
and U2504 (N_2504,N_2384,N_2169);
and U2505 (N_2505,N_1922,N_2074);
nor U2506 (N_2506,N_2297,N_2372);
and U2507 (N_2507,N_1942,N_2323);
or U2508 (N_2508,N_2335,N_2326);
nand U2509 (N_2509,N_2182,N_2217);
xnor U2510 (N_2510,N_1867,N_1920);
nand U2511 (N_2511,N_2162,N_1875);
nor U2512 (N_2512,N_2062,N_2373);
nand U2513 (N_2513,N_1987,N_2151);
nor U2514 (N_2514,N_2044,N_2388);
and U2515 (N_2515,N_1856,N_2050);
nor U2516 (N_2516,N_2353,N_1957);
or U2517 (N_2517,N_2399,N_1848);
nor U2518 (N_2518,N_2092,N_2188);
or U2519 (N_2519,N_2361,N_1876);
nor U2520 (N_2520,N_1912,N_2207);
or U2521 (N_2521,N_2056,N_2084);
and U2522 (N_2522,N_2320,N_2245);
or U2523 (N_2523,N_2377,N_2049);
nand U2524 (N_2524,N_2055,N_2053);
and U2525 (N_2525,N_2144,N_2293);
nand U2526 (N_2526,N_2314,N_2041);
or U2527 (N_2527,N_2288,N_2306);
nand U2528 (N_2528,N_2126,N_2296);
xor U2529 (N_2529,N_2103,N_2043);
nand U2530 (N_2530,N_1915,N_2216);
nand U2531 (N_2531,N_2309,N_2047);
nand U2532 (N_2532,N_2159,N_1836);
nor U2533 (N_2533,N_2375,N_1976);
and U2534 (N_2534,N_1866,N_2331);
xnor U2535 (N_2535,N_1948,N_1863);
nand U2536 (N_2536,N_2307,N_2275);
and U2537 (N_2537,N_2299,N_2308);
nor U2538 (N_2538,N_2386,N_1984);
nand U2539 (N_2539,N_1923,N_1806);
and U2540 (N_2540,N_1937,N_1908);
nand U2541 (N_2541,N_2370,N_1872);
and U2542 (N_2542,N_1877,N_1807);
xnor U2543 (N_2543,N_1831,N_2077);
and U2544 (N_2544,N_2195,N_1854);
nor U2545 (N_2545,N_2376,N_1829);
nor U2546 (N_2546,N_2155,N_2284);
or U2547 (N_2547,N_1861,N_1898);
or U2548 (N_2548,N_2206,N_1832);
or U2549 (N_2549,N_2337,N_1809);
nor U2550 (N_2550,N_2007,N_2290);
nand U2551 (N_2551,N_1982,N_1837);
or U2552 (N_2552,N_2091,N_2019);
nor U2553 (N_2553,N_2359,N_1974);
or U2554 (N_2554,N_2283,N_2324);
nand U2555 (N_2555,N_2010,N_2172);
xnor U2556 (N_2556,N_2031,N_2250);
and U2557 (N_2557,N_2298,N_2072);
nand U2558 (N_2558,N_1960,N_2003);
or U2559 (N_2559,N_2012,N_1909);
nor U2560 (N_2560,N_2261,N_2351);
and U2561 (N_2561,N_2215,N_2048);
nor U2562 (N_2562,N_2016,N_2392);
nand U2563 (N_2563,N_2287,N_2073);
nor U2564 (N_2564,N_2229,N_2076);
nor U2565 (N_2565,N_2253,N_1946);
nor U2566 (N_2566,N_2186,N_1943);
and U2567 (N_2567,N_2101,N_1962);
xnor U2568 (N_2568,N_2187,N_2279);
xnor U2569 (N_2569,N_2100,N_2098);
nand U2570 (N_2570,N_2201,N_2034);
nand U2571 (N_2571,N_1989,N_1955);
or U2572 (N_2572,N_2342,N_2271);
and U2573 (N_2573,N_2165,N_1849);
or U2574 (N_2574,N_2081,N_2269);
nand U2575 (N_2575,N_2203,N_1801);
and U2576 (N_2576,N_2347,N_1907);
nor U2577 (N_2577,N_1885,N_1985);
and U2578 (N_2578,N_1900,N_2029);
nor U2579 (N_2579,N_2093,N_2060);
and U2580 (N_2580,N_2220,N_1926);
nand U2581 (N_2581,N_2135,N_1871);
nor U2582 (N_2582,N_2317,N_2040);
nor U2583 (N_2583,N_1927,N_1966);
nor U2584 (N_2584,N_2037,N_1959);
nand U2585 (N_2585,N_2183,N_1925);
and U2586 (N_2586,N_1884,N_1981);
or U2587 (N_2587,N_2385,N_2235);
and U2588 (N_2588,N_2276,N_1949);
nor U2589 (N_2589,N_2295,N_2015);
nor U2590 (N_2590,N_1834,N_2355);
nand U2591 (N_2591,N_1983,N_2334);
nand U2592 (N_2592,N_2202,N_1828);
and U2593 (N_2593,N_2266,N_1967);
xor U2594 (N_2594,N_2116,N_1804);
nor U2595 (N_2595,N_2274,N_2149);
or U2596 (N_2596,N_2260,N_2300);
and U2597 (N_2597,N_1815,N_1822);
nor U2598 (N_2598,N_1843,N_1953);
nand U2599 (N_2599,N_1823,N_2125);
or U2600 (N_2600,N_1964,N_1868);
or U2601 (N_2601,N_2143,N_2282);
nor U2602 (N_2602,N_1929,N_1914);
xor U2603 (N_2603,N_2224,N_1940);
or U2604 (N_2604,N_2368,N_2102);
or U2605 (N_2605,N_1839,N_2014);
and U2606 (N_2606,N_2340,N_2210);
nor U2607 (N_2607,N_2277,N_2327);
nand U2608 (N_2608,N_1968,N_2110);
nand U2609 (N_2609,N_1919,N_2156);
and U2610 (N_2610,N_2111,N_2190);
nor U2611 (N_2611,N_2107,N_2248);
and U2612 (N_2612,N_2057,N_2189);
nand U2613 (N_2613,N_2154,N_2318);
or U2614 (N_2614,N_2177,N_2371);
and U2615 (N_2615,N_1935,N_2167);
or U2616 (N_2616,N_1911,N_1899);
and U2617 (N_2617,N_1846,N_1931);
and U2618 (N_2618,N_2362,N_2150);
nand U2619 (N_2619,N_2170,N_2305);
xor U2620 (N_2620,N_2294,N_1947);
nand U2621 (N_2621,N_2174,N_2079);
and U2622 (N_2622,N_1852,N_2349);
xor U2623 (N_2623,N_2262,N_2227);
nand U2624 (N_2624,N_1896,N_1965);
or U2625 (N_2625,N_1859,N_2336);
nand U2626 (N_2626,N_1952,N_2134);
and U2627 (N_2627,N_2364,N_2179);
or U2628 (N_2628,N_1821,N_1921);
or U2629 (N_2629,N_2228,N_2121);
and U2630 (N_2630,N_1816,N_2344);
or U2631 (N_2631,N_2211,N_2128);
nor U2632 (N_2632,N_1973,N_2366);
or U2633 (N_2633,N_1813,N_2200);
nor U2634 (N_2634,N_2234,N_2075);
nor U2635 (N_2635,N_2204,N_2218);
or U2636 (N_2636,N_1826,N_2380);
and U2637 (N_2637,N_2233,N_2301);
nand U2638 (N_2638,N_1917,N_2286);
nor U2639 (N_2639,N_2140,N_2114);
and U2640 (N_2640,N_1904,N_2180);
or U2641 (N_2641,N_1835,N_2000);
and U2642 (N_2642,N_2330,N_1883);
nand U2643 (N_2643,N_2069,N_1905);
nand U2644 (N_2644,N_2078,N_2232);
or U2645 (N_2645,N_1995,N_2054);
and U2646 (N_2646,N_2089,N_2113);
and U2647 (N_2647,N_2030,N_2258);
nor U2648 (N_2648,N_2087,N_2045);
nand U2649 (N_2649,N_2221,N_1811);
xor U2650 (N_2650,N_2365,N_1886);
xnor U2651 (N_2651,N_2181,N_2213);
nand U2652 (N_2652,N_2086,N_2367);
or U2653 (N_2653,N_1990,N_1956);
and U2654 (N_2654,N_2147,N_1897);
nor U2655 (N_2655,N_2379,N_2381);
or U2656 (N_2656,N_1845,N_1997);
or U2657 (N_2657,N_2070,N_2002);
nor U2658 (N_2658,N_2032,N_2272);
xnor U2659 (N_2659,N_1933,N_2219);
and U2660 (N_2660,N_2285,N_1993);
and U2661 (N_2661,N_1820,N_1994);
or U2662 (N_2662,N_2212,N_2246);
and U2663 (N_2663,N_1938,N_2137);
xor U2664 (N_2664,N_2158,N_1838);
nand U2665 (N_2665,N_2389,N_2146);
or U2666 (N_2666,N_2178,N_2061);
and U2667 (N_2667,N_1840,N_2357);
or U2668 (N_2668,N_1825,N_2067);
nand U2669 (N_2669,N_2104,N_2133);
and U2670 (N_2670,N_2005,N_2333);
and U2671 (N_2671,N_2322,N_1916);
nand U2672 (N_2672,N_1864,N_2230);
or U2673 (N_2673,N_2255,N_2242);
nor U2674 (N_2674,N_2096,N_2027);
nor U2675 (N_2675,N_2391,N_1878);
and U2676 (N_2676,N_2397,N_2316);
nand U2677 (N_2677,N_1892,N_2123);
or U2678 (N_2678,N_1894,N_2267);
xnor U2679 (N_2679,N_2009,N_2021);
nand U2680 (N_2680,N_2095,N_2240);
nor U2681 (N_2681,N_1930,N_2280);
or U2682 (N_2682,N_1869,N_2192);
nor U2683 (N_2683,N_1841,N_2315);
xnor U2684 (N_2684,N_2080,N_1882);
or U2685 (N_2685,N_2160,N_2236);
nor U2686 (N_2686,N_2390,N_2185);
or U2687 (N_2687,N_2278,N_2191);
and U2688 (N_2688,N_1950,N_2222);
or U2689 (N_2689,N_2184,N_2059);
nand U2690 (N_2690,N_2129,N_2176);
and U2691 (N_2691,N_1970,N_2360);
nor U2692 (N_2692,N_2291,N_2398);
and U2693 (N_2693,N_2356,N_2223);
nand U2694 (N_2694,N_1847,N_1932);
or U2695 (N_2695,N_2225,N_2063);
or U2696 (N_2696,N_1945,N_2145);
and U2697 (N_2697,N_1889,N_2214);
nand U2698 (N_2698,N_1988,N_2161);
nor U2699 (N_2699,N_1910,N_2198);
and U2700 (N_2700,N_1855,N_1912);
xnor U2701 (N_2701,N_2042,N_1972);
or U2702 (N_2702,N_2300,N_1893);
or U2703 (N_2703,N_1801,N_2090);
and U2704 (N_2704,N_1846,N_1869);
nand U2705 (N_2705,N_1964,N_2317);
or U2706 (N_2706,N_1911,N_2196);
or U2707 (N_2707,N_2147,N_2174);
and U2708 (N_2708,N_1952,N_2326);
or U2709 (N_2709,N_2155,N_2139);
and U2710 (N_2710,N_1916,N_2218);
and U2711 (N_2711,N_1927,N_2090);
nand U2712 (N_2712,N_2089,N_2086);
or U2713 (N_2713,N_2078,N_2046);
nand U2714 (N_2714,N_2016,N_2299);
nand U2715 (N_2715,N_2387,N_2158);
nand U2716 (N_2716,N_1990,N_1819);
or U2717 (N_2717,N_1987,N_2003);
xnor U2718 (N_2718,N_1995,N_2244);
nor U2719 (N_2719,N_2162,N_2233);
nand U2720 (N_2720,N_2146,N_2082);
and U2721 (N_2721,N_2014,N_2343);
nand U2722 (N_2722,N_2342,N_1811);
nor U2723 (N_2723,N_2055,N_1999);
nand U2724 (N_2724,N_2142,N_1896);
nand U2725 (N_2725,N_2274,N_2383);
nand U2726 (N_2726,N_2059,N_2265);
or U2727 (N_2727,N_1918,N_2176);
and U2728 (N_2728,N_2120,N_1965);
nand U2729 (N_2729,N_2388,N_1990);
xor U2730 (N_2730,N_2213,N_2152);
nand U2731 (N_2731,N_1888,N_1870);
nor U2732 (N_2732,N_2149,N_2355);
nor U2733 (N_2733,N_1992,N_2373);
and U2734 (N_2734,N_2125,N_2144);
and U2735 (N_2735,N_1904,N_2053);
and U2736 (N_2736,N_1830,N_2076);
or U2737 (N_2737,N_1821,N_1907);
nand U2738 (N_2738,N_1992,N_2061);
xnor U2739 (N_2739,N_1940,N_1893);
xor U2740 (N_2740,N_2336,N_2322);
nand U2741 (N_2741,N_2372,N_1847);
nor U2742 (N_2742,N_2061,N_2327);
xnor U2743 (N_2743,N_1869,N_2205);
nand U2744 (N_2744,N_2229,N_1905);
and U2745 (N_2745,N_2077,N_1924);
nor U2746 (N_2746,N_2202,N_1961);
xor U2747 (N_2747,N_1825,N_1913);
nand U2748 (N_2748,N_2035,N_1853);
nand U2749 (N_2749,N_1823,N_2013);
nor U2750 (N_2750,N_2134,N_1856);
xnor U2751 (N_2751,N_2057,N_2256);
or U2752 (N_2752,N_2121,N_1928);
nor U2753 (N_2753,N_1962,N_2246);
xor U2754 (N_2754,N_1854,N_2223);
and U2755 (N_2755,N_1960,N_2390);
nor U2756 (N_2756,N_2328,N_2108);
or U2757 (N_2757,N_2225,N_2106);
nor U2758 (N_2758,N_1872,N_2138);
or U2759 (N_2759,N_2315,N_2394);
or U2760 (N_2760,N_2209,N_2396);
xnor U2761 (N_2761,N_1956,N_1911);
nor U2762 (N_2762,N_1894,N_1843);
and U2763 (N_2763,N_2043,N_2178);
xor U2764 (N_2764,N_1851,N_2268);
or U2765 (N_2765,N_2105,N_2377);
or U2766 (N_2766,N_1938,N_2233);
nor U2767 (N_2767,N_2347,N_2171);
nand U2768 (N_2768,N_2071,N_1808);
nor U2769 (N_2769,N_2018,N_2227);
and U2770 (N_2770,N_2114,N_1868);
nor U2771 (N_2771,N_2222,N_1986);
nand U2772 (N_2772,N_2195,N_2031);
and U2773 (N_2773,N_2323,N_2029);
nor U2774 (N_2774,N_1972,N_2348);
and U2775 (N_2775,N_1915,N_1981);
and U2776 (N_2776,N_2152,N_2358);
or U2777 (N_2777,N_2372,N_2347);
nor U2778 (N_2778,N_2210,N_2141);
and U2779 (N_2779,N_2201,N_1919);
or U2780 (N_2780,N_2105,N_2309);
or U2781 (N_2781,N_2336,N_2180);
or U2782 (N_2782,N_2155,N_1880);
nand U2783 (N_2783,N_1980,N_2368);
and U2784 (N_2784,N_2104,N_1804);
and U2785 (N_2785,N_2024,N_1867);
and U2786 (N_2786,N_2221,N_2254);
nand U2787 (N_2787,N_2188,N_1932);
or U2788 (N_2788,N_1872,N_1881);
and U2789 (N_2789,N_2344,N_2212);
or U2790 (N_2790,N_2306,N_1863);
xnor U2791 (N_2791,N_2235,N_1883);
and U2792 (N_2792,N_1854,N_1971);
nor U2793 (N_2793,N_2056,N_2005);
or U2794 (N_2794,N_1879,N_1991);
and U2795 (N_2795,N_1879,N_2100);
xnor U2796 (N_2796,N_1993,N_1851);
nor U2797 (N_2797,N_1879,N_1935);
nand U2798 (N_2798,N_1960,N_1873);
or U2799 (N_2799,N_2081,N_2115);
and U2800 (N_2800,N_1856,N_2074);
or U2801 (N_2801,N_2172,N_2142);
nor U2802 (N_2802,N_2212,N_1937);
or U2803 (N_2803,N_2093,N_1933);
nand U2804 (N_2804,N_1877,N_1869);
or U2805 (N_2805,N_2191,N_1875);
nor U2806 (N_2806,N_2179,N_2074);
or U2807 (N_2807,N_2278,N_2322);
nor U2808 (N_2808,N_2154,N_2103);
nand U2809 (N_2809,N_1917,N_2151);
nand U2810 (N_2810,N_2215,N_2105);
xnor U2811 (N_2811,N_2319,N_1961);
nor U2812 (N_2812,N_2281,N_2010);
and U2813 (N_2813,N_1900,N_1871);
nand U2814 (N_2814,N_2154,N_1975);
nor U2815 (N_2815,N_2096,N_2393);
and U2816 (N_2816,N_1808,N_1959);
nor U2817 (N_2817,N_1927,N_2081);
xor U2818 (N_2818,N_2094,N_1981);
nand U2819 (N_2819,N_2324,N_2332);
xor U2820 (N_2820,N_2343,N_2008);
xnor U2821 (N_2821,N_1815,N_2196);
nand U2822 (N_2822,N_2028,N_1873);
and U2823 (N_2823,N_2081,N_2239);
nand U2824 (N_2824,N_1954,N_2222);
or U2825 (N_2825,N_2174,N_2378);
nand U2826 (N_2826,N_2153,N_2046);
nand U2827 (N_2827,N_2226,N_2092);
nor U2828 (N_2828,N_1991,N_2200);
or U2829 (N_2829,N_1955,N_1971);
nand U2830 (N_2830,N_1981,N_2335);
or U2831 (N_2831,N_2281,N_1930);
or U2832 (N_2832,N_2043,N_2088);
nand U2833 (N_2833,N_2050,N_2081);
nand U2834 (N_2834,N_2333,N_2360);
nand U2835 (N_2835,N_2354,N_2384);
or U2836 (N_2836,N_2015,N_2264);
or U2837 (N_2837,N_2043,N_2041);
or U2838 (N_2838,N_1902,N_1934);
nor U2839 (N_2839,N_2115,N_1908);
or U2840 (N_2840,N_2065,N_2398);
nor U2841 (N_2841,N_2386,N_2377);
nor U2842 (N_2842,N_2328,N_2162);
and U2843 (N_2843,N_2124,N_2054);
or U2844 (N_2844,N_2082,N_2285);
or U2845 (N_2845,N_2142,N_1814);
nor U2846 (N_2846,N_2158,N_2366);
or U2847 (N_2847,N_1866,N_2361);
xor U2848 (N_2848,N_1873,N_1888);
nand U2849 (N_2849,N_2364,N_1898);
or U2850 (N_2850,N_2365,N_2047);
nor U2851 (N_2851,N_2351,N_2318);
and U2852 (N_2852,N_2176,N_2339);
or U2853 (N_2853,N_1877,N_1885);
nand U2854 (N_2854,N_2292,N_2009);
and U2855 (N_2855,N_2328,N_1866);
or U2856 (N_2856,N_2222,N_1917);
nand U2857 (N_2857,N_1934,N_2163);
nor U2858 (N_2858,N_1865,N_2347);
xnor U2859 (N_2859,N_2261,N_2335);
nor U2860 (N_2860,N_2316,N_1829);
and U2861 (N_2861,N_1915,N_1828);
or U2862 (N_2862,N_2124,N_2301);
or U2863 (N_2863,N_1831,N_2004);
or U2864 (N_2864,N_2198,N_1967);
and U2865 (N_2865,N_2103,N_1926);
xnor U2866 (N_2866,N_1894,N_2231);
or U2867 (N_2867,N_2365,N_2364);
nor U2868 (N_2868,N_2193,N_1838);
nor U2869 (N_2869,N_1823,N_1983);
or U2870 (N_2870,N_2327,N_2117);
nand U2871 (N_2871,N_2326,N_2027);
nand U2872 (N_2872,N_1933,N_1960);
xor U2873 (N_2873,N_2004,N_1806);
nor U2874 (N_2874,N_2222,N_2282);
nor U2875 (N_2875,N_2359,N_2270);
xnor U2876 (N_2876,N_2052,N_2337);
or U2877 (N_2877,N_1854,N_1833);
nor U2878 (N_2878,N_2156,N_1934);
nand U2879 (N_2879,N_2348,N_2069);
or U2880 (N_2880,N_1915,N_2169);
xnor U2881 (N_2881,N_1813,N_2234);
xor U2882 (N_2882,N_2095,N_1898);
nor U2883 (N_2883,N_2388,N_2239);
nor U2884 (N_2884,N_2219,N_2225);
xnor U2885 (N_2885,N_2128,N_2258);
and U2886 (N_2886,N_2224,N_2090);
and U2887 (N_2887,N_2105,N_2175);
or U2888 (N_2888,N_2190,N_2218);
or U2889 (N_2889,N_2196,N_1872);
or U2890 (N_2890,N_2096,N_2299);
nand U2891 (N_2891,N_1953,N_2124);
nand U2892 (N_2892,N_2173,N_1924);
and U2893 (N_2893,N_2365,N_2301);
nor U2894 (N_2894,N_2204,N_2285);
nand U2895 (N_2895,N_2203,N_2366);
and U2896 (N_2896,N_2158,N_1941);
or U2897 (N_2897,N_1947,N_1917);
or U2898 (N_2898,N_2230,N_2293);
and U2899 (N_2899,N_1935,N_1884);
or U2900 (N_2900,N_1868,N_1899);
nor U2901 (N_2901,N_2274,N_1972);
nand U2902 (N_2902,N_2065,N_2136);
and U2903 (N_2903,N_2179,N_2082);
xor U2904 (N_2904,N_2248,N_2005);
and U2905 (N_2905,N_1948,N_2324);
xor U2906 (N_2906,N_2006,N_1874);
and U2907 (N_2907,N_1901,N_1942);
nand U2908 (N_2908,N_2036,N_2366);
and U2909 (N_2909,N_2319,N_1850);
nand U2910 (N_2910,N_1801,N_2291);
and U2911 (N_2911,N_2347,N_2014);
nand U2912 (N_2912,N_2164,N_2266);
or U2913 (N_2913,N_2262,N_2068);
xor U2914 (N_2914,N_1868,N_1906);
xor U2915 (N_2915,N_2364,N_1938);
nor U2916 (N_2916,N_1969,N_2074);
nor U2917 (N_2917,N_1825,N_2097);
xnor U2918 (N_2918,N_1940,N_2269);
nor U2919 (N_2919,N_2194,N_2101);
nand U2920 (N_2920,N_1969,N_2350);
nand U2921 (N_2921,N_2024,N_2156);
nand U2922 (N_2922,N_1951,N_2396);
xor U2923 (N_2923,N_1822,N_2318);
nor U2924 (N_2924,N_1853,N_2191);
or U2925 (N_2925,N_1888,N_2093);
or U2926 (N_2926,N_2015,N_1841);
and U2927 (N_2927,N_1918,N_2136);
nor U2928 (N_2928,N_2383,N_2077);
nor U2929 (N_2929,N_2028,N_2029);
and U2930 (N_2930,N_2071,N_2068);
and U2931 (N_2931,N_1894,N_2118);
nand U2932 (N_2932,N_1913,N_1920);
xnor U2933 (N_2933,N_2293,N_2332);
and U2934 (N_2934,N_2252,N_2294);
nor U2935 (N_2935,N_1829,N_1879);
nor U2936 (N_2936,N_1896,N_2158);
nand U2937 (N_2937,N_1854,N_1899);
and U2938 (N_2938,N_2380,N_2222);
nand U2939 (N_2939,N_1926,N_2280);
nand U2940 (N_2940,N_2246,N_1928);
and U2941 (N_2941,N_2388,N_2248);
and U2942 (N_2942,N_2104,N_2379);
and U2943 (N_2943,N_2369,N_1836);
nor U2944 (N_2944,N_2364,N_1835);
and U2945 (N_2945,N_1883,N_1982);
nand U2946 (N_2946,N_1903,N_1930);
nand U2947 (N_2947,N_2107,N_1990);
nor U2948 (N_2948,N_2378,N_1877);
nor U2949 (N_2949,N_2081,N_2217);
xor U2950 (N_2950,N_2111,N_2019);
nand U2951 (N_2951,N_1921,N_2096);
or U2952 (N_2952,N_2219,N_2349);
nand U2953 (N_2953,N_2266,N_2235);
nor U2954 (N_2954,N_2210,N_1915);
nor U2955 (N_2955,N_1986,N_2255);
nand U2956 (N_2956,N_1927,N_1843);
nand U2957 (N_2957,N_2191,N_2222);
nor U2958 (N_2958,N_2358,N_2253);
nor U2959 (N_2959,N_1955,N_2237);
and U2960 (N_2960,N_2131,N_2090);
nand U2961 (N_2961,N_2079,N_2265);
nand U2962 (N_2962,N_1996,N_2283);
and U2963 (N_2963,N_2098,N_2027);
and U2964 (N_2964,N_2036,N_2343);
xor U2965 (N_2965,N_1874,N_2111);
or U2966 (N_2966,N_1965,N_2145);
and U2967 (N_2967,N_2353,N_2236);
and U2968 (N_2968,N_1978,N_2297);
nor U2969 (N_2969,N_2323,N_2192);
and U2970 (N_2970,N_1949,N_1940);
and U2971 (N_2971,N_1945,N_1924);
xnor U2972 (N_2972,N_2240,N_2062);
nand U2973 (N_2973,N_2300,N_2083);
or U2974 (N_2974,N_2288,N_2340);
or U2975 (N_2975,N_2184,N_1939);
nor U2976 (N_2976,N_2182,N_2013);
xor U2977 (N_2977,N_2156,N_2060);
or U2978 (N_2978,N_1834,N_2305);
and U2979 (N_2979,N_2189,N_2324);
nor U2980 (N_2980,N_2000,N_2037);
or U2981 (N_2981,N_2114,N_1984);
nand U2982 (N_2982,N_2351,N_2109);
nand U2983 (N_2983,N_2228,N_2320);
nand U2984 (N_2984,N_2300,N_2333);
nand U2985 (N_2985,N_2242,N_2149);
or U2986 (N_2986,N_2276,N_2155);
or U2987 (N_2987,N_2145,N_1838);
or U2988 (N_2988,N_1935,N_2124);
nand U2989 (N_2989,N_2383,N_1875);
or U2990 (N_2990,N_2186,N_2203);
nor U2991 (N_2991,N_2193,N_2268);
nor U2992 (N_2992,N_2181,N_1854);
nor U2993 (N_2993,N_2139,N_1961);
or U2994 (N_2994,N_1834,N_2145);
and U2995 (N_2995,N_2089,N_2345);
or U2996 (N_2996,N_2261,N_2304);
or U2997 (N_2997,N_2060,N_1956);
and U2998 (N_2998,N_2306,N_2181);
xor U2999 (N_2999,N_2389,N_2209);
or UO_0 (O_0,N_2554,N_2752);
nand UO_1 (O_1,N_2601,N_2960);
or UO_2 (O_2,N_2481,N_2871);
or UO_3 (O_3,N_2518,N_2701);
nor UO_4 (O_4,N_2876,N_2593);
nand UO_5 (O_5,N_2462,N_2666);
nand UO_6 (O_6,N_2607,N_2543);
or UO_7 (O_7,N_2504,N_2927);
xnor UO_8 (O_8,N_2972,N_2477);
nor UO_9 (O_9,N_2842,N_2401);
xor UO_10 (O_10,N_2633,N_2721);
or UO_11 (O_11,N_2716,N_2758);
nor UO_12 (O_12,N_2637,N_2777);
or UO_13 (O_13,N_2761,N_2947);
or UO_14 (O_14,N_2614,N_2864);
xnor UO_15 (O_15,N_2743,N_2813);
nand UO_16 (O_16,N_2650,N_2836);
nor UO_17 (O_17,N_2403,N_2667);
nand UO_18 (O_18,N_2430,N_2949);
and UO_19 (O_19,N_2652,N_2923);
or UO_20 (O_20,N_2509,N_2683);
xnor UO_21 (O_21,N_2555,N_2682);
nand UO_22 (O_22,N_2793,N_2442);
or UO_23 (O_23,N_2575,N_2796);
nand UO_24 (O_24,N_2912,N_2724);
or UO_25 (O_25,N_2981,N_2723);
nor UO_26 (O_26,N_2645,N_2706);
nand UO_27 (O_27,N_2914,N_2558);
nor UO_28 (O_28,N_2431,N_2839);
or UO_29 (O_29,N_2475,N_2474);
nand UO_30 (O_30,N_2859,N_2885);
xor UO_31 (O_31,N_2797,N_2426);
or UO_32 (O_32,N_2454,N_2898);
nor UO_33 (O_33,N_2992,N_2974);
or UO_34 (O_34,N_2853,N_2616);
or UO_35 (O_35,N_2816,N_2953);
nand UO_36 (O_36,N_2862,N_2841);
nand UO_37 (O_37,N_2966,N_2515);
or UO_38 (O_38,N_2734,N_2902);
and UO_39 (O_39,N_2468,N_2817);
nor UO_40 (O_40,N_2609,N_2773);
nor UO_41 (O_41,N_2844,N_2566);
nand UO_42 (O_42,N_2651,N_2411);
nand UO_43 (O_43,N_2643,N_2684);
or UO_44 (O_44,N_2450,N_2417);
nand UO_45 (O_45,N_2603,N_2646);
and UO_46 (O_46,N_2897,N_2492);
and UO_47 (O_47,N_2409,N_2443);
and UO_48 (O_48,N_2828,N_2423);
or UO_49 (O_49,N_2771,N_2672);
and UO_50 (O_50,N_2869,N_2644);
nor UO_51 (O_51,N_2521,N_2970);
or UO_52 (O_52,N_2449,N_2808);
xor UO_53 (O_53,N_2501,N_2825);
or UO_54 (O_54,N_2438,N_2608);
and UO_55 (O_55,N_2563,N_2597);
nand UO_56 (O_56,N_2913,N_2460);
nand UO_57 (O_57,N_2617,N_2400);
or UO_58 (O_58,N_2804,N_2961);
nand UO_59 (O_59,N_2976,N_2964);
and UO_60 (O_60,N_2582,N_2886);
or UO_61 (O_61,N_2675,N_2639);
nand UO_62 (O_62,N_2707,N_2412);
xnor UO_63 (O_63,N_2704,N_2795);
xor UO_64 (O_64,N_2835,N_2562);
nor UO_65 (O_65,N_2516,N_2933);
nor UO_66 (O_66,N_2592,N_2879);
and UO_67 (O_67,N_2638,N_2679);
and UO_68 (O_68,N_2792,N_2730);
or UO_69 (O_69,N_2491,N_2801);
nor UO_70 (O_70,N_2720,N_2840);
nor UO_71 (O_71,N_2917,N_2785);
nand UO_72 (O_72,N_2975,N_2747);
or UO_73 (O_73,N_2647,N_2901);
or UO_74 (O_74,N_2494,N_2725);
nand UO_75 (O_75,N_2402,N_2738);
or UO_76 (O_76,N_2938,N_2416);
or UO_77 (O_77,N_2779,N_2822);
or UO_78 (O_78,N_2532,N_2506);
or UO_79 (O_79,N_2658,N_2447);
nand UO_80 (O_80,N_2588,N_2998);
nor UO_81 (O_81,N_2990,N_2894);
or UO_82 (O_82,N_2482,N_2620);
nor UO_83 (O_83,N_2728,N_2478);
or UO_84 (O_84,N_2594,N_2868);
or UO_85 (O_85,N_2674,N_2470);
and UO_86 (O_86,N_2753,N_2539);
xnor UO_87 (O_87,N_2687,N_2425);
and UO_88 (O_88,N_2663,N_2678);
and UO_89 (O_89,N_2484,N_2732);
xor UO_90 (O_90,N_2595,N_2439);
and UO_91 (O_91,N_2709,N_2433);
and UO_92 (O_92,N_2993,N_2987);
and UO_93 (O_93,N_2583,N_2548);
or UO_94 (O_94,N_2819,N_2769);
nor UO_95 (O_95,N_2692,N_2541);
xor UO_96 (O_96,N_2965,N_2551);
and UO_97 (O_97,N_2994,N_2668);
and UO_98 (O_98,N_2524,N_2549);
xor UO_99 (O_99,N_2452,N_2754);
and UO_100 (O_100,N_2415,N_2591);
nor UO_101 (O_101,N_2778,N_2843);
nor UO_102 (O_102,N_2556,N_2560);
or UO_103 (O_103,N_2969,N_2948);
nand UO_104 (O_104,N_2649,N_2744);
or UO_105 (O_105,N_2787,N_2500);
and UO_106 (O_106,N_2559,N_2435);
nand UO_107 (O_107,N_2580,N_2736);
nand UO_108 (O_108,N_2523,N_2669);
nand UO_109 (O_109,N_2453,N_2446);
and UO_110 (O_110,N_2479,N_2802);
or UO_111 (O_111,N_2847,N_2877);
nor UO_112 (O_112,N_2892,N_2888);
nand UO_113 (O_113,N_2550,N_2906);
or UO_114 (O_114,N_2708,N_2613);
or UO_115 (O_115,N_2745,N_2655);
nor UO_116 (O_116,N_2640,N_2852);
or UO_117 (O_117,N_2810,N_2887);
or UO_118 (O_118,N_2576,N_2574);
or UO_119 (O_119,N_2611,N_2820);
nand UO_120 (O_120,N_2542,N_2939);
and UO_121 (O_121,N_2823,N_2967);
nand UO_122 (O_122,N_2472,N_2765);
nand UO_123 (O_123,N_2424,N_2693);
nand UO_124 (O_124,N_2940,N_2610);
and UO_125 (O_125,N_2526,N_2767);
xnor UO_126 (O_126,N_2891,N_2552);
or UO_127 (O_127,N_2459,N_2729);
nand UO_128 (O_128,N_2890,N_2971);
and UO_129 (O_129,N_2671,N_2905);
or UO_130 (O_130,N_2731,N_2627);
nor UO_131 (O_131,N_2700,N_2957);
or UO_132 (O_132,N_2865,N_2636);
xor UO_133 (O_133,N_2641,N_2600);
xnor UO_134 (O_134,N_2855,N_2741);
nor UO_135 (O_135,N_2619,N_2826);
nor UO_136 (O_136,N_2444,N_2958);
and UO_137 (O_137,N_2455,N_2800);
nor UO_138 (O_138,N_2733,N_2831);
nand UO_139 (O_139,N_2705,N_2697);
nor UO_140 (O_140,N_2489,N_2480);
and UO_141 (O_141,N_2875,N_2832);
and UO_142 (O_142,N_2829,N_2686);
and UO_143 (O_143,N_2654,N_2851);
nor UO_144 (O_144,N_2952,N_2624);
xor UO_145 (O_145,N_2936,N_2937);
nand UO_146 (O_146,N_2712,N_2578);
or UO_147 (O_147,N_2568,N_2846);
and UO_148 (O_148,N_2904,N_2473);
and UO_149 (O_149,N_2856,N_2653);
nand UO_150 (O_150,N_2916,N_2534);
xor UO_151 (O_151,N_2996,N_2634);
xnor UO_152 (O_152,N_2485,N_2821);
and UO_153 (O_153,N_2907,N_2751);
nor UO_154 (O_154,N_2943,N_2922);
and UO_155 (O_155,N_2935,N_2861);
and UO_156 (O_156,N_2457,N_2919);
and UO_157 (O_157,N_2874,N_2579);
nand UO_158 (O_158,N_2628,N_2467);
nor UO_159 (O_159,N_2408,N_2698);
and UO_160 (O_160,N_2978,N_2929);
or UO_161 (O_161,N_2980,N_2977);
and UO_162 (O_162,N_2565,N_2547);
nor UO_163 (O_163,N_2776,N_2755);
and UO_164 (O_164,N_2714,N_2512);
and UO_165 (O_165,N_2955,N_2717);
or UO_166 (O_166,N_2989,N_2737);
nor UO_167 (O_167,N_2456,N_2858);
or UO_168 (O_168,N_2997,N_2931);
and UO_169 (O_169,N_2661,N_2872);
nand UO_170 (O_170,N_2882,N_2571);
and UO_171 (O_171,N_2428,N_2814);
xor UO_172 (O_172,N_2849,N_2405);
and UO_173 (O_173,N_2713,N_2437);
nor UO_174 (O_174,N_2794,N_2418);
and UO_175 (O_175,N_2807,N_2941);
nor UO_176 (O_176,N_2445,N_2854);
or UO_177 (O_177,N_2806,N_2419);
xnor UO_178 (O_178,N_2893,N_2680);
nand UO_179 (O_179,N_2632,N_2768);
nand UO_180 (O_180,N_2538,N_2621);
and UO_181 (O_181,N_2496,N_2791);
and UO_182 (O_182,N_2528,N_2903);
or UO_183 (O_183,N_2809,N_2530);
nor UO_184 (O_184,N_2766,N_2458);
nand UO_185 (O_185,N_2896,N_2803);
nand UO_186 (O_186,N_2488,N_2770);
nand UO_187 (O_187,N_2746,N_2845);
nor UO_188 (O_188,N_2799,N_2606);
and UO_189 (O_189,N_2464,N_2735);
and UO_190 (O_190,N_2763,N_2889);
nor UO_191 (O_191,N_2781,N_2909);
nor UO_192 (O_192,N_2469,N_2944);
or UO_193 (O_193,N_2465,N_2866);
nor UO_194 (O_194,N_2503,N_2699);
and UO_195 (O_195,N_2911,N_2900);
nor UO_196 (O_196,N_2883,N_2422);
xnor UO_197 (O_197,N_2589,N_2432);
and UO_198 (O_198,N_2921,N_2522);
and UO_199 (O_199,N_2584,N_2722);
nand UO_200 (O_200,N_2507,N_2838);
nand UO_201 (O_201,N_2696,N_2880);
or UO_202 (O_202,N_2662,N_2577);
nor UO_203 (O_203,N_2536,N_2727);
nand UO_204 (O_204,N_2915,N_2635);
xor UO_205 (O_205,N_2694,N_2519);
or UO_206 (O_206,N_2510,N_2740);
xor UO_207 (O_207,N_2573,N_2749);
nor UO_208 (O_208,N_2487,N_2585);
nor UO_209 (O_209,N_2895,N_2695);
and UO_210 (O_210,N_2673,N_2483);
nor UO_211 (O_211,N_2812,N_2567);
and UO_212 (O_212,N_2517,N_2780);
and UO_213 (O_213,N_2999,N_2789);
xor UO_214 (O_214,N_2715,N_2815);
or UO_215 (O_215,N_2991,N_2691);
or UO_216 (O_216,N_2448,N_2626);
or UO_217 (O_217,N_2604,N_2703);
nor UO_218 (O_218,N_2920,N_2490);
and UO_219 (O_219,N_2925,N_2407);
or UO_220 (O_220,N_2625,N_2973);
and UO_221 (O_221,N_2757,N_2502);
nor UO_222 (O_222,N_2954,N_2878);
nand UO_223 (O_223,N_2870,N_2984);
nand UO_224 (O_224,N_2615,N_2742);
or UO_225 (O_225,N_2544,N_2605);
xor UO_226 (O_226,N_2748,N_2834);
and UO_227 (O_227,N_2531,N_2629);
nor UO_228 (O_228,N_2739,N_2557);
or UO_229 (O_229,N_2928,N_2656);
and UO_230 (O_230,N_2962,N_2786);
nand UO_231 (O_231,N_2756,N_2463);
nand UO_232 (O_232,N_2587,N_2527);
and UO_233 (O_233,N_2676,N_2711);
nand UO_234 (O_234,N_2612,N_2908);
nor UO_235 (O_235,N_2790,N_2561);
nand UO_236 (O_236,N_2857,N_2677);
and UO_237 (O_237,N_2622,N_2505);
nor UO_238 (O_238,N_2884,N_2598);
nand UO_239 (O_239,N_2436,N_2586);
nand UO_240 (O_240,N_2410,N_2899);
or UO_241 (O_241,N_2618,N_2783);
nor UO_242 (O_242,N_2529,N_2533);
nand UO_243 (O_243,N_2486,N_2760);
and UO_244 (O_244,N_2985,N_2867);
nand UO_245 (O_245,N_2945,N_2833);
and UO_246 (O_246,N_2873,N_2553);
and UO_247 (O_247,N_2414,N_2498);
and UO_248 (O_248,N_2772,N_2762);
nor UO_249 (O_249,N_2540,N_2461);
and UO_250 (O_250,N_2811,N_2514);
and UO_251 (O_251,N_2429,N_2986);
nor UO_252 (O_252,N_2599,N_2421);
or UO_253 (O_253,N_2968,N_2982);
nor UO_254 (O_254,N_2545,N_2427);
or UO_255 (O_255,N_2631,N_2784);
xor UO_256 (O_256,N_2910,N_2942);
or UO_257 (O_257,N_2495,N_2520);
or UO_258 (O_258,N_2493,N_2926);
or UO_259 (O_259,N_2710,N_2659);
nor UO_260 (O_260,N_2818,N_2569);
and UO_261 (O_261,N_2688,N_2535);
nor UO_262 (O_262,N_2983,N_2979);
xnor UO_263 (O_263,N_2660,N_2956);
or UO_264 (O_264,N_2963,N_2642);
nor UO_265 (O_265,N_2782,N_2497);
nand UO_266 (O_266,N_2657,N_2932);
nand UO_267 (O_267,N_2950,N_2476);
or UO_268 (O_268,N_2681,N_2434);
nor UO_269 (O_269,N_2924,N_2988);
or UO_270 (O_270,N_2471,N_2726);
or UO_271 (O_271,N_2805,N_2525);
and UO_272 (O_272,N_2863,N_2959);
or UO_273 (O_273,N_2406,N_2596);
or UO_274 (O_274,N_2404,N_2798);
nand UO_275 (O_275,N_2918,N_2764);
or UO_276 (O_276,N_2788,N_2934);
and UO_277 (O_277,N_2750,N_2420);
or UO_278 (O_278,N_2830,N_2827);
nor UO_279 (O_279,N_2689,N_2513);
nand UO_280 (O_280,N_2511,N_2581);
nand UO_281 (O_281,N_2824,N_2690);
nor UO_282 (O_282,N_2718,N_2499);
and UO_283 (O_283,N_2665,N_2441);
and UO_284 (O_284,N_2451,N_2572);
or UO_285 (O_285,N_2951,N_2570);
xor UO_286 (O_286,N_2546,N_2466);
nand UO_287 (O_287,N_2440,N_2670);
and UO_288 (O_288,N_2623,N_2702);
nor UO_289 (O_289,N_2564,N_2685);
and UO_290 (O_290,N_2848,N_2537);
nor UO_291 (O_291,N_2850,N_2664);
nand UO_292 (O_292,N_2837,N_2759);
nand UO_293 (O_293,N_2719,N_2774);
nor UO_294 (O_294,N_2946,N_2602);
nand UO_295 (O_295,N_2860,N_2413);
nand UO_296 (O_296,N_2881,N_2775);
and UO_297 (O_297,N_2590,N_2630);
xor UO_298 (O_298,N_2648,N_2508);
nor UO_299 (O_299,N_2995,N_2930);
nand UO_300 (O_300,N_2585,N_2788);
nor UO_301 (O_301,N_2674,N_2695);
and UO_302 (O_302,N_2785,N_2765);
nand UO_303 (O_303,N_2622,N_2798);
nor UO_304 (O_304,N_2824,N_2736);
nor UO_305 (O_305,N_2854,N_2916);
and UO_306 (O_306,N_2502,N_2534);
and UO_307 (O_307,N_2490,N_2758);
nand UO_308 (O_308,N_2491,N_2966);
nand UO_309 (O_309,N_2808,N_2436);
or UO_310 (O_310,N_2411,N_2735);
nor UO_311 (O_311,N_2655,N_2698);
nand UO_312 (O_312,N_2767,N_2602);
nor UO_313 (O_313,N_2755,N_2632);
nor UO_314 (O_314,N_2692,N_2420);
nand UO_315 (O_315,N_2979,N_2959);
or UO_316 (O_316,N_2563,N_2575);
nor UO_317 (O_317,N_2844,N_2528);
nand UO_318 (O_318,N_2775,N_2827);
and UO_319 (O_319,N_2750,N_2856);
and UO_320 (O_320,N_2575,N_2808);
nor UO_321 (O_321,N_2972,N_2471);
nor UO_322 (O_322,N_2419,N_2496);
nand UO_323 (O_323,N_2872,N_2551);
or UO_324 (O_324,N_2518,N_2529);
nand UO_325 (O_325,N_2470,N_2896);
nor UO_326 (O_326,N_2981,N_2760);
nand UO_327 (O_327,N_2505,N_2727);
nand UO_328 (O_328,N_2566,N_2690);
nor UO_329 (O_329,N_2886,N_2894);
or UO_330 (O_330,N_2584,N_2527);
and UO_331 (O_331,N_2466,N_2419);
and UO_332 (O_332,N_2937,N_2541);
or UO_333 (O_333,N_2744,N_2557);
nor UO_334 (O_334,N_2932,N_2960);
nor UO_335 (O_335,N_2843,N_2471);
and UO_336 (O_336,N_2408,N_2771);
nand UO_337 (O_337,N_2539,N_2853);
nor UO_338 (O_338,N_2530,N_2513);
nor UO_339 (O_339,N_2816,N_2631);
nor UO_340 (O_340,N_2964,N_2795);
nor UO_341 (O_341,N_2809,N_2862);
or UO_342 (O_342,N_2784,N_2825);
and UO_343 (O_343,N_2862,N_2993);
nand UO_344 (O_344,N_2405,N_2838);
nor UO_345 (O_345,N_2406,N_2513);
nor UO_346 (O_346,N_2966,N_2992);
and UO_347 (O_347,N_2831,N_2460);
nand UO_348 (O_348,N_2459,N_2968);
nand UO_349 (O_349,N_2807,N_2838);
nor UO_350 (O_350,N_2747,N_2605);
or UO_351 (O_351,N_2424,N_2426);
or UO_352 (O_352,N_2448,N_2890);
nor UO_353 (O_353,N_2430,N_2893);
nand UO_354 (O_354,N_2827,N_2925);
nand UO_355 (O_355,N_2679,N_2894);
nand UO_356 (O_356,N_2856,N_2578);
xnor UO_357 (O_357,N_2432,N_2893);
and UO_358 (O_358,N_2606,N_2741);
nand UO_359 (O_359,N_2561,N_2588);
or UO_360 (O_360,N_2807,N_2619);
nor UO_361 (O_361,N_2477,N_2870);
or UO_362 (O_362,N_2567,N_2876);
or UO_363 (O_363,N_2999,N_2448);
nor UO_364 (O_364,N_2615,N_2689);
xor UO_365 (O_365,N_2788,N_2860);
or UO_366 (O_366,N_2530,N_2847);
and UO_367 (O_367,N_2590,N_2915);
nor UO_368 (O_368,N_2781,N_2485);
nor UO_369 (O_369,N_2719,N_2499);
or UO_370 (O_370,N_2905,N_2836);
or UO_371 (O_371,N_2566,N_2966);
or UO_372 (O_372,N_2922,N_2438);
nand UO_373 (O_373,N_2950,N_2623);
or UO_374 (O_374,N_2602,N_2628);
and UO_375 (O_375,N_2657,N_2794);
or UO_376 (O_376,N_2604,N_2690);
nor UO_377 (O_377,N_2682,N_2775);
and UO_378 (O_378,N_2521,N_2814);
nand UO_379 (O_379,N_2897,N_2536);
or UO_380 (O_380,N_2890,N_2616);
and UO_381 (O_381,N_2864,N_2868);
and UO_382 (O_382,N_2512,N_2944);
or UO_383 (O_383,N_2731,N_2718);
nor UO_384 (O_384,N_2820,N_2405);
or UO_385 (O_385,N_2642,N_2411);
nand UO_386 (O_386,N_2612,N_2501);
and UO_387 (O_387,N_2417,N_2999);
nor UO_388 (O_388,N_2471,N_2974);
and UO_389 (O_389,N_2723,N_2507);
nor UO_390 (O_390,N_2519,N_2904);
or UO_391 (O_391,N_2929,N_2844);
or UO_392 (O_392,N_2578,N_2483);
and UO_393 (O_393,N_2606,N_2492);
nor UO_394 (O_394,N_2717,N_2449);
or UO_395 (O_395,N_2606,N_2625);
nand UO_396 (O_396,N_2444,N_2474);
nor UO_397 (O_397,N_2535,N_2625);
and UO_398 (O_398,N_2728,N_2629);
xnor UO_399 (O_399,N_2456,N_2895);
and UO_400 (O_400,N_2656,N_2688);
nor UO_401 (O_401,N_2642,N_2973);
or UO_402 (O_402,N_2473,N_2982);
xor UO_403 (O_403,N_2523,N_2979);
or UO_404 (O_404,N_2709,N_2492);
xnor UO_405 (O_405,N_2928,N_2899);
nand UO_406 (O_406,N_2761,N_2502);
nand UO_407 (O_407,N_2870,N_2428);
or UO_408 (O_408,N_2686,N_2903);
nand UO_409 (O_409,N_2654,N_2969);
or UO_410 (O_410,N_2945,N_2442);
nand UO_411 (O_411,N_2489,N_2964);
nand UO_412 (O_412,N_2402,N_2866);
or UO_413 (O_413,N_2693,N_2856);
or UO_414 (O_414,N_2434,N_2991);
nor UO_415 (O_415,N_2605,N_2523);
xnor UO_416 (O_416,N_2680,N_2728);
xor UO_417 (O_417,N_2580,N_2598);
xnor UO_418 (O_418,N_2692,N_2865);
nor UO_419 (O_419,N_2735,N_2801);
or UO_420 (O_420,N_2879,N_2817);
and UO_421 (O_421,N_2754,N_2918);
or UO_422 (O_422,N_2924,N_2503);
xnor UO_423 (O_423,N_2727,N_2833);
or UO_424 (O_424,N_2803,N_2403);
nor UO_425 (O_425,N_2745,N_2581);
or UO_426 (O_426,N_2666,N_2628);
nor UO_427 (O_427,N_2509,N_2561);
nand UO_428 (O_428,N_2975,N_2646);
nor UO_429 (O_429,N_2858,N_2433);
nand UO_430 (O_430,N_2621,N_2923);
and UO_431 (O_431,N_2488,N_2422);
or UO_432 (O_432,N_2902,N_2430);
nand UO_433 (O_433,N_2709,N_2569);
nand UO_434 (O_434,N_2762,N_2699);
and UO_435 (O_435,N_2960,N_2954);
xnor UO_436 (O_436,N_2754,N_2464);
nand UO_437 (O_437,N_2415,N_2620);
and UO_438 (O_438,N_2794,N_2690);
nor UO_439 (O_439,N_2701,N_2495);
and UO_440 (O_440,N_2945,N_2814);
nand UO_441 (O_441,N_2788,N_2540);
xnor UO_442 (O_442,N_2538,N_2531);
nand UO_443 (O_443,N_2850,N_2548);
and UO_444 (O_444,N_2982,N_2616);
xnor UO_445 (O_445,N_2545,N_2893);
nand UO_446 (O_446,N_2786,N_2532);
or UO_447 (O_447,N_2533,N_2972);
xor UO_448 (O_448,N_2413,N_2538);
and UO_449 (O_449,N_2647,N_2993);
and UO_450 (O_450,N_2673,N_2533);
xor UO_451 (O_451,N_2802,N_2672);
or UO_452 (O_452,N_2540,N_2586);
xor UO_453 (O_453,N_2949,N_2603);
or UO_454 (O_454,N_2528,N_2887);
or UO_455 (O_455,N_2684,N_2627);
nor UO_456 (O_456,N_2954,N_2962);
and UO_457 (O_457,N_2553,N_2710);
or UO_458 (O_458,N_2456,N_2867);
xor UO_459 (O_459,N_2934,N_2705);
nor UO_460 (O_460,N_2774,N_2715);
nor UO_461 (O_461,N_2595,N_2627);
xnor UO_462 (O_462,N_2820,N_2986);
or UO_463 (O_463,N_2424,N_2957);
xor UO_464 (O_464,N_2511,N_2586);
nor UO_465 (O_465,N_2409,N_2991);
nor UO_466 (O_466,N_2726,N_2780);
and UO_467 (O_467,N_2462,N_2910);
or UO_468 (O_468,N_2510,N_2788);
nand UO_469 (O_469,N_2869,N_2960);
nand UO_470 (O_470,N_2655,N_2564);
nor UO_471 (O_471,N_2473,N_2582);
nand UO_472 (O_472,N_2912,N_2596);
nand UO_473 (O_473,N_2612,N_2492);
nand UO_474 (O_474,N_2807,N_2401);
nor UO_475 (O_475,N_2677,N_2631);
nand UO_476 (O_476,N_2974,N_2692);
nand UO_477 (O_477,N_2613,N_2792);
or UO_478 (O_478,N_2791,N_2604);
or UO_479 (O_479,N_2765,N_2873);
and UO_480 (O_480,N_2915,N_2997);
nand UO_481 (O_481,N_2628,N_2649);
nor UO_482 (O_482,N_2525,N_2890);
nand UO_483 (O_483,N_2735,N_2899);
and UO_484 (O_484,N_2902,N_2487);
nor UO_485 (O_485,N_2756,N_2952);
or UO_486 (O_486,N_2454,N_2810);
xnor UO_487 (O_487,N_2429,N_2881);
nor UO_488 (O_488,N_2821,N_2441);
xor UO_489 (O_489,N_2919,N_2672);
or UO_490 (O_490,N_2837,N_2926);
and UO_491 (O_491,N_2481,N_2873);
nand UO_492 (O_492,N_2824,N_2767);
or UO_493 (O_493,N_2560,N_2594);
nand UO_494 (O_494,N_2434,N_2534);
nor UO_495 (O_495,N_2991,N_2587);
or UO_496 (O_496,N_2516,N_2639);
and UO_497 (O_497,N_2805,N_2887);
nor UO_498 (O_498,N_2659,N_2409);
nand UO_499 (O_499,N_2521,N_2767);
endmodule