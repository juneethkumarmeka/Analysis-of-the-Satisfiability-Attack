module basic_3000_30000_3500_30_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_1928,In_1389);
nor U1 (N_1,In_1712,In_2753);
nand U2 (N_2,In_147,In_2859);
nor U3 (N_3,In_1784,In_1022);
nand U4 (N_4,In_1974,In_1726);
and U5 (N_5,In_2435,In_2697);
nand U6 (N_6,In_2870,In_396);
xor U7 (N_7,In_1522,In_523);
nand U8 (N_8,In_637,In_1417);
xor U9 (N_9,In_1869,In_2706);
nor U10 (N_10,In_839,In_2772);
xor U11 (N_11,In_179,In_691);
nor U12 (N_12,In_1880,In_1879);
nand U13 (N_13,In_267,In_2200);
xnor U14 (N_14,In_229,In_1893);
nand U15 (N_15,In_2548,In_1478);
or U16 (N_16,In_657,In_2925);
nand U17 (N_17,In_2114,In_2675);
nand U18 (N_18,In_1746,In_675);
nand U19 (N_19,In_269,In_1727);
and U20 (N_20,In_1519,In_1118);
and U21 (N_21,In_1601,In_1094);
nand U22 (N_22,In_2113,In_613);
nor U23 (N_23,In_601,In_444);
nor U24 (N_24,In_1590,In_912);
nor U25 (N_25,In_2845,In_1937);
nand U26 (N_26,In_1265,In_292);
nand U27 (N_27,In_706,In_832);
and U28 (N_28,In_2996,In_166);
or U29 (N_29,In_1402,In_1212);
xor U30 (N_30,In_2771,In_2539);
nand U31 (N_31,In_2705,In_632);
nand U32 (N_32,In_1592,In_735);
and U33 (N_33,In_988,In_299);
nor U34 (N_34,In_2401,In_2755);
nand U35 (N_35,In_1907,In_2045);
and U36 (N_36,In_2551,In_1385);
xor U37 (N_37,In_294,In_1273);
and U38 (N_38,In_2614,In_97);
or U39 (N_39,In_870,In_608);
xor U40 (N_40,In_2083,In_1698);
nand U41 (N_41,In_1939,In_289);
or U42 (N_42,In_1906,In_2838);
nor U43 (N_43,In_101,In_1454);
or U44 (N_44,In_1431,In_971);
nor U45 (N_45,In_1160,In_76);
or U46 (N_46,In_1918,In_1462);
or U47 (N_47,In_33,In_1322);
and U48 (N_48,In_1081,In_1681);
xnor U49 (N_49,In_1806,In_469);
or U50 (N_50,In_1466,In_1200);
nand U51 (N_51,In_1667,In_1315);
nor U52 (N_52,In_2280,In_2546);
nor U53 (N_53,In_1850,In_1499);
and U54 (N_54,In_2948,In_2277);
nand U55 (N_55,In_1832,In_2159);
xor U56 (N_56,In_2799,In_983);
nand U57 (N_57,In_771,In_2222);
or U58 (N_58,In_1734,In_1624);
xnor U59 (N_59,In_1891,In_216);
or U60 (N_60,In_712,In_1899);
or U61 (N_61,In_2575,In_2933);
or U62 (N_62,In_886,In_1044);
xnor U63 (N_63,In_961,In_1023);
nand U64 (N_64,In_11,In_2853);
nor U65 (N_65,In_2648,In_2993);
xor U66 (N_66,In_2020,In_2698);
or U67 (N_67,In_1070,In_1803);
nand U68 (N_68,In_81,In_2062);
nand U69 (N_69,In_29,In_681);
and U70 (N_70,In_1621,In_2515);
or U71 (N_71,In_848,In_1333);
and U72 (N_72,In_2734,In_2152);
xnor U73 (N_73,In_1556,In_1193);
nand U74 (N_74,In_2740,In_2470);
nand U75 (N_75,In_1532,In_2544);
and U76 (N_76,In_1537,In_30);
or U77 (N_77,In_2489,In_1905);
or U78 (N_78,In_2269,In_916);
nand U79 (N_79,In_2408,In_2966);
nor U80 (N_80,In_2228,In_346);
and U81 (N_81,In_2503,In_270);
or U82 (N_82,In_1946,In_1763);
and U83 (N_83,In_2813,In_734);
nand U84 (N_84,In_2709,In_160);
xor U85 (N_85,In_2794,In_1515);
or U86 (N_86,In_1640,In_2754);
and U87 (N_87,In_1046,In_2527);
nor U88 (N_88,In_555,In_1836);
nor U89 (N_89,In_2224,In_298);
nand U90 (N_90,In_2823,In_2673);
nand U91 (N_91,In_2008,In_2878);
nand U92 (N_92,In_312,In_2442);
nand U93 (N_93,In_416,In_1236);
xnor U94 (N_94,In_2054,In_2260);
nor U95 (N_95,In_742,In_2191);
and U96 (N_96,In_622,In_2559);
or U97 (N_97,In_1514,In_1352);
xnor U98 (N_98,In_471,In_598);
and U99 (N_99,In_2497,In_1630);
xnor U100 (N_100,In_1096,In_1429);
and U101 (N_101,In_1145,In_1544);
or U102 (N_102,In_1168,In_2148);
and U103 (N_103,In_755,In_2074);
and U104 (N_104,In_1473,In_2684);
xor U105 (N_105,In_110,In_909);
nand U106 (N_106,In_2413,In_2216);
nor U107 (N_107,In_2218,In_2031);
or U108 (N_108,In_628,In_656);
xnor U109 (N_109,In_689,In_562);
and U110 (N_110,In_2815,In_1877);
xor U111 (N_111,In_1314,In_2821);
nor U112 (N_112,In_922,In_2163);
nand U113 (N_113,In_1910,In_1816);
nand U114 (N_114,In_2596,In_667);
or U115 (N_115,In_1740,In_286);
or U116 (N_116,In_1670,In_2690);
nor U117 (N_117,In_1165,In_2025);
nand U118 (N_118,In_1255,In_715);
and U119 (N_119,In_2321,In_680);
or U120 (N_120,In_705,In_1393);
nor U121 (N_121,In_1881,In_700);
or U122 (N_122,In_1520,In_898);
nand U123 (N_123,In_1357,In_368);
xnor U124 (N_124,In_731,In_2909);
or U125 (N_125,In_478,In_957);
nand U126 (N_126,In_307,In_2582);
nor U127 (N_127,In_1468,In_1778);
nand U128 (N_128,In_1759,In_2434);
xor U129 (N_129,In_170,In_259);
and U130 (N_130,In_1350,In_84);
xor U131 (N_131,In_795,In_1755);
xor U132 (N_132,In_150,In_1310);
nor U133 (N_133,In_498,In_1767);
xnor U134 (N_134,In_2292,In_729);
xor U135 (N_135,In_173,In_1896);
nand U136 (N_136,In_685,In_1396);
xor U137 (N_137,In_1497,In_204);
xor U138 (N_138,In_1810,In_218);
xnor U139 (N_139,In_906,In_1364);
nand U140 (N_140,In_2383,In_2997);
xor U141 (N_141,In_1737,In_967);
nand U142 (N_142,In_1823,In_387);
nand U143 (N_143,In_2586,In_2495);
nand U144 (N_144,In_865,In_2855);
or U145 (N_145,In_573,In_1476);
and U146 (N_146,In_2556,In_2492);
nor U147 (N_147,In_2632,In_1442);
and U148 (N_148,In_1686,In_2379);
nor U149 (N_149,In_2214,In_2454);
and U150 (N_150,In_1410,In_1109);
xnor U151 (N_151,In_1294,In_353);
and U152 (N_152,In_2381,In_1078);
xor U153 (N_153,In_2276,In_920);
xor U154 (N_154,In_1733,In_2649);
or U155 (N_155,In_2249,In_2553);
xor U156 (N_156,In_1653,In_2959);
or U157 (N_157,In_2373,In_139);
and U158 (N_158,In_2954,In_558);
or U159 (N_159,In_2728,In_1471);
or U160 (N_160,In_747,In_381);
or U161 (N_161,In_180,In_445);
nor U162 (N_162,In_169,In_516);
nor U163 (N_163,In_798,In_1099);
xnor U164 (N_164,In_1090,In_794);
nand U165 (N_165,In_1676,In_648);
and U166 (N_166,In_435,In_694);
xor U167 (N_167,In_15,In_1969);
and U168 (N_168,In_2477,In_2095);
nand U169 (N_169,In_1422,In_0);
and U170 (N_170,In_1451,In_1925);
nand U171 (N_171,In_948,In_805);
nor U172 (N_172,In_1485,In_2980);
nand U173 (N_173,In_441,In_1239);
nor U174 (N_174,In_278,In_2721);
and U175 (N_175,In_1401,In_778);
or U176 (N_176,In_1040,In_708);
or U177 (N_177,In_65,In_1275);
and U178 (N_178,In_1517,In_2037);
or U179 (N_179,In_1944,In_2097);
and U180 (N_180,In_1056,In_385);
xnor U181 (N_181,In_2160,In_897);
nor U182 (N_182,In_371,In_1369);
nand U183 (N_183,In_2991,In_674);
and U184 (N_184,In_2407,In_111);
or U185 (N_185,In_2053,In_1004);
xnor U186 (N_186,In_1817,In_2136);
or U187 (N_187,In_393,In_2830);
nand U188 (N_188,In_2471,In_591);
nor U189 (N_189,In_2911,In_2938);
xnor U190 (N_190,In_2915,In_18);
nand U191 (N_191,In_1249,In_2463);
or U192 (N_192,In_374,In_842);
xnor U193 (N_193,In_1089,In_2776);
and U194 (N_194,In_2024,In_2588);
nor U195 (N_195,In_382,In_44);
nand U196 (N_196,In_1756,In_2978);
nor U197 (N_197,In_2341,In_2513);
xnor U198 (N_198,In_1814,In_1366);
or U199 (N_199,In_513,In_1516);
and U200 (N_200,In_1989,In_530);
or U201 (N_201,In_1133,In_2343);
nand U202 (N_202,In_9,In_2841);
nor U203 (N_203,In_1735,In_1710);
nor U204 (N_204,In_2060,In_2182);
and U205 (N_205,In_847,In_887);
xor U206 (N_206,In_1865,In_2668);
xnor U207 (N_207,In_2928,In_236);
xor U208 (N_208,In_793,In_1958);
nor U209 (N_209,In_1167,In_2485);
and U210 (N_210,In_237,In_360);
and U211 (N_211,In_1150,In_1194);
and U212 (N_212,In_1186,In_1487);
nor U213 (N_213,In_1392,In_2888);
nor U214 (N_214,In_2439,In_981);
or U215 (N_215,In_176,In_2038);
nand U216 (N_216,In_1453,In_1403);
and U217 (N_217,In_1649,In_2009);
or U218 (N_218,In_1020,In_846);
and U219 (N_219,In_2512,In_2749);
and U220 (N_220,In_1277,In_1845);
xnor U221 (N_221,In_1687,In_873);
nand U222 (N_222,In_224,In_2036);
nor U223 (N_223,In_941,In_272);
or U224 (N_224,In_2233,In_1965);
and U225 (N_225,In_1264,In_138);
nor U226 (N_226,In_436,In_2012);
xor U227 (N_227,In_1480,In_1587);
xnor U228 (N_228,In_459,In_2945);
nor U229 (N_229,In_2500,In_2761);
nand U230 (N_230,In_1950,In_1388);
nand U231 (N_231,In_1339,In_2677);
and U232 (N_232,In_2158,In_2636);
and U233 (N_233,In_1619,In_2579);
nor U234 (N_234,In_868,In_740);
or U235 (N_235,In_2969,In_363);
nand U236 (N_236,In_1146,In_1885);
nand U237 (N_237,In_1302,In_320);
or U238 (N_238,In_2727,In_902);
nand U239 (N_239,In_300,In_658);
or U240 (N_240,In_820,In_2412);
nand U241 (N_241,In_973,In_2899);
and U242 (N_242,In_593,In_1927);
nor U243 (N_243,In_2150,In_1419);
nor U244 (N_244,In_1503,In_2511);
and U245 (N_245,In_2528,In_668);
nor U246 (N_246,In_748,In_1585);
and U247 (N_247,In_537,In_944);
and U248 (N_248,In_2703,In_1890);
or U249 (N_249,In_2849,In_2328);
and U250 (N_250,In_905,In_2004);
and U251 (N_251,In_2059,In_2644);
and U252 (N_252,In_1943,In_305);
xor U253 (N_253,In_2699,In_2447);
and U254 (N_254,In_1644,In_2229);
nor U255 (N_255,In_806,In_2764);
xor U256 (N_256,In_1844,In_27);
nand U257 (N_257,In_2109,In_2493);
nand U258 (N_258,In_2883,In_409);
nor U259 (N_259,In_521,In_894);
xor U260 (N_260,In_1783,In_189);
and U261 (N_261,In_2898,In_2866);
xor U262 (N_262,In_1536,In_2161);
xor U263 (N_263,In_1608,In_1359);
nor U264 (N_264,In_670,In_2977);
nand U265 (N_265,In_750,In_2115);
or U266 (N_266,In_164,In_2048);
xnor U267 (N_267,In_1643,In_2580);
xnor U268 (N_268,In_1715,In_661);
xor U269 (N_269,In_824,In_2284);
nand U270 (N_270,In_2084,In_2430);
nor U271 (N_271,In_1589,In_2777);
nand U272 (N_272,In_1830,In_1084);
or U273 (N_273,In_1948,In_2930);
nor U274 (N_274,In_2758,In_117);
and U275 (N_275,In_2645,In_1208);
and U276 (N_276,In_238,In_114);
nand U277 (N_277,In_2605,In_1219);
xor U278 (N_278,In_2624,In_1280);
and U279 (N_279,In_1033,In_154);
nor U280 (N_280,In_654,In_1903);
nor U281 (N_281,In_1680,In_344);
xor U282 (N_282,In_1597,In_2459);
xnor U283 (N_283,In_1460,In_816);
or U284 (N_284,In_1518,In_407);
xnor U285 (N_285,In_1378,In_2329);
or U286 (N_286,In_2861,In_94);
or U287 (N_287,In_2934,In_2076);
or U288 (N_288,In_2968,In_502);
or U289 (N_289,In_541,In_2018);
nor U290 (N_290,In_2530,In_858);
and U291 (N_291,In_762,In_1005);
or U292 (N_292,In_251,In_2236);
or U293 (N_293,In_1338,In_349);
nand U294 (N_294,In_1661,In_2552);
and U295 (N_295,In_1873,In_2810);
and U296 (N_296,In_804,In_1964);
xnor U297 (N_297,In_1771,In_786);
xor U298 (N_298,In_2765,In_413);
and U299 (N_299,In_2804,In_1180);
nand U300 (N_300,In_1859,In_789);
and U301 (N_301,In_2143,In_1308);
or U302 (N_302,In_1149,In_1440);
or U303 (N_303,In_1444,In_2643);
and U304 (N_304,In_2127,In_2850);
xor U305 (N_305,In_143,In_2940);
nor U306 (N_306,In_1483,In_2710);
nand U307 (N_307,In_2431,In_1898);
nor U308 (N_308,In_1702,In_1951);
nor U309 (N_309,In_1260,In_1355);
xor U310 (N_310,In_1911,In_2067);
nand U311 (N_311,In_408,In_2380);
nand U312 (N_312,In_2891,In_188);
and U313 (N_313,In_1148,In_756);
nand U314 (N_314,In_1037,In_2390);
nand U315 (N_315,In_1615,In_2808);
or U316 (N_316,In_664,In_895);
and U317 (N_317,In_1252,In_1954);
xnor U318 (N_318,In_337,In_2029);
or U319 (N_319,In_2211,In_1818);
nand U320 (N_320,In_2679,In_1623);
nand U321 (N_321,In_2340,In_1691);
and U322 (N_322,In_2391,In_2723);
nand U323 (N_323,In_341,In_851);
and U324 (N_324,In_2812,In_2147);
xnor U325 (N_325,In_2735,In_1933);
nand U326 (N_326,In_1409,In_361);
nor U327 (N_327,In_161,In_2188);
and U328 (N_328,In_2906,In_1174);
and U329 (N_329,In_1128,In_547);
nor U330 (N_330,In_61,In_1210);
and U331 (N_331,In_1230,In_1805);
or U332 (N_332,In_775,In_596);
nand U333 (N_333,In_1305,In_669);
nand U334 (N_334,In_1365,In_2014);
and U335 (N_335,In_1085,In_666);
or U336 (N_336,In_1543,In_2212);
or U337 (N_337,In_1871,In_1293);
and U338 (N_338,In_2678,In_862);
nor U339 (N_339,In_2345,In_1656);
nand U340 (N_340,In_168,In_380);
and U341 (N_341,In_711,In_1018);
and U342 (N_342,In_1711,In_2350);
nand U343 (N_343,In_2016,In_106);
nand U344 (N_344,In_1479,In_2369);
nand U345 (N_345,In_1028,In_651);
nand U346 (N_346,In_19,In_1639);
nand U347 (N_347,In_12,In_1706);
xnor U348 (N_348,In_1721,In_334);
nor U349 (N_349,In_1450,In_508);
nand U350 (N_350,In_1434,In_2429);
and U351 (N_351,In_2642,In_1408);
and U352 (N_352,In_1674,In_2295);
nor U353 (N_353,In_607,In_2784);
xnor U354 (N_354,In_2738,In_1062);
or U355 (N_355,In_979,In_1102);
nand U356 (N_356,In_1611,In_487);
and U357 (N_357,In_2332,In_2173);
nand U358 (N_358,In_940,In_751);
and U359 (N_359,In_2300,In_2897);
xor U360 (N_360,In_1047,In_2985);
or U361 (N_361,In_2935,In_2221);
xnor U362 (N_362,In_2288,In_2577);
nand U363 (N_363,In_659,In_455);
and U364 (N_364,In_2490,In_1919);
xor U365 (N_365,In_1929,In_399);
xor U366 (N_366,In_1709,In_829);
xnor U367 (N_367,In_877,In_1183);
nand U368 (N_368,In_171,In_2676);
xor U369 (N_369,In_788,In_575);
or U370 (N_370,In_51,In_2090);
or U371 (N_371,In_69,In_2842);
and U372 (N_372,In_2460,In_871);
nand U373 (N_373,In_2438,In_317);
nor U374 (N_374,In_896,In_2183);
nor U375 (N_375,In_1579,In_1184);
nor U376 (N_376,In_301,In_1704);
nor U377 (N_377,In_780,In_1741);
or U378 (N_378,In_2879,In_1425);
nand U379 (N_379,In_115,In_539);
nand U380 (N_380,In_2205,In_1596);
and U381 (N_381,In_71,In_821);
or U382 (N_382,In_774,In_818);
nand U383 (N_383,In_463,In_205);
nand U384 (N_384,In_500,In_2733);
xnor U385 (N_385,In_1482,In_1016);
and U386 (N_386,In_2998,In_1934);
nand U387 (N_387,In_1531,In_1187);
nand U388 (N_388,In_1296,In_1481);
nand U389 (N_389,In_1664,In_2901);
and U390 (N_390,In_1942,In_1988);
and U391 (N_391,In_828,In_2405);
nor U392 (N_392,In_384,In_1106);
or U393 (N_393,In_1423,In_1141);
nand U394 (N_394,In_1622,In_642);
and U395 (N_395,In_2184,In_2333);
or U396 (N_396,In_2603,In_2667);
nand U397 (N_397,In_50,In_1742);
nor U398 (N_398,In_1012,In_2287);
xnor U399 (N_399,In_733,In_2086);
and U400 (N_400,In_1576,In_1703);
nor U401 (N_401,In_192,In_133);
and U402 (N_402,In_781,In_2137);
nor U403 (N_403,In_2308,In_2651);
and U404 (N_404,In_1984,In_1257);
xnor U405 (N_405,In_1383,In_2518);
nand U406 (N_406,In_102,In_2296);
xor U407 (N_407,In_1895,In_2078);
and U408 (N_408,In_1017,In_515);
or U409 (N_409,In_2741,In_2949);
nand U410 (N_410,In_1335,In_509);
and U411 (N_411,In_1231,In_693);
nand U412 (N_412,In_835,In_2394);
or U413 (N_413,In_2293,In_2529);
xnor U414 (N_414,In_273,In_440);
xor U415 (N_415,In_876,In_2789);
nor U416 (N_416,In_570,In_692);
nand U417 (N_417,In_1550,In_1566);
xnor U418 (N_418,In_2232,In_2298);
xnor U419 (N_419,In_2852,In_1535);
xor U420 (N_420,In_1572,In_2021);
nor U421 (N_421,In_2525,In_1779);
or U422 (N_422,In_1507,In_1281);
xor U423 (N_423,In_976,In_826);
and U424 (N_424,In_1826,In_2833);
xnor U425 (N_425,In_1731,In_1768);
or U426 (N_426,In_2768,In_2519);
xor U427 (N_427,In_1283,In_458);
nor U428 (N_428,In_2123,In_968);
xor U429 (N_429,In_1361,In_2342);
and U430 (N_430,In_1205,In_1699);
or U431 (N_431,In_2618,In_2669);
xor U432 (N_432,In_1326,In_2387);
nand U433 (N_433,In_1061,In_182);
xnor U434 (N_434,In_1999,In_38);
xnor U435 (N_435,In_1523,In_1125);
nor U436 (N_436,In_264,In_125);
nand U437 (N_437,In_2689,In_1775);
or U438 (N_438,In_2757,In_2905);
xor U439 (N_439,In_1801,In_1912);
and U440 (N_440,In_1351,In_370);
xor U441 (N_441,In_1430,In_2375);
nand U442 (N_442,In_1065,In_880);
or U443 (N_443,In_915,In_2167);
or U444 (N_444,In_293,In_1631);
or U445 (N_445,In_1508,In_2358);
or U446 (N_446,In_800,In_910);
or U447 (N_447,In_2658,In_1245);
and U448 (N_448,In_2103,In_1651);
or U449 (N_449,In_429,In_1059);
xor U450 (N_450,In_2615,In_181);
xnor U451 (N_451,In_724,In_243);
or U452 (N_452,In_844,In_2550);
and U453 (N_453,In_1011,In_439);
and U454 (N_454,In_79,In_1841);
nor U455 (N_455,In_2655,In_1051);
and U456 (N_456,In_2461,In_145);
xnor U457 (N_457,In_1334,In_567);
and U458 (N_458,In_2844,In_2540);
nand U459 (N_459,In_25,In_1714);
nor U460 (N_460,In_773,In_1324);
nand U461 (N_461,In_1557,In_2268);
or U462 (N_462,In_524,In_1435);
nand U463 (N_463,In_85,In_1015);
xor U464 (N_464,In_1837,In_1399);
nor U465 (N_465,In_536,In_2102);
nor U466 (N_466,In_1853,In_612);
nand U467 (N_467,In_1446,In_1511);
or U468 (N_468,In_1781,In_2234);
nor U469 (N_469,In_714,In_1506);
nor U470 (N_470,In_1021,In_113);
xnor U471 (N_471,In_1716,In_221);
nor U472 (N_472,In_605,In_2976);
and U473 (N_473,In_2876,In_1578);
xor U474 (N_474,In_903,In_260);
nor U475 (N_475,In_1732,In_813);
nor U476 (N_476,In_2252,In_2947);
or U477 (N_477,In_219,In_1135);
and U478 (N_478,In_2984,In_1382);
and U479 (N_479,In_2502,In_2595);
and U480 (N_480,In_1538,In_451);
and U481 (N_481,In_577,In_974);
and U482 (N_482,In_99,In_1421);
or U483 (N_483,In_290,In_1122);
nor U484 (N_484,In_2424,In_2116);
nor U485 (N_485,In_1376,In_768);
and U486 (N_486,In_52,In_579);
xnor U487 (N_487,In_1874,In_253);
xnor U488 (N_488,In_1496,In_1975);
nand U489 (N_489,In_891,In_2376);
and U490 (N_490,In_2432,In_723);
nand U491 (N_491,In_1226,In_1337);
nand U492 (N_492,In_1632,In_228);
and U493 (N_493,In_1120,In_2964);
xor U494 (N_494,In_1488,In_2426);
and U495 (N_495,In_364,In_2975);
or U496 (N_496,In_2465,In_982);
nor U497 (N_497,In_411,In_1744);
or U498 (N_498,In_2543,In_2065);
nand U499 (N_499,In_1838,In_54);
xnor U500 (N_500,In_13,In_355);
or U501 (N_501,In_45,In_1139);
or U502 (N_502,In_1307,In_564);
xnor U503 (N_503,In_2171,In_199);
nand U504 (N_504,In_635,In_178);
xnor U505 (N_505,In_1683,In_1562);
or U506 (N_506,In_1527,In_306);
or U507 (N_507,In_304,In_2960);
nand U508 (N_508,In_1981,In_2681);
or U509 (N_509,In_945,In_242);
nand U510 (N_510,In_2271,In_2104);
nand U511 (N_511,In_986,In_2175);
nor U512 (N_512,In_1107,In_630);
xor U513 (N_513,In_1822,In_797);
or U514 (N_514,In_1029,In_322);
nand U515 (N_515,In_354,In_1492);
nor U516 (N_516,In_1034,In_2043);
nand U517 (N_517,In_2745,In_2265);
or U518 (N_518,In_474,In_769);
and U519 (N_519,In_86,In_2524);
xnor U520 (N_520,In_1595,In_2731);
and U521 (N_521,In_566,In_2774);
nor U522 (N_522,In_2297,In_662);
and U523 (N_523,In_2592,In_2272);
nand U524 (N_524,In_2918,In_427);
and U525 (N_525,In_701,In_1941);
or U526 (N_526,In_1445,In_2357);
or U527 (N_527,In_8,In_1560);
nor U528 (N_528,In_972,In_2653);
nor U529 (N_529,In_2027,In_2763);
nand U530 (N_530,In_100,In_1030);
nor U531 (N_531,In_2132,In_2722);
nor U532 (N_532,In_1955,In_683);
xor U533 (N_533,In_2769,In_1427);
and U534 (N_534,In_1261,In_953);
or U535 (N_535,In_1297,In_586);
xnor U536 (N_536,In_2294,In_1987);
xor U537 (N_537,In_1164,In_2058);
and U538 (N_538,In_2965,In_2022);
xnor U539 (N_539,In_1512,In_2052);
xor U540 (N_540,In_2818,In_1143);
xor U541 (N_541,In_2261,In_1609);
or U542 (N_542,In_597,In_2953);
xor U543 (N_543,In_1833,In_131);
xnor U544 (N_544,In_250,In_790);
nor U545 (N_545,In_23,In_514);
nand U546 (N_546,In_2363,In_2663);
and U547 (N_547,In_2323,In_336);
and U548 (N_548,In_914,In_72);
nor U549 (N_549,In_191,In_830);
or U550 (N_550,In_324,In_1433);
xor U551 (N_551,In_2927,In_433);
xor U552 (N_552,In_2895,In_141);
or U553 (N_553,In_1795,In_869);
xor U554 (N_554,In_1884,In_87);
or U555 (N_555,In_1749,In_2640);
or U556 (N_556,In_1846,In_2943);
and U557 (N_557,In_2617,In_2779);
and U558 (N_558,In_2318,In_766);
xnor U559 (N_559,In_687,In_907);
nand U560 (N_560,In_966,In_1238);
nor U561 (N_561,In_375,In_1642);
xnor U562 (N_562,In_1209,In_1980);
and U563 (N_563,In_167,In_2542);
nor U564 (N_564,In_739,In_2055);
nand U565 (N_565,In_538,In_2428);
nand U566 (N_566,In_1175,In_1072);
and U567 (N_567,In_456,In_1799);
xor U568 (N_568,In_864,In_696);
nand U569 (N_569,In_126,In_1013);
or U570 (N_570,In_208,In_2661);
or U571 (N_571,In_1739,In_1675);
nand U572 (N_572,In_193,In_758);
xnor U573 (N_573,In_2811,In_450);
xor U574 (N_574,In_241,In_2718);
or U575 (N_575,In_1436,In_468);
nor U576 (N_576,In_2220,In_1404);
xor U577 (N_577,In_1138,In_2538);
nor U578 (N_578,In_41,In_1341);
xnor U579 (N_579,In_2006,In_1087);
xnor U580 (N_580,In_2433,In_2079);
nor U581 (N_581,In_1953,In_2063);
and U582 (N_582,In_365,In_2671);
nand U583 (N_583,In_226,In_990);
or U584 (N_584,In_339,In_1747);
nor U585 (N_585,In_351,In_1356);
nand U586 (N_586,In_486,In_1666);
and U587 (N_587,In_1197,In_2581);
nand U588 (N_588,In_883,In_2035);
and U589 (N_589,In_580,In_767);
xnor U590 (N_590,In_17,In_213);
nor U591 (N_591,In_489,In_1729);
and U592 (N_592,In_206,In_1688);
and U593 (N_593,In_2682,In_1224);
nor U594 (N_594,In_2869,In_2759);
nor U595 (N_595,In_2270,In_1130);
nand U596 (N_596,In_939,In_1045);
xor U597 (N_597,In_2564,In_1932);
and U598 (N_598,In_430,In_1633);
and U599 (N_599,In_825,In_2384);
and U600 (N_600,In_2275,In_2646);
xor U601 (N_601,In_1060,In_913);
xor U602 (N_602,In_2886,In_1792);
and U603 (N_603,In_2659,In_1708);
nand U604 (N_604,In_2843,In_342);
nand U605 (N_605,In_245,In_2312);
nor U606 (N_606,In_2414,In_202);
xor U607 (N_607,In_2194,In_484);
nand U608 (N_608,In_678,In_77);
nand U609 (N_609,In_534,In_310);
or U610 (N_610,In_2921,In_2989);
xor U611 (N_611,In_1663,In_1751);
nor U612 (N_612,In_2047,In_1003);
nand U613 (N_613,In_1963,In_285);
nor U614 (N_614,In_688,In_442);
nand U615 (N_615,In_911,In_2880);
nor U616 (N_616,In_2227,In_388);
xor U617 (N_617,In_1002,In_2486);
nand U618 (N_618,In_2956,In_962);
nand U619 (N_619,In_838,In_22);
xor U620 (N_620,In_1104,In_636);
nor U621 (N_621,In_1765,In_493);
or U622 (N_622,In_624,In_931);
or U623 (N_623,In_198,In_2441);
nor U624 (N_624,In_1213,In_1173);
and U625 (N_625,In_2650,In_1713);
xor U626 (N_626,In_390,In_652);
or U627 (N_627,In_889,In_625);
and U628 (N_628,In_960,In_1787);
and U629 (N_629,In_1997,In_2778);
nor U630 (N_630,In_1788,In_2696);
or U631 (N_631,In_908,In_1990);
and U632 (N_632,In_1019,In_1390);
and U633 (N_633,In_1521,In_759);
nor U634 (N_634,In_2190,In_1320);
and U635 (N_635,In_1620,In_2507);
or U636 (N_636,In_1692,In_1961);
nand U637 (N_637,In_1114,In_1221);
nand U638 (N_638,In_2273,In_587);
xnor U639 (N_639,In_1993,In_311);
nand U640 (N_640,In_277,In_819);
xnor U641 (N_641,In_1719,In_918);
nor U642 (N_642,In_1952,In_2170);
nand U643 (N_643,In_1707,In_2120);
or U644 (N_644,In_137,In_1750);
nand U645 (N_645,In_1486,In_1793);
xnor U646 (N_646,In_2361,In_148);
nor U647 (N_647,In_2744,In_2366);
and U648 (N_648,In_671,In_2064);
nand U649 (N_649,In_1284,In_1602);
or U650 (N_650,In_2416,In_2801);
and U651 (N_651,In_1876,In_520);
nand U652 (N_652,In_2071,In_2793);
or U653 (N_653,In_2118,In_2747);
nor U654 (N_654,In_1510,In_2467);
xnor U655 (N_655,In_2290,In_2309);
nor U656 (N_656,In_415,In_2611);
or U657 (N_657,In_857,In_1868);
xor U658 (N_658,In_796,In_2665);
or U659 (N_659,In_418,In_333);
and U660 (N_660,In_746,In_522);
nor U661 (N_661,In_629,In_501);
nand U662 (N_662,In_281,In_643);
and U663 (N_663,In_1368,In_938);
nor U664 (N_664,In_2139,In_2971);
xnor U665 (N_665,In_1857,In_2972);
or U666 (N_666,In_600,In_1725);
nor U667 (N_667,In_2767,In_2574);
and U668 (N_668,In_582,In_2446);
and U669 (N_669,In_546,In_1565);
nand U670 (N_670,In_1705,In_1607);
or U671 (N_671,In_1472,In_1278);
xnor U672 (N_672,In_2834,In_2326);
and U673 (N_673,In_1115,In_96);
nand U674 (N_674,In_999,In_2652);
or U675 (N_675,In_812,In_736);
or U676 (N_676,In_2291,In_975);
nor U677 (N_677,In_952,In_2398);
or U678 (N_678,In_2992,In_1494);
xor U679 (N_679,In_645,In_1465);
xnor U680 (N_680,In_1552,In_2347);
and U681 (N_681,In_2263,In_885);
or U682 (N_682,In_93,In_901);
and U683 (N_683,In_2482,In_207);
and U684 (N_684,In_1971,In_1490);
nor U685 (N_685,In_128,In_1437);
and U686 (N_686,In_836,In_1612);
xnor U687 (N_687,In_2466,In_2803);
and U688 (N_688,In_74,In_62);
xor U689 (N_689,In_1782,In_947);
xor U690 (N_690,In_1336,In_1233);
and U691 (N_691,In_162,In_2286);
nor U692 (N_692,In_1923,In_230);
and U693 (N_693,In_1548,In_1828);
nand U694 (N_694,In_810,In_1154);
xor U695 (N_695,In_67,In_481);
xnor U696 (N_696,In_1088,In_2420);
xor U697 (N_697,In_1617,In_2317);
nand U698 (N_698,In_2715,In_2942);
or U699 (N_699,In_2498,In_1424);
nand U700 (N_700,In_1459,In_2257);
nor U701 (N_701,In_1117,In_2141);
and U702 (N_702,In_2344,In_215);
nor U703 (N_703,In_1772,In_1291);
nand U704 (N_704,In_2231,In_2730);
xor U705 (N_705,In_2410,In_2623);
or U706 (N_706,In_677,In_1181);
xnor U707 (N_707,In_1387,In_2377);
nand U708 (N_708,In_1201,In_56);
nand U709 (N_709,In_104,In_2189);
nand U710 (N_710,In_1770,In_1126);
xor U711 (N_711,In_2448,In_2204);
nor U712 (N_712,In_1225,In_943);
or U713 (N_713,In_2258,In_1227);
and U714 (N_714,In_194,In_438);
or U715 (N_715,In_872,In_2683);
or U716 (N_716,In_831,In_2001);
xnor U717 (N_717,In_1864,In_1812);
and U718 (N_718,In_2070,In_722);
xnor U719 (N_719,In_1461,In_2638);
or U720 (N_720,In_1024,In_282);
and U721 (N_721,In_1840,In_2837);
and U722 (N_722,In_2100,In_1718);
or U723 (N_723,In_2105,In_921);
or U724 (N_724,In_37,In_2664);
nor U725 (N_725,In_2604,In_2185);
nand U726 (N_726,In_1648,In_2637);
nand U727 (N_727,In_764,In_802);
nor U728 (N_728,In_1701,In_1723);
xor U729 (N_729,In_2856,In_2537);
nor U730 (N_730,In_615,In_2283);
nand U731 (N_731,In_550,In_969);
nor U732 (N_732,In_1137,In_1802);
or U733 (N_733,In_1170,In_725);
nor U734 (N_734,In_646,In_470);
or U735 (N_735,In_2816,In_2081);
nand U736 (N_736,In_732,In_2600);
or U737 (N_737,In_1203,In_4);
and U738 (N_738,In_548,In_2421);
nand U739 (N_739,In_2450,In_1584);
and U740 (N_740,In_1829,In_2742);
xor U741 (N_741,In_1196,In_2066);
xnor U742 (N_742,In_995,In_2572);
nand U743 (N_743,In_2151,In_568);
or U744 (N_744,In_1900,In_1358);
nand U745 (N_745,In_201,In_419);
nor U746 (N_746,In_1915,In_996);
nand U747 (N_747,In_2256,In_553);
and U748 (N_748,In_2602,In_2629);
xnor U749 (N_749,In_994,In_1300);
nand U750 (N_750,In_485,In_1696);
or U751 (N_751,In_1689,In_75);
xor U752 (N_752,In_1894,In_2154);
xnor U753 (N_753,In_2462,In_88);
or U754 (N_754,In_1367,In_1972);
nor U755 (N_755,In_403,In_379);
nand U756 (N_756,In_1743,In_2633);
and U757 (N_757,In_1785,In_543);
or U758 (N_758,In_958,In_1534);
xnor U759 (N_759,In_2476,In_315);
nand U760 (N_760,In_297,In_1312);
and U761 (N_761,In_2628,In_2364);
and U762 (N_762,In_2000,In_2126);
and U763 (N_763,In_507,In_1752);
or U764 (N_764,In_697,In_942);
nand U765 (N_765,In_2936,In_690);
nand U766 (N_766,In_2807,In_373);
nor U767 (N_767,In_987,In_531);
xnor U768 (N_768,In_893,In_2451);
nand U769 (N_769,In_2311,In_2262);
or U770 (N_770,In_1259,In_1878);
nand U771 (N_771,In_472,In_223);
and U772 (N_772,In_2202,In_576);
and U773 (N_773,In_142,In_1276);
or U774 (N_774,In_2306,In_2701);
xor U775 (N_775,In_754,In_186);
nor U776 (N_776,In_2389,In_2092);
nand U777 (N_777,In_621,In_2199);
and U778 (N_778,In_1458,In_726);
nand U779 (N_779,In_1240,In_2957);
xnor U780 (N_780,In_153,In_665);
nand U781 (N_781,In_782,In_1524);
and U782 (N_782,In_1774,In_884);
xnor U783 (N_783,In_2877,In_980);
nand U784 (N_784,In_2562,In_497);
nand U785 (N_785,In_1054,In_1068);
or U786 (N_786,In_1204,In_540);
and U787 (N_787,In_432,In_452);
or U788 (N_788,In_1539,In_225);
nand U789 (N_789,In_965,In_1292);
or U790 (N_790,In_476,In_561);
and U791 (N_791,In_1132,In_510);
xnor U792 (N_792,In_1241,In_2187);
or U793 (N_793,In_710,In_1827);
nor U794 (N_794,In_604,In_149);
xnor U795 (N_795,In_412,In_165);
and U796 (N_796,In_1764,In_1025);
nand U797 (N_797,In_1108,In_1362);
and U798 (N_798,In_397,In_2647);
nand U799 (N_799,In_2798,In_332);
xor U800 (N_800,In_888,In_1374);
xor U801 (N_801,In_91,In_2209);
or U802 (N_802,In_2452,In_2907);
nand U803 (N_803,In_410,In_1395);
and U804 (N_804,In_2680,In_2266);
nand U805 (N_805,In_1027,In_1904);
and U806 (N_806,In_1796,In_1131);
nand U807 (N_807,In_35,In_569);
and U808 (N_808,In_2091,In_2080);
or U809 (N_809,In_676,In_1113);
nor U810 (N_810,In_2299,In_1924);
or U811 (N_811,In_1977,In_423);
nor U812 (N_812,In_850,In_1039);
nor U813 (N_813,In_348,In_483);
xnor U814 (N_814,In_2313,In_1558);
or U815 (N_815,In_1574,In_2359);
and U816 (N_816,In_1151,In_2922);
xnor U817 (N_817,In_2931,In_785);
xnor U818 (N_818,In_46,In_1014);
nor U819 (N_819,In_2320,In_2056);
nand U820 (N_820,In_2041,In_1901);
or U821 (N_821,In_1780,In_599);
or U822 (N_822,In_2917,In_1169);
or U823 (N_823,In_713,In_1007);
nor U824 (N_824,In_1962,In_2072);
and U825 (N_825,In_2217,In_2478);
nand U826 (N_826,In_2660,In_118);
and U827 (N_827,In_933,In_2932);
nor U828 (N_828,In_1207,In_1414);
or U829 (N_829,In_602,In_1220);
or U830 (N_830,In_2725,In_14);
and U831 (N_831,In_1573,In_1347);
nand U832 (N_832,In_2285,In_263);
nand U833 (N_833,In_1420,In_1474);
nor U834 (N_834,In_2026,In_1504);
xnor U835 (N_835,In_2890,In_2634);
nor U836 (N_836,In_1346,In_1647);
nor U837 (N_837,In_252,In_2822);
and U838 (N_838,In_801,In_1909);
nor U839 (N_839,In_158,In_2440);
or U840 (N_840,In_2089,In_1311);
and U841 (N_841,In_2444,In_1069);
xor U842 (N_842,In_1156,In_728);
or U843 (N_843,In_2657,In_2003);
or U844 (N_844,In_549,In_827);
and U845 (N_845,In_1509,In_2245);
and U846 (N_846,In_232,In_1247);
nand U847 (N_847,In_1237,In_2590);
nand U848 (N_848,In_776,In_2015);
and U849 (N_849,In_2887,In_2809);
nor U850 (N_850,In_749,In_1134);
nor U851 (N_851,In_1618,In_425);
nor U852 (N_852,In_2472,In_2226);
xnor U853 (N_853,In_2950,In_964);
nand U854 (N_854,In_2613,In_2112);
or U855 (N_855,In_1248,In_1246);
nor U856 (N_856,In_1635,In_2402);
nor U857 (N_857,In_1580,In_26);
nor U858 (N_858,In_279,In_32);
nor U859 (N_859,In_1604,In_1530);
or U860 (N_860,In_730,In_343);
and U861 (N_861,In_647,In_2138);
nor U862 (N_862,In_1158,In_1123);
nand U863 (N_863,In_1098,In_532);
nor U864 (N_864,In_7,In_998);
nand U865 (N_865,In_1053,In_1665);
xor U866 (N_866,In_2030,In_1456);
xnor U867 (N_867,In_2468,In_779);
or U868 (N_868,In_2506,In_2334);
nand U869 (N_869,In_1593,In_1282);
nor U870 (N_870,In_2750,In_2346);
and U871 (N_871,In_811,In_1645);
nor U872 (N_872,In_1586,In_1599);
or U873 (N_873,In_2981,In_1854);
nand U874 (N_874,In_1835,In_535);
nor U875 (N_875,In_505,In_1728);
nand U876 (N_876,In_1288,In_1063);
nor U877 (N_877,In_571,In_73);
nand U878 (N_878,In_2499,In_2702);
or U879 (N_879,In_2610,In_803);
or U880 (N_880,In_248,In_2494);
nand U881 (N_881,In_2351,In_1947);
nand U882 (N_882,In_274,In_1922);
xor U883 (N_883,In_196,In_2281);
xor U884 (N_884,In_2788,In_1855);
or U885 (N_885,In_2264,In_1057);
and U886 (N_886,In_1144,In_2314);
xnor U887 (N_887,In_2246,In_2419);
or U888 (N_888,In_2133,In_2213);
and U889 (N_889,In_2560,In_2165);
xnor U890 (N_890,In_90,In_716);
and U891 (N_891,In_2988,In_2536);
and U892 (N_892,In_682,In_262);
nor U893 (N_893,In_1867,In_465);
and U894 (N_894,In_1329,In_1274);
nand U895 (N_895,In_559,In_132);
nor U896 (N_896,In_1058,In_1176);
or U897 (N_897,In_326,In_1271);
nor U898 (N_898,In_900,In_1258);
nand U899 (N_899,In_2437,In_2692);
and U900 (N_900,In_2240,In_2088);
nand U901 (N_901,In_919,In_702);
or U902 (N_902,In_2598,In_2593);
nor U903 (N_903,In_2796,In_581);
xor U904 (N_904,In_358,In_2641);
or U905 (N_905,In_2267,In_1066);
or U906 (N_906,In_24,In_2674);
xor U907 (N_907,In_2,In_296);
or U908 (N_908,In_1851,In_2573);
nand U909 (N_909,In_2348,In_2814);
nand U910 (N_910,In_2716,In_89);
or U911 (N_911,In_1262,In_672);
nand U912 (N_912,In_2827,In_904);
and U913 (N_913,In_321,In_2739);
or U914 (N_914,In_1330,In_417);
nand U915 (N_915,In_1502,In_1163);
xor U916 (N_916,In_1161,In_2889);
or U917 (N_917,In_572,In_2144);
or U918 (N_918,In_1575,In_2106);
nand U919 (N_919,In_783,In_1171);
nand U920 (N_920,In_881,In_2301);
nor U921 (N_921,In_1866,In_2349);
nor U922 (N_922,In_464,In_175);
nand U923 (N_923,In_1077,In_2411);
nor U924 (N_924,In_155,In_2356);
nor U925 (N_925,In_956,In_2198);
and U926 (N_926,In_792,In_1657);
or U927 (N_927,In_1945,In_1992);
nand U928 (N_928,In_2487,In_43);
xnor U929 (N_929,In_1872,In_20);
xor U930 (N_930,In_2174,In_2162);
xor U931 (N_931,In_2310,In_2483);
nor U932 (N_932,In_1179,In_2400);
xnor U933 (N_933,In_1808,In_2903);
or U934 (N_934,In_1973,In_1103);
xnor U935 (N_935,In_2670,In_499);
nor U936 (N_936,In_2896,In_1381);
and U937 (N_937,In_1438,In_1501);
xnor U938 (N_938,In_737,In_1498);
and U939 (N_939,In_2941,In_1616);
or U940 (N_940,In_529,In_2578);
nand U941 (N_941,In_2382,In_2561);
or U942 (N_942,In_2900,In_172);
xor U943 (N_943,In_2146,In_1119);
and U944 (N_944,In_1055,In_2545);
nor U945 (N_945,In_2274,In_1797);
or U946 (N_946,In_2609,In_892);
xnor U947 (N_947,In_620,In_744);
and U948 (N_948,In_1121,In_1457);
or U949 (N_949,In_2374,In_1571);
and U950 (N_950,In_2481,In_406);
nand U951 (N_951,In_2169,In_2607);
xnor U952 (N_952,In_2145,In_340);
nand U953 (N_953,In_2279,In_2999);
nand U954 (N_954,In_2111,In_1902);
and U955 (N_955,In_2904,In_335);
and U956 (N_956,In_1159,In_763);
nand U957 (N_957,In_777,In_135);
nor U958 (N_958,In_1495,In_2324);
xor U959 (N_959,In_1568,In_627);
and U960 (N_960,In_1042,In_1863);
xnor U961 (N_961,In_2337,In_1452);
or U962 (N_962,In_2453,In_1610);
nand U963 (N_963,In_2101,In_177);
nor U964 (N_964,In_377,In_2967);
or U965 (N_965,In_2235,In_414);
and U966 (N_966,In_2780,In_1100);
nor U967 (N_967,In_2871,In_2418);
xor U968 (N_968,In_1477,In_1082);
nor U969 (N_969,In_2963,In_1888);
nor U970 (N_970,In_98,In_639);
xor U971 (N_971,In_328,In_822);
nor U972 (N_972,In_2608,In_2325);
nand U973 (N_973,In_1232,In_53);
nand U974 (N_974,In_1815,In_2415);
xnor U975 (N_975,In_400,In_1754);
or U976 (N_976,In_1684,In_2423);
xor U977 (N_977,In_2939,In_2688);
xnor U978 (N_978,In_2612,In_386);
or U979 (N_979,In_1672,In_2893);
or U980 (N_980,In_1263,In_1985);
xnor U981 (N_981,In_1354,In_1641);
nand U982 (N_982,In_2929,In_405);
nand U983 (N_983,In_1935,In_257);
or U984 (N_984,In_1662,In_398);
or U985 (N_985,In_1861,In_495);
and U986 (N_986,In_2875,In_163);
or U987 (N_987,In_590,In_2082);
xor U988 (N_988,In_2631,In_984);
or U989 (N_989,In_60,In_2568);
nor U990 (N_990,In_2186,In_318);
xnor U991 (N_991,In_1776,In_1809);
or U992 (N_992,In_120,In_526);
or U993 (N_993,In_2867,In_109);
or U994 (N_994,In_217,In_1031);
xnor U995 (N_995,In_1083,In_1443);
nand U996 (N_996,In_319,In_2178);
or U997 (N_997,In_95,In_1279);
or U998 (N_998,In_1856,In_761);
nor U999 (N_999,In_235,In_453);
nand U1000 (N_1000,In_2119,In_2427);
nor U1001 (N_1001,In_1697,In_2278);
nor U1002 (N_1002,In_1006,N_100);
or U1003 (N_1003,In_1528,N_674);
xnor U1004 (N_1004,In_1554,N_612);
nand U1005 (N_1005,In_1553,In_2456);
nor U1006 (N_1006,N_816,In_239);
or U1007 (N_1007,N_35,In_2571);
xor U1008 (N_1008,In_843,N_293);
and U1009 (N_1009,N_681,N_621);
or U1010 (N_1010,In_5,N_290);
or U1011 (N_1011,In_1105,In_2166);
or U1012 (N_1012,N_80,N_712);
nor U1013 (N_1013,In_1198,N_983);
and U1014 (N_1014,N_102,In_313);
and U1015 (N_1015,In_2365,N_867);
nor U1016 (N_1016,In_1860,N_845);
or U1017 (N_1017,N_153,In_963);
nand U1018 (N_1018,In_935,In_1577);
and U1019 (N_1019,N_512,In_2061);
nand U1020 (N_1020,N_36,In_544);
xnor U1021 (N_1021,N_302,N_518);
and U1022 (N_1022,In_1513,N_355);
nand U1023 (N_1023,N_658,N_65);
nand U1024 (N_1024,In_1825,In_1794);
nor U1025 (N_1025,In_1685,In_2908);
xnor U1026 (N_1026,In_2505,N_817);
nand U1027 (N_1027,N_317,N_428);
or U1028 (N_1028,N_743,N_170);
nor U1029 (N_1029,N_800,In_496);
or U1030 (N_1030,N_857,N_231);
and U1031 (N_1031,N_594,N_707);
nor U1032 (N_1032,N_142,In_614);
and U1033 (N_1033,N_641,N_4);
nor U1034 (N_1034,In_127,N_994);
or U1035 (N_1035,N_813,N_281);
nor U1036 (N_1036,N_502,In_2541);
and U1037 (N_1037,N_771,N_506);
and U1038 (N_1038,In_1379,In_1191);
xnor U1039 (N_1039,N_55,In_855);
nor U1040 (N_1040,In_2726,N_154);
nand U1041 (N_1041,N_308,In_70);
and U1042 (N_1042,N_378,In_2662);
nand U1043 (N_1043,N_94,N_832);
nor U1044 (N_1044,In_2534,N_866);
or U1045 (N_1045,In_928,In_2924);
nor U1046 (N_1046,In_1234,N_380);
nand U1047 (N_1047,N_559,N_461);
nor U1048 (N_1048,N_264,N_249);
nor U1049 (N_1049,N_573,N_396);
and U1050 (N_1050,N_890,In_2835);
or U1051 (N_1051,In_2196,In_2164);
nand U1052 (N_1052,N_721,In_2360);
xnor U1053 (N_1053,N_345,N_86);
and U1054 (N_1054,In_66,In_2033);
nor U1055 (N_1055,N_473,In_1695);
and U1056 (N_1056,In_985,N_495);
nor U1057 (N_1057,N_630,In_638);
xnor U1058 (N_1058,In_2032,In_303);
and U1059 (N_1059,In_1547,N_935);
or U1060 (N_1060,In_234,N_976);
or U1061 (N_1061,N_603,N_489);
nor U1062 (N_1062,In_2974,N_966);
nor U1063 (N_1063,In_330,N_894);
nand U1064 (N_1064,In_1316,In_2007);
nor U1065 (N_1065,In_2305,N_256);
nor U1066 (N_1066,In_2805,In_2338);
or U1067 (N_1067,In_934,N_487);
nor U1068 (N_1068,In_1162,N_24);
xor U1069 (N_1069,N_922,In_159);
and U1070 (N_1070,In_1475,N_953);
nor U1071 (N_1071,In_1242,N_638);
and U1072 (N_1072,In_1549,N_737);
xor U1073 (N_1073,N_454,In_34);
nand U1074 (N_1074,In_1594,N_118);
and U1075 (N_1075,In_2946,In_890);
nand U1076 (N_1076,N_323,N_401);
nor U1077 (N_1077,N_693,In_2520);
or U1078 (N_1078,In_753,N_583);
and U1079 (N_1079,N_62,N_7);
nand U1080 (N_1080,N_105,In_2436);
nand U1081 (N_1081,N_858,In_2128);
xnor U1082 (N_1082,In_254,In_1600);
or U1083 (N_1083,In_1652,N_887);
xor U1084 (N_1084,N_591,In_2691);
xnor U1085 (N_1085,In_457,In_525);
and U1086 (N_1086,In_1569,N_577);
nand U1087 (N_1087,In_2046,In_554);
xnor U1088 (N_1088,In_449,N_220);
and U1089 (N_1089,In_2181,In_1289);
nand U1090 (N_1090,In_1591,N_109);
xnor U1091 (N_1091,N_684,In_1439);
and U1092 (N_1092,N_400,In_1753);
and U1093 (N_1093,N_443,N_579);
nor U1094 (N_1094,In_1127,In_1076);
or U1095 (N_1095,N_955,N_695);
and U1096 (N_1096,In_1913,N_193);
xor U1097 (N_1097,N_811,N_337);
and U1098 (N_1098,N_79,In_2751);
or U1099 (N_1099,In_291,In_1629);
and U1100 (N_1100,In_2831,In_1995);
and U1101 (N_1101,N_213,N_554);
nand U1102 (N_1102,N_977,In_930);
nand U1103 (N_1103,N_251,N_141);
nand U1104 (N_1104,N_692,In_610);
xor U1105 (N_1105,N_725,N_644);
or U1106 (N_1106,N_675,N_654);
xnor U1107 (N_1107,N_710,In_1650);
and U1108 (N_1108,In_2737,N_783);
nor U1109 (N_1109,In_917,In_123);
or U1110 (N_1110,N_750,N_439);
xor U1111 (N_1111,N_860,N_223);
xnor U1112 (N_1112,In_1000,N_605);
xnor U1113 (N_1113,In_2193,In_2335);
nor U1114 (N_1114,N_344,N_758);
or U1115 (N_1115,N_430,N_802);
xor U1116 (N_1116,In_791,In_1188);
xor U1117 (N_1117,In_1978,In_383);
nand U1118 (N_1118,N_715,In_2762);
nor U1119 (N_1119,In_2847,In_852);
xor U1120 (N_1120,N_871,N_2);
or U1121 (N_1121,N_877,In_585);
nand U1122 (N_1122,In_1930,N_204);
nand U1123 (N_1123,In_2791,N_415);
or U1124 (N_1124,N_315,In_1157);
and U1125 (N_1125,N_23,In_2756);
nand U1126 (N_1126,N_185,N_57);
nand U1127 (N_1127,In_2225,In_347);
nand U1128 (N_1128,N_650,In_1700);
nand U1129 (N_1129,N_292,In_1266);
xnor U1130 (N_1130,N_600,In_2028);
nand U1131 (N_1131,N_910,N_107);
nor U1132 (N_1132,In_2635,In_2094);
and U1133 (N_1133,N_99,N_283);
nand U1134 (N_1134,In_2937,N_719);
nand U1135 (N_1135,N_726,N_215);
or U1136 (N_1136,N_305,N_490);
or U1137 (N_1137,N_838,N_150);
and U1138 (N_1138,In_2601,N_171);
xnor U1139 (N_1139,In_255,N_61);
and U1140 (N_1140,N_624,N_399);
and U1141 (N_1141,In_863,In_2397);
nor U1142 (N_1142,N_941,N_793);
nand U1143 (N_1143,N_766,N_818);
xor U1144 (N_1144,N_888,In_63);
nand U1145 (N_1145,In_357,In_592);
or U1146 (N_1146,In_1035,N_258);
nand U1147 (N_1147,N_884,N_85);
nand U1148 (N_1148,In_720,In_588);
or U1149 (N_1149,N_394,In_1638);
or U1150 (N_1150,In_2417,In_1331);
nor U1151 (N_1151,In_2836,In_222);
nor U1152 (N_1152,N_949,In_1075);
nand U1153 (N_1153,In_1398,N_348);
xnor U1154 (N_1154,In_1152,N_41);
xor U1155 (N_1155,In_650,N_286);
nand U1156 (N_1156,N_754,In_2894);
or U1157 (N_1157,In_1541,In_1655);
xor U1158 (N_1158,In_814,N_892);
nand U1159 (N_1159,N_22,In_119);
nand U1160 (N_1160,N_575,In_1268);
and U1161 (N_1161,N_421,In_2919);
xor U1162 (N_1162,In_533,In_1493);
and U1163 (N_1163,In_140,N_83);
nand U1164 (N_1164,In_2302,In_1917);
and U1165 (N_1165,In_1416,N_349);
nand U1166 (N_1166,N_613,In_2711);
nand U1167 (N_1167,N_374,In_703);
and U1168 (N_1168,N_581,N_797);
nor U1169 (N_1169,N_497,In_258);
and U1170 (N_1170,In_840,N_652);
nand U1171 (N_1171,N_938,In_2720);
xor U1172 (N_1172,In_1370,N_20);
or U1173 (N_1173,In_265,N_404);
and U1174 (N_1174,N_929,In_2654);
nor U1175 (N_1175,N_936,N_735);
and U1176 (N_1176,In_83,In_563);
or U1177 (N_1177,In_784,N_417);
and U1178 (N_1178,In_1730,N_601);
or U1179 (N_1179,N_311,In_1889);
nor U1180 (N_1180,In_1819,In_2885);
nor U1181 (N_1181,N_431,N_73);
xor U1182 (N_1182,N_503,In_2532);
nand U1183 (N_1183,In_1807,N_881);
nor U1184 (N_1184,In_1026,N_334);
and U1185 (N_1185,N_896,In_2587);
xnor U1186 (N_1186,In_1564,In_1914);
xnor U1187 (N_1187,N_160,In_2583);
xnor U1188 (N_1188,N_51,In_494);
or U1189 (N_1189,In_2197,N_757);
nor U1190 (N_1190,In_2962,N_143);
nand U1191 (N_1191,In_402,In_1384);
nor U1192 (N_1192,In_1769,In_2319);
nand U1193 (N_1193,In_2230,In_594);
nand U1194 (N_1194,N_151,In_1426);
xor U1195 (N_1195,N_633,In_1986);
and U1196 (N_1196,N_324,In_144);
or U1197 (N_1197,N_460,In_2172);
nand U1198 (N_1198,N_169,N_198);
xor U1199 (N_1199,In_350,N_739);
and U1200 (N_1200,In_327,N_263);
xnor U1201 (N_1201,In_1921,In_867);
or U1202 (N_1202,N_610,In_1309);
nand U1203 (N_1203,In_362,In_42);
or U1204 (N_1204,N_689,N_534);
nand U1205 (N_1205,In_1301,In_849);
nor U1206 (N_1206,In_1140,In_595);
and U1207 (N_1207,N_720,N_199);
or U1208 (N_1208,N_125,N_978);
or U1209 (N_1209,In_2666,In_2766);
xor U1210 (N_1210,In_1010,In_1344);
nor U1211 (N_1211,N_218,N_82);
or U1212 (N_1212,N_691,In_989);
and U1213 (N_1213,N_709,N_235);
or U1214 (N_1214,N_898,In_329);
nand U1215 (N_1215,In_359,In_36);
xnor U1216 (N_1216,In_2787,N_596);
xnor U1217 (N_1217,In_2639,N_916);
nand U1218 (N_1218,In_302,In_2625);
and U1219 (N_1219,N_851,N_452);
nor U1220 (N_1220,In_2829,N_98);
or U1221 (N_1221,N_243,In_129);
nor U1222 (N_1222,In_719,N_177);
nor U1223 (N_1223,N_951,N_724);
and U1224 (N_1224,N_42,In_2475);
nand U1225 (N_1225,In_2825,N_257);
nand U1226 (N_1226,In_1303,N_446);
and U1227 (N_1227,N_919,In_1211);
xor U1228 (N_1228,In_2108,N_493);
and U1229 (N_1229,N_276,N_456);
nand U1230 (N_1230,In_2135,N_216);
or U1231 (N_1231,In_1567,In_124);
or U1232 (N_1232,N_227,N_32);
or U1233 (N_1233,N_546,In_2156);
and U1234 (N_1234,In_1603,In_1559);
nand U1235 (N_1235,N_161,N_406);
nor U1236 (N_1236,N_555,N_934);
nand U1237 (N_1237,N_786,N_361);
xor U1238 (N_1238,N_318,N_217);
nor U1239 (N_1239,In_1551,N_694);
nor U1240 (N_1240,N_729,N_950);
nand U1241 (N_1241,In_924,In_443);
nor U1242 (N_1242,In_58,N_699);
and U1243 (N_1243,In_2782,In_462);
nand U1244 (N_1244,In_955,In_2315);
or U1245 (N_1245,In_1286,N_184);
xor U1246 (N_1246,In_1614,N_137);
nand U1247 (N_1247,N_368,N_532);
or U1248 (N_1248,In_1428,N_343);
and U1249 (N_1249,In_1206,In_923);
nor U1250 (N_1250,N_873,In_2982);
and U1251 (N_1251,In_2510,In_2627);
nor U1252 (N_1252,N_520,In_2370);
or U1253 (N_1253,N_874,In_1626);
or U1254 (N_1254,N_551,N_433);
or U1255 (N_1255,N_542,In_1317);
nor U1256 (N_1256,N_533,N_999);
nand U1257 (N_1257,N_104,In_1966);
nand U1258 (N_1258,N_672,N_360);
xnor U1259 (N_1259,N_425,N_882);
nor U1260 (N_1260,In_1745,In_1079);
or U1261 (N_1261,In_874,In_2630);
xnor U1262 (N_1262,In_506,N_72);
nand U1263 (N_1263,In_1074,In_2589);
or U1264 (N_1264,In_2860,In_121);
xor U1265 (N_1265,N_746,N_176);
or U1266 (N_1266,N_144,N_3);
xnor U1267 (N_1267,N_992,In_209);
nand U1268 (N_1268,In_460,In_2958);
and U1269 (N_1269,In_2585,N_434);
and U1270 (N_1270,N_278,N_56);
and U1271 (N_1271,In_2098,N_0);
xnor U1272 (N_1272,N_31,N_996);
nor U1273 (N_1273,In_1306,In_1581);
nor U1274 (N_1274,In_391,N_195);
nor U1275 (N_1275,N_78,N_440);
nand U1276 (N_1276,In_1897,In_1555);
and U1277 (N_1277,N_333,In_633);
nor U1278 (N_1278,In_772,In_1418);
xnor U1279 (N_1279,In_1469,In_1448);
xnor U1280 (N_1280,N_597,N_856);
nand U1281 (N_1281,N_498,In_2238);
and U1282 (N_1282,In_1637,In_2952);
nor U1283 (N_1283,N_623,N_885);
nor U1284 (N_1284,In_1110,In_1668);
nand U1285 (N_1285,N_505,N_165);
xor U1286 (N_1286,N_148,N_622);
nand U1287 (N_1287,In_2790,In_2606);
xor U1288 (N_1288,N_155,In_2707);
or U1289 (N_1289,In_59,N_298);
and U1290 (N_1290,N_736,N_408);
xnor U1291 (N_1291,N_212,In_2622);
and U1292 (N_1292,N_116,In_583);
and U1293 (N_1293,N_639,In_1153);
nand U1294 (N_1294,N_307,N_48);
xnor U1295 (N_1295,In_2840,In_1658);
xor U1296 (N_1296,In_6,In_2926);
xnor U1297 (N_1297,In_616,N_477);
nand U1298 (N_1298,In_2282,In_1678);
nand U1299 (N_1299,In_227,In_466);
nor U1300 (N_1300,N_321,In_2508);
nand U1301 (N_1301,N_145,N_112);
xnor U1302 (N_1302,N_167,In_1991);
and U1303 (N_1303,In_619,N_727);
nand U1304 (N_1304,N_273,N_588);
xor U1305 (N_1305,In_1172,In_2254);
or U1306 (N_1306,In_2752,In_116);
and U1307 (N_1307,N_548,In_1052);
xnor U1308 (N_1308,N_266,In_704);
and U1309 (N_1309,N_825,In_1875);
and U1310 (N_1310,In_1789,In_695);
xor U1311 (N_1311,N_162,N_335);
and U1312 (N_1312,In_421,N_312);
nor U1313 (N_1313,N_523,In_2121);
nor U1314 (N_1314,In_1540,N_226);
xnor U1315 (N_1315,In_2717,In_2533);
nand U1316 (N_1316,In_641,In_376);
nor U1317 (N_1317,In_2096,N_913);
nand U1318 (N_1318,In_152,In_1235);
xor U1319 (N_1319,In_927,In_2241);
and U1320 (N_1320,In_2781,In_634);
nor U1321 (N_1321,In_2075,In_1848);
and U1322 (N_1322,In_2023,N_722);
xor U1323 (N_1323,In_2824,N_453);
nor U1324 (N_1324,In_1463,In_475);
and U1325 (N_1325,N_937,In_1405);
nor U1326 (N_1326,N_981,In_2068);
nor U1327 (N_1327,N_111,N_560);
nand U1328 (N_1328,N_367,N_812);
xnor U1329 (N_1329,N_717,N_407);
xnor U1330 (N_1330,In_1067,In_2868);
nand U1331 (N_1331,In_2422,N_127);
or U1332 (N_1332,N_842,In_2378);
or U1333 (N_1333,N_465,In_1190);
or U1334 (N_1334,N_846,N_905);
nand U1335 (N_1335,N_69,N_429);
and U1336 (N_1336,In_1936,N_731);
and U1337 (N_1337,In_1267,In_519);
and U1338 (N_1338,N_481,N_186);
and U1339 (N_1339,In_552,N_526);
nand U1340 (N_1340,In_1967,N_636);
or U1341 (N_1341,In_316,In_1533);
nand U1342 (N_1342,In_461,N_110);
or U1343 (N_1343,In_699,N_87);
or U1344 (N_1344,N_15,In_1724);
or U1345 (N_1345,N_745,N_471);
and U1346 (N_1346,N_804,In_1673);
xnor U1347 (N_1347,In_1813,In_1811);
and U1348 (N_1348,In_2322,N_682);
xnor U1349 (N_1349,N_377,N_314);
nand U1350 (N_1350,In_2516,N_964);
xnor U1351 (N_1351,N_696,N_229);
nor U1352 (N_1352,N_920,In_653);
nor U1353 (N_1353,In_1862,N_664);
and U1354 (N_1354,N_66,In_1883);
and U1355 (N_1355,In_1295,N_174);
nor U1356 (N_1356,In_603,In_2039);
nand U1357 (N_1357,In_2044,N_187);
xnor U1358 (N_1358,In_356,N_210);
nor U1359 (N_1359,N_587,In_511);
nor U1360 (N_1360,N_422,In_1406);
and U1361 (N_1361,N_952,In_1251);
nor U1362 (N_1362,N_138,N_25);
nand U1363 (N_1363,In_490,In_1563);
nand U1364 (N_1364,In_1216,N_395);
and U1365 (N_1365,In_2069,In_2857);
xnor U1366 (N_1366,N_382,In_1983);
or U1367 (N_1367,In_557,In_560);
and U1368 (N_1368,In_372,N_798);
xnor U1369 (N_1369,In_551,N_975);
nand U1370 (N_1370,N_371,In_1345);
and U1371 (N_1371,In_2395,N_19);
or U1372 (N_1372,In_261,In_721);
nand U1373 (N_1373,N_232,N_595);
or U1374 (N_1374,N_982,N_59);
nand U1375 (N_1375,In_2599,In_2910);
or U1376 (N_1376,N_172,In_210);
nand U1377 (N_1377,N_755,N_807);
nor U1378 (N_1378,In_1189,N_826);
nor U1379 (N_1379,N_764,In_2157);
nand U1380 (N_1380,In_2851,In_314);
or U1381 (N_1381,In_480,N_680);
or U1382 (N_1382,N_28,In_1786);
or U1383 (N_1383,In_447,In_195);
or U1384 (N_1384,In_1349,N_790);
or U1385 (N_1385,In_565,In_244);
and U1386 (N_1386,N_346,In_1449);
and U1387 (N_1387,N_54,N_820);
xnor U1388 (N_1388,N_413,In_1290);
nand U1389 (N_1389,N_643,N_397);
xnor U1390 (N_1390,N_906,N_547);
xnor U1391 (N_1391,N_599,N_611);
nor U1392 (N_1392,N_960,In_617);
nor U1393 (N_1393,In_151,In_2864);
or U1394 (N_1394,N_646,N_509);
xnor U1395 (N_1395,In_190,N_49);
and U1396 (N_1396,N_540,In_2748);
nand U1397 (N_1397,In_157,In_2708);
nand U1398 (N_1398,N_618,In_1199);
nand U1399 (N_1399,N_84,In_1570);
xnor U1400 (N_1400,In_2195,N_995);
and U1401 (N_1401,N_987,N_524);
nand U1402 (N_1402,In_1693,N_760);
xnor U1403 (N_1403,In_1613,In_2549);
xor U1404 (N_1404,N_225,In_787);
nand U1405 (N_1405,In_187,In_770);
xor U1406 (N_1406,N_815,N_676);
nand U1407 (N_1407,N_246,N_219);
or U1408 (N_1408,N_925,In_2732);
or U1409 (N_1409,N_178,In_2567);
nor U1410 (N_1410,In_1373,In_1363);
or U1411 (N_1411,In_1001,In_1790);
or U1412 (N_1412,N_781,N_545);
nor U1413 (N_1413,In_2775,N_158);
nor U1414 (N_1414,In_2555,N_244);
or U1415 (N_1415,In_718,N_224);
nor U1416 (N_1416,In_2594,N_277);
xnor U1417 (N_1417,In_1545,In_611);
xor U1418 (N_1418,N_609,In_1080);
nand U1419 (N_1419,N_847,In_1093);
xnor U1420 (N_1420,N_656,In_211);
xor U1421 (N_1421,In_467,In_2547);
xnor U1422 (N_1422,N_146,In_808);
and U1423 (N_1423,In_92,N_844);
nor U1424 (N_1424,In_2140,In_2862);
or U1425 (N_1425,In_757,N_117);
nor U1426 (N_1426,N_991,N_634);
or U1427 (N_1427,N_961,N_663);
xnor U1428 (N_1428,N_801,In_679);
nor U1429 (N_1429,N_274,In_448);
xor U1430 (N_1430,N_275,In_2563);
nand U1431 (N_1431,In_1360,In_866);
xnor U1432 (N_1432,In_2013,In_1800);
and U1433 (N_1433,In_1455,N_558);
nor U1434 (N_1434,In_247,N_998);
nand U1435 (N_1435,In_1831,N_491);
nand U1436 (N_1436,In_492,In_698);
and U1437 (N_1437,In_2488,N_33);
or U1438 (N_1438,In_68,N_436);
nand U1439 (N_1439,N_432,N_209);
nand U1440 (N_1440,N_752,In_1136);
or U1441 (N_1441,In_2884,N_89);
nand U1442 (N_1442,In_424,N_854);
xnor U1443 (N_1443,In_1882,N_864);
nand U1444 (N_1444,N_879,In_2443);
xor U1445 (N_1445,N_233,N_147);
or U1446 (N_1446,N_747,N_921);
xor U1447 (N_1447,In_47,In_841);
nor U1448 (N_1448,In_853,N_859);
and U1449 (N_1449,In_2820,In_2469);
or U1450 (N_1450,In_977,N_480);
nor U1451 (N_1451,N_901,N_389);
or U1452 (N_1452,In_323,In_2192);
and U1453 (N_1453,N_140,N_569);
nand U1454 (N_1454,N_589,In_743);
and U1455 (N_1455,N_296,In_959);
and U1456 (N_1456,In_2826,N_900);
or U1457 (N_1457,N_530,In_1097);
nor U1458 (N_1458,In_231,N_565);
xnor U1459 (N_1459,In_1215,N_267);
nor U1460 (N_1460,N_88,N_188);
and U1461 (N_1461,In_1129,In_878);
and U1462 (N_1462,In_1321,N_386);
nand U1463 (N_1463,N_794,In_707);
xnor U1464 (N_1464,In_574,In_2223);
nor U1465 (N_1465,N_385,In_727);
nand U1466 (N_1466,N_778,N_34);
xnor U1467 (N_1467,In_1192,In_1926);
and U1468 (N_1468,N_862,N_124);
xor U1469 (N_1469,In_856,N_372);
and U1470 (N_1470,N_670,N_593);
nor U1471 (N_1471,N_50,N_527);
or U1472 (N_1472,In_2093,N_668);
and U1473 (N_1473,N_326,N_679);
nand U1474 (N_1474,N_427,In_929);
nor U1475 (N_1475,N_660,In_845);
nand U1476 (N_1476,In_1256,N_568);
or U1477 (N_1477,N_829,In_1253);
xnor U1478 (N_1478,In_57,N_853);
nand U1479 (N_1479,In_2514,N_27);
nand U1480 (N_1480,In_1218,N_592);
nand U1481 (N_1481,N_849,N_272);
or U1482 (N_1482,N_384,In_2713);
nor U1483 (N_1483,N_686,In_1285);
or U1484 (N_1484,In_1328,In_1415);
xnor U1485 (N_1485,In_709,In_80);
or U1486 (N_1486,In_1660,In_2832);
and U1487 (N_1487,N_713,In_1397);
nor U1488 (N_1488,In_2955,In_1411);
or U1489 (N_1489,In_1050,In_112);
xnor U1490 (N_1490,N_514,In_1908);
xnor U1491 (N_1491,N_972,In_2289);
xnor U1492 (N_1492,N_915,In_2153);
or U1493 (N_1493,In_1887,In_932);
and U1494 (N_1494,In_2117,In_1202);
xor U1495 (N_1495,N_75,N_482);
nand U1496 (N_1496,In_799,N_984);
nor U1497 (N_1497,In_2693,N_553);
nand U1498 (N_1498,N_269,N_511);
nor U1499 (N_1499,N_451,N_435);
xnor U1500 (N_1500,In_2250,In_1407);
or U1501 (N_1501,In_2253,N_827);
nor U1502 (N_1502,N_761,N_718);
nand U1503 (N_1503,In_997,N_259);
nand U1504 (N_1504,In_2576,N_521);
or U1505 (N_1505,In_1195,In_55);
or U1506 (N_1506,N_942,In_437);
and U1507 (N_1507,N_90,In_1318);
nand U1508 (N_1508,In_517,In_426);
nand U1509 (N_1509,In_2846,In_2073);
xnor U1510 (N_1510,In_926,N_954);
or U1511 (N_1511,In_2449,In_2523);
or U1512 (N_1512,N_784,N_485);
and U1513 (N_1513,N_476,N_130);
xnor U1514 (N_1514,N_309,N_208);
and U1515 (N_1515,N_957,In_899);
nand U1516 (N_1516,N_891,In_2509);
nor U1517 (N_1517,N_732,N_364);
nand U1518 (N_1518,In_1839,N_175);
nand U1519 (N_1519,In_2986,In_833);
and U1520 (N_1520,In_268,N_803);
xnor U1521 (N_1521,In_2399,N_702);
and U1522 (N_1522,N_458,N_53);
nand U1523 (N_1523,N_831,N_132);
or U1524 (N_1524,N_383,In_1646);
and U1525 (N_1525,In_2873,In_1842);
and U1526 (N_1526,N_280,In_663);
xor U1527 (N_1527,In_1738,N_529);
or U1528 (N_1528,In_1606,N_833);
nand U1529 (N_1529,N_627,In_684);
and U1530 (N_1530,N_683,N_767);
nand U1531 (N_1531,In_1332,N_850);
nand U1532 (N_1532,N_789,In_823);
nand U1533 (N_1533,N_206,N_580);
and U1534 (N_1534,N_234,N_418);
nand U1535 (N_1535,In_78,N_564);
and U1536 (N_1536,N_375,N_328);
nor U1537 (N_1537,In_1682,In_2979);
nor U1538 (N_1538,N_133,In_1489);
nor U1539 (N_1539,N_543,In_1994);
nor U1540 (N_1540,In_1998,In_631);
nor U1541 (N_1541,In_2704,In_1353);
or U1542 (N_1542,N_708,N_848);
nand U1543 (N_1543,In_434,In_1529);
xor U1544 (N_1544,N_248,In_446);
nor U1545 (N_1545,N_420,N_52);
nor U1546 (N_1546,N_799,In_2179);
and U1547 (N_1547,N_447,N_411);
or U1548 (N_1548,N_478,In_1413);
nand U1549 (N_1549,N_993,In_2724);
nor U1550 (N_1550,N_963,In_2201);
and U1551 (N_1551,In_655,N_241);
nand U1552 (N_1552,In_2215,N_93);
nor U1553 (N_1553,N_974,N_330);
and U1554 (N_1554,In_660,N_810);
nand U1555 (N_1555,N_134,N_742);
and U1556 (N_1556,In_2531,In_2425);
nand U1557 (N_1557,N_619,N_541);
nor U1558 (N_1558,In_2445,In_2504);
xor U1559 (N_1559,In_2367,N_470);
and U1560 (N_1560,In_1272,N_625);
or U1561 (N_1561,N_777,In_1791);
or U1562 (N_1562,N_63,N_123);
and U1563 (N_1563,In_2591,N_990);
or U1564 (N_1564,In_39,In_1);
xnor U1565 (N_1565,In_1843,In_2554);
and U1566 (N_1566,N_403,N_647);
and U1567 (N_1567,N_563,N_247);
xnor U1568 (N_1568,In_1583,N_340);
and U1569 (N_1569,N_252,N_806);
xor U1570 (N_1570,In_1892,In_392);
or U1571 (N_1571,In_2386,N_95);
nor U1572 (N_1572,In_1394,N_716);
xnor U1573 (N_1573,N_909,N_632);
and U1574 (N_1574,In_2902,N_586);
xor U1575 (N_1575,In_2712,In_105);
and U1576 (N_1576,In_686,N_115);
nor U1577 (N_1577,N_759,In_1032);
xor U1578 (N_1578,In_156,N_464);
and U1579 (N_1579,N_295,In_2122);
nor U1580 (N_1580,In_331,In_309);
nor U1581 (N_1581,N_18,N_897);
nand U1582 (N_1582,N_304,N_43);
xor U1583 (N_1583,In_2973,In_854);
xor U1584 (N_1584,In_1299,N_327);
and U1585 (N_1585,N_354,N_103);
or U1586 (N_1586,In_1287,N_902);
nand U1587 (N_1587,N_504,In_2392);
xnor U1588 (N_1588,N_410,N_129);
or U1589 (N_1589,N_828,N_669);
or U1590 (N_1590,N_352,In_3);
or U1591 (N_1591,N_119,In_2773);
or U1592 (N_1592,N_562,N_787);
nand U1593 (N_1593,In_1598,In_2626);
or U1594 (N_1594,N_294,N_886);
or U1595 (N_1595,In_395,N_661);
or U1596 (N_1596,N_701,In_40);
nor U1597 (N_1597,N_561,In_1071);
xnor U1598 (N_1598,N_287,In_1214);
and U1599 (N_1599,N_282,In_2685);
nor U1600 (N_1600,In_512,N_253);
and U1601 (N_1601,N_893,N_773);
and U1602 (N_1602,N_96,N_775);
xor U1603 (N_1603,In_1628,N_517);
or U1604 (N_1604,In_1343,N_365);
nand U1605 (N_1605,In_2331,N_245);
and U1606 (N_1606,N_336,In_367);
nand U1607 (N_1607,In_2208,N_642);
nor U1608 (N_1608,N_614,In_951);
xnor U1609 (N_1609,In_618,In_2839);
and U1610 (N_1610,N_837,N_262);
or U1611 (N_1611,N_830,In_2316);
and U1612 (N_1612,N_388,N_980);
nand U1613 (N_1613,In_2484,In_1762);
nor U1614 (N_1614,In_1996,N_332);
xnor U1615 (N_1615,In_2393,N_76);
and U1616 (N_1616,N_538,N_631);
or U1617 (N_1617,N_968,N_748);
and U1618 (N_1618,In_2858,In_271);
nand U1619 (N_1619,In_1627,N_338);
nand U1620 (N_1620,N_369,N_8);
xor U1621 (N_1621,N_191,In_2987);
or U1622 (N_1622,N_472,N_970);
or U1623 (N_1623,N_47,N_13);
nor U1624 (N_1624,In_1250,In_2239);
or U1625 (N_1625,In_1773,In_2248);
nor U1626 (N_1626,In_280,N_863);
or U1627 (N_1627,In_649,In_308);
and U1628 (N_1628,In_1229,N_519);
and U1629 (N_1629,N_617,N_391);
nand U1630 (N_1630,In_1116,N_319);
and U1631 (N_1631,In_1847,N_776);
and U1632 (N_1632,N_659,In_2327);
or U1633 (N_1633,In_431,N_576);
nor U1634 (N_1634,In_936,In_2584);
nor U1635 (N_1635,In_491,N_300);
xor U1636 (N_1636,N_299,N_899);
nor U1637 (N_1637,N_156,In_2034);
xnor U1638 (N_1638,N_821,In_2597);
or U1639 (N_1639,N_671,N_416);
nand U1640 (N_1640,In_197,In_1679);
xnor U1641 (N_1641,In_2736,N_353);
or U1642 (N_1642,In_389,N_381);
xnor U1643 (N_1643,In_1636,In_950);
xor U1644 (N_1644,N_779,In_1327);
nand U1645 (N_1645,In_2785,N_768);
xor U1646 (N_1646,N_200,In_174);
and U1647 (N_1647,N_402,N_762);
or U1648 (N_1648,In_2057,In_378);
and U1649 (N_1649,N_30,In_64);
and U1650 (N_1650,In_404,In_1243);
xnor U1651 (N_1651,N_450,In_504);
nand U1652 (N_1652,In_2019,In_2619);
and U1653 (N_1653,In_31,In_2800);
and U1654 (N_1654,In_2914,N_194);
nor U1655 (N_1655,In_2244,In_1223);
nor U1656 (N_1656,N_598,In_859);
nand U1657 (N_1657,N_44,In_345);
nor U1658 (N_1658,N_616,In_185);
xor U1659 (N_1659,In_1323,In_2124);
and U1660 (N_1660,In_837,In_879);
and U1661 (N_1661,In_2569,In_428);
xor U1662 (N_1662,In_1342,N_772);
nand U1663 (N_1663,N_749,N_685);
nor U1664 (N_1664,In_2797,In_2783);
xor U1665 (N_1665,N_139,In_2077);
and U1666 (N_1666,N_236,N_785);
nor U1667 (N_1667,N_424,N_516);
nor U1668 (N_1668,In_2458,N_149);
and U1669 (N_1669,N_932,In_640);
and U1670 (N_1670,In_1228,N_880);
nand U1671 (N_1671,In_2961,In_16);
and U1672 (N_1672,N_515,N_483);
and U1673 (N_1673,N_173,N_571);
nor U1674 (N_1674,N_791,In_1968);
xor U1675 (N_1675,N_769,N_409);
nor U1676 (N_1676,In_2496,In_1470);
nor U1677 (N_1677,In_2149,In_200);
nand U1678 (N_1678,N_255,N_131);
xnor U1679 (N_1679,N_626,In_1940);
xor U1680 (N_1680,In_2339,N_923);
xor U1681 (N_1681,N_740,N_753);
nand U1682 (N_1682,In_1720,In_2237);
or U1683 (N_1683,N_157,In_970);
and U1684 (N_1684,N_927,In_48);
and U1685 (N_1685,N_92,In_882);
or U1686 (N_1686,In_2176,In_2372);
and U1687 (N_1687,N_303,In_1526);
xnor U1688 (N_1688,N_60,In_2042);
or U1689 (N_1689,In_2304,In_1798);
nor U1690 (N_1690,In_2168,N_585);
and U1691 (N_1691,In_1804,N_114);
nand U1692 (N_1692,N_604,N_122);
xnor U1693 (N_1693,N_260,In_479);
nand U1694 (N_1694,In_925,In_2242);
and U1695 (N_1695,N_590,N_835);
or U1696 (N_1696,In_2786,N_912);
nor U1697 (N_1697,N_70,N_492);
nor U1698 (N_1698,In_1441,N_14);
and U1699 (N_1699,In_1542,In_1761);
nor U1700 (N_1700,In_2621,In_1870);
nor U1701 (N_1701,In_1690,In_2219);
or U1702 (N_1702,N_121,N_744);
or U1703 (N_1703,In_49,In_2210);
nand U1704 (N_1704,In_2457,In_2970);
and U1705 (N_1705,N_166,In_2983);
nor U1706 (N_1706,N_320,In_644);
or U1707 (N_1707,N_510,In_2944);
nor U1708 (N_1708,In_2792,In_366);
nand U1709 (N_1709,N_205,N_843);
xor U1710 (N_1710,N_582,In_212);
or U1711 (N_1711,N_872,N_865);
nor U1712 (N_1712,In_556,N_876);
nand U1713 (N_1713,N_163,In_1391);
or U1714 (N_1714,N_370,In_352);
xnor U1715 (N_1715,In_1938,In_1177);
nand U1716 (N_1716,In_1766,In_1124);
and U1717 (N_1717,In_1313,N_822);
xnor U1718 (N_1718,In_2243,N_97);
or U1719 (N_1719,N_653,In_1979);
and U1720 (N_1720,N_868,N_928);
nand U1721 (N_1721,N_108,N_462);
or U1722 (N_1722,N_10,N_733);
nand U1723 (N_1723,In_2863,N_271);
or U1724 (N_1724,N_943,In_2806);
nor U1725 (N_1725,N_640,In_325);
or U1726 (N_1726,N_557,N_347);
and U1727 (N_1727,In_2371,N_734);
nor U1728 (N_1728,N_878,N_306);
and U1729 (N_1729,In_1217,N_468);
nor U1730 (N_1730,N_552,In_1970);
and U1731 (N_1731,N_475,In_1185);
nor U1732 (N_1732,N_723,In_2177);
or U1733 (N_1733,N_40,N_459);
or U1734 (N_1734,In_2259,In_2616);
xnor U1735 (N_1735,N_500,In_2795);
xnor U1736 (N_1736,N_68,N_128);
nor U1737 (N_1737,In_609,In_2817);
and U1738 (N_1738,In_420,N_228);
nor U1739 (N_1739,In_146,N_449);
or U1740 (N_1740,N_437,N_792);
or U1741 (N_1741,In_2521,In_2990);
nor U1742 (N_1742,In_1325,N_351);
or U1743 (N_1743,In_2206,N_824);
xor U1744 (N_1744,In_246,N_706);
or U1745 (N_1745,N_423,N_180);
nand U1746 (N_1746,N_924,N_728);
xnor U1747 (N_1747,In_2526,In_2330);
nand U1748 (N_1748,N_819,In_249);
xnor U1749 (N_1749,N_357,In_28);
nand U1750 (N_1750,N_945,N_917);
xnor U1751 (N_1751,In_2474,N_285);
and U1752 (N_1752,In_626,In_752);
and U1753 (N_1753,In_2131,In_503);
or U1754 (N_1754,N_651,In_1142);
or U1755 (N_1755,In_82,In_183);
xnor U1756 (N_1756,N_291,In_1340);
and U1757 (N_1757,In_2854,N_64);
nor U1758 (N_1758,In_184,N_301);
and U1759 (N_1759,In_1041,N_628);
xnor U1760 (N_1760,In_473,In_10);
xor U1761 (N_1761,N_488,In_741);
nor U1762 (N_1762,N_101,N_197);
nor U1763 (N_1763,In_108,In_21);
and U1764 (N_1764,N_667,N_152);
and U1765 (N_1765,N_376,N_183);
or U1766 (N_1766,N_445,In_1886);
nand U1767 (N_1767,In_807,N_499);
xor U1768 (N_1768,N_796,N_238);
or U1769 (N_1769,N_242,In_1111);
and U1770 (N_1770,In_2473,In_1960);
nor U1771 (N_1771,In_1348,In_1625);
nor U1772 (N_1772,In_1582,In_1432);
xor U1773 (N_1773,In_1588,N_572);
or U1774 (N_1774,In_1982,In_488);
nor U1775 (N_1775,In_2207,In_1244);
nand U1776 (N_1776,N_190,N_947);
xnor U1777 (N_1777,In_817,In_1717);
or U1778 (N_1778,N_841,N_329);
xor U1779 (N_1779,In_1298,N_931);
nor U1780 (N_1780,In_2828,In_1956);
nand U1781 (N_1781,N_649,In_834);
nand U1782 (N_1782,N_214,N_635);
nor U1783 (N_1783,N_911,N_297);
and U1784 (N_1784,N_12,N_780);
and U1785 (N_1785,N_648,N_539);
or U1786 (N_1786,In_978,In_2155);
and U1787 (N_1787,In_1377,N_484);
xor U1788 (N_1788,N_239,In_717);
or U1789 (N_1789,In_1371,In_2686);
nor U1790 (N_1790,In_578,In_2881);
xor U1791 (N_1791,N_513,N_965);
or U1792 (N_1792,N_21,In_1375);
nor U1793 (N_1793,In_518,In_1464);
nor U1794 (N_1794,In_1748,N_918);
nand U1795 (N_1795,In_1043,In_2385);
or U1796 (N_1796,N_971,In_2303);
nor U1797 (N_1797,In_2570,N_985);
nand U1798 (N_1798,N_313,N_342);
nor U1799 (N_1799,N_730,N_608);
nor U1800 (N_1800,N_366,N_135);
or U1801 (N_1801,N_763,In_673);
nand U1802 (N_1802,N_522,In_214);
xor U1803 (N_1803,N_883,N_697);
nor U1804 (N_1804,In_2695,N_29);
or U1805 (N_1805,N_795,In_2522);
nor U1806 (N_1806,N_690,N_930);
and U1807 (N_1807,N_770,In_1447);
nand U1808 (N_1808,N_655,N_997);
nor U1809 (N_1809,N_288,N_46);
and U1810 (N_1810,In_1694,N_181);
xor U1811 (N_1811,In_2694,In_2501);
or U1812 (N_1812,N_363,N_159);
nor U1813 (N_1813,In_134,In_233);
nor U1814 (N_1814,In_2892,N_106);
xor U1815 (N_1815,In_2464,In_815);
xnor U1816 (N_1816,In_1722,N_58);
or U1817 (N_1817,In_1400,In_2951);
and U1818 (N_1818,In_2010,In_949);
nand U1819 (N_1819,In_1073,In_2558);
and U1820 (N_1820,N_549,N_438);
nor U1821 (N_1821,N_331,In_528);
nor U1822 (N_1822,N_508,In_1386);
nor U1823 (N_1823,In_860,In_256);
nor U1824 (N_1824,N_678,In_2409);
xnor U1825 (N_1825,N_765,In_1049);
nor U1826 (N_1826,In_1834,N_455);
nor U1827 (N_1827,In_2865,N_537);
or U1828 (N_1828,In_1178,In_2557);
or U1829 (N_1829,N_441,N_808);
xnor U1830 (N_1830,N_221,N_673);
or U1831 (N_1831,In_2180,In_2874);
or U1832 (N_1832,In_2396,N_189);
xor U1833 (N_1833,N_986,In_2819);
xor U1834 (N_1834,N_466,N_756);
or U1835 (N_1835,N_967,N_914);
nor U1836 (N_1836,In_1036,N_645);
or U1837 (N_1837,In_401,In_2455);
nor U1838 (N_1838,N_607,N_834);
nand U1839 (N_1839,N_316,In_527);
and U1840 (N_1840,In_1092,In_606);
xnor U1841 (N_1841,In_394,N_254);
and U1842 (N_1842,In_283,In_2491);
nand U1843 (N_1843,In_2085,N_805);
or U1844 (N_1844,In_2403,N_356);
xor U1845 (N_1845,In_1484,In_2110);
nand U1846 (N_1846,N_426,In_2620);
xor U1847 (N_1847,N_444,N_861);
and U1848 (N_1848,N_5,In_1605);
and U1849 (N_1849,In_2994,In_295);
nor U1850 (N_1850,In_2923,N_933);
nor U1851 (N_1851,In_2362,N_855);
nand U1852 (N_1852,N_358,In_276);
nand U1853 (N_1853,In_1525,N_265);
nand U1854 (N_1854,N_989,In_765);
xnor U1855 (N_1855,In_1112,N_113);
nand U1856 (N_1856,In_937,N_875);
or U1857 (N_1857,N_474,N_907);
nand U1858 (N_1858,N_751,In_1669);
nor U1859 (N_1859,In_477,N_284);
or U1860 (N_1860,N_657,N_405);
nor U1861 (N_1861,In_220,N_136);
nand U1862 (N_1862,N_398,In_2672);
nor U1863 (N_1863,In_2566,N_179);
xor U1864 (N_1864,N_387,In_338);
and U1865 (N_1865,N_393,In_1959);
and U1866 (N_1866,N_741,In_738);
and U1867 (N_1867,In_809,In_1916);
and U1868 (N_1868,N_120,N_944);
and U1869 (N_1869,In_1920,N_700);
nor U1870 (N_1870,N_889,In_2848);
or U1871 (N_1871,In_1760,In_288);
and U1872 (N_1872,In_2354,In_2002);
xnor U1873 (N_1873,In_2995,In_240);
and U1874 (N_1874,In_1634,In_2479);
nor U1875 (N_1875,N_230,N_494);
or U1876 (N_1876,N_956,In_2912);
nor U1877 (N_1877,In_2770,In_542);
nor U1878 (N_1878,N_602,In_1008);
nand U1879 (N_1879,N_414,In_2355);
nand U1880 (N_1880,N_26,In_2746);
xnor U1881 (N_1881,In_284,In_2336);
or U1882 (N_1882,N_240,In_861);
nand U1883 (N_1883,In_1757,In_2565);
and U1884 (N_1884,N_774,N_507);
xor U1885 (N_1885,In_993,In_482);
and U1886 (N_1886,N_486,N_988);
and U1887 (N_1887,In_1931,N_71);
xor U1888 (N_1888,In_545,In_1222);
nor U1889 (N_1889,N_469,In_2050);
and U1890 (N_1890,In_1254,In_1849);
and U1891 (N_1891,N_6,In_1957);
nor U1892 (N_1892,N_442,N_962);
and U1893 (N_1893,N_350,N_279);
xnor U1894 (N_1894,N_908,In_122);
nand U1895 (N_1895,In_991,In_584);
and U1896 (N_1896,N_620,N_77);
and U1897 (N_1897,N_711,N_339);
or U1898 (N_1898,N_688,In_2760);
nor U1899 (N_1899,N_556,N_852);
or U1900 (N_1900,In_1101,In_2005);
nand U1901 (N_1901,N_250,In_1095);
or U1902 (N_1902,N_531,In_1380);
nor U1903 (N_1903,In_2125,In_1858);
or U1904 (N_1904,In_454,N_979);
or U1905 (N_1905,N_196,N_81);
nor U1906 (N_1906,N_419,In_2130);
xor U1907 (N_1907,N_869,N_67);
nor U1908 (N_1908,N_182,In_760);
xnor U1909 (N_1909,In_1166,In_2255);
and U1910 (N_1910,N_615,N_895);
or U1911 (N_1911,In_1949,N_958);
xor U1912 (N_1912,In_2480,In_1086);
or U1913 (N_1913,N_16,N_325);
xnor U1914 (N_1914,N_939,In_2049);
nand U1915 (N_1915,In_2368,In_275);
and U1916 (N_1916,In_2913,N_310);
nor U1917 (N_1917,N_578,N_662);
xor U1918 (N_1918,N_973,N_168);
and U1919 (N_1919,In_992,In_1491);
and U1920 (N_1920,N_705,N_544);
and U1921 (N_1921,In_2203,In_2087);
xor U1922 (N_1922,In_2882,In_2011);
nand U1923 (N_1923,In_1500,In_623);
nand U1924 (N_1924,N_207,In_2099);
nor U1925 (N_1925,N_359,N_201);
xnor U1926 (N_1926,N_839,N_39);
nor U1927 (N_1927,N_948,In_1736);
nand U1928 (N_1928,N_606,N_379);
and U1929 (N_1929,In_2353,In_2051);
xnor U1930 (N_1930,In_1546,N_959);
nor U1931 (N_1931,In_2517,N_496);
and U1932 (N_1932,N_809,N_45);
and U1933 (N_1933,N_703,N_629);
nand U1934 (N_1934,In_1269,N_126);
nor U1935 (N_1935,N_192,In_2729);
nor U1936 (N_1936,N_823,In_745);
xnor U1937 (N_1937,In_1412,N_525);
nand U1938 (N_1938,N_270,In_1038);
and U1939 (N_1939,N_687,N_535);
nand U1940 (N_1940,N_392,In_2017);
or U1941 (N_1941,N_666,In_2388);
nor U1942 (N_1942,N_412,N_665);
xnor U1943 (N_1943,N_91,N_1);
xor U1944 (N_1944,In_266,In_2352);
xnor U1945 (N_1945,In_1064,N_222);
or U1946 (N_1946,N_903,In_2406);
xor U1947 (N_1947,N_164,In_203);
nor U1948 (N_1948,In_2700,N_37);
and U1949 (N_1949,In_1009,N_322);
or U1950 (N_1950,N_714,N_457);
or U1951 (N_1951,In_2535,In_946);
xnor U1952 (N_1952,N_570,N_584);
nor U1953 (N_1953,In_2802,N_289);
nand U1954 (N_1954,In_1182,N_341);
or U1955 (N_1955,N_203,N_237);
nand U1956 (N_1956,In_103,N_501);
xor U1957 (N_1957,N_567,In_2872);
nor U1958 (N_1958,N_479,N_814);
xnor U1959 (N_1959,N_704,N_74);
nand U1960 (N_1960,In_1758,N_202);
and U1961 (N_1961,N_17,In_2142);
and U1962 (N_1962,In_422,N_940);
and U1963 (N_1963,N_637,N_738);
and U1964 (N_1964,N_536,In_369);
nor U1965 (N_1965,N_870,In_2687);
or U1966 (N_1966,In_2719,In_875);
nor U1967 (N_1967,In_1467,In_2129);
xor U1968 (N_1968,N_362,In_2404);
or U1969 (N_1969,In_2743,N_566);
xor U1970 (N_1970,N_698,In_2714);
and U1971 (N_1971,N_946,N_788);
nand U1972 (N_1972,N_463,In_1147);
nor U1973 (N_1973,In_1048,N_448);
xnor U1974 (N_1974,In_107,In_1976);
xor U1975 (N_1975,In_1824,N_390);
and U1976 (N_1976,N_211,In_1372);
nand U1977 (N_1977,N_904,N_11);
nor U1978 (N_1978,In_2656,N_373);
xor U1979 (N_1979,In_2247,In_2040);
and U1980 (N_1980,In_1270,N_836);
or U1981 (N_1981,In_1821,In_1677);
or U1982 (N_1982,N_261,In_2307);
xor U1983 (N_1983,In_1155,In_1505);
and U1984 (N_1984,N_38,In_2107);
nand U1985 (N_1985,N_677,In_1852);
and U1986 (N_1986,In_136,N_268);
nand U1987 (N_1987,In_1561,In_1654);
or U1988 (N_1988,N_840,N_782);
and U1989 (N_1989,N_467,In_1659);
nor U1990 (N_1990,N_969,N_926);
xor U1991 (N_1991,In_1304,N_574);
nor U1992 (N_1992,In_589,In_954);
or U1993 (N_1993,In_2920,In_2916);
or U1994 (N_1994,In_1319,N_9);
and U1995 (N_1995,N_550,In_1777);
nand U1996 (N_1996,In_2134,N_528);
and U1997 (N_1997,In_1091,In_287);
nand U1998 (N_1998,In_1671,In_1820);
nor U1999 (N_1999,In_2251,In_130);
nor U2000 (N_2000,N_1332,N_1036);
and U2001 (N_2001,N_1380,N_1352);
nand U2002 (N_2002,N_1438,N_1231);
or U2003 (N_2003,N_1957,N_1168);
or U2004 (N_2004,N_1888,N_1034);
and U2005 (N_2005,N_1302,N_1011);
and U2006 (N_2006,N_1092,N_1254);
nor U2007 (N_2007,N_1341,N_1785);
or U2008 (N_2008,N_1658,N_1956);
nand U2009 (N_2009,N_1441,N_1026);
nand U2010 (N_2010,N_1997,N_1021);
xor U2011 (N_2011,N_1460,N_1239);
xnor U2012 (N_2012,N_1243,N_1445);
nand U2013 (N_2013,N_1753,N_1651);
nand U2014 (N_2014,N_1631,N_1701);
nor U2015 (N_2015,N_1087,N_1019);
nor U2016 (N_2016,N_1782,N_1462);
nor U2017 (N_2017,N_1298,N_1423);
nor U2018 (N_2018,N_1867,N_1280);
and U2019 (N_2019,N_1566,N_1284);
xnor U2020 (N_2020,N_1493,N_1094);
nor U2021 (N_2021,N_1550,N_1154);
or U2022 (N_2022,N_1077,N_1327);
and U2023 (N_2023,N_1503,N_1244);
or U2024 (N_2024,N_1303,N_1073);
or U2025 (N_2025,N_1805,N_1042);
nor U2026 (N_2026,N_1252,N_1938);
nand U2027 (N_2027,N_1098,N_1202);
nor U2028 (N_2028,N_1638,N_1541);
nand U2029 (N_2029,N_1727,N_1031);
nand U2030 (N_2030,N_1806,N_1055);
or U2031 (N_2031,N_1848,N_1232);
nand U2032 (N_2032,N_1839,N_1920);
or U2033 (N_2033,N_1457,N_1353);
xnor U2034 (N_2034,N_1770,N_1320);
xnor U2035 (N_2035,N_1109,N_1816);
nor U2036 (N_2036,N_1234,N_1266);
or U2037 (N_2037,N_1945,N_1050);
xnor U2038 (N_2038,N_1212,N_1847);
or U2039 (N_2039,N_1468,N_1836);
xnor U2040 (N_2040,N_1326,N_1429);
nor U2041 (N_2041,N_1113,N_1759);
nand U2042 (N_2042,N_1758,N_1869);
nor U2043 (N_2043,N_1907,N_1110);
and U2044 (N_2044,N_1630,N_1388);
nor U2045 (N_2045,N_1790,N_1307);
and U2046 (N_2046,N_1349,N_1435);
nand U2047 (N_2047,N_1742,N_1667);
xor U2048 (N_2048,N_1518,N_1600);
or U2049 (N_2049,N_1300,N_1842);
nand U2050 (N_2050,N_1028,N_1578);
nand U2051 (N_2051,N_1768,N_1364);
nand U2052 (N_2052,N_1817,N_1103);
xnor U2053 (N_2053,N_1661,N_1875);
and U2054 (N_2054,N_1463,N_1116);
xnor U2055 (N_2055,N_1653,N_1876);
and U2056 (N_2056,N_1972,N_1629);
xnor U2057 (N_2057,N_1844,N_1704);
xor U2058 (N_2058,N_1317,N_1650);
and U2059 (N_2059,N_1616,N_1012);
nor U2060 (N_2060,N_1866,N_1372);
and U2061 (N_2061,N_1292,N_1311);
nand U2062 (N_2062,N_1481,N_1647);
nor U2063 (N_2063,N_1365,N_1201);
or U2064 (N_2064,N_1579,N_1078);
nand U2065 (N_2065,N_1652,N_1835);
xor U2066 (N_2066,N_1786,N_1967);
nand U2067 (N_2067,N_1634,N_1729);
and U2068 (N_2068,N_1676,N_1175);
or U2069 (N_2069,N_1416,N_1863);
nand U2070 (N_2070,N_1067,N_1763);
xor U2071 (N_2071,N_1619,N_1649);
and U2072 (N_2072,N_1192,N_1333);
nand U2073 (N_2073,N_1296,N_1000);
nand U2074 (N_2074,N_1209,N_1166);
nor U2075 (N_2075,N_1030,N_1282);
or U2076 (N_2076,N_1060,N_1715);
and U2077 (N_2077,N_1536,N_1556);
xor U2078 (N_2078,N_1363,N_1703);
nor U2079 (N_2079,N_1024,N_1343);
or U2080 (N_2080,N_1123,N_1889);
and U2081 (N_2081,N_1414,N_1152);
nand U2082 (N_2082,N_1127,N_1724);
or U2083 (N_2083,N_1926,N_1115);
xnor U2084 (N_2084,N_1375,N_1147);
xnor U2085 (N_2085,N_1072,N_1378);
and U2086 (N_2086,N_1480,N_1017);
or U2087 (N_2087,N_1965,N_1524);
nand U2088 (N_2088,N_1752,N_1187);
and U2089 (N_2089,N_1797,N_1559);
nor U2090 (N_2090,N_1393,N_1891);
xor U2091 (N_2091,N_1814,N_1059);
or U2092 (N_2092,N_1063,N_1639);
nor U2093 (N_2093,N_1547,N_1775);
xor U2094 (N_2094,N_1452,N_1567);
and U2095 (N_2095,N_1301,N_1846);
nand U2096 (N_2096,N_1411,N_1265);
nand U2097 (N_2097,N_1189,N_1321);
nor U2098 (N_2098,N_1963,N_1684);
and U2099 (N_2099,N_1033,N_1360);
nand U2100 (N_2100,N_1792,N_1029);
nand U2101 (N_2101,N_1689,N_1004);
nand U2102 (N_2102,N_1155,N_1940);
xor U2103 (N_2103,N_1469,N_1855);
and U2104 (N_2104,N_1722,N_1058);
nor U2105 (N_2105,N_1596,N_1121);
and U2106 (N_2106,N_1685,N_1694);
and U2107 (N_2107,N_1278,N_1404);
xor U2108 (N_2108,N_1403,N_1096);
and U2109 (N_2109,N_1543,N_1777);
nor U2110 (N_2110,N_1958,N_1377);
xnor U2111 (N_2111,N_1673,N_1114);
nand U2112 (N_2112,N_1745,N_1126);
or U2113 (N_2113,N_1497,N_1613);
nor U2114 (N_2114,N_1761,N_1879);
and U2115 (N_2115,N_1432,N_1922);
or U2116 (N_2116,N_1084,N_1794);
and U2117 (N_2117,N_1720,N_1820);
nand U2118 (N_2118,N_1819,N_1617);
and U2119 (N_2119,N_1354,N_1350);
or U2120 (N_2120,N_1522,N_1996);
or U2121 (N_2121,N_1358,N_1229);
and U2122 (N_2122,N_1734,N_1853);
xnor U2123 (N_2123,N_1670,N_1609);
nand U2124 (N_2124,N_1682,N_1486);
nand U2125 (N_2125,N_1741,N_1539);
and U2126 (N_2126,N_1335,N_1800);
nor U2127 (N_2127,N_1890,N_1191);
and U2128 (N_2128,N_1571,N_1219);
or U2129 (N_2129,N_1796,N_1978);
and U2130 (N_2130,N_1743,N_1610);
and U2131 (N_2131,N_1558,N_1367);
xor U2132 (N_2132,N_1431,N_1331);
or U2133 (N_2133,N_1157,N_1923);
nor U2134 (N_2134,N_1508,N_1046);
xor U2135 (N_2135,N_1628,N_1771);
and U2136 (N_2136,N_1659,N_1730);
nand U2137 (N_2137,N_1502,N_1944);
and U2138 (N_2138,N_1799,N_1361);
and U2139 (N_2139,N_1160,N_1971);
xor U2140 (N_2140,N_1387,N_1041);
nor U2141 (N_2141,N_1974,N_1226);
xnor U2142 (N_2142,N_1756,N_1495);
or U2143 (N_2143,N_1677,N_1340);
nand U2144 (N_2144,N_1443,N_1632);
xnor U2145 (N_2145,N_1538,N_1089);
nand U2146 (N_2146,N_1315,N_1444);
xor U2147 (N_2147,N_1336,N_1749);
or U2148 (N_2148,N_1544,N_1313);
xor U2149 (N_2149,N_1319,N_1843);
or U2150 (N_2150,N_1295,N_1583);
xor U2151 (N_2151,N_1575,N_1289);
or U2152 (N_2152,N_1990,N_1500);
nor U2153 (N_2153,N_1285,N_1691);
xnor U2154 (N_2154,N_1385,N_1405);
or U2155 (N_2155,N_1993,N_1605);
and U2156 (N_2156,N_1516,N_1344);
nand U2157 (N_2157,N_1980,N_1862);
or U2158 (N_2158,N_1263,N_1672);
nor U2159 (N_2159,N_1664,N_1376);
nand U2160 (N_2160,N_1446,N_1754);
and U2161 (N_2161,N_1069,N_1645);
nor U2162 (N_2162,N_1735,N_1662);
nor U2163 (N_2163,N_1815,N_1456);
nand U2164 (N_2164,N_1953,N_1570);
and U2165 (N_2165,N_1016,N_1125);
xnor U2166 (N_2166,N_1856,N_1563);
nor U2167 (N_2167,N_1179,N_1080);
and U2168 (N_2168,N_1347,N_1531);
xnor U2169 (N_2169,N_1648,N_1608);
or U2170 (N_2170,N_1151,N_1408);
or U2171 (N_2171,N_1789,N_1475);
nor U2172 (N_2172,N_1721,N_1573);
xor U2173 (N_2173,N_1766,N_1681);
nor U2174 (N_2174,N_1379,N_1915);
or U2175 (N_2175,N_1395,N_1081);
xor U2176 (N_2176,N_1751,N_1176);
nand U2177 (N_2177,N_1299,N_1195);
nor U2178 (N_2178,N_1666,N_1040);
xnor U2179 (N_2179,N_1178,N_1827);
and U2180 (N_2180,N_1960,N_1764);
and U2181 (N_2181,N_1611,N_1359);
nor U2182 (N_2182,N_1865,N_1808);
nand U2183 (N_2183,N_1774,N_1561);
nand U2184 (N_2184,N_1874,N_1887);
nand U2185 (N_2185,N_1895,N_1622);
xor U2186 (N_2186,N_1213,N_1618);
nor U2187 (N_2187,N_1203,N_1112);
nand U2188 (N_2188,N_1051,N_1841);
xor U2189 (N_2189,N_1227,N_1472);
nor U2190 (N_2190,N_1052,N_1400);
and U2191 (N_2191,N_1504,N_1222);
or U2192 (N_2192,N_1644,N_1106);
nand U2193 (N_2193,N_1718,N_1450);
and U2194 (N_2194,N_1975,N_1801);
xor U2195 (N_2195,N_1656,N_1117);
nor U2196 (N_2196,N_1095,N_1470);
nor U2197 (N_2197,N_1439,N_1585);
nand U2198 (N_2198,N_1695,N_1308);
xor U2199 (N_2199,N_1906,N_1018);
nor U2200 (N_2200,N_1699,N_1240);
xor U2201 (N_2201,N_1318,N_1141);
and U2202 (N_2202,N_1275,N_1220);
nand U2203 (N_2203,N_1698,N_1198);
or U2204 (N_2204,N_1269,N_1700);
xnor U2205 (N_2205,N_1068,N_1124);
nand U2206 (N_2206,N_1409,N_1725);
and U2207 (N_2207,N_1513,N_1646);
xor U2208 (N_2208,N_1809,N_1401);
xor U2209 (N_2209,N_1877,N_1357);
xor U2210 (N_2210,N_1791,N_1690);
and U2211 (N_2211,N_1419,N_1802);
or U2212 (N_2212,N_1237,N_1546);
and U2213 (N_2213,N_1428,N_1330);
nand U2214 (N_2214,N_1101,N_1054);
nor U2215 (N_2215,N_1949,N_1453);
nand U2216 (N_2216,N_1737,N_1733);
or U2217 (N_2217,N_1498,N_1161);
or U2218 (N_2218,N_1509,N_1148);
nor U2219 (N_2219,N_1027,N_1128);
xnor U2220 (N_2220,N_1070,N_1591);
nand U2221 (N_2221,N_1913,N_1860);
nor U2222 (N_2222,N_1614,N_1257);
nor U2223 (N_2223,N_1976,N_1499);
and U2224 (N_2224,N_1693,N_1119);
xnor U2225 (N_2225,N_1342,N_1982);
nand U2226 (N_2226,N_1635,N_1717);
or U2227 (N_2227,N_1402,N_1399);
nor U2228 (N_2228,N_1549,N_1134);
xor U2229 (N_2229,N_1204,N_1142);
or U2230 (N_2230,N_1858,N_1838);
nor U2231 (N_2231,N_1345,N_1390);
xnor U2232 (N_2232,N_1413,N_1182);
or U2233 (N_2233,N_1417,N_1136);
nand U2234 (N_2234,N_1324,N_1249);
nand U2235 (N_2235,N_1449,N_1467);
nand U2236 (N_2236,N_1946,N_1813);
nand U2237 (N_2237,N_1276,N_1037);
nor U2238 (N_2238,N_1803,N_1248);
or U2239 (N_2239,N_1928,N_1593);
nand U2240 (N_2240,N_1702,N_1760);
and U2241 (N_2241,N_1821,N_1436);
nand U2242 (N_2242,N_1641,N_1746);
or U2243 (N_2243,N_1952,N_1983);
or U2244 (N_2244,N_1560,N_1942);
xor U2245 (N_2245,N_1038,N_1773);
and U2246 (N_2246,N_1130,N_1748);
or U2247 (N_2247,N_1007,N_1107);
xor U2248 (N_2248,N_1845,N_1908);
nor U2249 (N_2249,N_1880,N_1137);
or U2250 (N_2250,N_1484,N_1144);
and U2251 (N_2251,N_1274,N_1747);
xor U2252 (N_2252,N_1939,N_1001);
and U2253 (N_2253,N_1097,N_1071);
and U2254 (N_2254,N_1810,N_1159);
and U2255 (N_2255,N_1933,N_1104);
nand U2256 (N_2256,N_1169,N_1830);
xor U2257 (N_2257,N_1139,N_1167);
xor U2258 (N_2258,N_1005,N_1832);
or U2259 (N_2259,N_1892,N_1837);
xnor U2260 (N_2260,N_1950,N_1165);
nor U2261 (N_2261,N_1049,N_1918);
nand U2262 (N_2262,N_1074,N_1023);
or U2263 (N_2263,N_1262,N_1206);
xor U2264 (N_2264,N_1793,N_1286);
and U2265 (N_2265,N_1769,N_1478);
xor U2266 (N_2266,N_1533,N_1440);
nand U2267 (N_2267,N_1553,N_1824);
nand U2268 (N_2268,N_1568,N_1961);
nand U2269 (N_2269,N_1643,N_1986);
and U2270 (N_2270,N_1985,N_1250);
nor U2271 (N_2271,N_1371,N_1589);
nor U2272 (N_2272,N_1921,N_1305);
nor U2273 (N_2273,N_1555,N_1464);
nor U2274 (N_2274,N_1290,N_1989);
xor U2275 (N_2275,N_1479,N_1688);
or U2276 (N_2276,N_1461,N_1323);
and U2277 (N_2277,N_1857,N_1902);
xor U2278 (N_2278,N_1995,N_1009);
nand U2279 (N_2279,N_1588,N_1164);
or U2280 (N_2280,N_1309,N_1496);
xnor U2281 (N_2281,N_1186,N_1228);
nand U2282 (N_2282,N_1412,N_1581);
and U2283 (N_2283,N_1510,N_1894);
or U2284 (N_2284,N_1466,N_1199);
nand U2285 (N_2285,N_1482,N_1437);
nand U2286 (N_2286,N_1767,N_1962);
xnor U2287 (N_2287,N_1612,N_1697);
nand U2288 (N_2288,N_1987,N_1120);
and U2289 (N_2289,N_1032,N_1013);
nor U2290 (N_2290,N_1812,N_1185);
nor U2291 (N_2291,N_1304,N_1574);
nand U2292 (N_2292,N_1929,N_1406);
xnor U2293 (N_2293,N_1897,N_1277);
nor U2294 (N_2294,N_1757,N_1245);
and U2295 (N_2295,N_1968,N_1910);
or U2296 (N_2296,N_1133,N_1473);
and U2297 (N_2297,N_1736,N_1657);
xor U2298 (N_2298,N_1716,N_1163);
xor U2299 (N_2299,N_1362,N_1256);
and U2300 (N_2300,N_1881,N_1669);
nand U2301 (N_2301,N_1200,N_1964);
nand U2302 (N_2302,N_1825,N_1369);
or U2303 (N_2303,N_1765,N_1931);
or U2304 (N_2304,N_1183,N_1233);
nor U2305 (N_2305,N_1991,N_1795);
xor U2306 (N_2306,N_1132,N_1705);
xor U2307 (N_2307,N_1093,N_1994);
nand U2308 (N_2308,N_1602,N_1580);
nand U2309 (N_2309,N_1537,N_1590);
and U2310 (N_2310,N_1607,N_1287);
nand U2311 (N_2311,N_1852,N_1065);
nor U2312 (N_2312,N_1936,N_1615);
and U2313 (N_2313,N_1692,N_1270);
nand U2314 (N_2314,N_1675,N_1138);
nand U2315 (N_2315,N_1140,N_1582);
and U2316 (N_2316,N_1346,N_1787);
nor U2317 (N_2317,N_1418,N_1595);
or U2318 (N_2318,N_1061,N_1624);
or U2319 (N_2319,N_1442,N_1850);
xnor U2320 (N_2320,N_1122,N_1655);
nand U2321 (N_2321,N_1517,N_1740);
xor U2322 (N_2322,N_1337,N_1849);
nand U2323 (N_2323,N_1731,N_1057);
xor U2324 (N_2324,N_1512,N_1210);
nor U2325 (N_2325,N_1603,N_1919);
or U2326 (N_2326,N_1325,N_1224);
or U2327 (N_2327,N_1355,N_1893);
nand U2328 (N_2328,N_1750,N_1783);
xor U2329 (N_2329,N_1709,N_1914);
nand U2330 (N_2330,N_1083,N_1514);
or U2331 (N_2331,N_1100,N_1288);
nand U2332 (N_2332,N_1045,N_1912);
nand U2333 (N_2333,N_1977,N_1314);
xor U2334 (N_2334,N_1726,N_1506);
nor U2335 (N_2335,N_1898,N_1999);
or U2336 (N_2336,N_1082,N_1927);
nor U2337 (N_2337,N_1955,N_1519);
and U2338 (N_2338,N_1811,N_1525);
and U2339 (N_2339,N_1392,N_1181);
nand U2340 (N_2340,N_1218,N_1398);
nand U2341 (N_2341,N_1410,N_1872);
xor U2342 (N_2342,N_1238,N_1934);
nor U2343 (N_2343,N_1523,N_1015);
and U2344 (N_2344,N_1434,N_1494);
xnor U2345 (N_2345,N_1642,N_1328);
nor U2346 (N_2346,N_1878,N_1663);
and U2347 (N_2347,N_1719,N_1162);
xnor U2348 (N_2348,N_1708,N_1477);
and U2349 (N_2349,N_1707,N_1242);
nor U2350 (N_2350,N_1421,N_1884);
xor U2351 (N_2351,N_1235,N_1671);
xor U2352 (N_2352,N_1772,N_1217);
and U2353 (N_2353,N_1840,N_1279);
xor U2354 (N_2354,N_1492,N_1804);
nor U2355 (N_2355,N_1966,N_1885);
or U2356 (N_2356,N_1366,N_1025);
or U2357 (N_2357,N_1306,N_1633);
nor U2358 (N_2358,N_1158,N_1370);
nand U2359 (N_2359,N_1924,N_1135);
xor U2360 (N_2360,N_1102,N_1455);
nor U2361 (N_2361,N_1778,N_1584);
nand U2362 (N_2362,N_1592,N_1348);
nor U2363 (N_2363,N_1528,N_1091);
or U2364 (N_2364,N_1828,N_1621);
nand U2365 (N_2365,N_1451,N_1941);
nor U2366 (N_2366,N_1859,N_1973);
nor U2367 (N_2367,N_1088,N_1216);
and U2368 (N_2368,N_1654,N_1214);
and U2369 (N_2369,N_1992,N_1925);
nor U2370 (N_2370,N_1900,N_1904);
and U2371 (N_2371,N_1422,N_1686);
nor U2372 (N_2372,N_1679,N_1208);
xnor U2373 (N_2373,N_1788,N_1246);
nand U2374 (N_2374,N_1535,N_1329);
and U2375 (N_2375,N_1665,N_1491);
and U2376 (N_2376,N_1540,N_1447);
nor U2377 (N_2377,N_1551,N_1826);
nand U2378 (N_2378,N_1079,N_1283);
or U2379 (N_2379,N_1002,N_1268);
and U2380 (N_2380,N_1173,N_1732);
nor U2381 (N_2381,N_1177,N_1062);
nand U2382 (N_2382,N_1394,N_1738);
or U2383 (N_2383,N_1022,N_1086);
or U2384 (N_2384,N_1930,N_1565);
or U2385 (N_2385,N_1391,N_1970);
and U2386 (N_2386,N_1822,N_1871);
nor U2387 (N_2387,N_1744,N_1594);
or U2388 (N_2388,N_1981,N_1947);
or U2389 (N_2389,N_1954,N_1064);
and U2390 (N_2390,N_1520,N_1215);
and U2391 (N_2391,N_1236,N_1886);
nor U2392 (N_2392,N_1407,N_1784);
xnor U2393 (N_2393,N_1710,N_1587);
or U2394 (N_2394,N_1674,N_1683);
and U2395 (N_2395,N_1260,N_1310);
nand U2396 (N_2396,N_1515,N_1557);
or U2397 (N_2397,N_1272,N_1818);
or U2398 (N_2398,N_1714,N_1937);
nor U2399 (N_2399,N_1448,N_1488);
nor U2400 (N_2400,N_1542,N_1979);
xnor U2401 (N_2401,N_1626,N_1196);
xnor U2402 (N_2402,N_1948,N_1014);
nand U2403 (N_2403,N_1905,N_1149);
or U2404 (N_2404,N_1831,N_1471);
and U2405 (N_2405,N_1053,N_1396);
and U2406 (N_2406,N_1577,N_1529);
nor U2407 (N_2407,N_1273,N_1338);
or U2408 (N_2408,N_1969,N_1552);
or U2409 (N_2409,N_1264,N_1131);
xor U2410 (N_2410,N_1111,N_1188);
and U2411 (N_2411,N_1984,N_1660);
xor U2412 (N_2412,N_1668,N_1056);
xnor U2413 (N_2413,N_1190,N_1230);
xor U2414 (N_2414,N_1397,N_1006);
nor U2415 (N_2415,N_1564,N_1258);
and U2416 (N_2416,N_1490,N_1424);
or U2417 (N_2417,N_1489,N_1174);
xnor U2418 (N_2418,N_1003,N_1415);
or U2419 (N_2419,N_1267,N_1225);
or U2420 (N_2420,N_1755,N_1833);
or U2421 (N_2421,N_1193,N_1293);
nor U2422 (N_2422,N_1597,N_1780);
xnor U2423 (N_2423,N_1554,N_1951);
and U2424 (N_2424,N_1075,N_1501);
nand U2425 (N_2425,N_1207,N_1076);
xor U2426 (N_2426,N_1548,N_1426);
and U2427 (N_2427,N_1382,N_1146);
nand U2428 (N_2428,N_1427,N_1854);
nand U2429 (N_2429,N_1599,N_1129);
nand U2430 (N_2430,N_1039,N_1008);
nor U2431 (N_2431,N_1623,N_1762);
nand U2432 (N_2432,N_1172,N_1728);
nor U2433 (N_2433,N_1334,N_1194);
nor U2434 (N_2434,N_1988,N_1606);
nor U2435 (N_2435,N_1458,N_1916);
xor U2436 (N_2436,N_1454,N_1459);
or U2437 (N_2437,N_1389,N_1943);
xnor U2438 (N_2438,N_1253,N_1433);
nand U2439 (N_2439,N_1776,N_1627);
and U2440 (N_2440,N_1261,N_1882);
nand U2441 (N_2441,N_1145,N_1532);
or U2442 (N_2442,N_1598,N_1779);
and U2443 (N_2443,N_1184,N_1153);
xor U2444 (N_2444,N_1247,N_1180);
nand U2445 (N_2445,N_1339,N_1197);
nand U2446 (N_2446,N_1223,N_1883);
and U2447 (N_2447,N_1823,N_1316);
xor U2448 (N_2448,N_1108,N_1620);
or U2449 (N_2449,N_1291,N_1781);
nand U2450 (N_2450,N_1739,N_1998);
and U2451 (N_2451,N_1205,N_1043);
or U2452 (N_2452,N_1118,N_1221);
nor U2453 (N_2453,N_1873,N_1271);
or U2454 (N_2454,N_1711,N_1035);
and U2455 (N_2455,N_1381,N_1047);
xor U2456 (N_2456,N_1586,N_1911);
and U2457 (N_2457,N_1099,N_1932);
or U2458 (N_2458,N_1527,N_1903);
nor U2459 (N_2459,N_1430,N_1465);
and U2460 (N_2460,N_1476,N_1281);
and U2461 (N_2461,N_1143,N_1351);
nor U2462 (N_2462,N_1294,N_1896);
or U2463 (N_2463,N_1511,N_1861);
nor U2464 (N_2464,N_1864,N_1487);
nand U2465 (N_2465,N_1526,N_1569);
and U2466 (N_2466,N_1322,N_1066);
or U2467 (N_2467,N_1105,N_1909);
nor U2468 (N_2468,N_1572,N_1713);
and U2469 (N_2469,N_1259,N_1251);
nor U2470 (N_2470,N_1425,N_1297);
or U2471 (N_2471,N_1712,N_1150);
nand U2472 (N_2472,N_1534,N_1383);
nand U2473 (N_2473,N_1474,N_1680);
or U2474 (N_2474,N_1851,N_1899);
or U2475 (N_2475,N_1386,N_1637);
and U2476 (N_2476,N_1829,N_1687);
nor U2477 (N_2477,N_1834,N_1241);
xor U2478 (N_2478,N_1601,N_1483);
or U2479 (N_2479,N_1798,N_1640);
nor U2480 (N_2480,N_1485,N_1696);
and U2481 (N_2481,N_1090,N_1521);
nor U2482 (N_2482,N_1678,N_1870);
xnor U2483 (N_2483,N_1010,N_1507);
or U2484 (N_2484,N_1625,N_1356);
xnor U2485 (N_2485,N_1505,N_1807);
nor U2486 (N_2486,N_1020,N_1706);
and U2487 (N_2487,N_1384,N_1935);
and U2488 (N_2488,N_1211,N_1171);
nor U2489 (N_2489,N_1530,N_1255);
nand U2490 (N_2490,N_1959,N_1901);
nor U2491 (N_2491,N_1545,N_1636);
nand U2492 (N_2492,N_1044,N_1048);
and U2493 (N_2493,N_1374,N_1170);
nor U2494 (N_2494,N_1723,N_1604);
and U2495 (N_2495,N_1156,N_1373);
nor U2496 (N_2496,N_1368,N_1562);
and U2497 (N_2497,N_1085,N_1420);
xor U2498 (N_2498,N_1576,N_1868);
and U2499 (N_2499,N_1917,N_1312);
xnor U2500 (N_2500,N_1907,N_1643);
nor U2501 (N_2501,N_1668,N_1988);
or U2502 (N_2502,N_1375,N_1053);
nor U2503 (N_2503,N_1940,N_1288);
xnor U2504 (N_2504,N_1588,N_1985);
nor U2505 (N_2505,N_1133,N_1775);
and U2506 (N_2506,N_1942,N_1012);
or U2507 (N_2507,N_1810,N_1859);
nand U2508 (N_2508,N_1802,N_1098);
xnor U2509 (N_2509,N_1627,N_1176);
or U2510 (N_2510,N_1627,N_1835);
or U2511 (N_2511,N_1721,N_1827);
nor U2512 (N_2512,N_1797,N_1057);
nor U2513 (N_2513,N_1614,N_1010);
xor U2514 (N_2514,N_1986,N_1956);
nand U2515 (N_2515,N_1388,N_1464);
or U2516 (N_2516,N_1143,N_1909);
xnor U2517 (N_2517,N_1494,N_1945);
xnor U2518 (N_2518,N_1591,N_1652);
and U2519 (N_2519,N_1897,N_1975);
nor U2520 (N_2520,N_1879,N_1597);
or U2521 (N_2521,N_1624,N_1085);
nor U2522 (N_2522,N_1047,N_1897);
xnor U2523 (N_2523,N_1705,N_1031);
and U2524 (N_2524,N_1664,N_1286);
or U2525 (N_2525,N_1671,N_1986);
and U2526 (N_2526,N_1313,N_1336);
and U2527 (N_2527,N_1826,N_1642);
or U2528 (N_2528,N_1151,N_1161);
xnor U2529 (N_2529,N_1647,N_1091);
nand U2530 (N_2530,N_1150,N_1781);
and U2531 (N_2531,N_1163,N_1351);
and U2532 (N_2532,N_1532,N_1629);
and U2533 (N_2533,N_1995,N_1536);
or U2534 (N_2534,N_1141,N_1662);
or U2535 (N_2535,N_1675,N_1259);
nand U2536 (N_2536,N_1712,N_1646);
nor U2537 (N_2537,N_1279,N_1334);
nand U2538 (N_2538,N_1926,N_1478);
nor U2539 (N_2539,N_1882,N_1318);
and U2540 (N_2540,N_1410,N_1205);
nor U2541 (N_2541,N_1653,N_1200);
nand U2542 (N_2542,N_1845,N_1323);
nor U2543 (N_2543,N_1658,N_1837);
nand U2544 (N_2544,N_1623,N_1138);
nand U2545 (N_2545,N_1637,N_1826);
nor U2546 (N_2546,N_1057,N_1325);
and U2547 (N_2547,N_1320,N_1172);
and U2548 (N_2548,N_1208,N_1118);
or U2549 (N_2549,N_1549,N_1386);
or U2550 (N_2550,N_1074,N_1854);
nor U2551 (N_2551,N_1406,N_1262);
nand U2552 (N_2552,N_1272,N_1509);
xnor U2553 (N_2553,N_1640,N_1985);
nor U2554 (N_2554,N_1034,N_1450);
or U2555 (N_2555,N_1925,N_1626);
nand U2556 (N_2556,N_1788,N_1883);
or U2557 (N_2557,N_1455,N_1139);
nand U2558 (N_2558,N_1665,N_1823);
or U2559 (N_2559,N_1416,N_1536);
or U2560 (N_2560,N_1927,N_1767);
nor U2561 (N_2561,N_1539,N_1795);
or U2562 (N_2562,N_1178,N_1401);
nand U2563 (N_2563,N_1048,N_1877);
nand U2564 (N_2564,N_1255,N_1624);
nor U2565 (N_2565,N_1109,N_1202);
nand U2566 (N_2566,N_1484,N_1521);
xnor U2567 (N_2567,N_1011,N_1846);
or U2568 (N_2568,N_1098,N_1998);
nor U2569 (N_2569,N_1735,N_1503);
or U2570 (N_2570,N_1672,N_1897);
xor U2571 (N_2571,N_1533,N_1669);
or U2572 (N_2572,N_1699,N_1550);
xor U2573 (N_2573,N_1532,N_1470);
nand U2574 (N_2574,N_1852,N_1364);
nor U2575 (N_2575,N_1462,N_1682);
or U2576 (N_2576,N_1838,N_1430);
nor U2577 (N_2577,N_1824,N_1567);
or U2578 (N_2578,N_1379,N_1980);
xor U2579 (N_2579,N_1376,N_1573);
nor U2580 (N_2580,N_1244,N_1016);
and U2581 (N_2581,N_1240,N_1930);
or U2582 (N_2582,N_1976,N_1784);
or U2583 (N_2583,N_1112,N_1570);
or U2584 (N_2584,N_1428,N_1389);
nand U2585 (N_2585,N_1891,N_1817);
nand U2586 (N_2586,N_1015,N_1317);
nor U2587 (N_2587,N_1255,N_1867);
and U2588 (N_2588,N_1245,N_1510);
and U2589 (N_2589,N_1541,N_1511);
nand U2590 (N_2590,N_1796,N_1923);
nand U2591 (N_2591,N_1472,N_1242);
xnor U2592 (N_2592,N_1043,N_1913);
nand U2593 (N_2593,N_1807,N_1946);
nor U2594 (N_2594,N_1202,N_1658);
nor U2595 (N_2595,N_1356,N_1305);
or U2596 (N_2596,N_1654,N_1050);
or U2597 (N_2597,N_1686,N_1007);
nor U2598 (N_2598,N_1015,N_1104);
or U2599 (N_2599,N_1335,N_1454);
nor U2600 (N_2600,N_1438,N_1021);
and U2601 (N_2601,N_1383,N_1139);
nand U2602 (N_2602,N_1026,N_1025);
or U2603 (N_2603,N_1910,N_1569);
xor U2604 (N_2604,N_1537,N_1362);
nand U2605 (N_2605,N_1257,N_1467);
or U2606 (N_2606,N_1575,N_1326);
and U2607 (N_2607,N_1292,N_1956);
nand U2608 (N_2608,N_1158,N_1160);
or U2609 (N_2609,N_1883,N_1010);
xor U2610 (N_2610,N_1095,N_1553);
or U2611 (N_2611,N_1334,N_1256);
or U2612 (N_2612,N_1970,N_1405);
or U2613 (N_2613,N_1441,N_1608);
and U2614 (N_2614,N_1309,N_1386);
nor U2615 (N_2615,N_1845,N_1467);
nor U2616 (N_2616,N_1924,N_1143);
or U2617 (N_2617,N_1537,N_1560);
nand U2618 (N_2618,N_1471,N_1414);
nor U2619 (N_2619,N_1562,N_1446);
and U2620 (N_2620,N_1627,N_1255);
or U2621 (N_2621,N_1412,N_1478);
nor U2622 (N_2622,N_1107,N_1473);
xor U2623 (N_2623,N_1145,N_1777);
xor U2624 (N_2624,N_1439,N_1976);
and U2625 (N_2625,N_1405,N_1742);
xor U2626 (N_2626,N_1955,N_1804);
xnor U2627 (N_2627,N_1472,N_1822);
xnor U2628 (N_2628,N_1080,N_1863);
xor U2629 (N_2629,N_1258,N_1680);
nor U2630 (N_2630,N_1129,N_1039);
or U2631 (N_2631,N_1650,N_1995);
nor U2632 (N_2632,N_1688,N_1462);
and U2633 (N_2633,N_1422,N_1216);
or U2634 (N_2634,N_1342,N_1143);
nor U2635 (N_2635,N_1101,N_1275);
and U2636 (N_2636,N_1538,N_1858);
nor U2637 (N_2637,N_1310,N_1430);
nand U2638 (N_2638,N_1018,N_1311);
or U2639 (N_2639,N_1843,N_1620);
and U2640 (N_2640,N_1804,N_1730);
xor U2641 (N_2641,N_1694,N_1722);
or U2642 (N_2642,N_1239,N_1213);
and U2643 (N_2643,N_1554,N_1406);
nor U2644 (N_2644,N_1086,N_1710);
and U2645 (N_2645,N_1576,N_1982);
or U2646 (N_2646,N_1125,N_1833);
xnor U2647 (N_2647,N_1900,N_1477);
nor U2648 (N_2648,N_1798,N_1534);
xnor U2649 (N_2649,N_1665,N_1536);
or U2650 (N_2650,N_1486,N_1154);
or U2651 (N_2651,N_1267,N_1867);
nor U2652 (N_2652,N_1800,N_1115);
and U2653 (N_2653,N_1973,N_1789);
nor U2654 (N_2654,N_1678,N_1686);
nand U2655 (N_2655,N_1328,N_1715);
or U2656 (N_2656,N_1439,N_1616);
or U2657 (N_2657,N_1418,N_1293);
and U2658 (N_2658,N_1562,N_1570);
and U2659 (N_2659,N_1474,N_1872);
xnor U2660 (N_2660,N_1289,N_1581);
nor U2661 (N_2661,N_1066,N_1958);
nand U2662 (N_2662,N_1339,N_1183);
nor U2663 (N_2663,N_1273,N_1584);
and U2664 (N_2664,N_1496,N_1951);
and U2665 (N_2665,N_1447,N_1272);
or U2666 (N_2666,N_1779,N_1515);
nor U2667 (N_2667,N_1920,N_1962);
nand U2668 (N_2668,N_1077,N_1217);
nor U2669 (N_2669,N_1451,N_1632);
and U2670 (N_2670,N_1299,N_1524);
xor U2671 (N_2671,N_1749,N_1013);
or U2672 (N_2672,N_1842,N_1908);
or U2673 (N_2673,N_1145,N_1642);
nor U2674 (N_2674,N_1950,N_1648);
or U2675 (N_2675,N_1289,N_1164);
and U2676 (N_2676,N_1183,N_1582);
nor U2677 (N_2677,N_1099,N_1260);
xor U2678 (N_2678,N_1871,N_1631);
nand U2679 (N_2679,N_1185,N_1575);
or U2680 (N_2680,N_1211,N_1725);
xnor U2681 (N_2681,N_1886,N_1709);
or U2682 (N_2682,N_1718,N_1687);
and U2683 (N_2683,N_1623,N_1897);
and U2684 (N_2684,N_1739,N_1391);
or U2685 (N_2685,N_1280,N_1851);
and U2686 (N_2686,N_1163,N_1114);
nand U2687 (N_2687,N_1758,N_1867);
and U2688 (N_2688,N_1286,N_1121);
xnor U2689 (N_2689,N_1707,N_1887);
or U2690 (N_2690,N_1041,N_1915);
nor U2691 (N_2691,N_1467,N_1243);
xnor U2692 (N_2692,N_1871,N_1554);
nand U2693 (N_2693,N_1631,N_1184);
or U2694 (N_2694,N_1359,N_1229);
and U2695 (N_2695,N_1264,N_1366);
and U2696 (N_2696,N_1004,N_1724);
and U2697 (N_2697,N_1993,N_1564);
and U2698 (N_2698,N_1188,N_1673);
nand U2699 (N_2699,N_1031,N_1017);
nor U2700 (N_2700,N_1674,N_1710);
nor U2701 (N_2701,N_1002,N_1628);
xnor U2702 (N_2702,N_1053,N_1640);
or U2703 (N_2703,N_1872,N_1293);
nor U2704 (N_2704,N_1677,N_1413);
nand U2705 (N_2705,N_1028,N_1315);
and U2706 (N_2706,N_1836,N_1874);
nor U2707 (N_2707,N_1924,N_1095);
nor U2708 (N_2708,N_1060,N_1404);
nor U2709 (N_2709,N_1645,N_1071);
and U2710 (N_2710,N_1925,N_1616);
nand U2711 (N_2711,N_1768,N_1089);
nor U2712 (N_2712,N_1263,N_1426);
nand U2713 (N_2713,N_1254,N_1342);
nor U2714 (N_2714,N_1464,N_1248);
and U2715 (N_2715,N_1913,N_1440);
and U2716 (N_2716,N_1595,N_1189);
or U2717 (N_2717,N_1055,N_1881);
nor U2718 (N_2718,N_1902,N_1762);
nor U2719 (N_2719,N_1472,N_1475);
xor U2720 (N_2720,N_1788,N_1221);
or U2721 (N_2721,N_1562,N_1318);
nor U2722 (N_2722,N_1328,N_1193);
or U2723 (N_2723,N_1637,N_1447);
nand U2724 (N_2724,N_1308,N_1239);
and U2725 (N_2725,N_1933,N_1401);
nor U2726 (N_2726,N_1022,N_1795);
or U2727 (N_2727,N_1879,N_1218);
nand U2728 (N_2728,N_1133,N_1918);
nand U2729 (N_2729,N_1487,N_1369);
nand U2730 (N_2730,N_1363,N_1013);
and U2731 (N_2731,N_1183,N_1289);
xnor U2732 (N_2732,N_1068,N_1745);
nor U2733 (N_2733,N_1704,N_1295);
nor U2734 (N_2734,N_1430,N_1662);
xor U2735 (N_2735,N_1315,N_1876);
xnor U2736 (N_2736,N_1324,N_1305);
and U2737 (N_2737,N_1438,N_1736);
xor U2738 (N_2738,N_1457,N_1298);
nor U2739 (N_2739,N_1183,N_1757);
and U2740 (N_2740,N_1232,N_1104);
nor U2741 (N_2741,N_1815,N_1156);
and U2742 (N_2742,N_1080,N_1713);
nor U2743 (N_2743,N_1093,N_1194);
nor U2744 (N_2744,N_1589,N_1577);
nor U2745 (N_2745,N_1704,N_1734);
nand U2746 (N_2746,N_1692,N_1905);
xor U2747 (N_2747,N_1065,N_1798);
and U2748 (N_2748,N_1371,N_1622);
and U2749 (N_2749,N_1546,N_1084);
nor U2750 (N_2750,N_1296,N_1354);
and U2751 (N_2751,N_1138,N_1827);
nor U2752 (N_2752,N_1464,N_1905);
and U2753 (N_2753,N_1091,N_1486);
or U2754 (N_2754,N_1727,N_1287);
xnor U2755 (N_2755,N_1191,N_1361);
or U2756 (N_2756,N_1607,N_1095);
nand U2757 (N_2757,N_1676,N_1548);
and U2758 (N_2758,N_1644,N_1967);
and U2759 (N_2759,N_1067,N_1202);
xor U2760 (N_2760,N_1721,N_1279);
or U2761 (N_2761,N_1845,N_1960);
xnor U2762 (N_2762,N_1493,N_1754);
or U2763 (N_2763,N_1958,N_1592);
nor U2764 (N_2764,N_1658,N_1280);
or U2765 (N_2765,N_1110,N_1096);
or U2766 (N_2766,N_1920,N_1805);
nor U2767 (N_2767,N_1458,N_1210);
and U2768 (N_2768,N_1070,N_1192);
or U2769 (N_2769,N_1306,N_1134);
or U2770 (N_2770,N_1416,N_1356);
xnor U2771 (N_2771,N_1412,N_1148);
xor U2772 (N_2772,N_1310,N_1526);
nor U2773 (N_2773,N_1147,N_1430);
nor U2774 (N_2774,N_1383,N_1076);
xor U2775 (N_2775,N_1035,N_1171);
or U2776 (N_2776,N_1896,N_1065);
and U2777 (N_2777,N_1050,N_1144);
xnor U2778 (N_2778,N_1109,N_1866);
nor U2779 (N_2779,N_1429,N_1680);
xnor U2780 (N_2780,N_1594,N_1068);
or U2781 (N_2781,N_1163,N_1584);
and U2782 (N_2782,N_1191,N_1836);
or U2783 (N_2783,N_1724,N_1290);
xnor U2784 (N_2784,N_1857,N_1687);
nand U2785 (N_2785,N_1393,N_1575);
or U2786 (N_2786,N_1138,N_1658);
or U2787 (N_2787,N_1738,N_1756);
nor U2788 (N_2788,N_1285,N_1075);
or U2789 (N_2789,N_1447,N_1584);
and U2790 (N_2790,N_1868,N_1682);
nor U2791 (N_2791,N_1003,N_1383);
xnor U2792 (N_2792,N_1525,N_1258);
xor U2793 (N_2793,N_1431,N_1403);
nor U2794 (N_2794,N_1969,N_1850);
nand U2795 (N_2795,N_1262,N_1624);
xnor U2796 (N_2796,N_1829,N_1173);
nor U2797 (N_2797,N_1368,N_1866);
and U2798 (N_2798,N_1328,N_1781);
xor U2799 (N_2799,N_1619,N_1516);
and U2800 (N_2800,N_1352,N_1695);
nor U2801 (N_2801,N_1926,N_1261);
and U2802 (N_2802,N_1039,N_1729);
and U2803 (N_2803,N_1503,N_1480);
and U2804 (N_2804,N_1338,N_1513);
or U2805 (N_2805,N_1704,N_1152);
xor U2806 (N_2806,N_1706,N_1417);
xor U2807 (N_2807,N_1060,N_1718);
and U2808 (N_2808,N_1703,N_1455);
or U2809 (N_2809,N_1377,N_1603);
and U2810 (N_2810,N_1605,N_1603);
nor U2811 (N_2811,N_1574,N_1453);
nor U2812 (N_2812,N_1910,N_1943);
xnor U2813 (N_2813,N_1860,N_1179);
and U2814 (N_2814,N_1303,N_1208);
nand U2815 (N_2815,N_1656,N_1407);
and U2816 (N_2816,N_1456,N_1102);
and U2817 (N_2817,N_1487,N_1245);
nor U2818 (N_2818,N_1329,N_1092);
or U2819 (N_2819,N_1959,N_1985);
and U2820 (N_2820,N_1522,N_1588);
or U2821 (N_2821,N_1243,N_1570);
and U2822 (N_2822,N_1597,N_1761);
and U2823 (N_2823,N_1329,N_1428);
or U2824 (N_2824,N_1023,N_1148);
and U2825 (N_2825,N_1891,N_1087);
xnor U2826 (N_2826,N_1265,N_1642);
or U2827 (N_2827,N_1250,N_1634);
nor U2828 (N_2828,N_1582,N_1508);
nand U2829 (N_2829,N_1898,N_1841);
or U2830 (N_2830,N_1896,N_1118);
and U2831 (N_2831,N_1226,N_1048);
nand U2832 (N_2832,N_1450,N_1929);
or U2833 (N_2833,N_1656,N_1076);
xor U2834 (N_2834,N_1150,N_1399);
xnor U2835 (N_2835,N_1087,N_1875);
xor U2836 (N_2836,N_1886,N_1984);
or U2837 (N_2837,N_1356,N_1865);
xor U2838 (N_2838,N_1992,N_1285);
nor U2839 (N_2839,N_1999,N_1831);
xor U2840 (N_2840,N_1383,N_1145);
and U2841 (N_2841,N_1672,N_1681);
and U2842 (N_2842,N_1892,N_1987);
nor U2843 (N_2843,N_1283,N_1499);
and U2844 (N_2844,N_1394,N_1390);
nand U2845 (N_2845,N_1258,N_1708);
and U2846 (N_2846,N_1151,N_1038);
and U2847 (N_2847,N_1565,N_1977);
or U2848 (N_2848,N_1025,N_1672);
or U2849 (N_2849,N_1336,N_1159);
and U2850 (N_2850,N_1229,N_1951);
nor U2851 (N_2851,N_1407,N_1570);
xnor U2852 (N_2852,N_1285,N_1150);
xor U2853 (N_2853,N_1222,N_1420);
nand U2854 (N_2854,N_1557,N_1233);
and U2855 (N_2855,N_1134,N_1529);
and U2856 (N_2856,N_1750,N_1422);
and U2857 (N_2857,N_1737,N_1966);
xor U2858 (N_2858,N_1003,N_1099);
xor U2859 (N_2859,N_1167,N_1731);
or U2860 (N_2860,N_1637,N_1282);
or U2861 (N_2861,N_1445,N_1833);
xnor U2862 (N_2862,N_1761,N_1823);
xor U2863 (N_2863,N_1588,N_1406);
and U2864 (N_2864,N_1334,N_1039);
and U2865 (N_2865,N_1436,N_1303);
nand U2866 (N_2866,N_1370,N_1808);
and U2867 (N_2867,N_1367,N_1303);
or U2868 (N_2868,N_1684,N_1104);
or U2869 (N_2869,N_1397,N_1704);
nor U2870 (N_2870,N_1250,N_1471);
nor U2871 (N_2871,N_1407,N_1832);
and U2872 (N_2872,N_1670,N_1534);
nor U2873 (N_2873,N_1690,N_1650);
or U2874 (N_2874,N_1895,N_1005);
xor U2875 (N_2875,N_1363,N_1588);
nand U2876 (N_2876,N_1568,N_1557);
nand U2877 (N_2877,N_1112,N_1038);
or U2878 (N_2878,N_1794,N_1847);
nor U2879 (N_2879,N_1166,N_1280);
nand U2880 (N_2880,N_1037,N_1382);
nor U2881 (N_2881,N_1811,N_1960);
or U2882 (N_2882,N_1903,N_1535);
nor U2883 (N_2883,N_1740,N_1643);
xor U2884 (N_2884,N_1634,N_1484);
nor U2885 (N_2885,N_1960,N_1995);
or U2886 (N_2886,N_1852,N_1695);
nand U2887 (N_2887,N_1111,N_1230);
xnor U2888 (N_2888,N_1439,N_1796);
nand U2889 (N_2889,N_1149,N_1735);
and U2890 (N_2890,N_1800,N_1170);
nand U2891 (N_2891,N_1066,N_1591);
nand U2892 (N_2892,N_1087,N_1101);
or U2893 (N_2893,N_1977,N_1087);
and U2894 (N_2894,N_1374,N_1900);
or U2895 (N_2895,N_1162,N_1737);
and U2896 (N_2896,N_1763,N_1180);
xnor U2897 (N_2897,N_1591,N_1087);
nand U2898 (N_2898,N_1333,N_1076);
nor U2899 (N_2899,N_1304,N_1079);
nand U2900 (N_2900,N_1886,N_1041);
or U2901 (N_2901,N_1939,N_1526);
nand U2902 (N_2902,N_1687,N_1196);
and U2903 (N_2903,N_1796,N_1093);
and U2904 (N_2904,N_1701,N_1642);
nor U2905 (N_2905,N_1666,N_1502);
nand U2906 (N_2906,N_1247,N_1582);
and U2907 (N_2907,N_1076,N_1148);
or U2908 (N_2908,N_1395,N_1195);
nor U2909 (N_2909,N_1094,N_1419);
or U2910 (N_2910,N_1803,N_1114);
xnor U2911 (N_2911,N_1772,N_1824);
and U2912 (N_2912,N_1603,N_1150);
nand U2913 (N_2913,N_1381,N_1603);
and U2914 (N_2914,N_1401,N_1292);
xor U2915 (N_2915,N_1890,N_1979);
nor U2916 (N_2916,N_1023,N_1830);
xor U2917 (N_2917,N_1380,N_1763);
and U2918 (N_2918,N_1731,N_1502);
or U2919 (N_2919,N_1521,N_1625);
or U2920 (N_2920,N_1593,N_1256);
xnor U2921 (N_2921,N_1979,N_1158);
nand U2922 (N_2922,N_1120,N_1249);
nor U2923 (N_2923,N_1446,N_1280);
nor U2924 (N_2924,N_1986,N_1796);
and U2925 (N_2925,N_1977,N_1912);
xor U2926 (N_2926,N_1188,N_1372);
xor U2927 (N_2927,N_1004,N_1408);
or U2928 (N_2928,N_1282,N_1909);
and U2929 (N_2929,N_1649,N_1117);
and U2930 (N_2930,N_1992,N_1296);
or U2931 (N_2931,N_1318,N_1843);
and U2932 (N_2932,N_1457,N_1921);
or U2933 (N_2933,N_1753,N_1051);
and U2934 (N_2934,N_1684,N_1608);
nand U2935 (N_2935,N_1331,N_1429);
nor U2936 (N_2936,N_1210,N_1442);
nor U2937 (N_2937,N_1854,N_1586);
or U2938 (N_2938,N_1940,N_1315);
or U2939 (N_2939,N_1452,N_1247);
xor U2940 (N_2940,N_1283,N_1235);
and U2941 (N_2941,N_1730,N_1901);
and U2942 (N_2942,N_1576,N_1748);
nand U2943 (N_2943,N_1212,N_1999);
and U2944 (N_2944,N_1303,N_1336);
xnor U2945 (N_2945,N_1207,N_1730);
nand U2946 (N_2946,N_1417,N_1894);
and U2947 (N_2947,N_1304,N_1146);
xnor U2948 (N_2948,N_1759,N_1389);
xnor U2949 (N_2949,N_1836,N_1063);
or U2950 (N_2950,N_1342,N_1766);
or U2951 (N_2951,N_1781,N_1835);
and U2952 (N_2952,N_1917,N_1055);
and U2953 (N_2953,N_1869,N_1434);
and U2954 (N_2954,N_1315,N_1268);
and U2955 (N_2955,N_1174,N_1620);
nand U2956 (N_2956,N_1387,N_1184);
and U2957 (N_2957,N_1183,N_1820);
nand U2958 (N_2958,N_1075,N_1613);
xnor U2959 (N_2959,N_1203,N_1317);
or U2960 (N_2960,N_1632,N_1172);
xnor U2961 (N_2961,N_1349,N_1664);
or U2962 (N_2962,N_1195,N_1079);
and U2963 (N_2963,N_1270,N_1783);
xor U2964 (N_2964,N_1382,N_1579);
and U2965 (N_2965,N_1406,N_1819);
nor U2966 (N_2966,N_1083,N_1286);
nand U2967 (N_2967,N_1837,N_1825);
or U2968 (N_2968,N_1542,N_1836);
and U2969 (N_2969,N_1095,N_1679);
nor U2970 (N_2970,N_1623,N_1598);
nand U2971 (N_2971,N_1175,N_1063);
nor U2972 (N_2972,N_1098,N_1059);
nand U2973 (N_2973,N_1968,N_1655);
nand U2974 (N_2974,N_1840,N_1548);
and U2975 (N_2975,N_1694,N_1347);
and U2976 (N_2976,N_1551,N_1454);
and U2977 (N_2977,N_1999,N_1778);
and U2978 (N_2978,N_1956,N_1608);
xor U2979 (N_2979,N_1072,N_1532);
xor U2980 (N_2980,N_1830,N_1380);
and U2981 (N_2981,N_1011,N_1650);
nor U2982 (N_2982,N_1952,N_1647);
nor U2983 (N_2983,N_1323,N_1646);
and U2984 (N_2984,N_1485,N_1876);
and U2985 (N_2985,N_1066,N_1094);
nor U2986 (N_2986,N_1565,N_1805);
nor U2987 (N_2987,N_1021,N_1001);
nor U2988 (N_2988,N_1866,N_1103);
nor U2989 (N_2989,N_1145,N_1172);
or U2990 (N_2990,N_1055,N_1435);
nand U2991 (N_2991,N_1617,N_1511);
xnor U2992 (N_2992,N_1796,N_1517);
or U2993 (N_2993,N_1490,N_1150);
nand U2994 (N_2994,N_1754,N_1684);
nor U2995 (N_2995,N_1116,N_1916);
xnor U2996 (N_2996,N_1855,N_1417);
or U2997 (N_2997,N_1831,N_1569);
nor U2998 (N_2998,N_1421,N_1370);
nor U2999 (N_2999,N_1530,N_1762);
and U3000 (N_3000,N_2236,N_2461);
nand U3001 (N_3001,N_2128,N_2765);
nor U3002 (N_3002,N_2961,N_2436);
nand U3003 (N_3003,N_2039,N_2673);
nor U3004 (N_3004,N_2893,N_2248);
nand U3005 (N_3005,N_2363,N_2044);
nor U3006 (N_3006,N_2817,N_2570);
xor U3007 (N_3007,N_2987,N_2109);
and U3008 (N_3008,N_2352,N_2024);
nor U3009 (N_3009,N_2212,N_2845);
xor U3010 (N_3010,N_2833,N_2130);
or U3011 (N_3011,N_2976,N_2922);
nand U3012 (N_3012,N_2628,N_2739);
and U3013 (N_3013,N_2054,N_2207);
nand U3014 (N_3014,N_2177,N_2233);
xor U3015 (N_3015,N_2907,N_2521);
and U3016 (N_3016,N_2832,N_2558);
nand U3017 (N_3017,N_2600,N_2557);
xor U3018 (N_3018,N_2362,N_2438);
nand U3019 (N_3019,N_2528,N_2936);
xor U3020 (N_3020,N_2366,N_2573);
and U3021 (N_3021,N_2389,N_2283);
nor U3022 (N_3022,N_2234,N_2806);
nor U3023 (N_3023,N_2970,N_2382);
nand U3024 (N_3024,N_2854,N_2912);
nand U3025 (N_3025,N_2771,N_2019);
or U3026 (N_3026,N_2306,N_2149);
and U3027 (N_3027,N_2471,N_2873);
and U3028 (N_3028,N_2549,N_2770);
or U3029 (N_3029,N_2729,N_2105);
nor U3030 (N_3030,N_2371,N_2339);
and U3031 (N_3031,N_2006,N_2899);
and U3032 (N_3032,N_2435,N_2501);
xor U3033 (N_3033,N_2538,N_2626);
or U3034 (N_3034,N_2975,N_2107);
and U3035 (N_3035,N_2284,N_2768);
and U3036 (N_3036,N_2175,N_2955);
and U3037 (N_3037,N_2195,N_2048);
and U3038 (N_3038,N_2431,N_2217);
and U3039 (N_3039,N_2685,N_2712);
xor U3040 (N_3040,N_2202,N_2446);
nand U3041 (N_3041,N_2201,N_2088);
nand U3042 (N_3042,N_2657,N_2527);
nor U3043 (N_3043,N_2507,N_2848);
and U3044 (N_3044,N_2047,N_2835);
xor U3045 (N_3045,N_2933,N_2082);
nor U3046 (N_3046,N_2399,N_2273);
xnor U3047 (N_3047,N_2882,N_2486);
or U3048 (N_3048,N_2514,N_2485);
or U3049 (N_3049,N_2708,N_2827);
and U3050 (N_3050,N_2281,N_2151);
xor U3051 (N_3051,N_2780,N_2225);
nand U3052 (N_3052,N_2309,N_2153);
and U3053 (N_3053,N_2784,N_2635);
or U3054 (N_3054,N_2464,N_2322);
xor U3055 (N_3055,N_2404,N_2110);
and U3056 (N_3056,N_2851,N_2290);
nand U3057 (N_3057,N_2150,N_2026);
xor U3058 (N_3058,N_2740,N_2974);
xnor U3059 (N_3059,N_2748,N_2444);
and U3060 (N_3060,N_2682,N_2778);
or U3061 (N_3061,N_2226,N_2255);
xnor U3062 (N_3062,N_2242,N_2148);
xor U3063 (N_3063,N_2169,N_2658);
xor U3064 (N_3064,N_2895,N_2477);
nand U3065 (N_3065,N_2012,N_2689);
or U3066 (N_3066,N_2332,N_2228);
xor U3067 (N_3067,N_2119,N_2440);
nand U3068 (N_3068,N_2341,N_2564);
and U3069 (N_3069,N_2938,N_2167);
xor U3070 (N_3070,N_2286,N_2075);
xor U3071 (N_3071,N_2943,N_2911);
or U3072 (N_3072,N_2610,N_2822);
nor U3073 (N_3073,N_2831,N_2287);
nor U3074 (N_3074,N_2634,N_2468);
or U3075 (N_3075,N_2519,N_2947);
nor U3076 (N_3076,N_2040,N_2121);
nand U3077 (N_3077,N_2914,N_2072);
or U3078 (N_3078,N_2840,N_2722);
or U3079 (N_3079,N_2801,N_2454);
xnor U3080 (N_3080,N_2193,N_2419);
or U3081 (N_3081,N_2256,N_2918);
nand U3082 (N_3082,N_2750,N_2709);
nor U3083 (N_3083,N_2788,N_2354);
and U3084 (N_3084,N_2125,N_2876);
nand U3085 (N_3085,N_2434,N_2991);
nor U3086 (N_3086,N_2596,N_2022);
and U3087 (N_3087,N_2523,N_2364);
or U3088 (N_3088,N_2586,N_2651);
or U3089 (N_3089,N_2241,N_2483);
and U3090 (N_3090,N_2926,N_2868);
nor U3091 (N_3091,N_2578,N_2714);
xor U3092 (N_3092,N_2033,N_2409);
nand U3093 (N_3093,N_2526,N_2099);
and U3094 (N_3094,N_2412,N_2944);
nand U3095 (N_3095,N_2805,N_2867);
nor U3096 (N_3096,N_2551,N_2159);
or U3097 (N_3097,N_2157,N_2797);
or U3098 (N_3098,N_2553,N_2580);
and U3099 (N_3099,N_2718,N_2698);
or U3100 (N_3100,N_2945,N_2927);
nand U3101 (N_3101,N_2649,N_2257);
xor U3102 (N_3102,N_2762,N_2751);
nand U3103 (N_3103,N_2411,N_2396);
nand U3104 (N_3104,N_2823,N_2502);
or U3105 (N_3105,N_2869,N_2631);
nand U3106 (N_3106,N_2036,N_2213);
or U3107 (N_3107,N_2552,N_2803);
xor U3108 (N_3108,N_2422,N_2087);
xnor U3109 (N_3109,N_2081,N_2065);
xnor U3110 (N_3110,N_2323,N_2267);
nor U3111 (N_3111,N_2903,N_2491);
or U3112 (N_3112,N_2998,N_2999);
and U3113 (N_3113,N_2730,N_2497);
xor U3114 (N_3114,N_2367,N_2155);
nor U3115 (N_3115,N_2588,N_2016);
xor U3116 (N_3116,N_2478,N_2798);
or U3117 (N_3117,N_2102,N_2819);
nand U3118 (N_3118,N_2333,N_2214);
or U3119 (N_3119,N_2813,N_2078);
and U3120 (N_3120,N_2124,N_2014);
xor U3121 (N_3121,N_2162,N_2624);
nor U3122 (N_3122,N_2031,N_2381);
nor U3123 (N_3123,N_2199,N_2518);
nor U3124 (N_3124,N_2152,N_2074);
and U3125 (N_3125,N_2963,N_2802);
xor U3126 (N_3126,N_2327,N_2437);
xor U3127 (N_3127,N_2661,N_2258);
or U3128 (N_3128,N_2968,N_2053);
nand U3129 (N_3129,N_2244,N_2344);
nand U3130 (N_3130,N_2546,N_2433);
and U3131 (N_3131,N_2697,N_2844);
or U3132 (N_3132,N_2052,N_2539);
and U3133 (N_3133,N_2206,N_2316);
xnor U3134 (N_3134,N_2305,N_2189);
and U3135 (N_3135,N_2993,N_2337);
nor U3136 (N_3136,N_2676,N_2317);
and U3137 (N_3137,N_2475,N_2448);
or U3138 (N_3138,N_2632,N_2308);
nand U3139 (N_3139,N_2852,N_2766);
nor U3140 (N_3140,N_2706,N_2465);
nand U3141 (N_3141,N_2278,N_2856);
xnor U3142 (N_3142,N_2917,N_2935);
nand U3143 (N_3143,N_2745,N_2205);
or U3144 (N_3144,N_2674,N_2196);
xor U3145 (N_3145,N_2937,N_2656);
nand U3146 (N_3146,N_2544,N_2406);
or U3147 (N_3147,N_2601,N_2513);
nor U3148 (N_3148,N_2277,N_2408);
xor U3149 (N_3149,N_2321,N_2293);
xnor U3150 (N_3150,N_2260,N_2881);
nor U3151 (N_3151,N_2505,N_2240);
or U3152 (N_3152,N_2744,N_2599);
and U3153 (N_3153,N_2545,N_2146);
nand U3154 (N_3154,N_2210,N_2025);
or U3155 (N_3155,N_2787,N_2187);
and U3156 (N_3156,N_2776,N_2630);
nor U3157 (N_3157,N_2660,N_2007);
or U3158 (N_3158,N_2458,N_2716);
and U3159 (N_3159,N_2830,N_2418);
nand U3160 (N_3160,N_2427,N_2166);
nand U3161 (N_3161,N_2170,N_2400);
and U3162 (N_3162,N_2394,N_2401);
nand U3163 (N_3163,N_2948,N_2536);
nor U3164 (N_3164,N_2862,N_2295);
and U3165 (N_3165,N_2073,N_2351);
xor U3166 (N_3166,N_2550,N_2191);
nor U3167 (N_3167,N_2463,N_2220);
nor U3168 (N_3168,N_2731,N_2097);
or U3169 (N_3169,N_2183,N_2350);
xnor U3170 (N_3170,N_2828,N_2804);
xnor U3171 (N_3171,N_2772,N_2068);
and U3172 (N_3172,N_2061,N_2038);
nand U3173 (N_3173,N_2837,N_2756);
nor U3174 (N_3174,N_2836,N_2253);
xnor U3175 (N_3175,N_2481,N_2415);
nor U3176 (N_3176,N_2111,N_2931);
nand U3177 (N_3177,N_2930,N_2967);
xnor U3178 (N_3178,N_2541,N_2118);
nand U3179 (N_3179,N_2496,N_2623);
xnor U3180 (N_3180,N_2356,N_2884);
or U3181 (N_3181,N_2728,N_2958);
or U3182 (N_3182,N_2194,N_2878);
or U3183 (N_3183,N_2603,N_2383);
xnor U3184 (N_3184,N_2665,N_2636);
and U3185 (N_3185,N_2942,N_2793);
xnor U3186 (N_3186,N_2964,N_2959);
and U3187 (N_3187,N_2164,N_2678);
or U3188 (N_3188,N_2372,N_2488);
nand U3189 (N_3189,N_2227,N_2940);
nor U3190 (N_3190,N_2269,N_2981);
nand U3191 (N_3191,N_2452,N_2185);
xor U3192 (N_3192,N_2923,N_2161);
xor U3193 (N_3193,N_2897,N_2530);
nand U3194 (N_3194,N_2621,N_2863);
or U3195 (N_3195,N_2299,N_2971);
nand U3196 (N_3196,N_2066,N_2303);
or U3197 (N_3197,N_2037,N_2997);
nor U3198 (N_3198,N_2985,N_2849);
and U3199 (N_3199,N_2304,N_2171);
and U3200 (N_3200,N_2494,N_2272);
nor U3201 (N_3201,N_2059,N_2575);
or U3202 (N_3202,N_2640,N_2158);
and U3203 (N_3203,N_2537,N_2055);
or U3204 (N_3204,N_2338,N_2050);
nor U3205 (N_3205,N_2983,N_2915);
xor U3206 (N_3206,N_2652,N_2686);
and U3207 (N_3207,N_2021,N_2476);
or U3208 (N_3208,N_2100,N_2223);
nor U3209 (N_3209,N_2375,N_2783);
xor U3210 (N_3210,N_2866,N_2027);
or U3211 (N_3211,N_2810,N_2353);
or U3212 (N_3212,N_2913,N_2134);
and U3213 (N_3213,N_2349,N_2275);
nor U3214 (N_3214,N_2489,N_2120);
and U3215 (N_3215,N_2637,N_2368);
xor U3216 (N_3216,N_2613,N_2173);
nor U3217 (N_3217,N_2288,N_2548);
nand U3218 (N_3218,N_2949,N_2510);
or U3219 (N_3219,N_2547,N_2492);
xor U3220 (N_3220,N_2593,N_2654);
nor U3221 (N_3221,N_2049,N_2413);
and U3222 (N_3222,N_2064,N_2147);
and U3223 (N_3223,N_2713,N_2359);
nand U3224 (N_3224,N_2901,N_2500);
nor U3225 (N_3225,N_2165,N_2174);
and U3226 (N_3226,N_2680,N_2373);
xor U3227 (N_3227,N_2872,N_2369);
nor U3228 (N_3228,N_2924,N_2785);
nor U3229 (N_3229,N_2655,N_2280);
nor U3230 (N_3230,N_2182,N_2696);
and U3231 (N_3231,N_2051,N_2300);
nor U3232 (N_3232,N_2572,N_2115);
or U3233 (N_3233,N_2487,N_2126);
nand U3234 (N_3234,N_2137,N_2160);
and U3235 (N_3235,N_2681,N_2595);
and U3236 (N_3236,N_2972,N_2957);
xor U3237 (N_3237,N_2459,N_2015);
nand U3238 (N_3238,N_2390,N_2380);
nand U3239 (N_3239,N_2141,N_2896);
xnor U3240 (N_3240,N_2960,N_2753);
xnor U3241 (N_3241,N_2178,N_2466);
xor U3242 (N_3242,N_2532,N_2484);
xnor U3243 (N_3243,N_2442,N_2509);
and U3244 (N_3244,N_2559,N_2407);
nand U3245 (N_3245,N_2057,N_2606);
or U3246 (N_3246,N_2761,N_2758);
nor U3247 (N_3247,N_2816,N_2101);
and U3248 (N_3248,N_2347,N_2041);
or U3249 (N_3249,N_2346,N_2184);
nand U3250 (N_3250,N_2297,N_2754);
xor U3251 (N_3251,N_2786,N_2017);
xor U3252 (N_3252,N_2582,N_2140);
nand U3253 (N_3253,N_2749,N_2700);
or U3254 (N_3254,N_2920,N_2113);
nand U3255 (N_3255,N_2719,N_2525);
nand U3256 (N_3256,N_2707,N_2138);
or U3257 (N_3257,N_2336,N_2473);
nand U3258 (N_3258,N_2462,N_2671);
xnor U3259 (N_3259,N_2883,N_2585);
and U3260 (N_3260,N_2988,N_2659);
nand U3261 (N_3261,N_2825,N_2398);
and U3262 (N_3262,N_2232,N_2767);
xor U3263 (N_3263,N_2704,N_2123);
nand U3264 (N_3264,N_2329,N_2200);
nand U3265 (N_3265,N_2251,N_2800);
xnor U3266 (N_3266,N_2083,N_2853);
nor U3267 (N_3267,N_2560,N_2720);
xor U3268 (N_3268,N_2916,N_2060);
nor U3269 (N_3269,N_2430,N_2643);
and U3270 (N_3270,N_2870,N_2695);
or U3271 (N_3271,N_2262,N_2004);
nand U3272 (N_3272,N_2562,N_2414);
or U3273 (N_3273,N_2604,N_2887);
nor U3274 (N_3274,N_2313,N_2977);
xor U3275 (N_3275,N_2011,N_2741);
nand U3276 (N_3276,N_2715,N_2186);
xnor U3277 (N_3277,N_2535,N_2271);
nand U3278 (N_3278,N_2348,N_2743);
and U3279 (N_3279,N_2857,N_2633);
or U3280 (N_3280,N_2799,N_2221);
nand U3281 (N_3281,N_2030,N_2132);
and U3282 (N_3282,N_2112,N_2794);
nor U3283 (N_3283,N_2245,N_2777);
and U3284 (N_3284,N_2457,N_2180);
xor U3285 (N_3285,N_2378,N_2156);
or U3286 (N_3286,N_2067,N_2646);
and U3287 (N_3287,N_2737,N_2358);
nor U3288 (N_3288,N_2190,N_2423);
or U3289 (N_3289,N_2932,N_2426);
nor U3290 (N_3290,N_2919,N_2254);
and U3291 (N_3291,N_2990,N_2385);
nor U3292 (N_3292,N_2962,N_2984);
xnor U3293 (N_3293,N_2908,N_2108);
nor U3294 (N_3294,N_2208,N_2829);
or U3295 (N_3295,N_2734,N_2480);
or U3296 (N_3296,N_2516,N_2607);
or U3297 (N_3297,N_2773,N_2117);
or U3298 (N_3298,N_2469,N_2865);
nor U3299 (N_3299,N_2668,N_2219);
nand U3300 (N_3300,N_2261,N_2973);
nand U3301 (N_3301,N_2814,N_2095);
and U3302 (N_3302,N_2769,N_2215);
or U3303 (N_3303,N_2135,N_2569);
xnor U3304 (N_3304,N_2198,N_2237);
or U3305 (N_3305,N_2216,N_2474);
and U3306 (N_3306,N_2139,N_2395);
nand U3307 (N_3307,N_2608,N_2467);
nand U3308 (N_3308,N_2080,N_2402);
or U3309 (N_3309,N_2650,N_2605);
nor U3310 (N_3310,N_2265,N_2179);
xor U3311 (N_3311,N_2954,N_2889);
or U3312 (N_3312,N_2760,N_2843);
xnor U3313 (N_3313,N_2503,N_2763);
or U3314 (N_3314,N_2925,N_2859);
xor U3315 (N_3315,N_2966,N_2328);
or U3316 (N_3316,N_2711,N_2209);
nor U3317 (N_3317,N_2203,N_2342);
or U3318 (N_3318,N_2145,N_2291);
xnor U3319 (N_3319,N_2376,N_2370);
and U3320 (N_3320,N_2946,N_2592);
or U3321 (N_3321,N_2229,N_2264);
nor U3322 (N_3322,N_2428,N_2587);
nand U3323 (N_3323,N_2302,N_2952);
or U3324 (N_3324,N_2989,N_2790);
nand U3325 (N_3325,N_2644,N_2063);
or U3326 (N_3326,N_2629,N_2020);
or U3327 (N_3327,N_2090,N_2522);
xor U3328 (N_3328,N_2114,N_2450);
nor U3329 (N_3329,N_2133,N_2591);
xor U3330 (N_3330,N_2565,N_2238);
nand U3331 (N_3331,N_2702,N_2892);
nor U3332 (N_3332,N_2648,N_2292);
xnor U3333 (N_3333,N_2638,N_2574);
xnor U3334 (N_3334,N_2838,N_2641);
and U3335 (N_3335,N_2493,N_2517);
or U3336 (N_3336,N_2443,N_2699);
or U3337 (N_3337,N_2243,N_2058);
and U3338 (N_3338,N_2276,N_2609);
or U3339 (N_3339,N_2554,N_2667);
xnor U3340 (N_3340,N_2850,N_2764);
or U3341 (N_3341,N_2757,N_2318);
nor U3342 (N_3342,N_2619,N_2086);
nor U3343 (N_3343,N_2759,N_2994);
nor U3344 (N_3344,N_2089,N_2929);
nor U3345 (N_3345,N_2733,N_2417);
and U3346 (N_3346,N_2996,N_2555);
nor U3347 (N_3347,N_2252,N_2746);
nor U3348 (N_3348,N_2334,N_2579);
nand U3349 (N_3349,N_2791,N_2250);
nor U3350 (N_3350,N_2365,N_2432);
nand U3351 (N_3351,N_2343,N_2129);
nor U3352 (N_3352,N_2211,N_2249);
and U3353 (N_3353,N_2163,N_2902);
and U3354 (N_3354,N_2687,N_2703);
xnor U3355 (N_3355,N_2028,N_2688);
and U3356 (N_3356,N_2611,N_2531);
nand U3357 (N_3357,N_2397,N_2950);
and U3358 (N_3358,N_2460,N_2421);
and U3359 (N_3359,N_2782,N_2259);
nor U3360 (N_3360,N_2692,N_2310);
xor U3361 (N_3361,N_2906,N_2499);
xor U3362 (N_3362,N_2664,N_2670);
nor U3363 (N_3363,N_2724,N_2034);
and U3364 (N_3364,N_2796,N_2294);
nor U3365 (N_3365,N_2085,N_2391);
nand U3366 (N_3366,N_2441,N_2239);
or U3367 (N_3367,N_2735,N_2439);
nor U3368 (N_3368,N_2131,N_2472);
xor U3369 (N_3369,N_2934,N_2880);
nand U3370 (N_3370,N_2969,N_2324);
nor U3371 (N_3371,N_2826,N_2820);
nand U3372 (N_3372,N_2042,N_2921);
or U3373 (N_3373,N_2824,N_2841);
xnor U3374 (N_3374,N_2742,N_2694);
xnor U3375 (N_3375,N_2197,N_2314);
xor U3376 (N_3376,N_2639,N_2357);
and U3377 (N_3377,N_2965,N_2274);
and U3378 (N_3378,N_2614,N_2515);
or U3379 (N_3379,N_2144,N_2002);
xnor U3380 (N_3380,N_2490,N_2951);
nand U3381 (N_3381,N_2077,N_2116);
nor U3382 (N_3382,N_2821,N_2622);
xnor U3383 (N_3383,N_2263,N_2192);
and U3384 (N_3384,N_2098,N_2812);
nand U3385 (N_3385,N_2268,N_2279);
nand U3386 (N_3386,N_2717,N_2556);
or U3387 (N_3387,N_2312,N_2447);
or U3388 (N_3388,N_2142,N_2616);
nand U3389 (N_3389,N_2888,N_2747);
nor U3390 (N_3390,N_2384,N_2842);
nor U3391 (N_3391,N_2508,N_2789);
or U3392 (N_3392,N_2246,N_2886);
nor U3393 (N_3393,N_2891,N_2571);
or U3394 (N_3394,N_2235,N_2705);
and U3395 (N_3395,N_2995,N_2301);
nand U3396 (N_3396,N_2340,N_2666);
and U3397 (N_3397,N_2875,N_2424);
and U3398 (N_3398,N_2176,N_2331);
nand U3399 (N_3399,N_2690,N_2379);
xnor U3400 (N_3400,N_2684,N_2589);
nand U3401 (N_3401,N_2000,N_2023);
nand U3402 (N_3402,N_2445,N_2864);
xor U3403 (N_3403,N_2001,N_2029);
xor U3404 (N_3404,N_2627,N_2524);
nand U3405 (N_3405,N_2529,N_2345);
nor U3406 (N_3406,N_2127,N_2172);
and U3407 (N_3407,N_2727,N_2834);
or U3408 (N_3408,N_2045,N_2774);
nand U3409 (N_3409,N_2307,N_2986);
xor U3410 (N_3410,N_2726,N_2043);
and U3411 (N_3411,N_2890,N_2035);
xnor U3412 (N_3412,N_2425,N_2584);
and U3413 (N_3413,N_2091,N_2298);
nand U3414 (N_3414,N_2069,N_2533);
nor U3415 (N_3415,N_2939,N_2879);
xor U3416 (N_3416,N_2871,N_2860);
xnor U3417 (N_3417,N_2900,N_2567);
nand U3418 (N_3418,N_2512,N_2079);
nor U3419 (N_3419,N_2106,N_2071);
and U3420 (N_3420,N_2779,N_2675);
and U3421 (N_3421,N_2909,N_2320);
and U3422 (N_3422,N_2602,N_2732);
nand U3423 (N_3423,N_2710,N_2795);
xor U3424 (N_3424,N_2855,N_2846);
or U3425 (N_3425,N_2617,N_2807);
xor U3426 (N_3426,N_2330,N_2861);
nor U3427 (N_3427,N_2416,N_2096);
and U3428 (N_3428,N_2581,N_2679);
or U3429 (N_3429,N_2904,N_2410);
and U3430 (N_3430,N_2858,N_2092);
nand U3431 (N_3431,N_2449,N_2540);
nand U3432 (N_3432,N_2222,N_2752);
nor U3433 (N_3433,N_2103,N_2168);
nor U3434 (N_3434,N_2388,N_2725);
xor U3435 (N_3435,N_2326,N_2693);
nor U3436 (N_3436,N_2691,N_2285);
xor U3437 (N_3437,N_2576,N_2311);
nor U3438 (N_3438,N_2122,N_2566);
xnor U3439 (N_3439,N_2360,N_2669);
nand U3440 (N_3440,N_2542,N_2289);
or U3441 (N_3441,N_2910,N_2154);
nor U3442 (N_3442,N_2266,N_2736);
and U3443 (N_3443,N_2453,N_2181);
xnor U3444 (N_3444,N_2377,N_2093);
and U3445 (N_3445,N_2577,N_2982);
or U3446 (N_3446,N_2143,N_2429);
or U3447 (N_3447,N_2393,N_2642);
xnor U3448 (N_3448,N_2009,N_2953);
and U3449 (N_3449,N_2387,N_2662);
nor U3450 (N_3450,N_2218,N_2683);
xor U3451 (N_3451,N_2296,N_2612);
nor U3452 (N_3452,N_2470,N_2520);
or U3453 (N_3453,N_2620,N_2928);
xnor U3454 (N_3454,N_2046,N_2663);
and U3455 (N_3455,N_2809,N_2003);
nor U3456 (N_3456,N_2594,N_2839);
nor U3457 (N_3457,N_2645,N_2392);
or U3458 (N_3458,N_2755,N_2498);
xor U3459 (N_3459,N_2403,N_2405);
nand U3460 (N_3460,N_2231,N_2792);
xnor U3461 (N_3461,N_2084,N_2479);
nand U3462 (N_3462,N_2808,N_2598);
or U3463 (N_3463,N_2094,N_2247);
and U3464 (N_3464,N_2018,N_2885);
and U3465 (N_3465,N_2818,N_2456);
nor U3466 (N_3466,N_2361,N_2325);
nor U3467 (N_3467,N_2319,N_2230);
nor U3468 (N_3468,N_2076,N_2590);
xnor U3469 (N_3469,N_2723,N_2877);
and U3470 (N_3470,N_2775,N_2374);
and U3471 (N_3471,N_2534,N_2224);
xnor U3472 (N_3472,N_2506,N_2781);
nor U3473 (N_3473,N_2386,N_2677);
xor U3474 (N_3474,N_2978,N_2894);
xnor U3475 (N_3475,N_2568,N_2979);
nor U3476 (N_3476,N_2315,N_2941);
nor U3477 (N_3477,N_2270,N_2482);
nor U3478 (N_3478,N_2010,N_2282);
or U3479 (N_3479,N_2451,N_2905);
nand U3480 (N_3480,N_2511,N_2561);
nor U3481 (N_3481,N_2980,N_2811);
xnor U3482 (N_3482,N_2204,N_2136);
or U3483 (N_3483,N_2355,N_2625);
nor U3484 (N_3484,N_2543,N_2062);
xnor U3485 (N_3485,N_2815,N_2032);
xor U3486 (N_3486,N_2653,N_2005);
or U3487 (N_3487,N_2597,N_2056);
or U3488 (N_3488,N_2455,N_2013);
xnor U3489 (N_3489,N_2504,N_2738);
nor U3490 (N_3490,N_2583,N_2070);
or U3491 (N_3491,N_2615,N_2874);
nor U3492 (N_3492,N_2495,N_2992);
or U3493 (N_3493,N_2898,N_2647);
xor U3494 (N_3494,N_2847,N_2701);
xor U3495 (N_3495,N_2956,N_2188);
nor U3496 (N_3496,N_2104,N_2335);
and U3497 (N_3497,N_2563,N_2672);
xnor U3498 (N_3498,N_2721,N_2420);
and U3499 (N_3499,N_2618,N_2008);
nand U3500 (N_3500,N_2907,N_2211);
nand U3501 (N_3501,N_2804,N_2745);
xor U3502 (N_3502,N_2558,N_2864);
and U3503 (N_3503,N_2152,N_2499);
nand U3504 (N_3504,N_2897,N_2509);
xor U3505 (N_3505,N_2549,N_2238);
and U3506 (N_3506,N_2581,N_2985);
xnor U3507 (N_3507,N_2188,N_2568);
xnor U3508 (N_3508,N_2175,N_2525);
and U3509 (N_3509,N_2247,N_2570);
nor U3510 (N_3510,N_2115,N_2735);
or U3511 (N_3511,N_2243,N_2628);
or U3512 (N_3512,N_2318,N_2434);
or U3513 (N_3513,N_2660,N_2107);
xor U3514 (N_3514,N_2156,N_2947);
nor U3515 (N_3515,N_2334,N_2895);
nor U3516 (N_3516,N_2354,N_2973);
nand U3517 (N_3517,N_2954,N_2874);
and U3518 (N_3518,N_2553,N_2349);
xor U3519 (N_3519,N_2900,N_2660);
xor U3520 (N_3520,N_2626,N_2679);
or U3521 (N_3521,N_2907,N_2860);
and U3522 (N_3522,N_2310,N_2873);
nand U3523 (N_3523,N_2208,N_2926);
and U3524 (N_3524,N_2287,N_2520);
or U3525 (N_3525,N_2347,N_2352);
xor U3526 (N_3526,N_2570,N_2742);
nor U3527 (N_3527,N_2722,N_2321);
nor U3528 (N_3528,N_2849,N_2515);
nor U3529 (N_3529,N_2891,N_2763);
xnor U3530 (N_3530,N_2601,N_2198);
or U3531 (N_3531,N_2324,N_2630);
and U3532 (N_3532,N_2037,N_2549);
and U3533 (N_3533,N_2671,N_2197);
nor U3534 (N_3534,N_2225,N_2127);
xnor U3535 (N_3535,N_2674,N_2292);
nor U3536 (N_3536,N_2652,N_2898);
xor U3537 (N_3537,N_2240,N_2425);
nand U3538 (N_3538,N_2198,N_2077);
nand U3539 (N_3539,N_2186,N_2751);
xor U3540 (N_3540,N_2354,N_2719);
nand U3541 (N_3541,N_2809,N_2729);
and U3542 (N_3542,N_2324,N_2089);
or U3543 (N_3543,N_2709,N_2582);
and U3544 (N_3544,N_2150,N_2586);
xor U3545 (N_3545,N_2756,N_2962);
or U3546 (N_3546,N_2960,N_2284);
xnor U3547 (N_3547,N_2868,N_2828);
nand U3548 (N_3548,N_2233,N_2746);
xnor U3549 (N_3549,N_2474,N_2554);
or U3550 (N_3550,N_2338,N_2488);
and U3551 (N_3551,N_2300,N_2148);
or U3552 (N_3552,N_2400,N_2720);
and U3553 (N_3553,N_2438,N_2655);
nor U3554 (N_3554,N_2846,N_2018);
nor U3555 (N_3555,N_2240,N_2868);
nand U3556 (N_3556,N_2063,N_2026);
nand U3557 (N_3557,N_2461,N_2478);
nand U3558 (N_3558,N_2071,N_2460);
nand U3559 (N_3559,N_2916,N_2771);
xnor U3560 (N_3560,N_2485,N_2911);
and U3561 (N_3561,N_2713,N_2848);
nand U3562 (N_3562,N_2828,N_2262);
and U3563 (N_3563,N_2564,N_2422);
nand U3564 (N_3564,N_2218,N_2299);
or U3565 (N_3565,N_2856,N_2193);
xnor U3566 (N_3566,N_2080,N_2819);
xnor U3567 (N_3567,N_2280,N_2289);
nor U3568 (N_3568,N_2367,N_2940);
or U3569 (N_3569,N_2674,N_2765);
or U3570 (N_3570,N_2743,N_2682);
xor U3571 (N_3571,N_2883,N_2875);
xnor U3572 (N_3572,N_2492,N_2077);
nor U3573 (N_3573,N_2589,N_2763);
and U3574 (N_3574,N_2360,N_2657);
or U3575 (N_3575,N_2202,N_2820);
or U3576 (N_3576,N_2063,N_2361);
nand U3577 (N_3577,N_2777,N_2900);
and U3578 (N_3578,N_2344,N_2842);
nand U3579 (N_3579,N_2967,N_2909);
or U3580 (N_3580,N_2167,N_2336);
nor U3581 (N_3581,N_2009,N_2494);
and U3582 (N_3582,N_2615,N_2672);
nor U3583 (N_3583,N_2171,N_2971);
nand U3584 (N_3584,N_2837,N_2070);
nor U3585 (N_3585,N_2876,N_2085);
nand U3586 (N_3586,N_2156,N_2278);
or U3587 (N_3587,N_2707,N_2454);
xor U3588 (N_3588,N_2651,N_2539);
nand U3589 (N_3589,N_2524,N_2345);
xor U3590 (N_3590,N_2626,N_2083);
nor U3591 (N_3591,N_2027,N_2253);
nor U3592 (N_3592,N_2258,N_2610);
nor U3593 (N_3593,N_2640,N_2319);
and U3594 (N_3594,N_2450,N_2063);
and U3595 (N_3595,N_2766,N_2772);
xor U3596 (N_3596,N_2767,N_2850);
and U3597 (N_3597,N_2089,N_2753);
nor U3598 (N_3598,N_2114,N_2930);
and U3599 (N_3599,N_2627,N_2000);
nand U3600 (N_3600,N_2094,N_2712);
nor U3601 (N_3601,N_2266,N_2641);
and U3602 (N_3602,N_2250,N_2930);
nor U3603 (N_3603,N_2784,N_2493);
nor U3604 (N_3604,N_2536,N_2164);
and U3605 (N_3605,N_2679,N_2515);
xnor U3606 (N_3606,N_2517,N_2713);
or U3607 (N_3607,N_2966,N_2574);
nand U3608 (N_3608,N_2408,N_2483);
nor U3609 (N_3609,N_2592,N_2023);
and U3610 (N_3610,N_2620,N_2637);
nor U3611 (N_3611,N_2526,N_2830);
nand U3612 (N_3612,N_2722,N_2223);
xnor U3613 (N_3613,N_2407,N_2020);
xnor U3614 (N_3614,N_2234,N_2872);
nand U3615 (N_3615,N_2981,N_2952);
nor U3616 (N_3616,N_2303,N_2764);
and U3617 (N_3617,N_2720,N_2944);
or U3618 (N_3618,N_2977,N_2125);
nor U3619 (N_3619,N_2208,N_2968);
nor U3620 (N_3620,N_2332,N_2869);
xor U3621 (N_3621,N_2875,N_2423);
and U3622 (N_3622,N_2144,N_2577);
nor U3623 (N_3623,N_2779,N_2288);
nand U3624 (N_3624,N_2353,N_2874);
nand U3625 (N_3625,N_2625,N_2368);
and U3626 (N_3626,N_2301,N_2194);
and U3627 (N_3627,N_2447,N_2010);
xnor U3628 (N_3628,N_2939,N_2807);
xnor U3629 (N_3629,N_2177,N_2529);
and U3630 (N_3630,N_2011,N_2819);
nor U3631 (N_3631,N_2927,N_2485);
and U3632 (N_3632,N_2433,N_2082);
and U3633 (N_3633,N_2749,N_2602);
or U3634 (N_3634,N_2000,N_2568);
nor U3635 (N_3635,N_2040,N_2225);
nor U3636 (N_3636,N_2055,N_2079);
nand U3637 (N_3637,N_2599,N_2342);
nor U3638 (N_3638,N_2178,N_2139);
or U3639 (N_3639,N_2687,N_2488);
nor U3640 (N_3640,N_2521,N_2308);
or U3641 (N_3641,N_2048,N_2191);
nand U3642 (N_3642,N_2388,N_2773);
nor U3643 (N_3643,N_2721,N_2959);
and U3644 (N_3644,N_2840,N_2635);
nand U3645 (N_3645,N_2747,N_2768);
nor U3646 (N_3646,N_2445,N_2653);
xor U3647 (N_3647,N_2560,N_2367);
and U3648 (N_3648,N_2719,N_2480);
nor U3649 (N_3649,N_2151,N_2610);
nor U3650 (N_3650,N_2933,N_2948);
and U3651 (N_3651,N_2243,N_2688);
nand U3652 (N_3652,N_2736,N_2129);
xor U3653 (N_3653,N_2450,N_2641);
nor U3654 (N_3654,N_2190,N_2591);
nor U3655 (N_3655,N_2587,N_2968);
nor U3656 (N_3656,N_2022,N_2450);
xor U3657 (N_3657,N_2205,N_2254);
nor U3658 (N_3658,N_2075,N_2317);
nand U3659 (N_3659,N_2713,N_2660);
nand U3660 (N_3660,N_2751,N_2943);
xnor U3661 (N_3661,N_2824,N_2495);
or U3662 (N_3662,N_2574,N_2968);
xor U3663 (N_3663,N_2549,N_2518);
xnor U3664 (N_3664,N_2168,N_2999);
and U3665 (N_3665,N_2712,N_2936);
xnor U3666 (N_3666,N_2966,N_2593);
xnor U3667 (N_3667,N_2502,N_2907);
nor U3668 (N_3668,N_2328,N_2916);
nand U3669 (N_3669,N_2017,N_2267);
and U3670 (N_3670,N_2228,N_2340);
and U3671 (N_3671,N_2739,N_2364);
nor U3672 (N_3672,N_2423,N_2352);
xor U3673 (N_3673,N_2338,N_2646);
nand U3674 (N_3674,N_2738,N_2229);
and U3675 (N_3675,N_2730,N_2792);
and U3676 (N_3676,N_2433,N_2196);
xor U3677 (N_3677,N_2649,N_2856);
or U3678 (N_3678,N_2378,N_2675);
nand U3679 (N_3679,N_2177,N_2893);
xor U3680 (N_3680,N_2762,N_2686);
nor U3681 (N_3681,N_2715,N_2880);
or U3682 (N_3682,N_2641,N_2335);
nand U3683 (N_3683,N_2155,N_2701);
nor U3684 (N_3684,N_2442,N_2642);
or U3685 (N_3685,N_2965,N_2150);
nand U3686 (N_3686,N_2267,N_2023);
xnor U3687 (N_3687,N_2503,N_2298);
and U3688 (N_3688,N_2780,N_2099);
xor U3689 (N_3689,N_2035,N_2796);
nand U3690 (N_3690,N_2458,N_2781);
and U3691 (N_3691,N_2467,N_2299);
xnor U3692 (N_3692,N_2727,N_2868);
nor U3693 (N_3693,N_2024,N_2685);
xor U3694 (N_3694,N_2713,N_2675);
and U3695 (N_3695,N_2549,N_2129);
nor U3696 (N_3696,N_2566,N_2015);
or U3697 (N_3697,N_2197,N_2144);
or U3698 (N_3698,N_2415,N_2007);
nor U3699 (N_3699,N_2660,N_2459);
nand U3700 (N_3700,N_2152,N_2226);
xor U3701 (N_3701,N_2106,N_2983);
nand U3702 (N_3702,N_2864,N_2601);
xnor U3703 (N_3703,N_2150,N_2693);
xnor U3704 (N_3704,N_2512,N_2679);
or U3705 (N_3705,N_2824,N_2678);
nand U3706 (N_3706,N_2042,N_2058);
xor U3707 (N_3707,N_2325,N_2031);
and U3708 (N_3708,N_2820,N_2274);
or U3709 (N_3709,N_2514,N_2684);
xor U3710 (N_3710,N_2989,N_2793);
or U3711 (N_3711,N_2537,N_2946);
or U3712 (N_3712,N_2374,N_2178);
and U3713 (N_3713,N_2927,N_2838);
nand U3714 (N_3714,N_2811,N_2585);
nand U3715 (N_3715,N_2404,N_2486);
nand U3716 (N_3716,N_2642,N_2110);
and U3717 (N_3717,N_2033,N_2966);
or U3718 (N_3718,N_2014,N_2165);
and U3719 (N_3719,N_2690,N_2643);
nand U3720 (N_3720,N_2814,N_2283);
nand U3721 (N_3721,N_2152,N_2405);
and U3722 (N_3722,N_2893,N_2269);
nand U3723 (N_3723,N_2002,N_2151);
nor U3724 (N_3724,N_2128,N_2902);
and U3725 (N_3725,N_2706,N_2230);
nand U3726 (N_3726,N_2911,N_2926);
xor U3727 (N_3727,N_2554,N_2524);
or U3728 (N_3728,N_2981,N_2164);
nor U3729 (N_3729,N_2198,N_2432);
or U3730 (N_3730,N_2298,N_2089);
and U3731 (N_3731,N_2409,N_2818);
xnor U3732 (N_3732,N_2816,N_2062);
xnor U3733 (N_3733,N_2254,N_2793);
and U3734 (N_3734,N_2419,N_2451);
nor U3735 (N_3735,N_2453,N_2190);
nor U3736 (N_3736,N_2797,N_2605);
nand U3737 (N_3737,N_2356,N_2801);
nand U3738 (N_3738,N_2525,N_2767);
xor U3739 (N_3739,N_2224,N_2844);
or U3740 (N_3740,N_2987,N_2013);
or U3741 (N_3741,N_2858,N_2544);
xnor U3742 (N_3742,N_2509,N_2784);
nor U3743 (N_3743,N_2824,N_2809);
nand U3744 (N_3744,N_2573,N_2281);
or U3745 (N_3745,N_2558,N_2143);
xnor U3746 (N_3746,N_2111,N_2754);
nor U3747 (N_3747,N_2047,N_2108);
and U3748 (N_3748,N_2745,N_2007);
nand U3749 (N_3749,N_2595,N_2826);
nor U3750 (N_3750,N_2809,N_2877);
nand U3751 (N_3751,N_2644,N_2675);
and U3752 (N_3752,N_2168,N_2859);
nand U3753 (N_3753,N_2738,N_2082);
xor U3754 (N_3754,N_2157,N_2971);
and U3755 (N_3755,N_2642,N_2451);
nand U3756 (N_3756,N_2749,N_2842);
nor U3757 (N_3757,N_2139,N_2885);
nand U3758 (N_3758,N_2647,N_2358);
nand U3759 (N_3759,N_2117,N_2589);
nand U3760 (N_3760,N_2210,N_2645);
nor U3761 (N_3761,N_2768,N_2864);
and U3762 (N_3762,N_2931,N_2609);
nand U3763 (N_3763,N_2445,N_2088);
nor U3764 (N_3764,N_2361,N_2749);
or U3765 (N_3765,N_2301,N_2168);
nand U3766 (N_3766,N_2322,N_2071);
nand U3767 (N_3767,N_2072,N_2127);
and U3768 (N_3768,N_2746,N_2356);
nand U3769 (N_3769,N_2784,N_2820);
nor U3770 (N_3770,N_2208,N_2091);
nor U3771 (N_3771,N_2673,N_2273);
or U3772 (N_3772,N_2303,N_2393);
nor U3773 (N_3773,N_2402,N_2622);
and U3774 (N_3774,N_2746,N_2868);
nor U3775 (N_3775,N_2813,N_2873);
or U3776 (N_3776,N_2694,N_2337);
nor U3777 (N_3777,N_2020,N_2268);
nand U3778 (N_3778,N_2144,N_2686);
xnor U3779 (N_3779,N_2617,N_2996);
and U3780 (N_3780,N_2292,N_2243);
nor U3781 (N_3781,N_2871,N_2447);
or U3782 (N_3782,N_2496,N_2813);
or U3783 (N_3783,N_2743,N_2700);
xor U3784 (N_3784,N_2387,N_2855);
nand U3785 (N_3785,N_2122,N_2435);
nand U3786 (N_3786,N_2020,N_2650);
nand U3787 (N_3787,N_2076,N_2615);
nand U3788 (N_3788,N_2074,N_2446);
or U3789 (N_3789,N_2850,N_2801);
or U3790 (N_3790,N_2107,N_2722);
or U3791 (N_3791,N_2688,N_2303);
or U3792 (N_3792,N_2689,N_2223);
and U3793 (N_3793,N_2961,N_2645);
nor U3794 (N_3794,N_2717,N_2932);
and U3795 (N_3795,N_2525,N_2481);
nor U3796 (N_3796,N_2637,N_2558);
nor U3797 (N_3797,N_2906,N_2605);
nor U3798 (N_3798,N_2980,N_2886);
and U3799 (N_3799,N_2416,N_2542);
xnor U3800 (N_3800,N_2693,N_2724);
and U3801 (N_3801,N_2188,N_2508);
nor U3802 (N_3802,N_2846,N_2513);
nor U3803 (N_3803,N_2045,N_2594);
xnor U3804 (N_3804,N_2696,N_2724);
xnor U3805 (N_3805,N_2049,N_2755);
nand U3806 (N_3806,N_2949,N_2551);
xor U3807 (N_3807,N_2272,N_2888);
nand U3808 (N_3808,N_2396,N_2483);
nand U3809 (N_3809,N_2462,N_2769);
xor U3810 (N_3810,N_2294,N_2257);
xnor U3811 (N_3811,N_2398,N_2293);
nor U3812 (N_3812,N_2415,N_2170);
and U3813 (N_3813,N_2311,N_2550);
nor U3814 (N_3814,N_2582,N_2099);
xnor U3815 (N_3815,N_2693,N_2597);
nand U3816 (N_3816,N_2538,N_2466);
nand U3817 (N_3817,N_2864,N_2213);
and U3818 (N_3818,N_2222,N_2379);
and U3819 (N_3819,N_2838,N_2729);
nor U3820 (N_3820,N_2051,N_2617);
nand U3821 (N_3821,N_2675,N_2710);
and U3822 (N_3822,N_2872,N_2244);
or U3823 (N_3823,N_2372,N_2040);
nand U3824 (N_3824,N_2222,N_2092);
xnor U3825 (N_3825,N_2036,N_2078);
nand U3826 (N_3826,N_2042,N_2611);
nand U3827 (N_3827,N_2323,N_2191);
xnor U3828 (N_3828,N_2150,N_2903);
xor U3829 (N_3829,N_2886,N_2051);
and U3830 (N_3830,N_2803,N_2515);
xor U3831 (N_3831,N_2346,N_2918);
nand U3832 (N_3832,N_2200,N_2630);
xor U3833 (N_3833,N_2338,N_2335);
nor U3834 (N_3834,N_2916,N_2971);
nand U3835 (N_3835,N_2720,N_2609);
or U3836 (N_3836,N_2061,N_2489);
nor U3837 (N_3837,N_2041,N_2403);
nor U3838 (N_3838,N_2157,N_2354);
nand U3839 (N_3839,N_2228,N_2575);
nand U3840 (N_3840,N_2514,N_2827);
xnor U3841 (N_3841,N_2219,N_2712);
nand U3842 (N_3842,N_2735,N_2826);
and U3843 (N_3843,N_2815,N_2743);
or U3844 (N_3844,N_2789,N_2214);
xor U3845 (N_3845,N_2743,N_2186);
or U3846 (N_3846,N_2328,N_2610);
and U3847 (N_3847,N_2593,N_2752);
and U3848 (N_3848,N_2431,N_2283);
nand U3849 (N_3849,N_2024,N_2110);
nor U3850 (N_3850,N_2945,N_2733);
and U3851 (N_3851,N_2673,N_2728);
nand U3852 (N_3852,N_2413,N_2730);
or U3853 (N_3853,N_2323,N_2527);
nand U3854 (N_3854,N_2087,N_2555);
nand U3855 (N_3855,N_2646,N_2337);
or U3856 (N_3856,N_2925,N_2978);
nand U3857 (N_3857,N_2711,N_2944);
or U3858 (N_3858,N_2239,N_2103);
and U3859 (N_3859,N_2970,N_2828);
and U3860 (N_3860,N_2117,N_2580);
nand U3861 (N_3861,N_2213,N_2454);
nand U3862 (N_3862,N_2800,N_2948);
nand U3863 (N_3863,N_2591,N_2794);
nor U3864 (N_3864,N_2938,N_2697);
or U3865 (N_3865,N_2226,N_2589);
xor U3866 (N_3866,N_2655,N_2124);
and U3867 (N_3867,N_2640,N_2928);
nor U3868 (N_3868,N_2580,N_2641);
xor U3869 (N_3869,N_2577,N_2568);
and U3870 (N_3870,N_2981,N_2223);
nand U3871 (N_3871,N_2312,N_2210);
and U3872 (N_3872,N_2163,N_2034);
nand U3873 (N_3873,N_2146,N_2525);
nor U3874 (N_3874,N_2979,N_2612);
or U3875 (N_3875,N_2902,N_2551);
xnor U3876 (N_3876,N_2279,N_2252);
and U3877 (N_3877,N_2015,N_2157);
or U3878 (N_3878,N_2347,N_2608);
nor U3879 (N_3879,N_2924,N_2624);
xor U3880 (N_3880,N_2715,N_2233);
and U3881 (N_3881,N_2849,N_2918);
nor U3882 (N_3882,N_2073,N_2012);
or U3883 (N_3883,N_2747,N_2750);
nor U3884 (N_3884,N_2400,N_2469);
nand U3885 (N_3885,N_2006,N_2222);
nand U3886 (N_3886,N_2145,N_2319);
nor U3887 (N_3887,N_2194,N_2282);
nand U3888 (N_3888,N_2426,N_2302);
nor U3889 (N_3889,N_2788,N_2233);
nor U3890 (N_3890,N_2992,N_2453);
and U3891 (N_3891,N_2088,N_2863);
nor U3892 (N_3892,N_2585,N_2817);
xnor U3893 (N_3893,N_2210,N_2414);
nand U3894 (N_3894,N_2423,N_2463);
and U3895 (N_3895,N_2621,N_2425);
nor U3896 (N_3896,N_2048,N_2768);
nor U3897 (N_3897,N_2020,N_2226);
or U3898 (N_3898,N_2779,N_2718);
or U3899 (N_3899,N_2957,N_2120);
and U3900 (N_3900,N_2451,N_2918);
nor U3901 (N_3901,N_2823,N_2081);
nand U3902 (N_3902,N_2667,N_2127);
nand U3903 (N_3903,N_2160,N_2775);
xor U3904 (N_3904,N_2060,N_2494);
or U3905 (N_3905,N_2688,N_2709);
nor U3906 (N_3906,N_2694,N_2211);
xor U3907 (N_3907,N_2205,N_2529);
or U3908 (N_3908,N_2973,N_2922);
xor U3909 (N_3909,N_2476,N_2645);
and U3910 (N_3910,N_2974,N_2272);
or U3911 (N_3911,N_2807,N_2530);
or U3912 (N_3912,N_2723,N_2536);
xnor U3913 (N_3913,N_2184,N_2917);
xnor U3914 (N_3914,N_2481,N_2106);
and U3915 (N_3915,N_2357,N_2315);
and U3916 (N_3916,N_2281,N_2977);
or U3917 (N_3917,N_2374,N_2590);
nand U3918 (N_3918,N_2491,N_2093);
or U3919 (N_3919,N_2958,N_2393);
nor U3920 (N_3920,N_2888,N_2077);
and U3921 (N_3921,N_2076,N_2884);
xnor U3922 (N_3922,N_2395,N_2698);
nand U3923 (N_3923,N_2185,N_2445);
xnor U3924 (N_3924,N_2406,N_2594);
nand U3925 (N_3925,N_2967,N_2493);
nand U3926 (N_3926,N_2440,N_2078);
and U3927 (N_3927,N_2025,N_2731);
or U3928 (N_3928,N_2964,N_2633);
nor U3929 (N_3929,N_2894,N_2076);
or U3930 (N_3930,N_2837,N_2132);
or U3931 (N_3931,N_2685,N_2975);
nor U3932 (N_3932,N_2557,N_2169);
nor U3933 (N_3933,N_2960,N_2318);
nor U3934 (N_3934,N_2283,N_2184);
or U3935 (N_3935,N_2300,N_2514);
and U3936 (N_3936,N_2512,N_2204);
xnor U3937 (N_3937,N_2376,N_2952);
nand U3938 (N_3938,N_2563,N_2911);
nor U3939 (N_3939,N_2601,N_2377);
nand U3940 (N_3940,N_2894,N_2330);
xor U3941 (N_3941,N_2947,N_2008);
and U3942 (N_3942,N_2203,N_2879);
nor U3943 (N_3943,N_2237,N_2347);
nand U3944 (N_3944,N_2598,N_2637);
nor U3945 (N_3945,N_2120,N_2018);
and U3946 (N_3946,N_2697,N_2292);
and U3947 (N_3947,N_2759,N_2598);
xor U3948 (N_3948,N_2501,N_2378);
or U3949 (N_3949,N_2189,N_2097);
xnor U3950 (N_3950,N_2521,N_2377);
nand U3951 (N_3951,N_2343,N_2333);
xnor U3952 (N_3952,N_2744,N_2754);
nor U3953 (N_3953,N_2854,N_2892);
nand U3954 (N_3954,N_2269,N_2587);
nor U3955 (N_3955,N_2822,N_2992);
xnor U3956 (N_3956,N_2771,N_2039);
nand U3957 (N_3957,N_2147,N_2355);
xnor U3958 (N_3958,N_2135,N_2373);
nor U3959 (N_3959,N_2998,N_2847);
nand U3960 (N_3960,N_2626,N_2104);
and U3961 (N_3961,N_2444,N_2045);
nand U3962 (N_3962,N_2486,N_2033);
and U3963 (N_3963,N_2288,N_2789);
and U3964 (N_3964,N_2560,N_2990);
or U3965 (N_3965,N_2047,N_2691);
and U3966 (N_3966,N_2914,N_2375);
xor U3967 (N_3967,N_2429,N_2439);
xnor U3968 (N_3968,N_2472,N_2696);
xnor U3969 (N_3969,N_2584,N_2310);
nor U3970 (N_3970,N_2946,N_2161);
nand U3971 (N_3971,N_2672,N_2928);
nor U3972 (N_3972,N_2930,N_2352);
nor U3973 (N_3973,N_2838,N_2630);
and U3974 (N_3974,N_2348,N_2561);
xor U3975 (N_3975,N_2228,N_2144);
nor U3976 (N_3976,N_2151,N_2595);
nor U3977 (N_3977,N_2566,N_2330);
or U3978 (N_3978,N_2067,N_2214);
nand U3979 (N_3979,N_2721,N_2221);
and U3980 (N_3980,N_2775,N_2914);
or U3981 (N_3981,N_2107,N_2592);
xnor U3982 (N_3982,N_2739,N_2367);
or U3983 (N_3983,N_2457,N_2158);
xnor U3984 (N_3984,N_2466,N_2655);
and U3985 (N_3985,N_2234,N_2911);
nor U3986 (N_3986,N_2485,N_2666);
xnor U3987 (N_3987,N_2694,N_2599);
or U3988 (N_3988,N_2677,N_2283);
nand U3989 (N_3989,N_2584,N_2416);
nand U3990 (N_3990,N_2032,N_2698);
and U3991 (N_3991,N_2811,N_2548);
nor U3992 (N_3992,N_2202,N_2814);
or U3993 (N_3993,N_2389,N_2473);
nor U3994 (N_3994,N_2236,N_2224);
or U3995 (N_3995,N_2763,N_2016);
or U3996 (N_3996,N_2629,N_2359);
nand U3997 (N_3997,N_2423,N_2971);
nand U3998 (N_3998,N_2659,N_2632);
or U3999 (N_3999,N_2533,N_2999);
nor U4000 (N_4000,N_3914,N_3981);
or U4001 (N_4001,N_3975,N_3574);
and U4002 (N_4002,N_3749,N_3158);
nor U4003 (N_4003,N_3533,N_3220);
or U4004 (N_4004,N_3420,N_3812);
nor U4005 (N_4005,N_3897,N_3400);
or U4006 (N_4006,N_3935,N_3475);
xor U4007 (N_4007,N_3004,N_3484);
or U4008 (N_4008,N_3779,N_3537);
or U4009 (N_4009,N_3281,N_3328);
xor U4010 (N_4010,N_3211,N_3860);
or U4011 (N_4011,N_3809,N_3131);
or U4012 (N_4012,N_3839,N_3028);
nand U4013 (N_4013,N_3315,N_3480);
nand U4014 (N_4014,N_3938,N_3957);
nand U4015 (N_4015,N_3843,N_3609);
nor U4016 (N_4016,N_3447,N_3815);
xor U4017 (N_4017,N_3314,N_3289);
nand U4018 (N_4018,N_3240,N_3252);
nor U4019 (N_4019,N_3947,N_3376);
xor U4020 (N_4020,N_3494,N_3448);
and U4021 (N_4021,N_3081,N_3602);
or U4022 (N_4022,N_3991,N_3715);
nor U4023 (N_4023,N_3744,N_3671);
nand U4024 (N_4024,N_3139,N_3102);
xnor U4025 (N_4025,N_3697,N_3693);
nor U4026 (N_4026,N_3623,N_3942);
or U4027 (N_4027,N_3026,N_3463);
or U4028 (N_4028,N_3764,N_3456);
or U4029 (N_4029,N_3685,N_3755);
or U4030 (N_4030,N_3753,N_3011);
nand U4031 (N_4031,N_3237,N_3769);
or U4032 (N_4032,N_3021,N_3467);
or U4033 (N_4033,N_3301,N_3505);
nand U4034 (N_4034,N_3663,N_3302);
nor U4035 (N_4035,N_3312,N_3359);
xor U4036 (N_4036,N_3976,N_3655);
and U4037 (N_4037,N_3573,N_3527);
nand U4038 (N_4038,N_3255,N_3952);
nor U4039 (N_4039,N_3726,N_3037);
nor U4040 (N_4040,N_3873,N_3611);
or U4041 (N_4041,N_3725,N_3507);
or U4042 (N_4042,N_3740,N_3300);
xor U4043 (N_4043,N_3637,N_3063);
xor U4044 (N_4044,N_3486,N_3992);
and U4045 (N_4045,N_3250,N_3479);
or U4046 (N_4046,N_3035,N_3435);
xnor U4047 (N_4047,N_3858,N_3747);
and U4048 (N_4048,N_3822,N_3694);
or U4049 (N_4049,N_3896,N_3226);
nand U4050 (N_4050,N_3859,N_3188);
or U4051 (N_4051,N_3353,N_3895);
nor U4052 (N_4052,N_3422,N_3669);
xnor U4053 (N_4053,N_3391,N_3126);
nand U4054 (N_4054,N_3737,N_3612);
or U4055 (N_4055,N_3280,N_3856);
or U4056 (N_4056,N_3535,N_3418);
nor U4057 (N_4057,N_3890,N_3136);
nand U4058 (N_4058,N_3849,N_3325);
nor U4059 (N_4059,N_3679,N_3148);
nor U4060 (N_4060,N_3181,N_3069);
or U4061 (N_4061,N_3570,N_3683);
xnor U4062 (N_4062,N_3579,N_3603);
nor U4063 (N_4063,N_3443,N_3110);
or U4064 (N_4064,N_3831,N_3078);
xnor U4065 (N_4065,N_3855,N_3660);
nor U4066 (N_4066,N_3854,N_3294);
and U4067 (N_4067,N_3378,N_3525);
xnor U4068 (N_4068,N_3877,N_3375);
nor U4069 (N_4069,N_3712,N_3218);
xnor U4070 (N_4070,N_3259,N_3304);
and U4071 (N_4071,N_3521,N_3651);
xnor U4072 (N_4072,N_3275,N_3332);
and U4073 (N_4073,N_3150,N_3423);
and U4074 (N_4074,N_3646,N_3592);
or U4075 (N_4075,N_3515,N_3163);
xor U4076 (N_4076,N_3075,N_3024);
nor U4077 (N_4077,N_3607,N_3728);
nor U4078 (N_4078,N_3532,N_3056);
and U4079 (N_4079,N_3614,N_3362);
and U4080 (N_4080,N_3310,N_3550);
nor U4081 (N_4081,N_3911,N_3575);
nand U4082 (N_4082,N_3003,N_3595);
nor U4083 (N_4083,N_3930,N_3781);
or U4084 (N_4084,N_3395,N_3306);
nor U4085 (N_4085,N_3134,N_3182);
or U4086 (N_4086,N_3885,N_3120);
or U4087 (N_4087,N_3444,N_3900);
xor U4088 (N_4088,N_3374,N_3108);
xor U4089 (N_4089,N_3841,N_3705);
and U4090 (N_4090,N_3648,N_3932);
nand U4091 (N_4091,N_3939,N_3713);
nand U4092 (N_4092,N_3179,N_3977);
nand U4093 (N_4093,N_3266,N_3330);
nor U4094 (N_4094,N_3130,N_3888);
or U4095 (N_4095,N_3452,N_3185);
and U4096 (N_4096,N_3457,N_3702);
nand U4097 (N_4097,N_3904,N_3645);
and U4098 (N_4098,N_3785,N_3690);
nand U4099 (N_4099,N_3926,N_3222);
and U4100 (N_4100,N_3650,N_3263);
nand U4101 (N_4101,N_3284,N_3924);
and U4102 (N_4102,N_3239,N_3915);
nand U4103 (N_4103,N_3441,N_3514);
or U4104 (N_4104,N_3672,N_3208);
nor U4105 (N_4105,N_3765,N_3174);
xor U4106 (N_4106,N_3707,N_3331);
and U4107 (N_4107,N_3978,N_3879);
nor U4108 (N_4108,N_3937,N_3167);
nand U4109 (N_4109,N_3544,N_3397);
and U4110 (N_4110,N_3088,N_3960);
nand U4111 (N_4111,N_3161,N_3778);
nand U4112 (N_4112,N_3929,N_3333);
nor U4113 (N_4113,N_3996,N_3619);
xnor U4114 (N_4114,N_3054,N_3903);
nor U4115 (N_4115,N_3491,N_3825);
nor U4116 (N_4116,N_3988,N_3405);
or U4117 (N_4117,N_3554,N_3621);
xor U4118 (N_4118,N_3836,N_3349);
nor U4119 (N_4119,N_3582,N_3430);
or U4120 (N_4120,N_3461,N_3807);
and U4121 (N_4121,N_3216,N_3909);
nand U4122 (N_4122,N_3551,N_3913);
xnor U4123 (N_4123,N_3197,N_3070);
or U4124 (N_4124,N_3270,N_3268);
nor U4125 (N_4125,N_3170,N_3253);
and U4126 (N_4126,N_3092,N_3502);
nand U4127 (N_4127,N_3257,N_3708);
xnor U4128 (N_4128,N_3243,N_3203);
nor U4129 (N_4129,N_3656,N_3416);
xor U4130 (N_4130,N_3561,N_3387);
nand U4131 (N_4131,N_3659,N_3576);
xor U4132 (N_4132,N_3689,N_3066);
or U4133 (N_4133,N_3555,N_3305);
xor U4134 (N_4134,N_3661,N_3547);
nand U4135 (N_4135,N_3428,N_3691);
nor U4136 (N_4136,N_3347,N_3628);
nor U4137 (N_4137,N_3407,N_3048);
or U4138 (N_4138,N_3722,N_3756);
and U4139 (N_4139,N_3084,N_3039);
and U4140 (N_4140,N_3296,N_3385);
or U4141 (N_4141,N_3251,N_3086);
xor U4142 (N_4142,N_3558,N_3354);
and U4143 (N_4143,N_3380,N_3019);
xor U4144 (N_4144,N_3064,N_3973);
nand U4145 (N_4145,N_3238,N_3953);
xor U4146 (N_4146,N_3258,N_3427);
xnor U4147 (N_4147,N_3291,N_3020);
nand U4148 (N_4148,N_3090,N_3503);
and U4149 (N_4149,N_3927,N_3687);
and U4150 (N_4150,N_3233,N_3866);
nand U4151 (N_4151,N_3723,N_3225);
or U4152 (N_4152,N_3733,N_3307);
xnor U4153 (N_4153,N_3625,N_3639);
nand U4154 (N_4154,N_3762,N_3267);
nor U4155 (N_4155,N_3453,N_3217);
nor U4156 (N_4156,N_3759,N_3598);
xor U4157 (N_4157,N_3966,N_3523);
nand U4158 (N_4158,N_3971,N_3647);
nor U4159 (N_4159,N_3122,N_3360);
or U4160 (N_4160,N_3923,N_3559);
nand U4161 (N_4161,N_3089,N_3906);
nand U4162 (N_4162,N_3548,N_3638);
xor U4163 (N_4163,N_3792,N_3945);
nor U4164 (N_4164,N_3153,N_3506);
xnor U4165 (N_4165,N_3518,N_3326);
xnor U4166 (N_4166,N_3350,N_3589);
nor U4167 (N_4167,N_3664,N_3816);
and U4168 (N_4168,N_3470,N_3413);
nor U4169 (N_4169,N_3036,N_3847);
xnor U4170 (N_4170,N_3828,N_3076);
xor U4171 (N_4171,N_3264,N_3951);
xnor U4172 (N_4172,N_3630,N_3961);
nor U4173 (N_4173,N_3254,N_3445);
or U4174 (N_4174,N_3496,N_3442);
and U4175 (N_4175,N_3803,N_3113);
and U4176 (N_4176,N_3277,N_3365);
nand U4177 (N_4177,N_3994,N_3274);
or U4178 (N_4178,N_3204,N_3772);
or U4179 (N_4179,N_3499,N_3741);
nand U4180 (N_4180,N_3152,N_3487);
or U4181 (N_4181,N_3954,N_3049);
or U4182 (N_4182,N_3686,N_3142);
nand U4183 (N_4183,N_3958,N_3517);
or U4184 (N_4184,N_3286,N_3156);
nand U4185 (N_4185,N_3339,N_3419);
or U4186 (N_4186,N_3107,N_3446);
xnor U4187 (N_4187,N_3093,N_3543);
nor U4188 (N_4188,N_3177,N_3210);
nand U4189 (N_4189,N_3027,N_3869);
nand U4190 (N_4190,N_3531,N_3613);
xor U4191 (N_4191,N_3361,N_3770);
xnor U4192 (N_4192,N_3168,N_3288);
xor U4193 (N_4193,N_3393,N_3692);
nor U4194 (N_4194,N_3348,N_3119);
nand U4195 (N_4195,N_3223,N_3029);
or U4196 (N_4196,N_3928,N_3542);
nor U4197 (N_4197,N_3944,N_3017);
nand U4198 (N_4198,N_3043,N_3450);
nand U4199 (N_4199,N_3483,N_3481);
or U4200 (N_4200,N_3103,N_3172);
nand U4201 (N_4201,N_3941,N_3053);
nor U4202 (N_4202,N_3149,N_3501);
nor U4203 (N_4203,N_3867,N_3763);
xnor U4204 (N_4204,N_3817,N_3192);
nand U4205 (N_4205,N_3768,N_3553);
or U4206 (N_4206,N_3045,N_3833);
and U4207 (N_4207,N_3701,N_3845);
or U4208 (N_4208,N_3322,N_3371);
xnor U4209 (N_4209,N_3545,N_3460);
nand U4210 (N_4210,N_3106,N_3190);
nand U4211 (N_4211,N_3754,N_3529);
nand U4212 (N_4212,N_3449,N_3287);
nor U4213 (N_4213,N_3111,N_3196);
or U4214 (N_4214,N_3317,N_3015);
and U4215 (N_4215,N_3791,N_3183);
nand U4216 (N_4216,N_3321,N_3719);
or U4217 (N_4217,N_3808,N_3074);
nor U4218 (N_4218,N_3795,N_3802);
and U4219 (N_4219,N_3214,N_3616);
and U4220 (N_4220,N_3666,N_3293);
and U4221 (N_4221,N_3716,N_3104);
and U4222 (N_4222,N_3489,N_3097);
nor U4223 (N_4223,N_3844,N_3588);
nand U4224 (N_4224,N_3830,N_3827);
nor U4225 (N_4225,N_3285,N_3567);
nor U4226 (N_4226,N_3794,N_3584);
nand U4227 (N_4227,N_3654,N_3335);
or U4228 (N_4228,N_3571,N_3215);
nor U4229 (N_4229,N_3165,N_3230);
and U4230 (N_4230,N_3451,N_3193);
nor U4231 (N_4231,N_3364,N_3382);
nor U4232 (N_4232,N_3673,N_3946);
and U4233 (N_4233,N_3058,N_3112);
and U4234 (N_4234,N_3038,N_3983);
nor U4235 (N_4235,N_3721,N_3290);
or U4236 (N_4236,N_3783,N_3644);
nor U4237 (N_4237,N_3369,N_3246);
or U4238 (N_4238,N_3917,N_3062);
nand U4239 (N_4239,N_3292,N_3889);
xnor U4240 (N_4240,N_3956,N_3082);
nand U4241 (N_4241,N_3657,N_3546);
nor U4242 (N_4242,N_3200,N_3127);
and U4243 (N_4243,N_3739,N_3581);
and U4244 (N_4244,N_3396,N_3404);
xor U4245 (N_4245,N_3493,N_3851);
nor U4246 (N_4246,N_3878,N_3886);
nand U4247 (N_4247,N_3758,N_3746);
nand U4248 (N_4248,N_3796,N_3297);
or U4249 (N_4249,N_3970,N_3968);
nand U4250 (N_4250,N_3552,N_3585);
or U4251 (N_4251,N_3094,N_3863);
or U4252 (N_4252,N_3022,N_3509);
and U4253 (N_4253,N_3083,N_3114);
nor U4254 (N_4254,N_3566,N_3925);
nand U4255 (N_4255,N_3617,N_3633);
nor U4256 (N_4256,N_3133,N_3519);
xor U4257 (N_4257,N_3242,N_3209);
xor U4258 (N_4258,N_3569,N_3318);
and U4259 (N_4259,N_3891,N_3245);
or U4260 (N_4260,N_3643,N_3351);
nor U4261 (N_4261,N_3100,N_3984);
or U4262 (N_4262,N_3044,N_3205);
xnor U4263 (N_4263,N_3718,N_3751);
nand U4264 (N_4264,N_3597,N_3227);
nand U4265 (N_4265,N_3437,N_3649);
and U4266 (N_4266,N_3823,N_3256);
or U4267 (N_4267,N_3098,N_3670);
xnor U4268 (N_4268,N_3774,N_3539);
and U4269 (N_4269,N_3124,N_3135);
or U4270 (N_4270,N_3832,N_3875);
or U4271 (N_4271,N_3560,N_3080);
nor U4272 (N_4272,N_3469,N_3436);
nand U4273 (N_4273,N_3363,N_3144);
and U4274 (N_4274,N_3343,N_3383);
nand U4275 (N_4275,N_3231,N_3853);
or U4276 (N_4276,N_3116,N_3408);
or U4277 (N_4277,N_3714,N_3260);
nand U4278 (N_4278,N_3207,N_3141);
or U4279 (N_4279,N_3433,N_3308);
or U4280 (N_4280,N_3101,N_3600);
or U4281 (N_4281,N_3272,N_3700);
or U4282 (N_4282,N_3757,N_3894);
or U4283 (N_4283,N_3596,N_3872);
nor U4284 (N_4284,N_3990,N_3025);
nand U4285 (N_4285,N_3276,N_3010);
xor U4286 (N_4286,N_3736,N_3987);
and U4287 (N_4287,N_3249,N_3191);
nand U4288 (N_4288,N_3392,N_3032);
xor U4289 (N_4289,N_3730,N_3228);
nor U4290 (N_4290,N_3536,N_3474);
xnor U4291 (N_4291,N_3580,N_3282);
or U4292 (N_4292,N_3511,N_3040);
or U4293 (N_4293,N_3563,N_3234);
or U4294 (N_4294,N_3154,N_3432);
or U4295 (N_4295,N_3018,N_3206);
nand U4296 (N_4296,N_3009,N_3732);
xor U4297 (N_4297,N_3950,N_3959);
or U4298 (N_4298,N_3381,N_3398);
xnor U4299 (N_4299,N_3640,N_3417);
nand U4300 (N_4300,N_3390,N_3782);
nor U4301 (N_4301,N_3578,N_3704);
or U4302 (N_4302,N_3176,N_3005);
and U4303 (N_4303,N_3464,N_3346);
nand U4304 (N_4304,N_3247,N_3265);
nor U4305 (N_4305,N_3115,N_3674);
nor U4306 (N_4306,N_3837,N_3949);
xnor U4307 (N_4307,N_3980,N_3882);
and U4308 (N_4308,N_3169,N_3834);
nor U4309 (N_4309,N_3273,N_3261);
and U4310 (N_4310,N_3818,N_3504);
xnor U4311 (N_4311,N_3406,N_3892);
or U4312 (N_4312,N_3695,N_3901);
xor U4313 (N_4313,N_3344,N_3121);
nand U4314 (N_4314,N_3626,N_3235);
nand U4315 (N_4315,N_3077,N_3309);
nor U4316 (N_4316,N_3710,N_3151);
xnor U4317 (N_4317,N_3846,N_3810);
xnor U4318 (N_4318,N_3199,N_3411);
nor U4319 (N_4319,N_3166,N_3379);
or U4320 (N_4320,N_3155,N_3319);
or U4321 (N_4321,N_3425,N_3972);
xnor U4322 (N_4322,N_3224,N_3013);
nand U4323 (N_4323,N_3688,N_3711);
nand U4324 (N_4324,N_3316,N_3402);
nor U4325 (N_4325,N_3157,N_3997);
nand U4326 (N_4326,N_3618,N_3403);
nor U4327 (N_4327,N_3784,N_3916);
nor U4328 (N_4328,N_3790,N_3138);
or U4329 (N_4329,N_3989,N_3244);
and U4330 (N_4330,N_3229,N_3933);
or U4331 (N_4331,N_3488,N_3508);
or U4332 (N_4332,N_3835,N_3164);
nand U4333 (N_4333,N_3738,N_3175);
xnor U4334 (N_4334,N_3336,N_3061);
and U4335 (N_4335,N_3524,N_3132);
xnor U4336 (N_4336,N_3128,N_3629);
xnor U4337 (N_4337,N_3955,N_3590);
and U4338 (N_4338,N_3034,N_3667);
or U4339 (N_4339,N_3516,N_3813);
xnor U4340 (N_4340,N_3995,N_3171);
nand U4341 (N_4341,N_3658,N_3880);
xnor U4342 (N_4342,N_3780,N_3767);
nor U4343 (N_4343,N_3720,N_3194);
nor U4344 (N_4344,N_3180,N_3556);
and U4345 (N_4345,N_3202,N_3677);
xor U4346 (N_4346,N_3868,N_3033);
xor U4347 (N_4347,N_3299,N_3967);
or U4348 (N_4348,N_3500,N_3963);
xnor U4349 (N_4349,N_3965,N_3936);
nand U4350 (N_4350,N_3368,N_3001);
xor U4351 (N_4351,N_3438,N_3068);
nand U4352 (N_4352,N_3060,N_3538);
xnor U4353 (N_4353,N_3041,N_3412);
nor U4354 (N_4354,N_3874,N_3377);
nand U4355 (N_4355,N_3703,N_3352);
nand U4356 (N_4356,N_3742,N_3125);
nand U4357 (N_4357,N_3680,N_3462);
xor U4358 (N_4358,N_3071,N_3599);
nor U4359 (N_4359,N_3698,N_3313);
nand U4360 (N_4360,N_3472,N_3096);
or U4361 (N_4361,N_3775,N_3789);
and U4362 (N_4362,N_3320,N_3342);
nand U4363 (N_4363,N_3861,N_3717);
and U4364 (N_4364,N_3137,N_3857);
and U4365 (N_4365,N_3345,N_3549);
and U4366 (N_4366,N_3099,N_3476);
nand U4367 (N_4367,N_3143,N_3145);
and U4368 (N_4368,N_3898,N_3440);
and U4369 (N_4369,N_3526,N_3384);
nor U4370 (N_4370,N_3439,N_3824);
or U4371 (N_4371,N_3870,N_3323);
or U4372 (N_4372,N_3682,N_3642);
xor U4373 (N_4373,N_3681,N_3840);
nor U4374 (N_4374,N_3850,N_3372);
xor U4375 (N_4375,N_3492,N_3557);
xnor U4376 (N_4376,N_3786,N_3811);
or U4377 (N_4377,N_3006,N_3458);
xnor U4378 (N_4378,N_3777,N_3605);
xnor U4379 (N_4379,N_3907,N_3793);
xor U4380 (N_4380,N_3819,N_3059);
xnor U4381 (N_4381,N_3198,N_3324);
or U4382 (N_4382,N_3471,N_3761);
and U4383 (N_4383,N_3806,N_3871);
or U4384 (N_4384,N_3338,N_3962);
nor U4385 (N_4385,N_3386,N_3178);
nand U4386 (N_4386,N_3221,N_3095);
nor U4387 (N_4387,N_3776,N_3283);
xor U4388 (N_4388,N_3140,N_3373);
or U4389 (N_4389,N_3920,N_3341);
and U4390 (N_4390,N_3766,N_3974);
xnor U4391 (N_4391,N_3173,N_3248);
xnor U4392 (N_4392,N_3482,N_3495);
or U4393 (N_4393,N_3884,N_3998);
nand U4394 (N_4394,N_3805,N_3921);
and U4395 (N_4395,N_3985,N_3601);
nor U4396 (N_4396,N_3520,N_3012);
and U4397 (N_4397,N_3073,N_3160);
or U4398 (N_4398,N_3606,N_3727);
nor U4399 (N_4399,N_3236,N_3278);
and U4400 (N_4400,N_3067,N_3634);
nor U4401 (N_4401,N_3902,N_3399);
and U4402 (N_4402,N_3184,N_3541);
or U4403 (N_4403,N_3030,N_3979);
or U4404 (N_4404,N_3105,N_3587);
or U4405 (N_4405,N_3865,N_3743);
and U4406 (N_4406,N_3522,N_3652);
nand U4407 (N_4407,N_3409,N_3478);
or U4408 (N_4408,N_3232,N_3540);
nor U4409 (N_4409,N_3653,N_3838);
xnor U4410 (N_4410,N_3513,N_3271);
and U4411 (N_4411,N_3031,N_3724);
nor U4412 (N_4412,N_3109,N_3940);
xor U4413 (N_4413,N_3636,N_3002);
and U4414 (N_4414,N_3610,N_3485);
nand U4415 (N_4415,N_3943,N_3147);
and U4416 (N_4416,N_3748,N_3731);
nor U4417 (N_4417,N_3016,N_3042);
and U4418 (N_4418,N_3477,N_3577);
nand U4419 (N_4419,N_3186,N_3918);
and U4420 (N_4420,N_3213,N_3922);
or U4421 (N_4421,N_3908,N_3468);
xor U4422 (N_4422,N_3565,N_3999);
nor U4423 (N_4423,N_3424,N_3303);
xor U4424 (N_4424,N_3969,N_3340);
nor U4425 (N_4425,N_3820,N_3787);
nand U4426 (N_4426,N_3201,N_3534);
or U4427 (N_4427,N_3117,N_3512);
nand U4428 (N_4428,N_3356,N_3881);
nand U4429 (N_4429,N_3189,N_3510);
and U4430 (N_4430,N_3752,N_3212);
or U4431 (N_4431,N_3269,N_3814);
xor U4432 (N_4432,N_3298,N_3615);
xnor U4433 (N_4433,N_3635,N_3455);
xor U4434 (N_4434,N_3414,N_3593);
xor U4435 (N_4435,N_3848,N_3055);
and U4436 (N_4436,N_3497,N_3964);
nand U4437 (N_4437,N_3014,N_3568);
xnor U4438 (N_4438,N_3745,N_3051);
nor U4439 (N_4439,N_3431,N_3641);
or U4440 (N_4440,N_3622,N_3388);
or U4441 (N_4441,N_3295,N_3490);
and U4442 (N_4442,N_3311,N_3821);
and U4443 (N_4443,N_3684,N_3586);
or U4444 (N_4444,N_3023,N_3773);
or U4445 (N_4445,N_3662,N_3241);
nor U4446 (N_4446,N_3394,N_3072);
nor U4447 (N_4447,N_3583,N_3528);
nand U4448 (N_4448,N_3862,N_3887);
nor U4449 (N_4449,N_3159,N_3668);
nor U4450 (N_4450,N_3146,N_3337);
xnor U4451 (N_4451,N_3091,N_3804);
or U4452 (N_4452,N_3864,N_3760);
xnor U4453 (N_4453,N_3279,N_3771);
nor U4454 (N_4454,N_3530,N_3334);
nand U4455 (N_4455,N_3735,N_3696);
and U4456 (N_4456,N_3948,N_3919);
nor U4457 (N_4457,N_3624,N_3087);
and U4458 (N_4458,N_3000,N_3594);
nand U4459 (N_4459,N_3366,N_3910);
xor U4460 (N_4460,N_3608,N_3466);
or U4461 (N_4461,N_3459,N_3798);
or U4462 (N_4462,N_3632,N_3620);
or U4463 (N_4463,N_3982,N_3434);
nor U4464 (N_4464,N_3993,N_3262);
xor U4465 (N_4465,N_3799,N_3627);
and U4466 (N_4466,N_3057,N_3415);
nand U4467 (N_4467,N_3065,N_3007);
xor U4468 (N_4468,N_3734,N_3912);
nand U4469 (N_4469,N_3675,N_3801);
and U4470 (N_4470,N_3562,N_3085);
and U4471 (N_4471,N_3370,N_3047);
nor U4472 (N_4472,N_3358,N_3564);
or U4473 (N_4473,N_3162,N_3389);
and U4474 (N_4474,N_3852,N_3367);
nand U4475 (N_4475,N_3591,N_3905);
and U4476 (N_4476,N_3052,N_3329);
nor U4477 (N_4477,N_3473,N_3826);
nor U4478 (N_4478,N_3426,N_3572);
and U4479 (N_4479,N_3129,N_3678);
nor U4480 (N_4480,N_3429,N_3676);
and U4481 (N_4481,N_3665,N_3986);
nor U4482 (N_4482,N_3706,N_3876);
nor U4483 (N_4483,N_3934,N_3800);
or U4484 (N_4484,N_3118,N_3788);
nor U4485 (N_4485,N_3729,N_3355);
xor U4486 (N_4486,N_3410,N_3893);
and U4487 (N_4487,N_3829,N_3465);
and U4488 (N_4488,N_3931,N_3498);
nor U4489 (N_4489,N_3046,N_3631);
xnor U4490 (N_4490,N_3050,N_3842);
and U4491 (N_4491,N_3750,N_3187);
nand U4492 (N_4492,N_3327,N_3401);
or U4493 (N_4493,N_3454,N_3008);
nor U4494 (N_4494,N_3699,N_3357);
nand U4495 (N_4495,N_3079,N_3797);
xor U4496 (N_4496,N_3899,N_3883);
nand U4497 (N_4497,N_3123,N_3709);
nand U4498 (N_4498,N_3195,N_3604);
and U4499 (N_4499,N_3421,N_3219);
and U4500 (N_4500,N_3312,N_3971);
nand U4501 (N_4501,N_3379,N_3294);
nor U4502 (N_4502,N_3434,N_3198);
nand U4503 (N_4503,N_3524,N_3072);
xor U4504 (N_4504,N_3106,N_3906);
nor U4505 (N_4505,N_3950,N_3565);
and U4506 (N_4506,N_3909,N_3744);
nand U4507 (N_4507,N_3102,N_3844);
nor U4508 (N_4508,N_3453,N_3710);
or U4509 (N_4509,N_3734,N_3867);
nor U4510 (N_4510,N_3333,N_3160);
xnor U4511 (N_4511,N_3972,N_3335);
or U4512 (N_4512,N_3267,N_3626);
xor U4513 (N_4513,N_3383,N_3381);
nor U4514 (N_4514,N_3298,N_3147);
and U4515 (N_4515,N_3218,N_3122);
and U4516 (N_4516,N_3695,N_3847);
xor U4517 (N_4517,N_3840,N_3754);
xnor U4518 (N_4518,N_3601,N_3440);
nand U4519 (N_4519,N_3402,N_3626);
or U4520 (N_4520,N_3807,N_3292);
or U4521 (N_4521,N_3546,N_3841);
nand U4522 (N_4522,N_3064,N_3139);
nor U4523 (N_4523,N_3385,N_3973);
xnor U4524 (N_4524,N_3136,N_3475);
and U4525 (N_4525,N_3091,N_3935);
or U4526 (N_4526,N_3916,N_3818);
nor U4527 (N_4527,N_3128,N_3228);
or U4528 (N_4528,N_3827,N_3214);
nand U4529 (N_4529,N_3665,N_3450);
nor U4530 (N_4530,N_3737,N_3371);
nand U4531 (N_4531,N_3520,N_3369);
or U4532 (N_4532,N_3624,N_3924);
nand U4533 (N_4533,N_3279,N_3259);
and U4534 (N_4534,N_3112,N_3215);
nand U4535 (N_4535,N_3064,N_3684);
or U4536 (N_4536,N_3483,N_3112);
nor U4537 (N_4537,N_3764,N_3607);
nand U4538 (N_4538,N_3145,N_3425);
or U4539 (N_4539,N_3368,N_3941);
nor U4540 (N_4540,N_3916,N_3241);
nand U4541 (N_4541,N_3733,N_3213);
or U4542 (N_4542,N_3380,N_3562);
nor U4543 (N_4543,N_3000,N_3611);
nand U4544 (N_4544,N_3768,N_3301);
and U4545 (N_4545,N_3224,N_3380);
xnor U4546 (N_4546,N_3976,N_3675);
nor U4547 (N_4547,N_3884,N_3821);
xor U4548 (N_4548,N_3089,N_3257);
and U4549 (N_4549,N_3051,N_3695);
nand U4550 (N_4550,N_3565,N_3657);
or U4551 (N_4551,N_3791,N_3029);
and U4552 (N_4552,N_3368,N_3495);
and U4553 (N_4553,N_3183,N_3292);
nand U4554 (N_4554,N_3610,N_3548);
and U4555 (N_4555,N_3271,N_3796);
xor U4556 (N_4556,N_3627,N_3468);
xor U4557 (N_4557,N_3650,N_3577);
or U4558 (N_4558,N_3304,N_3299);
xnor U4559 (N_4559,N_3248,N_3700);
nor U4560 (N_4560,N_3198,N_3250);
xnor U4561 (N_4561,N_3303,N_3260);
or U4562 (N_4562,N_3780,N_3575);
nand U4563 (N_4563,N_3454,N_3131);
xor U4564 (N_4564,N_3483,N_3969);
nor U4565 (N_4565,N_3355,N_3027);
and U4566 (N_4566,N_3521,N_3922);
nand U4567 (N_4567,N_3711,N_3533);
and U4568 (N_4568,N_3175,N_3000);
nand U4569 (N_4569,N_3449,N_3103);
nand U4570 (N_4570,N_3767,N_3645);
and U4571 (N_4571,N_3997,N_3916);
and U4572 (N_4572,N_3030,N_3156);
or U4573 (N_4573,N_3386,N_3857);
and U4574 (N_4574,N_3893,N_3272);
and U4575 (N_4575,N_3362,N_3329);
nor U4576 (N_4576,N_3384,N_3603);
and U4577 (N_4577,N_3635,N_3777);
nand U4578 (N_4578,N_3395,N_3553);
xor U4579 (N_4579,N_3052,N_3402);
or U4580 (N_4580,N_3550,N_3069);
xnor U4581 (N_4581,N_3664,N_3764);
or U4582 (N_4582,N_3897,N_3961);
nand U4583 (N_4583,N_3798,N_3756);
xnor U4584 (N_4584,N_3047,N_3168);
nand U4585 (N_4585,N_3656,N_3379);
xnor U4586 (N_4586,N_3969,N_3812);
xor U4587 (N_4587,N_3904,N_3304);
nand U4588 (N_4588,N_3277,N_3312);
nand U4589 (N_4589,N_3103,N_3076);
nand U4590 (N_4590,N_3635,N_3789);
xnor U4591 (N_4591,N_3368,N_3510);
and U4592 (N_4592,N_3837,N_3975);
or U4593 (N_4593,N_3271,N_3847);
xnor U4594 (N_4594,N_3200,N_3779);
nor U4595 (N_4595,N_3388,N_3470);
and U4596 (N_4596,N_3867,N_3865);
nor U4597 (N_4597,N_3028,N_3578);
xor U4598 (N_4598,N_3481,N_3631);
nor U4599 (N_4599,N_3956,N_3805);
nand U4600 (N_4600,N_3412,N_3234);
and U4601 (N_4601,N_3536,N_3519);
or U4602 (N_4602,N_3706,N_3862);
xnor U4603 (N_4603,N_3939,N_3168);
or U4604 (N_4604,N_3014,N_3366);
and U4605 (N_4605,N_3107,N_3290);
nor U4606 (N_4606,N_3528,N_3002);
nand U4607 (N_4607,N_3116,N_3163);
nand U4608 (N_4608,N_3430,N_3076);
and U4609 (N_4609,N_3848,N_3038);
and U4610 (N_4610,N_3859,N_3335);
xor U4611 (N_4611,N_3945,N_3294);
xor U4612 (N_4612,N_3907,N_3435);
or U4613 (N_4613,N_3272,N_3611);
and U4614 (N_4614,N_3277,N_3850);
or U4615 (N_4615,N_3236,N_3674);
nor U4616 (N_4616,N_3847,N_3936);
or U4617 (N_4617,N_3780,N_3065);
and U4618 (N_4618,N_3830,N_3139);
nand U4619 (N_4619,N_3674,N_3261);
and U4620 (N_4620,N_3535,N_3412);
nand U4621 (N_4621,N_3375,N_3828);
xnor U4622 (N_4622,N_3040,N_3973);
xor U4623 (N_4623,N_3755,N_3579);
nand U4624 (N_4624,N_3414,N_3370);
nand U4625 (N_4625,N_3149,N_3976);
nor U4626 (N_4626,N_3983,N_3389);
or U4627 (N_4627,N_3207,N_3061);
nor U4628 (N_4628,N_3782,N_3096);
and U4629 (N_4629,N_3678,N_3225);
nand U4630 (N_4630,N_3870,N_3185);
or U4631 (N_4631,N_3721,N_3801);
xnor U4632 (N_4632,N_3836,N_3224);
and U4633 (N_4633,N_3949,N_3803);
or U4634 (N_4634,N_3741,N_3964);
and U4635 (N_4635,N_3520,N_3668);
and U4636 (N_4636,N_3406,N_3786);
nand U4637 (N_4637,N_3273,N_3085);
nor U4638 (N_4638,N_3313,N_3654);
nor U4639 (N_4639,N_3154,N_3004);
or U4640 (N_4640,N_3611,N_3953);
nand U4641 (N_4641,N_3852,N_3552);
and U4642 (N_4642,N_3892,N_3774);
xor U4643 (N_4643,N_3173,N_3324);
xnor U4644 (N_4644,N_3385,N_3366);
xnor U4645 (N_4645,N_3450,N_3762);
nor U4646 (N_4646,N_3080,N_3568);
and U4647 (N_4647,N_3812,N_3083);
or U4648 (N_4648,N_3432,N_3234);
xor U4649 (N_4649,N_3922,N_3556);
xnor U4650 (N_4650,N_3107,N_3967);
nor U4651 (N_4651,N_3937,N_3513);
or U4652 (N_4652,N_3054,N_3214);
and U4653 (N_4653,N_3565,N_3990);
nand U4654 (N_4654,N_3367,N_3339);
or U4655 (N_4655,N_3791,N_3319);
and U4656 (N_4656,N_3084,N_3210);
nor U4657 (N_4657,N_3833,N_3066);
nor U4658 (N_4658,N_3231,N_3242);
and U4659 (N_4659,N_3420,N_3913);
and U4660 (N_4660,N_3478,N_3405);
nor U4661 (N_4661,N_3298,N_3884);
xnor U4662 (N_4662,N_3759,N_3407);
xor U4663 (N_4663,N_3126,N_3774);
xor U4664 (N_4664,N_3970,N_3330);
xor U4665 (N_4665,N_3837,N_3738);
nor U4666 (N_4666,N_3627,N_3013);
nand U4667 (N_4667,N_3360,N_3968);
nand U4668 (N_4668,N_3823,N_3772);
or U4669 (N_4669,N_3342,N_3343);
nand U4670 (N_4670,N_3974,N_3808);
xor U4671 (N_4671,N_3401,N_3424);
nand U4672 (N_4672,N_3079,N_3636);
or U4673 (N_4673,N_3354,N_3823);
or U4674 (N_4674,N_3029,N_3081);
nand U4675 (N_4675,N_3023,N_3738);
nor U4676 (N_4676,N_3137,N_3418);
or U4677 (N_4677,N_3224,N_3912);
nand U4678 (N_4678,N_3280,N_3759);
xor U4679 (N_4679,N_3864,N_3180);
nor U4680 (N_4680,N_3465,N_3909);
or U4681 (N_4681,N_3118,N_3295);
or U4682 (N_4682,N_3470,N_3393);
xnor U4683 (N_4683,N_3179,N_3660);
nor U4684 (N_4684,N_3912,N_3273);
and U4685 (N_4685,N_3863,N_3565);
nor U4686 (N_4686,N_3654,N_3808);
nor U4687 (N_4687,N_3503,N_3443);
nor U4688 (N_4688,N_3769,N_3579);
nor U4689 (N_4689,N_3607,N_3477);
nor U4690 (N_4690,N_3051,N_3179);
or U4691 (N_4691,N_3008,N_3448);
nor U4692 (N_4692,N_3108,N_3211);
nor U4693 (N_4693,N_3374,N_3459);
nor U4694 (N_4694,N_3937,N_3882);
xor U4695 (N_4695,N_3367,N_3443);
xnor U4696 (N_4696,N_3510,N_3051);
xor U4697 (N_4697,N_3228,N_3324);
and U4698 (N_4698,N_3488,N_3928);
xor U4699 (N_4699,N_3194,N_3732);
nor U4700 (N_4700,N_3092,N_3202);
xnor U4701 (N_4701,N_3746,N_3248);
and U4702 (N_4702,N_3702,N_3682);
nor U4703 (N_4703,N_3020,N_3268);
or U4704 (N_4704,N_3796,N_3275);
nor U4705 (N_4705,N_3204,N_3709);
nor U4706 (N_4706,N_3407,N_3108);
xor U4707 (N_4707,N_3948,N_3079);
nor U4708 (N_4708,N_3721,N_3280);
nor U4709 (N_4709,N_3897,N_3071);
nor U4710 (N_4710,N_3343,N_3509);
xnor U4711 (N_4711,N_3447,N_3963);
or U4712 (N_4712,N_3249,N_3816);
nand U4713 (N_4713,N_3638,N_3625);
xnor U4714 (N_4714,N_3570,N_3756);
nor U4715 (N_4715,N_3904,N_3188);
or U4716 (N_4716,N_3835,N_3501);
or U4717 (N_4717,N_3852,N_3891);
nand U4718 (N_4718,N_3436,N_3539);
or U4719 (N_4719,N_3157,N_3015);
nor U4720 (N_4720,N_3380,N_3468);
nor U4721 (N_4721,N_3746,N_3234);
or U4722 (N_4722,N_3508,N_3958);
and U4723 (N_4723,N_3572,N_3276);
nor U4724 (N_4724,N_3853,N_3168);
xnor U4725 (N_4725,N_3892,N_3217);
and U4726 (N_4726,N_3937,N_3798);
or U4727 (N_4727,N_3528,N_3059);
nand U4728 (N_4728,N_3769,N_3482);
or U4729 (N_4729,N_3691,N_3987);
xnor U4730 (N_4730,N_3513,N_3099);
nand U4731 (N_4731,N_3089,N_3254);
and U4732 (N_4732,N_3199,N_3756);
or U4733 (N_4733,N_3562,N_3604);
nor U4734 (N_4734,N_3210,N_3124);
and U4735 (N_4735,N_3029,N_3905);
nand U4736 (N_4736,N_3479,N_3007);
or U4737 (N_4737,N_3091,N_3354);
nor U4738 (N_4738,N_3745,N_3277);
xor U4739 (N_4739,N_3524,N_3285);
nand U4740 (N_4740,N_3796,N_3357);
xor U4741 (N_4741,N_3623,N_3617);
or U4742 (N_4742,N_3316,N_3874);
xnor U4743 (N_4743,N_3064,N_3096);
and U4744 (N_4744,N_3137,N_3091);
nand U4745 (N_4745,N_3202,N_3498);
nand U4746 (N_4746,N_3654,N_3756);
and U4747 (N_4747,N_3170,N_3258);
nor U4748 (N_4748,N_3925,N_3820);
xor U4749 (N_4749,N_3301,N_3285);
and U4750 (N_4750,N_3044,N_3198);
and U4751 (N_4751,N_3821,N_3986);
xnor U4752 (N_4752,N_3199,N_3240);
nand U4753 (N_4753,N_3302,N_3942);
and U4754 (N_4754,N_3868,N_3699);
xnor U4755 (N_4755,N_3025,N_3976);
and U4756 (N_4756,N_3350,N_3896);
or U4757 (N_4757,N_3412,N_3227);
xor U4758 (N_4758,N_3225,N_3606);
nor U4759 (N_4759,N_3641,N_3198);
nor U4760 (N_4760,N_3484,N_3700);
nor U4761 (N_4761,N_3403,N_3203);
and U4762 (N_4762,N_3078,N_3308);
and U4763 (N_4763,N_3647,N_3201);
and U4764 (N_4764,N_3347,N_3842);
xnor U4765 (N_4765,N_3053,N_3733);
nor U4766 (N_4766,N_3730,N_3798);
nand U4767 (N_4767,N_3461,N_3232);
xor U4768 (N_4768,N_3204,N_3207);
nand U4769 (N_4769,N_3661,N_3991);
nor U4770 (N_4770,N_3269,N_3117);
nor U4771 (N_4771,N_3140,N_3613);
or U4772 (N_4772,N_3478,N_3931);
nor U4773 (N_4773,N_3582,N_3215);
nand U4774 (N_4774,N_3802,N_3170);
nor U4775 (N_4775,N_3501,N_3850);
or U4776 (N_4776,N_3164,N_3369);
nand U4777 (N_4777,N_3321,N_3560);
xnor U4778 (N_4778,N_3679,N_3040);
nand U4779 (N_4779,N_3214,N_3332);
or U4780 (N_4780,N_3443,N_3233);
or U4781 (N_4781,N_3328,N_3384);
nand U4782 (N_4782,N_3468,N_3082);
nor U4783 (N_4783,N_3555,N_3093);
and U4784 (N_4784,N_3791,N_3134);
xor U4785 (N_4785,N_3754,N_3061);
and U4786 (N_4786,N_3177,N_3628);
or U4787 (N_4787,N_3175,N_3550);
nor U4788 (N_4788,N_3579,N_3453);
nand U4789 (N_4789,N_3520,N_3897);
xor U4790 (N_4790,N_3426,N_3570);
and U4791 (N_4791,N_3437,N_3329);
nand U4792 (N_4792,N_3430,N_3602);
nand U4793 (N_4793,N_3996,N_3036);
nand U4794 (N_4794,N_3988,N_3674);
nand U4795 (N_4795,N_3756,N_3827);
xor U4796 (N_4796,N_3983,N_3613);
xor U4797 (N_4797,N_3621,N_3328);
and U4798 (N_4798,N_3679,N_3163);
nor U4799 (N_4799,N_3110,N_3464);
and U4800 (N_4800,N_3935,N_3411);
xor U4801 (N_4801,N_3156,N_3935);
nand U4802 (N_4802,N_3504,N_3958);
nand U4803 (N_4803,N_3973,N_3606);
xnor U4804 (N_4804,N_3955,N_3485);
nor U4805 (N_4805,N_3036,N_3534);
and U4806 (N_4806,N_3231,N_3009);
nor U4807 (N_4807,N_3288,N_3913);
xnor U4808 (N_4808,N_3520,N_3851);
and U4809 (N_4809,N_3644,N_3205);
xor U4810 (N_4810,N_3087,N_3200);
or U4811 (N_4811,N_3083,N_3431);
xnor U4812 (N_4812,N_3438,N_3686);
or U4813 (N_4813,N_3264,N_3830);
and U4814 (N_4814,N_3407,N_3880);
xnor U4815 (N_4815,N_3009,N_3966);
or U4816 (N_4816,N_3099,N_3933);
nand U4817 (N_4817,N_3870,N_3454);
or U4818 (N_4818,N_3808,N_3022);
xnor U4819 (N_4819,N_3481,N_3737);
and U4820 (N_4820,N_3784,N_3998);
nand U4821 (N_4821,N_3902,N_3591);
xnor U4822 (N_4822,N_3135,N_3462);
and U4823 (N_4823,N_3200,N_3580);
nor U4824 (N_4824,N_3818,N_3820);
xor U4825 (N_4825,N_3305,N_3059);
and U4826 (N_4826,N_3882,N_3078);
nor U4827 (N_4827,N_3879,N_3258);
and U4828 (N_4828,N_3587,N_3607);
nand U4829 (N_4829,N_3290,N_3347);
or U4830 (N_4830,N_3020,N_3161);
nand U4831 (N_4831,N_3433,N_3398);
and U4832 (N_4832,N_3420,N_3908);
and U4833 (N_4833,N_3388,N_3739);
xnor U4834 (N_4834,N_3048,N_3883);
nor U4835 (N_4835,N_3213,N_3119);
nor U4836 (N_4836,N_3454,N_3425);
or U4837 (N_4837,N_3086,N_3302);
and U4838 (N_4838,N_3346,N_3853);
nor U4839 (N_4839,N_3503,N_3270);
nor U4840 (N_4840,N_3471,N_3057);
nand U4841 (N_4841,N_3523,N_3896);
or U4842 (N_4842,N_3799,N_3909);
nand U4843 (N_4843,N_3532,N_3271);
nor U4844 (N_4844,N_3662,N_3428);
nand U4845 (N_4845,N_3457,N_3801);
nor U4846 (N_4846,N_3614,N_3441);
nand U4847 (N_4847,N_3894,N_3006);
nand U4848 (N_4848,N_3746,N_3092);
nor U4849 (N_4849,N_3405,N_3739);
or U4850 (N_4850,N_3605,N_3365);
nand U4851 (N_4851,N_3519,N_3114);
nand U4852 (N_4852,N_3356,N_3458);
or U4853 (N_4853,N_3929,N_3795);
xnor U4854 (N_4854,N_3121,N_3470);
or U4855 (N_4855,N_3914,N_3839);
nor U4856 (N_4856,N_3847,N_3473);
nor U4857 (N_4857,N_3701,N_3165);
nor U4858 (N_4858,N_3429,N_3094);
or U4859 (N_4859,N_3335,N_3779);
nand U4860 (N_4860,N_3462,N_3688);
or U4861 (N_4861,N_3726,N_3464);
xor U4862 (N_4862,N_3594,N_3046);
xnor U4863 (N_4863,N_3660,N_3757);
xnor U4864 (N_4864,N_3990,N_3042);
nand U4865 (N_4865,N_3936,N_3176);
nor U4866 (N_4866,N_3870,N_3105);
nand U4867 (N_4867,N_3147,N_3281);
nor U4868 (N_4868,N_3949,N_3600);
and U4869 (N_4869,N_3582,N_3431);
nor U4870 (N_4870,N_3683,N_3001);
nand U4871 (N_4871,N_3536,N_3446);
xor U4872 (N_4872,N_3799,N_3860);
nor U4873 (N_4873,N_3887,N_3345);
nand U4874 (N_4874,N_3054,N_3821);
nor U4875 (N_4875,N_3393,N_3239);
nor U4876 (N_4876,N_3573,N_3365);
or U4877 (N_4877,N_3054,N_3203);
nor U4878 (N_4878,N_3084,N_3249);
nor U4879 (N_4879,N_3825,N_3878);
and U4880 (N_4880,N_3245,N_3058);
nand U4881 (N_4881,N_3411,N_3921);
xor U4882 (N_4882,N_3351,N_3767);
or U4883 (N_4883,N_3526,N_3674);
and U4884 (N_4884,N_3608,N_3147);
nor U4885 (N_4885,N_3715,N_3930);
nor U4886 (N_4886,N_3921,N_3863);
and U4887 (N_4887,N_3500,N_3034);
or U4888 (N_4888,N_3362,N_3778);
xnor U4889 (N_4889,N_3083,N_3924);
or U4890 (N_4890,N_3311,N_3704);
or U4891 (N_4891,N_3006,N_3553);
nand U4892 (N_4892,N_3334,N_3911);
xnor U4893 (N_4893,N_3895,N_3667);
and U4894 (N_4894,N_3159,N_3637);
nand U4895 (N_4895,N_3984,N_3742);
nor U4896 (N_4896,N_3979,N_3203);
nand U4897 (N_4897,N_3578,N_3606);
nand U4898 (N_4898,N_3099,N_3841);
nor U4899 (N_4899,N_3430,N_3334);
or U4900 (N_4900,N_3290,N_3970);
nand U4901 (N_4901,N_3482,N_3652);
and U4902 (N_4902,N_3041,N_3695);
and U4903 (N_4903,N_3380,N_3222);
nor U4904 (N_4904,N_3347,N_3818);
nand U4905 (N_4905,N_3419,N_3858);
xnor U4906 (N_4906,N_3127,N_3829);
and U4907 (N_4907,N_3126,N_3784);
nor U4908 (N_4908,N_3918,N_3473);
and U4909 (N_4909,N_3473,N_3154);
nand U4910 (N_4910,N_3697,N_3650);
nand U4911 (N_4911,N_3948,N_3273);
nand U4912 (N_4912,N_3922,N_3898);
nor U4913 (N_4913,N_3012,N_3133);
nor U4914 (N_4914,N_3221,N_3568);
nand U4915 (N_4915,N_3085,N_3877);
xnor U4916 (N_4916,N_3269,N_3002);
nor U4917 (N_4917,N_3981,N_3427);
xor U4918 (N_4918,N_3243,N_3678);
xor U4919 (N_4919,N_3226,N_3048);
xnor U4920 (N_4920,N_3977,N_3513);
nand U4921 (N_4921,N_3587,N_3392);
xor U4922 (N_4922,N_3929,N_3114);
nand U4923 (N_4923,N_3582,N_3183);
nand U4924 (N_4924,N_3281,N_3457);
xnor U4925 (N_4925,N_3082,N_3628);
xor U4926 (N_4926,N_3833,N_3209);
xnor U4927 (N_4927,N_3857,N_3928);
xor U4928 (N_4928,N_3157,N_3888);
and U4929 (N_4929,N_3186,N_3973);
xnor U4930 (N_4930,N_3895,N_3270);
nand U4931 (N_4931,N_3205,N_3103);
or U4932 (N_4932,N_3499,N_3664);
nor U4933 (N_4933,N_3923,N_3855);
nor U4934 (N_4934,N_3726,N_3687);
and U4935 (N_4935,N_3080,N_3276);
nand U4936 (N_4936,N_3769,N_3120);
nand U4937 (N_4937,N_3519,N_3200);
nand U4938 (N_4938,N_3068,N_3034);
and U4939 (N_4939,N_3062,N_3794);
and U4940 (N_4940,N_3982,N_3289);
or U4941 (N_4941,N_3841,N_3469);
nor U4942 (N_4942,N_3659,N_3836);
nand U4943 (N_4943,N_3664,N_3249);
and U4944 (N_4944,N_3075,N_3067);
xnor U4945 (N_4945,N_3404,N_3071);
or U4946 (N_4946,N_3154,N_3827);
xor U4947 (N_4947,N_3648,N_3275);
nor U4948 (N_4948,N_3023,N_3841);
or U4949 (N_4949,N_3767,N_3400);
xnor U4950 (N_4950,N_3506,N_3458);
nand U4951 (N_4951,N_3437,N_3006);
and U4952 (N_4952,N_3231,N_3672);
or U4953 (N_4953,N_3354,N_3482);
or U4954 (N_4954,N_3279,N_3437);
and U4955 (N_4955,N_3834,N_3142);
and U4956 (N_4956,N_3127,N_3195);
nor U4957 (N_4957,N_3993,N_3458);
nand U4958 (N_4958,N_3933,N_3717);
nor U4959 (N_4959,N_3901,N_3121);
xor U4960 (N_4960,N_3492,N_3414);
or U4961 (N_4961,N_3525,N_3076);
or U4962 (N_4962,N_3155,N_3339);
and U4963 (N_4963,N_3818,N_3385);
and U4964 (N_4964,N_3164,N_3529);
nand U4965 (N_4965,N_3247,N_3592);
nand U4966 (N_4966,N_3001,N_3209);
and U4967 (N_4967,N_3154,N_3980);
and U4968 (N_4968,N_3502,N_3160);
nand U4969 (N_4969,N_3090,N_3664);
and U4970 (N_4970,N_3327,N_3728);
nand U4971 (N_4971,N_3169,N_3578);
or U4972 (N_4972,N_3560,N_3381);
and U4973 (N_4973,N_3270,N_3858);
or U4974 (N_4974,N_3065,N_3634);
nor U4975 (N_4975,N_3848,N_3290);
nand U4976 (N_4976,N_3459,N_3627);
and U4977 (N_4977,N_3544,N_3250);
or U4978 (N_4978,N_3432,N_3995);
and U4979 (N_4979,N_3368,N_3902);
nand U4980 (N_4980,N_3945,N_3717);
or U4981 (N_4981,N_3447,N_3362);
xnor U4982 (N_4982,N_3156,N_3686);
nor U4983 (N_4983,N_3207,N_3262);
xnor U4984 (N_4984,N_3829,N_3454);
nand U4985 (N_4985,N_3169,N_3708);
nand U4986 (N_4986,N_3166,N_3447);
and U4987 (N_4987,N_3665,N_3445);
xor U4988 (N_4988,N_3928,N_3974);
or U4989 (N_4989,N_3438,N_3582);
nand U4990 (N_4990,N_3029,N_3322);
and U4991 (N_4991,N_3635,N_3798);
xor U4992 (N_4992,N_3250,N_3887);
nor U4993 (N_4993,N_3246,N_3124);
nand U4994 (N_4994,N_3641,N_3259);
and U4995 (N_4995,N_3958,N_3101);
nand U4996 (N_4996,N_3705,N_3786);
or U4997 (N_4997,N_3968,N_3103);
or U4998 (N_4998,N_3520,N_3137);
xor U4999 (N_4999,N_3913,N_3405);
and U5000 (N_5000,N_4820,N_4100);
nor U5001 (N_5001,N_4049,N_4396);
or U5002 (N_5002,N_4409,N_4404);
or U5003 (N_5003,N_4014,N_4304);
and U5004 (N_5004,N_4452,N_4330);
or U5005 (N_5005,N_4983,N_4532);
or U5006 (N_5006,N_4564,N_4589);
nor U5007 (N_5007,N_4126,N_4852);
and U5008 (N_5008,N_4981,N_4553);
and U5009 (N_5009,N_4137,N_4345);
or U5010 (N_5010,N_4988,N_4869);
nand U5011 (N_5011,N_4075,N_4847);
nor U5012 (N_5012,N_4510,N_4406);
or U5013 (N_5013,N_4633,N_4459);
and U5014 (N_5014,N_4796,N_4332);
and U5015 (N_5015,N_4756,N_4766);
and U5016 (N_5016,N_4210,N_4809);
nand U5017 (N_5017,N_4355,N_4397);
xnor U5018 (N_5018,N_4993,N_4176);
nor U5019 (N_5019,N_4753,N_4867);
xor U5020 (N_5020,N_4090,N_4307);
nand U5021 (N_5021,N_4819,N_4623);
or U5022 (N_5022,N_4393,N_4688);
and U5023 (N_5023,N_4036,N_4260);
xnor U5024 (N_5024,N_4984,N_4389);
nand U5025 (N_5025,N_4377,N_4177);
nand U5026 (N_5026,N_4838,N_4598);
xnor U5027 (N_5027,N_4431,N_4597);
nand U5028 (N_5028,N_4798,N_4654);
xor U5029 (N_5029,N_4708,N_4735);
nand U5030 (N_5030,N_4773,N_4799);
and U5031 (N_5031,N_4777,N_4349);
and U5032 (N_5032,N_4618,N_4804);
xnor U5033 (N_5033,N_4845,N_4987);
nand U5034 (N_5034,N_4982,N_4353);
or U5035 (N_5035,N_4682,N_4270);
nor U5036 (N_5036,N_4932,N_4506);
or U5037 (N_5037,N_4939,N_4687);
nor U5038 (N_5038,N_4060,N_4175);
or U5039 (N_5039,N_4219,N_4944);
and U5040 (N_5040,N_4976,N_4134);
nand U5041 (N_5041,N_4830,N_4476);
nor U5042 (N_5042,N_4948,N_4681);
or U5043 (N_5043,N_4061,N_4817);
xnor U5044 (N_5044,N_4964,N_4733);
xnor U5045 (N_5045,N_4354,N_4627);
xnor U5046 (N_5046,N_4447,N_4956);
or U5047 (N_5047,N_4474,N_4356);
xor U5048 (N_5048,N_4823,N_4325);
or U5049 (N_5049,N_4873,N_4123);
and U5050 (N_5050,N_4818,N_4555);
and U5051 (N_5051,N_4664,N_4466);
and U5052 (N_5052,N_4376,N_4714);
xnor U5053 (N_5053,N_4395,N_4016);
nor U5054 (N_5054,N_4001,N_4770);
nor U5055 (N_5055,N_4346,N_4730);
or U5056 (N_5056,N_4684,N_4585);
nand U5057 (N_5057,N_4509,N_4430);
nand U5058 (N_5058,N_4282,N_4755);
and U5059 (N_5059,N_4563,N_4054);
nor U5060 (N_5060,N_4806,N_4924);
and U5061 (N_5061,N_4294,N_4569);
xnor U5062 (N_5062,N_4504,N_4583);
nor U5063 (N_5063,N_4386,N_4243);
nand U5064 (N_5064,N_4212,N_4401);
nand U5065 (N_5065,N_4518,N_4275);
xor U5066 (N_5066,N_4320,N_4704);
or U5067 (N_5067,N_4158,N_4925);
or U5068 (N_5068,N_4043,N_4870);
nor U5069 (N_5069,N_4846,N_4696);
or U5070 (N_5070,N_4881,N_4022);
xnor U5071 (N_5071,N_4234,N_4534);
or U5072 (N_5072,N_4482,N_4199);
and U5073 (N_5073,N_4239,N_4822);
and U5074 (N_5074,N_4003,N_4029);
and U5075 (N_5075,N_4827,N_4266);
and U5076 (N_5076,N_4667,N_4642);
nor U5077 (N_5077,N_4550,N_4237);
xor U5078 (N_5078,N_4183,N_4146);
nor U5079 (N_5079,N_4306,N_4546);
and U5080 (N_5080,N_4006,N_4295);
nand U5081 (N_5081,N_4094,N_4596);
or U5082 (N_5082,N_4473,N_4480);
xnor U5083 (N_5083,N_4200,N_4505);
or U5084 (N_5084,N_4858,N_4617);
or U5085 (N_5085,N_4138,N_4762);
or U5086 (N_5086,N_4971,N_4256);
nand U5087 (N_5087,N_4497,N_4795);
nand U5088 (N_5088,N_4802,N_4500);
and U5089 (N_5089,N_4740,N_4368);
xor U5090 (N_5090,N_4685,N_4771);
or U5091 (N_5091,N_4197,N_4025);
xnor U5092 (N_5092,N_4917,N_4539);
nand U5093 (N_5093,N_4188,N_4149);
nand U5094 (N_5094,N_4267,N_4233);
or U5095 (N_5095,N_4050,N_4615);
and U5096 (N_5096,N_4652,N_4910);
nand U5097 (N_5097,N_4141,N_4666);
xor U5098 (N_5098,N_4039,N_4861);
or U5099 (N_5099,N_4479,N_4659);
nand U5100 (N_5100,N_4384,N_4454);
nand U5101 (N_5101,N_4651,N_4579);
nand U5102 (N_5102,N_4463,N_4276);
nor U5103 (N_5103,N_4637,N_4879);
and U5104 (N_5104,N_4350,N_4220);
or U5105 (N_5105,N_4783,N_4545);
and U5106 (N_5106,N_4883,N_4201);
or U5107 (N_5107,N_4106,N_4418);
and U5108 (N_5108,N_4030,N_4400);
or U5109 (N_5109,N_4966,N_4736);
nor U5110 (N_5110,N_4876,N_4706);
nand U5111 (N_5111,N_4725,N_4182);
or U5112 (N_5112,N_4274,N_4731);
nor U5113 (N_5113,N_4033,N_4127);
nand U5114 (N_5114,N_4607,N_4992);
or U5115 (N_5115,N_4528,N_4957);
nand U5116 (N_5116,N_4168,N_4660);
or U5117 (N_5117,N_4411,N_4339);
and U5118 (N_5118,N_4655,N_4118);
xor U5119 (N_5119,N_4573,N_4859);
or U5120 (N_5120,N_4602,N_4414);
nand U5121 (N_5121,N_4161,N_4457);
xnor U5122 (N_5122,N_4021,N_4702);
or U5123 (N_5123,N_4460,N_4135);
nor U5124 (N_5124,N_4842,N_4192);
xnor U5125 (N_5125,N_4507,N_4568);
or U5126 (N_5126,N_4890,N_4228);
and U5127 (N_5127,N_4405,N_4235);
nor U5128 (N_5128,N_4906,N_4741);
and U5129 (N_5129,N_4698,N_4156);
nand U5130 (N_5130,N_4211,N_4631);
and U5131 (N_5131,N_4040,N_4011);
nand U5132 (N_5132,N_4378,N_4997);
or U5133 (N_5133,N_4429,N_4467);
or U5134 (N_5134,N_4793,N_4899);
nand U5135 (N_5135,N_4882,N_4348);
or U5136 (N_5136,N_4171,N_4104);
and U5137 (N_5137,N_4347,N_4609);
xor U5138 (N_5138,N_4752,N_4689);
or U5139 (N_5139,N_4031,N_4630);
and U5140 (N_5140,N_4716,N_4903);
and U5141 (N_5141,N_4365,N_4595);
and U5142 (N_5142,N_4340,N_4225);
or U5143 (N_5143,N_4835,N_4693);
nand U5144 (N_5144,N_4301,N_4492);
nor U5145 (N_5145,N_4247,N_4259);
and U5146 (N_5146,N_4481,N_4311);
nor U5147 (N_5147,N_4581,N_4136);
nor U5148 (N_5148,N_4117,N_4187);
or U5149 (N_5149,N_4485,N_4162);
xor U5150 (N_5150,N_4972,N_4814);
or U5151 (N_5151,N_4871,N_4748);
xnor U5152 (N_5152,N_4337,N_4815);
xnor U5153 (N_5153,N_4483,N_4262);
xnor U5154 (N_5154,N_4229,N_4283);
xor U5155 (N_5155,N_4512,N_4811);
nor U5156 (N_5156,N_4372,N_4665);
nand U5157 (N_5157,N_4214,N_4734);
and U5158 (N_5158,N_4165,N_4991);
xnor U5159 (N_5159,N_4745,N_4709);
or U5160 (N_5160,N_4934,N_4190);
and U5161 (N_5161,N_4526,N_4331);
nor U5162 (N_5162,N_4035,N_4000);
xor U5163 (N_5163,N_4921,N_4231);
or U5164 (N_5164,N_4985,N_4812);
and U5165 (N_5165,N_4769,N_4624);
and U5166 (N_5166,N_4565,N_4763);
nor U5167 (N_5167,N_4787,N_4077);
or U5168 (N_5168,N_4611,N_4821);
nand U5169 (N_5169,N_4765,N_4503);
nor U5170 (N_5170,N_4962,N_4278);
or U5171 (N_5171,N_4556,N_4855);
nor U5172 (N_5172,N_4831,N_4236);
nor U5173 (N_5173,N_4625,N_4712);
or U5174 (N_5174,N_4729,N_4329);
or U5175 (N_5175,N_4608,N_4399);
nor U5176 (N_5176,N_4860,N_4408);
and U5177 (N_5177,N_4290,N_4501);
xor U5178 (N_5178,N_4105,N_4264);
and U5179 (N_5179,N_4132,N_4475);
or U5180 (N_5180,N_4241,N_4195);
and U5181 (N_5181,N_4490,N_4172);
or U5182 (N_5182,N_4453,N_4251);
and U5183 (N_5183,N_4002,N_4907);
or U5184 (N_5184,N_4101,N_4059);
nor U5185 (N_5185,N_4515,N_4455);
or U5186 (N_5186,N_4207,N_4677);
or U5187 (N_5187,N_4066,N_4244);
nand U5188 (N_5188,N_4125,N_4647);
xnor U5189 (N_5189,N_4759,N_4005);
and U5190 (N_5190,N_4697,N_4420);
or U5191 (N_5191,N_4439,N_4477);
nor U5192 (N_5192,N_4661,N_4407);
or U5193 (N_5193,N_4544,N_4152);
xnor U5194 (N_5194,N_4468,N_4548);
nand U5195 (N_5195,N_4854,N_4484);
or U5196 (N_5196,N_4242,N_4604);
xor U5197 (N_5197,N_4163,N_4949);
and U5198 (N_5198,N_4374,N_4415);
nand U5199 (N_5199,N_4670,N_4315);
nand U5200 (N_5200,N_4635,N_4367);
or U5201 (N_5201,N_4621,N_4542);
or U5202 (N_5202,N_4916,N_4754);
or U5203 (N_5203,N_4760,N_4428);
or U5204 (N_5204,N_4284,N_4786);
nand U5205 (N_5205,N_4394,N_4213);
or U5206 (N_5206,N_4690,N_4517);
nor U5207 (N_5207,N_4761,N_4965);
or U5208 (N_5208,N_4967,N_4832);
and U5209 (N_5209,N_4513,N_4326);
xor U5210 (N_5210,N_4551,N_4519);
nand U5211 (N_5211,N_4742,N_4788);
and U5212 (N_5212,N_4286,N_4034);
or U5213 (N_5213,N_4224,N_4416);
or U5214 (N_5214,N_4574,N_4464);
xnor U5215 (N_5215,N_4946,N_4092);
xor U5216 (N_5216,N_4801,N_4606);
xnor U5217 (N_5217,N_4888,N_4252);
xnor U5218 (N_5218,N_4114,N_4851);
nand U5219 (N_5219,N_4221,N_4099);
xnor U5220 (N_5220,N_4778,N_4361);
nand U5221 (N_5221,N_4085,N_4605);
xnor U5222 (N_5222,N_4371,N_4923);
and U5223 (N_5223,N_4810,N_4790);
and U5224 (N_5224,N_4710,N_4829);
nand U5225 (N_5225,N_4281,N_4913);
nor U5226 (N_5226,N_4065,N_4462);
or U5227 (N_5227,N_4064,N_4673);
nor U5228 (N_5228,N_4216,N_4246);
and U5229 (N_5229,N_4896,N_4849);
xnor U5230 (N_5230,N_4516,N_4184);
xnor U5231 (N_5231,N_4531,N_4728);
nor U5232 (N_5232,N_4908,N_4634);
xor U5233 (N_5233,N_4711,N_4558);
or U5234 (N_5234,N_4757,N_4930);
or U5235 (N_5235,N_4952,N_4719);
or U5236 (N_5236,N_4557,N_4028);
nor U5237 (N_5237,N_4864,N_4646);
nand U5238 (N_5238,N_4344,N_4198);
and U5239 (N_5239,N_4767,N_4538);
and U5240 (N_5240,N_4784,N_4857);
or U5241 (N_5241,N_4525,N_4324);
nand U5242 (N_5242,N_4079,N_4586);
nor U5243 (N_5243,N_4437,N_4387);
nor U5244 (N_5244,N_4073,N_4576);
nor U5245 (N_5245,N_4904,N_4095);
nor U5246 (N_5246,N_4076,N_4222);
and U5247 (N_5247,N_4657,N_4450);
nand U5248 (N_5248,N_4575,N_4413);
nor U5249 (N_5249,N_4261,N_4298);
or U5250 (N_5250,N_4980,N_4045);
and U5251 (N_5251,N_4258,N_4425);
xor U5252 (N_5252,N_4836,N_4470);
or U5253 (N_5253,N_4561,N_4686);
nand U5254 (N_5254,N_4323,N_4808);
or U5255 (N_5255,N_4383,N_4695);
or U5256 (N_5256,N_4813,N_4537);
xnor U5257 (N_5257,N_4058,N_4253);
and U5258 (N_5258,N_4780,N_4498);
xnor U5259 (N_5259,N_4044,N_4865);
nand U5260 (N_5260,N_4717,N_4392);
nand U5261 (N_5261,N_4699,N_4417);
nor U5262 (N_5262,N_4587,N_4886);
nand U5263 (N_5263,N_4421,N_4194);
nand U5264 (N_5264,N_4375,N_4174);
xor U5265 (N_5265,N_4626,N_4974);
xor U5266 (N_5266,N_4639,N_4732);
nand U5267 (N_5267,N_4335,N_4230);
xnor U5268 (N_5268,N_4273,N_4700);
nand U5269 (N_5269,N_4426,N_4359);
and U5270 (N_5270,N_4446,N_4995);
or U5271 (N_5271,N_4268,N_4920);
nor U5272 (N_5272,N_4047,N_4391);
or U5273 (N_5273,N_4317,N_4691);
xnor U5274 (N_5274,N_4616,N_4072);
and U5275 (N_5275,N_4305,N_4789);
xnor U5276 (N_5276,N_4204,N_4063);
or U5277 (N_5277,N_4902,N_4433);
xnor U5278 (N_5278,N_4128,N_4310);
nand U5279 (N_5279,N_4178,N_4600);
nor U5280 (N_5280,N_4940,N_4203);
or U5281 (N_5281,N_4848,N_4185);
and U5282 (N_5282,N_4215,N_4520);
xor U5283 (N_5283,N_4297,N_4772);
nor U5284 (N_5284,N_4472,N_4422);
nand U5285 (N_5285,N_4785,N_4540);
nor U5286 (N_5286,N_4638,N_4672);
xor U5287 (N_5287,N_4549,N_4622);
xnor U5288 (N_5288,N_4958,N_4071);
nor U5289 (N_5289,N_4202,N_4658);
xnor U5290 (N_5290,N_4115,N_4720);
nor U5291 (N_5291,N_4254,N_4656);
nor U5292 (N_5292,N_4680,N_4889);
nor U5293 (N_5293,N_4108,N_4139);
and U5294 (N_5294,N_4032,N_4678);
and U5295 (N_5295,N_4048,N_4436);
and U5296 (N_5296,N_4328,N_4078);
or U5297 (N_5297,N_4291,N_4692);
or U5298 (N_5298,N_4379,N_4083);
xnor U5299 (N_5299,N_4893,N_4938);
or U5300 (N_5300,N_4679,N_4352);
and U5301 (N_5301,N_4018,N_4166);
nor U5302 (N_5302,N_4758,N_4508);
nor U5303 (N_5303,N_4150,N_4552);
nand U5304 (N_5304,N_4496,N_4091);
nor U5305 (N_5305,N_4943,N_4289);
and U5306 (N_5306,N_4056,N_4826);
and U5307 (N_5307,N_4444,N_4590);
nor U5308 (N_5308,N_4919,N_4341);
xor U5309 (N_5309,N_4333,N_4293);
or U5310 (N_5310,N_4314,N_4279);
nand U5311 (N_5311,N_4448,N_4088);
and U5312 (N_5312,N_4739,N_4743);
and U5313 (N_5313,N_4160,N_4794);
or U5314 (N_5314,N_4316,N_4449);
nand U5315 (N_5315,N_4905,N_4017);
nand U5316 (N_5316,N_4937,N_4232);
and U5317 (N_5317,N_4322,N_4866);
nand U5318 (N_5318,N_4465,N_4764);
xnor U5319 (N_5319,N_4914,N_4385);
or U5320 (N_5320,N_4173,N_4362);
or U5321 (N_5321,N_4456,N_4901);
xnor U5322 (N_5322,N_4004,N_4435);
or U5323 (N_5323,N_4196,N_4942);
and U5324 (N_5324,N_4434,N_4441);
and U5325 (N_5325,N_4023,N_4388);
xor U5326 (N_5326,N_4189,N_4724);
and U5327 (N_5327,N_4559,N_4300);
nor U5328 (N_5328,N_4302,N_4062);
nor U5329 (N_5329,N_4098,N_4102);
or U5330 (N_5330,N_4037,N_4628);
and U5331 (N_5331,N_4653,N_4933);
and U5332 (N_5332,N_4303,N_4588);
xor U5333 (N_5333,N_4238,N_4493);
xnor U5334 (N_5334,N_4954,N_4594);
nand U5335 (N_5335,N_4986,N_4797);
nand U5336 (N_5336,N_4928,N_4955);
and U5337 (N_5337,N_4272,N_4959);
nor U5338 (N_5338,N_4872,N_4012);
nand U5339 (N_5339,N_4746,N_4360);
nand U5340 (N_5340,N_4792,N_4931);
and U5341 (N_5341,N_4113,N_4833);
xor U5342 (N_5342,N_4929,N_4989);
nor U5343 (N_5343,N_4461,N_4255);
xor U5344 (N_5344,N_4683,N_4601);
xor U5345 (N_5345,N_4768,N_4926);
nand U5346 (N_5346,N_4577,N_4834);
or U5347 (N_5347,N_4313,N_4841);
and U5348 (N_5348,N_4119,N_4338);
nand U5349 (N_5349,N_4245,N_4775);
nand U5350 (N_5350,N_4248,N_4535);
xor U5351 (N_5351,N_4038,N_4703);
or U5352 (N_5352,N_4950,N_4180);
or U5353 (N_5353,N_4945,N_4478);
and U5354 (N_5354,N_4523,N_4363);
nor U5355 (N_5355,N_4824,N_4541);
nor U5356 (N_5356,N_4390,N_4327);
nand U5357 (N_5357,N_4791,N_4124);
nand U5358 (N_5358,N_4342,N_4206);
and U5359 (N_5359,N_4850,N_4055);
or U5360 (N_5360,N_4915,N_4081);
nor U5361 (N_5361,N_4880,N_4024);
and U5362 (N_5362,N_4007,N_4911);
nand U5363 (N_5363,N_4632,N_4805);
xor U5364 (N_5364,N_4612,N_4514);
or U5365 (N_5365,N_4107,N_4427);
and U5366 (N_5366,N_4718,N_4469);
nand U5367 (N_5367,N_4990,N_4445);
and U5368 (N_5368,N_4977,N_4186);
nor U5369 (N_5369,N_4144,N_4529);
xnor U5370 (N_5370,N_4026,N_4705);
or U5371 (N_5371,N_4381,N_4662);
xor U5372 (N_5372,N_4082,N_4580);
and U5373 (N_5373,N_4053,N_4084);
or U5374 (N_5374,N_4285,N_4380);
nand U5375 (N_5375,N_4321,N_4069);
or U5376 (N_5376,N_4998,N_4521);
xor U5377 (N_5377,N_4419,N_4130);
and U5378 (N_5378,N_4856,N_4994);
and U5379 (N_5379,N_4721,N_4727);
xor U5380 (N_5380,N_4636,N_4008);
nand U5381 (N_5381,N_4410,N_4582);
or U5382 (N_5382,N_4089,N_4676);
nor U5383 (N_5383,N_4271,N_4862);
or U5384 (N_5384,N_4975,N_4674);
or U5385 (N_5385,N_4193,N_4951);
nand U5386 (N_5386,N_4853,N_4319);
nor U5387 (N_5387,N_4154,N_4153);
or U5388 (N_5388,N_4837,N_4280);
nand U5389 (N_5389,N_4898,N_4209);
xor U5390 (N_5390,N_4935,N_4620);
nor U5391 (N_5391,N_4067,N_4068);
and U5392 (N_5392,N_4840,N_4843);
nor U5393 (N_5393,N_4649,N_4776);
and U5394 (N_5394,N_4423,N_4779);
xnor U5395 (N_5395,N_4825,N_4351);
or U5396 (N_5396,N_4968,N_4020);
and U5397 (N_5397,N_4257,N_4364);
xnor U5398 (N_5398,N_4013,N_4440);
xor U5399 (N_5399,N_4533,N_4599);
and U5400 (N_5400,N_4249,N_4960);
xor U5401 (N_5401,N_4491,N_4015);
nor U5402 (N_5402,N_4309,N_4969);
and U5403 (N_5403,N_4227,N_4292);
nor U5404 (N_5404,N_4343,N_4057);
nor U5405 (N_5405,N_4308,N_4143);
nand U5406 (N_5406,N_4800,N_4640);
nand U5407 (N_5407,N_4641,N_4191);
nor U5408 (N_5408,N_4218,N_4489);
nor U5409 (N_5409,N_4087,N_4179);
xor U5410 (N_5410,N_4159,N_4884);
xor U5411 (N_5411,N_4722,N_4121);
nand U5412 (N_5412,N_4358,N_4663);
nor U5413 (N_5413,N_4807,N_4675);
nor U5414 (N_5414,N_4751,N_4694);
xnor U5415 (N_5415,N_4499,N_4412);
or U5416 (N_5416,N_4155,N_4277);
nor U5417 (N_5417,N_4205,N_4878);
xor U5418 (N_5418,N_4131,N_4750);
and U5419 (N_5419,N_4424,N_4471);
xor U5420 (N_5420,N_4978,N_4643);
nor U5421 (N_5421,N_4263,N_4614);
or U5422 (N_5422,N_4167,N_4895);
or U5423 (N_5423,N_4370,N_4120);
nand U5424 (N_5424,N_4299,N_4458);
nor U5425 (N_5425,N_4562,N_4336);
nor U5426 (N_5426,N_4129,N_4543);
nor U5427 (N_5427,N_4547,N_4603);
nor U5428 (N_5428,N_4487,N_4669);
nor U5429 (N_5429,N_4715,N_4074);
xor U5430 (N_5430,N_4312,N_4142);
or U5431 (N_5431,N_4208,N_4524);
or U5432 (N_5432,N_4738,N_4963);
nand U5433 (N_5433,N_4877,N_4900);
or U5434 (N_5434,N_4567,N_4027);
or U5435 (N_5435,N_4918,N_4782);
nand U5436 (N_5436,N_4701,N_4296);
nand U5437 (N_5437,N_4897,N_4650);
and U5438 (N_5438,N_4885,N_4240);
nor U5439 (N_5439,N_4530,N_4560);
nand U5440 (N_5440,N_4443,N_4723);
nor U5441 (N_5441,N_4671,N_4046);
nand U5442 (N_5442,N_4403,N_4874);
nand U5443 (N_5443,N_4922,N_4584);
xnor U5444 (N_5444,N_4828,N_4527);
xnor U5445 (N_5445,N_4170,N_4287);
nor U5446 (N_5446,N_4522,N_4042);
nor U5447 (N_5447,N_4145,N_4488);
or U5448 (N_5448,N_4645,N_4116);
xnor U5449 (N_5449,N_4953,N_4041);
nand U5450 (N_5450,N_4096,N_4570);
nand U5451 (N_5451,N_4164,N_4648);
nand U5452 (N_5452,N_4973,N_4494);
nor U5453 (N_5453,N_4140,N_4070);
or U5454 (N_5454,N_4382,N_4571);
xnor U5455 (N_5455,N_4438,N_4109);
or U5456 (N_5456,N_4844,N_4536);
or U5457 (N_5457,N_4010,N_4644);
xor U5458 (N_5458,N_4133,N_4912);
xnor U5459 (N_5459,N_4894,N_4398);
or U5460 (N_5460,N_4269,N_4086);
or U5461 (N_5461,N_4774,N_4442);
and U5462 (N_5462,N_4891,N_4936);
or U5463 (N_5463,N_4110,N_4019);
and U5464 (N_5464,N_4875,N_4613);
nor U5465 (N_5465,N_4970,N_4927);
or U5466 (N_5466,N_4147,N_4863);
xor U5467 (N_5467,N_4868,N_4803);
or U5468 (N_5468,N_4502,N_4181);
xor U5469 (N_5469,N_4217,N_4369);
nor U5470 (N_5470,N_4250,N_4892);
nand U5471 (N_5471,N_4288,N_4103);
or U5472 (N_5472,N_4572,N_4629);
xor U5473 (N_5473,N_4052,N_4357);
nand U5474 (N_5474,N_4941,N_4909);
nand U5475 (N_5475,N_4373,N_4947);
and U5476 (N_5476,N_4747,N_4781);
xor U5477 (N_5477,N_4996,N_4265);
or U5478 (N_5478,N_4080,N_4707);
and U5479 (N_5479,N_4334,N_4979);
nand U5480 (N_5480,N_4668,N_4111);
xnor U5481 (N_5481,N_4511,N_4097);
nor U5482 (N_5482,N_4713,N_4226);
and U5483 (N_5483,N_4112,N_4151);
and U5484 (N_5484,N_4591,N_4887);
or U5485 (N_5485,N_4051,N_4999);
nor U5486 (N_5486,N_4169,N_4961);
xor U5487 (N_5487,N_4451,N_4009);
nor U5488 (N_5488,N_4432,N_4157);
nand U5489 (N_5489,N_4749,N_4122);
nand U5490 (N_5490,N_4093,N_4619);
xor U5491 (N_5491,N_4578,N_4726);
or U5492 (N_5492,N_4318,N_4402);
xnor U5493 (N_5493,N_4148,N_4554);
nor U5494 (N_5494,N_4223,N_4592);
nor U5495 (N_5495,N_4566,N_4610);
and U5496 (N_5496,N_4839,N_4744);
xnor U5497 (N_5497,N_4816,N_4495);
or U5498 (N_5498,N_4486,N_4366);
or U5499 (N_5499,N_4737,N_4593);
xnor U5500 (N_5500,N_4318,N_4771);
and U5501 (N_5501,N_4918,N_4431);
nand U5502 (N_5502,N_4864,N_4042);
and U5503 (N_5503,N_4525,N_4597);
xnor U5504 (N_5504,N_4212,N_4432);
xnor U5505 (N_5505,N_4154,N_4263);
xnor U5506 (N_5506,N_4426,N_4543);
or U5507 (N_5507,N_4654,N_4396);
xor U5508 (N_5508,N_4745,N_4555);
nor U5509 (N_5509,N_4563,N_4808);
xnor U5510 (N_5510,N_4081,N_4467);
and U5511 (N_5511,N_4871,N_4882);
nand U5512 (N_5512,N_4776,N_4047);
or U5513 (N_5513,N_4374,N_4273);
xnor U5514 (N_5514,N_4376,N_4696);
and U5515 (N_5515,N_4349,N_4034);
and U5516 (N_5516,N_4091,N_4523);
nand U5517 (N_5517,N_4996,N_4962);
nor U5518 (N_5518,N_4189,N_4558);
nor U5519 (N_5519,N_4746,N_4289);
or U5520 (N_5520,N_4703,N_4600);
and U5521 (N_5521,N_4406,N_4807);
or U5522 (N_5522,N_4417,N_4206);
nand U5523 (N_5523,N_4061,N_4649);
and U5524 (N_5524,N_4760,N_4682);
xnor U5525 (N_5525,N_4612,N_4292);
nand U5526 (N_5526,N_4927,N_4835);
nand U5527 (N_5527,N_4518,N_4572);
xnor U5528 (N_5528,N_4914,N_4477);
nor U5529 (N_5529,N_4935,N_4443);
nand U5530 (N_5530,N_4891,N_4419);
nand U5531 (N_5531,N_4594,N_4209);
and U5532 (N_5532,N_4459,N_4201);
and U5533 (N_5533,N_4081,N_4859);
xnor U5534 (N_5534,N_4963,N_4374);
or U5535 (N_5535,N_4032,N_4639);
nand U5536 (N_5536,N_4753,N_4907);
and U5537 (N_5537,N_4249,N_4467);
nor U5538 (N_5538,N_4007,N_4208);
xor U5539 (N_5539,N_4241,N_4042);
nand U5540 (N_5540,N_4321,N_4922);
xor U5541 (N_5541,N_4107,N_4202);
and U5542 (N_5542,N_4112,N_4554);
and U5543 (N_5543,N_4714,N_4014);
or U5544 (N_5544,N_4425,N_4900);
nor U5545 (N_5545,N_4681,N_4582);
or U5546 (N_5546,N_4001,N_4820);
nor U5547 (N_5547,N_4553,N_4666);
nand U5548 (N_5548,N_4943,N_4841);
or U5549 (N_5549,N_4610,N_4365);
or U5550 (N_5550,N_4178,N_4729);
nor U5551 (N_5551,N_4482,N_4944);
or U5552 (N_5552,N_4936,N_4303);
nand U5553 (N_5553,N_4578,N_4888);
xor U5554 (N_5554,N_4522,N_4965);
nand U5555 (N_5555,N_4710,N_4665);
and U5556 (N_5556,N_4560,N_4877);
nand U5557 (N_5557,N_4891,N_4548);
or U5558 (N_5558,N_4111,N_4316);
nand U5559 (N_5559,N_4876,N_4764);
nand U5560 (N_5560,N_4148,N_4324);
or U5561 (N_5561,N_4975,N_4814);
and U5562 (N_5562,N_4832,N_4926);
and U5563 (N_5563,N_4777,N_4471);
nor U5564 (N_5564,N_4851,N_4941);
xor U5565 (N_5565,N_4996,N_4032);
and U5566 (N_5566,N_4353,N_4029);
and U5567 (N_5567,N_4050,N_4844);
xor U5568 (N_5568,N_4479,N_4064);
nand U5569 (N_5569,N_4683,N_4603);
xor U5570 (N_5570,N_4827,N_4726);
nor U5571 (N_5571,N_4818,N_4552);
nand U5572 (N_5572,N_4966,N_4558);
and U5573 (N_5573,N_4164,N_4383);
nor U5574 (N_5574,N_4693,N_4076);
or U5575 (N_5575,N_4764,N_4654);
or U5576 (N_5576,N_4411,N_4367);
nor U5577 (N_5577,N_4604,N_4963);
nor U5578 (N_5578,N_4692,N_4549);
or U5579 (N_5579,N_4564,N_4424);
and U5580 (N_5580,N_4429,N_4274);
nor U5581 (N_5581,N_4919,N_4878);
xnor U5582 (N_5582,N_4819,N_4217);
xor U5583 (N_5583,N_4528,N_4663);
xor U5584 (N_5584,N_4999,N_4858);
or U5585 (N_5585,N_4063,N_4185);
and U5586 (N_5586,N_4692,N_4196);
nand U5587 (N_5587,N_4508,N_4931);
nor U5588 (N_5588,N_4167,N_4610);
and U5589 (N_5589,N_4062,N_4030);
and U5590 (N_5590,N_4603,N_4613);
or U5591 (N_5591,N_4671,N_4770);
nor U5592 (N_5592,N_4330,N_4183);
xor U5593 (N_5593,N_4844,N_4231);
and U5594 (N_5594,N_4923,N_4737);
and U5595 (N_5595,N_4582,N_4851);
nand U5596 (N_5596,N_4762,N_4123);
nand U5597 (N_5597,N_4614,N_4082);
or U5598 (N_5598,N_4742,N_4389);
nand U5599 (N_5599,N_4719,N_4663);
or U5600 (N_5600,N_4438,N_4550);
xnor U5601 (N_5601,N_4250,N_4081);
and U5602 (N_5602,N_4808,N_4930);
nor U5603 (N_5603,N_4513,N_4811);
xnor U5604 (N_5604,N_4094,N_4304);
nor U5605 (N_5605,N_4280,N_4464);
nand U5606 (N_5606,N_4665,N_4371);
and U5607 (N_5607,N_4272,N_4503);
nor U5608 (N_5608,N_4102,N_4081);
xor U5609 (N_5609,N_4569,N_4499);
or U5610 (N_5610,N_4677,N_4251);
or U5611 (N_5611,N_4152,N_4169);
nand U5612 (N_5612,N_4502,N_4471);
or U5613 (N_5613,N_4894,N_4986);
xor U5614 (N_5614,N_4091,N_4796);
or U5615 (N_5615,N_4208,N_4246);
xor U5616 (N_5616,N_4576,N_4542);
and U5617 (N_5617,N_4195,N_4857);
nand U5618 (N_5618,N_4471,N_4993);
nor U5619 (N_5619,N_4159,N_4942);
xor U5620 (N_5620,N_4650,N_4585);
or U5621 (N_5621,N_4866,N_4282);
xnor U5622 (N_5622,N_4124,N_4962);
nand U5623 (N_5623,N_4231,N_4837);
xnor U5624 (N_5624,N_4094,N_4390);
nand U5625 (N_5625,N_4557,N_4610);
xnor U5626 (N_5626,N_4421,N_4913);
or U5627 (N_5627,N_4326,N_4987);
and U5628 (N_5628,N_4521,N_4287);
xnor U5629 (N_5629,N_4038,N_4137);
or U5630 (N_5630,N_4307,N_4546);
nand U5631 (N_5631,N_4693,N_4615);
nand U5632 (N_5632,N_4880,N_4729);
xor U5633 (N_5633,N_4910,N_4234);
or U5634 (N_5634,N_4899,N_4990);
xnor U5635 (N_5635,N_4692,N_4996);
nand U5636 (N_5636,N_4097,N_4387);
or U5637 (N_5637,N_4021,N_4475);
xor U5638 (N_5638,N_4558,N_4129);
or U5639 (N_5639,N_4519,N_4184);
and U5640 (N_5640,N_4680,N_4036);
nand U5641 (N_5641,N_4621,N_4261);
nor U5642 (N_5642,N_4891,N_4473);
and U5643 (N_5643,N_4087,N_4641);
and U5644 (N_5644,N_4083,N_4213);
and U5645 (N_5645,N_4818,N_4073);
nand U5646 (N_5646,N_4037,N_4722);
or U5647 (N_5647,N_4692,N_4126);
or U5648 (N_5648,N_4669,N_4591);
xnor U5649 (N_5649,N_4139,N_4272);
nor U5650 (N_5650,N_4352,N_4116);
and U5651 (N_5651,N_4366,N_4991);
nor U5652 (N_5652,N_4901,N_4598);
nand U5653 (N_5653,N_4795,N_4258);
or U5654 (N_5654,N_4994,N_4687);
or U5655 (N_5655,N_4599,N_4304);
nand U5656 (N_5656,N_4900,N_4634);
nor U5657 (N_5657,N_4770,N_4319);
xor U5658 (N_5658,N_4892,N_4159);
or U5659 (N_5659,N_4949,N_4220);
and U5660 (N_5660,N_4013,N_4770);
nand U5661 (N_5661,N_4041,N_4989);
and U5662 (N_5662,N_4568,N_4506);
nor U5663 (N_5663,N_4891,N_4392);
and U5664 (N_5664,N_4573,N_4357);
xor U5665 (N_5665,N_4386,N_4355);
xnor U5666 (N_5666,N_4997,N_4807);
nand U5667 (N_5667,N_4894,N_4679);
and U5668 (N_5668,N_4380,N_4064);
and U5669 (N_5669,N_4674,N_4760);
or U5670 (N_5670,N_4603,N_4101);
xnor U5671 (N_5671,N_4759,N_4586);
nand U5672 (N_5672,N_4379,N_4017);
or U5673 (N_5673,N_4132,N_4918);
xnor U5674 (N_5674,N_4430,N_4625);
and U5675 (N_5675,N_4970,N_4294);
and U5676 (N_5676,N_4313,N_4562);
xor U5677 (N_5677,N_4941,N_4773);
nor U5678 (N_5678,N_4570,N_4268);
and U5679 (N_5679,N_4939,N_4936);
nor U5680 (N_5680,N_4604,N_4628);
xor U5681 (N_5681,N_4826,N_4270);
xnor U5682 (N_5682,N_4981,N_4731);
xnor U5683 (N_5683,N_4454,N_4000);
and U5684 (N_5684,N_4161,N_4249);
nand U5685 (N_5685,N_4543,N_4008);
or U5686 (N_5686,N_4277,N_4262);
nand U5687 (N_5687,N_4864,N_4743);
nand U5688 (N_5688,N_4830,N_4707);
and U5689 (N_5689,N_4896,N_4123);
nand U5690 (N_5690,N_4533,N_4581);
nor U5691 (N_5691,N_4622,N_4930);
nand U5692 (N_5692,N_4288,N_4048);
xnor U5693 (N_5693,N_4822,N_4830);
and U5694 (N_5694,N_4719,N_4411);
nand U5695 (N_5695,N_4261,N_4882);
xor U5696 (N_5696,N_4374,N_4558);
xnor U5697 (N_5697,N_4598,N_4822);
and U5698 (N_5698,N_4743,N_4066);
and U5699 (N_5699,N_4111,N_4121);
nand U5700 (N_5700,N_4770,N_4078);
nand U5701 (N_5701,N_4312,N_4699);
or U5702 (N_5702,N_4448,N_4886);
nor U5703 (N_5703,N_4335,N_4982);
and U5704 (N_5704,N_4219,N_4517);
nor U5705 (N_5705,N_4692,N_4509);
xnor U5706 (N_5706,N_4802,N_4252);
xnor U5707 (N_5707,N_4846,N_4525);
and U5708 (N_5708,N_4310,N_4166);
nor U5709 (N_5709,N_4811,N_4681);
nor U5710 (N_5710,N_4047,N_4211);
xor U5711 (N_5711,N_4635,N_4869);
xnor U5712 (N_5712,N_4290,N_4929);
nor U5713 (N_5713,N_4567,N_4247);
and U5714 (N_5714,N_4874,N_4370);
xnor U5715 (N_5715,N_4526,N_4715);
and U5716 (N_5716,N_4626,N_4813);
and U5717 (N_5717,N_4230,N_4896);
or U5718 (N_5718,N_4625,N_4698);
or U5719 (N_5719,N_4335,N_4562);
nand U5720 (N_5720,N_4736,N_4441);
nor U5721 (N_5721,N_4811,N_4311);
or U5722 (N_5722,N_4416,N_4653);
and U5723 (N_5723,N_4881,N_4168);
xor U5724 (N_5724,N_4058,N_4966);
or U5725 (N_5725,N_4380,N_4605);
and U5726 (N_5726,N_4505,N_4344);
xnor U5727 (N_5727,N_4937,N_4335);
xor U5728 (N_5728,N_4450,N_4361);
nand U5729 (N_5729,N_4744,N_4464);
nor U5730 (N_5730,N_4245,N_4089);
xor U5731 (N_5731,N_4680,N_4454);
xor U5732 (N_5732,N_4018,N_4659);
nand U5733 (N_5733,N_4687,N_4439);
and U5734 (N_5734,N_4937,N_4402);
nand U5735 (N_5735,N_4575,N_4746);
or U5736 (N_5736,N_4528,N_4694);
nand U5737 (N_5737,N_4462,N_4760);
nand U5738 (N_5738,N_4620,N_4173);
and U5739 (N_5739,N_4778,N_4926);
xnor U5740 (N_5740,N_4356,N_4939);
or U5741 (N_5741,N_4991,N_4628);
nor U5742 (N_5742,N_4541,N_4128);
xnor U5743 (N_5743,N_4378,N_4931);
xor U5744 (N_5744,N_4443,N_4875);
nand U5745 (N_5745,N_4387,N_4829);
or U5746 (N_5746,N_4578,N_4380);
xnor U5747 (N_5747,N_4216,N_4574);
xor U5748 (N_5748,N_4143,N_4362);
and U5749 (N_5749,N_4015,N_4570);
and U5750 (N_5750,N_4699,N_4188);
xor U5751 (N_5751,N_4369,N_4777);
or U5752 (N_5752,N_4384,N_4295);
xnor U5753 (N_5753,N_4236,N_4436);
or U5754 (N_5754,N_4754,N_4868);
nand U5755 (N_5755,N_4745,N_4225);
and U5756 (N_5756,N_4342,N_4326);
and U5757 (N_5757,N_4394,N_4630);
xnor U5758 (N_5758,N_4016,N_4977);
nor U5759 (N_5759,N_4124,N_4829);
or U5760 (N_5760,N_4893,N_4161);
or U5761 (N_5761,N_4996,N_4269);
nor U5762 (N_5762,N_4913,N_4171);
nor U5763 (N_5763,N_4850,N_4150);
nand U5764 (N_5764,N_4082,N_4924);
or U5765 (N_5765,N_4444,N_4091);
xor U5766 (N_5766,N_4238,N_4877);
and U5767 (N_5767,N_4166,N_4842);
or U5768 (N_5768,N_4473,N_4590);
nand U5769 (N_5769,N_4649,N_4385);
nand U5770 (N_5770,N_4495,N_4432);
and U5771 (N_5771,N_4839,N_4105);
or U5772 (N_5772,N_4619,N_4919);
nand U5773 (N_5773,N_4095,N_4217);
and U5774 (N_5774,N_4322,N_4356);
or U5775 (N_5775,N_4116,N_4186);
xor U5776 (N_5776,N_4978,N_4617);
xnor U5777 (N_5777,N_4814,N_4442);
nand U5778 (N_5778,N_4965,N_4752);
xnor U5779 (N_5779,N_4568,N_4380);
and U5780 (N_5780,N_4275,N_4198);
xnor U5781 (N_5781,N_4196,N_4160);
or U5782 (N_5782,N_4083,N_4195);
xnor U5783 (N_5783,N_4306,N_4632);
or U5784 (N_5784,N_4569,N_4060);
xor U5785 (N_5785,N_4095,N_4391);
or U5786 (N_5786,N_4027,N_4778);
xnor U5787 (N_5787,N_4420,N_4920);
nor U5788 (N_5788,N_4547,N_4604);
and U5789 (N_5789,N_4941,N_4189);
or U5790 (N_5790,N_4392,N_4901);
xnor U5791 (N_5791,N_4429,N_4336);
or U5792 (N_5792,N_4589,N_4422);
nand U5793 (N_5793,N_4399,N_4483);
and U5794 (N_5794,N_4219,N_4582);
nand U5795 (N_5795,N_4653,N_4704);
and U5796 (N_5796,N_4101,N_4142);
nor U5797 (N_5797,N_4217,N_4627);
nand U5798 (N_5798,N_4512,N_4802);
nand U5799 (N_5799,N_4821,N_4120);
and U5800 (N_5800,N_4628,N_4567);
or U5801 (N_5801,N_4181,N_4254);
and U5802 (N_5802,N_4632,N_4360);
nor U5803 (N_5803,N_4470,N_4491);
or U5804 (N_5804,N_4894,N_4332);
or U5805 (N_5805,N_4195,N_4457);
xnor U5806 (N_5806,N_4869,N_4634);
and U5807 (N_5807,N_4912,N_4503);
or U5808 (N_5808,N_4740,N_4656);
or U5809 (N_5809,N_4510,N_4980);
xnor U5810 (N_5810,N_4897,N_4299);
xnor U5811 (N_5811,N_4737,N_4120);
nand U5812 (N_5812,N_4430,N_4131);
nor U5813 (N_5813,N_4113,N_4146);
nor U5814 (N_5814,N_4870,N_4164);
or U5815 (N_5815,N_4555,N_4225);
nor U5816 (N_5816,N_4768,N_4367);
xor U5817 (N_5817,N_4973,N_4278);
xor U5818 (N_5818,N_4595,N_4447);
and U5819 (N_5819,N_4973,N_4664);
nor U5820 (N_5820,N_4113,N_4687);
nand U5821 (N_5821,N_4135,N_4915);
nand U5822 (N_5822,N_4342,N_4934);
xnor U5823 (N_5823,N_4112,N_4036);
nand U5824 (N_5824,N_4960,N_4910);
nor U5825 (N_5825,N_4539,N_4829);
nor U5826 (N_5826,N_4516,N_4342);
or U5827 (N_5827,N_4628,N_4760);
and U5828 (N_5828,N_4378,N_4576);
or U5829 (N_5829,N_4970,N_4662);
nor U5830 (N_5830,N_4190,N_4896);
nand U5831 (N_5831,N_4495,N_4505);
or U5832 (N_5832,N_4666,N_4262);
nor U5833 (N_5833,N_4075,N_4619);
or U5834 (N_5834,N_4318,N_4081);
or U5835 (N_5835,N_4115,N_4455);
nor U5836 (N_5836,N_4376,N_4698);
xor U5837 (N_5837,N_4740,N_4842);
nand U5838 (N_5838,N_4332,N_4531);
or U5839 (N_5839,N_4461,N_4261);
and U5840 (N_5840,N_4365,N_4332);
and U5841 (N_5841,N_4511,N_4392);
nor U5842 (N_5842,N_4828,N_4469);
nand U5843 (N_5843,N_4817,N_4006);
and U5844 (N_5844,N_4466,N_4124);
nor U5845 (N_5845,N_4324,N_4516);
nor U5846 (N_5846,N_4072,N_4055);
nor U5847 (N_5847,N_4208,N_4188);
xnor U5848 (N_5848,N_4939,N_4828);
or U5849 (N_5849,N_4754,N_4160);
xor U5850 (N_5850,N_4750,N_4222);
nor U5851 (N_5851,N_4225,N_4139);
nor U5852 (N_5852,N_4567,N_4060);
and U5853 (N_5853,N_4947,N_4074);
and U5854 (N_5854,N_4946,N_4197);
nor U5855 (N_5855,N_4577,N_4502);
and U5856 (N_5856,N_4503,N_4419);
xor U5857 (N_5857,N_4465,N_4964);
nor U5858 (N_5858,N_4621,N_4507);
xor U5859 (N_5859,N_4652,N_4408);
nand U5860 (N_5860,N_4409,N_4656);
xnor U5861 (N_5861,N_4655,N_4451);
xnor U5862 (N_5862,N_4655,N_4458);
nor U5863 (N_5863,N_4463,N_4944);
nand U5864 (N_5864,N_4559,N_4292);
nor U5865 (N_5865,N_4192,N_4559);
xnor U5866 (N_5866,N_4659,N_4156);
or U5867 (N_5867,N_4687,N_4664);
or U5868 (N_5868,N_4833,N_4082);
nor U5869 (N_5869,N_4160,N_4734);
xnor U5870 (N_5870,N_4703,N_4149);
and U5871 (N_5871,N_4426,N_4549);
nand U5872 (N_5872,N_4290,N_4808);
and U5873 (N_5873,N_4193,N_4183);
or U5874 (N_5874,N_4088,N_4456);
nor U5875 (N_5875,N_4366,N_4458);
or U5876 (N_5876,N_4356,N_4117);
nand U5877 (N_5877,N_4277,N_4390);
or U5878 (N_5878,N_4975,N_4741);
and U5879 (N_5879,N_4376,N_4230);
and U5880 (N_5880,N_4223,N_4237);
xnor U5881 (N_5881,N_4589,N_4122);
nand U5882 (N_5882,N_4089,N_4140);
nand U5883 (N_5883,N_4052,N_4783);
and U5884 (N_5884,N_4324,N_4219);
or U5885 (N_5885,N_4208,N_4567);
xnor U5886 (N_5886,N_4443,N_4625);
or U5887 (N_5887,N_4739,N_4486);
xor U5888 (N_5888,N_4860,N_4294);
nand U5889 (N_5889,N_4628,N_4742);
or U5890 (N_5890,N_4638,N_4309);
and U5891 (N_5891,N_4165,N_4952);
nor U5892 (N_5892,N_4203,N_4225);
xor U5893 (N_5893,N_4099,N_4558);
and U5894 (N_5894,N_4320,N_4316);
xor U5895 (N_5895,N_4584,N_4911);
nor U5896 (N_5896,N_4032,N_4232);
and U5897 (N_5897,N_4365,N_4958);
and U5898 (N_5898,N_4937,N_4220);
or U5899 (N_5899,N_4075,N_4621);
and U5900 (N_5900,N_4877,N_4809);
nand U5901 (N_5901,N_4980,N_4015);
nand U5902 (N_5902,N_4044,N_4357);
and U5903 (N_5903,N_4328,N_4278);
nand U5904 (N_5904,N_4300,N_4037);
xnor U5905 (N_5905,N_4229,N_4671);
and U5906 (N_5906,N_4977,N_4825);
or U5907 (N_5907,N_4983,N_4447);
nand U5908 (N_5908,N_4701,N_4048);
and U5909 (N_5909,N_4766,N_4064);
xnor U5910 (N_5910,N_4960,N_4052);
xnor U5911 (N_5911,N_4316,N_4663);
or U5912 (N_5912,N_4721,N_4088);
nor U5913 (N_5913,N_4151,N_4347);
nand U5914 (N_5914,N_4370,N_4463);
and U5915 (N_5915,N_4516,N_4080);
nor U5916 (N_5916,N_4988,N_4736);
nor U5917 (N_5917,N_4970,N_4215);
and U5918 (N_5918,N_4626,N_4319);
and U5919 (N_5919,N_4513,N_4246);
or U5920 (N_5920,N_4315,N_4858);
or U5921 (N_5921,N_4907,N_4932);
or U5922 (N_5922,N_4743,N_4843);
nor U5923 (N_5923,N_4094,N_4365);
nor U5924 (N_5924,N_4468,N_4630);
or U5925 (N_5925,N_4425,N_4439);
nor U5926 (N_5926,N_4805,N_4406);
or U5927 (N_5927,N_4080,N_4380);
nor U5928 (N_5928,N_4068,N_4012);
or U5929 (N_5929,N_4709,N_4864);
nand U5930 (N_5930,N_4020,N_4026);
or U5931 (N_5931,N_4014,N_4423);
or U5932 (N_5932,N_4052,N_4214);
nand U5933 (N_5933,N_4150,N_4204);
nand U5934 (N_5934,N_4764,N_4012);
nor U5935 (N_5935,N_4036,N_4181);
or U5936 (N_5936,N_4675,N_4210);
xor U5937 (N_5937,N_4565,N_4859);
or U5938 (N_5938,N_4954,N_4208);
xor U5939 (N_5939,N_4989,N_4078);
nand U5940 (N_5940,N_4601,N_4463);
or U5941 (N_5941,N_4791,N_4432);
xor U5942 (N_5942,N_4903,N_4629);
or U5943 (N_5943,N_4624,N_4104);
nor U5944 (N_5944,N_4347,N_4350);
xnor U5945 (N_5945,N_4541,N_4732);
xor U5946 (N_5946,N_4143,N_4029);
and U5947 (N_5947,N_4723,N_4390);
nor U5948 (N_5948,N_4786,N_4085);
xnor U5949 (N_5949,N_4871,N_4026);
nand U5950 (N_5950,N_4586,N_4443);
xnor U5951 (N_5951,N_4540,N_4500);
or U5952 (N_5952,N_4953,N_4939);
nor U5953 (N_5953,N_4706,N_4159);
and U5954 (N_5954,N_4710,N_4482);
nor U5955 (N_5955,N_4272,N_4692);
or U5956 (N_5956,N_4510,N_4419);
nor U5957 (N_5957,N_4791,N_4528);
or U5958 (N_5958,N_4151,N_4536);
nand U5959 (N_5959,N_4083,N_4298);
nand U5960 (N_5960,N_4973,N_4360);
or U5961 (N_5961,N_4874,N_4527);
nand U5962 (N_5962,N_4734,N_4929);
nor U5963 (N_5963,N_4674,N_4239);
and U5964 (N_5964,N_4566,N_4167);
and U5965 (N_5965,N_4014,N_4055);
nor U5966 (N_5966,N_4808,N_4058);
and U5967 (N_5967,N_4090,N_4626);
and U5968 (N_5968,N_4601,N_4984);
or U5969 (N_5969,N_4781,N_4273);
nand U5970 (N_5970,N_4151,N_4586);
or U5971 (N_5971,N_4344,N_4416);
nor U5972 (N_5972,N_4176,N_4073);
nand U5973 (N_5973,N_4512,N_4703);
and U5974 (N_5974,N_4547,N_4544);
or U5975 (N_5975,N_4984,N_4896);
and U5976 (N_5976,N_4665,N_4773);
xnor U5977 (N_5977,N_4242,N_4399);
nand U5978 (N_5978,N_4644,N_4258);
or U5979 (N_5979,N_4177,N_4643);
nand U5980 (N_5980,N_4921,N_4830);
nor U5981 (N_5981,N_4793,N_4086);
or U5982 (N_5982,N_4714,N_4613);
xor U5983 (N_5983,N_4567,N_4156);
nor U5984 (N_5984,N_4731,N_4750);
xnor U5985 (N_5985,N_4827,N_4500);
xnor U5986 (N_5986,N_4068,N_4337);
xor U5987 (N_5987,N_4425,N_4896);
nand U5988 (N_5988,N_4940,N_4046);
xnor U5989 (N_5989,N_4112,N_4079);
xor U5990 (N_5990,N_4262,N_4663);
nor U5991 (N_5991,N_4920,N_4010);
nor U5992 (N_5992,N_4974,N_4120);
xnor U5993 (N_5993,N_4076,N_4402);
nand U5994 (N_5994,N_4100,N_4447);
nand U5995 (N_5995,N_4758,N_4830);
nand U5996 (N_5996,N_4131,N_4217);
nand U5997 (N_5997,N_4279,N_4391);
xnor U5998 (N_5998,N_4443,N_4177);
nor U5999 (N_5999,N_4504,N_4032);
nor U6000 (N_6000,N_5790,N_5113);
nand U6001 (N_6001,N_5632,N_5678);
xor U6002 (N_6002,N_5134,N_5718);
and U6003 (N_6003,N_5128,N_5847);
xnor U6004 (N_6004,N_5116,N_5147);
nor U6005 (N_6005,N_5643,N_5644);
or U6006 (N_6006,N_5458,N_5984);
xnor U6007 (N_6007,N_5019,N_5293);
nor U6008 (N_6008,N_5685,N_5303);
or U6009 (N_6009,N_5357,N_5805);
or U6010 (N_6010,N_5951,N_5641);
nor U6011 (N_6011,N_5390,N_5036);
xor U6012 (N_6012,N_5658,N_5075);
nor U6013 (N_6013,N_5343,N_5689);
nor U6014 (N_6014,N_5832,N_5270);
nor U6015 (N_6015,N_5364,N_5345);
nor U6016 (N_6016,N_5577,N_5629);
and U6017 (N_6017,N_5592,N_5513);
or U6018 (N_6018,N_5903,N_5563);
xor U6019 (N_6019,N_5891,N_5415);
or U6020 (N_6020,N_5675,N_5776);
or U6021 (N_6021,N_5500,N_5013);
or U6022 (N_6022,N_5322,N_5898);
xnor U6023 (N_6023,N_5088,N_5107);
nand U6024 (N_6024,N_5872,N_5058);
nor U6025 (N_6025,N_5713,N_5591);
or U6026 (N_6026,N_5759,N_5924);
nand U6027 (N_6027,N_5203,N_5727);
xor U6028 (N_6028,N_5065,N_5835);
xnor U6029 (N_6029,N_5717,N_5647);
nand U6030 (N_6030,N_5138,N_5325);
xnor U6031 (N_6031,N_5876,N_5905);
xor U6032 (N_6032,N_5286,N_5981);
nor U6033 (N_6033,N_5849,N_5761);
nor U6034 (N_6034,N_5318,N_5613);
xor U6035 (N_6035,N_5089,N_5139);
xnor U6036 (N_6036,N_5901,N_5758);
or U6037 (N_6037,N_5086,N_5267);
nor U6038 (N_6038,N_5947,N_5277);
or U6039 (N_6039,N_5460,N_5804);
nor U6040 (N_6040,N_5782,N_5480);
and U6041 (N_6041,N_5608,N_5908);
xor U6042 (N_6042,N_5423,N_5968);
xnor U6043 (N_6043,N_5550,N_5229);
and U6044 (N_6044,N_5998,N_5562);
and U6045 (N_6045,N_5187,N_5186);
or U6046 (N_6046,N_5218,N_5823);
or U6047 (N_6047,N_5320,N_5828);
or U6048 (N_6048,N_5056,N_5929);
and U6049 (N_6049,N_5255,N_5261);
nor U6050 (N_6050,N_5022,N_5389);
nor U6051 (N_6051,N_5911,N_5543);
and U6052 (N_6052,N_5886,N_5475);
or U6053 (N_6053,N_5661,N_5739);
or U6054 (N_6054,N_5774,N_5117);
or U6055 (N_6055,N_5080,N_5416);
nor U6056 (N_6056,N_5413,N_5171);
and U6057 (N_6057,N_5370,N_5939);
or U6058 (N_6058,N_5624,N_5446);
nor U6059 (N_6059,N_5582,N_5795);
xnor U6060 (N_6060,N_5424,N_5940);
and U6061 (N_6061,N_5735,N_5109);
nor U6062 (N_6062,N_5917,N_5972);
nand U6063 (N_6063,N_5983,N_5481);
nor U6064 (N_6064,N_5792,N_5771);
nand U6065 (N_6065,N_5395,N_5596);
xor U6066 (N_6066,N_5800,N_5396);
nor U6067 (N_6067,N_5476,N_5837);
xor U6068 (N_6068,N_5967,N_5544);
nand U6069 (N_6069,N_5944,N_5451);
nand U6070 (N_6070,N_5611,N_5857);
or U6071 (N_6071,N_5173,N_5160);
nor U6072 (N_6072,N_5575,N_5422);
nand U6073 (N_6073,N_5433,N_5851);
and U6074 (N_6074,N_5970,N_5846);
nor U6075 (N_6075,N_5928,N_5031);
nand U6076 (N_6076,N_5786,N_5175);
and U6077 (N_6077,N_5540,N_5992);
nor U6078 (N_6078,N_5214,N_5656);
xor U6079 (N_6079,N_5141,N_5402);
xnor U6080 (N_6080,N_5071,N_5299);
or U6081 (N_6081,N_5617,N_5262);
xnor U6082 (N_6082,N_5266,N_5537);
nand U6083 (N_6083,N_5288,N_5838);
or U6084 (N_6084,N_5765,N_5275);
nor U6085 (N_6085,N_5720,N_5677);
nand U6086 (N_6086,N_5131,N_5378);
xnor U6087 (N_6087,N_5816,N_5140);
nand U6088 (N_6088,N_5397,N_5290);
or U6089 (N_6089,N_5244,N_5174);
and U6090 (N_6090,N_5220,N_5772);
nor U6091 (N_6091,N_5964,N_5406);
and U6092 (N_6092,N_5902,N_5637);
nand U6093 (N_6093,N_5383,N_5887);
nor U6094 (N_6094,N_5646,N_5166);
xnor U6095 (N_6095,N_5309,N_5279);
xnor U6096 (N_6096,N_5826,N_5979);
nor U6097 (N_6097,N_5843,N_5040);
or U6098 (N_6098,N_5512,N_5502);
xor U6099 (N_6099,N_5530,N_5963);
nand U6100 (N_6100,N_5194,N_5606);
nand U6101 (N_6101,N_5009,N_5733);
or U6102 (N_6102,N_5815,N_5457);
or U6103 (N_6103,N_5878,N_5927);
xor U6104 (N_6104,N_5285,N_5912);
nor U6105 (N_6105,N_5007,N_5344);
or U6106 (N_6106,N_5687,N_5976);
nand U6107 (N_6107,N_5148,N_5483);
nor U6108 (N_6108,N_5030,N_5354);
and U6109 (N_6109,N_5111,N_5412);
and U6110 (N_6110,N_5690,N_5841);
nor U6111 (N_6111,N_5260,N_5265);
xor U6112 (N_6112,N_5743,N_5462);
or U6113 (N_6113,N_5788,N_5645);
xor U6114 (N_6114,N_5193,N_5133);
and U6115 (N_6115,N_5163,N_5698);
and U6116 (N_6116,N_5410,N_5503);
nor U6117 (N_6117,N_5149,N_5867);
or U6118 (N_6118,N_5465,N_5315);
nor U6119 (N_6119,N_5338,N_5565);
nand U6120 (N_6120,N_5794,N_5352);
nor U6121 (N_6121,N_5185,N_5329);
xnor U6122 (N_6122,N_5559,N_5313);
nand U6123 (N_6123,N_5292,N_5625);
or U6124 (N_6124,N_5978,N_5877);
nand U6125 (N_6125,N_5797,N_5047);
and U6126 (N_6126,N_5135,N_5479);
xnor U6127 (N_6127,N_5635,N_5369);
nand U6128 (N_6128,N_5538,N_5327);
or U6129 (N_6129,N_5074,N_5312);
nand U6130 (N_6130,N_5861,N_5589);
and U6131 (N_6131,N_5616,N_5232);
or U6132 (N_6132,N_5243,N_5051);
or U6133 (N_6133,N_5361,N_5210);
nand U6134 (N_6134,N_5283,N_5836);
nand U6135 (N_6135,N_5914,N_5524);
and U6136 (N_6136,N_5399,N_5767);
or U6137 (N_6137,N_5226,N_5156);
nor U6138 (N_6138,N_5280,N_5798);
and U6139 (N_6139,N_5568,N_5817);
nand U6140 (N_6140,N_5385,N_5747);
nand U6141 (N_6141,N_5235,N_5558);
nor U6142 (N_6142,N_5862,N_5418);
xnor U6143 (N_6143,N_5623,N_5557);
nor U6144 (N_6144,N_5222,N_5434);
xor U6145 (N_6145,N_5427,N_5291);
or U6146 (N_6146,N_5102,N_5182);
xnor U6147 (N_6147,N_5578,N_5249);
or U6148 (N_6148,N_5556,N_5868);
or U6149 (N_6149,N_5010,N_5554);
and U6150 (N_6150,N_5489,N_5000);
and U6151 (N_6151,N_5494,N_5918);
nand U6152 (N_6152,N_5725,N_5948);
nand U6153 (N_6153,N_5365,N_5549);
and U6154 (N_6154,N_5583,N_5620);
nor U6155 (N_6155,N_5098,N_5337);
and U6156 (N_6156,N_5428,N_5570);
nand U6157 (N_6157,N_5042,N_5848);
xor U6158 (N_6158,N_5411,N_5094);
nor U6159 (N_6159,N_5989,N_5982);
or U6160 (N_6160,N_5707,N_5959);
or U6161 (N_6161,N_5551,N_5899);
nand U6162 (N_6162,N_5207,N_5311);
and U6163 (N_6163,N_5432,N_5517);
and U6164 (N_6164,N_5969,N_5850);
nor U6165 (N_6165,N_5587,N_5618);
xor U6166 (N_6166,N_5119,N_5704);
and U6167 (N_6167,N_5026,N_5223);
and U6168 (N_6168,N_5663,N_5356);
nand U6169 (N_6169,N_5200,N_5332);
xor U6170 (N_6170,N_5062,N_5821);
nand U6171 (N_6171,N_5038,N_5242);
xor U6172 (N_6172,N_5097,N_5638);
xor U6173 (N_6173,N_5904,N_5431);
or U6174 (N_6174,N_5648,N_5414);
nor U6175 (N_6175,N_5688,N_5977);
nand U6176 (N_6176,N_5037,N_5137);
nand U6177 (N_6177,N_5784,N_5189);
xnor U6178 (N_6178,N_5971,N_5110);
or U6179 (N_6179,N_5372,N_5447);
nand U6180 (N_6180,N_5238,N_5334);
or U6181 (N_6181,N_5335,N_5183);
nand U6182 (N_6182,N_5787,N_5768);
nand U6183 (N_6183,N_5691,N_5032);
or U6184 (N_6184,N_5374,N_5775);
nand U6185 (N_6185,N_5770,N_5525);
xor U6186 (N_6186,N_5514,N_5323);
and U6187 (N_6187,N_5615,N_5409);
nor U6188 (N_6188,N_5586,N_5161);
xor U6189 (N_6189,N_5087,N_5342);
or U6190 (N_6190,N_5392,N_5715);
or U6191 (N_6191,N_5831,N_5162);
and U6192 (N_6192,N_5310,N_5581);
nor U6193 (N_6193,N_5178,N_5858);
xnor U6194 (N_6194,N_5806,N_5024);
nor U6195 (N_6195,N_5781,N_5990);
nor U6196 (N_6196,N_5225,N_5934);
or U6197 (N_6197,N_5692,N_5588);
xor U6198 (N_6198,N_5241,N_5566);
or U6199 (N_6199,N_5803,N_5073);
or U6200 (N_6200,N_5076,N_5885);
xnor U6201 (N_6201,N_5272,N_5740);
and U6202 (N_6202,N_5671,N_5333);
xor U6203 (N_6203,N_5003,N_5965);
and U6204 (N_6204,N_5916,N_5498);
or U6205 (N_6205,N_5751,N_5555);
xor U6206 (N_6206,N_5937,N_5529);
xor U6207 (N_6207,N_5305,N_5705);
and U6208 (N_6208,N_5453,N_5239);
or U6209 (N_6209,N_5213,N_5144);
or U6210 (N_6210,N_5880,N_5486);
nand U6211 (N_6211,N_5980,N_5221);
or U6212 (N_6212,N_5321,N_5384);
or U6213 (N_6213,N_5282,N_5470);
xnor U6214 (N_6214,N_5854,N_5693);
xor U6215 (N_6215,N_5943,N_5973);
nor U6216 (N_6216,N_5463,N_5029);
and U6217 (N_6217,N_5264,N_5005);
and U6218 (N_6218,N_5179,N_5340);
nor U6219 (N_6219,N_5840,N_5996);
xor U6220 (N_6220,N_5741,N_5442);
nand U6221 (N_6221,N_5523,N_5441);
nand U6222 (N_6222,N_5206,N_5752);
xnor U6223 (N_6223,N_5492,N_5104);
or U6224 (N_6224,N_5716,N_5468);
nand U6225 (N_6225,N_5533,N_5676);
nand U6226 (N_6226,N_5719,N_5350);
or U6227 (N_6227,N_5501,N_5896);
xor U6228 (N_6228,N_5339,N_5952);
and U6229 (N_6229,N_5728,N_5197);
nor U6230 (N_6230,N_5257,N_5619);
nor U6231 (N_6231,N_5505,N_5686);
or U6232 (N_6232,N_5027,N_5108);
or U6233 (N_6233,N_5825,N_5477);
xnor U6234 (N_6234,N_5473,N_5793);
xnor U6235 (N_6235,N_5789,N_5136);
nand U6236 (N_6236,N_5077,N_5381);
xor U6237 (N_6237,N_5809,N_5394);
nor U6238 (N_6238,N_5694,N_5778);
nor U6239 (N_6239,N_5039,N_5855);
nor U6240 (N_6240,N_5511,N_5067);
nor U6241 (N_6241,N_5923,N_5177);
nand U6242 (N_6242,N_5584,N_5628);
or U6243 (N_6243,N_5373,N_5769);
nand U6244 (N_6244,N_5304,N_5932);
nand U6245 (N_6245,N_5994,N_5126);
and U6246 (N_6246,N_5362,N_5054);
and U6247 (N_6247,N_5254,N_5231);
or U6248 (N_6248,N_5375,N_5035);
nor U6249 (N_6249,N_5742,N_5127);
xnor U6250 (N_6250,N_5496,N_5259);
xnor U6251 (N_6251,N_5330,N_5281);
nand U6252 (N_6252,N_5004,N_5961);
and U6253 (N_6253,N_5531,N_5407);
and U6254 (N_6254,N_5985,N_5856);
nand U6255 (N_6255,N_5534,N_5573);
nand U6256 (N_6256,N_5371,N_5301);
xor U6257 (N_6257,N_5873,N_5008);
xor U6258 (N_6258,N_5942,N_5763);
xor U6259 (N_6259,N_5124,N_5801);
xnor U6260 (N_6260,N_5063,N_5745);
and U6261 (N_6261,N_5724,N_5467);
xnor U6262 (N_6262,N_5152,N_5023);
nor U6263 (N_6263,N_5240,N_5118);
or U6264 (N_6264,N_5545,N_5892);
or U6265 (N_6265,N_5820,N_5382);
and U6266 (N_6266,N_5659,N_5188);
nand U6267 (N_6267,N_5539,N_5308);
nand U6268 (N_6268,N_5945,N_5700);
nor U6269 (N_6269,N_5975,N_5660);
nor U6270 (N_6270,N_5358,N_5602);
xnor U6271 (N_6271,N_5180,N_5360);
or U6272 (N_6272,N_5070,N_5597);
nor U6273 (N_6273,N_5184,N_5316);
nand U6274 (N_6274,N_5276,N_5702);
and U6275 (N_6275,N_5561,N_5256);
xnor U6276 (N_6276,N_5510,N_5749);
nor U6277 (N_6277,N_5653,N_5199);
or U6278 (N_6278,N_5757,N_5493);
nor U6279 (N_6279,N_5145,N_5734);
nand U6280 (N_6280,N_5552,N_5082);
or U6281 (N_6281,N_5580,N_5456);
xnor U6282 (N_6282,N_5379,N_5634);
or U6283 (N_6283,N_5096,N_5122);
nand U6284 (N_6284,N_5112,N_5445);
nand U6285 (N_6285,N_5170,N_5488);
and U6286 (N_6286,N_5553,N_5014);
xor U6287 (N_6287,N_5437,N_5478);
and U6288 (N_6288,N_5509,N_5930);
xor U6289 (N_6289,N_5773,N_5012);
xor U6290 (N_6290,N_5541,N_5101);
or U6291 (N_6291,N_5610,N_5018);
xor U6292 (N_6292,N_5449,N_5609);
xor U6293 (N_6293,N_5936,N_5954);
and U6294 (N_6294,N_5865,N_5664);
and U6295 (N_6295,N_5655,N_5683);
or U6296 (N_6296,N_5324,N_5211);
or U6297 (N_6297,N_5827,N_5895);
xnor U6298 (N_6298,N_5667,N_5485);
and U6299 (N_6299,N_5426,N_5251);
or U6300 (N_6300,N_5506,N_5627);
and U6301 (N_6301,N_5949,N_5125);
or U6302 (N_6302,N_5995,N_5755);
and U6303 (N_6303,N_5154,N_5237);
nor U6304 (N_6304,N_5654,N_5710);
nand U6305 (N_6305,N_5461,N_5839);
or U6306 (N_6306,N_5649,N_5866);
nand U6307 (N_6307,N_5106,N_5603);
or U6308 (N_6308,N_5296,N_5662);
or U6309 (N_6309,N_5906,N_5520);
xor U6310 (N_6310,N_5712,N_5595);
nand U6311 (N_6311,N_5234,N_5695);
and U6312 (N_6312,N_5810,N_5205);
or U6313 (N_6313,N_5326,N_5811);
and U6314 (N_6314,N_5287,N_5567);
xnor U6315 (N_6315,N_5050,N_5738);
and U6316 (N_6316,N_5933,N_5960);
xor U6317 (N_6317,N_5363,N_5889);
or U6318 (N_6318,N_5860,N_5732);
xor U6319 (N_6319,N_5701,N_5879);
nor U6320 (N_6320,N_5668,N_5103);
nor U6321 (N_6321,N_5670,N_5017);
nand U6322 (N_6322,N_5910,N_5722);
or U6323 (N_6323,N_5897,N_5380);
nor U6324 (N_6324,N_5092,N_5388);
nor U6325 (N_6325,N_5258,N_5650);
xnor U6326 (N_6326,N_5314,N_5289);
nor U6327 (N_6327,N_5736,N_5044);
nor U6328 (N_6328,N_5753,N_5348);
xnor U6329 (N_6329,N_5504,N_5614);
nor U6330 (N_6330,N_5900,N_5153);
xnor U6331 (N_6331,N_5535,N_5780);
or U6332 (N_6332,N_5673,N_5150);
nor U6333 (N_6333,N_5521,N_5926);
and U6334 (N_6334,N_5863,N_5176);
or U6335 (N_6335,N_5622,N_5066);
and U6336 (N_6336,N_5393,N_5726);
or U6337 (N_6337,N_5190,N_5215);
nand U6338 (N_6338,N_5404,N_5869);
nor U6339 (N_6339,N_5355,N_5359);
and U6340 (N_6340,N_5057,N_5053);
nor U6341 (N_6341,N_5439,N_5665);
nand U6342 (N_6342,N_5682,N_5853);
xor U6343 (N_6343,N_5547,N_5429);
or U6344 (N_6344,N_5915,N_5572);
nor U6345 (N_6345,N_5401,N_5955);
xnor U6346 (N_6346,N_5123,N_5590);
nor U6347 (N_6347,N_5061,N_5099);
or U6348 (N_6348,N_5852,N_5120);
nor U6349 (N_6349,N_5737,N_5208);
or U6350 (N_6350,N_5909,N_5950);
and U6351 (N_6351,N_5052,N_5224);
nand U6352 (N_6352,N_5630,N_5386);
nand U6353 (N_6353,N_5430,N_5294);
xnor U6354 (N_6354,N_5452,N_5469);
xnor U6355 (N_6355,N_5349,N_5158);
xnor U6356 (N_6356,N_5248,N_5146);
nand U6357 (N_6357,N_5723,N_5130);
or U6358 (N_6358,N_5571,N_5020);
and U6359 (N_6359,N_5958,N_5699);
nor U6360 (N_6360,N_5585,N_5974);
nor U6361 (N_6361,N_5230,N_5672);
and U6362 (N_6362,N_5564,N_5756);
and U6363 (N_6363,N_5167,N_5060);
nand U6364 (N_6364,N_5202,N_5708);
nand U6365 (N_6365,N_5444,N_5920);
or U6366 (N_6366,N_5181,N_5165);
nor U6367 (N_6367,N_5986,N_5093);
or U6368 (N_6368,N_5791,N_5499);
and U6369 (N_6369,N_5919,N_5844);
or U6370 (N_6370,N_5870,N_5021);
nand U6371 (N_6371,N_5048,N_5997);
and U6372 (N_6372,N_5814,N_5762);
nand U6373 (N_6373,N_5247,N_5651);
or U6374 (N_6374,N_5459,N_5443);
nand U6375 (N_6375,N_5245,N_5890);
or U6376 (N_6376,N_5487,N_5263);
xor U6377 (N_6377,N_5729,N_5819);
and U6378 (N_6378,N_5420,N_5528);
and U6379 (N_6379,N_5495,N_5864);
xor U6380 (N_6380,N_5631,N_5605);
nor U6381 (N_6381,N_5435,N_5522);
or U6382 (N_6382,N_5888,N_5941);
and U6383 (N_6383,N_5079,N_5217);
nand U6384 (N_6384,N_5471,N_5336);
nand U6385 (N_6385,N_5607,N_5807);
xor U6386 (N_6386,N_5569,N_5599);
and U6387 (N_6387,N_5957,N_5016);
nand U6388 (N_6388,N_5041,N_5894);
nor U6389 (N_6389,N_5198,N_5696);
or U6390 (N_6390,N_5143,N_5730);
or U6391 (N_6391,N_5069,N_5626);
nand U6392 (N_6392,N_5367,N_5155);
nand U6393 (N_6393,N_5883,N_5002);
and U6394 (N_6394,N_5347,N_5490);
xnor U6395 (N_6395,N_5331,N_5812);
nand U6396 (N_6396,N_5802,N_5464);
nand U6397 (N_6397,N_5652,N_5548);
nor U6398 (N_6398,N_5068,N_5842);
or U6399 (N_6399,N_5250,N_5151);
nand U6400 (N_6400,N_5542,N_5497);
nand U6401 (N_6401,N_5808,N_5921);
nand U6402 (N_6402,N_5172,N_5448);
nor U6403 (N_6403,N_5129,N_5192);
xor U6404 (N_6404,N_5421,N_5204);
nand U6405 (N_6405,N_5300,N_5640);
nand U6406 (N_6406,N_5049,N_5440);
nor U6407 (N_6407,N_5913,N_5195);
xor U6408 (N_6408,N_5657,N_5766);
nand U6409 (N_6409,N_5594,N_5091);
xnor U6410 (N_6410,N_5799,N_5679);
and U6411 (N_6411,N_5988,N_5600);
nand U6412 (N_6412,N_5881,N_5425);
nor U6413 (N_6413,N_5191,N_5882);
or U6414 (N_6414,N_5400,N_5081);
and U6415 (N_6415,N_5526,N_5233);
nand U6416 (N_6416,N_5011,N_5884);
xor U6417 (N_6417,N_5777,N_5907);
or U6418 (N_6418,N_5946,N_5674);
and U6419 (N_6419,N_5391,N_5228);
and U6420 (N_6420,N_5925,N_5824);
and U6421 (N_6421,N_5472,N_5830);
nor U6422 (N_6422,N_5466,N_5253);
or U6423 (N_6423,N_5142,N_5121);
or U6424 (N_6424,N_5621,N_5006);
nor U6425 (N_6425,N_5376,N_5368);
and U6426 (N_6426,N_5201,N_5633);
or U6427 (N_6427,N_5474,N_5822);
and U6428 (N_6428,N_5612,N_5938);
xnor U6429 (N_6429,N_5859,N_5532);
nor U6430 (N_6430,N_5168,N_5307);
and U6431 (N_6431,N_5083,N_5209);
nand U6432 (N_6432,N_5636,N_5764);
or U6433 (N_6433,N_5055,N_5987);
and U6434 (N_6434,N_5482,N_5405);
and U6435 (N_6435,N_5346,N_5871);
nand U6436 (N_6436,N_5164,N_5779);
xor U6437 (N_6437,N_5159,N_5703);
and U6438 (N_6438,N_5398,N_5519);
nand U6439 (N_6439,N_5721,N_5450);
and U6440 (N_6440,N_5252,N_5993);
and U6441 (N_6441,N_5078,N_5875);
and U6442 (N_6442,N_5518,N_5845);
nand U6443 (N_6443,N_5072,N_5576);
nor U6444 (N_6444,N_5034,N_5025);
and U6445 (N_6445,N_5454,N_5278);
xnor U6446 (N_6446,N_5681,N_5403);
xor U6447 (N_6447,N_5711,N_5033);
and U6448 (N_6448,N_5100,N_5246);
or U6449 (N_6449,N_5196,N_5601);
nand U6450 (N_6450,N_5419,N_5377);
nor U6451 (N_6451,N_5090,N_5297);
xor U6452 (N_6452,N_5064,N_5298);
xnor U6453 (N_6453,N_5302,N_5706);
nor U6454 (N_6454,N_5922,N_5748);
nor U6455 (N_6455,N_5115,N_5408);
xor U6456 (N_6456,N_5527,N_5574);
or U6457 (N_6457,N_5680,N_5833);
xor U6458 (N_6458,N_5085,N_5484);
nor U6459 (N_6459,N_5760,N_5604);
nand U6460 (N_6460,N_5059,N_5507);
nand U6461 (N_6461,N_5169,N_5560);
xnor U6462 (N_6462,N_5455,N_5105);
xnor U6463 (N_6463,N_5697,N_5731);
and U6464 (N_6464,N_5001,N_5317);
nand U6465 (N_6465,N_5508,N_5666);
or U6466 (N_6466,N_5268,N_5966);
nor U6467 (N_6467,N_5935,N_5212);
nand U6468 (N_6468,N_5999,N_5387);
nor U6469 (N_6469,N_5236,N_5028);
nand U6470 (N_6470,N_5754,N_5893);
or U6471 (N_6471,N_5593,N_5813);
nor U6472 (N_6472,N_5015,N_5785);
nand U6473 (N_6473,N_5438,N_5319);
and U6474 (N_6474,N_5043,N_5709);
or U6475 (N_6475,N_5642,N_5750);
nor U6476 (N_6476,N_5157,N_5095);
nor U6477 (N_6477,N_5219,N_5669);
nand U6478 (N_6478,N_5295,N_5274);
and U6479 (N_6479,N_5956,N_5284);
nor U6480 (N_6480,N_5598,N_5046);
or U6481 (N_6481,N_5744,N_5953);
or U6482 (N_6482,N_5874,N_5783);
nand U6483 (N_6483,N_5269,N_5328);
nand U6484 (N_6484,N_5834,N_5962);
or U6485 (N_6485,N_5045,N_5714);
or U6486 (N_6486,N_5796,N_5684);
xnor U6487 (N_6487,N_5639,N_5931);
or U6488 (N_6488,N_5417,N_5516);
nor U6489 (N_6489,N_5818,N_5306);
and U6490 (N_6490,N_5353,N_5084);
and U6491 (N_6491,N_5515,N_5991);
nand U6492 (N_6492,N_5216,N_5546);
nor U6493 (N_6493,N_5341,N_5829);
nor U6494 (N_6494,N_5273,N_5114);
nor U6495 (N_6495,N_5491,N_5579);
nand U6496 (N_6496,N_5536,N_5227);
or U6497 (N_6497,N_5271,N_5366);
or U6498 (N_6498,N_5746,N_5132);
nand U6499 (N_6499,N_5436,N_5351);
nand U6500 (N_6500,N_5026,N_5460);
nand U6501 (N_6501,N_5132,N_5062);
or U6502 (N_6502,N_5878,N_5594);
nor U6503 (N_6503,N_5127,N_5256);
and U6504 (N_6504,N_5459,N_5487);
xnor U6505 (N_6505,N_5071,N_5505);
nand U6506 (N_6506,N_5295,N_5147);
nand U6507 (N_6507,N_5802,N_5506);
nand U6508 (N_6508,N_5060,N_5455);
nand U6509 (N_6509,N_5014,N_5706);
or U6510 (N_6510,N_5904,N_5269);
and U6511 (N_6511,N_5018,N_5438);
xnor U6512 (N_6512,N_5327,N_5878);
nand U6513 (N_6513,N_5416,N_5660);
and U6514 (N_6514,N_5930,N_5412);
xor U6515 (N_6515,N_5640,N_5701);
and U6516 (N_6516,N_5486,N_5477);
and U6517 (N_6517,N_5472,N_5040);
or U6518 (N_6518,N_5271,N_5602);
and U6519 (N_6519,N_5642,N_5423);
or U6520 (N_6520,N_5149,N_5360);
nor U6521 (N_6521,N_5409,N_5522);
and U6522 (N_6522,N_5950,N_5966);
xnor U6523 (N_6523,N_5516,N_5997);
and U6524 (N_6524,N_5630,N_5584);
nor U6525 (N_6525,N_5927,N_5368);
or U6526 (N_6526,N_5435,N_5851);
nor U6527 (N_6527,N_5890,N_5519);
nor U6528 (N_6528,N_5661,N_5599);
nor U6529 (N_6529,N_5851,N_5090);
and U6530 (N_6530,N_5591,N_5780);
or U6531 (N_6531,N_5814,N_5162);
nor U6532 (N_6532,N_5831,N_5662);
xor U6533 (N_6533,N_5380,N_5519);
or U6534 (N_6534,N_5209,N_5495);
nand U6535 (N_6535,N_5970,N_5502);
and U6536 (N_6536,N_5193,N_5256);
xor U6537 (N_6537,N_5011,N_5845);
or U6538 (N_6538,N_5071,N_5613);
nand U6539 (N_6539,N_5067,N_5320);
or U6540 (N_6540,N_5839,N_5066);
nand U6541 (N_6541,N_5445,N_5858);
nand U6542 (N_6542,N_5817,N_5188);
nand U6543 (N_6543,N_5076,N_5322);
xnor U6544 (N_6544,N_5026,N_5584);
xor U6545 (N_6545,N_5639,N_5572);
or U6546 (N_6546,N_5359,N_5267);
xor U6547 (N_6547,N_5796,N_5802);
and U6548 (N_6548,N_5235,N_5884);
nor U6549 (N_6549,N_5010,N_5692);
and U6550 (N_6550,N_5888,N_5390);
nand U6551 (N_6551,N_5335,N_5936);
nor U6552 (N_6552,N_5828,N_5319);
nor U6553 (N_6553,N_5995,N_5090);
nand U6554 (N_6554,N_5752,N_5708);
or U6555 (N_6555,N_5585,N_5092);
and U6556 (N_6556,N_5530,N_5918);
nand U6557 (N_6557,N_5402,N_5917);
nor U6558 (N_6558,N_5718,N_5750);
nor U6559 (N_6559,N_5890,N_5807);
nand U6560 (N_6560,N_5216,N_5084);
nand U6561 (N_6561,N_5487,N_5773);
nand U6562 (N_6562,N_5165,N_5059);
and U6563 (N_6563,N_5258,N_5402);
or U6564 (N_6564,N_5135,N_5952);
nor U6565 (N_6565,N_5594,N_5220);
nor U6566 (N_6566,N_5302,N_5517);
nor U6567 (N_6567,N_5305,N_5092);
nor U6568 (N_6568,N_5797,N_5128);
nand U6569 (N_6569,N_5215,N_5266);
xnor U6570 (N_6570,N_5410,N_5444);
or U6571 (N_6571,N_5052,N_5423);
nand U6572 (N_6572,N_5021,N_5249);
nand U6573 (N_6573,N_5770,N_5091);
and U6574 (N_6574,N_5561,N_5012);
xnor U6575 (N_6575,N_5538,N_5418);
nand U6576 (N_6576,N_5576,N_5520);
nor U6577 (N_6577,N_5933,N_5067);
or U6578 (N_6578,N_5312,N_5990);
xor U6579 (N_6579,N_5631,N_5659);
and U6580 (N_6580,N_5723,N_5056);
or U6581 (N_6581,N_5041,N_5794);
or U6582 (N_6582,N_5323,N_5502);
nand U6583 (N_6583,N_5935,N_5622);
or U6584 (N_6584,N_5484,N_5340);
nor U6585 (N_6585,N_5381,N_5736);
or U6586 (N_6586,N_5598,N_5573);
nand U6587 (N_6587,N_5247,N_5600);
and U6588 (N_6588,N_5192,N_5286);
and U6589 (N_6589,N_5736,N_5255);
nor U6590 (N_6590,N_5239,N_5655);
and U6591 (N_6591,N_5424,N_5502);
xnor U6592 (N_6592,N_5554,N_5119);
xnor U6593 (N_6593,N_5215,N_5685);
nor U6594 (N_6594,N_5290,N_5648);
or U6595 (N_6595,N_5158,N_5532);
nor U6596 (N_6596,N_5490,N_5476);
nand U6597 (N_6597,N_5713,N_5757);
or U6598 (N_6598,N_5469,N_5361);
xnor U6599 (N_6599,N_5094,N_5643);
nor U6600 (N_6600,N_5338,N_5841);
xnor U6601 (N_6601,N_5209,N_5823);
and U6602 (N_6602,N_5748,N_5849);
and U6603 (N_6603,N_5628,N_5185);
nand U6604 (N_6604,N_5397,N_5100);
nand U6605 (N_6605,N_5945,N_5892);
nor U6606 (N_6606,N_5533,N_5601);
or U6607 (N_6607,N_5310,N_5602);
or U6608 (N_6608,N_5344,N_5695);
xor U6609 (N_6609,N_5098,N_5536);
nand U6610 (N_6610,N_5927,N_5868);
and U6611 (N_6611,N_5698,N_5831);
and U6612 (N_6612,N_5210,N_5766);
nand U6613 (N_6613,N_5871,N_5893);
xnor U6614 (N_6614,N_5818,N_5694);
xor U6615 (N_6615,N_5837,N_5811);
xor U6616 (N_6616,N_5030,N_5445);
and U6617 (N_6617,N_5601,N_5929);
nor U6618 (N_6618,N_5169,N_5316);
xor U6619 (N_6619,N_5393,N_5285);
and U6620 (N_6620,N_5556,N_5461);
and U6621 (N_6621,N_5555,N_5408);
nor U6622 (N_6622,N_5782,N_5023);
and U6623 (N_6623,N_5103,N_5123);
or U6624 (N_6624,N_5472,N_5967);
or U6625 (N_6625,N_5561,N_5577);
nor U6626 (N_6626,N_5902,N_5850);
xor U6627 (N_6627,N_5136,N_5545);
nand U6628 (N_6628,N_5797,N_5848);
or U6629 (N_6629,N_5545,N_5967);
and U6630 (N_6630,N_5099,N_5780);
or U6631 (N_6631,N_5843,N_5007);
nor U6632 (N_6632,N_5608,N_5812);
xnor U6633 (N_6633,N_5600,N_5349);
xor U6634 (N_6634,N_5768,N_5452);
or U6635 (N_6635,N_5638,N_5210);
nor U6636 (N_6636,N_5111,N_5929);
and U6637 (N_6637,N_5751,N_5008);
nand U6638 (N_6638,N_5527,N_5044);
nand U6639 (N_6639,N_5655,N_5083);
xnor U6640 (N_6640,N_5386,N_5754);
nand U6641 (N_6641,N_5082,N_5727);
or U6642 (N_6642,N_5074,N_5635);
nand U6643 (N_6643,N_5705,N_5577);
xor U6644 (N_6644,N_5572,N_5015);
nor U6645 (N_6645,N_5025,N_5541);
or U6646 (N_6646,N_5499,N_5226);
nor U6647 (N_6647,N_5396,N_5529);
or U6648 (N_6648,N_5419,N_5710);
nand U6649 (N_6649,N_5243,N_5798);
nand U6650 (N_6650,N_5875,N_5657);
nor U6651 (N_6651,N_5824,N_5901);
xor U6652 (N_6652,N_5112,N_5111);
nor U6653 (N_6653,N_5153,N_5384);
and U6654 (N_6654,N_5107,N_5309);
nand U6655 (N_6655,N_5687,N_5152);
and U6656 (N_6656,N_5894,N_5630);
and U6657 (N_6657,N_5912,N_5252);
nand U6658 (N_6658,N_5004,N_5626);
xnor U6659 (N_6659,N_5354,N_5656);
nand U6660 (N_6660,N_5211,N_5201);
or U6661 (N_6661,N_5371,N_5411);
xor U6662 (N_6662,N_5101,N_5118);
nand U6663 (N_6663,N_5065,N_5745);
and U6664 (N_6664,N_5561,N_5098);
xor U6665 (N_6665,N_5991,N_5498);
nand U6666 (N_6666,N_5938,N_5941);
nand U6667 (N_6667,N_5530,N_5614);
nand U6668 (N_6668,N_5702,N_5077);
xor U6669 (N_6669,N_5868,N_5061);
nor U6670 (N_6670,N_5634,N_5505);
and U6671 (N_6671,N_5978,N_5857);
or U6672 (N_6672,N_5547,N_5503);
nor U6673 (N_6673,N_5289,N_5883);
nand U6674 (N_6674,N_5561,N_5866);
nor U6675 (N_6675,N_5587,N_5839);
and U6676 (N_6676,N_5935,N_5220);
xor U6677 (N_6677,N_5028,N_5582);
nand U6678 (N_6678,N_5704,N_5164);
and U6679 (N_6679,N_5366,N_5463);
nor U6680 (N_6680,N_5029,N_5266);
xnor U6681 (N_6681,N_5168,N_5863);
and U6682 (N_6682,N_5695,N_5798);
nor U6683 (N_6683,N_5660,N_5519);
or U6684 (N_6684,N_5201,N_5824);
nor U6685 (N_6685,N_5295,N_5413);
xnor U6686 (N_6686,N_5863,N_5463);
nor U6687 (N_6687,N_5908,N_5276);
xnor U6688 (N_6688,N_5284,N_5010);
nand U6689 (N_6689,N_5807,N_5864);
or U6690 (N_6690,N_5621,N_5795);
or U6691 (N_6691,N_5148,N_5710);
nor U6692 (N_6692,N_5070,N_5676);
nor U6693 (N_6693,N_5878,N_5887);
or U6694 (N_6694,N_5506,N_5568);
nor U6695 (N_6695,N_5901,N_5650);
or U6696 (N_6696,N_5694,N_5985);
nor U6697 (N_6697,N_5564,N_5562);
xnor U6698 (N_6698,N_5004,N_5766);
and U6699 (N_6699,N_5659,N_5806);
nor U6700 (N_6700,N_5531,N_5184);
nand U6701 (N_6701,N_5910,N_5977);
or U6702 (N_6702,N_5065,N_5837);
xnor U6703 (N_6703,N_5148,N_5162);
nor U6704 (N_6704,N_5458,N_5420);
or U6705 (N_6705,N_5315,N_5097);
nor U6706 (N_6706,N_5197,N_5368);
and U6707 (N_6707,N_5004,N_5213);
or U6708 (N_6708,N_5091,N_5694);
xor U6709 (N_6709,N_5044,N_5555);
nand U6710 (N_6710,N_5044,N_5731);
nor U6711 (N_6711,N_5265,N_5505);
or U6712 (N_6712,N_5121,N_5702);
or U6713 (N_6713,N_5675,N_5523);
xnor U6714 (N_6714,N_5466,N_5270);
and U6715 (N_6715,N_5750,N_5708);
or U6716 (N_6716,N_5017,N_5617);
or U6717 (N_6717,N_5248,N_5630);
xor U6718 (N_6718,N_5248,N_5160);
or U6719 (N_6719,N_5702,N_5617);
or U6720 (N_6720,N_5353,N_5664);
or U6721 (N_6721,N_5463,N_5361);
or U6722 (N_6722,N_5584,N_5565);
nor U6723 (N_6723,N_5559,N_5806);
and U6724 (N_6724,N_5516,N_5684);
and U6725 (N_6725,N_5669,N_5721);
xor U6726 (N_6726,N_5002,N_5621);
xor U6727 (N_6727,N_5769,N_5623);
or U6728 (N_6728,N_5020,N_5878);
nand U6729 (N_6729,N_5658,N_5163);
xnor U6730 (N_6730,N_5452,N_5247);
xnor U6731 (N_6731,N_5868,N_5272);
or U6732 (N_6732,N_5280,N_5059);
or U6733 (N_6733,N_5045,N_5048);
or U6734 (N_6734,N_5260,N_5692);
xnor U6735 (N_6735,N_5587,N_5573);
or U6736 (N_6736,N_5311,N_5644);
and U6737 (N_6737,N_5060,N_5597);
and U6738 (N_6738,N_5402,N_5405);
nand U6739 (N_6739,N_5463,N_5277);
nor U6740 (N_6740,N_5722,N_5459);
xor U6741 (N_6741,N_5813,N_5242);
xor U6742 (N_6742,N_5223,N_5454);
xnor U6743 (N_6743,N_5715,N_5279);
or U6744 (N_6744,N_5211,N_5113);
nand U6745 (N_6745,N_5986,N_5013);
nand U6746 (N_6746,N_5477,N_5523);
or U6747 (N_6747,N_5995,N_5657);
nor U6748 (N_6748,N_5930,N_5042);
and U6749 (N_6749,N_5578,N_5726);
and U6750 (N_6750,N_5741,N_5097);
or U6751 (N_6751,N_5658,N_5025);
nand U6752 (N_6752,N_5124,N_5614);
or U6753 (N_6753,N_5021,N_5996);
nor U6754 (N_6754,N_5532,N_5291);
and U6755 (N_6755,N_5683,N_5390);
nor U6756 (N_6756,N_5741,N_5016);
nand U6757 (N_6757,N_5122,N_5313);
nand U6758 (N_6758,N_5748,N_5098);
nand U6759 (N_6759,N_5364,N_5158);
and U6760 (N_6760,N_5458,N_5073);
xor U6761 (N_6761,N_5182,N_5470);
and U6762 (N_6762,N_5627,N_5523);
or U6763 (N_6763,N_5095,N_5519);
nor U6764 (N_6764,N_5324,N_5990);
and U6765 (N_6765,N_5498,N_5147);
xnor U6766 (N_6766,N_5392,N_5805);
and U6767 (N_6767,N_5174,N_5726);
and U6768 (N_6768,N_5173,N_5718);
xor U6769 (N_6769,N_5138,N_5265);
xor U6770 (N_6770,N_5320,N_5117);
and U6771 (N_6771,N_5615,N_5547);
nand U6772 (N_6772,N_5212,N_5444);
xnor U6773 (N_6773,N_5297,N_5177);
xnor U6774 (N_6774,N_5448,N_5585);
nor U6775 (N_6775,N_5980,N_5941);
nor U6776 (N_6776,N_5612,N_5743);
nand U6777 (N_6777,N_5601,N_5288);
and U6778 (N_6778,N_5350,N_5068);
nand U6779 (N_6779,N_5679,N_5409);
nor U6780 (N_6780,N_5447,N_5803);
nor U6781 (N_6781,N_5458,N_5931);
nor U6782 (N_6782,N_5435,N_5905);
nand U6783 (N_6783,N_5894,N_5109);
and U6784 (N_6784,N_5110,N_5323);
or U6785 (N_6785,N_5644,N_5972);
xor U6786 (N_6786,N_5712,N_5491);
nor U6787 (N_6787,N_5373,N_5980);
nand U6788 (N_6788,N_5096,N_5008);
or U6789 (N_6789,N_5788,N_5221);
nand U6790 (N_6790,N_5718,N_5388);
or U6791 (N_6791,N_5964,N_5046);
nor U6792 (N_6792,N_5691,N_5308);
xor U6793 (N_6793,N_5841,N_5342);
or U6794 (N_6794,N_5236,N_5135);
nand U6795 (N_6795,N_5271,N_5203);
nand U6796 (N_6796,N_5459,N_5688);
and U6797 (N_6797,N_5733,N_5085);
nor U6798 (N_6798,N_5434,N_5715);
or U6799 (N_6799,N_5581,N_5928);
xnor U6800 (N_6800,N_5372,N_5109);
xor U6801 (N_6801,N_5055,N_5999);
xor U6802 (N_6802,N_5347,N_5101);
and U6803 (N_6803,N_5544,N_5774);
and U6804 (N_6804,N_5447,N_5080);
xnor U6805 (N_6805,N_5643,N_5427);
xor U6806 (N_6806,N_5182,N_5312);
nand U6807 (N_6807,N_5158,N_5429);
or U6808 (N_6808,N_5567,N_5827);
or U6809 (N_6809,N_5578,N_5931);
nand U6810 (N_6810,N_5717,N_5294);
and U6811 (N_6811,N_5257,N_5521);
nor U6812 (N_6812,N_5599,N_5488);
nor U6813 (N_6813,N_5461,N_5147);
nand U6814 (N_6814,N_5652,N_5476);
xor U6815 (N_6815,N_5150,N_5514);
nand U6816 (N_6816,N_5182,N_5564);
xor U6817 (N_6817,N_5226,N_5346);
and U6818 (N_6818,N_5097,N_5839);
nand U6819 (N_6819,N_5810,N_5037);
or U6820 (N_6820,N_5385,N_5390);
or U6821 (N_6821,N_5226,N_5021);
and U6822 (N_6822,N_5081,N_5782);
nand U6823 (N_6823,N_5917,N_5184);
nor U6824 (N_6824,N_5891,N_5596);
and U6825 (N_6825,N_5031,N_5491);
nand U6826 (N_6826,N_5640,N_5318);
and U6827 (N_6827,N_5056,N_5985);
or U6828 (N_6828,N_5476,N_5377);
or U6829 (N_6829,N_5466,N_5823);
nor U6830 (N_6830,N_5718,N_5517);
nand U6831 (N_6831,N_5036,N_5118);
nand U6832 (N_6832,N_5733,N_5954);
nand U6833 (N_6833,N_5644,N_5717);
or U6834 (N_6834,N_5029,N_5630);
nor U6835 (N_6835,N_5973,N_5039);
xnor U6836 (N_6836,N_5748,N_5674);
nand U6837 (N_6837,N_5819,N_5744);
nor U6838 (N_6838,N_5028,N_5248);
xnor U6839 (N_6839,N_5981,N_5905);
nand U6840 (N_6840,N_5662,N_5652);
and U6841 (N_6841,N_5583,N_5859);
or U6842 (N_6842,N_5875,N_5679);
and U6843 (N_6843,N_5821,N_5858);
and U6844 (N_6844,N_5185,N_5682);
nor U6845 (N_6845,N_5211,N_5517);
nand U6846 (N_6846,N_5604,N_5399);
xor U6847 (N_6847,N_5078,N_5997);
nand U6848 (N_6848,N_5629,N_5443);
xnor U6849 (N_6849,N_5458,N_5567);
xor U6850 (N_6850,N_5243,N_5947);
xor U6851 (N_6851,N_5094,N_5265);
nand U6852 (N_6852,N_5496,N_5080);
xor U6853 (N_6853,N_5870,N_5492);
nor U6854 (N_6854,N_5214,N_5674);
or U6855 (N_6855,N_5646,N_5645);
xor U6856 (N_6856,N_5937,N_5707);
nand U6857 (N_6857,N_5483,N_5634);
and U6858 (N_6858,N_5251,N_5125);
nor U6859 (N_6859,N_5478,N_5398);
nor U6860 (N_6860,N_5734,N_5113);
nor U6861 (N_6861,N_5981,N_5338);
and U6862 (N_6862,N_5794,N_5693);
xnor U6863 (N_6863,N_5615,N_5725);
or U6864 (N_6864,N_5854,N_5453);
nand U6865 (N_6865,N_5526,N_5654);
nand U6866 (N_6866,N_5050,N_5538);
nor U6867 (N_6867,N_5247,N_5599);
nand U6868 (N_6868,N_5033,N_5163);
nand U6869 (N_6869,N_5856,N_5122);
and U6870 (N_6870,N_5714,N_5838);
nand U6871 (N_6871,N_5451,N_5412);
and U6872 (N_6872,N_5287,N_5839);
nor U6873 (N_6873,N_5249,N_5927);
nor U6874 (N_6874,N_5432,N_5053);
nor U6875 (N_6875,N_5187,N_5890);
nor U6876 (N_6876,N_5068,N_5642);
and U6877 (N_6877,N_5674,N_5960);
xnor U6878 (N_6878,N_5710,N_5400);
and U6879 (N_6879,N_5591,N_5585);
and U6880 (N_6880,N_5437,N_5758);
nand U6881 (N_6881,N_5010,N_5676);
or U6882 (N_6882,N_5852,N_5819);
xnor U6883 (N_6883,N_5502,N_5450);
xor U6884 (N_6884,N_5724,N_5781);
or U6885 (N_6885,N_5031,N_5941);
or U6886 (N_6886,N_5481,N_5717);
nand U6887 (N_6887,N_5496,N_5003);
xnor U6888 (N_6888,N_5009,N_5164);
or U6889 (N_6889,N_5185,N_5243);
and U6890 (N_6890,N_5740,N_5235);
or U6891 (N_6891,N_5124,N_5380);
nand U6892 (N_6892,N_5447,N_5232);
and U6893 (N_6893,N_5782,N_5899);
or U6894 (N_6894,N_5874,N_5113);
nor U6895 (N_6895,N_5204,N_5360);
nand U6896 (N_6896,N_5097,N_5291);
nand U6897 (N_6897,N_5429,N_5882);
nor U6898 (N_6898,N_5670,N_5393);
xnor U6899 (N_6899,N_5068,N_5531);
nand U6900 (N_6900,N_5536,N_5217);
nor U6901 (N_6901,N_5891,N_5104);
or U6902 (N_6902,N_5791,N_5196);
nor U6903 (N_6903,N_5648,N_5745);
nand U6904 (N_6904,N_5652,N_5970);
nand U6905 (N_6905,N_5618,N_5916);
and U6906 (N_6906,N_5298,N_5987);
nand U6907 (N_6907,N_5857,N_5619);
nand U6908 (N_6908,N_5241,N_5476);
nor U6909 (N_6909,N_5469,N_5335);
or U6910 (N_6910,N_5005,N_5366);
nand U6911 (N_6911,N_5877,N_5672);
and U6912 (N_6912,N_5068,N_5100);
nor U6913 (N_6913,N_5353,N_5335);
and U6914 (N_6914,N_5025,N_5750);
nand U6915 (N_6915,N_5636,N_5248);
or U6916 (N_6916,N_5970,N_5314);
xnor U6917 (N_6917,N_5423,N_5908);
or U6918 (N_6918,N_5671,N_5101);
and U6919 (N_6919,N_5141,N_5859);
nor U6920 (N_6920,N_5398,N_5788);
or U6921 (N_6921,N_5472,N_5802);
or U6922 (N_6922,N_5380,N_5532);
or U6923 (N_6923,N_5803,N_5003);
and U6924 (N_6924,N_5571,N_5010);
xnor U6925 (N_6925,N_5508,N_5989);
nand U6926 (N_6926,N_5674,N_5553);
or U6927 (N_6927,N_5896,N_5676);
xnor U6928 (N_6928,N_5091,N_5405);
nor U6929 (N_6929,N_5830,N_5902);
nor U6930 (N_6930,N_5805,N_5518);
xor U6931 (N_6931,N_5742,N_5855);
nand U6932 (N_6932,N_5381,N_5342);
and U6933 (N_6933,N_5984,N_5582);
nor U6934 (N_6934,N_5103,N_5460);
nand U6935 (N_6935,N_5081,N_5427);
nand U6936 (N_6936,N_5018,N_5913);
nor U6937 (N_6937,N_5207,N_5043);
or U6938 (N_6938,N_5256,N_5515);
nand U6939 (N_6939,N_5431,N_5271);
nand U6940 (N_6940,N_5611,N_5100);
nand U6941 (N_6941,N_5031,N_5572);
nand U6942 (N_6942,N_5298,N_5789);
nor U6943 (N_6943,N_5657,N_5580);
or U6944 (N_6944,N_5591,N_5647);
nand U6945 (N_6945,N_5547,N_5356);
and U6946 (N_6946,N_5407,N_5765);
or U6947 (N_6947,N_5899,N_5119);
or U6948 (N_6948,N_5042,N_5889);
or U6949 (N_6949,N_5564,N_5602);
or U6950 (N_6950,N_5202,N_5768);
nand U6951 (N_6951,N_5935,N_5301);
xnor U6952 (N_6952,N_5011,N_5521);
xor U6953 (N_6953,N_5859,N_5137);
and U6954 (N_6954,N_5421,N_5771);
or U6955 (N_6955,N_5127,N_5416);
and U6956 (N_6956,N_5217,N_5011);
or U6957 (N_6957,N_5630,N_5825);
xnor U6958 (N_6958,N_5411,N_5079);
nand U6959 (N_6959,N_5166,N_5351);
and U6960 (N_6960,N_5434,N_5063);
and U6961 (N_6961,N_5545,N_5093);
xor U6962 (N_6962,N_5939,N_5104);
or U6963 (N_6963,N_5179,N_5669);
and U6964 (N_6964,N_5227,N_5458);
or U6965 (N_6965,N_5890,N_5147);
nor U6966 (N_6966,N_5407,N_5744);
or U6967 (N_6967,N_5134,N_5997);
xnor U6968 (N_6968,N_5013,N_5533);
and U6969 (N_6969,N_5819,N_5512);
xor U6970 (N_6970,N_5451,N_5488);
xor U6971 (N_6971,N_5684,N_5279);
or U6972 (N_6972,N_5401,N_5885);
nand U6973 (N_6973,N_5211,N_5288);
or U6974 (N_6974,N_5654,N_5881);
or U6975 (N_6975,N_5316,N_5910);
nand U6976 (N_6976,N_5702,N_5055);
or U6977 (N_6977,N_5088,N_5370);
and U6978 (N_6978,N_5015,N_5723);
nor U6979 (N_6979,N_5854,N_5469);
or U6980 (N_6980,N_5957,N_5303);
or U6981 (N_6981,N_5788,N_5635);
and U6982 (N_6982,N_5449,N_5765);
nand U6983 (N_6983,N_5265,N_5657);
nor U6984 (N_6984,N_5746,N_5249);
xnor U6985 (N_6985,N_5410,N_5495);
nand U6986 (N_6986,N_5784,N_5197);
nand U6987 (N_6987,N_5823,N_5192);
and U6988 (N_6988,N_5120,N_5660);
nand U6989 (N_6989,N_5349,N_5552);
nor U6990 (N_6990,N_5847,N_5427);
or U6991 (N_6991,N_5544,N_5489);
and U6992 (N_6992,N_5767,N_5987);
nor U6993 (N_6993,N_5981,N_5014);
or U6994 (N_6994,N_5561,N_5611);
or U6995 (N_6995,N_5919,N_5888);
or U6996 (N_6996,N_5701,N_5403);
and U6997 (N_6997,N_5204,N_5523);
and U6998 (N_6998,N_5923,N_5468);
or U6999 (N_6999,N_5839,N_5286);
xnor U7000 (N_7000,N_6621,N_6868);
xor U7001 (N_7001,N_6610,N_6581);
nor U7002 (N_7002,N_6889,N_6335);
and U7003 (N_7003,N_6405,N_6729);
nor U7004 (N_7004,N_6428,N_6858);
xnor U7005 (N_7005,N_6835,N_6568);
xnor U7006 (N_7006,N_6271,N_6305);
nand U7007 (N_7007,N_6480,N_6855);
nand U7008 (N_7008,N_6218,N_6642);
nor U7009 (N_7009,N_6607,N_6413);
nand U7010 (N_7010,N_6631,N_6167);
nand U7011 (N_7011,N_6865,N_6069);
nand U7012 (N_7012,N_6301,N_6102);
nand U7013 (N_7013,N_6742,N_6478);
xor U7014 (N_7014,N_6692,N_6286);
xor U7015 (N_7015,N_6974,N_6097);
and U7016 (N_7016,N_6222,N_6947);
or U7017 (N_7017,N_6163,N_6110);
and U7018 (N_7018,N_6664,N_6346);
xor U7019 (N_7019,N_6202,N_6979);
nand U7020 (N_7020,N_6613,N_6698);
nor U7021 (N_7021,N_6980,N_6015);
and U7022 (N_7022,N_6871,N_6825);
xnor U7023 (N_7023,N_6806,N_6074);
xnor U7024 (N_7024,N_6040,N_6997);
and U7025 (N_7025,N_6052,N_6216);
xor U7026 (N_7026,N_6454,N_6598);
nand U7027 (N_7027,N_6616,N_6435);
xor U7028 (N_7028,N_6433,N_6994);
xnor U7029 (N_7029,N_6025,N_6922);
xor U7030 (N_7030,N_6063,N_6768);
or U7031 (N_7031,N_6227,N_6936);
and U7032 (N_7032,N_6911,N_6123);
or U7033 (N_7033,N_6733,N_6961);
and U7034 (N_7034,N_6907,N_6763);
and U7035 (N_7035,N_6141,N_6067);
nand U7036 (N_7036,N_6073,N_6691);
nor U7037 (N_7037,N_6426,N_6926);
xnor U7038 (N_7038,N_6430,N_6471);
xnor U7039 (N_7039,N_6467,N_6668);
and U7040 (N_7040,N_6627,N_6963);
nand U7041 (N_7041,N_6185,N_6432);
and U7042 (N_7042,N_6001,N_6279);
and U7043 (N_7043,N_6083,N_6045);
or U7044 (N_7044,N_6233,N_6542);
or U7045 (N_7045,N_6833,N_6557);
nand U7046 (N_7046,N_6887,N_6162);
and U7047 (N_7047,N_6132,N_6814);
nor U7048 (N_7048,N_6283,N_6658);
nand U7049 (N_7049,N_6470,N_6273);
nor U7050 (N_7050,N_6869,N_6601);
nand U7051 (N_7051,N_6131,N_6453);
nand U7052 (N_7052,N_6307,N_6217);
nor U7053 (N_7053,N_6295,N_6574);
nor U7054 (N_7054,N_6489,N_6314);
and U7055 (N_7055,N_6700,N_6731);
and U7056 (N_7056,N_6367,N_6565);
nor U7057 (N_7057,N_6164,N_6970);
xor U7058 (N_7058,N_6502,N_6127);
or U7059 (N_7059,N_6667,N_6014);
xor U7060 (N_7060,N_6894,N_6673);
nor U7061 (N_7061,N_6312,N_6382);
and U7062 (N_7062,N_6925,N_6477);
nor U7063 (N_7063,N_6678,N_6751);
or U7064 (N_7064,N_6065,N_6674);
and U7065 (N_7065,N_6860,N_6340);
and U7066 (N_7066,N_6921,N_6807);
nor U7067 (N_7067,N_6361,N_6856);
nor U7068 (N_7068,N_6559,N_6089);
and U7069 (N_7069,N_6838,N_6836);
or U7070 (N_7070,N_6122,N_6830);
or U7071 (N_7071,N_6289,N_6592);
and U7072 (N_7072,N_6403,N_6615);
and U7073 (N_7073,N_6583,N_6517);
nand U7074 (N_7074,N_6696,N_6969);
or U7075 (N_7075,N_6495,N_6804);
xnor U7076 (N_7076,N_6556,N_6735);
xnor U7077 (N_7077,N_6369,N_6626);
or U7078 (N_7078,N_6038,N_6705);
nor U7079 (N_7079,N_6421,N_6659);
nor U7080 (N_7080,N_6447,N_6680);
nand U7081 (N_7081,N_6212,N_6445);
and U7082 (N_7082,N_6460,N_6910);
xnor U7083 (N_7083,N_6928,N_6986);
xor U7084 (N_7084,N_6945,N_6012);
xnor U7085 (N_7085,N_6180,N_6396);
nor U7086 (N_7086,N_6114,N_6165);
xnor U7087 (N_7087,N_6573,N_6579);
or U7088 (N_7088,N_6042,N_6812);
xor U7089 (N_7089,N_6635,N_6550);
nor U7090 (N_7090,N_6702,N_6071);
xnor U7091 (N_7091,N_6389,N_6727);
and U7092 (N_7092,N_6618,N_6243);
nor U7093 (N_7093,N_6786,N_6844);
and U7094 (N_7094,N_6656,N_6646);
or U7095 (N_7095,N_6126,N_6750);
or U7096 (N_7096,N_6490,N_6730);
and U7097 (N_7097,N_6684,N_6745);
and U7098 (N_7098,N_6602,N_6992);
and U7099 (N_7099,N_6140,N_6157);
xnor U7100 (N_7100,N_6739,N_6561);
and U7101 (N_7101,N_6420,N_6117);
nor U7102 (N_7102,N_6917,N_6004);
or U7103 (N_7103,N_6996,N_6541);
and U7104 (N_7104,N_6189,N_6406);
nor U7105 (N_7105,N_6670,N_6688);
or U7106 (N_7106,N_6983,N_6087);
and U7107 (N_7107,N_6138,N_6210);
nand U7108 (N_7108,N_6535,N_6054);
nand U7109 (N_7109,N_6392,N_6240);
and U7110 (N_7110,N_6169,N_6133);
or U7111 (N_7111,N_6538,N_6712);
xnor U7112 (N_7112,N_6451,N_6563);
nand U7113 (N_7113,N_6029,N_6000);
nor U7114 (N_7114,N_6671,N_6266);
or U7115 (N_7115,N_6352,N_6913);
xnor U7116 (N_7116,N_6802,N_6046);
nor U7117 (N_7117,N_6755,N_6648);
and U7118 (N_7118,N_6724,N_6205);
nor U7119 (N_7119,N_6519,N_6024);
nor U7120 (N_7120,N_6697,N_6575);
and U7121 (N_7121,N_6251,N_6619);
xnor U7122 (N_7122,N_6297,N_6510);
nor U7123 (N_7123,N_6170,N_6603);
or U7124 (N_7124,N_6766,N_6899);
nor U7125 (N_7125,N_6515,N_6640);
nand U7126 (N_7126,N_6867,N_6360);
xor U7127 (N_7127,N_6417,N_6546);
or U7128 (N_7128,N_6896,N_6407);
xnor U7129 (N_7129,N_6683,N_6919);
xnor U7130 (N_7130,N_6752,N_6155);
and U7131 (N_7131,N_6672,N_6070);
or U7132 (N_7132,N_6274,N_6225);
or U7133 (N_7133,N_6464,N_6773);
nor U7134 (N_7134,N_6657,N_6077);
or U7135 (N_7135,N_6456,N_6508);
and U7136 (N_7136,N_6675,N_6325);
nor U7137 (N_7137,N_6713,N_6536);
xor U7138 (N_7138,N_6452,N_6881);
nor U7139 (N_7139,N_6181,N_6522);
nand U7140 (N_7140,N_6507,N_6422);
nor U7141 (N_7141,N_6061,N_6245);
or U7142 (N_7142,N_6566,N_6577);
or U7143 (N_7143,N_6606,N_6687);
or U7144 (N_7144,N_6008,N_6526);
or U7145 (N_7145,N_6689,N_6144);
nor U7146 (N_7146,N_6135,N_6770);
and U7147 (N_7147,N_6484,N_6736);
and U7148 (N_7148,N_6803,N_6857);
or U7149 (N_7149,N_6436,N_6638);
or U7150 (N_7150,N_6021,N_6861);
nand U7151 (N_7151,N_6831,N_6439);
nor U7152 (N_7152,N_6438,N_6588);
xnor U7153 (N_7153,N_6322,N_6387);
or U7154 (N_7154,N_6296,N_6118);
and U7155 (N_7155,N_6381,N_6234);
and U7156 (N_7156,N_6115,N_6554);
nand U7157 (N_7157,N_6570,N_6954);
or U7158 (N_7158,N_6276,N_6278);
nand U7159 (N_7159,N_6875,N_6419);
and U7160 (N_7160,N_6776,N_6832);
nand U7161 (N_7161,N_6820,N_6036);
nand U7162 (N_7162,N_6548,N_6564);
xnor U7163 (N_7163,N_6028,N_6319);
xnor U7164 (N_7164,N_6043,N_6524);
nand U7165 (N_7165,N_6842,N_6347);
nand U7166 (N_7166,N_6125,N_6909);
or U7167 (N_7167,N_6794,N_6874);
nand U7168 (N_7168,N_6280,N_6553);
nor U7169 (N_7169,N_6142,N_6800);
xnor U7170 (N_7170,N_6264,N_6967);
nand U7171 (N_7171,N_6330,N_6878);
and U7172 (N_7172,N_6385,N_6375);
and U7173 (N_7173,N_6408,N_6946);
xor U7174 (N_7174,N_6487,N_6754);
xnor U7175 (N_7175,N_6081,N_6402);
and U7176 (N_7176,N_6549,N_6977);
or U7177 (N_7177,N_6275,N_6300);
xor U7178 (N_7178,N_6509,N_6262);
nand U7179 (N_7179,N_6174,N_6989);
or U7180 (N_7180,N_6485,N_6044);
or U7181 (N_7181,N_6840,N_6308);
and U7182 (N_7182,N_6746,N_6728);
nand U7183 (N_7183,N_6363,N_6242);
or U7184 (N_7184,N_6187,N_6531);
xnor U7185 (N_7185,N_6228,N_6810);
nor U7186 (N_7186,N_6639,N_6533);
and U7187 (N_7187,N_6379,N_6993);
or U7188 (N_7188,N_6176,N_6192);
nor U7189 (N_7189,N_6323,N_6320);
xor U7190 (N_7190,N_6152,N_6383);
nor U7191 (N_7191,N_6186,N_6207);
xor U7192 (N_7192,N_6666,N_6331);
nand U7193 (N_7193,N_6523,N_6771);
nand U7194 (N_7194,N_6950,N_6880);
or U7195 (N_7195,N_6194,N_6787);
nor U7196 (N_7196,N_6269,N_6545);
or U7197 (N_7197,N_6514,N_6235);
xor U7198 (N_7198,N_6748,N_6605);
and U7199 (N_7199,N_6551,N_6534);
nand U7200 (N_7200,N_6364,N_6304);
xor U7201 (N_7201,N_6372,N_6769);
xnor U7202 (N_7202,N_6350,N_6654);
and U7203 (N_7203,N_6898,N_6962);
nor U7204 (N_7204,N_6356,N_6968);
xnor U7205 (N_7205,N_6411,N_6665);
nor U7206 (N_7206,N_6506,N_6050);
xor U7207 (N_7207,N_6359,N_6255);
nor U7208 (N_7208,N_6048,N_6410);
nor U7209 (N_7209,N_6734,N_6529);
or U7210 (N_7210,N_6294,N_6645);
nor U7211 (N_7211,N_6394,N_6175);
xor U7212 (N_7212,N_6013,N_6003);
nor U7213 (N_7213,N_6516,N_6572);
and U7214 (N_7214,N_6608,N_6846);
or U7215 (N_7215,N_6479,N_6850);
nand U7216 (N_7216,N_6595,N_6412);
nor U7217 (N_7217,N_6512,N_6075);
nand U7218 (N_7218,N_6253,N_6571);
nor U7219 (N_7219,N_6504,N_6448);
nor U7220 (N_7220,N_6808,N_6941);
nand U7221 (N_7221,N_6384,N_6064);
nand U7222 (N_7222,N_6877,N_6111);
nand U7223 (N_7223,N_6079,N_6791);
and U7224 (N_7224,N_6332,N_6316);
or U7225 (N_7225,N_6298,N_6034);
nor U7226 (N_7226,N_6268,N_6190);
nand U7227 (N_7227,N_6873,N_6890);
nand U7228 (N_7228,N_6895,N_6530);
nor U7229 (N_7229,N_6146,N_6722);
and U7230 (N_7230,N_6468,N_6982);
or U7231 (N_7231,N_6465,N_6520);
and U7232 (N_7232,N_6972,N_6472);
nand U7233 (N_7233,N_6906,N_6441);
or U7234 (N_7234,N_6965,N_6695);
xor U7235 (N_7235,N_6784,N_6197);
or U7236 (N_7236,N_6949,N_6912);
xnor U7237 (N_7237,N_6237,N_6976);
or U7238 (N_7238,N_6981,N_6049);
nand U7239 (N_7239,N_6072,N_6578);
xor U7240 (N_7240,N_6953,N_6344);
or U7241 (N_7241,N_6703,N_6885);
nor U7242 (N_7242,N_6397,N_6096);
or U7243 (N_7243,N_6938,N_6153);
or U7244 (N_7244,N_6208,N_6261);
or U7245 (N_7245,N_6196,N_6782);
and U7246 (N_7246,N_6555,N_6476);
nor U7247 (N_7247,N_6562,N_6931);
xor U7248 (N_7248,N_6811,N_6685);
or U7249 (N_7249,N_6622,N_6457);
and U7250 (N_7250,N_6277,N_6492);
and U7251 (N_7251,N_6446,N_6018);
nand U7252 (N_7252,N_6929,N_6129);
or U7253 (N_7253,N_6358,N_6783);
or U7254 (N_7254,N_6845,N_6749);
nor U7255 (N_7255,N_6005,N_6991);
and U7256 (N_7256,N_6777,N_6033);
or U7257 (N_7257,N_6220,N_6112);
nand U7258 (N_7258,N_6414,N_6537);
nand U7259 (N_7259,N_6518,N_6371);
and U7260 (N_7260,N_6796,N_6120);
nor U7261 (N_7261,N_6918,N_6552);
and U7262 (N_7262,N_6416,N_6247);
and U7263 (N_7263,N_6876,N_6539);
xnor U7264 (N_7264,N_6341,N_6183);
xnor U7265 (N_7265,N_6738,N_6145);
xor U7266 (N_7266,N_6952,N_6104);
or U7267 (N_7267,N_6740,N_6136);
nor U7268 (N_7268,N_6368,N_6299);
and U7269 (N_7269,N_6985,N_6852);
xnor U7270 (N_7270,N_6409,N_6023);
and U7271 (N_7271,N_6569,N_6282);
and U7272 (N_7272,N_6124,N_6055);
or U7273 (N_7273,N_6828,N_6444);
or U7274 (N_7274,N_6099,N_6415);
and U7275 (N_7275,N_6288,N_6310);
and U7276 (N_7276,N_6254,N_6824);
nor U7277 (N_7277,N_6498,N_6815);
nor U7278 (N_7278,N_6652,N_6693);
xnor U7279 (N_7279,N_6707,N_6503);
nor U7280 (N_7280,N_6790,N_6179);
and U7281 (N_7281,N_6249,N_6362);
or U7282 (N_7282,N_6978,N_6474);
nor U7283 (N_7283,N_6429,N_6851);
or U7284 (N_7284,N_6848,N_6257);
nand U7285 (N_7285,N_6351,N_6604);
or U7286 (N_7286,N_6213,N_6944);
or U7287 (N_7287,N_6826,N_6026);
and U7288 (N_7288,N_6427,N_6720);
nand U7289 (N_7289,N_6171,N_6580);
xor U7290 (N_7290,N_6892,N_6287);
or U7291 (N_7291,N_6558,N_6263);
and U7292 (N_7292,N_6883,N_6178);
or U7293 (N_7293,N_6647,N_6098);
and U7294 (N_7294,N_6191,N_6374);
xnor U7295 (N_7295,N_6306,N_6173);
nor U7296 (N_7296,N_6440,N_6291);
nor U7297 (N_7297,N_6349,N_6841);
nor U7298 (N_7298,N_6653,N_6475);
xor U7299 (N_7299,N_6849,N_6501);
xnor U7300 (N_7300,N_6085,N_6463);
nor U7301 (N_7301,N_6400,N_6354);
or U7302 (N_7302,N_6094,N_6076);
and U7303 (N_7303,N_6789,N_6376);
nor U7304 (N_7304,N_6650,N_6500);
and U7305 (N_7305,N_6393,N_6971);
nand U7306 (N_7306,N_6057,N_6955);
and U7307 (N_7307,N_6011,N_6258);
nand U7308 (N_7308,N_6357,N_6188);
or U7309 (N_7309,N_6311,N_6821);
and U7310 (N_7310,N_6161,N_6747);
nand U7311 (N_7311,N_6884,N_6915);
nor U7312 (N_7312,N_6843,N_6107);
or U7313 (N_7313,N_6139,N_6716);
nor U7314 (N_7314,N_6450,N_6816);
nor U7315 (N_7315,N_6143,N_6966);
or U7316 (N_7316,N_6780,N_6960);
and U7317 (N_7317,N_6121,N_6035);
nand U7318 (N_7318,N_6732,N_6644);
xnor U7319 (N_7319,N_6204,N_6951);
nand U7320 (N_7320,N_6158,N_6937);
xor U7321 (N_7321,N_6792,N_6223);
or U7322 (N_7322,N_6704,N_6221);
or U7323 (N_7323,N_6482,N_6019);
nand U7324 (N_7324,N_6589,N_6365);
or U7325 (N_7325,N_6995,N_6775);
nor U7326 (N_7326,N_6611,N_6973);
nand U7327 (N_7327,N_6339,N_6437);
or U7328 (N_7328,N_6010,N_6741);
nor U7329 (N_7329,N_6086,N_6404);
nor U7330 (N_7330,N_6781,N_6051);
nor U7331 (N_7331,N_6499,N_6134);
nor U7332 (N_7332,N_6547,N_6398);
and U7333 (N_7333,N_6270,N_6779);
or U7334 (N_7334,N_6334,N_6246);
or U7335 (N_7335,N_6930,N_6629);
and U7336 (N_7336,N_6725,N_6032);
or U7337 (N_7337,N_6100,N_6544);
nand U7338 (N_7338,N_6060,N_6758);
nor U7339 (N_7339,N_6020,N_6765);
or U7340 (N_7340,N_6904,N_6238);
or U7341 (N_7341,N_6998,N_6256);
or U7342 (N_7342,N_6431,N_6721);
nor U7343 (N_7343,N_6328,N_6027);
nand U7344 (N_7344,N_6764,N_6401);
xor U7345 (N_7345,N_6859,N_6116);
nand U7346 (N_7346,N_6302,N_6582);
xnor U7347 (N_7347,N_6923,N_6723);
and U7348 (N_7348,N_6793,N_6957);
nor U7349 (N_7349,N_6649,N_6483);
or U7350 (N_7350,N_6637,N_6290);
nand U7351 (N_7351,N_6059,N_6853);
nor U7352 (N_7352,N_6560,N_6630);
nor U7353 (N_7353,N_6902,N_6866);
nand U7354 (N_7354,N_6105,N_6718);
nor U7355 (N_7355,N_6743,N_6056);
nand U7356 (N_7356,N_6609,N_6443);
xor U7357 (N_7357,N_6708,N_6068);
and U7358 (N_7358,N_6744,N_6914);
or U7359 (N_7359,N_6711,N_6798);
xnor U7360 (N_7360,N_6600,N_6511);
nor U7361 (N_7361,N_6182,N_6596);
nand U7362 (N_7362,N_6466,N_6676);
and U7363 (N_7363,N_6199,N_6091);
xor U7364 (N_7364,N_6888,N_6759);
and U7365 (N_7365,N_6757,N_6617);
nand U7366 (N_7366,N_6625,N_6505);
xor U7367 (N_7367,N_6399,N_6920);
nor U7368 (N_7368,N_6370,N_6897);
nor U7369 (N_7369,N_6459,N_6154);
xnor U7370 (N_7370,N_6799,N_6905);
or U7371 (N_7371,N_6232,N_6494);
nor U7372 (N_7372,N_6681,N_6293);
or U7373 (N_7373,N_6643,N_6395);
and U7374 (N_7374,N_6373,N_6203);
nor U7375 (N_7375,N_6236,N_6066);
and U7376 (N_7376,N_6473,N_6847);
nor U7377 (N_7377,N_6903,N_6496);
or U7378 (N_7378,N_6829,N_6281);
xor U7379 (N_7379,N_6088,N_6984);
nand U7380 (N_7380,N_6872,N_6797);
and U7381 (N_7381,N_6927,N_6080);
nor U7382 (N_7382,N_6092,N_6193);
xnor U7383 (N_7383,N_6488,N_6822);
or U7384 (N_7384,N_6567,N_6461);
or U7385 (N_7385,N_6948,N_6239);
xnor U7386 (N_7386,N_6224,N_6893);
xnor U7387 (N_7387,N_6378,N_6214);
nand U7388 (N_7388,N_6206,N_6106);
nor U7389 (N_7389,N_6813,N_6327);
nand U7390 (N_7390,N_6101,N_6788);
or U7391 (N_7391,N_6377,N_6543);
and U7392 (N_7392,N_6458,N_6423);
nand U7393 (N_7393,N_6584,N_6315);
xnor U7394 (N_7394,N_6706,N_6137);
nor U7395 (N_7395,N_6908,N_6624);
and U7396 (N_7396,N_6677,N_6634);
and U7397 (N_7397,N_6882,N_6380);
nand U7398 (N_7398,N_6756,N_6958);
xor U7399 (N_7399,N_6201,N_6195);
nor U7400 (N_7400,N_6762,N_6886);
nor U7401 (N_7401,N_6039,N_6149);
nand U7402 (N_7402,N_6329,N_6682);
or U7403 (N_7403,N_6839,N_6219);
nor U7404 (N_7404,N_6128,N_6651);
or U7405 (N_7405,N_6661,N_6891);
nand U7406 (N_7406,N_6587,N_6699);
and U7407 (N_7407,N_6260,N_6834);
nand U7408 (N_7408,N_6486,N_6309);
and U7409 (N_7409,N_6455,N_6939);
or U7410 (N_7410,N_6321,N_6229);
xnor U7411 (N_7411,N_6108,N_6313);
or U7412 (N_7412,N_6863,N_6576);
or U7413 (N_7413,N_6701,N_6988);
or U7414 (N_7414,N_6119,N_6022);
nor U7415 (N_7415,N_6662,N_6292);
xnor U7416 (N_7416,N_6801,N_6386);
or U7417 (N_7417,N_6200,N_6864);
xnor U7418 (N_7418,N_6959,N_6031);
nand U7419 (N_7419,N_6774,N_6956);
nor U7420 (N_7420,N_6760,N_6540);
xor U7421 (N_7421,N_6924,N_6525);
nand U7422 (N_7422,N_6932,N_6002);
nand U7423 (N_7423,N_6184,N_6147);
or U7424 (N_7424,N_6900,N_6663);
nand U7425 (N_7425,N_6062,N_6148);
xor U7426 (N_7426,N_6809,N_6521);
or U7427 (N_7427,N_6391,N_6113);
and U7428 (N_7428,N_6940,N_6355);
or U7429 (N_7429,N_6284,N_6818);
xnor U7430 (N_7430,N_6016,N_6150);
xor U7431 (N_7431,N_6493,N_6669);
or U7432 (N_7432,N_6943,N_6686);
or U7433 (N_7433,N_6532,N_6597);
xor U7434 (N_7434,N_6715,N_6151);
xnor U7435 (N_7435,N_6272,N_6726);
nand U7436 (N_7436,N_6230,N_6710);
or U7437 (N_7437,N_6772,N_6336);
or U7438 (N_7438,N_6047,N_6244);
xor U7439 (N_7439,N_6481,N_6017);
xor U7440 (N_7440,N_6303,N_6241);
and U7441 (N_7441,N_6058,N_6333);
nand U7442 (N_7442,N_6337,N_6823);
or U7443 (N_7443,N_6390,N_6623);
nand U7444 (N_7444,N_6660,N_6916);
nor U7445 (N_7445,N_6819,N_6795);
nand U7446 (N_7446,N_6078,N_6030);
and U7447 (N_7447,N_6987,N_6714);
or U7448 (N_7448,N_6252,N_6612);
xnor U7449 (N_7449,N_6785,N_6198);
nor U7450 (N_7450,N_6641,N_6215);
and U7451 (N_7451,N_6964,N_6497);
nand U7452 (N_7452,N_6449,N_6166);
nand U7453 (N_7453,N_6177,N_6285);
nor U7454 (N_7454,N_6778,N_6037);
nor U7455 (N_7455,N_6767,N_6593);
xnor U7456 (N_7456,N_6599,N_6343);
and U7457 (N_7457,N_6156,N_6090);
and U7458 (N_7458,N_6418,N_6694);
and U7459 (N_7459,N_6614,N_6109);
nor U7460 (N_7460,N_6805,N_6424);
and U7461 (N_7461,N_6348,N_6209);
xor U7462 (N_7462,N_6942,N_6719);
xor U7463 (N_7463,N_6345,N_6679);
and U7464 (N_7464,N_6633,N_6761);
nor U7465 (N_7465,N_6231,N_6093);
and U7466 (N_7466,N_6082,N_6053);
or U7467 (N_7467,N_6434,N_6265);
and U7468 (N_7468,N_6591,N_6259);
or U7469 (N_7469,N_6827,N_6935);
xor U7470 (N_7470,N_6342,N_6753);
nand U7471 (N_7471,N_6388,N_6211);
or U7472 (N_7472,N_6318,N_6159);
or U7473 (N_7473,N_6425,N_6338);
and U7474 (N_7474,N_6628,N_6103);
nand U7475 (N_7475,N_6528,N_6006);
nor U7476 (N_7476,N_6267,N_6366);
and U7477 (N_7477,N_6095,N_6854);
nand U7478 (N_7478,N_6690,N_6901);
xnor U7479 (N_7479,N_6632,N_6009);
or U7480 (N_7480,N_6620,N_6324);
nor U7481 (N_7481,N_6933,N_6084);
and U7482 (N_7482,N_6636,N_6879);
and U7483 (N_7483,N_6469,N_6862);
and U7484 (N_7484,N_6837,N_6041);
nor U7485 (N_7485,N_6870,N_6737);
or U7486 (N_7486,N_6317,N_6160);
and U7487 (N_7487,N_6655,N_6585);
xnor U7488 (N_7488,N_6172,N_6527);
xor U7489 (N_7489,N_6586,N_6462);
nor U7490 (N_7490,N_6491,N_6934);
nand U7491 (N_7491,N_6130,N_6007);
xnor U7492 (N_7492,N_6817,N_6442);
nor U7493 (N_7493,N_6226,N_6590);
or U7494 (N_7494,N_6248,N_6250);
nand U7495 (N_7495,N_6999,N_6975);
nor U7496 (N_7496,N_6709,N_6594);
xor U7497 (N_7497,N_6990,N_6326);
xnor U7498 (N_7498,N_6353,N_6717);
and U7499 (N_7499,N_6513,N_6168);
and U7500 (N_7500,N_6620,N_6698);
nand U7501 (N_7501,N_6879,N_6672);
nand U7502 (N_7502,N_6183,N_6104);
nor U7503 (N_7503,N_6191,N_6993);
or U7504 (N_7504,N_6268,N_6056);
xor U7505 (N_7505,N_6925,N_6311);
and U7506 (N_7506,N_6356,N_6518);
xnor U7507 (N_7507,N_6244,N_6163);
or U7508 (N_7508,N_6598,N_6826);
or U7509 (N_7509,N_6442,N_6742);
or U7510 (N_7510,N_6629,N_6389);
xnor U7511 (N_7511,N_6198,N_6841);
nand U7512 (N_7512,N_6930,N_6205);
and U7513 (N_7513,N_6570,N_6565);
nand U7514 (N_7514,N_6927,N_6189);
nor U7515 (N_7515,N_6795,N_6694);
nor U7516 (N_7516,N_6798,N_6616);
and U7517 (N_7517,N_6708,N_6271);
nor U7518 (N_7518,N_6093,N_6171);
nor U7519 (N_7519,N_6115,N_6358);
nor U7520 (N_7520,N_6305,N_6492);
and U7521 (N_7521,N_6202,N_6389);
nor U7522 (N_7522,N_6238,N_6644);
nor U7523 (N_7523,N_6332,N_6683);
nor U7524 (N_7524,N_6753,N_6183);
nor U7525 (N_7525,N_6399,N_6747);
or U7526 (N_7526,N_6261,N_6378);
nor U7527 (N_7527,N_6835,N_6854);
and U7528 (N_7528,N_6491,N_6938);
or U7529 (N_7529,N_6124,N_6260);
or U7530 (N_7530,N_6076,N_6021);
nor U7531 (N_7531,N_6766,N_6199);
nor U7532 (N_7532,N_6619,N_6872);
xnor U7533 (N_7533,N_6956,N_6469);
nand U7534 (N_7534,N_6294,N_6785);
xnor U7535 (N_7535,N_6009,N_6362);
and U7536 (N_7536,N_6131,N_6416);
and U7537 (N_7537,N_6625,N_6301);
xor U7538 (N_7538,N_6379,N_6064);
xor U7539 (N_7539,N_6131,N_6230);
or U7540 (N_7540,N_6498,N_6484);
nor U7541 (N_7541,N_6278,N_6888);
nor U7542 (N_7542,N_6926,N_6618);
nor U7543 (N_7543,N_6069,N_6281);
xnor U7544 (N_7544,N_6221,N_6259);
nor U7545 (N_7545,N_6270,N_6175);
and U7546 (N_7546,N_6883,N_6833);
and U7547 (N_7547,N_6395,N_6121);
or U7548 (N_7548,N_6493,N_6417);
or U7549 (N_7549,N_6090,N_6362);
or U7550 (N_7550,N_6963,N_6243);
nand U7551 (N_7551,N_6632,N_6850);
or U7552 (N_7552,N_6588,N_6393);
nor U7553 (N_7553,N_6789,N_6308);
xnor U7554 (N_7554,N_6691,N_6579);
xnor U7555 (N_7555,N_6321,N_6313);
or U7556 (N_7556,N_6173,N_6053);
nor U7557 (N_7557,N_6430,N_6243);
nor U7558 (N_7558,N_6552,N_6139);
or U7559 (N_7559,N_6013,N_6970);
xnor U7560 (N_7560,N_6258,N_6420);
xor U7561 (N_7561,N_6237,N_6788);
nand U7562 (N_7562,N_6384,N_6247);
nor U7563 (N_7563,N_6365,N_6161);
nand U7564 (N_7564,N_6885,N_6081);
and U7565 (N_7565,N_6435,N_6350);
or U7566 (N_7566,N_6472,N_6331);
nor U7567 (N_7567,N_6663,N_6241);
nand U7568 (N_7568,N_6443,N_6346);
nor U7569 (N_7569,N_6359,N_6578);
nor U7570 (N_7570,N_6821,N_6637);
or U7571 (N_7571,N_6021,N_6335);
or U7572 (N_7572,N_6323,N_6351);
xnor U7573 (N_7573,N_6003,N_6944);
or U7574 (N_7574,N_6899,N_6289);
or U7575 (N_7575,N_6800,N_6245);
and U7576 (N_7576,N_6482,N_6070);
and U7577 (N_7577,N_6107,N_6958);
nor U7578 (N_7578,N_6787,N_6790);
and U7579 (N_7579,N_6737,N_6079);
and U7580 (N_7580,N_6159,N_6705);
and U7581 (N_7581,N_6038,N_6138);
xor U7582 (N_7582,N_6837,N_6132);
or U7583 (N_7583,N_6520,N_6308);
nand U7584 (N_7584,N_6341,N_6376);
nand U7585 (N_7585,N_6415,N_6181);
or U7586 (N_7586,N_6183,N_6625);
nor U7587 (N_7587,N_6917,N_6352);
nor U7588 (N_7588,N_6263,N_6859);
xor U7589 (N_7589,N_6728,N_6546);
and U7590 (N_7590,N_6197,N_6936);
or U7591 (N_7591,N_6907,N_6146);
or U7592 (N_7592,N_6188,N_6288);
nor U7593 (N_7593,N_6327,N_6438);
xnor U7594 (N_7594,N_6341,N_6009);
and U7595 (N_7595,N_6466,N_6121);
or U7596 (N_7596,N_6586,N_6858);
xor U7597 (N_7597,N_6150,N_6320);
or U7598 (N_7598,N_6852,N_6393);
nand U7599 (N_7599,N_6861,N_6023);
nor U7600 (N_7600,N_6061,N_6254);
and U7601 (N_7601,N_6133,N_6875);
nand U7602 (N_7602,N_6857,N_6292);
and U7603 (N_7603,N_6589,N_6068);
xnor U7604 (N_7604,N_6248,N_6429);
xor U7605 (N_7605,N_6458,N_6981);
xnor U7606 (N_7606,N_6877,N_6248);
nor U7607 (N_7607,N_6897,N_6963);
or U7608 (N_7608,N_6344,N_6952);
and U7609 (N_7609,N_6021,N_6477);
nor U7610 (N_7610,N_6606,N_6363);
xor U7611 (N_7611,N_6927,N_6069);
xnor U7612 (N_7612,N_6864,N_6519);
and U7613 (N_7613,N_6653,N_6058);
nand U7614 (N_7614,N_6827,N_6103);
and U7615 (N_7615,N_6406,N_6957);
xor U7616 (N_7616,N_6849,N_6050);
nand U7617 (N_7617,N_6340,N_6982);
nor U7618 (N_7618,N_6666,N_6646);
and U7619 (N_7619,N_6046,N_6868);
or U7620 (N_7620,N_6176,N_6046);
nand U7621 (N_7621,N_6899,N_6395);
xnor U7622 (N_7622,N_6744,N_6328);
xor U7623 (N_7623,N_6588,N_6330);
nand U7624 (N_7624,N_6279,N_6998);
and U7625 (N_7625,N_6779,N_6781);
xnor U7626 (N_7626,N_6624,N_6275);
xnor U7627 (N_7627,N_6784,N_6821);
xnor U7628 (N_7628,N_6378,N_6535);
nand U7629 (N_7629,N_6726,N_6782);
nor U7630 (N_7630,N_6428,N_6808);
or U7631 (N_7631,N_6805,N_6888);
and U7632 (N_7632,N_6175,N_6557);
xnor U7633 (N_7633,N_6847,N_6149);
xor U7634 (N_7634,N_6077,N_6961);
or U7635 (N_7635,N_6030,N_6837);
and U7636 (N_7636,N_6525,N_6119);
nor U7637 (N_7637,N_6350,N_6552);
nor U7638 (N_7638,N_6850,N_6796);
nand U7639 (N_7639,N_6384,N_6303);
and U7640 (N_7640,N_6577,N_6196);
xor U7641 (N_7641,N_6286,N_6991);
nand U7642 (N_7642,N_6810,N_6029);
nand U7643 (N_7643,N_6322,N_6017);
or U7644 (N_7644,N_6536,N_6589);
or U7645 (N_7645,N_6645,N_6899);
xnor U7646 (N_7646,N_6124,N_6624);
and U7647 (N_7647,N_6208,N_6918);
nand U7648 (N_7648,N_6945,N_6408);
nand U7649 (N_7649,N_6108,N_6717);
and U7650 (N_7650,N_6882,N_6973);
nor U7651 (N_7651,N_6729,N_6599);
xor U7652 (N_7652,N_6775,N_6962);
nand U7653 (N_7653,N_6903,N_6818);
nand U7654 (N_7654,N_6737,N_6032);
nor U7655 (N_7655,N_6344,N_6649);
or U7656 (N_7656,N_6830,N_6158);
nor U7657 (N_7657,N_6082,N_6930);
nand U7658 (N_7658,N_6255,N_6402);
xnor U7659 (N_7659,N_6586,N_6297);
nand U7660 (N_7660,N_6726,N_6096);
or U7661 (N_7661,N_6535,N_6318);
and U7662 (N_7662,N_6878,N_6074);
or U7663 (N_7663,N_6937,N_6966);
and U7664 (N_7664,N_6724,N_6188);
and U7665 (N_7665,N_6179,N_6822);
nor U7666 (N_7666,N_6131,N_6810);
and U7667 (N_7667,N_6487,N_6570);
nand U7668 (N_7668,N_6617,N_6806);
or U7669 (N_7669,N_6767,N_6391);
and U7670 (N_7670,N_6145,N_6324);
xor U7671 (N_7671,N_6269,N_6255);
xor U7672 (N_7672,N_6340,N_6149);
and U7673 (N_7673,N_6366,N_6879);
nor U7674 (N_7674,N_6805,N_6665);
and U7675 (N_7675,N_6253,N_6936);
nand U7676 (N_7676,N_6859,N_6965);
or U7677 (N_7677,N_6315,N_6018);
and U7678 (N_7678,N_6942,N_6785);
or U7679 (N_7679,N_6910,N_6847);
or U7680 (N_7680,N_6679,N_6453);
and U7681 (N_7681,N_6109,N_6736);
nor U7682 (N_7682,N_6244,N_6032);
or U7683 (N_7683,N_6284,N_6896);
and U7684 (N_7684,N_6906,N_6555);
nand U7685 (N_7685,N_6710,N_6195);
and U7686 (N_7686,N_6189,N_6688);
nand U7687 (N_7687,N_6590,N_6303);
and U7688 (N_7688,N_6482,N_6954);
xor U7689 (N_7689,N_6549,N_6835);
and U7690 (N_7690,N_6235,N_6759);
or U7691 (N_7691,N_6991,N_6887);
nor U7692 (N_7692,N_6973,N_6035);
or U7693 (N_7693,N_6299,N_6987);
nor U7694 (N_7694,N_6909,N_6243);
nand U7695 (N_7695,N_6986,N_6684);
nor U7696 (N_7696,N_6978,N_6181);
and U7697 (N_7697,N_6908,N_6013);
xnor U7698 (N_7698,N_6129,N_6109);
nand U7699 (N_7699,N_6160,N_6039);
xnor U7700 (N_7700,N_6377,N_6868);
or U7701 (N_7701,N_6655,N_6475);
nand U7702 (N_7702,N_6671,N_6398);
and U7703 (N_7703,N_6600,N_6234);
and U7704 (N_7704,N_6405,N_6901);
and U7705 (N_7705,N_6109,N_6443);
xor U7706 (N_7706,N_6408,N_6312);
nor U7707 (N_7707,N_6604,N_6271);
or U7708 (N_7708,N_6923,N_6710);
or U7709 (N_7709,N_6666,N_6661);
nand U7710 (N_7710,N_6305,N_6974);
and U7711 (N_7711,N_6734,N_6867);
xor U7712 (N_7712,N_6527,N_6618);
nand U7713 (N_7713,N_6174,N_6643);
nor U7714 (N_7714,N_6934,N_6984);
or U7715 (N_7715,N_6792,N_6524);
and U7716 (N_7716,N_6652,N_6980);
or U7717 (N_7717,N_6518,N_6825);
and U7718 (N_7718,N_6241,N_6025);
and U7719 (N_7719,N_6957,N_6188);
nor U7720 (N_7720,N_6726,N_6434);
or U7721 (N_7721,N_6471,N_6519);
and U7722 (N_7722,N_6580,N_6892);
xor U7723 (N_7723,N_6754,N_6467);
or U7724 (N_7724,N_6901,N_6149);
nor U7725 (N_7725,N_6136,N_6361);
nand U7726 (N_7726,N_6859,N_6680);
nand U7727 (N_7727,N_6784,N_6701);
or U7728 (N_7728,N_6551,N_6890);
nand U7729 (N_7729,N_6660,N_6849);
xnor U7730 (N_7730,N_6324,N_6130);
nor U7731 (N_7731,N_6140,N_6484);
and U7732 (N_7732,N_6981,N_6506);
nor U7733 (N_7733,N_6924,N_6602);
or U7734 (N_7734,N_6699,N_6131);
or U7735 (N_7735,N_6283,N_6947);
or U7736 (N_7736,N_6674,N_6020);
and U7737 (N_7737,N_6277,N_6932);
xnor U7738 (N_7738,N_6657,N_6975);
xor U7739 (N_7739,N_6289,N_6601);
or U7740 (N_7740,N_6836,N_6757);
or U7741 (N_7741,N_6964,N_6549);
nand U7742 (N_7742,N_6161,N_6417);
nor U7743 (N_7743,N_6890,N_6383);
and U7744 (N_7744,N_6921,N_6658);
xnor U7745 (N_7745,N_6274,N_6270);
and U7746 (N_7746,N_6633,N_6788);
and U7747 (N_7747,N_6843,N_6941);
or U7748 (N_7748,N_6070,N_6742);
xnor U7749 (N_7749,N_6246,N_6241);
xor U7750 (N_7750,N_6101,N_6580);
xnor U7751 (N_7751,N_6817,N_6126);
nor U7752 (N_7752,N_6057,N_6117);
or U7753 (N_7753,N_6993,N_6653);
xor U7754 (N_7754,N_6822,N_6077);
nor U7755 (N_7755,N_6726,N_6739);
or U7756 (N_7756,N_6155,N_6756);
xnor U7757 (N_7757,N_6311,N_6532);
xnor U7758 (N_7758,N_6172,N_6684);
xor U7759 (N_7759,N_6716,N_6486);
or U7760 (N_7760,N_6924,N_6442);
nand U7761 (N_7761,N_6571,N_6089);
nor U7762 (N_7762,N_6814,N_6436);
and U7763 (N_7763,N_6179,N_6240);
and U7764 (N_7764,N_6581,N_6498);
nand U7765 (N_7765,N_6218,N_6766);
nor U7766 (N_7766,N_6568,N_6074);
xnor U7767 (N_7767,N_6709,N_6035);
nand U7768 (N_7768,N_6874,N_6087);
or U7769 (N_7769,N_6172,N_6168);
or U7770 (N_7770,N_6153,N_6691);
and U7771 (N_7771,N_6609,N_6242);
and U7772 (N_7772,N_6900,N_6528);
nor U7773 (N_7773,N_6616,N_6976);
nand U7774 (N_7774,N_6784,N_6797);
nor U7775 (N_7775,N_6949,N_6506);
nand U7776 (N_7776,N_6700,N_6673);
and U7777 (N_7777,N_6417,N_6273);
or U7778 (N_7778,N_6651,N_6630);
nand U7779 (N_7779,N_6767,N_6756);
or U7780 (N_7780,N_6577,N_6038);
or U7781 (N_7781,N_6065,N_6696);
or U7782 (N_7782,N_6936,N_6678);
xor U7783 (N_7783,N_6951,N_6456);
or U7784 (N_7784,N_6106,N_6205);
nor U7785 (N_7785,N_6366,N_6774);
nor U7786 (N_7786,N_6009,N_6700);
and U7787 (N_7787,N_6515,N_6300);
or U7788 (N_7788,N_6090,N_6982);
and U7789 (N_7789,N_6716,N_6138);
or U7790 (N_7790,N_6141,N_6687);
and U7791 (N_7791,N_6953,N_6549);
nand U7792 (N_7792,N_6511,N_6905);
nor U7793 (N_7793,N_6089,N_6946);
nor U7794 (N_7794,N_6699,N_6168);
xor U7795 (N_7795,N_6717,N_6071);
nand U7796 (N_7796,N_6818,N_6714);
xnor U7797 (N_7797,N_6197,N_6235);
xor U7798 (N_7798,N_6046,N_6399);
and U7799 (N_7799,N_6390,N_6955);
and U7800 (N_7800,N_6210,N_6035);
xnor U7801 (N_7801,N_6862,N_6706);
and U7802 (N_7802,N_6642,N_6540);
nor U7803 (N_7803,N_6741,N_6144);
or U7804 (N_7804,N_6336,N_6223);
nand U7805 (N_7805,N_6245,N_6408);
nand U7806 (N_7806,N_6740,N_6188);
and U7807 (N_7807,N_6413,N_6927);
nand U7808 (N_7808,N_6449,N_6685);
xnor U7809 (N_7809,N_6689,N_6796);
nand U7810 (N_7810,N_6511,N_6278);
xor U7811 (N_7811,N_6534,N_6681);
nand U7812 (N_7812,N_6790,N_6050);
nor U7813 (N_7813,N_6052,N_6714);
nand U7814 (N_7814,N_6971,N_6293);
nand U7815 (N_7815,N_6711,N_6634);
or U7816 (N_7816,N_6338,N_6098);
or U7817 (N_7817,N_6549,N_6321);
xnor U7818 (N_7818,N_6239,N_6861);
xnor U7819 (N_7819,N_6388,N_6714);
nor U7820 (N_7820,N_6354,N_6974);
and U7821 (N_7821,N_6411,N_6601);
nor U7822 (N_7822,N_6100,N_6061);
nand U7823 (N_7823,N_6830,N_6092);
or U7824 (N_7824,N_6064,N_6979);
xor U7825 (N_7825,N_6253,N_6202);
nor U7826 (N_7826,N_6869,N_6501);
nor U7827 (N_7827,N_6149,N_6191);
nor U7828 (N_7828,N_6928,N_6049);
or U7829 (N_7829,N_6161,N_6648);
nand U7830 (N_7830,N_6064,N_6536);
xor U7831 (N_7831,N_6385,N_6659);
nand U7832 (N_7832,N_6630,N_6067);
xnor U7833 (N_7833,N_6439,N_6450);
xnor U7834 (N_7834,N_6562,N_6024);
nor U7835 (N_7835,N_6542,N_6895);
nand U7836 (N_7836,N_6176,N_6923);
and U7837 (N_7837,N_6764,N_6633);
or U7838 (N_7838,N_6814,N_6956);
and U7839 (N_7839,N_6862,N_6279);
and U7840 (N_7840,N_6380,N_6154);
nand U7841 (N_7841,N_6434,N_6414);
nor U7842 (N_7842,N_6298,N_6831);
nand U7843 (N_7843,N_6868,N_6646);
and U7844 (N_7844,N_6433,N_6588);
nor U7845 (N_7845,N_6552,N_6964);
nand U7846 (N_7846,N_6054,N_6680);
nor U7847 (N_7847,N_6322,N_6551);
and U7848 (N_7848,N_6471,N_6756);
nor U7849 (N_7849,N_6180,N_6349);
and U7850 (N_7850,N_6313,N_6604);
xor U7851 (N_7851,N_6993,N_6195);
nor U7852 (N_7852,N_6950,N_6260);
xor U7853 (N_7853,N_6083,N_6637);
nor U7854 (N_7854,N_6272,N_6231);
or U7855 (N_7855,N_6907,N_6607);
xor U7856 (N_7856,N_6324,N_6772);
or U7857 (N_7857,N_6847,N_6556);
and U7858 (N_7858,N_6606,N_6154);
and U7859 (N_7859,N_6268,N_6042);
and U7860 (N_7860,N_6141,N_6604);
nor U7861 (N_7861,N_6738,N_6903);
nor U7862 (N_7862,N_6325,N_6986);
and U7863 (N_7863,N_6079,N_6761);
nor U7864 (N_7864,N_6015,N_6587);
or U7865 (N_7865,N_6084,N_6953);
or U7866 (N_7866,N_6551,N_6401);
nand U7867 (N_7867,N_6162,N_6174);
or U7868 (N_7868,N_6770,N_6760);
or U7869 (N_7869,N_6107,N_6509);
nand U7870 (N_7870,N_6993,N_6368);
nor U7871 (N_7871,N_6546,N_6392);
xor U7872 (N_7872,N_6700,N_6086);
nor U7873 (N_7873,N_6062,N_6459);
nand U7874 (N_7874,N_6647,N_6014);
nor U7875 (N_7875,N_6035,N_6217);
or U7876 (N_7876,N_6737,N_6354);
nor U7877 (N_7877,N_6741,N_6708);
nand U7878 (N_7878,N_6525,N_6918);
xor U7879 (N_7879,N_6122,N_6563);
nand U7880 (N_7880,N_6509,N_6860);
nand U7881 (N_7881,N_6072,N_6859);
nor U7882 (N_7882,N_6473,N_6543);
nor U7883 (N_7883,N_6232,N_6376);
and U7884 (N_7884,N_6145,N_6399);
xnor U7885 (N_7885,N_6734,N_6108);
xor U7886 (N_7886,N_6121,N_6064);
nand U7887 (N_7887,N_6452,N_6061);
nand U7888 (N_7888,N_6432,N_6735);
xnor U7889 (N_7889,N_6480,N_6703);
nor U7890 (N_7890,N_6638,N_6071);
xor U7891 (N_7891,N_6599,N_6228);
xnor U7892 (N_7892,N_6757,N_6814);
nand U7893 (N_7893,N_6298,N_6670);
nor U7894 (N_7894,N_6591,N_6511);
nor U7895 (N_7895,N_6001,N_6364);
nand U7896 (N_7896,N_6743,N_6210);
xor U7897 (N_7897,N_6624,N_6997);
or U7898 (N_7898,N_6042,N_6265);
nand U7899 (N_7899,N_6786,N_6693);
xnor U7900 (N_7900,N_6840,N_6011);
nor U7901 (N_7901,N_6966,N_6463);
or U7902 (N_7902,N_6093,N_6341);
or U7903 (N_7903,N_6125,N_6013);
and U7904 (N_7904,N_6849,N_6534);
nor U7905 (N_7905,N_6858,N_6556);
or U7906 (N_7906,N_6704,N_6073);
or U7907 (N_7907,N_6600,N_6868);
nand U7908 (N_7908,N_6434,N_6024);
and U7909 (N_7909,N_6152,N_6586);
nand U7910 (N_7910,N_6155,N_6834);
nand U7911 (N_7911,N_6921,N_6900);
or U7912 (N_7912,N_6471,N_6657);
nand U7913 (N_7913,N_6495,N_6857);
nand U7914 (N_7914,N_6916,N_6086);
xor U7915 (N_7915,N_6698,N_6664);
xnor U7916 (N_7916,N_6238,N_6416);
xor U7917 (N_7917,N_6112,N_6406);
and U7918 (N_7918,N_6463,N_6373);
or U7919 (N_7919,N_6451,N_6560);
and U7920 (N_7920,N_6384,N_6859);
nand U7921 (N_7921,N_6334,N_6372);
or U7922 (N_7922,N_6457,N_6387);
xor U7923 (N_7923,N_6147,N_6867);
nor U7924 (N_7924,N_6421,N_6433);
and U7925 (N_7925,N_6171,N_6636);
nand U7926 (N_7926,N_6646,N_6910);
nand U7927 (N_7927,N_6506,N_6799);
xor U7928 (N_7928,N_6714,N_6994);
and U7929 (N_7929,N_6790,N_6818);
nand U7930 (N_7930,N_6636,N_6424);
or U7931 (N_7931,N_6219,N_6951);
and U7932 (N_7932,N_6974,N_6183);
xnor U7933 (N_7933,N_6112,N_6491);
and U7934 (N_7934,N_6049,N_6985);
xnor U7935 (N_7935,N_6278,N_6427);
or U7936 (N_7936,N_6699,N_6580);
or U7937 (N_7937,N_6956,N_6614);
xor U7938 (N_7938,N_6582,N_6985);
nand U7939 (N_7939,N_6879,N_6634);
and U7940 (N_7940,N_6294,N_6381);
nor U7941 (N_7941,N_6485,N_6802);
nand U7942 (N_7942,N_6906,N_6325);
or U7943 (N_7943,N_6871,N_6975);
nor U7944 (N_7944,N_6925,N_6002);
or U7945 (N_7945,N_6899,N_6366);
xnor U7946 (N_7946,N_6043,N_6554);
xnor U7947 (N_7947,N_6052,N_6119);
nand U7948 (N_7948,N_6416,N_6271);
xor U7949 (N_7949,N_6252,N_6722);
xor U7950 (N_7950,N_6156,N_6206);
and U7951 (N_7951,N_6209,N_6912);
nand U7952 (N_7952,N_6421,N_6419);
or U7953 (N_7953,N_6807,N_6816);
and U7954 (N_7954,N_6349,N_6253);
and U7955 (N_7955,N_6701,N_6351);
or U7956 (N_7956,N_6208,N_6925);
or U7957 (N_7957,N_6359,N_6373);
xnor U7958 (N_7958,N_6239,N_6872);
and U7959 (N_7959,N_6933,N_6273);
nor U7960 (N_7960,N_6188,N_6778);
and U7961 (N_7961,N_6087,N_6534);
and U7962 (N_7962,N_6917,N_6210);
and U7963 (N_7963,N_6156,N_6865);
and U7964 (N_7964,N_6122,N_6508);
nand U7965 (N_7965,N_6139,N_6525);
nor U7966 (N_7966,N_6217,N_6431);
xor U7967 (N_7967,N_6103,N_6716);
xnor U7968 (N_7968,N_6491,N_6956);
or U7969 (N_7969,N_6386,N_6151);
xor U7970 (N_7970,N_6498,N_6111);
and U7971 (N_7971,N_6886,N_6223);
xor U7972 (N_7972,N_6790,N_6884);
and U7973 (N_7973,N_6255,N_6655);
xor U7974 (N_7974,N_6905,N_6810);
and U7975 (N_7975,N_6541,N_6276);
nand U7976 (N_7976,N_6487,N_6233);
nand U7977 (N_7977,N_6772,N_6234);
nand U7978 (N_7978,N_6283,N_6251);
and U7979 (N_7979,N_6321,N_6072);
nor U7980 (N_7980,N_6850,N_6837);
nor U7981 (N_7981,N_6054,N_6964);
xnor U7982 (N_7982,N_6665,N_6490);
nor U7983 (N_7983,N_6233,N_6297);
and U7984 (N_7984,N_6681,N_6295);
nor U7985 (N_7985,N_6203,N_6097);
or U7986 (N_7986,N_6020,N_6401);
and U7987 (N_7987,N_6638,N_6093);
nand U7988 (N_7988,N_6763,N_6261);
or U7989 (N_7989,N_6122,N_6218);
nor U7990 (N_7990,N_6477,N_6012);
xnor U7991 (N_7991,N_6847,N_6954);
or U7992 (N_7992,N_6606,N_6804);
nor U7993 (N_7993,N_6224,N_6490);
and U7994 (N_7994,N_6199,N_6830);
or U7995 (N_7995,N_6484,N_6077);
or U7996 (N_7996,N_6849,N_6377);
nor U7997 (N_7997,N_6648,N_6268);
or U7998 (N_7998,N_6448,N_6192);
and U7999 (N_7999,N_6261,N_6613);
and U8000 (N_8000,N_7480,N_7913);
nor U8001 (N_8001,N_7000,N_7532);
nor U8002 (N_8002,N_7168,N_7378);
and U8003 (N_8003,N_7051,N_7384);
nand U8004 (N_8004,N_7368,N_7283);
xor U8005 (N_8005,N_7839,N_7096);
nand U8006 (N_8006,N_7521,N_7109);
or U8007 (N_8007,N_7766,N_7273);
or U8008 (N_8008,N_7530,N_7652);
nor U8009 (N_8009,N_7185,N_7202);
and U8010 (N_8010,N_7927,N_7563);
and U8011 (N_8011,N_7551,N_7830);
nand U8012 (N_8012,N_7523,N_7298);
xor U8013 (N_8013,N_7812,N_7498);
nor U8014 (N_8014,N_7990,N_7760);
nand U8015 (N_8015,N_7325,N_7542);
nand U8016 (N_8016,N_7092,N_7166);
nand U8017 (N_8017,N_7441,N_7969);
or U8018 (N_8018,N_7728,N_7123);
xnor U8019 (N_8019,N_7741,N_7395);
or U8020 (N_8020,N_7949,N_7677);
xnor U8021 (N_8021,N_7425,N_7831);
nand U8022 (N_8022,N_7189,N_7948);
nand U8023 (N_8023,N_7186,N_7516);
and U8024 (N_8024,N_7914,N_7783);
or U8025 (N_8025,N_7009,N_7377);
nand U8026 (N_8026,N_7869,N_7991);
xnor U8027 (N_8027,N_7236,N_7287);
nand U8028 (N_8028,N_7014,N_7788);
nor U8029 (N_8029,N_7928,N_7689);
nor U8030 (N_8030,N_7870,N_7450);
or U8031 (N_8031,N_7187,N_7809);
and U8032 (N_8032,N_7538,N_7278);
and U8033 (N_8033,N_7912,N_7889);
nor U8034 (N_8034,N_7755,N_7505);
nand U8035 (N_8035,N_7258,N_7864);
or U8036 (N_8036,N_7041,N_7672);
and U8037 (N_8037,N_7122,N_7796);
nand U8038 (N_8038,N_7445,N_7940);
or U8039 (N_8039,N_7644,N_7238);
xor U8040 (N_8040,N_7178,N_7686);
or U8041 (N_8041,N_7607,N_7582);
or U8042 (N_8042,N_7827,N_7408);
xnor U8043 (N_8043,N_7054,N_7294);
nand U8044 (N_8044,N_7348,N_7361);
nand U8045 (N_8045,N_7331,N_7112);
nand U8046 (N_8046,N_7555,N_7793);
xor U8047 (N_8047,N_7587,N_7265);
nor U8048 (N_8048,N_7225,N_7194);
and U8049 (N_8049,N_7808,N_7525);
or U8050 (N_8050,N_7289,N_7110);
nor U8051 (N_8051,N_7872,N_7972);
nor U8052 (N_8052,N_7782,N_7873);
nand U8053 (N_8053,N_7199,N_7806);
nand U8054 (N_8054,N_7321,N_7704);
or U8055 (N_8055,N_7860,N_7547);
or U8056 (N_8056,N_7753,N_7814);
and U8057 (N_8057,N_7739,N_7623);
or U8058 (N_8058,N_7577,N_7581);
xnor U8059 (N_8059,N_7127,N_7633);
nand U8060 (N_8060,N_7917,N_7039);
nand U8061 (N_8061,N_7299,N_7107);
nand U8062 (N_8062,N_7443,N_7971);
and U8063 (N_8063,N_7130,N_7825);
and U8064 (N_8064,N_7217,N_7484);
nor U8065 (N_8065,N_7897,N_7098);
and U8066 (N_8066,N_7879,N_7787);
or U8067 (N_8067,N_7474,N_7459);
or U8068 (N_8068,N_7124,N_7192);
nor U8069 (N_8069,N_7144,N_7430);
or U8070 (N_8070,N_7863,N_7619);
and U8071 (N_8071,N_7550,N_7664);
nand U8072 (N_8072,N_7399,N_7492);
or U8073 (N_8073,N_7257,N_7841);
and U8074 (N_8074,N_7737,N_7840);
nand U8075 (N_8075,N_7218,N_7875);
nand U8076 (N_8076,N_7167,N_7013);
or U8077 (N_8077,N_7479,N_7026);
or U8078 (N_8078,N_7993,N_7336);
nand U8079 (N_8079,N_7703,N_7763);
and U8080 (N_8080,N_7434,N_7502);
nand U8081 (N_8081,N_7485,N_7506);
nand U8082 (N_8082,N_7093,N_7082);
nand U8083 (N_8083,N_7409,N_7277);
and U8084 (N_8084,N_7680,N_7396);
nor U8085 (N_8085,N_7132,N_7345);
xnor U8086 (N_8086,N_7081,N_7919);
or U8087 (N_8087,N_7922,N_7779);
nor U8088 (N_8088,N_7557,N_7448);
xor U8089 (N_8089,N_7416,N_7161);
or U8090 (N_8090,N_7822,N_7259);
xnor U8091 (N_8091,N_7031,N_7747);
and U8092 (N_8092,N_7648,N_7269);
or U8093 (N_8093,N_7180,N_7835);
xnor U8094 (N_8094,N_7805,N_7744);
nor U8095 (N_8095,N_7359,N_7250);
and U8096 (N_8096,N_7526,N_7926);
and U8097 (N_8097,N_7973,N_7529);
nor U8098 (N_8098,N_7415,N_7335);
and U8099 (N_8099,N_7288,N_7896);
nand U8100 (N_8100,N_7383,N_7137);
xnor U8101 (N_8101,N_7233,N_7791);
xor U8102 (N_8102,N_7893,N_7354);
or U8103 (N_8103,N_7169,N_7007);
nand U8104 (N_8104,N_7309,N_7724);
nand U8105 (N_8105,N_7438,N_7757);
and U8106 (N_8106,N_7956,N_7876);
nor U8107 (N_8107,N_7346,N_7905);
or U8108 (N_8108,N_7702,N_7540);
and U8109 (N_8109,N_7967,N_7586);
or U8110 (N_8110,N_7908,N_7799);
xor U8111 (N_8111,N_7726,N_7121);
nor U8112 (N_8112,N_7952,N_7073);
xnor U8113 (N_8113,N_7074,N_7100);
and U8114 (N_8114,N_7979,N_7866);
xnor U8115 (N_8115,N_7861,N_7413);
nor U8116 (N_8116,N_7997,N_7018);
and U8117 (N_8117,N_7235,N_7903);
or U8118 (N_8118,N_7360,N_7155);
or U8119 (N_8119,N_7291,N_7974);
and U8120 (N_8120,N_7575,N_7646);
nand U8121 (N_8121,N_7695,N_7609);
xnor U8122 (N_8122,N_7823,N_7687);
nor U8123 (N_8123,N_7011,N_7647);
nand U8124 (N_8124,N_7350,N_7950);
nor U8125 (N_8125,N_7770,N_7135);
or U8126 (N_8126,N_7150,N_7153);
and U8127 (N_8127,N_7171,N_7848);
xor U8128 (N_8128,N_7663,N_7820);
xor U8129 (N_8129,N_7397,N_7337);
nand U8130 (N_8130,N_7320,N_7691);
nor U8131 (N_8131,N_7314,N_7639);
nor U8132 (N_8132,N_7865,N_7804);
nor U8133 (N_8133,N_7732,N_7572);
and U8134 (N_8134,N_7426,N_7427);
nor U8135 (N_8135,N_7157,N_7198);
or U8136 (N_8136,N_7482,N_7892);
and U8137 (N_8137,N_7057,N_7936);
and U8138 (N_8138,N_7855,N_7681);
nor U8139 (N_8139,N_7115,N_7069);
nor U8140 (N_8140,N_7232,N_7548);
nor U8141 (N_8141,N_7945,N_7984);
nor U8142 (N_8142,N_7877,N_7583);
xnor U8143 (N_8143,N_7419,N_7570);
or U8144 (N_8144,N_7898,N_7657);
nand U8145 (N_8145,N_7992,N_7758);
nor U8146 (N_8146,N_7802,N_7683);
and U8147 (N_8147,N_7684,N_7352);
nor U8148 (N_8148,N_7095,N_7671);
and U8149 (N_8149,N_7666,N_7735);
xor U8150 (N_8150,N_7608,N_7322);
xnor U8151 (N_8151,N_7565,N_7637);
nor U8152 (N_8152,N_7669,N_7097);
nor U8153 (N_8153,N_7446,N_7519);
nand U8154 (N_8154,N_7227,N_7676);
and U8155 (N_8155,N_7906,N_7264);
or U8156 (N_8156,N_7308,N_7980);
and U8157 (N_8157,N_7837,N_7078);
or U8158 (N_8158,N_7317,N_7491);
and U8159 (N_8159,N_7296,N_7718);
or U8160 (N_8160,N_7181,N_7206);
xnor U8161 (N_8161,N_7310,N_7544);
or U8162 (N_8162,N_7024,N_7182);
and U8163 (N_8163,N_7595,N_7602);
nand U8164 (N_8164,N_7077,N_7442);
and U8165 (N_8165,N_7094,N_7696);
nand U8166 (N_8166,N_7151,N_7414);
or U8167 (N_8167,N_7716,N_7638);
and U8168 (N_8168,N_7773,N_7590);
and U8169 (N_8169,N_7566,N_7088);
or U8170 (N_8170,N_7392,N_7966);
or U8171 (N_8171,N_7968,N_7142);
nand U8172 (N_8172,N_7549,N_7842);
and U8173 (N_8173,N_7759,N_7931);
xor U8174 (N_8174,N_7829,N_7072);
xor U8175 (N_8175,N_7909,N_7682);
nor U8176 (N_8176,N_7154,N_7133);
nand U8177 (N_8177,N_7473,N_7915);
nand U8178 (N_8178,N_7522,N_7003);
nand U8179 (N_8179,N_7164,N_7247);
and U8180 (N_8180,N_7828,N_7868);
and U8181 (N_8181,N_7622,N_7105);
nand U8182 (N_8182,N_7838,N_7483);
nand U8183 (N_8183,N_7528,N_7047);
xor U8184 (N_8184,N_7036,N_7929);
nor U8185 (N_8185,N_7748,N_7836);
or U8186 (N_8186,N_7537,N_7674);
or U8187 (N_8187,N_7717,N_7811);
nor U8188 (N_8188,N_7636,N_7297);
nor U8189 (N_8189,N_7162,N_7103);
nor U8190 (N_8190,N_7500,N_7784);
and U8191 (N_8191,N_7319,N_7601);
nor U8192 (N_8192,N_7710,N_7947);
or U8193 (N_8193,N_7813,N_7719);
or U8194 (N_8194,N_7375,N_7714);
nand U8195 (N_8195,N_7824,N_7944);
xnor U8196 (N_8196,N_7631,N_7785);
and U8197 (N_8197,N_7561,N_7329);
xor U8198 (N_8198,N_7670,N_7571);
nand U8199 (N_8199,N_7721,N_7497);
nand U8200 (N_8200,N_7584,N_7412);
or U8201 (N_8201,N_7251,N_7025);
xnor U8202 (N_8202,N_7934,N_7776);
nor U8203 (N_8203,N_7985,N_7501);
nor U8204 (N_8204,N_7079,N_7156);
or U8205 (N_8205,N_7006,N_7986);
and U8206 (N_8206,N_7274,N_7351);
nor U8207 (N_8207,N_7918,N_7372);
and U8208 (N_8208,N_7055,N_7578);
or U8209 (N_8209,N_7076,N_7645);
nor U8210 (N_8210,N_7270,N_7790);
nor U8211 (N_8211,N_7514,N_7001);
nand U8212 (N_8212,N_7699,N_7859);
nor U8213 (N_8213,N_7512,N_7111);
nand U8214 (N_8214,N_7675,N_7924);
xnor U8215 (N_8215,N_7508,N_7205);
xor U8216 (N_8216,N_7316,N_7126);
and U8217 (N_8217,N_7567,N_7761);
xor U8218 (N_8218,N_7116,N_7436);
nor U8219 (N_8219,N_7624,N_7471);
nor U8220 (N_8220,N_7428,N_7208);
and U8221 (N_8221,N_7874,N_7685);
xnor U8222 (N_8222,N_7052,N_7955);
xnor U8223 (N_8223,N_7226,N_7780);
xnor U8224 (N_8224,N_7883,N_7534);
nand U8225 (N_8225,N_7307,N_7743);
or U8226 (N_8226,N_7102,N_7768);
nand U8227 (N_8227,N_7580,N_7313);
xnor U8228 (N_8228,N_7511,N_7649);
nand U8229 (N_8229,N_7941,N_7591);
nand U8230 (N_8230,N_7943,N_7422);
xnor U8231 (N_8231,N_7745,N_7546);
nor U8232 (N_8232,N_7851,N_7452);
nor U8233 (N_8233,N_7708,N_7598);
nand U8234 (N_8234,N_7630,N_7890);
nor U8235 (N_8235,N_7911,N_7464);
nor U8236 (N_8236,N_7463,N_7230);
nor U8237 (N_8237,N_7460,N_7461);
and U8238 (N_8238,N_7810,N_7343);
nand U8239 (N_8239,N_7533,N_7056);
nor U8240 (N_8240,N_7362,N_7276);
xor U8241 (N_8241,N_7679,N_7946);
or U8242 (N_8242,N_7357,N_7754);
or U8243 (N_8243,N_7641,N_7113);
and U8244 (N_8244,N_7462,N_7794);
and U8245 (N_8245,N_7120,N_7900);
xnor U8246 (N_8246,N_7170,N_7381);
nor U8247 (N_8247,N_7020,N_7141);
xor U8248 (N_8248,N_7290,N_7267);
or U8249 (N_8249,N_7959,N_7494);
xor U8250 (N_8250,N_7282,N_7213);
xnor U8251 (N_8251,N_7970,N_7256);
nor U8252 (N_8252,N_7370,N_7140);
or U8253 (N_8253,N_7365,N_7531);
nor U8254 (N_8254,N_7059,N_7777);
and U8255 (N_8255,N_7191,N_7600);
xnor U8256 (N_8256,N_7742,N_7019);
nand U8257 (N_8257,N_7803,N_7261);
nand U8258 (N_8258,N_7035,N_7603);
or U8259 (N_8259,N_7939,N_7470);
nor U8260 (N_8260,N_7469,N_7173);
nand U8261 (N_8261,N_7423,N_7240);
nand U8262 (N_8262,N_7216,N_7618);
or U8263 (N_8263,N_7552,N_7148);
nand U8264 (N_8264,N_7143,N_7243);
nand U8265 (N_8265,N_7032,N_7962);
xor U8266 (N_8266,N_7465,N_7882);
nand U8267 (N_8267,N_7987,N_7615);
nor U8268 (N_8268,N_7612,N_7106);
nor U8269 (N_8269,N_7579,N_7064);
or U8270 (N_8270,N_7209,N_7040);
and U8271 (N_8271,N_7885,N_7751);
nor U8272 (N_8272,N_7342,N_7499);
nand U8273 (N_8273,N_7231,N_7517);
or U8274 (N_8274,N_7543,N_7453);
nor U8275 (N_8275,N_7058,N_7574);
xor U8276 (N_8276,N_7978,N_7087);
nand U8277 (N_8277,N_7789,N_7312);
nand U8278 (N_8278,N_7108,N_7027);
nand U8279 (N_8279,N_7190,N_7203);
and U8280 (N_8280,N_7010,N_7642);
nand U8281 (N_8281,N_7017,N_7400);
and U8282 (N_8282,N_7042,N_7136);
or U8283 (N_8283,N_7558,N_7275);
and U8284 (N_8284,N_7228,N_7736);
and U8285 (N_8285,N_7858,N_7439);
nor U8286 (N_8286,N_7028,N_7844);
or U8287 (N_8287,N_7705,N_7589);
nand U8288 (N_8288,N_7196,N_7495);
xnor U8289 (N_8289,N_7421,N_7305);
nor U8290 (N_8290,N_7467,N_7300);
or U8291 (N_8291,N_7627,N_7099);
and U8292 (N_8292,N_7725,N_7071);
or U8293 (N_8293,N_7662,N_7921);
nand U8294 (N_8294,N_7070,N_7188);
nor U8295 (N_8295,N_7323,N_7554);
nor U8296 (N_8296,N_7746,N_7369);
and U8297 (N_8297,N_7951,N_7772);
nor U8298 (N_8298,N_7244,N_7435);
xor U8299 (N_8299,N_7617,N_7573);
and U8300 (N_8300,N_7472,N_7665);
or U8301 (N_8301,N_7061,N_7285);
xor U8302 (N_8302,N_7925,N_7424);
and U8303 (N_8303,N_7722,N_7458);
nor U8304 (N_8304,N_7324,N_7887);
nor U8305 (N_8305,N_7129,N_7286);
xor U8306 (N_8306,N_7701,N_7326);
and U8307 (N_8307,N_7711,N_7177);
or U8308 (N_8308,N_7393,N_7340);
and U8309 (N_8309,N_7447,N_7338);
nor U8310 (N_8310,N_7795,N_7653);
or U8311 (N_8311,N_7786,N_7332);
and U8312 (N_8312,N_7149,N_7847);
xnor U8313 (N_8313,N_7935,N_7139);
xor U8314 (N_8314,N_7594,N_7295);
xnor U8315 (N_8315,N_7654,N_7692);
or U8316 (N_8316,N_7084,N_7688);
nand U8317 (N_8317,N_7404,N_7886);
and U8318 (N_8318,N_7697,N_7698);
nor U8319 (N_8319,N_7942,N_7016);
nand U8320 (N_8320,N_7706,N_7049);
or U8321 (N_8321,N_7303,N_7128);
xor U8322 (N_8322,N_7431,N_7327);
or U8323 (N_8323,N_7733,N_7729);
nand U8324 (N_8324,N_7085,N_7982);
nor U8325 (N_8325,N_7576,N_7060);
or U8326 (N_8326,N_7953,N_7756);
nor U8327 (N_8327,N_7643,N_7988);
nor U8328 (N_8328,N_7388,N_7960);
nand U8329 (N_8329,N_7659,N_7560);
or U8330 (N_8330,N_7008,N_7596);
nor U8331 (N_8331,N_7819,N_7610);
xor U8332 (N_8332,N_7302,N_7311);
and U8333 (N_8333,N_7389,N_7373);
and U8334 (N_8334,N_7175,N_7901);
nand U8335 (N_8335,N_7067,N_7229);
or U8336 (N_8336,N_7660,N_7559);
xnor U8337 (N_8337,N_7632,N_7850);
and U8338 (N_8338,N_7403,N_7476);
nor U8339 (N_8339,N_7849,N_7138);
xnor U8340 (N_8340,N_7954,N_7260);
nor U8341 (N_8341,N_7821,N_7222);
nand U8342 (N_8342,N_7043,N_7564);
nand U8343 (N_8343,N_7486,N_7080);
nand U8344 (N_8344,N_7406,N_7268);
and U8345 (N_8345,N_7834,N_7022);
nand U8346 (N_8346,N_7158,N_7852);
or U8347 (N_8347,N_7998,N_7668);
xnor U8348 (N_8348,N_7355,N_7568);
and U8349 (N_8349,N_7983,N_7401);
xor U8350 (N_8350,N_7266,N_7380);
xnor U8351 (N_8351,N_7902,N_7503);
xor U8352 (N_8352,N_7449,N_7815);
nor U8353 (N_8353,N_7588,N_7977);
and U8354 (N_8354,N_7731,N_7493);
or U8355 (N_8355,N_7816,N_7005);
nand U8356 (N_8356,N_7881,N_7367);
and U8357 (N_8357,N_7920,N_7700);
nand U8358 (N_8358,N_7545,N_7125);
xnor U8359 (N_8359,N_7249,N_7147);
or U8360 (N_8360,N_7599,N_7239);
and U8361 (N_8361,N_7193,N_7817);
xnor U8362 (N_8362,N_7455,N_7690);
or U8363 (N_8363,N_7976,N_7002);
xnor U8364 (N_8364,N_7030,N_7650);
nor U8365 (N_8365,N_7541,N_7957);
xor U8366 (N_8366,N_7301,N_7279);
nand U8367 (N_8367,N_7363,N_7605);
xnor U8368 (N_8368,N_7798,N_7101);
and U8369 (N_8369,N_7775,N_7062);
and U8370 (N_8370,N_7224,N_7709);
and U8371 (N_8371,N_7723,N_7620);
xnor U8372 (N_8372,N_7520,N_7496);
and U8373 (N_8373,N_7242,N_7515);
nand U8374 (N_8374,N_7871,N_7562);
or U8375 (N_8375,N_7961,N_7420);
nor U8376 (N_8376,N_7195,N_7635);
or U8377 (N_8377,N_7488,N_7454);
nand U8378 (N_8378,N_7916,N_7904);
and U8379 (N_8379,N_7923,N_7104);
nand U8380 (N_8380,N_7958,N_7184);
nor U8381 (N_8381,N_7341,N_7767);
and U8382 (N_8382,N_7315,N_7405);
or U8383 (N_8383,N_7853,N_7214);
or U8384 (N_8384,N_7707,N_7801);
nor U8385 (N_8385,N_7625,N_7667);
or U8386 (N_8386,N_7174,N_7749);
and U8387 (N_8387,N_7457,N_7220);
and U8388 (N_8388,N_7781,N_7075);
xor U8389 (N_8389,N_7411,N_7163);
and U8390 (N_8390,N_7661,N_7524);
or U8391 (N_8391,N_7066,N_7366);
nor U8392 (N_8392,N_7358,N_7065);
xor U8393 (N_8393,N_7995,N_7390);
nand U8394 (N_8394,N_7353,N_7626);
or U8395 (N_8395,N_7328,N_7160);
nor U8396 (N_8396,N_7614,N_7539);
and U8397 (N_8397,N_7429,N_7179);
or U8398 (N_8398,N_7730,N_7857);
or U8399 (N_8399,N_7994,N_7629);
nand U8400 (N_8400,N_7818,N_7765);
xor U8401 (N_8401,N_7306,N_7391);
or U8402 (N_8402,N_7086,N_7553);
nor U8403 (N_8403,N_7255,N_7963);
and U8404 (N_8404,N_7262,N_7487);
or U8405 (N_8405,N_7234,N_7048);
nand U8406 (N_8406,N_7204,N_7063);
and U8407 (N_8407,N_7176,N_7930);
nor U8408 (N_8408,N_7621,N_7854);
nor U8409 (N_8409,N_7478,N_7693);
xnor U8410 (N_8410,N_7410,N_7440);
or U8411 (N_8411,N_7398,N_7527);
nand U8412 (N_8412,N_7907,N_7371);
and U8413 (N_8413,N_7826,N_7044);
and U8414 (N_8414,N_7089,N_7034);
nor U8415 (N_8415,N_7418,N_7385);
nor U8416 (N_8416,N_7867,N_7880);
xor U8417 (N_8417,N_7800,N_7715);
nand U8418 (N_8418,N_7933,N_7004);
nand U8419 (N_8419,N_7975,N_7432);
and U8420 (N_8420,N_7280,N_7640);
and U8421 (N_8421,N_7386,N_7509);
xor U8422 (N_8422,N_7965,N_7037);
or U8423 (N_8423,N_7376,N_7604);
nand U8424 (N_8424,N_7613,N_7658);
xnor U8425 (N_8425,N_7284,N_7489);
nor U8426 (N_8426,N_7253,N_7856);
nand U8427 (N_8427,N_7507,N_7475);
or U8428 (N_8428,N_7764,N_7333);
or U8429 (N_8429,N_7159,N_7845);
xor U8430 (N_8430,N_7263,N_7330);
nor U8431 (N_8431,N_7938,N_7029);
or U8432 (N_8432,N_7888,N_7752);
nor U8433 (N_8433,N_7021,N_7535);
or U8434 (N_8434,N_7556,N_7727);
nand U8435 (N_8435,N_7334,N_7481);
xor U8436 (N_8436,N_7884,N_7628);
nand U8437 (N_8437,N_7518,N_7083);
or U8438 (N_8438,N_7068,N_7281);
nand U8439 (N_8439,N_7797,N_7878);
or U8440 (N_8440,N_7114,N_7152);
and U8441 (N_8441,N_7616,N_7846);
nand U8442 (N_8442,N_7012,N_7349);
nand U8443 (N_8443,N_7272,N_7513);
or U8444 (N_8444,N_7510,N_7504);
and U8445 (N_8445,N_7477,N_7197);
nand U8446 (N_8446,N_7964,N_7118);
nor U8447 (N_8447,N_7678,N_7862);
xor U8448 (N_8448,N_7712,N_7091);
xor U8449 (N_8449,N_7145,N_7593);
and U8450 (N_8450,N_7356,N_7592);
and U8451 (N_8451,N_7673,N_7304);
nor U8452 (N_8452,N_7134,N_7932);
or U8453 (N_8453,N_7212,N_7651);
nand U8454 (N_8454,N_7117,N_7394);
or U8455 (N_8455,N_7456,N_7015);
nand U8456 (N_8456,N_7762,N_7750);
and U8457 (N_8457,N_7536,N_7387);
nor U8458 (N_8458,N_7292,N_7165);
nand U8459 (N_8459,N_7937,N_7146);
or U8460 (N_8460,N_7769,N_7221);
or U8461 (N_8461,N_7569,N_7910);
nor U8462 (N_8462,N_7891,N_7045);
nor U8463 (N_8463,N_7466,N_7339);
and U8464 (N_8464,N_7451,N_7713);
xnor U8465 (N_8465,N_7740,N_7252);
and U8466 (N_8466,N_7248,N_7038);
and U8467 (N_8467,N_7597,N_7417);
xnor U8468 (N_8468,N_7437,N_7843);
nand U8469 (N_8469,N_7254,N_7364);
nor U8470 (N_8470,N_7201,N_7899);
or U8471 (N_8471,N_7738,N_7271);
nor U8472 (N_8472,N_7090,N_7606);
xnor U8473 (N_8473,N_7407,N_7694);
nand U8474 (N_8474,N_7807,N_7382);
nand U8475 (N_8475,N_7119,N_7468);
or U8476 (N_8476,N_7611,N_7050);
nor U8477 (N_8477,N_7792,N_7379);
xor U8478 (N_8478,N_7245,N_7293);
nor U8479 (N_8479,N_7237,N_7344);
and U8480 (N_8480,N_7200,N_7246);
or U8481 (N_8481,N_7634,N_7046);
and U8482 (N_8482,N_7734,N_7223);
and U8483 (N_8483,N_7215,N_7778);
xor U8484 (N_8484,N_7207,N_7219);
nand U8485 (N_8485,N_7989,N_7490);
nand U8486 (N_8486,N_7895,N_7433);
xnor U8487 (N_8487,N_7832,N_7656);
and U8488 (N_8488,N_7241,N_7774);
xnor U8489 (N_8489,N_7347,N_7720);
nor U8490 (N_8490,N_7833,N_7211);
nand U8491 (N_8491,N_7655,N_7183);
or U8492 (N_8492,N_7131,N_7053);
nand U8493 (N_8493,N_7981,N_7771);
or U8494 (N_8494,N_7999,N_7374);
nor U8495 (N_8495,N_7318,N_7172);
nand U8496 (N_8496,N_7210,N_7585);
or U8497 (N_8497,N_7033,N_7023);
nand U8498 (N_8498,N_7996,N_7444);
nor U8499 (N_8499,N_7402,N_7894);
or U8500 (N_8500,N_7085,N_7800);
or U8501 (N_8501,N_7456,N_7159);
nand U8502 (N_8502,N_7077,N_7007);
and U8503 (N_8503,N_7308,N_7235);
xnor U8504 (N_8504,N_7615,N_7261);
xor U8505 (N_8505,N_7999,N_7893);
nor U8506 (N_8506,N_7131,N_7816);
nor U8507 (N_8507,N_7412,N_7380);
nor U8508 (N_8508,N_7622,N_7099);
and U8509 (N_8509,N_7450,N_7877);
xor U8510 (N_8510,N_7535,N_7413);
or U8511 (N_8511,N_7003,N_7807);
and U8512 (N_8512,N_7865,N_7349);
or U8513 (N_8513,N_7297,N_7548);
nand U8514 (N_8514,N_7901,N_7012);
and U8515 (N_8515,N_7751,N_7998);
nand U8516 (N_8516,N_7164,N_7894);
xnor U8517 (N_8517,N_7711,N_7078);
nand U8518 (N_8518,N_7671,N_7301);
and U8519 (N_8519,N_7343,N_7998);
nand U8520 (N_8520,N_7683,N_7649);
and U8521 (N_8521,N_7455,N_7963);
and U8522 (N_8522,N_7398,N_7409);
nor U8523 (N_8523,N_7709,N_7584);
nand U8524 (N_8524,N_7793,N_7902);
and U8525 (N_8525,N_7413,N_7858);
xor U8526 (N_8526,N_7880,N_7050);
or U8527 (N_8527,N_7459,N_7923);
or U8528 (N_8528,N_7631,N_7541);
nor U8529 (N_8529,N_7865,N_7193);
nand U8530 (N_8530,N_7201,N_7651);
and U8531 (N_8531,N_7978,N_7385);
and U8532 (N_8532,N_7301,N_7207);
nor U8533 (N_8533,N_7006,N_7276);
nor U8534 (N_8534,N_7302,N_7295);
or U8535 (N_8535,N_7749,N_7102);
and U8536 (N_8536,N_7023,N_7120);
xnor U8537 (N_8537,N_7522,N_7215);
nor U8538 (N_8538,N_7319,N_7245);
nand U8539 (N_8539,N_7757,N_7659);
nor U8540 (N_8540,N_7582,N_7683);
xnor U8541 (N_8541,N_7657,N_7414);
and U8542 (N_8542,N_7209,N_7934);
nand U8543 (N_8543,N_7087,N_7875);
and U8544 (N_8544,N_7967,N_7862);
nand U8545 (N_8545,N_7670,N_7563);
nor U8546 (N_8546,N_7210,N_7127);
and U8547 (N_8547,N_7301,N_7663);
nor U8548 (N_8548,N_7574,N_7557);
xnor U8549 (N_8549,N_7647,N_7534);
nor U8550 (N_8550,N_7405,N_7725);
and U8551 (N_8551,N_7747,N_7555);
or U8552 (N_8552,N_7037,N_7296);
xor U8553 (N_8553,N_7754,N_7544);
or U8554 (N_8554,N_7383,N_7600);
nor U8555 (N_8555,N_7656,N_7841);
nor U8556 (N_8556,N_7089,N_7790);
nor U8557 (N_8557,N_7741,N_7383);
nand U8558 (N_8558,N_7494,N_7608);
or U8559 (N_8559,N_7836,N_7408);
xor U8560 (N_8560,N_7086,N_7697);
and U8561 (N_8561,N_7085,N_7323);
or U8562 (N_8562,N_7805,N_7537);
and U8563 (N_8563,N_7196,N_7458);
xor U8564 (N_8564,N_7131,N_7448);
or U8565 (N_8565,N_7021,N_7989);
or U8566 (N_8566,N_7446,N_7947);
nand U8567 (N_8567,N_7903,N_7286);
or U8568 (N_8568,N_7803,N_7509);
xor U8569 (N_8569,N_7966,N_7004);
nand U8570 (N_8570,N_7803,N_7281);
nand U8571 (N_8571,N_7270,N_7211);
xnor U8572 (N_8572,N_7709,N_7019);
and U8573 (N_8573,N_7041,N_7441);
xor U8574 (N_8574,N_7181,N_7284);
and U8575 (N_8575,N_7482,N_7588);
nand U8576 (N_8576,N_7267,N_7156);
and U8577 (N_8577,N_7208,N_7627);
xnor U8578 (N_8578,N_7366,N_7933);
nand U8579 (N_8579,N_7920,N_7137);
xor U8580 (N_8580,N_7051,N_7589);
nand U8581 (N_8581,N_7094,N_7114);
nor U8582 (N_8582,N_7583,N_7710);
xnor U8583 (N_8583,N_7332,N_7989);
nand U8584 (N_8584,N_7627,N_7920);
nand U8585 (N_8585,N_7431,N_7410);
nor U8586 (N_8586,N_7921,N_7475);
nand U8587 (N_8587,N_7244,N_7834);
and U8588 (N_8588,N_7925,N_7556);
nor U8589 (N_8589,N_7572,N_7149);
nor U8590 (N_8590,N_7278,N_7886);
and U8591 (N_8591,N_7869,N_7609);
and U8592 (N_8592,N_7484,N_7461);
and U8593 (N_8593,N_7385,N_7559);
and U8594 (N_8594,N_7777,N_7249);
and U8595 (N_8595,N_7416,N_7660);
xnor U8596 (N_8596,N_7405,N_7958);
xnor U8597 (N_8597,N_7778,N_7021);
nor U8598 (N_8598,N_7041,N_7249);
or U8599 (N_8599,N_7469,N_7239);
xnor U8600 (N_8600,N_7645,N_7341);
or U8601 (N_8601,N_7449,N_7474);
and U8602 (N_8602,N_7843,N_7269);
and U8603 (N_8603,N_7879,N_7815);
xor U8604 (N_8604,N_7884,N_7183);
and U8605 (N_8605,N_7220,N_7115);
and U8606 (N_8606,N_7571,N_7065);
nor U8607 (N_8607,N_7195,N_7308);
nor U8608 (N_8608,N_7807,N_7445);
xnor U8609 (N_8609,N_7958,N_7079);
and U8610 (N_8610,N_7086,N_7477);
nand U8611 (N_8611,N_7252,N_7121);
xor U8612 (N_8612,N_7801,N_7884);
nor U8613 (N_8613,N_7176,N_7469);
and U8614 (N_8614,N_7070,N_7220);
nand U8615 (N_8615,N_7318,N_7699);
nand U8616 (N_8616,N_7651,N_7323);
and U8617 (N_8617,N_7396,N_7931);
xnor U8618 (N_8618,N_7012,N_7469);
nand U8619 (N_8619,N_7023,N_7965);
and U8620 (N_8620,N_7715,N_7637);
nor U8621 (N_8621,N_7603,N_7516);
and U8622 (N_8622,N_7197,N_7304);
or U8623 (N_8623,N_7763,N_7556);
nor U8624 (N_8624,N_7737,N_7978);
or U8625 (N_8625,N_7734,N_7930);
or U8626 (N_8626,N_7376,N_7205);
nor U8627 (N_8627,N_7894,N_7531);
or U8628 (N_8628,N_7265,N_7248);
nor U8629 (N_8629,N_7546,N_7748);
nor U8630 (N_8630,N_7582,N_7823);
xnor U8631 (N_8631,N_7710,N_7763);
nand U8632 (N_8632,N_7179,N_7207);
or U8633 (N_8633,N_7204,N_7980);
nand U8634 (N_8634,N_7772,N_7393);
xor U8635 (N_8635,N_7327,N_7292);
xnor U8636 (N_8636,N_7227,N_7575);
or U8637 (N_8637,N_7296,N_7554);
xor U8638 (N_8638,N_7822,N_7675);
xor U8639 (N_8639,N_7031,N_7431);
nand U8640 (N_8640,N_7928,N_7364);
or U8641 (N_8641,N_7610,N_7130);
and U8642 (N_8642,N_7343,N_7547);
nand U8643 (N_8643,N_7834,N_7786);
nand U8644 (N_8644,N_7786,N_7840);
xor U8645 (N_8645,N_7563,N_7937);
or U8646 (N_8646,N_7246,N_7285);
and U8647 (N_8647,N_7766,N_7101);
nor U8648 (N_8648,N_7076,N_7605);
xor U8649 (N_8649,N_7449,N_7126);
and U8650 (N_8650,N_7022,N_7793);
and U8651 (N_8651,N_7658,N_7902);
or U8652 (N_8652,N_7092,N_7491);
or U8653 (N_8653,N_7651,N_7816);
xnor U8654 (N_8654,N_7256,N_7124);
xor U8655 (N_8655,N_7538,N_7589);
nor U8656 (N_8656,N_7794,N_7953);
and U8657 (N_8657,N_7674,N_7199);
xor U8658 (N_8658,N_7401,N_7334);
or U8659 (N_8659,N_7927,N_7454);
nand U8660 (N_8660,N_7222,N_7608);
or U8661 (N_8661,N_7142,N_7709);
nand U8662 (N_8662,N_7028,N_7544);
xor U8663 (N_8663,N_7074,N_7446);
nand U8664 (N_8664,N_7932,N_7319);
nand U8665 (N_8665,N_7855,N_7115);
xnor U8666 (N_8666,N_7647,N_7238);
nor U8667 (N_8667,N_7277,N_7489);
nor U8668 (N_8668,N_7903,N_7083);
and U8669 (N_8669,N_7659,N_7073);
nor U8670 (N_8670,N_7199,N_7943);
nand U8671 (N_8671,N_7063,N_7402);
xnor U8672 (N_8672,N_7205,N_7519);
xor U8673 (N_8673,N_7751,N_7788);
or U8674 (N_8674,N_7477,N_7790);
and U8675 (N_8675,N_7628,N_7036);
or U8676 (N_8676,N_7334,N_7134);
or U8677 (N_8677,N_7155,N_7458);
or U8678 (N_8678,N_7859,N_7260);
or U8679 (N_8679,N_7016,N_7712);
xor U8680 (N_8680,N_7329,N_7581);
or U8681 (N_8681,N_7792,N_7538);
nand U8682 (N_8682,N_7873,N_7100);
xor U8683 (N_8683,N_7572,N_7137);
xnor U8684 (N_8684,N_7494,N_7225);
nor U8685 (N_8685,N_7219,N_7201);
nand U8686 (N_8686,N_7094,N_7271);
and U8687 (N_8687,N_7171,N_7609);
xor U8688 (N_8688,N_7982,N_7781);
nand U8689 (N_8689,N_7964,N_7159);
nand U8690 (N_8690,N_7992,N_7665);
nor U8691 (N_8691,N_7400,N_7518);
or U8692 (N_8692,N_7831,N_7489);
and U8693 (N_8693,N_7267,N_7853);
nand U8694 (N_8694,N_7724,N_7177);
or U8695 (N_8695,N_7060,N_7500);
or U8696 (N_8696,N_7279,N_7959);
nor U8697 (N_8697,N_7512,N_7412);
xor U8698 (N_8698,N_7975,N_7116);
and U8699 (N_8699,N_7210,N_7674);
and U8700 (N_8700,N_7994,N_7256);
and U8701 (N_8701,N_7026,N_7533);
and U8702 (N_8702,N_7671,N_7851);
xor U8703 (N_8703,N_7963,N_7112);
nor U8704 (N_8704,N_7626,N_7694);
nor U8705 (N_8705,N_7417,N_7150);
nor U8706 (N_8706,N_7403,N_7799);
nand U8707 (N_8707,N_7351,N_7880);
nand U8708 (N_8708,N_7229,N_7439);
or U8709 (N_8709,N_7474,N_7140);
nor U8710 (N_8710,N_7996,N_7285);
or U8711 (N_8711,N_7452,N_7204);
nand U8712 (N_8712,N_7131,N_7016);
and U8713 (N_8713,N_7146,N_7524);
xnor U8714 (N_8714,N_7849,N_7194);
or U8715 (N_8715,N_7635,N_7834);
and U8716 (N_8716,N_7443,N_7812);
nand U8717 (N_8717,N_7280,N_7822);
or U8718 (N_8718,N_7380,N_7585);
nor U8719 (N_8719,N_7415,N_7559);
xor U8720 (N_8720,N_7701,N_7778);
xor U8721 (N_8721,N_7896,N_7789);
and U8722 (N_8722,N_7333,N_7789);
nand U8723 (N_8723,N_7340,N_7729);
nand U8724 (N_8724,N_7112,N_7351);
and U8725 (N_8725,N_7829,N_7448);
or U8726 (N_8726,N_7149,N_7576);
or U8727 (N_8727,N_7134,N_7959);
nor U8728 (N_8728,N_7531,N_7847);
or U8729 (N_8729,N_7333,N_7558);
or U8730 (N_8730,N_7771,N_7046);
nand U8731 (N_8731,N_7759,N_7677);
nand U8732 (N_8732,N_7267,N_7384);
and U8733 (N_8733,N_7574,N_7400);
nand U8734 (N_8734,N_7585,N_7557);
nand U8735 (N_8735,N_7876,N_7450);
and U8736 (N_8736,N_7531,N_7473);
and U8737 (N_8737,N_7346,N_7898);
xnor U8738 (N_8738,N_7881,N_7957);
or U8739 (N_8739,N_7562,N_7625);
xor U8740 (N_8740,N_7762,N_7656);
nand U8741 (N_8741,N_7759,N_7888);
and U8742 (N_8742,N_7789,N_7373);
xor U8743 (N_8743,N_7221,N_7308);
and U8744 (N_8744,N_7202,N_7231);
xor U8745 (N_8745,N_7288,N_7974);
and U8746 (N_8746,N_7478,N_7880);
nor U8747 (N_8747,N_7694,N_7365);
nor U8748 (N_8748,N_7912,N_7278);
or U8749 (N_8749,N_7202,N_7282);
or U8750 (N_8750,N_7915,N_7369);
or U8751 (N_8751,N_7665,N_7596);
xnor U8752 (N_8752,N_7498,N_7391);
or U8753 (N_8753,N_7825,N_7788);
xnor U8754 (N_8754,N_7289,N_7111);
nand U8755 (N_8755,N_7552,N_7136);
nor U8756 (N_8756,N_7589,N_7699);
nor U8757 (N_8757,N_7715,N_7270);
nor U8758 (N_8758,N_7640,N_7657);
nor U8759 (N_8759,N_7412,N_7402);
nor U8760 (N_8760,N_7025,N_7620);
and U8761 (N_8761,N_7887,N_7261);
xor U8762 (N_8762,N_7201,N_7392);
nor U8763 (N_8763,N_7115,N_7723);
nor U8764 (N_8764,N_7485,N_7279);
or U8765 (N_8765,N_7619,N_7606);
xnor U8766 (N_8766,N_7823,N_7192);
and U8767 (N_8767,N_7774,N_7175);
or U8768 (N_8768,N_7966,N_7015);
or U8769 (N_8769,N_7373,N_7452);
xnor U8770 (N_8770,N_7265,N_7934);
or U8771 (N_8771,N_7037,N_7478);
and U8772 (N_8772,N_7772,N_7218);
nor U8773 (N_8773,N_7944,N_7992);
nor U8774 (N_8774,N_7001,N_7951);
or U8775 (N_8775,N_7151,N_7390);
or U8776 (N_8776,N_7705,N_7107);
and U8777 (N_8777,N_7141,N_7004);
nor U8778 (N_8778,N_7573,N_7802);
xor U8779 (N_8779,N_7266,N_7927);
or U8780 (N_8780,N_7337,N_7929);
and U8781 (N_8781,N_7972,N_7529);
nor U8782 (N_8782,N_7070,N_7293);
and U8783 (N_8783,N_7030,N_7202);
xnor U8784 (N_8784,N_7428,N_7854);
and U8785 (N_8785,N_7084,N_7326);
and U8786 (N_8786,N_7945,N_7979);
and U8787 (N_8787,N_7004,N_7591);
nor U8788 (N_8788,N_7799,N_7842);
xor U8789 (N_8789,N_7842,N_7455);
xor U8790 (N_8790,N_7527,N_7319);
nor U8791 (N_8791,N_7422,N_7243);
nand U8792 (N_8792,N_7970,N_7480);
nand U8793 (N_8793,N_7179,N_7931);
nand U8794 (N_8794,N_7626,N_7770);
and U8795 (N_8795,N_7508,N_7208);
or U8796 (N_8796,N_7354,N_7439);
nor U8797 (N_8797,N_7825,N_7633);
nor U8798 (N_8798,N_7989,N_7739);
nand U8799 (N_8799,N_7650,N_7608);
and U8800 (N_8800,N_7654,N_7382);
and U8801 (N_8801,N_7420,N_7013);
nor U8802 (N_8802,N_7915,N_7816);
nand U8803 (N_8803,N_7447,N_7642);
nor U8804 (N_8804,N_7470,N_7801);
xnor U8805 (N_8805,N_7817,N_7367);
or U8806 (N_8806,N_7930,N_7413);
xnor U8807 (N_8807,N_7830,N_7884);
and U8808 (N_8808,N_7236,N_7054);
nor U8809 (N_8809,N_7729,N_7372);
and U8810 (N_8810,N_7587,N_7452);
xnor U8811 (N_8811,N_7292,N_7529);
xor U8812 (N_8812,N_7623,N_7134);
nand U8813 (N_8813,N_7558,N_7745);
nand U8814 (N_8814,N_7337,N_7663);
nand U8815 (N_8815,N_7936,N_7625);
and U8816 (N_8816,N_7685,N_7411);
or U8817 (N_8817,N_7784,N_7060);
or U8818 (N_8818,N_7099,N_7977);
nor U8819 (N_8819,N_7283,N_7479);
nor U8820 (N_8820,N_7538,N_7822);
xor U8821 (N_8821,N_7095,N_7306);
or U8822 (N_8822,N_7174,N_7426);
and U8823 (N_8823,N_7966,N_7705);
nand U8824 (N_8824,N_7988,N_7210);
nand U8825 (N_8825,N_7624,N_7529);
nand U8826 (N_8826,N_7956,N_7011);
xor U8827 (N_8827,N_7772,N_7080);
nor U8828 (N_8828,N_7085,N_7488);
nand U8829 (N_8829,N_7248,N_7494);
xnor U8830 (N_8830,N_7206,N_7353);
or U8831 (N_8831,N_7199,N_7559);
xnor U8832 (N_8832,N_7181,N_7831);
nand U8833 (N_8833,N_7829,N_7589);
nor U8834 (N_8834,N_7445,N_7394);
and U8835 (N_8835,N_7396,N_7470);
xnor U8836 (N_8836,N_7735,N_7566);
or U8837 (N_8837,N_7545,N_7450);
xor U8838 (N_8838,N_7559,N_7804);
or U8839 (N_8839,N_7606,N_7754);
and U8840 (N_8840,N_7428,N_7559);
xnor U8841 (N_8841,N_7030,N_7518);
xor U8842 (N_8842,N_7484,N_7370);
nand U8843 (N_8843,N_7554,N_7960);
nand U8844 (N_8844,N_7373,N_7757);
and U8845 (N_8845,N_7683,N_7131);
nor U8846 (N_8846,N_7556,N_7699);
xor U8847 (N_8847,N_7633,N_7408);
or U8848 (N_8848,N_7802,N_7240);
or U8849 (N_8849,N_7426,N_7894);
nand U8850 (N_8850,N_7696,N_7851);
or U8851 (N_8851,N_7635,N_7273);
xnor U8852 (N_8852,N_7914,N_7042);
nor U8853 (N_8853,N_7306,N_7385);
or U8854 (N_8854,N_7885,N_7272);
or U8855 (N_8855,N_7104,N_7481);
or U8856 (N_8856,N_7252,N_7426);
xor U8857 (N_8857,N_7080,N_7679);
nor U8858 (N_8858,N_7644,N_7126);
nor U8859 (N_8859,N_7542,N_7516);
nand U8860 (N_8860,N_7769,N_7731);
or U8861 (N_8861,N_7482,N_7341);
xor U8862 (N_8862,N_7203,N_7088);
nand U8863 (N_8863,N_7940,N_7315);
or U8864 (N_8864,N_7724,N_7637);
or U8865 (N_8865,N_7207,N_7791);
xnor U8866 (N_8866,N_7663,N_7718);
xnor U8867 (N_8867,N_7594,N_7500);
and U8868 (N_8868,N_7575,N_7182);
xor U8869 (N_8869,N_7301,N_7874);
nand U8870 (N_8870,N_7215,N_7371);
xor U8871 (N_8871,N_7225,N_7806);
xnor U8872 (N_8872,N_7776,N_7930);
nand U8873 (N_8873,N_7126,N_7687);
nor U8874 (N_8874,N_7667,N_7609);
xnor U8875 (N_8875,N_7588,N_7010);
or U8876 (N_8876,N_7014,N_7028);
nor U8877 (N_8877,N_7125,N_7171);
and U8878 (N_8878,N_7366,N_7217);
and U8879 (N_8879,N_7944,N_7833);
and U8880 (N_8880,N_7982,N_7360);
nand U8881 (N_8881,N_7563,N_7130);
nand U8882 (N_8882,N_7300,N_7335);
nor U8883 (N_8883,N_7385,N_7345);
and U8884 (N_8884,N_7748,N_7674);
xor U8885 (N_8885,N_7041,N_7647);
nor U8886 (N_8886,N_7531,N_7362);
nor U8887 (N_8887,N_7557,N_7048);
or U8888 (N_8888,N_7732,N_7464);
and U8889 (N_8889,N_7250,N_7760);
and U8890 (N_8890,N_7563,N_7788);
xnor U8891 (N_8891,N_7447,N_7166);
or U8892 (N_8892,N_7599,N_7532);
and U8893 (N_8893,N_7999,N_7968);
or U8894 (N_8894,N_7487,N_7223);
nand U8895 (N_8895,N_7549,N_7880);
or U8896 (N_8896,N_7456,N_7042);
nand U8897 (N_8897,N_7658,N_7482);
nand U8898 (N_8898,N_7618,N_7581);
or U8899 (N_8899,N_7313,N_7924);
nor U8900 (N_8900,N_7449,N_7189);
xor U8901 (N_8901,N_7672,N_7228);
nand U8902 (N_8902,N_7114,N_7201);
xor U8903 (N_8903,N_7952,N_7557);
and U8904 (N_8904,N_7816,N_7183);
xor U8905 (N_8905,N_7504,N_7641);
nor U8906 (N_8906,N_7333,N_7733);
nand U8907 (N_8907,N_7832,N_7354);
xor U8908 (N_8908,N_7843,N_7543);
or U8909 (N_8909,N_7309,N_7767);
nand U8910 (N_8910,N_7609,N_7088);
nand U8911 (N_8911,N_7132,N_7250);
nand U8912 (N_8912,N_7714,N_7144);
xnor U8913 (N_8913,N_7596,N_7018);
nand U8914 (N_8914,N_7510,N_7123);
xor U8915 (N_8915,N_7522,N_7939);
nand U8916 (N_8916,N_7807,N_7684);
nor U8917 (N_8917,N_7007,N_7301);
xnor U8918 (N_8918,N_7458,N_7861);
nand U8919 (N_8919,N_7041,N_7309);
nand U8920 (N_8920,N_7921,N_7838);
nand U8921 (N_8921,N_7188,N_7217);
and U8922 (N_8922,N_7098,N_7232);
xnor U8923 (N_8923,N_7736,N_7264);
xnor U8924 (N_8924,N_7933,N_7658);
nand U8925 (N_8925,N_7956,N_7310);
xnor U8926 (N_8926,N_7392,N_7210);
nand U8927 (N_8927,N_7738,N_7668);
xor U8928 (N_8928,N_7260,N_7517);
nor U8929 (N_8929,N_7693,N_7524);
nand U8930 (N_8930,N_7648,N_7966);
or U8931 (N_8931,N_7093,N_7345);
nand U8932 (N_8932,N_7653,N_7989);
xnor U8933 (N_8933,N_7289,N_7753);
nand U8934 (N_8934,N_7355,N_7971);
and U8935 (N_8935,N_7742,N_7256);
nor U8936 (N_8936,N_7997,N_7705);
xnor U8937 (N_8937,N_7851,N_7112);
nor U8938 (N_8938,N_7348,N_7236);
nor U8939 (N_8939,N_7410,N_7784);
nand U8940 (N_8940,N_7385,N_7051);
xnor U8941 (N_8941,N_7645,N_7946);
or U8942 (N_8942,N_7891,N_7271);
nor U8943 (N_8943,N_7364,N_7776);
nand U8944 (N_8944,N_7672,N_7660);
or U8945 (N_8945,N_7500,N_7702);
nand U8946 (N_8946,N_7105,N_7801);
and U8947 (N_8947,N_7924,N_7292);
nor U8948 (N_8948,N_7216,N_7226);
and U8949 (N_8949,N_7304,N_7140);
or U8950 (N_8950,N_7188,N_7344);
nand U8951 (N_8951,N_7933,N_7123);
xnor U8952 (N_8952,N_7694,N_7309);
and U8953 (N_8953,N_7371,N_7889);
xnor U8954 (N_8954,N_7919,N_7443);
nand U8955 (N_8955,N_7796,N_7261);
nor U8956 (N_8956,N_7708,N_7124);
nand U8957 (N_8957,N_7090,N_7452);
and U8958 (N_8958,N_7963,N_7892);
nor U8959 (N_8959,N_7706,N_7490);
nor U8960 (N_8960,N_7185,N_7115);
xnor U8961 (N_8961,N_7205,N_7799);
nand U8962 (N_8962,N_7192,N_7024);
xnor U8963 (N_8963,N_7115,N_7836);
nand U8964 (N_8964,N_7037,N_7621);
and U8965 (N_8965,N_7887,N_7161);
nor U8966 (N_8966,N_7777,N_7166);
or U8967 (N_8967,N_7436,N_7295);
nand U8968 (N_8968,N_7422,N_7102);
xor U8969 (N_8969,N_7510,N_7747);
and U8970 (N_8970,N_7583,N_7613);
nor U8971 (N_8971,N_7594,N_7866);
xor U8972 (N_8972,N_7599,N_7477);
nand U8973 (N_8973,N_7629,N_7752);
nor U8974 (N_8974,N_7238,N_7677);
and U8975 (N_8975,N_7069,N_7914);
or U8976 (N_8976,N_7923,N_7773);
nor U8977 (N_8977,N_7663,N_7680);
and U8978 (N_8978,N_7317,N_7959);
nor U8979 (N_8979,N_7724,N_7007);
nand U8980 (N_8980,N_7879,N_7436);
or U8981 (N_8981,N_7641,N_7782);
xnor U8982 (N_8982,N_7170,N_7456);
nor U8983 (N_8983,N_7116,N_7221);
nand U8984 (N_8984,N_7656,N_7797);
nand U8985 (N_8985,N_7967,N_7729);
xnor U8986 (N_8986,N_7326,N_7615);
nor U8987 (N_8987,N_7358,N_7934);
and U8988 (N_8988,N_7731,N_7734);
or U8989 (N_8989,N_7086,N_7300);
or U8990 (N_8990,N_7023,N_7937);
nor U8991 (N_8991,N_7213,N_7329);
or U8992 (N_8992,N_7295,N_7490);
xnor U8993 (N_8993,N_7506,N_7409);
and U8994 (N_8994,N_7422,N_7674);
and U8995 (N_8995,N_7630,N_7213);
xnor U8996 (N_8996,N_7630,N_7095);
nor U8997 (N_8997,N_7187,N_7548);
or U8998 (N_8998,N_7528,N_7559);
and U8999 (N_8999,N_7984,N_7997);
xnor U9000 (N_9000,N_8133,N_8480);
nand U9001 (N_9001,N_8045,N_8606);
nor U9002 (N_9002,N_8981,N_8583);
and U9003 (N_9003,N_8800,N_8705);
and U9004 (N_9004,N_8811,N_8877);
xnor U9005 (N_9005,N_8665,N_8476);
and U9006 (N_9006,N_8332,N_8706);
nor U9007 (N_9007,N_8451,N_8502);
nand U9008 (N_9008,N_8531,N_8396);
and U9009 (N_9009,N_8536,N_8679);
xor U9010 (N_9010,N_8419,N_8026);
nor U9011 (N_9011,N_8720,N_8612);
nand U9012 (N_9012,N_8319,N_8103);
and U9013 (N_9013,N_8915,N_8182);
nor U9014 (N_9014,N_8237,N_8604);
nor U9015 (N_9015,N_8382,N_8986);
and U9016 (N_9016,N_8433,N_8163);
and U9017 (N_9017,N_8173,N_8972);
xor U9018 (N_9018,N_8749,N_8539);
or U9019 (N_9019,N_8183,N_8513);
xor U9020 (N_9020,N_8700,N_8895);
and U9021 (N_9021,N_8509,N_8709);
xnor U9022 (N_9022,N_8731,N_8358);
nand U9023 (N_9023,N_8534,N_8410);
or U9024 (N_9024,N_8269,N_8184);
or U9025 (N_9025,N_8590,N_8758);
or U9026 (N_9026,N_8384,N_8324);
or U9027 (N_9027,N_8096,N_8175);
and U9028 (N_9028,N_8345,N_8444);
or U9029 (N_9029,N_8858,N_8381);
or U9030 (N_9030,N_8992,N_8389);
nor U9031 (N_9031,N_8646,N_8864);
and U9032 (N_9032,N_8478,N_8687);
xor U9033 (N_9033,N_8769,N_8870);
nand U9034 (N_9034,N_8714,N_8938);
or U9035 (N_9035,N_8690,N_8941);
nor U9036 (N_9036,N_8072,N_8862);
or U9037 (N_9037,N_8686,N_8420);
or U9038 (N_9038,N_8934,N_8998);
nand U9039 (N_9039,N_8655,N_8960);
and U9040 (N_9040,N_8848,N_8892);
xnor U9041 (N_9041,N_8178,N_8947);
and U9042 (N_9042,N_8458,N_8727);
nor U9043 (N_9043,N_8076,N_8568);
and U9044 (N_9044,N_8985,N_8212);
and U9045 (N_9045,N_8219,N_8192);
or U9046 (N_9046,N_8233,N_8157);
and U9047 (N_9047,N_8819,N_8553);
or U9048 (N_9048,N_8701,N_8397);
or U9049 (N_9049,N_8284,N_8028);
and U9050 (N_9050,N_8274,N_8452);
or U9051 (N_9051,N_8311,N_8744);
nand U9052 (N_9052,N_8684,N_8979);
and U9053 (N_9053,N_8473,N_8555);
nand U9054 (N_9054,N_8429,N_8414);
xnor U9055 (N_9055,N_8369,N_8780);
and U9056 (N_9056,N_8794,N_8147);
or U9057 (N_9057,N_8334,N_8627);
nand U9058 (N_9058,N_8678,N_8089);
or U9059 (N_9059,N_8065,N_8398);
xor U9060 (N_9060,N_8196,N_8785);
nand U9061 (N_9061,N_8543,N_8786);
nand U9062 (N_9062,N_8748,N_8626);
and U9063 (N_9063,N_8850,N_8151);
and U9064 (N_9064,N_8106,N_8812);
nor U9065 (N_9065,N_8847,N_8077);
xor U9066 (N_9066,N_8620,N_8120);
xnor U9067 (N_9067,N_8214,N_8246);
xor U9068 (N_9068,N_8408,N_8060);
nand U9069 (N_9069,N_8017,N_8660);
and U9070 (N_9070,N_8517,N_8712);
and U9071 (N_9071,N_8697,N_8841);
xnor U9072 (N_9072,N_8359,N_8362);
xnor U9073 (N_9073,N_8418,N_8708);
nor U9074 (N_9074,N_8238,N_8263);
xnor U9075 (N_9075,N_8716,N_8383);
nor U9076 (N_9076,N_8771,N_8088);
and U9077 (N_9077,N_8518,N_8411);
xnor U9078 (N_9078,N_8625,N_8501);
and U9079 (N_9079,N_8961,N_8789);
nor U9080 (N_9080,N_8462,N_8011);
nor U9081 (N_9081,N_8868,N_8307);
nor U9082 (N_9082,N_8589,N_8181);
and U9083 (N_9083,N_8019,N_8622);
or U9084 (N_9084,N_8931,N_8240);
and U9085 (N_9085,N_8942,N_8461);
or U9086 (N_9086,N_8888,N_8587);
nand U9087 (N_9087,N_8000,N_8857);
xor U9088 (N_9088,N_8043,N_8025);
nor U9089 (N_9089,N_8217,N_8730);
nand U9090 (N_9090,N_8865,N_8576);
or U9091 (N_9091,N_8609,N_8556);
nor U9092 (N_9092,N_8245,N_8668);
nand U9093 (N_9093,N_8260,N_8601);
nor U9094 (N_9094,N_8965,N_8884);
nand U9095 (N_9095,N_8453,N_8953);
xnor U9096 (N_9096,N_8613,N_8838);
nand U9097 (N_9097,N_8897,N_8547);
and U9098 (N_9098,N_8628,N_8399);
nand U9099 (N_9099,N_8649,N_8887);
nor U9100 (N_9100,N_8236,N_8891);
nand U9101 (N_9101,N_8228,N_8216);
nor U9102 (N_9102,N_8797,N_8680);
and U9103 (N_9103,N_8067,N_8034);
xnor U9104 (N_9104,N_8044,N_8978);
nand U9105 (N_9105,N_8929,N_8764);
nand U9106 (N_9106,N_8801,N_8405);
or U9107 (N_9107,N_8357,N_8940);
or U9108 (N_9108,N_8943,N_8899);
nand U9109 (N_9109,N_8252,N_8928);
and U9110 (N_9110,N_8251,N_8851);
nor U9111 (N_9111,N_8958,N_8293);
or U9112 (N_9112,N_8933,N_8097);
nor U9113 (N_9113,N_8361,N_8138);
nor U9114 (N_9114,N_8050,N_8202);
nand U9115 (N_9115,N_8492,N_8346);
and U9116 (N_9116,N_8991,N_8787);
and U9117 (N_9117,N_8520,N_8290);
or U9118 (N_9118,N_8835,N_8894);
or U9119 (N_9119,N_8790,N_8530);
or U9120 (N_9120,N_8842,N_8339);
and U9121 (N_9121,N_8258,N_8071);
or U9122 (N_9122,N_8316,N_8285);
nor U9123 (N_9123,N_8693,N_8839);
and U9124 (N_9124,N_8921,N_8306);
nor U9125 (N_9125,N_8742,N_8936);
and U9126 (N_9126,N_8149,N_8909);
xor U9127 (N_9127,N_8195,N_8598);
xor U9128 (N_9128,N_8828,N_8308);
nand U9129 (N_9129,N_8635,N_8463);
nor U9130 (N_9130,N_8738,N_8289);
and U9131 (N_9131,N_8296,N_8494);
xor U9132 (N_9132,N_8910,N_8107);
nand U9133 (N_9133,N_8564,N_8248);
nand U9134 (N_9134,N_8728,N_8683);
or U9135 (N_9135,N_8090,N_8600);
xnor U9136 (N_9136,N_8641,N_8846);
or U9137 (N_9137,N_8618,N_8695);
xor U9138 (N_9138,N_8187,N_8803);
nor U9139 (N_9139,N_8393,N_8437);
and U9140 (N_9140,N_8087,N_8578);
or U9141 (N_9141,N_8834,N_8804);
xor U9142 (N_9142,N_8012,N_8400);
and U9143 (N_9143,N_8596,N_8924);
xor U9144 (N_9144,N_8733,N_8566);
or U9145 (N_9145,N_8669,N_8014);
and U9146 (N_9146,N_8310,N_8752);
or U9147 (N_9147,N_8432,N_8439);
nand U9148 (N_9148,N_8468,N_8372);
nand U9149 (N_9149,N_8853,N_8854);
nand U9150 (N_9150,N_8337,N_8951);
nand U9151 (N_9151,N_8599,N_8482);
or U9152 (N_9152,N_8220,N_8507);
xor U9153 (N_9153,N_8917,N_8715);
xnor U9154 (N_9154,N_8230,N_8360);
xor U9155 (N_9155,N_8079,N_8760);
nor U9156 (N_9156,N_8591,N_8484);
nand U9157 (N_9157,N_8352,N_8755);
xor U9158 (N_9158,N_8373,N_8557);
nand U9159 (N_9159,N_8863,N_8488);
xnor U9160 (N_9160,N_8465,N_8585);
nor U9161 (N_9161,N_8412,N_8820);
or U9162 (N_9162,N_8867,N_8882);
nor U9163 (N_9163,N_8002,N_8351);
and U9164 (N_9164,N_8843,N_8648);
and U9165 (N_9165,N_8559,N_8350);
or U9166 (N_9166,N_8191,N_8676);
and U9167 (N_9167,N_8213,N_8464);
nand U9168 (N_9168,N_8605,N_8487);
nor U9169 (N_9169,N_8747,N_8869);
nor U9170 (N_9170,N_8996,N_8529);
and U9171 (N_9171,N_8784,N_8443);
nor U9172 (N_9172,N_8018,N_8336);
or U9173 (N_9173,N_8554,N_8662);
nor U9174 (N_9174,N_8793,N_8344);
xor U9175 (N_9175,N_8190,N_8579);
nand U9176 (N_9176,N_8836,N_8431);
nand U9177 (N_9177,N_8390,N_8833);
or U9178 (N_9178,N_8244,N_8082);
xor U9179 (N_9179,N_8225,N_8922);
xnor U9180 (N_9180,N_8713,N_8912);
or U9181 (N_9181,N_8914,N_8881);
and U9182 (N_9182,N_8644,N_8435);
or U9183 (N_9183,N_8394,N_8615);
nand U9184 (N_9184,N_8282,N_8723);
nor U9185 (N_9185,N_8541,N_8407);
nand U9186 (N_9186,N_8112,N_8234);
and U9187 (N_9187,N_8905,N_8313);
nand U9188 (N_9188,N_8856,N_8058);
nor U9189 (N_9189,N_8831,N_8124);
nor U9190 (N_9190,N_8540,N_8736);
or U9191 (N_9191,N_8292,N_8342);
nor U9192 (N_9192,N_8078,N_8973);
xor U9193 (N_9193,N_8253,N_8855);
xnor U9194 (N_9194,N_8607,N_8526);
nor U9195 (N_9195,N_8340,N_8218);
and U9196 (N_9196,N_8732,N_8490);
xor U9197 (N_9197,N_8229,N_8276);
or U9198 (N_9198,N_8907,N_8059);
nor U9199 (N_9199,N_8805,N_8094);
xor U9200 (N_9200,N_8073,N_8015);
nor U9201 (N_9201,N_8001,N_8164);
nand U9202 (N_9202,N_8904,N_8677);
and U9203 (N_9203,N_8481,N_8279);
nand U9204 (N_9204,N_8469,N_8242);
nor U9205 (N_9205,N_8348,N_8172);
and U9206 (N_9206,N_8634,N_8257);
or U9207 (N_9207,N_8778,N_8883);
xor U9208 (N_9208,N_8954,N_8535);
nand U9209 (N_9209,N_8122,N_8699);
xor U9210 (N_9210,N_8170,N_8798);
nand U9211 (N_9211,N_8528,N_8673);
nor U9212 (N_9212,N_8523,N_8637);
xor U9213 (N_9213,N_8425,N_8250);
nand U9214 (N_9214,N_8654,N_8406);
and U9215 (N_9215,N_8074,N_8491);
nor U9216 (N_9216,N_8594,N_8134);
and U9217 (N_9217,N_8117,N_8208);
xor U9218 (N_9218,N_8524,N_8466);
nand U9219 (N_9219,N_8142,N_8624);
xor U9220 (N_9220,N_8066,N_8971);
or U9221 (N_9221,N_8436,N_8670);
xor U9222 (N_9222,N_8572,N_8156);
nand U9223 (N_9223,N_8499,N_8664);
and U9224 (N_9224,N_8982,N_8199);
nand U9225 (N_9225,N_8514,N_8809);
nand U9226 (N_9226,N_8141,N_8321);
or U9227 (N_9227,N_8674,N_8860);
and U9228 (N_9228,N_8113,N_8763);
or U9229 (N_9229,N_8631,N_8546);
nand U9230 (N_9230,N_8084,N_8969);
nand U9231 (N_9231,N_8180,N_8168);
or U9232 (N_9232,N_8303,N_8022);
and U9233 (N_9233,N_8003,N_8560);
nand U9234 (N_9234,N_8256,N_8186);
nor U9235 (N_9235,N_8685,N_8203);
xnor U9236 (N_9236,N_8108,N_8054);
and U9237 (N_9237,N_8404,N_8696);
or U9238 (N_9238,N_8448,N_8967);
or U9239 (N_9239,N_8966,N_8949);
nor U9240 (N_9240,N_8923,N_8368);
and U9241 (N_9241,N_8266,N_8725);
xor U9242 (N_9242,N_8243,N_8745);
nor U9243 (N_9243,N_8807,N_8051);
nor U9244 (N_9244,N_8642,N_8302);
and U9245 (N_9245,N_8057,N_8055);
or U9246 (N_9246,N_8756,N_8287);
and U9247 (N_9247,N_8675,N_8667);
nand U9248 (N_9248,N_8379,N_8896);
and U9249 (N_9249,N_8765,N_8314);
and U9250 (N_9250,N_8185,N_8355);
and U9251 (N_9251,N_8750,N_8416);
xnor U9252 (N_9252,N_8166,N_8584);
nor U9253 (N_9253,N_8827,N_8385);
or U9254 (N_9254,N_8273,N_8574);
nand U9255 (N_9255,N_8875,N_8254);
xor U9256 (N_9256,N_8861,N_8879);
nand U9257 (N_9257,N_8092,N_8571);
nor U9258 (N_9258,N_8544,N_8401);
xor U9259 (N_9259,N_8061,N_8046);
nand U9260 (N_9260,N_8768,N_8030);
nand U9261 (N_9261,N_8048,N_8698);
nand U9262 (N_9262,N_8146,N_8040);
nor U9263 (N_9263,N_8866,N_8131);
and U9264 (N_9264,N_8945,N_8197);
nor U9265 (N_9265,N_8630,N_8563);
and U9266 (N_9266,N_8957,N_8995);
nor U9267 (N_9267,N_8927,N_8160);
or U9268 (N_9268,N_8610,N_8322);
nand U9269 (N_9269,N_8286,N_8455);
nand U9270 (N_9270,N_8633,N_8671);
xor U9271 (N_9271,N_8512,N_8063);
xnor U9272 (N_9272,N_8315,N_8415);
nand U9273 (N_9273,N_8154,N_8999);
and U9274 (N_9274,N_8496,N_8140);
nor U9275 (N_9275,N_8013,N_8659);
nor U9276 (N_9276,N_8817,N_8643);
nor U9277 (N_9277,N_8886,N_8329);
and U9278 (N_9278,N_8719,N_8277);
or U9279 (N_9279,N_8532,N_8037);
and U9280 (N_9280,N_8300,N_8586);
xor U9281 (N_9281,N_8323,N_8459);
or U9282 (N_9282,N_8136,N_8349);
xnor U9283 (N_9283,N_8268,N_8911);
xnor U9284 (N_9284,N_8333,N_8221);
nor U9285 (N_9285,N_8483,N_8295);
and U9286 (N_9286,N_8118,N_8153);
nand U9287 (N_9287,N_8479,N_8663);
nor U9288 (N_9288,N_8597,N_8849);
xor U9289 (N_9289,N_8740,N_8005);
nor U9290 (N_9290,N_8110,N_8485);
or U9291 (N_9291,N_8388,N_8987);
xnor U9292 (N_9292,N_8903,N_8171);
xnor U9293 (N_9293,N_8188,N_8109);
and U9294 (N_9294,N_8522,N_8165);
or U9295 (N_9295,N_8537,N_8511);
or U9296 (N_9296,N_8751,N_8467);
or U9297 (N_9297,N_8457,N_8162);
nor U9298 (N_9298,N_8666,N_8611);
or U9299 (N_9299,N_8975,N_8796);
nor U9300 (N_9300,N_8049,N_8021);
nor U9301 (N_9301,N_8504,N_8772);
nor U9302 (N_9302,N_8033,N_8006);
nand U9303 (N_9303,N_8901,N_8261);
nor U9304 (N_9304,N_8977,N_8215);
nand U9305 (N_9305,N_8746,N_8737);
xnor U9306 (N_9306,N_8224,N_8493);
and U9307 (N_9307,N_8262,N_8691);
and U9308 (N_9308,N_8791,N_8515);
and U9309 (N_9309,N_8460,N_8100);
and U9310 (N_9310,N_8569,N_8211);
nor U9311 (N_9311,N_8232,N_8356);
nor U9312 (N_9312,N_8375,N_8688);
nand U9313 (N_9313,N_8830,N_8438);
or U9314 (N_9314,N_8328,N_8580);
and U9315 (N_9315,N_8792,N_8226);
nor U9316 (N_9316,N_8064,N_8454);
nor U9317 (N_9317,N_8291,N_8148);
and U9318 (N_9318,N_8024,N_8711);
or U9319 (N_9319,N_8083,N_8976);
and U9320 (N_9320,N_8813,N_8689);
xnor U9321 (N_9321,N_8085,N_8395);
nand U9322 (N_9322,N_8761,N_8354);
or U9323 (N_9323,N_8086,N_8821);
nand U9324 (N_9324,N_8994,N_8421);
or U9325 (N_9325,N_8091,N_8826);
or U9326 (N_9326,N_8980,N_8471);
or U9327 (N_9327,N_8781,N_8150);
nor U9328 (N_9328,N_8353,N_8900);
xnor U9329 (N_9329,N_8814,N_8053);
xor U9330 (N_9330,N_8710,N_8298);
or U9331 (N_9331,N_8505,N_8010);
or U9332 (N_9332,N_8155,N_8770);
nor U9333 (N_9333,N_8029,N_8130);
and U9334 (N_9334,N_8145,N_8486);
nor U9335 (N_9335,N_8309,N_8326);
nor U9336 (N_9336,N_8962,N_8939);
and U9337 (N_9337,N_8636,N_8516);
nor U9338 (N_9338,N_8222,N_8623);
or U9339 (N_9339,N_8702,N_8423);
xnor U9340 (N_9340,N_8325,N_8020);
and U9341 (N_9341,N_8189,N_8510);
or U9342 (N_9342,N_8080,N_8859);
nor U9343 (N_9343,N_8128,N_8272);
xnor U9344 (N_9344,N_8602,N_8341);
nand U9345 (N_9345,N_8717,N_8653);
nand U9346 (N_9346,N_8152,N_8824);
or U9347 (N_9347,N_8417,N_8852);
and U9348 (N_9348,N_8950,N_8776);
nand U9349 (N_9349,N_8402,N_8317);
and U9350 (N_9350,N_8593,N_8194);
and U9351 (N_9351,N_8176,N_8038);
nor U9352 (N_9352,N_8878,N_8426);
or U9353 (N_9353,N_8721,N_8158);
xor U9354 (N_9354,N_8829,N_8205);
xnor U9355 (N_9355,N_8521,N_8925);
nor U9356 (N_9356,N_8027,N_8906);
or U9357 (N_9357,N_8449,N_8582);
nor U9358 (N_9358,N_8632,N_8565);
nand U9359 (N_9359,N_8231,N_8657);
nor U9360 (N_9360,N_8802,N_8647);
or U9361 (N_9361,N_8808,N_8200);
and U9362 (N_9362,N_8409,N_8739);
xor U9363 (N_9363,N_8239,N_8447);
or U9364 (N_9364,N_8392,N_8004);
nor U9365 (N_9365,N_8111,N_8095);
or U9366 (N_9366,N_8549,N_8235);
and U9367 (N_9367,N_8595,N_8068);
nand U9368 (N_9368,N_8391,N_8270);
or U9369 (N_9369,N_8729,N_8380);
xor U9370 (N_9370,N_8081,N_8757);
xor U9371 (N_9371,N_8041,N_8508);
nor U9372 (N_9372,N_8387,N_8312);
xnor U9373 (N_9373,N_8127,N_8070);
nor U9374 (N_9374,N_8161,N_8031);
xnor U9375 (N_9375,N_8795,N_8363);
nand U9376 (N_9376,N_8959,N_8890);
xor U9377 (N_9377,N_8264,N_8989);
nor U9378 (N_9378,N_8335,N_8265);
and U9379 (N_9379,N_8777,N_8301);
nand U9380 (N_9380,N_8343,N_8658);
xor U9381 (N_9381,N_8428,N_8042);
nand U9382 (N_9382,N_8629,N_8874);
nor U9383 (N_9383,N_8588,N_8902);
nand U9384 (N_9384,N_8434,N_8413);
xor U9385 (N_9385,N_8008,N_8937);
or U9386 (N_9386,N_8993,N_8970);
and U9387 (N_9387,N_8114,N_8788);
nor U9388 (N_9388,N_8825,N_8159);
or U9389 (N_9389,N_8016,N_8919);
or U9390 (N_9390,N_8498,N_8652);
or U9391 (N_9391,N_8371,N_8871);
or U9392 (N_9392,N_8876,N_8093);
nand U9393 (N_9393,N_8774,N_8617);
or U9394 (N_9394,N_8545,N_8920);
nor U9395 (N_9395,N_8552,N_8682);
nand U9396 (N_9396,N_8614,N_8639);
or U9397 (N_9397,N_8944,N_8767);
nor U9398 (N_9398,N_8575,N_8032);
xnor U9399 (N_9399,N_8227,N_8893);
nor U9400 (N_9400,N_8427,N_8577);
nor U9401 (N_9401,N_8707,N_8773);
nand U9402 (N_9402,N_8946,N_8338);
nor U9403 (N_9403,N_8880,N_8538);
and U9404 (N_9404,N_8984,N_8143);
xnor U9405 (N_9405,N_8551,N_8062);
xor U9406 (N_9406,N_8259,N_8174);
xnor U9407 (N_9407,N_8320,N_8477);
nor U9408 (N_9408,N_8422,N_8818);
or U9409 (N_9409,N_8592,N_8898);
nor U9410 (N_9410,N_8640,N_8783);
or U9411 (N_9411,N_8281,N_8844);
and U9412 (N_9412,N_8386,N_8567);
xnor U9413 (N_9413,N_8023,N_8327);
nand U9414 (N_9414,N_8241,N_8249);
or U9415 (N_9415,N_8169,N_8956);
and U9416 (N_9416,N_8075,N_8204);
nand U9417 (N_9417,N_8519,N_8036);
nand U9418 (N_9418,N_8926,N_8288);
nor U9419 (N_9419,N_8822,N_8207);
or U9420 (N_9420,N_8983,N_8271);
nand U9421 (N_9421,N_8206,N_8470);
xor U9422 (N_9422,N_8446,N_8570);
xnor U9423 (N_9423,N_8661,N_8845);
nand U9424 (N_9424,N_8974,N_8775);
and U9425 (N_9425,N_8672,N_8370);
nor U9426 (N_9426,N_8503,N_8734);
nor U9427 (N_9427,N_8440,N_8815);
nor U9428 (N_9428,N_8681,N_8283);
xor U9429 (N_9429,N_8116,N_8115);
xnor U9430 (N_9430,N_8119,N_8366);
or U9431 (N_9431,N_8365,N_8456);
nand U9432 (N_9432,N_8935,N_8330);
or U9433 (N_9433,N_8210,N_8988);
nor U9434 (N_9434,N_8766,N_8275);
nand U9435 (N_9435,N_8889,N_8558);
nand U9436 (N_9436,N_8527,N_8616);
nor U9437 (N_9437,N_8299,N_8799);
and U9438 (N_9438,N_8374,N_8489);
xor U9439 (N_9439,N_8990,N_8608);
nand U9440 (N_9440,N_8816,N_8137);
and U9441 (N_9441,N_8823,N_8840);
and U9442 (N_9442,N_8377,N_8297);
nor U9443 (N_9443,N_8500,N_8952);
and U9444 (N_9444,N_8704,N_8121);
nor U9445 (N_9445,N_8474,N_8873);
or U9446 (N_9446,N_8722,N_8167);
or U9447 (N_9447,N_8495,N_8741);
xnor U9448 (N_9448,N_8305,N_8039);
and U9449 (N_9449,N_8193,N_8135);
xnor U9450 (N_9450,N_8638,N_8506);
or U9451 (N_9451,N_8318,N_8105);
nor U9452 (N_9452,N_8179,N_8581);
nor U9453 (N_9453,N_8123,N_8562);
xor U9454 (N_9454,N_8692,N_8198);
xnor U9455 (N_9455,N_8144,N_8102);
nand U9456 (N_9456,N_8009,N_8548);
and U9457 (N_9457,N_8525,N_8908);
xor U9458 (N_9458,N_8347,N_8126);
nor U9459 (N_9459,N_8209,N_8650);
nand U9460 (N_9460,N_8278,N_8280);
xor U9461 (N_9461,N_8651,N_8255);
nand U9462 (N_9462,N_8533,N_8304);
or U9463 (N_9463,N_8056,N_8450);
and U9464 (N_9464,N_8753,N_8367);
nand U9465 (N_9465,N_8645,N_8441);
or U9466 (N_9466,N_8762,N_8561);
or U9467 (N_9467,N_8099,N_8724);
or U9468 (N_9468,N_8101,N_8694);
and U9469 (N_9469,N_8472,N_8916);
or U9470 (N_9470,N_8759,N_8424);
or U9471 (N_9471,N_8782,N_8997);
xnor U9472 (N_9472,N_8132,N_8932);
nand U9473 (N_9473,N_8497,N_8619);
nor U9474 (N_9474,N_8069,N_8403);
nand U9475 (N_9475,N_8267,N_8223);
and U9476 (N_9476,N_8550,N_8810);
xnor U9477 (N_9477,N_8963,N_8779);
or U9478 (N_9478,N_8735,N_8331);
and U9479 (N_9479,N_8573,N_8378);
nor U9480 (N_9480,N_8139,N_8964);
nand U9481 (N_9481,N_8656,N_8955);
and U9482 (N_9482,N_8098,N_8445);
nand U9483 (N_9483,N_8718,N_8918);
xnor U9484 (N_9484,N_8035,N_8052);
or U9485 (N_9485,N_8125,N_8913);
or U9486 (N_9486,N_8837,N_8621);
xor U9487 (N_9487,N_8603,N_8968);
nor U9488 (N_9488,N_8885,N_8104);
nand U9489 (N_9489,N_8442,N_8430);
nand U9490 (N_9490,N_8475,N_8726);
or U9491 (N_9491,N_8832,N_8948);
or U9492 (N_9492,N_8364,N_8806);
nor U9493 (N_9493,N_8247,N_8872);
xnor U9494 (N_9494,N_8177,N_8930);
nand U9495 (N_9495,N_8376,N_8754);
nor U9496 (N_9496,N_8542,N_8294);
nor U9497 (N_9497,N_8703,N_8047);
or U9498 (N_9498,N_8743,N_8129);
and U9499 (N_9499,N_8201,N_8007);
and U9500 (N_9500,N_8395,N_8688);
nand U9501 (N_9501,N_8864,N_8743);
nand U9502 (N_9502,N_8653,N_8606);
nand U9503 (N_9503,N_8844,N_8664);
and U9504 (N_9504,N_8215,N_8035);
and U9505 (N_9505,N_8167,N_8338);
and U9506 (N_9506,N_8291,N_8009);
xnor U9507 (N_9507,N_8246,N_8563);
nand U9508 (N_9508,N_8472,N_8313);
and U9509 (N_9509,N_8263,N_8961);
nand U9510 (N_9510,N_8925,N_8306);
nand U9511 (N_9511,N_8886,N_8098);
or U9512 (N_9512,N_8048,N_8750);
or U9513 (N_9513,N_8873,N_8874);
or U9514 (N_9514,N_8500,N_8593);
or U9515 (N_9515,N_8108,N_8933);
xnor U9516 (N_9516,N_8849,N_8730);
nor U9517 (N_9517,N_8682,N_8127);
and U9518 (N_9518,N_8978,N_8004);
or U9519 (N_9519,N_8102,N_8282);
and U9520 (N_9520,N_8470,N_8385);
or U9521 (N_9521,N_8596,N_8249);
or U9522 (N_9522,N_8810,N_8904);
and U9523 (N_9523,N_8016,N_8042);
nand U9524 (N_9524,N_8189,N_8091);
and U9525 (N_9525,N_8004,N_8892);
nor U9526 (N_9526,N_8182,N_8352);
and U9527 (N_9527,N_8424,N_8943);
nor U9528 (N_9528,N_8958,N_8254);
nor U9529 (N_9529,N_8402,N_8408);
or U9530 (N_9530,N_8152,N_8860);
nor U9531 (N_9531,N_8448,N_8610);
nand U9532 (N_9532,N_8813,N_8850);
xor U9533 (N_9533,N_8515,N_8034);
and U9534 (N_9534,N_8196,N_8696);
xnor U9535 (N_9535,N_8723,N_8130);
nor U9536 (N_9536,N_8545,N_8728);
or U9537 (N_9537,N_8247,N_8780);
and U9538 (N_9538,N_8617,N_8755);
or U9539 (N_9539,N_8510,N_8243);
or U9540 (N_9540,N_8981,N_8906);
nor U9541 (N_9541,N_8768,N_8182);
nand U9542 (N_9542,N_8788,N_8235);
xnor U9543 (N_9543,N_8565,N_8431);
nor U9544 (N_9544,N_8579,N_8007);
or U9545 (N_9545,N_8685,N_8239);
nand U9546 (N_9546,N_8552,N_8090);
and U9547 (N_9547,N_8156,N_8548);
or U9548 (N_9548,N_8993,N_8064);
nand U9549 (N_9549,N_8936,N_8481);
or U9550 (N_9550,N_8572,N_8197);
or U9551 (N_9551,N_8120,N_8567);
and U9552 (N_9552,N_8961,N_8610);
xor U9553 (N_9553,N_8537,N_8715);
and U9554 (N_9554,N_8527,N_8894);
nand U9555 (N_9555,N_8517,N_8454);
and U9556 (N_9556,N_8811,N_8126);
nor U9557 (N_9557,N_8761,N_8153);
xnor U9558 (N_9558,N_8930,N_8343);
and U9559 (N_9559,N_8332,N_8231);
or U9560 (N_9560,N_8371,N_8034);
nand U9561 (N_9561,N_8238,N_8308);
nand U9562 (N_9562,N_8531,N_8454);
nand U9563 (N_9563,N_8028,N_8957);
xnor U9564 (N_9564,N_8360,N_8558);
nor U9565 (N_9565,N_8338,N_8983);
and U9566 (N_9566,N_8018,N_8349);
nor U9567 (N_9567,N_8864,N_8678);
nand U9568 (N_9568,N_8603,N_8191);
xor U9569 (N_9569,N_8243,N_8723);
nor U9570 (N_9570,N_8003,N_8195);
and U9571 (N_9571,N_8303,N_8361);
xor U9572 (N_9572,N_8724,N_8552);
xor U9573 (N_9573,N_8060,N_8094);
xor U9574 (N_9574,N_8620,N_8819);
nor U9575 (N_9575,N_8140,N_8324);
nor U9576 (N_9576,N_8280,N_8708);
xnor U9577 (N_9577,N_8920,N_8863);
nor U9578 (N_9578,N_8644,N_8243);
and U9579 (N_9579,N_8518,N_8531);
and U9580 (N_9580,N_8045,N_8313);
xor U9581 (N_9581,N_8105,N_8013);
nor U9582 (N_9582,N_8725,N_8805);
xor U9583 (N_9583,N_8390,N_8731);
and U9584 (N_9584,N_8008,N_8018);
nor U9585 (N_9585,N_8175,N_8593);
and U9586 (N_9586,N_8569,N_8381);
and U9587 (N_9587,N_8908,N_8423);
nand U9588 (N_9588,N_8226,N_8286);
nor U9589 (N_9589,N_8810,N_8382);
nor U9590 (N_9590,N_8281,N_8645);
and U9591 (N_9591,N_8080,N_8210);
nor U9592 (N_9592,N_8369,N_8924);
or U9593 (N_9593,N_8684,N_8750);
or U9594 (N_9594,N_8780,N_8889);
and U9595 (N_9595,N_8819,N_8932);
and U9596 (N_9596,N_8450,N_8974);
nand U9597 (N_9597,N_8396,N_8297);
and U9598 (N_9598,N_8266,N_8863);
and U9599 (N_9599,N_8796,N_8806);
xnor U9600 (N_9600,N_8718,N_8249);
xnor U9601 (N_9601,N_8323,N_8116);
nand U9602 (N_9602,N_8032,N_8975);
nor U9603 (N_9603,N_8887,N_8201);
nand U9604 (N_9604,N_8270,N_8907);
nor U9605 (N_9605,N_8419,N_8184);
or U9606 (N_9606,N_8996,N_8763);
nor U9607 (N_9607,N_8808,N_8494);
xnor U9608 (N_9608,N_8936,N_8295);
nand U9609 (N_9609,N_8701,N_8962);
nor U9610 (N_9610,N_8635,N_8515);
or U9611 (N_9611,N_8197,N_8005);
nand U9612 (N_9612,N_8745,N_8799);
or U9613 (N_9613,N_8823,N_8043);
nand U9614 (N_9614,N_8297,N_8664);
and U9615 (N_9615,N_8038,N_8690);
nand U9616 (N_9616,N_8412,N_8622);
and U9617 (N_9617,N_8927,N_8174);
xnor U9618 (N_9618,N_8977,N_8199);
or U9619 (N_9619,N_8601,N_8642);
nor U9620 (N_9620,N_8689,N_8896);
nor U9621 (N_9621,N_8854,N_8634);
or U9622 (N_9622,N_8560,N_8806);
xnor U9623 (N_9623,N_8258,N_8941);
xnor U9624 (N_9624,N_8389,N_8153);
and U9625 (N_9625,N_8826,N_8336);
or U9626 (N_9626,N_8730,N_8603);
nand U9627 (N_9627,N_8320,N_8148);
nand U9628 (N_9628,N_8096,N_8253);
or U9629 (N_9629,N_8938,N_8811);
nand U9630 (N_9630,N_8182,N_8756);
and U9631 (N_9631,N_8064,N_8387);
and U9632 (N_9632,N_8536,N_8988);
or U9633 (N_9633,N_8714,N_8704);
nor U9634 (N_9634,N_8377,N_8089);
nor U9635 (N_9635,N_8262,N_8318);
or U9636 (N_9636,N_8552,N_8487);
and U9637 (N_9637,N_8122,N_8323);
and U9638 (N_9638,N_8760,N_8040);
xnor U9639 (N_9639,N_8332,N_8432);
xnor U9640 (N_9640,N_8694,N_8996);
nand U9641 (N_9641,N_8621,N_8612);
xor U9642 (N_9642,N_8940,N_8968);
xor U9643 (N_9643,N_8263,N_8120);
nor U9644 (N_9644,N_8259,N_8659);
or U9645 (N_9645,N_8587,N_8382);
xor U9646 (N_9646,N_8874,N_8760);
nor U9647 (N_9647,N_8194,N_8745);
nor U9648 (N_9648,N_8476,N_8489);
xnor U9649 (N_9649,N_8161,N_8511);
nor U9650 (N_9650,N_8427,N_8552);
nor U9651 (N_9651,N_8770,N_8896);
xnor U9652 (N_9652,N_8777,N_8065);
or U9653 (N_9653,N_8005,N_8220);
nor U9654 (N_9654,N_8036,N_8471);
nand U9655 (N_9655,N_8216,N_8650);
nand U9656 (N_9656,N_8873,N_8542);
xor U9657 (N_9657,N_8684,N_8439);
and U9658 (N_9658,N_8752,N_8517);
or U9659 (N_9659,N_8239,N_8439);
xnor U9660 (N_9660,N_8086,N_8167);
nor U9661 (N_9661,N_8122,N_8005);
xor U9662 (N_9662,N_8122,N_8076);
nand U9663 (N_9663,N_8403,N_8405);
nand U9664 (N_9664,N_8283,N_8404);
nand U9665 (N_9665,N_8469,N_8545);
xnor U9666 (N_9666,N_8665,N_8708);
nand U9667 (N_9667,N_8132,N_8645);
nand U9668 (N_9668,N_8492,N_8734);
nand U9669 (N_9669,N_8688,N_8611);
xor U9670 (N_9670,N_8173,N_8710);
nand U9671 (N_9671,N_8752,N_8103);
nor U9672 (N_9672,N_8234,N_8724);
or U9673 (N_9673,N_8362,N_8811);
nor U9674 (N_9674,N_8504,N_8051);
or U9675 (N_9675,N_8212,N_8723);
xor U9676 (N_9676,N_8684,N_8198);
nand U9677 (N_9677,N_8504,N_8882);
nor U9678 (N_9678,N_8959,N_8501);
xnor U9679 (N_9679,N_8274,N_8242);
nand U9680 (N_9680,N_8852,N_8047);
or U9681 (N_9681,N_8881,N_8162);
and U9682 (N_9682,N_8936,N_8184);
nand U9683 (N_9683,N_8088,N_8442);
nand U9684 (N_9684,N_8229,N_8745);
or U9685 (N_9685,N_8755,N_8438);
or U9686 (N_9686,N_8550,N_8302);
or U9687 (N_9687,N_8946,N_8009);
nand U9688 (N_9688,N_8916,N_8786);
nor U9689 (N_9689,N_8197,N_8041);
nor U9690 (N_9690,N_8940,N_8156);
or U9691 (N_9691,N_8326,N_8109);
nand U9692 (N_9692,N_8349,N_8877);
and U9693 (N_9693,N_8319,N_8575);
xnor U9694 (N_9694,N_8250,N_8854);
or U9695 (N_9695,N_8455,N_8090);
nand U9696 (N_9696,N_8012,N_8974);
xnor U9697 (N_9697,N_8582,N_8371);
xnor U9698 (N_9698,N_8828,N_8612);
or U9699 (N_9699,N_8841,N_8180);
or U9700 (N_9700,N_8833,N_8444);
and U9701 (N_9701,N_8091,N_8497);
and U9702 (N_9702,N_8396,N_8349);
and U9703 (N_9703,N_8700,N_8179);
xnor U9704 (N_9704,N_8622,N_8920);
nor U9705 (N_9705,N_8685,N_8042);
nor U9706 (N_9706,N_8023,N_8671);
or U9707 (N_9707,N_8822,N_8945);
or U9708 (N_9708,N_8500,N_8331);
xor U9709 (N_9709,N_8652,N_8975);
and U9710 (N_9710,N_8418,N_8069);
or U9711 (N_9711,N_8893,N_8593);
or U9712 (N_9712,N_8596,N_8956);
nor U9713 (N_9713,N_8863,N_8531);
nor U9714 (N_9714,N_8327,N_8205);
or U9715 (N_9715,N_8916,N_8691);
nand U9716 (N_9716,N_8674,N_8952);
nand U9717 (N_9717,N_8152,N_8783);
nor U9718 (N_9718,N_8695,N_8944);
and U9719 (N_9719,N_8800,N_8691);
nor U9720 (N_9720,N_8651,N_8824);
nor U9721 (N_9721,N_8933,N_8959);
xor U9722 (N_9722,N_8332,N_8900);
nor U9723 (N_9723,N_8866,N_8745);
nor U9724 (N_9724,N_8815,N_8940);
nor U9725 (N_9725,N_8709,N_8555);
nand U9726 (N_9726,N_8721,N_8227);
and U9727 (N_9727,N_8976,N_8113);
xor U9728 (N_9728,N_8016,N_8083);
nor U9729 (N_9729,N_8013,N_8621);
nor U9730 (N_9730,N_8696,N_8977);
and U9731 (N_9731,N_8109,N_8575);
and U9732 (N_9732,N_8461,N_8212);
xnor U9733 (N_9733,N_8452,N_8116);
xor U9734 (N_9734,N_8192,N_8862);
nand U9735 (N_9735,N_8089,N_8207);
nand U9736 (N_9736,N_8572,N_8451);
or U9737 (N_9737,N_8224,N_8074);
nor U9738 (N_9738,N_8272,N_8718);
nor U9739 (N_9739,N_8046,N_8520);
and U9740 (N_9740,N_8319,N_8274);
xor U9741 (N_9741,N_8730,N_8964);
nand U9742 (N_9742,N_8914,N_8789);
nor U9743 (N_9743,N_8511,N_8693);
nor U9744 (N_9744,N_8141,N_8364);
xnor U9745 (N_9745,N_8943,N_8211);
xor U9746 (N_9746,N_8800,N_8710);
xor U9747 (N_9747,N_8463,N_8478);
and U9748 (N_9748,N_8079,N_8705);
nor U9749 (N_9749,N_8515,N_8735);
or U9750 (N_9750,N_8827,N_8133);
xnor U9751 (N_9751,N_8774,N_8772);
or U9752 (N_9752,N_8186,N_8947);
nor U9753 (N_9753,N_8638,N_8670);
and U9754 (N_9754,N_8108,N_8371);
xnor U9755 (N_9755,N_8365,N_8847);
nor U9756 (N_9756,N_8002,N_8517);
nand U9757 (N_9757,N_8548,N_8088);
or U9758 (N_9758,N_8698,N_8388);
nand U9759 (N_9759,N_8268,N_8744);
nor U9760 (N_9760,N_8105,N_8048);
xor U9761 (N_9761,N_8777,N_8321);
and U9762 (N_9762,N_8355,N_8685);
or U9763 (N_9763,N_8592,N_8658);
xor U9764 (N_9764,N_8533,N_8450);
xnor U9765 (N_9765,N_8736,N_8358);
or U9766 (N_9766,N_8040,N_8801);
nand U9767 (N_9767,N_8570,N_8995);
and U9768 (N_9768,N_8175,N_8289);
or U9769 (N_9769,N_8082,N_8607);
nand U9770 (N_9770,N_8992,N_8009);
xnor U9771 (N_9771,N_8854,N_8237);
nor U9772 (N_9772,N_8375,N_8089);
or U9773 (N_9773,N_8162,N_8929);
xnor U9774 (N_9774,N_8132,N_8084);
xnor U9775 (N_9775,N_8015,N_8922);
nand U9776 (N_9776,N_8474,N_8030);
xor U9777 (N_9777,N_8173,N_8015);
nand U9778 (N_9778,N_8201,N_8727);
nand U9779 (N_9779,N_8762,N_8043);
xor U9780 (N_9780,N_8333,N_8129);
xnor U9781 (N_9781,N_8034,N_8459);
xor U9782 (N_9782,N_8649,N_8794);
or U9783 (N_9783,N_8230,N_8794);
and U9784 (N_9784,N_8126,N_8859);
nor U9785 (N_9785,N_8732,N_8306);
nor U9786 (N_9786,N_8791,N_8811);
nor U9787 (N_9787,N_8202,N_8121);
nor U9788 (N_9788,N_8125,N_8838);
and U9789 (N_9789,N_8397,N_8912);
and U9790 (N_9790,N_8090,N_8172);
xor U9791 (N_9791,N_8637,N_8781);
and U9792 (N_9792,N_8875,N_8995);
xnor U9793 (N_9793,N_8816,N_8604);
and U9794 (N_9794,N_8472,N_8861);
or U9795 (N_9795,N_8224,N_8315);
and U9796 (N_9796,N_8430,N_8641);
nand U9797 (N_9797,N_8916,N_8893);
and U9798 (N_9798,N_8931,N_8605);
xnor U9799 (N_9799,N_8424,N_8464);
nand U9800 (N_9800,N_8403,N_8974);
nand U9801 (N_9801,N_8102,N_8517);
and U9802 (N_9802,N_8518,N_8817);
nand U9803 (N_9803,N_8307,N_8107);
or U9804 (N_9804,N_8081,N_8734);
or U9805 (N_9805,N_8210,N_8012);
nor U9806 (N_9806,N_8266,N_8422);
and U9807 (N_9807,N_8085,N_8900);
and U9808 (N_9808,N_8184,N_8780);
xor U9809 (N_9809,N_8121,N_8078);
nor U9810 (N_9810,N_8128,N_8421);
nor U9811 (N_9811,N_8406,N_8763);
nand U9812 (N_9812,N_8012,N_8938);
and U9813 (N_9813,N_8847,N_8277);
and U9814 (N_9814,N_8120,N_8292);
nor U9815 (N_9815,N_8795,N_8378);
nand U9816 (N_9816,N_8498,N_8926);
xor U9817 (N_9817,N_8564,N_8829);
nand U9818 (N_9818,N_8108,N_8104);
nor U9819 (N_9819,N_8408,N_8269);
nand U9820 (N_9820,N_8867,N_8997);
xnor U9821 (N_9821,N_8586,N_8858);
nor U9822 (N_9822,N_8482,N_8942);
xor U9823 (N_9823,N_8822,N_8167);
nor U9824 (N_9824,N_8360,N_8116);
or U9825 (N_9825,N_8262,N_8584);
nor U9826 (N_9826,N_8174,N_8309);
or U9827 (N_9827,N_8970,N_8575);
or U9828 (N_9828,N_8251,N_8400);
nand U9829 (N_9829,N_8592,N_8574);
nand U9830 (N_9830,N_8540,N_8217);
nand U9831 (N_9831,N_8896,N_8390);
and U9832 (N_9832,N_8064,N_8702);
xor U9833 (N_9833,N_8177,N_8789);
xnor U9834 (N_9834,N_8629,N_8096);
or U9835 (N_9835,N_8284,N_8489);
xor U9836 (N_9836,N_8681,N_8600);
nand U9837 (N_9837,N_8668,N_8801);
nand U9838 (N_9838,N_8186,N_8068);
or U9839 (N_9839,N_8322,N_8288);
xor U9840 (N_9840,N_8557,N_8253);
nand U9841 (N_9841,N_8344,N_8207);
nand U9842 (N_9842,N_8337,N_8741);
nor U9843 (N_9843,N_8658,N_8906);
xor U9844 (N_9844,N_8300,N_8579);
and U9845 (N_9845,N_8314,N_8793);
nand U9846 (N_9846,N_8389,N_8600);
nand U9847 (N_9847,N_8060,N_8757);
or U9848 (N_9848,N_8296,N_8941);
xnor U9849 (N_9849,N_8405,N_8037);
xor U9850 (N_9850,N_8548,N_8311);
nand U9851 (N_9851,N_8503,N_8516);
xnor U9852 (N_9852,N_8336,N_8982);
nand U9853 (N_9853,N_8835,N_8887);
nand U9854 (N_9854,N_8421,N_8299);
or U9855 (N_9855,N_8346,N_8221);
or U9856 (N_9856,N_8576,N_8446);
and U9857 (N_9857,N_8329,N_8944);
and U9858 (N_9858,N_8035,N_8585);
nand U9859 (N_9859,N_8577,N_8957);
nor U9860 (N_9860,N_8525,N_8670);
and U9861 (N_9861,N_8965,N_8943);
or U9862 (N_9862,N_8919,N_8185);
nand U9863 (N_9863,N_8881,N_8435);
xor U9864 (N_9864,N_8422,N_8173);
xor U9865 (N_9865,N_8115,N_8055);
xor U9866 (N_9866,N_8774,N_8585);
xor U9867 (N_9867,N_8825,N_8753);
nand U9868 (N_9868,N_8365,N_8167);
nand U9869 (N_9869,N_8408,N_8737);
and U9870 (N_9870,N_8561,N_8706);
nand U9871 (N_9871,N_8274,N_8178);
nor U9872 (N_9872,N_8322,N_8163);
nor U9873 (N_9873,N_8378,N_8458);
xnor U9874 (N_9874,N_8317,N_8846);
or U9875 (N_9875,N_8747,N_8464);
and U9876 (N_9876,N_8049,N_8709);
and U9877 (N_9877,N_8029,N_8538);
and U9878 (N_9878,N_8006,N_8995);
or U9879 (N_9879,N_8891,N_8926);
nor U9880 (N_9880,N_8761,N_8137);
nand U9881 (N_9881,N_8665,N_8797);
nand U9882 (N_9882,N_8480,N_8749);
nor U9883 (N_9883,N_8878,N_8009);
nand U9884 (N_9884,N_8877,N_8443);
or U9885 (N_9885,N_8861,N_8189);
nor U9886 (N_9886,N_8700,N_8757);
nand U9887 (N_9887,N_8776,N_8611);
xor U9888 (N_9888,N_8527,N_8231);
and U9889 (N_9889,N_8429,N_8718);
xor U9890 (N_9890,N_8300,N_8473);
xnor U9891 (N_9891,N_8483,N_8707);
and U9892 (N_9892,N_8744,N_8826);
and U9893 (N_9893,N_8171,N_8324);
xnor U9894 (N_9894,N_8181,N_8225);
or U9895 (N_9895,N_8762,N_8922);
nand U9896 (N_9896,N_8701,N_8271);
nand U9897 (N_9897,N_8424,N_8491);
or U9898 (N_9898,N_8873,N_8860);
nor U9899 (N_9899,N_8837,N_8520);
xnor U9900 (N_9900,N_8391,N_8819);
nand U9901 (N_9901,N_8941,N_8486);
nor U9902 (N_9902,N_8163,N_8308);
nand U9903 (N_9903,N_8941,N_8978);
nand U9904 (N_9904,N_8362,N_8028);
nor U9905 (N_9905,N_8003,N_8844);
nor U9906 (N_9906,N_8160,N_8766);
or U9907 (N_9907,N_8605,N_8248);
or U9908 (N_9908,N_8405,N_8689);
or U9909 (N_9909,N_8021,N_8383);
nand U9910 (N_9910,N_8726,N_8471);
or U9911 (N_9911,N_8669,N_8327);
or U9912 (N_9912,N_8987,N_8188);
nor U9913 (N_9913,N_8005,N_8006);
nor U9914 (N_9914,N_8382,N_8966);
and U9915 (N_9915,N_8658,N_8634);
nand U9916 (N_9916,N_8808,N_8239);
nor U9917 (N_9917,N_8611,N_8599);
and U9918 (N_9918,N_8508,N_8299);
or U9919 (N_9919,N_8908,N_8719);
nand U9920 (N_9920,N_8570,N_8135);
nand U9921 (N_9921,N_8296,N_8473);
or U9922 (N_9922,N_8604,N_8651);
nand U9923 (N_9923,N_8115,N_8571);
and U9924 (N_9924,N_8523,N_8030);
nand U9925 (N_9925,N_8939,N_8187);
xnor U9926 (N_9926,N_8768,N_8763);
xor U9927 (N_9927,N_8764,N_8758);
nand U9928 (N_9928,N_8144,N_8872);
nand U9929 (N_9929,N_8540,N_8255);
xnor U9930 (N_9930,N_8011,N_8779);
xor U9931 (N_9931,N_8089,N_8116);
or U9932 (N_9932,N_8085,N_8648);
nor U9933 (N_9933,N_8604,N_8804);
nor U9934 (N_9934,N_8800,N_8804);
nor U9935 (N_9935,N_8142,N_8694);
and U9936 (N_9936,N_8517,N_8240);
nand U9937 (N_9937,N_8203,N_8967);
and U9938 (N_9938,N_8528,N_8373);
nand U9939 (N_9939,N_8614,N_8954);
and U9940 (N_9940,N_8332,N_8863);
or U9941 (N_9941,N_8781,N_8400);
nand U9942 (N_9942,N_8623,N_8075);
or U9943 (N_9943,N_8159,N_8941);
and U9944 (N_9944,N_8410,N_8725);
nand U9945 (N_9945,N_8560,N_8406);
and U9946 (N_9946,N_8470,N_8093);
nor U9947 (N_9947,N_8761,N_8306);
nand U9948 (N_9948,N_8892,N_8124);
and U9949 (N_9949,N_8361,N_8417);
and U9950 (N_9950,N_8155,N_8782);
nand U9951 (N_9951,N_8974,N_8718);
and U9952 (N_9952,N_8462,N_8693);
nand U9953 (N_9953,N_8059,N_8872);
nand U9954 (N_9954,N_8323,N_8639);
nor U9955 (N_9955,N_8081,N_8036);
or U9956 (N_9956,N_8304,N_8950);
or U9957 (N_9957,N_8001,N_8633);
nor U9958 (N_9958,N_8370,N_8612);
and U9959 (N_9959,N_8821,N_8599);
nand U9960 (N_9960,N_8713,N_8022);
nor U9961 (N_9961,N_8008,N_8678);
and U9962 (N_9962,N_8334,N_8785);
or U9963 (N_9963,N_8298,N_8552);
xor U9964 (N_9964,N_8231,N_8559);
xor U9965 (N_9965,N_8412,N_8851);
xnor U9966 (N_9966,N_8440,N_8402);
and U9967 (N_9967,N_8772,N_8157);
or U9968 (N_9968,N_8417,N_8365);
nand U9969 (N_9969,N_8774,N_8426);
nor U9970 (N_9970,N_8525,N_8891);
nor U9971 (N_9971,N_8244,N_8366);
nand U9972 (N_9972,N_8842,N_8589);
or U9973 (N_9973,N_8446,N_8575);
and U9974 (N_9974,N_8218,N_8579);
or U9975 (N_9975,N_8990,N_8841);
nor U9976 (N_9976,N_8334,N_8624);
xor U9977 (N_9977,N_8447,N_8287);
nand U9978 (N_9978,N_8763,N_8924);
xnor U9979 (N_9979,N_8039,N_8901);
nand U9980 (N_9980,N_8878,N_8362);
or U9981 (N_9981,N_8213,N_8893);
xor U9982 (N_9982,N_8221,N_8140);
xnor U9983 (N_9983,N_8153,N_8965);
nor U9984 (N_9984,N_8278,N_8419);
xnor U9985 (N_9985,N_8815,N_8826);
xor U9986 (N_9986,N_8746,N_8780);
or U9987 (N_9987,N_8825,N_8254);
nand U9988 (N_9988,N_8848,N_8199);
or U9989 (N_9989,N_8277,N_8707);
or U9990 (N_9990,N_8305,N_8114);
nand U9991 (N_9991,N_8489,N_8070);
xnor U9992 (N_9992,N_8570,N_8895);
nor U9993 (N_9993,N_8162,N_8167);
xor U9994 (N_9994,N_8889,N_8591);
xnor U9995 (N_9995,N_8760,N_8895);
nand U9996 (N_9996,N_8209,N_8957);
and U9997 (N_9997,N_8076,N_8420);
nor U9998 (N_9998,N_8957,N_8906);
or U9999 (N_9999,N_8602,N_8182);
xnor U10000 (N_10000,N_9109,N_9203);
or U10001 (N_10001,N_9172,N_9750);
xnor U10002 (N_10002,N_9018,N_9191);
nand U10003 (N_10003,N_9804,N_9965);
and U10004 (N_10004,N_9884,N_9133);
xor U10005 (N_10005,N_9800,N_9945);
nand U10006 (N_10006,N_9959,N_9817);
xor U10007 (N_10007,N_9230,N_9140);
nor U10008 (N_10008,N_9051,N_9815);
nand U10009 (N_10009,N_9714,N_9485);
nor U10010 (N_10010,N_9527,N_9591);
and U10011 (N_10011,N_9154,N_9881);
nand U10012 (N_10012,N_9869,N_9196);
xnor U10013 (N_10013,N_9859,N_9938);
or U10014 (N_10014,N_9032,N_9242);
or U10015 (N_10015,N_9093,N_9941);
xnor U10016 (N_10016,N_9743,N_9098);
or U10017 (N_10017,N_9440,N_9165);
nor U10018 (N_10018,N_9180,N_9977);
nor U10019 (N_10019,N_9736,N_9957);
nand U10020 (N_10020,N_9946,N_9807);
nor U10021 (N_10021,N_9808,N_9811);
xnor U10022 (N_10022,N_9748,N_9919);
xnor U10023 (N_10023,N_9495,N_9390);
xor U10024 (N_10024,N_9183,N_9323);
nand U10025 (N_10025,N_9371,N_9512);
xnor U10026 (N_10026,N_9972,N_9711);
nor U10027 (N_10027,N_9548,N_9339);
and U10028 (N_10028,N_9493,N_9353);
nand U10029 (N_10029,N_9901,N_9491);
or U10030 (N_10030,N_9231,N_9094);
nand U10031 (N_10031,N_9691,N_9052);
nor U10032 (N_10032,N_9973,N_9505);
and U10033 (N_10033,N_9064,N_9215);
xnor U10034 (N_10034,N_9818,N_9653);
and U10035 (N_10035,N_9942,N_9129);
and U10036 (N_10036,N_9741,N_9664);
nor U10037 (N_10037,N_9651,N_9606);
or U10038 (N_10038,N_9749,N_9697);
nor U10039 (N_10039,N_9285,N_9223);
nand U10040 (N_10040,N_9274,N_9541);
xnor U10041 (N_10041,N_9333,N_9564);
nand U10042 (N_10042,N_9663,N_9236);
nor U10043 (N_10043,N_9668,N_9074);
xor U10044 (N_10044,N_9650,N_9515);
and U10045 (N_10045,N_9991,N_9783);
or U10046 (N_10046,N_9506,N_9825);
nor U10047 (N_10047,N_9526,N_9683);
or U10048 (N_10048,N_9772,N_9602);
xnor U10049 (N_10049,N_9598,N_9906);
nand U10050 (N_10050,N_9717,N_9573);
or U10051 (N_10051,N_9954,N_9028);
xnor U10052 (N_10052,N_9340,N_9089);
or U10053 (N_10053,N_9923,N_9571);
xor U10054 (N_10054,N_9304,N_9417);
and U10055 (N_10055,N_9130,N_9226);
nand U10056 (N_10056,N_9213,N_9368);
xnor U10057 (N_10057,N_9587,N_9160);
nand U10058 (N_10058,N_9570,N_9559);
nand U10059 (N_10059,N_9656,N_9331);
nor U10060 (N_10060,N_9135,N_9915);
and U10061 (N_10061,N_9712,N_9574);
xor U10062 (N_10062,N_9473,N_9828);
nor U10063 (N_10063,N_9674,N_9437);
nor U10064 (N_10064,N_9284,N_9354);
nor U10065 (N_10065,N_9292,N_9062);
and U10066 (N_10066,N_9856,N_9855);
and U10067 (N_10067,N_9747,N_9418);
xor U10068 (N_10068,N_9734,N_9289);
and U10069 (N_10069,N_9100,N_9806);
xor U10070 (N_10070,N_9115,N_9192);
nor U10071 (N_10071,N_9532,N_9374);
or U10072 (N_10072,N_9561,N_9623);
nor U10073 (N_10073,N_9426,N_9775);
nand U10074 (N_10074,N_9865,N_9410);
nor U10075 (N_10075,N_9551,N_9150);
nor U10076 (N_10076,N_9534,N_9763);
nand U10077 (N_10077,N_9992,N_9194);
xor U10078 (N_10078,N_9488,N_9083);
xnor U10079 (N_10079,N_9731,N_9258);
and U10080 (N_10080,N_9975,N_9005);
or U10081 (N_10081,N_9886,N_9301);
nor U10082 (N_10082,N_9517,N_9634);
and U10083 (N_10083,N_9812,N_9720);
xor U10084 (N_10084,N_9852,N_9389);
xor U10085 (N_10085,N_9616,N_9842);
nor U10086 (N_10086,N_9398,N_9281);
nor U10087 (N_10087,N_9306,N_9680);
and U10088 (N_10088,N_9829,N_9609);
nor U10089 (N_10089,N_9890,N_9250);
or U10090 (N_10090,N_9996,N_9948);
and U10091 (N_10091,N_9696,N_9624);
or U10092 (N_10092,N_9268,N_9472);
nand U10093 (N_10093,N_9703,N_9466);
and U10094 (N_10094,N_9672,N_9279);
and U10095 (N_10095,N_9420,N_9006);
or U10096 (N_10096,N_9630,N_9900);
nor U10097 (N_10097,N_9603,N_9294);
or U10098 (N_10098,N_9214,N_9404);
or U10099 (N_10099,N_9413,N_9873);
and U10100 (N_10100,N_9197,N_9518);
and U10101 (N_10101,N_9536,N_9332);
nand U10102 (N_10102,N_9870,N_9102);
and U10103 (N_10103,N_9091,N_9361);
and U10104 (N_10104,N_9228,N_9670);
nor U10105 (N_10105,N_9925,N_9516);
xnor U10106 (N_10106,N_9839,N_9117);
or U10107 (N_10107,N_9928,N_9047);
or U10108 (N_10108,N_9406,N_9146);
and U10109 (N_10109,N_9500,N_9016);
or U10110 (N_10110,N_9202,N_9246);
and U10111 (N_10111,N_9845,N_9857);
and U10112 (N_10112,N_9464,N_9320);
xnor U10113 (N_10113,N_9070,N_9953);
and U10114 (N_10114,N_9921,N_9468);
nand U10115 (N_10115,N_9907,N_9759);
xnor U10116 (N_10116,N_9378,N_9805);
and U10117 (N_10117,N_9596,N_9365);
or U10118 (N_10118,N_9955,N_9127);
xor U10119 (N_10119,N_9438,N_9308);
or U10120 (N_10120,N_9586,N_9987);
or U10121 (N_10121,N_9694,N_9961);
or U10122 (N_10122,N_9029,N_9357);
nor U10123 (N_10123,N_9513,N_9033);
xnor U10124 (N_10124,N_9163,N_9756);
and U10125 (N_10125,N_9964,N_9732);
and U10126 (N_10126,N_9958,N_9317);
nor U10127 (N_10127,N_9178,N_9055);
nor U10128 (N_10128,N_9065,N_9677);
nand U10129 (N_10129,N_9531,N_9833);
nor U10130 (N_10130,N_9004,N_9036);
xor U10131 (N_10131,N_9187,N_9729);
and U10132 (N_10132,N_9208,N_9170);
nand U10133 (N_10133,N_9695,N_9045);
nor U10134 (N_10134,N_9034,N_9142);
or U10135 (N_10135,N_9149,N_9988);
or U10136 (N_10136,N_9261,N_9621);
nand U10137 (N_10137,N_9580,N_9793);
or U10138 (N_10138,N_9899,N_9782);
nand U10139 (N_10139,N_9200,N_9579);
nor U10140 (N_10140,N_9897,N_9838);
nor U10141 (N_10141,N_9158,N_9847);
nor U10142 (N_10142,N_9380,N_9421);
nand U10143 (N_10143,N_9066,N_9943);
xor U10144 (N_10144,N_9244,N_9479);
xnor U10145 (N_10145,N_9920,N_9400);
xor U10146 (N_10146,N_9902,N_9787);
nand U10147 (N_10147,N_9940,N_9199);
and U10148 (N_10148,N_9983,N_9903);
and U10149 (N_10149,N_9085,N_9742);
and U10150 (N_10150,N_9038,N_9792);
xnor U10151 (N_10151,N_9234,N_9665);
xnor U10152 (N_10152,N_9978,N_9644);
nand U10153 (N_10153,N_9131,N_9309);
and U10154 (N_10154,N_9022,N_9666);
xor U10155 (N_10155,N_9872,N_9264);
and U10156 (N_10156,N_9416,N_9824);
nor U10157 (N_10157,N_9757,N_9726);
nand U10158 (N_10158,N_9046,N_9635);
and U10159 (N_10159,N_9166,N_9583);
or U10160 (N_10160,N_9898,N_9463);
and U10161 (N_10161,N_9471,N_9728);
or U10162 (N_10162,N_9201,N_9222);
xnor U10163 (N_10163,N_9467,N_9990);
and U10164 (N_10164,N_9862,N_9615);
and U10165 (N_10165,N_9498,N_9851);
nand U10166 (N_10166,N_9181,N_9090);
xor U10167 (N_10167,N_9311,N_9409);
nand U10168 (N_10168,N_9642,N_9056);
nand U10169 (N_10169,N_9751,N_9871);
and U10170 (N_10170,N_9015,N_9917);
nor U10171 (N_10171,N_9545,N_9275);
nand U10172 (N_10172,N_9342,N_9701);
and U10173 (N_10173,N_9947,N_9295);
nor U10174 (N_10174,N_9290,N_9359);
or U10175 (N_10175,N_9575,N_9071);
or U10176 (N_10176,N_9069,N_9027);
xnor U10177 (N_10177,N_9486,N_9931);
xor U10178 (N_10178,N_9894,N_9888);
nor U10179 (N_10179,N_9622,N_9522);
xor U10180 (N_10180,N_9219,N_9985);
or U10181 (N_10181,N_9177,N_9989);
or U10182 (N_10182,N_9533,N_9584);
nand U10183 (N_10183,N_9648,N_9709);
or U10184 (N_10184,N_9235,N_9278);
and U10185 (N_10185,N_9035,N_9567);
xnor U10186 (N_10186,N_9879,N_9174);
xor U10187 (N_10187,N_9224,N_9451);
and U10188 (N_10188,N_9723,N_9162);
and U10189 (N_10189,N_9073,N_9023);
and U10190 (N_10190,N_9009,N_9998);
or U10191 (N_10191,N_9831,N_9684);
xnor U10192 (N_10192,N_9153,N_9040);
nand U10193 (N_10193,N_9508,N_9067);
xnor U10194 (N_10194,N_9535,N_9576);
nor U10195 (N_10195,N_9863,N_9492);
and U10196 (N_10196,N_9474,N_9511);
nor U10197 (N_10197,N_9362,N_9003);
or U10198 (N_10198,N_9537,N_9169);
and U10199 (N_10199,N_9735,N_9345);
or U10200 (N_10200,N_9552,N_9314);
nor U10201 (N_10201,N_9446,N_9976);
and U10202 (N_10202,N_9654,N_9351);
and U10203 (N_10203,N_9692,N_9316);
nand U10204 (N_10204,N_9685,N_9277);
or U10205 (N_10205,N_9509,N_9381);
or U10206 (N_10206,N_9836,N_9913);
nand U10207 (N_10207,N_9218,N_9179);
or U10208 (N_10208,N_9761,N_9360);
nor U10209 (N_10209,N_9638,N_9072);
xor U10210 (N_10210,N_9053,N_9352);
nor U10211 (N_10211,N_9819,N_9452);
and U10212 (N_10212,N_9786,N_9103);
nand U10213 (N_10213,N_9627,N_9001);
nand U10214 (N_10214,N_9568,N_9893);
and U10215 (N_10215,N_9427,N_9781);
or U10216 (N_10216,N_9119,N_9594);
nand U10217 (N_10217,N_9335,N_9408);
and U10218 (N_10218,N_9713,N_9929);
or U10219 (N_10219,N_9291,N_9245);
xnor U10220 (N_10220,N_9431,N_9675);
nor U10221 (N_10221,N_9021,N_9844);
and U10222 (N_10222,N_9265,N_9979);
nor U10223 (N_10223,N_9254,N_9415);
xnor U10224 (N_10224,N_9789,N_9303);
nand U10225 (N_10225,N_9676,N_9765);
nor U10226 (N_10226,N_9671,N_9971);
and U10227 (N_10227,N_9310,N_9126);
nor U10228 (N_10228,N_9962,N_9529);
nor U10229 (N_10229,N_9096,N_9758);
nor U10230 (N_10230,N_9106,N_9966);
or U10231 (N_10231,N_9762,N_9496);
xor U10232 (N_10232,N_9601,N_9367);
nor U10233 (N_10233,N_9049,N_9356);
or U10234 (N_10234,N_9784,N_9476);
and U10235 (N_10235,N_9041,N_9521);
or U10236 (N_10236,N_9547,N_9514);
xor U10237 (N_10237,N_9530,N_9257);
or U10238 (N_10238,N_9061,N_9443);
nand U10239 (N_10239,N_9739,N_9950);
nor U10240 (N_10240,N_9483,N_9539);
nor U10241 (N_10241,N_9210,N_9746);
or U10242 (N_10242,N_9502,N_9614);
xor U10243 (N_10243,N_9707,N_9995);
nor U10244 (N_10244,N_9039,N_9827);
and U10245 (N_10245,N_9436,N_9263);
xor U10246 (N_10246,N_9058,N_9708);
and U10247 (N_10247,N_9366,N_9050);
or U10248 (N_10248,N_9444,N_9148);
nand U10249 (N_10249,N_9841,N_9935);
and U10250 (N_10250,N_9075,N_9937);
and U10251 (N_10251,N_9850,N_9233);
nand U10252 (N_10252,N_9867,N_9424);
nor U10253 (N_10253,N_9113,N_9286);
nor U10254 (N_10254,N_9114,N_9910);
nand U10255 (N_10255,N_9092,N_9132);
nor U10256 (N_10256,N_9974,N_9271);
xnor U10257 (N_10257,N_9143,N_9689);
or U10258 (N_10258,N_9462,N_9877);
xor U10259 (N_10259,N_9253,N_9249);
nand U10260 (N_10260,N_9791,N_9423);
xnor U10261 (N_10261,N_9324,N_9853);
or U10262 (N_10262,N_9889,N_9608);
nand U10263 (N_10263,N_9704,N_9188);
or U10264 (N_10264,N_9549,N_9956);
nor U10265 (N_10265,N_9328,N_9382);
xnor U10266 (N_10266,N_9364,N_9840);
or U10267 (N_10267,N_9737,N_9101);
and U10268 (N_10268,N_9238,N_9814);
or U10269 (N_10269,N_9702,N_9383);
or U10270 (N_10270,N_9318,N_9076);
xnor U10271 (N_10271,N_9330,N_9740);
nor U10272 (N_10272,N_9391,N_9315);
or U10273 (N_10273,N_9725,N_9002);
or U10274 (N_10274,N_9984,N_9393);
xor U10275 (N_10275,N_9283,N_9010);
nor U10276 (N_10276,N_9540,N_9087);
nand U10277 (N_10277,N_9667,N_9459);
and U10278 (N_10278,N_9256,N_9399);
nand U10279 (N_10279,N_9447,N_9754);
xor U10280 (N_10280,N_9497,N_9456);
or U10281 (N_10281,N_9885,N_9874);
or U10282 (N_10282,N_9661,N_9428);
nor U10283 (N_10283,N_9110,N_9487);
or U10284 (N_10284,N_9773,N_9790);
nor U10285 (N_10285,N_9585,N_9013);
nand U10286 (N_10286,N_9625,N_9293);
xor U10287 (N_10287,N_9057,N_9590);
nor U10288 (N_10288,N_9730,N_9597);
and U10289 (N_10289,N_9240,N_9217);
or U10290 (N_10290,N_9878,N_9123);
xnor U10291 (N_10291,N_9569,N_9429);
or U10292 (N_10292,N_9344,N_9558);
xor U10293 (N_10293,N_9449,N_9599);
and U10294 (N_10294,N_9700,N_9933);
or U10295 (N_10295,N_9771,N_9255);
and U10296 (N_10296,N_9718,N_9024);
and U10297 (N_10297,N_9422,N_9876);
xnor U10298 (N_10298,N_9305,N_9145);
xor U10299 (N_10299,N_9124,N_9760);
xor U10300 (N_10300,N_9312,N_9523);
nand U10301 (N_10301,N_9778,N_9767);
nor U10302 (N_10302,N_9280,N_9394);
xnor U10303 (N_10303,N_9430,N_9849);
and U10304 (N_10304,N_9252,N_9669);
nor U10305 (N_10305,N_9647,N_9403);
nor U10306 (N_10306,N_9078,N_9116);
and U10307 (N_10307,N_9626,N_9068);
xor U10308 (N_10308,N_9823,N_9780);
or U10309 (N_10309,N_9134,N_9733);
nand U10310 (N_10310,N_9769,N_9572);
or U10311 (N_10311,N_9593,N_9875);
nand U10312 (N_10312,N_9081,N_9809);
or U10313 (N_10313,N_9402,N_9544);
nor U10314 (N_10314,N_9588,N_9682);
nand U10315 (N_10315,N_9348,N_9225);
and U10316 (N_10316,N_9337,N_9450);
nand U10317 (N_10317,N_9396,N_9721);
and U10318 (N_10318,N_9138,N_9826);
xor U10319 (N_10319,N_9205,N_9848);
nand U10320 (N_10320,N_9846,N_9543);
nor U10321 (N_10321,N_9097,N_9834);
nor U10322 (N_10322,N_9813,N_9687);
or U10323 (N_10323,N_9031,N_9026);
or U10324 (N_10324,N_9980,N_9017);
nand U10325 (N_10325,N_9952,N_9916);
and U10326 (N_10326,N_9538,N_9141);
nor U10327 (N_10327,N_9908,N_9611);
xor U10328 (N_10328,N_9195,N_9397);
nand U10329 (N_10329,N_9457,N_9193);
and U10330 (N_10330,N_9854,N_9475);
xor U10331 (N_10331,N_9722,N_9930);
nor U10332 (N_10332,N_9128,N_9059);
nor U10333 (N_10333,N_9560,N_9477);
nand U10334 (N_10334,N_9470,N_9414);
nand U10335 (N_10335,N_9649,N_9307);
nand U10336 (N_10336,N_9904,N_9241);
or U10337 (N_10337,N_9122,N_9358);
and U10338 (N_10338,N_9745,N_9489);
or U10339 (N_10339,N_9341,N_9251);
and U10340 (N_10340,N_9273,N_9816);
and U10341 (N_10341,N_9678,N_9657);
or U10342 (N_10342,N_9830,N_9288);
nor U10343 (N_10343,N_9768,N_9715);
nor U10344 (N_10344,N_9296,N_9607);
xnor U10345 (N_10345,N_9433,N_9997);
nand U10346 (N_10346,N_9519,N_9660);
xor U10347 (N_10347,N_9080,N_9788);
nand U10348 (N_10348,N_9764,N_9484);
or U10349 (N_10349,N_9243,N_9555);
or U10350 (N_10350,N_9581,N_9799);
xnor U10351 (N_10351,N_9480,N_9088);
xor U10352 (N_10352,N_9125,N_9982);
and U10353 (N_10353,N_9465,N_9266);
and U10354 (N_10354,N_9766,N_9895);
xnor U10355 (N_10355,N_9460,N_9355);
xor U10356 (N_10356,N_9776,N_9944);
or U10357 (N_10357,N_9699,N_9151);
nand U10358 (N_10358,N_9777,N_9774);
nand U10359 (N_10359,N_9453,N_9633);
and U10360 (N_10360,N_9372,N_9343);
and U10361 (N_10361,N_9710,N_9168);
xor U10362 (N_10362,N_9395,N_9407);
and U10363 (N_10363,N_9167,N_9753);
nor U10364 (N_10364,N_9628,N_9282);
and U10365 (N_10365,N_9891,N_9461);
nor U10366 (N_10366,N_9173,N_9385);
nor U10367 (N_10367,N_9880,N_9896);
xor U10368 (N_10368,N_9120,N_9785);
xor U10369 (N_10369,N_9619,N_9797);
nand U10370 (N_10370,N_9688,N_9375);
nand U10371 (N_10371,N_9629,N_9719);
and U10372 (N_10372,N_9520,N_9229);
xor U10373 (N_10373,N_9198,N_9686);
nand U10374 (N_10374,N_9155,N_9000);
nor U10375 (N_10375,N_9562,N_9969);
nor U10376 (N_10376,N_9137,N_9993);
xor U10377 (N_10377,N_9297,N_9970);
xor U10378 (N_10378,N_9209,N_9801);
or U10379 (N_10379,N_9239,N_9837);
nor U10380 (N_10380,N_9216,N_9860);
or U10381 (N_10381,N_9190,N_9963);
or U10382 (N_10382,N_9269,N_9868);
or U10383 (N_10383,N_9960,N_9706);
or U10384 (N_10384,N_9350,N_9442);
or U10385 (N_10385,N_9951,N_9652);
nand U10386 (N_10386,N_9905,N_9858);
or U10387 (N_10387,N_9260,N_9392);
and U10388 (N_10388,N_9600,N_9439);
or U10389 (N_10389,N_9152,N_9206);
nor U10390 (N_10390,N_9327,N_9504);
xor U10391 (N_10391,N_9503,N_9557);
nand U10392 (N_10392,N_9690,N_9159);
and U10393 (N_10393,N_9589,N_9738);
nand U10394 (N_10394,N_9909,N_9104);
nand U10395 (N_10395,N_9025,N_9379);
nand U10396 (N_10396,N_9363,N_9802);
or U10397 (N_10397,N_9482,N_9405);
and U10398 (N_10398,N_9147,N_9144);
nand U10399 (N_10399,N_9646,N_9175);
nor U10400 (N_10400,N_9441,N_9582);
nand U10401 (N_10401,N_9387,N_9967);
or U10402 (N_10402,N_9613,N_9912);
xor U10403 (N_10403,N_9432,N_9752);
nor U10404 (N_10404,N_9820,N_9986);
or U10405 (N_10405,N_9949,N_9086);
nor U10406 (N_10406,N_9319,N_9118);
or U10407 (N_10407,N_9079,N_9556);
xor U10408 (N_10408,N_9494,N_9042);
and U10409 (N_10409,N_9007,N_9563);
and U10410 (N_10410,N_9445,N_9994);
nand U10411 (N_10411,N_9448,N_9554);
nor U10412 (N_10412,N_9592,N_9204);
xnor U10413 (N_10413,N_9370,N_9501);
or U10414 (N_10414,N_9247,N_9546);
nand U10415 (N_10415,N_9645,N_9605);
xor U10416 (N_10416,N_9054,N_9469);
xor U10417 (N_10417,N_9926,N_9156);
nand U10418 (N_10418,N_9866,N_9349);
or U10419 (N_10419,N_9112,N_9161);
xnor U10420 (N_10420,N_9577,N_9048);
xor U10421 (N_10421,N_9412,N_9553);
nor U10422 (N_10422,N_9716,N_9184);
or U10423 (N_10423,N_9099,N_9662);
xor U10424 (N_10424,N_9659,N_9550);
xor U10425 (N_10425,N_9082,N_9302);
xnor U10426 (N_10426,N_9157,N_9227);
nor U10427 (N_10427,N_9211,N_9107);
xor U10428 (N_10428,N_9388,N_9121);
nor U10429 (N_10429,N_9481,N_9454);
nand U10430 (N_10430,N_9139,N_9105);
nand U10431 (N_10431,N_9639,N_9681);
or U10432 (N_10432,N_9435,N_9267);
nand U10433 (N_10433,N_9864,N_9207);
nor U10434 (N_10434,N_9861,N_9595);
xor U10435 (N_10435,N_9369,N_9655);
nor U10436 (N_10436,N_9111,N_9455);
nor U10437 (N_10437,N_9313,N_9610);
or U10438 (N_10438,N_9636,N_9336);
or U10439 (N_10439,N_9914,N_9658);
xnor U10440 (N_10440,N_9237,N_9164);
xor U10441 (N_10441,N_9248,N_9835);
and U10442 (N_10442,N_9321,N_9011);
or U10443 (N_10443,N_9329,N_9287);
or U10444 (N_10444,N_9542,N_9300);
nor U10445 (N_10445,N_9999,N_9220);
xnor U10446 (N_10446,N_9095,N_9510);
nand U10447 (N_10447,N_9186,N_9185);
nand U10448 (N_10448,N_9376,N_9566);
nand U10449 (N_10449,N_9617,N_9744);
nor U10450 (N_10450,N_9770,N_9171);
nor U10451 (N_10451,N_9565,N_9968);
nand U10452 (N_10452,N_9020,N_9641);
nor U10453 (N_10453,N_9924,N_9262);
nor U10454 (N_10454,N_9528,N_9892);
nor U10455 (N_10455,N_9060,N_9419);
nor U10456 (N_10456,N_9384,N_9981);
and U10457 (N_10457,N_9347,N_9637);
xnor U10458 (N_10458,N_9044,N_9136);
nor U10459 (N_10459,N_9338,N_9727);
or U10460 (N_10460,N_9612,N_9922);
and U10461 (N_10461,N_9631,N_9822);
and U10462 (N_10462,N_9936,N_9377);
and U10463 (N_10463,N_9298,N_9401);
nand U10464 (N_10464,N_9063,N_9346);
nor U10465 (N_10465,N_9724,N_9524);
xor U10466 (N_10466,N_9705,N_9084);
xor U10467 (N_10467,N_9259,N_9019);
nand U10468 (N_10468,N_9373,N_9276);
and U10469 (N_10469,N_9643,N_9821);
nor U10470 (N_10470,N_9934,N_9832);
nand U10471 (N_10471,N_9911,N_9212);
and U10472 (N_10472,N_9810,N_9883);
nor U10473 (N_10473,N_9299,N_9325);
and U10474 (N_10474,N_9673,N_9490);
xnor U10475 (N_10475,N_9458,N_9882);
xnor U10476 (N_10476,N_9232,N_9326);
and U10477 (N_10477,N_9108,N_9008);
or U10478 (N_10478,N_9618,N_9918);
and U10479 (N_10479,N_9779,N_9794);
and U10480 (N_10480,N_9322,N_9679);
or U10481 (N_10481,N_9499,N_9189);
and U10482 (N_10482,N_9927,N_9221);
nor U10483 (N_10483,N_9578,N_9640);
or U10484 (N_10484,N_9803,N_9270);
nand U10485 (N_10485,N_9037,N_9796);
and U10486 (N_10486,N_9014,N_9693);
or U10487 (N_10487,N_9843,N_9077);
nor U10488 (N_10488,N_9795,N_9604);
nor U10489 (N_10489,N_9334,N_9272);
and U10490 (N_10490,N_9632,N_9620);
and U10491 (N_10491,N_9043,N_9798);
nand U10492 (N_10492,N_9386,N_9525);
and U10493 (N_10493,N_9012,N_9887);
and U10494 (N_10494,N_9932,N_9939);
and U10495 (N_10495,N_9411,N_9478);
nor U10496 (N_10496,N_9698,N_9030);
xor U10497 (N_10497,N_9176,N_9507);
nand U10498 (N_10498,N_9425,N_9182);
xnor U10499 (N_10499,N_9755,N_9434);
and U10500 (N_10500,N_9728,N_9742);
xnor U10501 (N_10501,N_9877,N_9723);
nand U10502 (N_10502,N_9381,N_9882);
nor U10503 (N_10503,N_9405,N_9606);
nand U10504 (N_10504,N_9586,N_9576);
nand U10505 (N_10505,N_9567,N_9987);
and U10506 (N_10506,N_9835,N_9527);
nor U10507 (N_10507,N_9754,N_9496);
nor U10508 (N_10508,N_9010,N_9760);
xnor U10509 (N_10509,N_9288,N_9665);
and U10510 (N_10510,N_9402,N_9055);
or U10511 (N_10511,N_9332,N_9115);
nor U10512 (N_10512,N_9965,N_9653);
and U10513 (N_10513,N_9060,N_9769);
xnor U10514 (N_10514,N_9318,N_9870);
xor U10515 (N_10515,N_9267,N_9655);
nand U10516 (N_10516,N_9370,N_9312);
or U10517 (N_10517,N_9671,N_9907);
xor U10518 (N_10518,N_9702,N_9127);
nand U10519 (N_10519,N_9343,N_9132);
nor U10520 (N_10520,N_9727,N_9948);
xor U10521 (N_10521,N_9545,N_9071);
nand U10522 (N_10522,N_9242,N_9877);
xor U10523 (N_10523,N_9175,N_9287);
nand U10524 (N_10524,N_9833,N_9038);
nor U10525 (N_10525,N_9445,N_9824);
nand U10526 (N_10526,N_9655,N_9763);
nand U10527 (N_10527,N_9505,N_9256);
xor U10528 (N_10528,N_9442,N_9451);
or U10529 (N_10529,N_9173,N_9162);
nand U10530 (N_10530,N_9940,N_9639);
or U10531 (N_10531,N_9759,N_9967);
nand U10532 (N_10532,N_9315,N_9826);
nor U10533 (N_10533,N_9482,N_9032);
nand U10534 (N_10534,N_9701,N_9474);
or U10535 (N_10535,N_9831,N_9330);
nor U10536 (N_10536,N_9663,N_9621);
nor U10537 (N_10537,N_9513,N_9873);
nand U10538 (N_10538,N_9079,N_9632);
nand U10539 (N_10539,N_9975,N_9635);
and U10540 (N_10540,N_9596,N_9515);
or U10541 (N_10541,N_9992,N_9592);
nor U10542 (N_10542,N_9849,N_9129);
xor U10543 (N_10543,N_9373,N_9539);
nor U10544 (N_10544,N_9331,N_9361);
or U10545 (N_10545,N_9185,N_9684);
and U10546 (N_10546,N_9541,N_9189);
and U10547 (N_10547,N_9593,N_9247);
nand U10548 (N_10548,N_9993,N_9789);
nand U10549 (N_10549,N_9964,N_9347);
nand U10550 (N_10550,N_9842,N_9402);
or U10551 (N_10551,N_9706,N_9533);
nand U10552 (N_10552,N_9792,N_9139);
xor U10553 (N_10553,N_9139,N_9020);
nor U10554 (N_10554,N_9729,N_9346);
xor U10555 (N_10555,N_9495,N_9021);
xnor U10556 (N_10556,N_9183,N_9303);
or U10557 (N_10557,N_9638,N_9940);
nand U10558 (N_10558,N_9842,N_9568);
xor U10559 (N_10559,N_9487,N_9523);
or U10560 (N_10560,N_9374,N_9592);
xor U10561 (N_10561,N_9147,N_9724);
xor U10562 (N_10562,N_9954,N_9447);
or U10563 (N_10563,N_9228,N_9360);
and U10564 (N_10564,N_9066,N_9664);
and U10565 (N_10565,N_9464,N_9013);
or U10566 (N_10566,N_9877,N_9994);
xor U10567 (N_10567,N_9351,N_9860);
and U10568 (N_10568,N_9320,N_9659);
nor U10569 (N_10569,N_9614,N_9207);
or U10570 (N_10570,N_9844,N_9886);
xor U10571 (N_10571,N_9624,N_9418);
or U10572 (N_10572,N_9960,N_9061);
nand U10573 (N_10573,N_9210,N_9303);
nand U10574 (N_10574,N_9515,N_9062);
nor U10575 (N_10575,N_9442,N_9660);
and U10576 (N_10576,N_9580,N_9192);
or U10577 (N_10577,N_9414,N_9112);
nor U10578 (N_10578,N_9669,N_9240);
or U10579 (N_10579,N_9422,N_9779);
nand U10580 (N_10580,N_9029,N_9335);
or U10581 (N_10581,N_9919,N_9485);
xnor U10582 (N_10582,N_9082,N_9508);
nor U10583 (N_10583,N_9095,N_9270);
or U10584 (N_10584,N_9296,N_9756);
and U10585 (N_10585,N_9331,N_9815);
nand U10586 (N_10586,N_9611,N_9866);
nand U10587 (N_10587,N_9805,N_9064);
and U10588 (N_10588,N_9258,N_9761);
and U10589 (N_10589,N_9550,N_9939);
or U10590 (N_10590,N_9605,N_9851);
and U10591 (N_10591,N_9527,N_9661);
xor U10592 (N_10592,N_9594,N_9831);
and U10593 (N_10593,N_9159,N_9750);
nand U10594 (N_10594,N_9010,N_9845);
xor U10595 (N_10595,N_9139,N_9635);
and U10596 (N_10596,N_9091,N_9400);
or U10597 (N_10597,N_9738,N_9196);
nor U10598 (N_10598,N_9669,N_9220);
nand U10599 (N_10599,N_9535,N_9277);
xor U10600 (N_10600,N_9710,N_9737);
xor U10601 (N_10601,N_9297,N_9652);
and U10602 (N_10602,N_9077,N_9343);
nand U10603 (N_10603,N_9802,N_9075);
and U10604 (N_10604,N_9190,N_9367);
xor U10605 (N_10605,N_9218,N_9067);
and U10606 (N_10606,N_9149,N_9469);
nand U10607 (N_10607,N_9465,N_9673);
and U10608 (N_10608,N_9039,N_9521);
and U10609 (N_10609,N_9073,N_9462);
nor U10610 (N_10610,N_9193,N_9100);
or U10611 (N_10611,N_9666,N_9875);
or U10612 (N_10612,N_9118,N_9639);
or U10613 (N_10613,N_9593,N_9389);
xor U10614 (N_10614,N_9435,N_9203);
and U10615 (N_10615,N_9165,N_9287);
or U10616 (N_10616,N_9760,N_9281);
nor U10617 (N_10617,N_9027,N_9849);
nor U10618 (N_10618,N_9177,N_9845);
nor U10619 (N_10619,N_9980,N_9552);
nor U10620 (N_10620,N_9290,N_9183);
nand U10621 (N_10621,N_9618,N_9847);
nor U10622 (N_10622,N_9044,N_9279);
nand U10623 (N_10623,N_9116,N_9962);
xnor U10624 (N_10624,N_9322,N_9512);
nor U10625 (N_10625,N_9133,N_9212);
xor U10626 (N_10626,N_9405,N_9609);
xor U10627 (N_10627,N_9649,N_9857);
and U10628 (N_10628,N_9011,N_9024);
xnor U10629 (N_10629,N_9467,N_9983);
xor U10630 (N_10630,N_9715,N_9438);
xor U10631 (N_10631,N_9528,N_9264);
nor U10632 (N_10632,N_9136,N_9795);
xnor U10633 (N_10633,N_9885,N_9921);
nand U10634 (N_10634,N_9385,N_9270);
nor U10635 (N_10635,N_9256,N_9236);
nor U10636 (N_10636,N_9940,N_9136);
nor U10637 (N_10637,N_9272,N_9049);
nand U10638 (N_10638,N_9636,N_9390);
xor U10639 (N_10639,N_9562,N_9508);
xnor U10640 (N_10640,N_9661,N_9581);
xnor U10641 (N_10641,N_9183,N_9739);
or U10642 (N_10642,N_9750,N_9790);
or U10643 (N_10643,N_9923,N_9831);
and U10644 (N_10644,N_9860,N_9073);
xnor U10645 (N_10645,N_9984,N_9650);
or U10646 (N_10646,N_9494,N_9179);
and U10647 (N_10647,N_9204,N_9419);
or U10648 (N_10648,N_9867,N_9045);
xnor U10649 (N_10649,N_9344,N_9494);
and U10650 (N_10650,N_9206,N_9388);
and U10651 (N_10651,N_9905,N_9173);
nor U10652 (N_10652,N_9567,N_9167);
nor U10653 (N_10653,N_9518,N_9666);
xnor U10654 (N_10654,N_9268,N_9894);
or U10655 (N_10655,N_9116,N_9439);
or U10656 (N_10656,N_9879,N_9960);
or U10657 (N_10657,N_9289,N_9844);
xnor U10658 (N_10658,N_9195,N_9992);
or U10659 (N_10659,N_9724,N_9651);
or U10660 (N_10660,N_9994,N_9860);
nand U10661 (N_10661,N_9667,N_9630);
nand U10662 (N_10662,N_9664,N_9494);
xnor U10663 (N_10663,N_9913,N_9052);
nand U10664 (N_10664,N_9669,N_9786);
or U10665 (N_10665,N_9106,N_9856);
xnor U10666 (N_10666,N_9926,N_9887);
or U10667 (N_10667,N_9391,N_9564);
nor U10668 (N_10668,N_9232,N_9104);
xnor U10669 (N_10669,N_9316,N_9921);
or U10670 (N_10670,N_9152,N_9499);
xor U10671 (N_10671,N_9568,N_9986);
xnor U10672 (N_10672,N_9925,N_9598);
xnor U10673 (N_10673,N_9069,N_9563);
nand U10674 (N_10674,N_9166,N_9785);
nand U10675 (N_10675,N_9200,N_9986);
xor U10676 (N_10676,N_9747,N_9915);
nor U10677 (N_10677,N_9269,N_9287);
and U10678 (N_10678,N_9705,N_9462);
nor U10679 (N_10679,N_9242,N_9281);
and U10680 (N_10680,N_9494,N_9731);
or U10681 (N_10681,N_9904,N_9621);
nor U10682 (N_10682,N_9887,N_9812);
xnor U10683 (N_10683,N_9686,N_9018);
or U10684 (N_10684,N_9834,N_9913);
and U10685 (N_10685,N_9383,N_9061);
or U10686 (N_10686,N_9124,N_9175);
and U10687 (N_10687,N_9112,N_9389);
nand U10688 (N_10688,N_9945,N_9677);
and U10689 (N_10689,N_9579,N_9400);
xor U10690 (N_10690,N_9517,N_9462);
nor U10691 (N_10691,N_9820,N_9950);
xor U10692 (N_10692,N_9148,N_9084);
nor U10693 (N_10693,N_9737,N_9624);
or U10694 (N_10694,N_9433,N_9298);
nor U10695 (N_10695,N_9569,N_9743);
and U10696 (N_10696,N_9003,N_9122);
and U10697 (N_10697,N_9117,N_9863);
nor U10698 (N_10698,N_9153,N_9600);
nor U10699 (N_10699,N_9939,N_9673);
nand U10700 (N_10700,N_9443,N_9407);
nor U10701 (N_10701,N_9570,N_9243);
or U10702 (N_10702,N_9700,N_9052);
and U10703 (N_10703,N_9912,N_9655);
or U10704 (N_10704,N_9999,N_9229);
nor U10705 (N_10705,N_9138,N_9230);
xnor U10706 (N_10706,N_9051,N_9141);
nor U10707 (N_10707,N_9035,N_9977);
or U10708 (N_10708,N_9329,N_9839);
or U10709 (N_10709,N_9383,N_9001);
xor U10710 (N_10710,N_9817,N_9368);
or U10711 (N_10711,N_9763,N_9799);
and U10712 (N_10712,N_9553,N_9098);
nor U10713 (N_10713,N_9847,N_9165);
nand U10714 (N_10714,N_9223,N_9837);
and U10715 (N_10715,N_9505,N_9946);
or U10716 (N_10716,N_9697,N_9882);
or U10717 (N_10717,N_9442,N_9044);
and U10718 (N_10718,N_9470,N_9463);
or U10719 (N_10719,N_9591,N_9779);
nor U10720 (N_10720,N_9092,N_9977);
and U10721 (N_10721,N_9253,N_9196);
and U10722 (N_10722,N_9569,N_9888);
nand U10723 (N_10723,N_9563,N_9077);
nand U10724 (N_10724,N_9684,N_9795);
nand U10725 (N_10725,N_9570,N_9113);
and U10726 (N_10726,N_9274,N_9248);
or U10727 (N_10727,N_9097,N_9491);
and U10728 (N_10728,N_9050,N_9270);
and U10729 (N_10729,N_9616,N_9277);
nand U10730 (N_10730,N_9351,N_9567);
nor U10731 (N_10731,N_9146,N_9719);
nand U10732 (N_10732,N_9990,N_9624);
and U10733 (N_10733,N_9397,N_9027);
or U10734 (N_10734,N_9228,N_9230);
xnor U10735 (N_10735,N_9355,N_9453);
nor U10736 (N_10736,N_9804,N_9622);
and U10737 (N_10737,N_9359,N_9988);
nor U10738 (N_10738,N_9989,N_9604);
or U10739 (N_10739,N_9077,N_9558);
or U10740 (N_10740,N_9624,N_9671);
nor U10741 (N_10741,N_9107,N_9138);
or U10742 (N_10742,N_9330,N_9207);
xor U10743 (N_10743,N_9276,N_9043);
nor U10744 (N_10744,N_9650,N_9982);
nor U10745 (N_10745,N_9848,N_9745);
nand U10746 (N_10746,N_9656,N_9513);
xor U10747 (N_10747,N_9360,N_9271);
and U10748 (N_10748,N_9795,N_9750);
nand U10749 (N_10749,N_9598,N_9632);
and U10750 (N_10750,N_9728,N_9081);
nand U10751 (N_10751,N_9914,N_9105);
or U10752 (N_10752,N_9457,N_9868);
nand U10753 (N_10753,N_9566,N_9782);
nor U10754 (N_10754,N_9315,N_9292);
nor U10755 (N_10755,N_9853,N_9055);
and U10756 (N_10756,N_9230,N_9126);
nor U10757 (N_10757,N_9937,N_9123);
or U10758 (N_10758,N_9519,N_9365);
nor U10759 (N_10759,N_9733,N_9598);
xor U10760 (N_10760,N_9550,N_9206);
nand U10761 (N_10761,N_9340,N_9652);
nor U10762 (N_10762,N_9871,N_9881);
xnor U10763 (N_10763,N_9393,N_9641);
or U10764 (N_10764,N_9590,N_9124);
xor U10765 (N_10765,N_9631,N_9851);
and U10766 (N_10766,N_9207,N_9694);
xnor U10767 (N_10767,N_9011,N_9876);
xnor U10768 (N_10768,N_9206,N_9974);
nor U10769 (N_10769,N_9322,N_9003);
xnor U10770 (N_10770,N_9332,N_9540);
xnor U10771 (N_10771,N_9481,N_9717);
xnor U10772 (N_10772,N_9261,N_9338);
nor U10773 (N_10773,N_9227,N_9886);
and U10774 (N_10774,N_9369,N_9763);
xor U10775 (N_10775,N_9007,N_9237);
xor U10776 (N_10776,N_9471,N_9359);
xor U10777 (N_10777,N_9077,N_9791);
nor U10778 (N_10778,N_9029,N_9022);
and U10779 (N_10779,N_9347,N_9044);
or U10780 (N_10780,N_9957,N_9275);
and U10781 (N_10781,N_9119,N_9007);
and U10782 (N_10782,N_9710,N_9487);
or U10783 (N_10783,N_9270,N_9646);
and U10784 (N_10784,N_9997,N_9248);
or U10785 (N_10785,N_9056,N_9984);
or U10786 (N_10786,N_9335,N_9988);
or U10787 (N_10787,N_9335,N_9098);
and U10788 (N_10788,N_9201,N_9509);
nand U10789 (N_10789,N_9676,N_9033);
or U10790 (N_10790,N_9764,N_9964);
nand U10791 (N_10791,N_9239,N_9629);
or U10792 (N_10792,N_9228,N_9344);
and U10793 (N_10793,N_9404,N_9905);
nor U10794 (N_10794,N_9607,N_9582);
nor U10795 (N_10795,N_9836,N_9283);
xnor U10796 (N_10796,N_9490,N_9519);
xor U10797 (N_10797,N_9469,N_9209);
nand U10798 (N_10798,N_9016,N_9655);
xnor U10799 (N_10799,N_9099,N_9912);
xnor U10800 (N_10800,N_9738,N_9510);
xor U10801 (N_10801,N_9978,N_9847);
or U10802 (N_10802,N_9249,N_9490);
nand U10803 (N_10803,N_9519,N_9699);
or U10804 (N_10804,N_9861,N_9891);
and U10805 (N_10805,N_9524,N_9219);
xnor U10806 (N_10806,N_9746,N_9762);
xnor U10807 (N_10807,N_9777,N_9069);
and U10808 (N_10808,N_9300,N_9124);
xnor U10809 (N_10809,N_9262,N_9116);
nor U10810 (N_10810,N_9030,N_9756);
nor U10811 (N_10811,N_9183,N_9709);
and U10812 (N_10812,N_9336,N_9018);
nand U10813 (N_10813,N_9907,N_9950);
and U10814 (N_10814,N_9212,N_9606);
nor U10815 (N_10815,N_9365,N_9324);
xnor U10816 (N_10816,N_9135,N_9971);
xnor U10817 (N_10817,N_9450,N_9935);
and U10818 (N_10818,N_9526,N_9008);
xnor U10819 (N_10819,N_9888,N_9428);
and U10820 (N_10820,N_9784,N_9261);
xor U10821 (N_10821,N_9404,N_9598);
xor U10822 (N_10822,N_9606,N_9940);
and U10823 (N_10823,N_9114,N_9451);
or U10824 (N_10824,N_9943,N_9166);
nor U10825 (N_10825,N_9413,N_9949);
xor U10826 (N_10826,N_9949,N_9381);
or U10827 (N_10827,N_9208,N_9464);
and U10828 (N_10828,N_9240,N_9296);
or U10829 (N_10829,N_9622,N_9730);
xor U10830 (N_10830,N_9880,N_9481);
and U10831 (N_10831,N_9362,N_9854);
xor U10832 (N_10832,N_9391,N_9717);
nor U10833 (N_10833,N_9913,N_9506);
nand U10834 (N_10834,N_9719,N_9560);
nand U10835 (N_10835,N_9097,N_9198);
or U10836 (N_10836,N_9804,N_9290);
and U10837 (N_10837,N_9581,N_9705);
nand U10838 (N_10838,N_9887,N_9654);
nor U10839 (N_10839,N_9851,N_9936);
and U10840 (N_10840,N_9116,N_9644);
and U10841 (N_10841,N_9103,N_9313);
xnor U10842 (N_10842,N_9247,N_9462);
and U10843 (N_10843,N_9832,N_9082);
and U10844 (N_10844,N_9289,N_9168);
or U10845 (N_10845,N_9160,N_9525);
or U10846 (N_10846,N_9279,N_9664);
and U10847 (N_10847,N_9912,N_9446);
nand U10848 (N_10848,N_9138,N_9367);
or U10849 (N_10849,N_9252,N_9226);
nand U10850 (N_10850,N_9107,N_9309);
or U10851 (N_10851,N_9086,N_9859);
nor U10852 (N_10852,N_9000,N_9365);
nand U10853 (N_10853,N_9728,N_9879);
nand U10854 (N_10854,N_9886,N_9708);
or U10855 (N_10855,N_9732,N_9511);
or U10856 (N_10856,N_9767,N_9757);
xnor U10857 (N_10857,N_9816,N_9672);
and U10858 (N_10858,N_9763,N_9301);
nor U10859 (N_10859,N_9723,N_9026);
xor U10860 (N_10860,N_9532,N_9951);
xnor U10861 (N_10861,N_9438,N_9705);
and U10862 (N_10862,N_9225,N_9784);
nor U10863 (N_10863,N_9334,N_9253);
or U10864 (N_10864,N_9137,N_9608);
and U10865 (N_10865,N_9539,N_9406);
nand U10866 (N_10866,N_9805,N_9178);
or U10867 (N_10867,N_9111,N_9103);
nand U10868 (N_10868,N_9523,N_9365);
nand U10869 (N_10869,N_9608,N_9291);
xor U10870 (N_10870,N_9938,N_9679);
nor U10871 (N_10871,N_9135,N_9449);
and U10872 (N_10872,N_9341,N_9079);
xor U10873 (N_10873,N_9500,N_9077);
xnor U10874 (N_10874,N_9885,N_9986);
or U10875 (N_10875,N_9861,N_9813);
nand U10876 (N_10876,N_9601,N_9902);
xor U10877 (N_10877,N_9223,N_9270);
xor U10878 (N_10878,N_9179,N_9588);
xor U10879 (N_10879,N_9566,N_9595);
xnor U10880 (N_10880,N_9392,N_9447);
xnor U10881 (N_10881,N_9401,N_9933);
or U10882 (N_10882,N_9388,N_9603);
xnor U10883 (N_10883,N_9941,N_9290);
xnor U10884 (N_10884,N_9883,N_9554);
nand U10885 (N_10885,N_9563,N_9978);
nor U10886 (N_10886,N_9965,N_9676);
nand U10887 (N_10887,N_9601,N_9523);
nand U10888 (N_10888,N_9716,N_9288);
and U10889 (N_10889,N_9054,N_9194);
and U10890 (N_10890,N_9960,N_9008);
and U10891 (N_10891,N_9818,N_9264);
or U10892 (N_10892,N_9820,N_9322);
nor U10893 (N_10893,N_9468,N_9675);
nand U10894 (N_10894,N_9181,N_9021);
or U10895 (N_10895,N_9747,N_9771);
or U10896 (N_10896,N_9602,N_9068);
or U10897 (N_10897,N_9534,N_9471);
xor U10898 (N_10898,N_9705,N_9608);
xnor U10899 (N_10899,N_9990,N_9823);
or U10900 (N_10900,N_9004,N_9569);
nand U10901 (N_10901,N_9922,N_9030);
and U10902 (N_10902,N_9223,N_9822);
xor U10903 (N_10903,N_9306,N_9060);
xnor U10904 (N_10904,N_9349,N_9631);
nand U10905 (N_10905,N_9612,N_9919);
and U10906 (N_10906,N_9244,N_9690);
xor U10907 (N_10907,N_9847,N_9215);
or U10908 (N_10908,N_9118,N_9771);
or U10909 (N_10909,N_9906,N_9803);
nand U10910 (N_10910,N_9576,N_9447);
or U10911 (N_10911,N_9669,N_9491);
nor U10912 (N_10912,N_9971,N_9023);
and U10913 (N_10913,N_9604,N_9307);
xor U10914 (N_10914,N_9170,N_9068);
nor U10915 (N_10915,N_9550,N_9627);
xnor U10916 (N_10916,N_9685,N_9939);
nor U10917 (N_10917,N_9711,N_9482);
nor U10918 (N_10918,N_9488,N_9135);
nor U10919 (N_10919,N_9055,N_9601);
and U10920 (N_10920,N_9233,N_9197);
nand U10921 (N_10921,N_9864,N_9309);
xnor U10922 (N_10922,N_9479,N_9352);
and U10923 (N_10923,N_9053,N_9642);
xor U10924 (N_10924,N_9340,N_9689);
nand U10925 (N_10925,N_9557,N_9724);
xnor U10926 (N_10926,N_9601,N_9677);
nand U10927 (N_10927,N_9690,N_9654);
nand U10928 (N_10928,N_9536,N_9143);
or U10929 (N_10929,N_9550,N_9997);
nand U10930 (N_10930,N_9028,N_9846);
xor U10931 (N_10931,N_9234,N_9146);
or U10932 (N_10932,N_9008,N_9761);
xnor U10933 (N_10933,N_9973,N_9249);
and U10934 (N_10934,N_9062,N_9944);
xor U10935 (N_10935,N_9269,N_9378);
and U10936 (N_10936,N_9445,N_9275);
and U10937 (N_10937,N_9130,N_9762);
and U10938 (N_10938,N_9524,N_9747);
nor U10939 (N_10939,N_9547,N_9327);
nor U10940 (N_10940,N_9576,N_9559);
nand U10941 (N_10941,N_9618,N_9795);
nand U10942 (N_10942,N_9372,N_9711);
and U10943 (N_10943,N_9985,N_9503);
nor U10944 (N_10944,N_9669,N_9417);
or U10945 (N_10945,N_9370,N_9150);
xor U10946 (N_10946,N_9241,N_9626);
nand U10947 (N_10947,N_9964,N_9573);
nor U10948 (N_10948,N_9736,N_9745);
and U10949 (N_10949,N_9080,N_9666);
or U10950 (N_10950,N_9413,N_9241);
nand U10951 (N_10951,N_9038,N_9730);
nand U10952 (N_10952,N_9397,N_9322);
xnor U10953 (N_10953,N_9436,N_9202);
nor U10954 (N_10954,N_9257,N_9628);
or U10955 (N_10955,N_9233,N_9331);
nor U10956 (N_10956,N_9363,N_9584);
or U10957 (N_10957,N_9006,N_9172);
and U10958 (N_10958,N_9342,N_9150);
and U10959 (N_10959,N_9004,N_9003);
nand U10960 (N_10960,N_9890,N_9885);
or U10961 (N_10961,N_9313,N_9336);
or U10962 (N_10962,N_9456,N_9496);
nor U10963 (N_10963,N_9943,N_9088);
nor U10964 (N_10964,N_9332,N_9457);
nand U10965 (N_10965,N_9047,N_9784);
xnor U10966 (N_10966,N_9972,N_9719);
or U10967 (N_10967,N_9400,N_9698);
xnor U10968 (N_10968,N_9552,N_9202);
xnor U10969 (N_10969,N_9911,N_9774);
nor U10970 (N_10970,N_9777,N_9684);
and U10971 (N_10971,N_9447,N_9838);
or U10972 (N_10972,N_9623,N_9050);
nand U10973 (N_10973,N_9997,N_9390);
and U10974 (N_10974,N_9701,N_9230);
nand U10975 (N_10975,N_9405,N_9345);
and U10976 (N_10976,N_9742,N_9387);
xor U10977 (N_10977,N_9098,N_9154);
nor U10978 (N_10978,N_9556,N_9439);
or U10979 (N_10979,N_9678,N_9333);
and U10980 (N_10980,N_9321,N_9783);
or U10981 (N_10981,N_9742,N_9493);
nor U10982 (N_10982,N_9175,N_9129);
nand U10983 (N_10983,N_9089,N_9504);
xor U10984 (N_10984,N_9897,N_9294);
and U10985 (N_10985,N_9222,N_9335);
nand U10986 (N_10986,N_9286,N_9838);
and U10987 (N_10987,N_9726,N_9688);
or U10988 (N_10988,N_9422,N_9687);
or U10989 (N_10989,N_9789,N_9588);
nor U10990 (N_10990,N_9480,N_9273);
nand U10991 (N_10991,N_9505,N_9184);
xnor U10992 (N_10992,N_9357,N_9880);
or U10993 (N_10993,N_9149,N_9733);
nand U10994 (N_10994,N_9790,N_9170);
nor U10995 (N_10995,N_9430,N_9491);
nor U10996 (N_10996,N_9653,N_9261);
or U10997 (N_10997,N_9856,N_9099);
nor U10998 (N_10998,N_9448,N_9424);
and U10999 (N_10999,N_9653,N_9086);
nor U11000 (N_11000,N_10439,N_10604);
xnor U11001 (N_11001,N_10412,N_10758);
nor U11002 (N_11002,N_10383,N_10969);
xor U11003 (N_11003,N_10314,N_10180);
nand U11004 (N_11004,N_10676,N_10086);
nand U11005 (N_11005,N_10992,N_10560);
nor U11006 (N_11006,N_10428,N_10380);
nor U11007 (N_11007,N_10612,N_10082);
xnor U11008 (N_11008,N_10952,N_10065);
or U11009 (N_11009,N_10799,N_10983);
xnor U11010 (N_11010,N_10045,N_10092);
and U11011 (N_11011,N_10597,N_10582);
nor U11012 (N_11012,N_10779,N_10066);
and U11013 (N_11013,N_10624,N_10694);
and U11014 (N_11014,N_10640,N_10410);
or U11015 (N_11015,N_10498,N_10618);
or U11016 (N_11016,N_10042,N_10685);
or U11017 (N_11017,N_10321,N_10932);
nor U11018 (N_11018,N_10921,N_10872);
xnor U11019 (N_11019,N_10525,N_10474);
xor U11020 (N_11020,N_10977,N_10368);
nand U11021 (N_11021,N_10577,N_10129);
or U11022 (N_11022,N_10344,N_10654);
or U11023 (N_11023,N_10530,N_10208);
nor U11024 (N_11024,N_10851,N_10834);
and U11025 (N_11025,N_10709,N_10285);
or U11026 (N_11026,N_10827,N_10449);
nor U11027 (N_11027,N_10912,N_10088);
nand U11028 (N_11028,N_10081,N_10602);
xnor U11029 (N_11029,N_10935,N_10950);
and U11030 (N_11030,N_10219,N_10537);
xor U11031 (N_11031,N_10951,N_10480);
xor U11032 (N_11032,N_10677,N_10581);
xnor U11033 (N_11033,N_10293,N_10179);
or U11034 (N_11034,N_10578,N_10083);
nor U11035 (N_11035,N_10854,N_10810);
nor U11036 (N_11036,N_10615,N_10980);
xor U11037 (N_11037,N_10975,N_10069);
or U11038 (N_11038,N_10242,N_10524);
xnor U11039 (N_11039,N_10215,N_10232);
or U11040 (N_11040,N_10097,N_10998);
xnor U11041 (N_11041,N_10073,N_10135);
nand U11042 (N_11042,N_10606,N_10011);
nor U11043 (N_11043,N_10408,N_10771);
nand U11044 (N_11044,N_10649,N_10448);
nand U11045 (N_11045,N_10387,N_10189);
nor U11046 (N_11046,N_10866,N_10101);
nor U11047 (N_11047,N_10322,N_10005);
nor U11048 (N_11048,N_10887,N_10468);
xnor U11049 (N_11049,N_10460,N_10919);
xnor U11050 (N_11050,N_10857,N_10328);
xor U11051 (N_11051,N_10148,N_10643);
nand U11052 (N_11052,N_10305,N_10499);
and U11053 (N_11053,N_10304,N_10164);
nor U11054 (N_11054,N_10890,N_10197);
xnor U11055 (N_11055,N_10588,N_10868);
nor U11056 (N_11056,N_10829,N_10382);
nand U11057 (N_11057,N_10120,N_10263);
nor U11058 (N_11058,N_10715,N_10220);
nor U11059 (N_11059,N_10331,N_10905);
xor U11060 (N_11060,N_10748,N_10824);
nand U11061 (N_11061,N_10021,N_10355);
and U11062 (N_11062,N_10347,N_10006);
nor U11063 (N_11063,N_10586,N_10417);
and U11064 (N_11064,N_10497,N_10707);
nand U11065 (N_11065,N_10405,N_10451);
or U11066 (N_11066,N_10716,N_10636);
nand U11067 (N_11067,N_10348,N_10956);
and U11068 (N_11068,N_10399,N_10031);
nand U11069 (N_11069,N_10398,N_10822);
nor U11070 (N_11070,N_10652,N_10443);
or U11071 (N_11071,N_10634,N_10161);
xor U11072 (N_11072,N_10297,N_10972);
nor U11073 (N_11073,N_10240,N_10349);
xnor U11074 (N_11074,N_10703,N_10472);
nor U11075 (N_11075,N_10697,N_10743);
nor U11076 (N_11076,N_10084,N_10378);
nand U11077 (N_11077,N_10999,N_10358);
nor U11078 (N_11078,N_10024,N_10646);
xnor U11079 (N_11079,N_10218,N_10450);
or U11080 (N_11080,N_10641,N_10736);
nand U11081 (N_11081,N_10807,N_10249);
and U11082 (N_11082,N_10510,N_10243);
and U11083 (N_11083,N_10786,N_10264);
nand U11084 (N_11084,N_10223,N_10632);
or U11085 (N_11085,N_10713,N_10843);
xnor U11086 (N_11086,N_10416,N_10421);
nand U11087 (N_11087,N_10257,N_10711);
nor U11088 (N_11088,N_10205,N_10067);
or U11089 (N_11089,N_10267,N_10727);
nor U11090 (N_11090,N_10766,N_10914);
xor U11091 (N_11091,N_10605,N_10596);
nand U11092 (N_11092,N_10201,N_10216);
or U11093 (N_11093,N_10751,N_10491);
nor U11094 (N_11094,N_10192,N_10319);
nand U11095 (N_11095,N_10049,N_10522);
and U11096 (N_11096,N_10052,N_10268);
nor U11097 (N_11097,N_10313,N_10246);
xnor U11098 (N_11098,N_10139,N_10486);
nor U11099 (N_11099,N_10995,N_10623);
xor U11100 (N_11100,N_10169,N_10312);
nor U11101 (N_11101,N_10241,N_10206);
nand U11102 (N_11102,N_10761,N_10942);
or U11103 (N_11103,N_10365,N_10885);
xor U11104 (N_11104,N_10104,N_10102);
nand U11105 (N_11105,N_10376,N_10362);
nand U11106 (N_11106,N_10311,N_10533);
and U11107 (N_11107,N_10424,N_10106);
nor U11108 (N_11108,N_10431,N_10607);
or U11109 (N_11109,N_10819,N_10704);
xor U11110 (N_11110,N_10603,N_10238);
nand U11111 (N_11111,N_10453,N_10515);
nand U11112 (N_11112,N_10444,N_10258);
xor U11113 (N_11113,N_10611,N_10846);
nor U11114 (N_11114,N_10070,N_10513);
or U11115 (N_11115,N_10411,N_10361);
and U11116 (N_11116,N_10911,N_10369);
and U11117 (N_11117,N_10837,N_10260);
nor U11118 (N_11118,N_10392,N_10274);
or U11119 (N_11119,N_10823,N_10543);
and U11120 (N_11120,N_10955,N_10842);
and U11121 (N_11121,N_10953,N_10063);
nand U11122 (N_11122,N_10630,N_10136);
xor U11123 (N_11123,N_10883,N_10683);
nor U11124 (N_11124,N_10419,N_10173);
xor U11125 (N_11125,N_10592,N_10788);
xnor U11126 (N_11126,N_10898,N_10360);
and U11127 (N_11127,N_10200,N_10796);
or U11128 (N_11128,N_10036,N_10818);
or U11129 (N_11129,N_10617,N_10891);
or U11130 (N_11130,N_10939,N_10534);
nor U11131 (N_11131,N_10740,N_10339);
and U11132 (N_11132,N_10813,N_10318);
xnor U11133 (N_11133,N_10627,N_10295);
or U11134 (N_11134,N_10859,N_10458);
xnor U11135 (N_11135,N_10541,N_10591);
and U11136 (N_11136,N_10307,N_10839);
xnor U11137 (N_11137,N_10023,N_10565);
or U11138 (N_11138,N_10929,N_10255);
or U11139 (N_11139,N_10462,N_10688);
and U11140 (N_11140,N_10874,N_10126);
xnor U11141 (N_11141,N_10769,N_10504);
or U11142 (N_11142,N_10664,N_10809);
nand U11143 (N_11143,N_10131,N_10356);
nand U11144 (N_11144,N_10876,N_10107);
and U11145 (N_11145,N_10217,N_10836);
nand U11146 (N_11146,N_10281,N_10529);
and U11147 (N_11147,N_10714,N_10384);
nor U11148 (N_11148,N_10115,N_10946);
nand U11149 (N_11149,N_10732,N_10210);
nor U11150 (N_11150,N_10826,N_10695);
or U11151 (N_11151,N_10767,N_10559);
and U11152 (N_11152,N_10787,N_10614);
xnor U11153 (N_11153,N_10982,N_10375);
nand U11154 (N_11154,N_10712,N_10168);
and U11155 (N_11155,N_10792,N_10095);
nor U11156 (N_11156,N_10269,N_10841);
or U11157 (N_11157,N_10968,N_10233);
xor U11158 (N_11158,N_10401,N_10390);
nand U11159 (N_11159,N_10579,N_10265);
nor U11160 (N_11160,N_10108,N_10090);
nand U11161 (N_11161,N_10734,N_10058);
nand U11162 (N_11162,N_10487,N_10973);
xnor U11163 (N_11163,N_10985,N_10686);
nand U11164 (N_11164,N_10760,N_10296);
nand U11165 (N_11165,N_10237,N_10888);
nor U11166 (N_11166,N_10064,N_10178);
xor U11167 (N_11167,N_10132,N_10454);
xor U11168 (N_11168,N_10961,N_10523);
xnor U11169 (N_11169,N_10072,N_10802);
or U11170 (N_11170,N_10418,N_10558);
or U11171 (N_11171,N_10004,N_10464);
or U11172 (N_11172,N_10554,N_10954);
nand U11173 (N_11173,N_10330,N_10445);
and U11174 (N_11174,N_10928,N_10367);
nand U11175 (N_11175,N_10655,N_10414);
nand U11176 (N_11176,N_10186,N_10459);
nor U11177 (N_11177,N_10693,N_10144);
nor U11178 (N_11178,N_10409,N_10395);
xnor U11179 (N_11179,N_10724,N_10551);
and U11180 (N_11180,N_10167,N_10133);
nand U11181 (N_11181,N_10001,N_10811);
nand U11182 (N_11182,N_10284,N_10680);
nor U11183 (N_11183,N_10645,N_10035);
and U11184 (N_11184,N_10061,N_10849);
nand U11185 (N_11185,N_10053,N_10234);
and U11186 (N_11186,N_10231,N_10723);
or U11187 (N_11187,N_10508,N_10987);
or U11188 (N_11188,N_10917,N_10739);
or U11189 (N_11189,N_10032,N_10926);
nand U11190 (N_11190,N_10209,N_10698);
xor U11191 (N_11191,N_10770,N_10960);
and U11192 (N_11192,N_10119,N_10177);
xnor U11193 (N_11193,N_10324,N_10589);
xnor U11194 (N_11194,N_10991,N_10741);
nor U11195 (N_11195,N_10043,N_10622);
nor U11196 (N_11196,N_10286,N_10496);
xor U11197 (N_11197,N_10722,N_10549);
nor U11198 (N_11198,N_10039,N_10316);
nor U11199 (N_11199,N_10336,N_10153);
xnor U11200 (N_11200,N_10423,N_10665);
xor U11201 (N_11201,N_10520,N_10909);
or U11202 (N_11202,N_10661,N_10765);
and U11203 (N_11203,N_10374,N_10400);
nand U11204 (N_11204,N_10923,N_10310);
or U11205 (N_11205,N_10145,N_10521);
xnor U11206 (N_11206,N_10396,N_10574);
or U11207 (N_11207,N_10143,N_10294);
or U11208 (N_11208,N_10718,N_10130);
nand U11209 (N_11209,N_10873,N_10762);
or U11210 (N_11210,N_10555,N_10934);
nand U11211 (N_11211,N_10546,N_10291);
nand U11212 (N_11212,N_10068,N_10947);
or U11213 (N_11213,N_10403,N_10340);
or U11214 (N_11214,N_10354,N_10880);
and U11215 (N_11215,N_10385,N_10198);
xor U11216 (N_11216,N_10341,N_10469);
nand U11217 (N_11217,N_10165,N_10172);
and U11218 (N_11218,N_10270,N_10759);
nor U11219 (N_11219,N_10276,N_10601);
or U11220 (N_11220,N_10147,N_10548);
and U11221 (N_11221,N_10441,N_10783);
and U11222 (N_11222,N_10575,N_10283);
and U11223 (N_11223,N_10393,N_10278);
and U11224 (N_11224,N_10320,N_10158);
or U11225 (N_11225,N_10878,N_10584);
xnor U11226 (N_11226,N_10511,N_10301);
xor U11227 (N_11227,N_10227,N_10725);
or U11228 (N_11228,N_10920,N_10027);
nor U11229 (N_11229,N_10432,N_10871);
nand U11230 (N_11230,N_10211,N_10275);
and U11231 (N_11231,N_10726,N_10228);
and U11232 (N_11232,N_10389,N_10900);
and U11233 (N_11233,N_10828,N_10552);
xnor U11234 (N_11234,N_10113,N_10673);
nand U11235 (N_11235,N_10670,N_10930);
nor U11236 (N_11236,N_10048,N_10853);
and U11237 (N_11237,N_10473,N_10803);
or U11238 (N_11238,N_10886,N_10059);
nand U11239 (N_11239,N_10706,N_10138);
nand U11240 (N_11240,N_10895,N_10774);
and U11241 (N_11241,N_10465,N_10728);
nand U11242 (N_11242,N_10671,N_10185);
xnor U11243 (N_11243,N_10742,N_10492);
and U11244 (N_11244,N_10309,N_10794);
nand U11245 (N_11245,N_10705,N_10567);
or U11246 (N_11246,N_10600,N_10117);
nand U11247 (N_11247,N_10658,N_10816);
or U11248 (N_11248,N_10651,N_10800);
and U11249 (N_11249,N_10338,N_10572);
nor U11250 (N_11250,N_10166,N_10879);
xnor U11251 (N_11251,N_10187,N_10038);
nor U11252 (N_11252,N_10327,N_10008);
or U11253 (N_11253,N_10966,N_10544);
and U11254 (N_11254,N_10924,N_10100);
nand U11255 (N_11255,N_10160,N_10861);
xor U11256 (N_11256,N_10855,N_10815);
nor U11257 (N_11257,N_10745,N_10207);
xnor U11258 (N_11258,N_10044,N_10154);
or U11259 (N_11259,N_10778,N_10343);
nor U11260 (N_11260,N_10323,N_10894);
xnor U11261 (N_11261,N_10755,N_10657);
xnor U11262 (N_11262,N_10337,N_10110);
or U11263 (N_11263,N_10175,N_10884);
xor U11264 (N_11264,N_10248,N_10483);
and U11265 (N_11265,N_10812,N_10221);
xor U11266 (N_11266,N_10236,N_10467);
and U11267 (N_11267,N_10481,N_10832);
nor U11268 (N_11268,N_10682,N_10763);
nand U11269 (N_11269,N_10239,N_10094);
and U11270 (N_11270,N_10542,N_10346);
nand U11271 (N_11271,N_10162,N_10037);
nand U11272 (N_11272,N_10570,N_10940);
nand U11273 (N_11273,N_10245,N_10502);
nor U11274 (N_11274,N_10701,N_10302);
nor U11275 (N_11275,N_10964,N_10620);
xnor U11276 (N_11276,N_10118,N_10626);
and U11277 (N_11277,N_10157,N_10287);
xnor U11278 (N_11278,N_10003,N_10252);
and U11279 (N_11279,N_10470,N_10026);
xor U11280 (N_11280,N_10500,N_10225);
or U11281 (N_11281,N_10494,N_10493);
or U11282 (N_11282,N_10867,N_10943);
nor U11283 (N_11283,N_10013,N_10730);
or U11284 (N_11284,N_10817,N_10616);
or U11285 (N_11285,N_10422,N_10583);
nor U11286 (N_11286,N_10244,N_10625);
xnor U11287 (N_11287,N_10754,N_10332);
and U11288 (N_11288,N_10194,N_10351);
nand U11289 (N_11289,N_10290,N_10080);
and U11290 (N_11290,N_10253,N_10089);
or U11291 (N_11291,N_10435,N_10994);
nor U11292 (N_11292,N_10116,N_10566);
nand U11293 (N_11293,N_10060,N_10780);
or U11294 (N_11294,N_10941,N_10516);
and U11295 (N_11295,N_10282,N_10055);
or U11296 (N_11296,N_10087,N_10931);
nand U11297 (N_11297,N_10580,N_10028);
and U11298 (N_11298,N_10863,N_10495);
and U11299 (N_11299,N_10700,N_10518);
nand U11300 (N_11300,N_10528,N_10557);
or U11301 (N_11301,N_10430,N_10717);
nand U11302 (N_11302,N_10599,N_10689);
or U11303 (N_11303,N_10669,N_10808);
nand U11304 (N_11304,N_10913,N_10798);
xor U11305 (N_11305,N_10226,N_10466);
or U11306 (N_11306,N_10394,N_10333);
and U11307 (N_11307,N_10420,N_10016);
nand U11308 (N_11308,N_10479,N_10413);
nor U11309 (N_11309,N_10750,N_10532);
nor U11310 (N_11310,N_10289,N_10353);
nor U11311 (N_11311,N_10550,N_10638);
or U11312 (N_11312,N_10672,N_10903);
nor U11313 (N_11313,N_10509,N_10539);
or U11314 (N_11314,N_10292,N_10644);
nor U11315 (N_11315,N_10949,N_10125);
xor U11316 (N_11316,N_10804,N_10938);
and U11317 (N_11317,N_10182,N_10288);
and U11318 (N_11318,N_10897,N_10907);
nand U11319 (N_11319,N_10864,N_10124);
xor U11320 (N_11320,N_10015,N_10391);
nand U11321 (N_11321,N_10034,N_10993);
or U11322 (N_11322,N_10610,N_10370);
and U11323 (N_11323,N_10076,N_10047);
nand U11324 (N_11324,N_10545,N_10128);
nand U11325 (N_11325,N_10379,N_10373);
or U11326 (N_11326,N_10326,N_10948);
xor U11327 (N_11327,N_10699,N_10345);
nor U11328 (N_11328,N_10825,N_10335);
nor U11329 (N_11329,N_10105,N_10096);
nand U11330 (N_11330,N_10254,N_10631);
xor U11331 (N_11331,N_10025,N_10156);
nor U11332 (N_11332,N_10662,N_10137);
and U11333 (N_11333,N_10054,N_10062);
nor U11334 (N_11334,N_10456,N_10564);
or U11335 (N_11335,N_10757,N_10204);
nor U11336 (N_11336,N_10461,N_10325);
nand U11337 (N_11337,N_10442,N_10438);
nand U11338 (N_11338,N_10598,N_10519);
or U11339 (N_11339,N_10971,N_10489);
or U11340 (N_11340,N_10170,N_10679);
xor U11341 (N_11341,N_10140,N_10127);
nand U11342 (N_11342,N_10865,N_10359);
nor U11343 (N_11343,N_10918,N_10768);
nand U11344 (N_11344,N_10196,N_10915);
nand U11345 (N_11345,N_10446,N_10896);
or U11346 (N_11346,N_10988,N_10656);
and U11347 (N_11347,N_10785,N_10010);
xor U11348 (N_11348,N_10174,N_10563);
or U11349 (N_11349,N_10777,N_10642);
or U11350 (N_11350,N_10970,N_10261);
or U11351 (N_11351,N_10773,N_10041);
and U11352 (N_11352,N_10406,N_10789);
nor U11353 (N_11353,N_10568,N_10925);
nand U11354 (N_11354,N_10075,N_10587);
nor U11355 (N_11355,N_10363,N_10916);
nor U11356 (N_11356,N_10277,N_10753);
nand U11357 (N_11357,N_10019,N_10111);
and U11358 (N_11358,N_10556,N_10463);
and U11359 (N_11359,N_10280,N_10250);
or U11360 (N_11360,N_10710,N_10621);
and U11361 (N_11361,N_10959,N_10476);
and U11362 (N_11362,N_10099,N_10012);
and U11363 (N_11363,N_10908,N_10247);
nand U11364 (N_11364,N_10573,N_10990);
or U11365 (N_11365,N_10224,N_10485);
and U11366 (N_11366,N_10562,N_10553);
and U11367 (N_11367,N_10790,N_10256);
nand U11368 (N_11368,N_10945,N_10381);
xor U11369 (N_11369,N_10576,N_10927);
and U11370 (N_11370,N_10152,N_10404);
and U11371 (N_11371,N_10214,N_10910);
or U11372 (N_11372,N_10889,N_10017);
nand U11373 (N_11373,N_10585,N_10814);
and U11374 (N_11374,N_10482,N_10440);
xor U11375 (N_11375,N_10212,N_10114);
or U11376 (N_11376,N_10775,N_10526);
nor U11377 (N_11377,N_10764,N_10531);
and U11378 (N_11378,N_10273,N_10831);
nand U11379 (N_11379,N_10478,N_10334);
nand U11380 (N_11380,N_10112,N_10820);
nor U11381 (N_11381,N_10922,N_10862);
and U11382 (N_11382,N_10350,N_10436);
nor U11383 (N_11383,N_10203,N_10142);
and U11384 (N_11384,N_10434,N_10877);
nor U11385 (N_11385,N_10447,N_10653);
nand U11386 (N_11386,N_10029,N_10678);
nand U11387 (N_11387,N_10648,N_10425);
nand U11388 (N_11388,N_10681,N_10149);
and U11389 (N_11389,N_10051,N_10906);
and U11390 (N_11390,N_10471,N_10266);
nand U11391 (N_11391,N_10569,N_10437);
xnor U11392 (N_11392,N_10547,N_10213);
and U11393 (N_11393,N_10860,N_10300);
and U11394 (N_11394,N_10833,N_10317);
nand U11395 (N_11395,N_10720,N_10882);
nor U11396 (N_11396,N_10506,N_10427);
nor U11397 (N_11397,N_10181,N_10503);
or U11398 (N_11398,N_10372,N_10738);
and U11399 (N_11399,N_10364,N_10869);
nor U11400 (N_11400,N_10452,N_10002);
xor U11401 (N_11401,N_10608,N_10962);
nand U11402 (N_11402,N_10772,N_10571);
xor U11403 (N_11403,N_10077,N_10974);
xnor U11404 (N_11404,N_10892,N_10965);
nand U11405 (N_11405,N_10195,N_10687);
nor U11406 (N_11406,N_10979,N_10329);
or U11407 (N_11407,N_10901,N_10271);
nor U11408 (N_11408,N_10262,N_10595);
nand U11409 (N_11409,N_10046,N_10904);
nand U11410 (N_11410,N_10986,N_10171);
nand U11411 (N_11411,N_10667,N_10074);
xor U11412 (N_11412,N_10791,N_10490);
xor U11413 (N_11413,N_10666,N_10590);
and U11414 (N_11414,N_10609,N_10821);
nor U11415 (N_11415,N_10407,N_10835);
xnor U11416 (N_11416,N_10033,N_10801);
nand U11417 (N_11417,N_10989,N_10303);
or U11418 (N_11418,N_10366,N_10684);
xnor U11419 (N_11419,N_10199,N_10477);
xnor U11420 (N_11420,N_10731,N_10009);
nand U11421 (N_11421,N_10749,N_10737);
and U11422 (N_11422,N_10536,N_10752);
xor U11423 (N_11423,N_10719,N_10776);
nor U11424 (N_11424,N_10230,N_10235);
or U11425 (N_11425,N_10650,N_10647);
or U11426 (N_11426,N_10455,N_10141);
nor U11427 (N_11427,N_10729,N_10619);
nor U11428 (N_11428,N_10488,N_10306);
or U11429 (N_11429,N_10976,N_10377);
and U11430 (N_11430,N_10708,N_10830);
and U11431 (N_11431,N_10635,N_10902);
or U11432 (N_11432,N_10517,N_10702);
and U11433 (N_11433,N_10457,N_10967);
nor U11434 (N_11434,N_10540,N_10388);
and U11435 (N_11435,N_10845,N_10936);
nor U11436 (N_11436,N_10996,N_10018);
or U11437 (N_11437,N_10085,N_10014);
and U11438 (N_11438,N_10997,N_10793);
xor U11439 (N_11439,N_10415,N_10781);
xor U11440 (N_11440,N_10933,N_10020);
nor U11441 (N_11441,N_10628,N_10978);
or U11442 (N_11442,N_10594,N_10279);
nand U11443 (N_11443,N_10944,N_10782);
nand U11444 (N_11444,N_10981,N_10512);
nor U11445 (N_11445,N_10639,N_10251);
xor U11446 (N_11446,N_10690,N_10386);
nor U11447 (N_11447,N_10259,N_10746);
nand U11448 (N_11448,N_10071,N_10692);
and U11449 (N_11449,N_10030,N_10298);
nand U11450 (N_11450,N_10022,N_10668);
and U11451 (N_11451,N_10958,N_10183);
or U11452 (N_11452,N_10484,N_10963);
nor U11453 (N_11453,N_10696,N_10795);
and U11454 (N_11454,N_10299,N_10184);
or U11455 (N_11455,N_10191,N_10308);
xnor U11456 (N_11456,N_10507,N_10163);
xor U11457 (N_11457,N_10629,N_10040);
nand U11458 (N_11458,N_10838,N_10151);
or U11459 (N_11459,N_10561,N_10357);
and U11460 (N_11460,N_10613,N_10535);
and U11461 (N_11461,N_10079,N_10848);
nand U11462 (N_11462,N_10797,N_10155);
nor U11463 (N_11463,N_10747,N_10475);
and U11464 (N_11464,N_10850,N_10744);
or U11465 (N_11465,N_10505,N_10984);
nand U11466 (N_11466,N_10538,N_10501);
and U11467 (N_11467,N_10937,N_10202);
xnor U11468 (N_11468,N_10193,N_10840);
or U11469 (N_11469,N_10844,N_10272);
nand U11470 (N_11470,N_10660,N_10057);
nor U11471 (N_11471,N_10659,N_10222);
xor U11472 (N_11472,N_10433,N_10007);
and U11473 (N_11473,N_10721,N_10093);
nor U11474 (N_11474,N_10103,N_10852);
and U11475 (N_11475,N_10188,N_10122);
nor U11476 (N_11476,N_10806,N_10352);
xor U11477 (N_11477,N_10134,N_10784);
nand U11478 (N_11478,N_10633,N_10109);
and U11479 (N_11479,N_10735,N_10691);
and U11480 (N_11480,N_10856,N_10397);
nor U11481 (N_11481,N_10858,N_10674);
xor U11482 (N_11482,N_10159,N_10315);
nor U11483 (N_11483,N_10593,N_10050);
nand U11484 (N_11484,N_10091,N_10899);
and U11485 (N_11485,N_10371,N_10875);
nand U11486 (N_11486,N_10870,N_10733);
nand U11487 (N_11487,N_10663,N_10000);
nand U11488 (N_11488,N_10847,N_10121);
nand U11489 (N_11489,N_10190,N_10637);
nand U11490 (N_11490,N_10123,N_10429);
or U11491 (N_11491,N_10229,N_10056);
nand U11492 (N_11492,N_10527,N_10756);
nor U11493 (N_11493,N_10675,N_10514);
xor U11494 (N_11494,N_10426,N_10098);
xnor U11495 (N_11495,N_10893,N_10805);
nand U11496 (N_11496,N_10957,N_10078);
nand U11497 (N_11497,N_10402,N_10146);
nand U11498 (N_11498,N_10342,N_10176);
and U11499 (N_11499,N_10150,N_10881);
or U11500 (N_11500,N_10388,N_10839);
nor U11501 (N_11501,N_10253,N_10180);
or U11502 (N_11502,N_10846,N_10899);
nand U11503 (N_11503,N_10376,N_10656);
nand U11504 (N_11504,N_10257,N_10723);
or U11505 (N_11505,N_10195,N_10430);
nor U11506 (N_11506,N_10228,N_10733);
and U11507 (N_11507,N_10212,N_10730);
nor U11508 (N_11508,N_10439,N_10253);
nand U11509 (N_11509,N_10195,N_10228);
nor U11510 (N_11510,N_10027,N_10314);
nor U11511 (N_11511,N_10599,N_10011);
nor U11512 (N_11512,N_10949,N_10241);
or U11513 (N_11513,N_10405,N_10813);
xor U11514 (N_11514,N_10386,N_10031);
or U11515 (N_11515,N_10187,N_10449);
or U11516 (N_11516,N_10903,N_10019);
and U11517 (N_11517,N_10383,N_10261);
xor U11518 (N_11518,N_10891,N_10799);
or U11519 (N_11519,N_10668,N_10380);
and U11520 (N_11520,N_10176,N_10311);
and U11521 (N_11521,N_10534,N_10469);
nor U11522 (N_11522,N_10322,N_10636);
or U11523 (N_11523,N_10406,N_10590);
nor U11524 (N_11524,N_10297,N_10815);
nor U11525 (N_11525,N_10570,N_10101);
and U11526 (N_11526,N_10358,N_10423);
or U11527 (N_11527,N_10757,N_10636);
nor U11528 (N_11528,N_10421,N_10210);
xnor U11529 (N_11529,N_10488,N_10277);
xor U11530 (N_11530,N_10778,N_10673);
nand U11531 (N_11531,N_10993,N_10129);
nand U11532 (N_11532,N_10299,N_10575);
nor U11533 (N_11533,N_10080,N_10550);
and U11534 (N_11534,N_10017,N_10241);
and U11535 (N_11535,N_10377,N_10945);
and U11536 (N_11536,N_10094,N_10119);
xnor U11537 (N_11537,N_10430,N_10592);
nand U11538 (N_11538,N_10383,N_10898);
xor U11539 (N_11539,N_10657,N_10540);
xnor U11540 (N_11540,N_10422,N_10624);
or U11541 (N_11541,N_10588,N_10322);
and U11542 (N_11542,N_10819,N_10894);
or U11543 (N_11543,N_10280,N_10831);
nand U11544 (N_11544,N_10138,N_10341);
and U11545 (N_11545,N_10229,N_10241);
nand U11546 (N_11546,N_10304,N_10468);
and U11547 (N_11547,N_10150,N_10980);
and U11548 (N_11548,N_10519,N_10285);
or U11549 (N_11549,N_10293,N_10600);
nor U11550 (N_11550,N_10665,N_10648);
or U11551 (N_11551,N_10220,N_10689);
xnor U11552 (N_11552,N_10287,N_10824);
nor U11553 (N_11553,N_10188,N_10894);
and U11554 (N_11554,N_10626,N_10387);
xor U11555 (N_11555,N_10309,N_10379);
xnor U11556 (N_11556,N_10025,N_10465);
xor U11557 (N_11557,N_10036,N_10948);
nand U11558 (N_11558,N_10963,N_10878);
xor U11559 (N_11559,N_10351,N_10963);
nand U11560 (N_11560,N_10744,N_10984);
nand U11561 (N_11561,N_10069,N_10104);
nor U11562 (N_11562,N_10436,N_10029);
or U11563 (N_11563,N_10599,N_10445);
xor U11564 (N_11564,N_10010,N_10850);
or U11565 (N_11565,N_10229,N_10118);
and U11566 (N_11566,N_10888,N_10906);
nor U11567 (N_11567,N_10910,N_10195);
and U11568 (N_11568,N_10824,N_10461);
nor U11569 (N_11569,N_10146,N_10483);
and U11570 (N_11570,N_10631,N_10417);
and U11571 (N_11571,N_10404,N_10436);
nor U11572 (N_11572,N_10195,N_10773);
or U11573 (N_11573,N_10229,N_10703);
and U11574 (N_11574,N_10379,N_10344);
or U11575 (N_11575,N_10094,N_10593);
nor U11576 (N_11576,N_10666,N_10669);
and U11577 (N_11577,N_10610,N_10237);
nor U11578 (N_11578,N_10316,N_10550);
xor U11579 (N_11579,N_10509,N_10461);
nand U11580 (N_11580,N_10739,N_10599);
and U11581 (N_11581,N_10392,N_10772);
xnor U11582 (N_11582,N_10558,N_10237);
nor U11583 (N_11583,N_10624,N_10699);
xnor U11584 (N_11584,N_10821,N_10499);
and U11585 (N_11585,N_10368,N_10888);
and U11586 (N_11586,N_10751,N_10099);
or U11587 (N_11587,N_10861,N_10954);
and U11588 (N_11588,N_10325,N_10607);
and U11589 (N_11589,N_10527,N_10602);
and U11590 (N_11590,N_10047,N_10656);
nand U11591 (N_11591,N_10907,N_10168);
nand U11592 (N_11592,N_10865,N_10084);
xnor U11593 (N_11593,N_10218,N_10224);
nor U11594 (N_11594,N_10470,N_10253);
and U11595 (N_11595,N_10840,N_10880);
xnor U11596 (N_11596,N_10749,N_10150);
or U11597 (N_11597,N_10859,N_10849);
and U11598 (N_11598,N_10846,N_10570);
xnor U11599 (N_11599,N_10977,N_10317);
and U11600 (N_11600,N_10506,N_10437);
or U11601 (N_11601,N_10548,N_10907);
nand U11602 (N_11602,N_10206,N_10663);
xnor U11603 (N_11603,N_10940,N_10122);
xor U11604 (N_11604,N_10339,N_10775);
nor U11605 (N_11605,N_10483,N_10102);
nor U11606 (N_11606,N_10887,N_10040);
nand U11607 (N_11607,N_10461,N_10053);
nor U11608 (N_11608,N_10122,N_10698);
nand U11609 (N_11609,N_10014,N_10348);
or U11610 (N_11610,N_10597,N_10835);
nand U11611 (N_11611,N_10386,N_10813);
nor U11612 (N_11612,N_10764,N_10067);
and U11613 (N_11613,N_10472,N_10079);
and U11614 (N_11614,N_10969,N_10090);
nand U11615 (N_11615,N_10700,N_10091);
nor U11616 (N_11616,N_10912,N_10446);
xnor U11617 (N_11617,N_10384,N_10747);
or U11618 (N_11618,N_10781,N_10916);
and U11619 (N_11619,N_10129,N_10013);
xnor U11620 (N_11620,N_10607,N_10632);
nor U11621 (N_11621,N_10422,N_10872);
or U11622 (N_11622,N_10192,N_10891);
nand U11623 (N_11623,N_10924,N_10756);
nand U11624 (N_11624,N_10989,N_10747);
or U11625 (N_11625,N_10006,N_10772);
nand U11626 (N_11626,N_10748,N_10416);
and U11627 (N_11627,N_10424,N_10989);
nor U11628 (N_11628,N_10113,N_10978);
nor U11629 (N_11629,N_10827,N_10185);
nand U11630 (N_11630,N_10178,N_10090);
nor U11631 (N_11631,N_10850,N_10555);
nand U11632 (N_11632,N_10140,N_10527);
nand U11633 (N_11633,N_10188,N_10251);
or U11634 (N_11634,N_10776,N_10420);
nand U11635 (N_11635,N_10920,N_10679);
xnor U11636 (N_11636,N_10181,N_10363);
and U11637 (N_11637,N_10190,N_10209);
and U11638 (N_11638,N_10689,N_10618);
xnor U11639 (N_11639,N_10345,N_10432);
xnor U11640 (N_11640,N_10981,N_10757);
nor U11641 (N_11641,N_10095,N_10645);
or U11642 (N_11642,N_10751,N_10883);
xnor U11643 (N_11643,N_10029,N_10411);
and U11644 (N_11644,N_10367,N_10282);
or U11645 (N_11645,N_10123,N_10358);
nand U11646 (N_11646,N_10330,N_10769);
nand U11647 (N_11647,N_10122,N_10208);
or U11648 (N_11648,N_10545,N_10877);
or U11649 (N_11649,N_10564,N_10639);
and U11650 (N_11650,N_10691,N_10676);
nor U11651 (N_11651,N_10438,N_10889);
nand U11652 (N_11652,N_10477,N_10675);
nor U11653 (N_11653,N_10143,N_10926);
nand U11654 (N_11654,N_10279,N_10963);
nor U11655 (N_11655,N_10940,N_10196);
xor U11656 (N_11656,N_10135,N_10104);
and U11657 (N_11657,N_10053,N_10598);
nor U11658 (N_11658,N_10665,N_10716);
and U11659 (N_11659,N_10061,N_10778);
nor U11660 (N_11660,N_10207,N_10246);
and U11661 (N_11661,N_10773,N_10073);
nand U11662 (N_11662,N_10422,N_10017);
xor U11663 (N_11663,N_10606,N_10216);
nand U11664 (N_11664,N_10083,N_10111);
nand U11665 (N_11665,N_10718,N_10836);
or U11666 (N_11666,N_10569,N_10699);
or U11667 (N_11667,N_10882,N_10527);
xor U11668 (N_11668,N_10999,N_10091);
nor U11669 (N_11669,N_10548,N_10564);
xnor U11670 (N_11670,N_10008,N_10629);
nor U11671 (N_11671,N_10277,N_10843);
or U11672 (N_11672,N_10114,N_10784);
xnor U11673 (N_11673,N_10831,N_10859);
or U11674 (N_11674,N_10860,N_10794);
nand U11675 (N_11675,N_10380,N_10459);
nand U11676 (N_11676,N_10270,N_10533);
nand U11677 (N_11677,N_10143,N_10538);
nor U11678 (N_11678,N_10840,N_10487);
and U11679 (N_11679,N_10913,N_10367);
nand U11680 (N_11680,N_10108,N_10278);
and U11681 (N_11681,N_10096,N_10760);
nand U11682 (N_11682,N_10092,N_10512);
xor U11683 (N_11683,N_10741,N_10775);
or U11684 (N_11684,N_10725,N_10270);
and U11685 (N_11685,N_10201,N_10848);
nor U11686 (N_11686,N_10390,N_10886);
xor U11687 (N_11687,N_10604,N_10375);
or U11688 (N_11688,N_10384,N_10005);
xor U11689 (N_11689,N_10215,N_10107);
and U11690 (N_11690,N_10741,N_10517);
nor U11691 (N_11691,N_10369,N_10936);
or U11692 (N_11692,N_10984,N_10036);
and U11693 (N_11693,N_10164,N_10955);
and U11694 (N_11694,N_10239,N_10909);
nor U11695 (N_11695,N_10578,N_10807);
nor U11696 (N_11696,N_10840,N_10396);
nor U11697 (N_11697,N_10194,N_10258);
or U11698 (N_11698,N_10295,N_10158);
or U11699 (N_11699,N_10069,N_10447);
nand U11700 (N_11700,N_10031,N_10892);
nand U11701 (N_11701,N_10864,N_10309);
or U11702 (N_11702,N_10115,N_10180);
nand U11703 (N_11703,N_10829,N_10356);
nand U11704 (N_11704,N_10284,N_10474);
nor U11705 (N_11705,N_10625,N_10848);
nand U11706 (N_11706,N_10296,N_10052);
xnor U11707 (N_11707,N_10501,N_10894);
and U11708 (N_11708,N_10613,N_10038);
and U11709 (N_11709,N_10883,N_10287);
or U11710 (N_11710,N_10947,N_10024);
and U11711 (N_11711,N_10564,N_10824);
nand U11712 (N_11712,N_10740,N_10791);
nand U11713 (N_11713,N_10491,N_10604);
or U11714 (N_11714,N_10195,N_10054);
and U11715 (N_11715,N_10692,N_10969);
nor U11716 (N_11716,N_10952,N_10129);
and U11717 (N_11717,N_10667,N_10606);
or U11718 (N_11718,N_10051,N_10327);
nor U11719 (N_11719,N_10513,N_10421);
and U11720 (N_11720,N_10866,N_10081);
xnor U11721 (N_11721,N_10463,N_10797);
or U11722 (N_11722,N_10197,N_10120);
xnor U11723 (N_11723,N_10469,N_10830);
and U11724 (N_11724,N_10414,N_10723);
and U11725 (N_11725,N_10123,N_10061);
or U11726 (N_11726,N_10526,N_10421);
xor U11727 (N_11727,N_10734,N_10011);
or U11728 (N_11728,N_10273,N_10054);
nand U11729 (N_11729,N_10687,N_10752);
and U11730 (N_11730,N_10024,N_10064);
xor U11731 (N_11731,N_10775,N_10343);
nand U11732 (N_11732,N_10432,N_10295);
xor U11733 (N_11733,N_10937,N_10244);
or U11734 (N_11734,N_10743,N_10148);
nand U11735 (N_11735,N_10534,N_10590);
xnor U11736 (N_11736,N_10588,N_10332);
or U11737 (N_11737,N_10955,N_10462);
or U11738 (N_11738,N_10942,N_10736);
nor U11739 (N_11739,N_10234,N_10063);
and U11740 (N_11740,N_10821,N_10533);
nand U11741 (N_11741,N_10863,N_10467);
or U11742 (N_11742,N_10660,N_10529);
nand U11743 (N_11743,N_10079,N_10592);
or U11744 (N_11744,N_10905,N_10038);
or U11745 (N_11745,N_10469,N_10558);
xnor U11746 (N_11746,N_10405,N_10775);
nand U11747 (N_11747,N_10190,N_10491);
and U11748 (N_11748,N_10251,N_10683);
and U11749 (N_11749,N_10220,N_10456);
xor U11750 (N_11750,N_10749,N_10242);
and U11751 (N_11751,N_10459,N_10141);
or U11752 (N_11752,N_10060,N_10580);
or U11753 (N_11753,N_10867,N_10684);
or U11754 (N_11754,N_10297,N_10932);
nand U11755 (N_11755,N_10680,N_10049);
nand U11756 (N_11756,N_10229,N_10952);
nor U11757 (N_11757,N_10273,N_10572);
xnor U11758 (N_11758,N_10274,N_10780);
nor U11759 (N_11759,N_10596,N_10484);
nor U11760 (N_11760,N_10336,N_10254);
xnor U11761 (N_11761,N_10815,N_10623);
and U11762 (N_11762,N_10920,N_10183);
and U11763 (N_11763,N_10860,N_10683);
xnor U11764 (N_11764,N_10498,N_10603);
and U11765 (N_11765,N_10170,N_10018);
nand U11766 (N_11766,N_10042,N_10005);
xor U11767 (N_11767,N_10399,N_10489);
and U11768 (N_11768,N_10542,N_10309);
or U11769 (N_11769,N_10463,N_10788);
xnor U11770 (N_11770,N_10997,N_10595);
xor U11771 (N_11771,N_10358,N_10200);
and U11772 (N_11772,N_10187,N_10550);
or U11773 (N_11773,N_10812,N_10805);
nand U11774 (N_11774,N_10420,N_10240);
or U11775 (N_11775,N_10256,N_10457);
nor U11776 (N_11776,N_10863,N_10257);
or U11777 (N_11777,N_10593,N_10549);
and U11778 (N_11778,N_10617,N_10910);
and U11779 (N_11779,N_10878,N_10812);
or U11780 (N_11780,N_10172,N_10350);
and U11781 (N_11781,N_10148,N_10042);
and U11782 (N_11782,N_10085,N_10480);
and U11783 (N_11783,N_10956,N_10195);
or U11784 (N_11784,N_10898,N_10030);
nor U11785 (N_11785,N_10370,N_10350);
or U11786 (N_11786,N_10902,N_10783);
nand U11787 (N_11787,N_10157,N_10783);
nor U11788 (N_11788,N_10354,N_10516);
and U11789 (N_11789,N_10079,N_10088);
nand U11790 (N_11790,N_10663,N_10719);
and U11791 (N_11791,N_10337,N_10107);
xor U11792 (N_11792,N_10778,N_10634);
xor U11793 (N_11793,N_10269,N_10460);
nand U11794 (N_11794,N_10730,N_10199);
nand U11795 (N_11795,N_10265,N_10556);
and U11796 (N_11796,N_10696,N_10248);
nand U11797 (N_11797,N_10982,N_10282);
nor U11798 (N_11798,N_10938,N_10520);
nor U11799 (N_11799,N_10170,N_10927);
nand U11800 (N_11800,N_10134,N_10206);
nand U11801 (N_11801,N_10529,N_10005);
nand U11802 (N_11802,N_10910,N_10679);
nor U11803 (N_11803,N_10506,N_10860);
or U11804 (N_11804,N_10645,N_10116);
nand U11805 (N_11805,N_10058,N_10752);
xor U11806 (N_11806,N_10179,N_10024);
or U11807 (N_11807,N_10642,N_10443);
xor U11808 (N_11808,N_10282,N_10210);
xnor U11809 (N_11809,N_10377,N_10856);
or U11810 (N_11810,N_10269,N_10598);
nand U11811 (N_11811,N_10739,N_10420);
or U11812 (N_11812,N_10284,N_10184);
and U11813 (N_11813,N_10096,N_10489);
nand U11814 (N_11814,N_10930,N_10560);
or U11815 (N_11815,N_10838,N_10824);
and U11816 (N_11816,N_10508,N_10372);
nand U11817 (N_11817,N_10473,N_10894);
or U11818 (N_11818,N_10691,N_10473);
xnor U11819 (N_11819,N_10808,N_10347);
nand U11820 (N_11820,N_10190,N_10242);
nand U11821 (N_11821,N_10135,N_10116);
nand U11822 (N_11822,N_10631,N_10876);
and U11823 (N_11823,N_10113,N_10824);
nand U11824 (N_11824,N_10846,N_10395);
nor U11825 (N_11825,N_10484,N_10081);
nor U11826 (N_11826,N_10053,N_10120);
nor U11827 (N_11827,N_10489,N_10080);
nor U11828 (N_11828,N_10677,N_10902);
nor U11829 (N_11829,N_10836,N_10016);
nand U11830 (N_11830,N_10723,N_10842);
nor U11831 (N_11831,N_10992,N_10193);
and U11832 (N_11832,N_10577,N_10606);
or U11833 (N_11833,N_10423,N_10610);
nor U11834 (N_11834,N_10363,N_10892);
nand U11835 (N_11835,N_10867,N_10893);
nor U11836 (N_11836,N_10185,N_10439);
nand U11837 (N_11837,N_10751,N_10933);
and U11838 (N_11838,N_10147,N_10528);
nand U11839 (N_11839,N_10971,N_10079);
nor U11840 (N_11840,N_10142,N_10870);
or U11841 (N_11841,N_10420,N_10888);
or U11842 (N_11842,N_10177,N_10667);
xnor U11843 (N_11843,N_10944,N_10292);
or U11844 (N_11844,N_10386,N_10623);
or U11845 (N_11845,N_10043,N_10053);
nor U11846 (N_11846,N_10425,N_10300);
xnor U11847 (N_11847,N_10379,N_10985);
xnor U11848 (N_11848,N_10300,N_10304);
xor U11849 (N_11849,N_10861,N_10116);
nand U11850 (N_11850,N_10965,N_10863);
xnor U11851 (N_11851,N_10132,N_10344);
or U11852 (N_11852,N_10430,N_10045);
nor U11853 (N_11853,N_10012,N_10837);
and U11854 (N_11854,N_10654,N_10012);
nor U11855 (N_11855,N_10559,N_10759);
xnor U11856 (N_11856,N_10330,N_10362);
and U11857 (N_11857,N_10354,N_10779);
nand U11858 (N_11858,N_10050,N_10237);
or U11859 (N_11859,N_10771,N_10827);
nand U11860 (N_11860,N_10857,N_10874);
or U11861 (N_11861,N_10800,N_10730);
xor U11862 (N_11862,N_10026,N_10343);
and U11863 (N_11863,N_10665,N_10123);
nand U11864 (N_11864,N_10122,N_10688);
nor U11865 (N_11865,N_10066,N_10358);
nand U11866 (N_11866,N_10100,N_10589);
and U11867 (N_11867,N_10715,N_10735);
nor U11868 (N_11868,N_10422,N_10314);
nor U11869 (N_11869,N_10504,N_10238);
nand U11870 (N_11870,N_10525,N_10350);
and U11871 (N_11871,N_10322,N_10690);
or U11872 (N_11872,N_10247,N_10556);
or U11873 (N_11873,N_10282,N_10225);
and U11874 (N_11874,N_10389,N_10868);
and U11875 (N_11875,N_10717,N_10243);
or U11876 (N_11876,N_10178,N_10097);
xnor U11877 (N_11877,N_10441,N_10944);
xor U11878 (N_11878,N_10228,N_10301);
xnor U11879 (N_11879,N_10572,N_10002);
and U11880 (N_11880,N_10080,N_10937);
or U11881 (N_11881,N_10706,N_10128);
and U11882 (N_11882,N_10535,N_10299);
and U11883 (N_11883,N_10998,N_10385);
nor U11884 (N_11884,N_10390,N_10221);
or U11885 (N_11885,N_10037,N_10519);
nor U11886 (N_11886,N_10490,N_10190);
xnor U11887 (N_11887,N_10055,N_10337);
or U11888 (N_11888,N_10228,N_10124);
and U11889 (N_11889,N_10301,N_10693);
nand U11890 (N_11890,N_10516,N_10294);
xnor U11891 (N_11891,N_10222,N_10592);
or U11892 (N_11892,N_10922,N_10274);
and U11893 (N_11893,N_10813,N_10781);
nand U11894 (N_11894,N_10264,N_10878);
nor U11895 (N_11895,N_10548,N_10849);
and U11896 (N_11896,N_10314,N_10488);
and U11897 (N_11897,N_10579,N_10886);
xnor U11898 (N_11898,N_10040,N_10544);
nand U11899 (N_11899,N_10742,N_10207);
and U11900 (N_11900,N_10594,N_10458);
xor U11901 (N_11901,N_10167,N_10358);
nand U11902 (N_11902,N_10128,N_10567);
nand U11903 (N_11903,N_10034,N_10327);
xnor U11904 (N_11904,N_10085,N_10442);
xor U11905 (N_11905,N_10502,N_10612);
nor U11906 (N_11906,N_10277,N_10961);
nor U11907 (N_11907,N_10363,N_10558);
nand U11908 (N_11908,N_10063,N_10008);
xor U11909 (N_11909,N_10027,N_10347);
xor U11910 (N_11910,N_10043,N_10633);
xor U11911 (N_11911,N_10540,N_10428);
or U11912 (N_11912,N_10071,N_10300);
and U11913 (N_11913,N_10249,N_10641);
and U11914 (N_11914,N_10114,N_10108);
nand U11915 (N_11915,N_10131,N_10926);
nand U11916 (N_11916,N_10278,N_10603);
xor U11917 (N_11917,N_10699,N_10077);
nor U11918 (N_11918,N_10470,N_10166);
xnor U11919 (N_11919,N_10502,N_10447);
and U11920 (N_11920,N_10719,N_10796);
nor U11921 (N_11921,N_10598,N_10000);
and U11922 (N_11922,N_10881,N_10148);
or U11923 (N_11923,N_10269,N_10341);
nor U11924 (N_11924,N_10384,N_10750);
or U11925 (N_11925,N_10357,N_10634);
nand U11926 (N_11926,N_10278,N_10302);
and U11927 (N_11927,N_10125,N_10070);
or U11928 (N_11928,N_10107,N_10431);
or U11929 (N_11929,N_10733,N_10700);
nand U11930 (N_11930,N_10413,N_10511);
or U11931 (N_11931,N_10881,N_10289);
xor U11932 (N_11932,N_10486,N_10790);
xor U11933 (N_11933,N_10814,N_10445);
or U11934 (N_11934,N_10007,N_10516);
nand U11935 (N_11935,N_10072,N_10327);
or U11936 (N_11936,N_10006,N_10038);
nand U11937 (N_11937,N_10306,N_10293);
and U11938 (N_11938,N_10227,N_10364);
nand U11939 (N_11939,N_10327,N_10605);
or U11940 (N_11940,N_10988,N_10677);
nor U11941 (N_11941,N_10628,N_10511);
or U11942 (N_11942,N_10467,N_10202);
and U11943 (N_11943,N_10161,N_10515);
nor U11944 (N_11944,N_10879,N_10310);
nor U11945 (N_11945,N_10753,N_10609);
and U11946 (N_11946,N_10231,N_10015);
and U11947 (N_11947,N_10706,N_10344);
nor U11948 (N_11948,N_10073,N_10115);
nor U11949 (N_11949,N_10566,N_10257);
and U11950 (N_11950,N_10875,N_10597);
or U11951 (N_11951,N_10101,N_10397);
nand U11952 (N_11952,N_10311,N_10361);
and U11953 (N_11953,N_10029,N_10515);
and U11954 (N_11954,N_10997,N_10735);
nand U11955 (N_11955,N_10728,N_10789);
xnor U11956 (N_11956,N_10141,N_10665);
or U11957 (N_11957,N_10734,N_10151);
or U11958 (N_11958,N_10379,N_10728);
or U11959 (N_11959,N_10372,N_10183);
nand U11960 (N_11960,N_10993,N_10214);
and U11961 (N_11961,N_10620,N_10821);
nand U11962 (N_11962,N_10294,N_10566);
xor U11963 (N_11963,N_10545,N_10145);
or U11964 (N_11964,N_10084,N_10167);
and U11965 (N_11965,N_10212,N_10413);
nand U11966 (N_11966,N_10527,N_10177);
nor U11967 (N_11967,N_10979,N_10176);
nand U11968 (N_11968,N_10505,N_10349);
or U11969 (N_11969,N_10403,N_10782);
xor U11970 (N_11970,N_10567,N_10841);
nor U11971 (N_11971,N_10339,N_10834);
xnor U11972 (N_11972,N_10820,N_10023);
xnor U11973 (N_11973,N_10613,N_10196);
xnor U11974 (N_11974,N_10291,N_10673);
or U11975 (N_11975,N_10379,N_10664);
or U11976 (N_11976,N_10200,N_10801);
nor U11977 (N_11977,N_10078,N_10122);
nor U11978 (N_11978,N_10489,N_10095);
and U11979 (N_11979,N_10791,N_10047);
nor U11980 (N_11980,N_10667,N_10662);
or U11981 (N_11981,N_10248,N_10552);
nor U11982 (N_11982,N_10323,N_10239);
nor U11983 (N_11983,N_10100,N_10023);
nand U11984 (N_11984,N_10565,N_10867);
or U11985 (N_11985,N_10341,N_10385);
nor U11986 (N_11986,N_10101,N_10743);
and U11987 (N_11987,N_10255,N_10744);
nand U11988 (N_11988,N_10082,N_10241);
nand U11989 (N_11989,N_10781,N_10370);
xor U11990 (N_11990,N_10139,N_10349);
nor U11991 (N_11991,N_10547,N_10206);
nor U11992 (N_11992,N_10334,N_10301);
xnor U11993 (N_11993,N_10071,N_10416);
nand U11994 (N_11994,N_10273,N_10647);
or U11995 (N_11995,N_10394,N_10917);
nor U11996 (N_11996,N_10027,N_10243);
nor U11997 (N_11997,N_10351,N_10813);
nor U11998 (N_11998,N_10738,N_10893);
nor U11999 (N_11999,N_10591,N_10415);
or U12000 (N_12000,N_11285,N_11804);
and U12001 (N_12001,N_11210,N_11503);
nand U12002 (N_12002,N_11510,N_11987);
or U12003 (N_12003,N_11824,N_11003);
and U12004 (N_12004,N_11640,N_11175);
or U12005 (N_12005,N_11363,N_11538);
nor U12006 (N_12006,N_11414,N_11269);
or U12007 (N_12007,N_11726,N_11975);
or U12008 (N_12008,N_11055,N_11806);
nand U12009 (N_12009,N_11309,N_11189);
nor U12010 (N_12010,N_11877,N_11536);
xnor U12011 (N_12011,N_11662,N_11511);
nor U12012 (N_12012,N_11650,N_11761);
nor U12013 (N_12013,N_11360,N_11765);
xor U12014 (N_12014,N_11995,N_11386);
or U12015 (N_12015,N_11322,N_11502);
and U12016 (N_12016,N_11951,N_11289);
nor U12017 (N_12017,N_11604,N_11950);
nand U12018 (N_12018,N_11695,N_11678);
nor U12019 (N_12019,N_11953,N_11149);
nor U12020 (N_12020,N_11153,N_11395);
and U12021 (N_12021,N_11193,N_11145);
nor U12022 (N_12022,N_11571,N_11310);
nand U12023 (N_12023,N_11264,N_11708);
nand U12024 (N_12024,N_11667,N_11833);
nand U12025 (N_12025,N_11434,N_11711);
nand U12026 (N_12026,N_11181,N_11487);
nand U12027 (N_12027,N_11431,N_11560);
and U12028 (N_12028,N_11301,N_11859);
nand U12029 (N_12029,N_11334,N_11092);
and U12030 (N_12030,N_11446,N_11702);
or U12031 (N_12031,N_11074,N_11735);
xnor U12032 (N_12032,N_11519,N_11687);
or U12033 (N_12033,N_11323,N_11663);
nand U12034 (N_12034,N_11023,N_11771);
nand U12035 (N_12035,N_11298,N_11040);
nand U12036 (N_12036,N_11991,N_11682);
or U12037 (N_12037,N_11148,N_11842);
nor U12038 (N_12038,N_11306,N_11076);
xnor U12039 (N_12039,N_11444,N_11154);
or U12040 (N_12040,N_11686,N_11647);
nor U12041 (N_12041,N_11295,N_11960);
nand U12042 (N_12042,N_11930,N_11531);
xnor U12043 (N_12043,N_11988,N_11794);
xnor U12044 (N_12044,N_11331,N_11247);
xor U12045 (N_12045,N_11245,N_11151);
nor U12046 (N_12046,N_11954,N_11225);
and U12047 (N_12047,N_11773,N_11392);
and U12048 (N_12048,N_11525,N_11004);
or U12049 (N_12049,N_11753,N_11863);
and U12050 (N_12050,N_11411,N_11905);
xnor U12051 (N_12051,N_11948,N_11177);
xnor U12052 (N_12052,N_11373,N_11768);
and U12053 (N_12053,N_11106,N_11160);
nand U12054 (N_12054,N_11522,N_11978);
xor U12055 (N_12055,N_11020,N_11209);
and U12056 (N_12056,N_11613,N_11451);
nor U12057 (N_12057,N_11828,N_11725);
or U12058 (N_12058,N_11653,N_11913);
nand U12059 (N_12059,N_11450,N_11752);
or U12060 (N_12060,N_11772,N_11214);
and U12061 (N_12061,N_11815,N_11250);
and U12062 (N_12062,N_11565,N_11699);
nor U12063 (N_12063,N_11294,N_11164);
nor U12064 (N_12064,N_11595,N_11024);
or U12065 (N_12065,N_11258,N_11848);
xnor U12066 (N_12066,N_11559,N_11195);
nor U12067 (N_12067,N_11675,N_11637);
xor U12068 (N_12068,N_11071,N_11933);
xnor U12069 (N_12069,N_11758,N_11775);
and U12070 (N_12070,N_11038,N_11066);
xnor U12071 (N_12071,N_11688,N_11564);
nor U12072 (N_12072,N_11410,N_11255);
xnor U12073 (N_12073,N_11015,N_11664);
and U12074 (N_12074,N_11671,N_11769);
nand U12075 (N_12075,N_11485,N_11293);
nor U12076 (N_12076,N_11856,N_11219);
or U12077 (N_12077,N_11308,N_11589);
nor U12078 (N_12078,N_11998,N_11129);
and U12079 (N_12079,N_11563,N_11982);
and U12080 (N_12080,N_11469,N_11047);
or U12081 (N_12081,N_11277,N_11412);
or U12082 (N_12082,N_11871,N_11555);
or U12083 (N_12083,N_11803,N_11025);
xor U12084 (N_12084,N_11668,N_11914);
or U12085 (N_12085,N_11173,N_11026);
nor U12086 (N_12086,N_11719,N_11490);
nand U12087 (N_12087,N_11528,N_11078);
and U12088 (N_12088,N_11496,N_11939);
or U12089 (N_12089,N_11603,N_11121);
xnor U12090 (N_12090,N_11032,N_11862);
xor U12091 (N_12091,N_11442,N_11353);
or U12092 (N_12092,N_11274,N_11578);
and U12093 (N_12093,N_11095,N_11657);
or U12094 (N_12094,N_11103,N_11002);
and U12095 (N_12095,N_11669,N_11826);
or U12096 (N_12096,N_11275,N_11986);
and U12097 (N_12097,N_11072,N_11733);
nor U12098 (N_12098,N_11116,N_11260);
or U12099 (N_12099,N_11415,N_11413);
xor U12100 (N_12100,N_11248,N_11529);
and U12101 (N_12101,N_11350,N_11318);
xnor U12102 (N_12102,N_11198,N_11498);
and U12103 (N_12103,N_11229,N_11608);
or U12104 (N_12104,N_11419,N_11867);
or U12105 (N_12105,N_11718,N_11906);
nand U12106 (N_12106,N_11601,N_11847);
xor U12107 (N_12107,N_11272,N_11408);
and U12108 (N_12108,N_11019,N_11981);
nand U12109 (N_12109,N_11463,N_11377);
nand U12110 (N_12110,N_11741,N_11850);
nand U12111 (N_12111,N_11748,N_11985);
and U12112 (N_12112,N_11369,N_11455);
and U12113 (N_12113,N_11259,N_11715);
nand U12114 (N_12114,N_11633,N_11799);
and U12115 (N_12115,N_11812,N_11213);
nor U12116 (N_12116,N_11174,N_11468);
nor U12117 (N_12117,N_11261,N_11287);
nand U12118 (N_12118,N_11556,N_11014);
and U12119 (N_12119,N_11792,N_11119);
and U12120 (N_12120,N_11239,N_11888);
nor U12121 (N_12121,N_11049,N_11453);
nor U12122 (N_12122,N_11027,N_11409);
nor U12123 (N_12123,N_11537,N_11892);
nand U12124 (N_12124,N_11626,N_11944);
nor U12125 (N_12125,N_11817,N_11013);
and U12126 (N_12126,N_11482,N_11827);
xor U12127 (N_12127,N_11325,N_11146);
or U12128 (N_12128,N_11227,N_11231);
nor U12129 (N_12129,N_11838,N_11832);
nor U12130 (N_12130,N_11479,N_11574);
and U12131 (N_12131,N_11391,N_11441);
or U12132 (N_12132,N_11314,N_11628);
or U12133 (N_12133,N_11139,N_11232);
or U12134 (N_12134,N_11253,N_11355);
and U12135 (N_12135,N_11852,N_11062);
and U12136 (N_12136,N_11836,N_11632);
xor U12137 (N_12137,N_11242,N_11083);
xnor U12138 (N_12138,N_11330,N_11104);
xor U12139 (N_12139,N_11235,N_11897);
nor U12140 (N_12140,N_11730,N_11790);
and U12141 (N_12141,N_11512,N_11100);
or U12142 (N_12142,N_11869,N_11202);
or U12143 (N_12143,N_11418,N_11620);
nor U12144 (N_12144,N_11224,N_11102);
xor U12145 (N_12145,N_11581,N_11236);
nand U12146 (N_12146,N_11857,N_11120);
nor U12147 (N_12147,N_11138,N_11636);
or U12148 (N_12148,N_11456,N_11327);
or U12149 (N_12149,N_11825,N_11185);
or U12150 (N_12150,N_11720,N_11966);
xnor U12151 (N_12151,N_11739,N_11118);
nor U12152 (N_12152,N_11263,N_11942);
nand U12153 (N_12153,N_11732,N_11683);
nor U12154 (N_12154,N_11370,N_11801);
and U12155 (N_12155,N_11142,N_11917);
or U12156 (N_12156,N_11839,N_11477);
nor U12157 (N_12157,N_11679,N_11648);
or U12158 (N_12158,N_11738,N_11473);
xor U12159 (N_12159,N_11197,N_11305);
xnor U12160 (N_12160,N_11467,N_11627);
nor U12161 (N_12161,N_11896,N_11459);
or U12162 (N_12162,N_11539,N_11816);
or U12163 (N_12163,N_11465,N_11449);
nand U12164 (N_12164,N_11217,N_11329);
or U12165 (N_12165,N_11523,N_11124);
and U12166 (N_12166,N_11883,N_11976);
and U12167 (N_12167,N_11374,N_11929);
nor U12168 (N_12168,N_11313,N_11935);
nand U12169 (N_12169,N_11461,N_11706);
xnor U12170 (N_12170,N_11077,N_11553);
and U12171 (N_12171,N_11656,N_11721);
nand U12172 (N_12172,N_11508,N_11005);
xnor U12173 (N_12173,N_11271,N_11596);
nand U12174 (N_12174,N_11705,N_11171);
nor U12175 (N_12175,N_11584,N_11182);
nand U12176 (N_12176,N_11882,N_11407);
xnor U12177 (N_12177,N_11364,N_11915);
nand U12178 (N_12178,N_11290,N_11051);
or U12179 (N_12179,N_11088,N_11167);
or U12180 (N_12180,N_11731,N_11776);
and U12181 (N_12181,N_11616,N_11190);
nand U12182 (N_12182,N_11552,N_11952);
and U12183 (N_12183,N_11244,N_11048);
xor U12184 (N_12184,N_11107,N_11033);
nand U12185 (N_12185,N_11136,N_11543);
and U12186 (N_12186,N_11932,N_11056);
or U12187 (N_12187,N_11911,N_11743);
xnor U12188 (N_12188,N_11516,N_11645);
nor U12189 (N_12189,N_11110,N_11159);
and U12190 (N_12190,N_11868,N_11387);
xor U12191 (N_12191,N_11054,N_11416);
nand U12192 (N_12192,N_11090,N_11689);
nand U12193 (N_12193,N_11751,N_11297);
xor U12194 (N_12194,N_11349,N_11215);
or U12195 (N_12195,N_11432,N_11494);
and U12196 (N_12196,N_11381,N_11423);
and U12197 (N_12197,N_11226,N_11569);
and U12198 (N_12198,N_11646,N_11317);
nor U12199 (N_12199,N_11017,N_11524);
or U12200 (N_12200,N_11240,N_11813);
nor U12201 (N_12201,N_11207,N_11782);
nand U12202 (N_12202,N_11841,N_11440);
xor U12203 (N_12203,N_11938,N_11161);
xor U12204 (N_12204,N_11874,N_11001);
or U12205 (N_12205,N_11729,N_11899);
nand U12206 (N_12206,N_11582,N_11819);
and U12207 (N_12207,N_11808,N_11814);
xnor U12208 (N_12208,N_11094,N_11820);
and U12209 (N_12209,N_11784,N_11457);
or U12210 (N_12210,N_11818,N_11402);
nand U12211 (N_12211,N_11396,N_11375);
nor U12212 (N_12212,N_11143,N_11478);
nor U12213 (N_12213,N_11372,N_11172);
nand U12214 (N_12214,N_11362,N_11131);
xor U12215 (N_12215,N_11117,N_11504);
or U12216 (N_12216,N_11579,N_11879);
or U12217 (N_12217,N_11105,N_11714);
nand U12218 (N_12218,N_11918,N_11891);
nand U12219 (N_12219,N_11521,N_11787);
xnor U12220 (N_12220,N_11204,N_11368);
or U12221 (N_12221,N_11141,N_11974);
xnor U12222 (N_12222,N_11400,N_11111);
xnor U12223 (N_12223,N_11216,N_11576);
or U12224 (N_12224,N_11534,N_11357);
and U12225 (N_12225,N_11041,N_11351);
and U12226 (N_12226,N_11922,N_11946);
nand U12227 (N_12227,N_11475,N_11831);
and U12228 (N_12228,N_11320,N_11108);
xnor U12229 (N_12229,N_11061,N_11619);
nor U12230 (N_12230,N_11973,N_11977);
nor U12231 (N_12231,N_11727,N_11070);
xnor U12232 (N_12232,N_11670,N_11462);
and U12233 (N_12233,N_11635,N_11542);
xor U12234 (N_12234,N_11588,N_11992);
nor U12235 (N_12235,N_11065,N_11540);
or U12236 (N_12236,N_11179,N_11053);
xor U12237 (N_12237,N_11163,N_11520);
nor U12238 (N_12238,N_11900,N_11747);
xor U12239 (N_12239,N_11218,N_11898);
or U12240 (N_12240,N_11749,N_11166);
xor U12241 (N_12241,N_11677,N_11492);
xor U12242 (N_12242,N_11507,N_11655);
or U12243 (N_12243,N_11445,N_11886);
and U12244 (N_12244,N_11925,N_11499);
nand U12245 (N_12245,N_11389,N_11694);
or U12246 (N_12246,N_11183,N_11889);
nand U12247 (N_12247,N_11592,N_11428);
nand U12248 (N_12248,N_11967,N_11266);
nor U12249 (N_12249,N_11280,N_11007);
or U12250 (N_12250,N_11703,N_11319);
and U12251 (N_12251,N_11821,N_11602);
nand U12252 (N_12252,N_11237,N_11672);
xor U12253 (N_12253,N_11756,N_11777);
xnor U12254 (N_12254,N_11165,N_11222);
nor U12255 (N_12255,N_11211,N_11354);
and U12256 (N_12256,N_11780,N_11567);
and U12257 (N_12257,N_11957,N_11379);
nor U12258 (N_12258,N_11380,N_11435);
and U12259 (N_12259,N_11779,N_11958);
xnor U12260 (N_12260,N_11760,N_11403);
or U12261 (N_12261,N_11994,N_11358);
and U12262 (N_12262,N_11610,N_11846);
xnor U12263 (N_12263,N_11778,N_11206);
and U12264 (N_12264,N_11367,N_11547);
and U12265 (N_12265,N_11843,N_11770);
or U12266 (N_12266,N_11554,N_11470);
or U12267 (N_12267,N_11698,N_11132);
nor U12268 (N_12268,N_11430,N_11447);
xor U12269 (N_12269,N_11249,N_11844);
and U12270 (N_12270,N_11388,N_11965);
nand U12271 (N_12271,N_11223,N_11279);
and U12272 (N_12272,N_11234,N_11904);
or U12273 (N_12273,N_11737,N_11155);
xnor U12274 (N_12274,N_11979,N_11800);
or U12275 (N_12275,N_11028,N_11359);
xnor U12276 (N_12276,N_11724,N_11058);
nor U12277 (N_12277,N_11178,N_11692);
nand U12278 (N_12278,N_11199,N_11654);
or U12279 (N_12279,N_11972,N_11681);
nand U12280 (N_12280,N_11561,N_11805);
and U12281 (N_12281,N_11057,N_11580);
nor U12282 (N_12282,N_11039,N_11937);
nor U12283 (N_12283,N_11858,N_11684);
or U12284 (N_12284,N_11191,N_11282);
and U12285 (N_12285,N_11383,N_11855);
and U12286 (N_12286,N_11866,N_11212);
nand U12287 (N_12287,N_11208,N_11625);
xnor U12288 (N_12288,N_11949,N_11114);
nand U12289 (N_12289,N_11587,N_11332);
xnor U12290 (N_12290,N_11876,N_11097);
nand U12291 (N_12291,N_11546,N_11658);
xor U12292 (N_12292,N_11638,N_11283);
or U12293 (N_12293,N_11068,N_11067);
xnor U12294 (N_12294,N_11575,N_11042);
and U12295 (N_12295,N_11600,N_11623);
and U12296 (N_12296,N_11940,N_11811);
xnor U12297 (N_12297,N_11085,N_11113);
xor U12298 (N_12298,N_11716,N_11962);
or U12299 (N_12299,N_11674,N_11754);
xor U12300 (N_12300,N_11505,N_11016);
nor U12301 (N_12301,N_11486,N_11109);
nand U12302 (N_12302,N_11927,N_11018);
and U12303 (N_12303,N_11059,N_11481);
nor U12304 (N_12304,N_11156,N_11452);
nor U12305 (N_12305,N_11073,N_11276);
and U12306 (N_12306,N_11562,N_11810);
nor U12307 (N_12307,N_11880,N_11609);
and U12308 (N_12308,N_11887,N_11598);
nand U12309 (N_12309,N_11786,N_11643);
nand U12310 (N_12310,N_11630,N_11194);
nand U12311 (N_12311,N_11712,N_11956);
xor U12312 (N_12312,N_11781,N_11541);
nand U12313 (N_12313,N_11926,N_11518);
and U12314 (N_12314,N_11570,N_11284);
nand U12315 (N_12315,N_11338,N_11493);
and U12316 (N_12316,N_11000,N_11286);
and U12317 (N_12317,N_11734,N_11710);
nor U12318 (N_12318,N_11251,N_11125);
nand U12319 (N_12319,N_11500,N_11809);
and U12320 (N_12320,N_11081,N_11795);
nand U12321 (N_12321,N_11851,N_11115);
nand U12322 (N_12322,N_11495,N_11659);
nor U12323 (N_12323,N_11513,N_11312);
nor U12324 (N_12324,N_11509,N_11928);
nor U12325 (N_12325,N_11082,N_11265);
and U12326 (N_12326,N_11728,N_11168);
or U12327 (N_12327,N_11797,N_11586);
nor U12328 (N_12328,N_11093,N_11943);
nor U12329 (N_12329,N_11220,N_11549);
nand U12330 (N_12330,N_11759,N_11573);
nand U12331 (N_12331,N_11134,N_11947);
xor U12332 (N_12332,N_11558,N_11910);
or U12333 (N_12333,N_11750,N_11830);
or U12334 (N_12334,N_11158,N_11079);
and U12335 (N_12335,N_11064,N_11696);
xnor U12336 (N_12336,N_11270,N_11834);
nor U12337 (N_12337,N_11321,N_11180);
and U12338 (N_12338,N_11384,N_11624);
and U12339 (N_12339,N_11989,N_11955);
or U12340 (N_12340,N_11766,N_11717);
and U12341 (N_12341,N_11621,N_11983);
nand U12342 (N_12342,N_11346,N_11599);
nand U12343 (N_12343,N_11527,N_11029);
or U12344 (N_12344,N_11660,N_11009);
nor U12345 (N_12345,N_11371,N_11326);
xor U12346 (N_12346,N_11366,N_11590);
nand U12347 (N_12347,N_11228,N_11789);
nor U12348 (N_12348,N_11533,N_11902);
or U12349 (N_12349,N_11112,N_11012);
xnor U12350 (N_12350,N_11673,N_11288);
and U12351 (N_12351,N_11666,N_11031);
or U12352 (N_12352,N_11488,N_11837);
or U12353 (N_12353,N_11652,N_11438);
or U12354 (N_12354,N_11568,N_11709);
xnor U12355 (N_12355,N_11256,N_11884);
and U12356 (N_12356,N_11936,N_11087);
nor U12357 (N_12357,N_11639,N_11304);
or U12358 (N_12358,N_11996,N_11548);
or U12359 (N_12359,N_11514,N_11680);
or U12360 (N_12360,N_11091,N_11861);
or U12361 (N_12361,N_11740,N_11333);
or U12362 (N_12362,N_11458,N_11895);
nand U12363 (N_12363,N_11420,N_11931);
nor U12364 (N_12364,N_11894,N_11075);
xor U12365 (N_12365,N_11634,N_11422);
nor U12366 (N_12366,N_11483,N_11835);
and U12367 (N_12367,N_11722,N_11744);
nor U12368 (N_12368,N_11909,N_11133);
or U12369 (N_12369,N_11296,N_11480);
xnor U12370 (N_12370,N_11267,N_11292);
nand U12371 (N_12371,N_11901,N_11170);
nor U12372 (N_12372,N_11631,N_11060);
and U12373 (N_12373,N_11397,N_11299);
nand U12374 (N_12374,N_11169,N_11959);
or U12375 (N_12375,N_11890,N_11200);
and U12376 (N_12376,N_11783,N_11745);
or U12377 (N_12377,N_11893,N_11829);
and U12378 (N_12378,N_11424,N_11532);
nor U12379 (N_12379,N_11788,N_11390);
or U12380 (N_12380,N_11572,N_11585);
or U12381 (N_12381,N_11970,N_11315);
nor U12382 (N_12382,N_11046,N_11137);
nor U12383 (N_12383,N_11466,N_11594);
and U12384 (N_12384,N_11644,N_11437);
nand U12385 (N_12385,N_11152,N_11324);
or U12386 (N_12386,N_11063,N_11617);
xor U12387 (N_12387,N_11035,N_11961);
and U12388 (N_12388,N_11096,N_11484);
nand U12389 (N_12389,N_11089,N_11622);
nand U12390 (N_12390,N_11147,N_11246);
nor U12391 (N_12391,N_11941,N_11454);
xnor U12392 (N_12392,N_11713,N_11685);
xnor U12393 (N_12393,N_11690,N_11188);
nor U12394 (N_12394,N_11036,N_11997);
xnor U12395 (N_12395,N_11291,N_11238);
and U12396 (N_12396,N_11629,N_11870);
nor U12397 (N_12397,N_11340,N_11881);
or U12398 (N_12398,N_11394,N_11405);
xnor U12399 (N_12399,N_11262,N_11807);
xnor U12400 (N_12400,N_11385,N_11421);
nand U12401 (N_12401,N_11593,N_11281);
or U12402 (N_12402,N_11489,N_11607);
nor U12403 (N_12403,N_11924,N_11872);
nand U12404 (N_12404,N_11615,N_11257);
and U12405 (N_12405,N_11971,N_11404);
xor U12406 (N_12406,N_11964,N_11885);
or U12407 (N_12407,N_11642,N_11530);
nand U12408 (N_12408,N_11126,N_11535);
and U12409 (N_12409,N_11436,N_11127);
nand U12410 (N_12410,N_11551,N_11614);
nand U12411 (N_12411,N_11343,N_11550);
xor U12412 (N_12412,N_11597,N_11853);
nand U12413 (N_12413,N_11476,N_11921);
nand U12414 (N_12414,N_11448,N_11908);
xnor U12415 (N_12415,N_11796,N_11344);
or U12416 (N_12416,N_11854,N_11365);
xnor U12417 (N_12417,N_11472,N_11187);
xnor U12418 (N_12418,N_11241,N_11864);
xnor U12419 (N_12419,N_11471,N_11798);
or U12420 (N_12420,N_11665,N_11254);
nand U12421 (N_12421,N_11612,N_11425);
or U12422 (N_12422,N_11393,N_11491);
or U12423 (N_12423,N_11316,N_11865);
or U12424 (N_12424,N_11157,N_11707);
and U12425 (N_12425,N_11268,N_11044);
and U12426 (N_12426,N_11591,N_11767);
nand U12427 (N_12427,N_11583,N_11378);
nand U12428 (N_12428,N_11233,N_11526);
or U12429 (N_12429,N_11774,N_11348);
and U12430 (N_12430,N_11205,N_11460);
and U12431 (N_12431,N_11221,N_11086);
and U12432 (N_12432,N_11878,N_11045);
nand U12433 (N_12433,N_11544,N_11907);
or U12434 (N_12434,N_11736,N_11356);
nor U12435 (N_12435,N_11080,N_11150);
and U12436 (N_12436,N_11341,N_11618);
or U12437 (N_12437,N_11515,N_11243);
xor U12438 (N_12438,N_11201,N_11700);
and U12439 (N_12439,N_11037,N_11676);
xnor U12440 (N_12440,N_11300,N_11697);
nor U12441 (N_12441,N_11566,N_11920);
or U12442 (N_12442,N_11984,N_11873);
nand U12443 (N_12443,N_11345,N_11693);
nand U12444 (N_12444,N_11969,N_11130);
and U12445 (N_12445,N_11605,N_11849);
nand U12446 (N_12446,N_11135,N_11303);
nor U12447 (N_12447,N_11822,N_11649);
or U12448 (N_12448,N_11651,N_11742);
xnor U12449 (N_12449,N_11845,N_11577);
xnor U12450 (N_12450,N_11361,N_11474);
and U12451 (N_12451,N_11443,N_11429);
and U12452 (N_12452,N_11517,N_11802);
xor U12453 (N_12453,N_11339,N_11328);
xor U12454 (N_12454,N_11030,N_11793);
nor U12455 (N_12455,N_11144,N_11050);
and U12456 (N_12456,N_11426,N_11433);
and U12457 (N_12457,N_11764,N_11501);
and U12458 (N_12458,N_11034,N_11311);
or U12459 (N_12459,N_11337,N_11439);
or U12460 (N_12460,N_11382,N_11762);
nor U12461 (N_12461,N_11335,N_11043);
nand U12462 (N_12462,N_11008,N_11427);
nand U12463 (N_12463,N_11184,N_11230);
nand U12464 (N_12464,N_11763,N_11860);
xnor U12465 (N_12465,N_11342,N_11123);
xnor U12466 (N_12466,N_11176,N_11347);
nand U12467 (N_12467,N_11376,N_11011);
nand U12468 (N_12468,N_11785,N_11999);
nand U12469 (N_12469,N_11606,N_11022);
nor U12470 (N_12470,N_11307,N_11140);
nand U12471 (N_12471,N_11723,N_11192);
or U12472 (N_12472,N_11757,N_11464);
xor U12473 (N_12473,N_11401,N_11691);
and U12474 (N_12474,N_11398,N_11968);
and U12475 (N_12475,N_11203,N_11196);
nand U12476 (N_12476,N_11084,N_11010);
or U12477 (N_12477,N_11641,N_11912);
xor U12478 (N_12478,N_11352,N_11052);
nor U12479 (N_12479,N_11661,N_11122);
xnor U12480 (N_12480,N_11098,N_11336);
xor U12481 (N_12481,N_11945,N_11823);
and U12482 (N_12482,N_11923,N_11916);
or U12483 (N_12483,N_11990,N_11497);
nor U12484 (N_12484,N_11099,N_11278);
nor U12485 (N_12485,N_11101,N_11021);
or U12486 (N_12486,N_11128,N_11701);
and U12487 (N_12487,N_11934,N_11302);
nand U12488 (N_12488,N_11746,N_11506);
nor U12489 (N_12489,N_11252,N_11704);
or U12490 (N_12490,N_11186,N_11993);
nand U12491 (N_12491,N_11417,N_11840);
nor U12492 (N_12492,N_11875,N_11006);
nor U12493 (N_12493,N_11162,N_11557);
xor U12494 (N_12494,N_11545,N_11406);
xor U12495 (N_12495,N_11069,N_11903);
nand U12496 (N_12496,N_11611,N_11980);
or U12497 (N_12497,N_11791,N_11273);
xnor U12498 (N_12498,N_11399,N_11963);
and U12499 (N_12499,N_11755,N_11919);
nor U12500 (N_12500,N_11084,N_11240);
or U12501 (N_12501,N_11276,N_11811);
nor U12502 (N_12502,N_11021,N_11128);
and U12503 (N_12503,N_11374,N_11456);
xor U12504 (N_12504,N_11842,N_11936);
nor U12505 (N_12505,N_11526,N_11142);
nor U12506 (N_12506,N_11587,N_11842);
and U12507 (N_12507,N_11946,N_11167);
or U12508 (N_12508,N_11894,N_11586);
nor U12509 (N_12509,N_11937,N_11759);
xor U12510 (N_12510,N_11601,N_11945);
or U12511 (N_12511,N_11070,N_11721);
nand U12512 (N_12512,N_11676,N_11496);
or U12513 (N_12513,N_11805,N_11401);
nand U12514 (N_12514,N_11676,N_11234);
xnor U12515 (N_12515,N_11964,N_11222);
or U12516 (N_12516,N_11528,N_11209);
or U12517 (N_12517,N_11172,N_11735);
or U12518 (N_12518,N_11028,N_11518);
nor U12519 (N_12519,N_11884,N_11616);
nor U12520 (N_12520,N_11457,N_11370);
xor U12521 (N_12521,N_11757,N_11861);
nand U12522 (N_12522,N_11482,N_11431);
or U12523 (N_12523,N_11652,N_11637);
nor U12524 (N_12524,N_11645,N_11529);
nor U12525 (N_12525,N_11010,N_11778);
or U12526 (N_12526,N_11598,N_11955);
nor U12527 (N_12527,N_11099,N_11441);
nor U12528 (N_12528,N_11134,N_11127);
xnor U12529 (N_12529,N_11009,N_11301);
nor U12530 (N_12530,N_11835,N_11798);
or U12531 (N_12531,N_11595,N_11489);
nand U12532 (N_12532,N_11186,N_11719);
nor U12533 (N_12533,N_11687,N_11978);
nand U12534 (N_12534,N_11137,N_11266);
nand U12535 (N_12535,N_11985,N_11453);
or U12536 (N_12536,N_11134,N_11714);
nor U12537 (N_12537,N_11474,N_11619);
nand U12538 (N_12538,N_11553,N_11471);
and U12539 (N_12539,N_11686,N_11344);
nand U12540 (N_12540,N_11636,N_11187);
and U12541 (N_12541,N_11585,N_11953);
or U12542 (N_12542,N_11918,N_11388);
nor U12543 (N_12543,N_11803,N_11097);
or U12544 (N_12544,N_11252,N_11539);
xnor U12545 (N_12545,N_11456,N_11306);
xnor U12546 (N_12546,N_11723,N_11365);
and U12547 (N_12547,N_11367,N_11863);
or U12548 (N_12548,N_11393,N_11721);
and U12549 (N_12549,N_11451,N_11919);
or U12550 (N_12550,N_11809,N_11097);
nor U12551 (N_12551,N_11054,N_11791);
and U12552 (N_12552,N_11439,N_11382);
and U12553 (N_12553,N_11987,N_11862);
nor U12554 (N_12554,N_11939,N_11632);
xnor U12555 (N_12555,N_11366,N_11584);
nor U12556 (N_12556,N_11395,N_11686);
nand U12557 (N_12557,N_11717,N_11202);
xnor U12558 (N_12558,N_11421,N_11234);
and U12559 (N_12559,N_11987,N_11134);
xnor U12560 (N_12560,N_11690,N_11587);
nand U12561 (N_12561,N_11086,N_11005);
nor U12562 (N_12562,N_11596,N_11876);
and U12563 (N_12563,N_11015,N_11575);
nor U12564 (N_12564,N_11180,N_11950);
and U12565 (N_12565,N_11677,N_11827);
nand U12566 (N_12566,N_11175,N_11832);
xnor U12567 (N_12567,N_11032,N_11804);
nand U12568 (N_12568,N_11683,N_11073);
and U12569 (N_12569,N_11289,N_11467);
xnor U12570 (N_12570,N_11249,N_11444);
or U12571 (N_12571,N_11501,N_11731);
or U12572 (N_12572,N_11086,N_11885);
nand U12573 (N_12573,N_11041,N_11714);
nand U12574 (N_12574,N_11632,N_11518);
and U12575 (N_12575,N_11613,N_11133);
and U12576 (N_12576,N_11000,N_11565);
nor U12577 (N_12577,N_11879,N_11432);
xnor U12578 (N_12578,N_11855,N_11823);
or U12579 (N_12579,N_11618,N_11022);
nand U12580 (N_12580,N_11802,N_11322);
nor U12581 (N_12581,N_11791,N_11242);
nand U12582 (N_12582,N_11421,N_11771);
xor U12583 (N_12583,N_11952,N_11550);
nand U12584 (N_12584,N_11643,N_11749);
or U12585 (N_12585,N_11570,N_11400);
nand U12586 (N_12586,N_11947,N_11196);
and U12587 (N_12587,N_11176,N_11963);
nor U12588 (N_12588,N_11082,N_11222);
xnor U12589 (N_12589,N_11000,N_11577);
xor U12590 (N_12590,N_11913,N_11602);
nor U12591 (N_12591,N_11598,N_11481);
and U12592 (N_12592,N_11856,N_11741);
xnor U12593 (N_12593,N_11535,N_11898);
or U12594 (N_12594,N_11965,N_11274);
xor U12595 (N_12595,N_11043,N_11049);
and U12596 (N_12596,N_11932,N_11509);
and U12597 (N_12597,N_11901,N_11293);
and U12598 (N_12598,N_11448,N_11422);
or U12599 (N_12599,N_11768,N_11978);
or U12600 (N_12600,N_11366,N_11024);
and U12601 (N_12601,N_11602,N_11491);
or U12602 (N_12602,N_11676,N_11590);
or U12603 (N_12603,N_11149,N_11363);
or U12604 (N_12604,N_11150,N_11383);
or U12605 (N_12605,N_11945,N_11493);
nand U12606 (N_12606,N_11607,N_11535);
and U12607 (N_12607,N_11826,N_11117);
nand U12608 (N_12608,N_11042,N_11839);
or U12609 (N_12609,N_11535,N_11560);
xnor U12610 (N_12610,N_11256,N_11246);
xnor U12611 (N_12611,N_11891,N_11060);
nor U12612 (N_12612,N_11123,N_11057);
nand U12613 (N_12613,N_11599,N_11975);
and U12614 (N_12614,N_11045,N_11847);
and U12615 (N_12615,N_11755,N_11814);
or U12616 (N_12616,N_11112,N_11226);
and U12617 (N_12617,N_11541,N_11102);
nor U12618 (N_12618,N_11195,N_11306);
xor U12619 (N_12619,N_11384,N_11584);
xor U12620 (N_12620,N_11864,N_11520);
nor U12621 (N_12621,N_11735,N_11528);
and U12622 (N_12622,N_11879,N_11037);
xnor U12623 (N_12623,N_11184,N_11604);
or U12624 (N_12624,N_11057,N_11372);
and U12625 (N_12625,N_11800,N_11017);
xor U12626 (N_12626,N_11004,N_11935);
nand U12627 (N_12627,N_11726,N_11307);
nor U12628 (N_12628,N_11471,N_11700);
and U12629 (N_12629,N_11148,N_11224);
nand U12630 (N_12630,N_11950,N_11727);
or U12631 (N_12631,N_11329,N_11514);
nand U12632 (N_12632,N_11775,N_11517);
and U12633 (N_12633,N_11256,N_11398);
and U12634 (N_12634,N_11415,N_11064);
and U12635 (N_12635,N_11631,N_11053);
nor U12636 (N_12636,N_11116,N_11397);
or U12637 (N_12637,N_11017,N_11600);
nand U12638 (N_12638,N_11397,N_11876);
xor U12639 (N_12639,N_11081,N_11005);
nand U12640 (N_12640,N_11339,N_11083);
xnor U12641 (N_12641,N_11680,N_11401);
nand U12642 (N_12642,N_11220,N_11790);
or U12643 (N_12643,N_11717,N_11103);
nor U12644 (N_12644,N_11791,N_11820);
nand U12645 (N_12645,N_11466,N_11141);
nand U12646 (N_12646,N_11401,N_11508);
nor U12647 (N_12647,N_11783,N_11974);
nand U12648 (N_12648,N_11179,N_11115);
nor U12649 (N_12649,N_11266,N_11084);
and U12650 (N_12650,N_11566,N_11926);
xor U12651 (N_12651,N_11027,N_11540);
xor U12652 (N_12652,N_11857,N_11345);
nand U12653 (N_12653,N_11074,N_11730);
nor U12654 (N_12654,N_11831,N_11244);
and U12655 (N_12655,N_11518,N_11757);
xnor U12656 (N_12656,N_11164,N_11009);
xnor U12657 (N_12657,N_11501,N_11898);
xor U12658 (N_12658,N_11955,N_11772);
nand U12659 (N_12659,N_11981,N_11088);
and U12660 (N_12660,N_11903,N_11401);
and U12661 (N_12661,N_11943,N_11389);
nor U12662 (N_12662,N_11715,N_11638);
xnor U12663 (N_12663,N_11881,N_11190);
nand U12664 (N_12664,N_11679,N_11321);
nand U12665 (N_12665,N_11444,N_11665);
xor U12666 (N_12666,N_11035,N_11108);
and U12667 (N_12667,N_11163,N_11318);
or U12668 (N_12668,N_11250,N_11233);
and U12669 (N_12669,N_11325,N_11208);
or U12670 (N_12670,N_11686,N_11781);
and U12671 (N_12671,N_11999,N_11534);
and U12672 (N_12672,N_11301,N_11452);
nor U12673 (N_12673,N_11488,N_11519);
nor U12674 (N_12674,N_11849,N_11032);
xnor U12675 (N_12675,N_11185,N_11772);
or U12676 (N_12676,N_11036,N_11368);
xor U12677 (N_12677,N_11081,N_11750);
xnor U12678 (N_12678,N_11535,N_11477);
nand U12679 (N_12679,N_11873,N_11409);
xor U12680 (N_12680,N_11714,N_11156);
nor U12681 (N_12681,N_11346,N_11370);
xnor U12682 (N_12682,N_11739,N_11134);
nor U12683 (N_12683,N_11728,N_11839);
and U12684 (N_12684,N_11107,N_11833);
and U12685 (N_12685,N_11314,N_11654);
and U12686 (N_12686,N_11468,N_11022);
nor U12687 (N_12687,N_11445,N_11988);
and U12688 (N_12688,N_11903,N_11712);
and U12689 (N_12689,N_11176,N_11268);
nor U12690 (N_12690,N_11698,N_11244);
nor U12691 (N_12691,N_11799,N_11153);
or U12692 (N_12692,N_11704,N_11730);
xor U12693 (N_12693,N_11479,N_11056);
nand U12694 (N_12694,N_11650,N_11943);
and U12695 (N_12695,N_11797,N_11424);
nand U12696 (N_12696,N_11540,N_11592);
or U12697 (N_12697,N_11380,N_11416);
nand U12698 (N_12698,N_11763,N_11824);
xnor U12699 (N_12699,N_11110,N_11794);
xnor U12700 (N_12700,N_11168,N_11892);
or U12701 (N_12701,N_11812,N_11773);
nor U12702 (N_12702,N_11383,N_11943);
and U12703 (N_12703,N_11679,N_11928);
xnor U12704 (N_12704,N_11593,N_11547);
or U12705 (N_12705,N_11213,N_11266);
xor U12706 (N_12706,N_11422,N_11451);
and U12707 (N_12707,N_11301,N_11117);
and U12708 (N_12708,N_11942,N_11226);
nand U12709 (N_12709,N_11757,N_11835);
xor U12710 (N_12710,N_11321,N_11591);
nand U12711 (N_12711,N_11973,N_11846);
nor U12712 (N_12712,N_11007,N_11021);
or U12713 (N_12713,N_11819,N_11875);
or U12714 (N_12714,N_11539,N_11583);
xnor U12715 (N_12715,N_11073,N_11301);
nand U12716 (N_12716,N_11774,N_11294);
or U12717 (N_12717,N_11306,N_11865);
or U12718 (N_12718,N_11694,N_11057);
xnor U12719 (N_12719,N_11041,N_11746);
or U12720 (N_12720,N_11489,N_11628);
xnor U12721 (N_12721,N_11351,N_11544);
xnor U12722 (N_12722,N_11898,N_11724);
nor U12723 (N_12723,N_11472,N_11914);
or U12724 (N_12724,N_11157,N_11032);
or U12725 (N_12725,N_11215,N_11978);
xnor U12726 (N_12726,N_11877,N_11174);
and U12727 (N_12727,N_11668,N_11971);
nor U12728 (N_12728,N_11807,N_11059);
nand U12729 (N_12729,N_11628,N_11370);
nand U12730 (N_12730,N_11681,N_11437);
and U12731 (N_12731,N_11643,N_11538);
nand U12732 (N_12732,N_11294,N_11625);
and U12733 (N_12733,N_11070,N_11851);
or U12734 (N_12734,N_11953,N_11199);
or U12735 (N_12735,N_11773,N_11642);
nand U12736 (N_12736,N_11198,N_11970);
nand U12737 (N_12737,N_11581,N_11633);
nor U12738 (N_12738,N_11176,N_11937);
and U12739 (N_12739,N_11440,N_11935);
nor U12740 (N_12740,N_11008,N_11308);
or U12741 (N_12741,N_11061,N_11158);
nor U12742 (N_12742,N_11126,N_11528);
or U12743 (N_12743,N_11600,N_11419);
or U12744 (N_12744,N_11322,N_11539);
xor U12745 (N_12745,N_11349,N_11252);
or U12746 (N_12746,N_11970,N_11709);
xnor U12747 (N_12747,N_11223,N_11571);
or U12748 (N_12748,N_11553,N_11075);
nand U12749 (N_12749,N_11084,N_11064);
xor U12750 (N_12750,N_11946,N_11596);
or U12751 (N_12751,N_11633,N_11693);
or U12752 (N_12752,N_11372,N_11676);
nor U12753 (N_12753,N_11360,N_11529);
nand U12754 (N_12754,N_11132,N_11895);
nor U12755 (N_12755,N_11917,N_11780);
nand U12756 (N_12756,N_11019,N_11380);
and U12757 (N_12757,N_11607,N_11608);
nor U12758 (N_12758,N_11723,N_11030);
or U12759 (N_12759,N_11947,N_11830);
or U12760 (N_12760,N_11462,N_11974);
nor U12761 (N_12761,N_11649,N_11570);
nand U12762 (N_12762,N_11108,N_11256);
and U12763 (N_12763,N_11869,N_11093);
nor U12764 (N_12764,N_11543,N_11402);
and U12765 (N_12765,N_11735,N_11164);
or U12766 (N_12766,N_11255,N_11775);
nand U12767 (N_12767,N_11633,N_11610);
xor U12768 (N_12768,N_11099,N_11781);
xnor U12769 (N_12769,N_11188,N_11634);
and U12770 (N_12770,N_11811,N_11233);
nand U12771 (N_12771,N_11242,N_11315);
xnor U12772 (N_12772,N_11957,N_11822);
nand U12773 (N_12773,N_11191,N_11148);
xnor U12774 (N_12774,N_11481,N_11733);
nand U12775 (N_12775,N_11309,N_11473);
nand U12776 (N_12776,N_11128,N_11621);
or U12777 (N_12777,N_11784,N_11673);
nor U12778 (N_12778,N_11386,N_11780);
xor U12779 (N_12779,N_11527,N_11142);
nand U12780 (N_12780,N_11017,N_11356);
or U12781 (N_12781,N_11979,N_11403);
and U12782 (N_12782,N_11208,N_11975);
nor U12783 (N_12783,N_11774,N_11134);
xor U12784 (N_12784,N_11555,N_11391);
nor U12785 (N_12785,N_11524,N_11501);
xor U12786 (N_12786,N_11423,N_11196);
or U12787 (N_12787,N_11189,N_11299);
and U12788 (N_12788,N_11575,N_11825);
xnor U12789 (N_12789,N_11895,N_11164);
and U12790 (N_12790,N_11588,N_11686);
xnor U12791 (N_12791,N_11215,N_11520);
and U12792 (N_12792,N_11314,N_11361);
xnor U12793 (N_12793,N_11609,N_11217);
or U12794 (N_12794,N_11736,N_11408);
nand U12795 (N_12795,N_11061,N_11360);
xor U12796 (N_12796,N_11552,N_11653);
or U12797 (N_12797,N_11152,N_11910);
xnor U12798 (N_12798,N_11263,N_11888);
xor U12799 (N_12799,N_11676,N_11398);
and U12800 (N_12800,N_11918,N_11222);
xor U12801 (N_12801,N_11066,N_11611);
xor U12802 (N_12802,N_11242,N_11022);
nor U12803 (N_12803,N_11328,N_11836);
and U12804 (N_12804,N_11838,N_11621);
xnor U12805 (N_12805,N_11542,N_11274);
xor U12806 (N_12806,N_11640,N_11989);
or U12807 (N_12807,N_11179,N_11116);
or U12808 (N_12808,N_11741,N_11341);
and U12809 (N_12809,N_11107,N_11305);
xnor U12810 (N_12810,N_11748,N_11778);
nand U12811 (N_12811,N_11875,N_11499);
xnor U12812 (N_12812,N_11844,N_11269);
nor U12813 (N_12813,N_11595,N_11621);
and U12814 (N_12814,N_11080,N_11677);
or U12815 (N_12815,N_11480,N_11474);
nor U12816 (N_12816,N_11721,N_11094);
or U12817 (N_12817,N_11416,N_11953);
nor U12818 (N_12818,N_11832,N_11816);
nor U12819 (N_12819,N_11354,N_11837);
or U12820 (N_12820,N_11561,N_11617);
xor U12821 (N_12821,N_11476,N_11501);
nor U12822 (N_12822,N_11835,N_11527);
xor U12823 (N_12823,N_11289,N_11481);
nor U12824 (N_12824,N_11062,N_11178);
nor U12825 (N_12825,N_11677,N_11865);
xnor U12826 (N_12826,N_11581,N_11886);
nand U12827 (N_12827,N_11031,N_11797);
and U12828 (N_12828,N_11044,N_11653);
nor U12829 (N_12829,N_11556,N_11338);
nand U12830 (N_12830,N_11513,N_11767);
or U12831 (N_12831,N_11095,N_11594);
or U12832 (N_12832,N_11603,N_11165);
nor U12833 (N_12833,N_11057,N_11864);
nand U12834 (N_12834,N_11127,N_11357);
and U12835 (N_12835,N_11390,N_11466);
nor U12836 (N_12836,N_11112,N_11938);
xor U12837 (N_12837,N_11774,N_11035);
or U12838 (N_12838,N_11796,N_11453);
and U12839 (N_12839,N_11416,N_11480);
xnor U12840 (N_12840,N_11796,N_11920);
nand U12841 (N_12841,N_11305,N_11662);
xor U12842 (N_12842,N_11030,N_11421);
nand U12843 (N_12843,N_11058,N_11822);
nand U12844 (N_12844,N_11747,N_11027);
nor U12845 (N_12845,N_11016,N_11713);
nor U12846 (N_12846,N_11151,N_11619);
or U12847 (N_12847,N_11953,N_11066);
nor U12848 (N_12848,N_11581,N_11945);
or U12849 (N_12849,N_11538,N_11323);
or U12850 (N_12850,N_11013,N_11885);
or U12851 (N_12851,N_11327,N_11914);
and U12852 (N_12852,N_11783,N_11502);
and U12853 (N_12853,N_11974,N_11397);
and U12854 (N_12854,N_11737,N_11538);
and U12855 (N_12855,N_11570,N_11159);
or U12856 (N_12856,N_11538,N_11739);
nor U12857 (N_12857,N_11675,N_11331);
xor U12858 (N_12858,N_11770,N_11133);
nor U12859 (N_12859,N_11175,N_11629);
nor U12860 (N_12860,N_11322,N_11979);
xnor U12861 (N_12861,N_11393,N_11884);
nand U12862 (N_12862,N_11613,N_11313);
or U12863 (N_12863,N_11977,N_11254);
xor U12864 (N_12864,N_11020,N_11319);
or U12865 (N_12865,N_11040,N_11481);
and U12866 (N_12866,N_11082,N_11873);
and U12867 (N_12867,N_11325,N_11126);
or U12868 (N_12868,N_11093,N_11996);
and U12869 (N_12869,N_11683,N_11807);
xor U12870 (N_12870,N_11370,N_11982);
xnor U12871 (N_12871,N_11656,N_11404);
nor U12872 (N_12872,N_11742,N_11266);
nand U12873 (N_12873,N_11240,N_11593);
and U12874 (N_12874,N_11605,N_11407);
nand U12875 (N_12875,N_11694,N_11439);
and U12876 (N_12876,N_11823,N_11683);
or U12877 (N_12877,N_11370,N_11070);
nor U12878 (N_12878,N_11046,N_11331);
and U12879 (N_12879,N_11407,N_11204);
or U12880 (N_12880,N_11165,N_11187);
or U12881 (N_12881,N_11749,N_11420);
or U12882 (N_12882,N_11685,N_11131);
and U12883 (N_12883,N_11929,N_11571);
or U12884 (N_12884,N_11236,N_11264);
xor U12885 (N_12885,N_11273,N_11269);
nand U12886 (N_12886,N_11827,N_11522);
xnor U12887 (N_12887,N_11093,N_11405);
xor U12888 (N_12888,N_11279,N_11345);
nand U12889 (N_12889,N_11901,N_11896);
and U12890 (N_12890,N_11532,N_11885);
nand U12891 (N_12891,N_11878,N_11916);
xnor U12892 (N_12892,N_11690,N_11189);
nor U12893 (N_12893,N_11352,N_11230);
nand U12894 (N_12894,N_11702,N_11413);
nor U12895 (N_12895,N_11145,N_11377);
nor U12896 (N_12896,N_11507,N_11845);
xnor U12897 (N_12897,N_11661,N_11178);
nand U12898 (N_12898,N_11554,N_11439);
or U12899 (N_12899,N_11067,N_11899);
nor U12900 (N_12900,N_11671,N_11890);
or U12901 (N_12901,N_11480,N_11081);
xnor U12902 (N_12902,N_11971,N_11031);
nand U12903 (N_12903,N_11730,N_11638);
and U12904 (N_12904,N_11851,N_11198);
nand U12905 (N_12905,N_11489,N_11985);
nand U12906 (N_12906,N_11415,N_11162);
nand U12907 (N_12907,N_11729,N_11394);
or U12908 (N_12908,N_11253,N_11660);
nand U12909 (N_12909,N_11471,N_11375);
nor U12910 (N_12910,N_11665,N_11632);
or U12911 (N_12911,N_11457,N_11537);
or U12912 (N_12912,N_11403,N_11834);
or U12913 (N_12913,N_11594,N_11072);
and U12914 (N_12914,N_11788,N_11837);
xor U12915 (N_12915,N_11944,N_11486);
xnor U12916 (N_12916,N_11295,N_11388);
nor U12917 (N_12917,N_11662,N_11779);
or U12918 (N_12918,N_11671,N_11997);
or U12919 (N_12919,N_11730,N_11197);
and U12920 (N_12920,N_11910,N_11762);
nor U12921 (N_12921,N_11568,N_11116);
nor U12922 (N_12922,N_11586,N_11355);
and U12923 (N_12923,N_11215,N_11040);
or U12924 (N_12924,N_11023,N_11259);
nand U12925 (N_12925,N_11591,N_11506);
nand U12926 (N_12926,N_11307,N_11723);
xor U12927 (N_12927,N_11026,N_11105);
and U12928 (N_12928,N_11602,N_11481);
and U12929 (N_12929,N_11172,N_11864);
and U12930 (N_12930,N_11210,N_11096);
nand U12931 (N_12931,N_11360,N_11386);
nand U12932 (N_12932,N_11054,N_11467);
xor U12933 (N_12933,N_11783,N_11132);
or U12934 (N_12934,N_11025,N_11260);
nand U12935 (N_12935,N_11937,N_11308);
xor U12936 (N_12936,N_11355,N_11473);
or U12937 (N_12937,N_11150,N_11622);
or U12938 (N_12938,N_11054,N_11858);
nand U12939 (N_12939,N_11880,N_11648);
nand U12940 (N_12940,N_11684,N_11520);
nand U12941 (N_12941,N_11911,N_11014);
xnor U12942 (N_12942,N_11241,N_11170);
and U12943 (N_12943,N_11393,N_11944);
and U12944 (N_12944,N_11856,N_11123);
nor U12945 (N_12945,N_11136,N_11327);
nand U12946 (N_12946,N_11759,N_11985);
xnor U12947 (N_12947,N_11599,N_11045);
nor U12948 (N_12948,N_11711,N_11491);
nand U12949 (N_12949,N_11425,N_11912);
nand U12950 (N_12950,N_11351,N_11904);
or U12951 (N_12951,N_11058,N_11538);
and U12952 (N_12952,N_11195,N_11662);
xor U12953 (N_12953,N_11401,N_11084);
nor U12954 (N_12954,N_11023,N_11751);
xor U12955 (N_12955,N_11674,N_11863);
nand U12956 (N_12956,N_11383,N_11453);
and U12957 (N_12957,N_11132,N_11329);
nand U12958 (N_12958,N_11013,N_11649);
xnor U12959 (N_12959,N_11913,N_11328);
nand U12960 (N_12960,N_11500,N_11093);
and U12961 (N_12961,N_11414,N_11230);
nor U12962 (N_12962,N_11160,N_11568);
or U12963 (N_12963,N_11875,N_11055);
nand U12964 (N_12964,N_11011,N_11044);
xnor U12965 (N_12965,N_11567,N_11971);
and U12966 (N_12966,N_11051,N_11000);
xnor U12967 (N_12967,N_11913,N_11607);
nand U12968 (N_12968,N_11385,N_11037);
or U12969 (N_12969,N_11693,N_11495);
or U12970 (N_12970,N_11429,N_11544);
nor U12971 (N_12971,N_11425,N_11443);
or U12972 (N_12972,N_11067,N_11677);
or U12973 (N_12973,N_11307,N_11361);
and U12974 (N_12974,N_11273,N_11822);
xor U12975 (N_12975,N_11280,N_11566);
and U12976 (N_12976,N_11809,N_11314);
and U12977 (N_12977,N_11278,N_11682);
nor U12978 (N_12978,N_11335,N_11554);
or U12979 (N_12979,N_11188,N_11758);
xor U12980 (N_12980,N_11675,N_11326);
nor U12981 (N_12981,N_11676,N_11057);
xnor U12982 (N_12982,N_11924,N_11497);
and U12983 (N_12983,N_11505,N_11904);
or U12984 (N_12984,N_11938,N_11642);
or U12985 (N_12985,N_11798,N_11352);
xnor U12986 (N_12986,N_11906,N_11139);
nor U12987 (N_12987,N_11918,N_11510);
nand U12988 (N_12988,N_11780,N_11044);
or U12989 (N_12989,N_11655,N_11627);
nor U12990 (N_12990,N_11346,N_11944);
nand U12991 (N_12991,N_11794,N_11140);
nor U12992 (N_12992,N_11215,N_11874);
xnor U12993 (N_12993,N_11761,N_11162);
or U12994 (N_12994,N_11261,N_11705);
or U12995 (N_12995,N_11847,N_11565);
nor U12996 (N_12996,N_11467,N_11074);
or U12997 (N_12997,N_11400,N_11399);
nand U12998 (N_12998,N_11684,N_11742);
xor U12999 (N_12999,N_11575,N_11999);
nor U13000 (N_13000,N_12860,N_12614);
or U13001 (N_13001,N_12078,N_12779);
and U13002 (N_13002,N_12071,N_12205);
and U13003 (N_13003,N_12488,N_12380);
or U13004 (N_13004,N_12930,N_12715);
and U13005 (N_13005,N_12076,N_12894);
nor U13006 (N_13006,N_12199,N_12829);
or U13007 (N_13007,N_12814,N_12274);
nor U13008 (N_13008,N_12867,N_12469);
xor U13009 (N_13009,N_12815,N_12887);
and U13010 (N_13010,N_12929,N_12838);
or U13011 (N_13011,N_12408,N_12223);
xnor U13012 (N_13012,N_12377,N_12140);
xnor U13013 (N_13013,N_12917,N_12703);
nor U13014 (N_13014,N_12508,N_12214);
nor U13015 (N_13015,N_12372,N_12483);
or U13016 (N_13016,N_12624,N_12954);
or U13017 (N_13017,N_12901,N_12858);
xnor U13018 (N_13018,N_12869,N_12203);
or U13019 (N_13019,N_12177,N_12899);
and U13020 (N_13020,N_12077,N_12880);
or U13021 (N_13021,N_12861,N_12857);
or U13022 (N_13022,N_12485,N_12403);
and U13023 (N_13023,N_12603,N_12760);
nand U13024 (N_13024,N_12597,N_12415);
and U13025 (N_13025,N_12632,N_12583);
xnor U13026 (N_13026,N_12547,N_12736);
nor U13027 (N_13027,N_12472,N_12315);
xor U13028 (N_13028,N_12619,N_12280);
or U13029 (N_13029,N_12184,N_12623);
nor U13030 (N_13030,N_12376,N_12594);
or U13031 (N_13031,N_12176,N_12863);
and U13032 (N_13032,N_12119,N_12093);
or U13033 (N_13033,N_12981,N_12672);
or U13034 (N_13034,N_12246,N_12748);
or U13035 (N_13035,N_12367,N_12729);
or U13036 (N_13036,N_12254,N_12724);
or U13037 (N_13037,N_12806,N_12505);
nor U13038 (N_13038,N_12731,N_12757);
and U13039 (N_13039,N_12633,N_12875);
nor U13040 (N_13040,N_12573,N_12166);
or U13041 (N_13041,N_12978,N_12965);
nand U13042 (N_13042,N_12397,N_12790);
nand U13043 (N_13043,N_12097,N_12892);
nand U13044 (N_13044,N_12481,N_12183);
nor U13045 (N_13045,N_12523,N_12443);
nand U13046 (N_13046,N_12865,N_12781);
or U13047 (N_13047,N_12296,N_12771);
nor U13048 (N_13048,N_12522,N_12253);
nand U13049 (N_13049,N_12299,N_12088);
nand U13050 (N_13050,N_12373,N_12359);
or U13051 (N_13051,N_12992,N_12767);
nand U13052 (N_13052,N_12264,N_12019);
xor U13053 (N_13053,N_12031,N_12144);
nor U13054 (N_13054,N_12318,N_12425);
nand U13055 (N_13055,N_12646,N_12255);
nand U13056 (N_13056,N_12354,N_12514);
and U13057 (N_13057,N_12083,N_12162);
xor U13058 (N_13058,N_12292,N_12655);
or U13059 (N_13059,N_12566,N_12378);
and U13060 (N_13060,N_12035,N_12947);
and U13061 (N_13061,N_12284,N_12471);
and U13062 (N_13062,N_12329,N_12711);
and U13063 (N_13063,N_12922,N_12555);
nor U13064 (N_13064,N_12404,N_12651);
and U13065 (N_13065,N_12700,N_12387);
xor U13066 (N_13066,N_12540,N_12448);
or U13067 (N_13067,N_12449,N_12761);
nand U13068 (N_13068,N_12504,N_12942);
and U13069 (N_13069,N_12568,N_12009);
nand U13070 (N_13070,N_12098,N_12730);
nor U13071 (N_13071,N_12828,N_12155);
or U13072 (N_13072,N_12052,N_12844);
and U13073 (N_13073,N_12014,N_12147);
nor U13074 (N_13074,N_12412,N_12371);
or U13075 (N_13075,N_12734,N_12741);
nand U13076 (N_13076,N_12985,N_12440);
nand U13077 (N_13077,N_12447,N_12805);
or U13078 (N_13078,N_12626,N_12820);
or U13079 (N_13079,N_12532,N_12972);
nand U13080 (N_13080,N_12392,N_12735);
or U13081 (N_13081,N_12721,N_12245);
or U13082 (N_13082,N_12324,N_12200);
nor U13083 (N_13083,N_12021,N_12989);
or U13084 (N_13084,N_12285,N_12435);
xor U13085 (N_13085,N_12773,N_12780);
nor U13086 (N_13086,N_12852,N_12235);
and U13087 (N_13087,N_12219,N_12596);
nand U13088 (N_13088,N_12821,N_12466);
nor U13089 (N_13089,N_12610,N_12365);
or U13090 (N_13090,N_12634,N_12968);
and U13091 (N_13091,N_12710,N_12616);
and U13092 (N_13092,N_12990,N_12146);
xor U13093 (N_13093,N_12690,N_12240);
xnor U13094 (N_13094,N_12565,N_12525);
or U13095 (N_13095,N_12552,N_12537);
or U13096 (N_13096,N_12092,N_12158);
or U13097 (N_13097,N_12490,N_12178);
or U13098 (N_13098,N_12231,N_12502);
xor U13099 (N_13099,N_12360,N_12074);
or U13100 (N_13100,N_12313,N_12227);
xor U13101 (N_13101,N_12928,N_12430);
and U13102 (N_13102,N_12062,N_12452);
and U13103 (N_13103,N_12055,N_12800);
or U13104 (N_13104,N_12694,N_12840);
nand U13105 (N_13105,N_12749,N_12496);
and U13106 (N_13106,N_12519,N_12333);
nor U13107 (N_13107,N_12289,N_12298);
nand U13108 (N_13108,N_12370,N_12001);
xnor U13109 (N_13109,N_12418,N_12453);
nor U13110 (N_13110,N_12139,N_12629);
xnor U13111 (N_13111,N_12004,N_12877);
or U13112 (N_13112,N_12163,N_12334);
nor U13113 (N_13113,N_12216,N_12669);
xor U13114 (N_13114,N_12770,N_12718);
nor U13115 (N_13115,N_12266,N_12919);
nor U13116 (N_13116,N_12667,N_12520);
and U13117 (N_13117,N_12966,N_12516);
nand U13118 (N_13118,N_12218,N_12916);
nor U13119 (N_13119,N_12217,N_12132);
nor U13120 (N_13120,N_12808,N_12862);
nor U13121 (N_13121,N_12643,N_12664);
nor U13122 (N_13122,N_12560,N_12906);
nand U13123 (N_13123,N_12924,N_12192);
and U13124 (N_13124,N_12891,N_12524);
and U13125 (N_13125,N_12799,N_12578);
or U13126 (N_13126,N_12382,N_12189);
or U13127 (N_13127,N_12586,N_12866);
nor U13128 (N_13128,N_12048,N_12512);
nor U13129 (N_13129,N_12982,N_12356);
xnor U13130 (N_13130,N_12394,N_12258);
nor U13131 (N_13131,N_12951,N_12259);
nand U13132 (N_13132,N_12558,N_12889);
xor U13133 (N_13133,N_12641,N_12445);
and U13134 (N_13134,N_12131,N_12903);
nor U13135 (N_13135,N_12243,N_12225);
and U13136 (N_13136,N_12328,N_12503);
nand U13137 (N_13137,N_12959,N_12896);
and U13138 (N_13138,N_12247,N_12495);
or U13139 (N_13139,N_12263,N_12104);
xnor U13140 (N_13140,N_12340,N_12708);
nor U13141 (N_13141,N_12347,N_12389);
nand U13142 (N_13142,N_12918,N_12213);
xnor U13143 (N_13143,N_12087,N_12234);
and U13144 (N_13144,N_12618,N_12036);
and U13145 (N_13145,N_12644,N_12434);
nor U13146 (N_13146,N_12145,N_12539);
or U13147 (N_13147,N_12744,N_12383);
or U13148 (N_13148,N_12794,N_12701);
nand U13149 (N_13149,N_12513,N_12493);
or U13150 (N_13150,N_12498,N_12697);
or U13151 (N_13151,N_12257,N_12769);
and U13152 (N_13152,N_12677,N_12095);
nor U13153 (N_13153,N_12117,N_12268);
and U13154 (N_13154,N_12294,N_12474);
xor U13155 (N_13155,N_12832,N_12997);
nor U13156 (N_13156,N_12330,N_12134);
nand U13157 (N_13157,N_12937,N_12043);
and U13158 (N_13158,N_12311,N_12826);
nor U13159 (N_13159,N_12952,N_12393);
and U13160 (N_13160,N_12720,N_12327);
nand U13161 (N_13161,N_12108,N_12676);
and U13162 (N_13162,N_12706,N_12229);
nor U13163 (N_13163,N_12886,N_12625);
and U13164 (N_13164,N_12303,N_12556);
and U13165 (N_13165,N_12116,N_12705);
nand U13166 (N_13166,N_12237,N_12511);
nand U13167 (N_13167,N_12172,N_12999);
or U13168 (N_13168,N_12000,N_12346);
or U13169 (N_13169,N_12421,N_12692);
and U13170 (N_13170,N_12409,N_12517);
or U13171 (N_13171,N_12920,N_12368);
and U13172 (N_13172,N_12550,N_12286);
or U13173 (N_13173,N_12441,N_12492);
nor U13174 (N_13174,N_12058,N_12288);
nand U13175 (N_13175,N_12535,N_12196);
xor U13176 (N_13176,N_12064,N_12910);
or U13177 (N_13177,N_12369,N_12739);
nor U13178 (N_13178,N_12126,N_12529);
and U13179 (N_13179,N_12044,N_12657);
xor U13180 (N_13180,N_12956,N_12233);
nand U13181 (N_13181,N_12282,N_12656);
or U13182 (N_13182,N_12591,N_12079);
and U13183 (N_13183,N_12785,N_12198);
xnor U13184 (N_13184,N_12080,N_12849);
or U13185 (N_13185,N_12979,N_12827);
and U13186 (N_13186,N_12987,N_12228);
or U13187 (N_13187,N_12506,N_12762);
nor U13188 (N_13188,N_12312,N_12766);
nand U13189 (N_13189,N_12410,N_12142);
or U13190 (N_13190,N_12883,N_12823);
nand U13191 (N_13191,N_12467,N_12260);
and U13192 (N_13192,N_12545,N_12355);
or U13193 (N_13193,N_12465,N_12949);
nand U13194 (N_13194,N_12348,N_12940);
xnor U13195 (N_13195,N_12615,N_12463);
and U13196 (N_13196,N_12774,N_12622);
nand U13197 (N_13197,N_12442,N_12893);
nor U13198 (N_13198,N_12357,N_12637);
nor U13199 (N_13199,N_12293,N_12755);
and U13200 (N_13200,N_12460,N_12682);
nor U13201 (N_13201,N_12938,N_12400);
nor U13202 (N_13202,N_12436,N_12109);
xor U13203 (N_13203,N_12604,N_12642);
nand U13204 (N_13204,N_12630,N_12750);
and U13205 (N_13205,N_12349,N_12598);
xnor U13206 (N_13206,N_12070,N_12819);
nand U13207 (N_13207,N_12017,N_12559);
xnor U13208 (N_13208,N_12322,N_12592);
xnor U13209 (N_13209,N_12847,N_12691);
nand U13210 (N_13210,N_12699,N_12124);
nor U13211 (N_13211,N_12156,N_12335);
xnor U13212 (N_13212,N_12961,N_12932);
nand U13213 (N_13213,N_12845,N_12812);
nor U13214 (N_13214,N_12232,N_12673);
xor U13215 (N_13215,N_12008,N_12572);
xnor U13216 (N_13216,N_12745,N_12160);
and U13217 (N_13217,N_12548,N_12996);
and U13218 (N_13218,N_12281,N_12912);
and U13219 (N_13219,N_12605,N_12476);
nor U13220 (N_13220,N_12053,N_12607);
or U13221 (N_13221,N_12226,N_12390);
nor U13222 (N_13222,N_12791,N_12830);
nand U13223 (N_13223,N_12628,N_12544);
or U13224 (N_13224,N_12754,N_12149);
and U13225 (N_13225,N_12038,N_12181);
nand U13226 (N_13226,N_12003,N_12732);
nor U13227 (N_13227,N_12265,N_12837);
nor U13228 (N_13228,N_12722,N_12613);
xor U13229 (N_13229,N_12122,N_12331);
or U13230 (N_13230,N_12143,N_12332);
xor U13231 (N_13231,N_12551,N_12752);
and U13232 (N_13232,N_12738,N_12553);
xor U13233 (N_13233,N_12963,N_12120);
nor U13234 (N_13234,N_12685,N_12169);
or U13235 (N_13235,N_12659,N_12890);
and U13236 (N_13236,N_12168,N_12509);
nand U13237 (N_13237,N_12151,N_12416);
nand U13238 (N_13238,N_12206,N_12015);
nand U13239 (N_13239,N_12925,N_12171);
and U13240 (N_13240,N_12564,N_12859);
or U13241 (N_13241,N_12709,N_12675);
nor U13242 (N_13242,N_12479,N_12627);
nor U13243 (N_13243,N_12101,N_12895);
nor U13244 (N_13244,N_12765,N_12023);
xor U13245 (N_13245,N_12193,N_12581);
nand U13246 (N_13246,N_12510,N_12967);
xnor U13247 (N_13247,N_12068,N_12300);
and U13248 (N_13248,N_12927,N_12662);
and U13249 (N_13249,N_12816,N_12475);
and U13250 (N_13250,N_12945,N_12687);
xnor U13251 (N_13251,N_12497,N_12631);
or U13252 (N_13252,N_12879,N_12661);
and U13253 (N_13253,N_12702,N_12121);
nand U13254 (N_13254,N_12980,N_12679);
xnor U13255 (N_13255,N_12670,N_12939);
or U13256 (N_13256,N_12316,N_12114);
nand U13257 (N_13257,N_12305,N_12194);
nand U13258 (N_13258,N_12841,N_12577);
or U13259 (N_13259,N_12955,N_12457);
nand U13260 (N_13260,N_12777,N_12640);
xor U13261 (N_13261,N_12536,N_12417);
and U13262 (N_13262,N_12005,N_12907);
or U13263 (N_13263,N_12273,N_12526);
and U13264 (N_13264,N_12432,N_12252);
nor U13265 (N_13265,N_12420,N_12150);
xor U13266 (N_13266,N_12494,N_12319);
nor U13267 (N_13267,N_12606,N_12251);
or U13268 (N_13268,N_12825,N_12527);
nand U13269 (N_13269,N_12962,N_12668);
nand U13270 (N_13270,N_12431,N_12188);
xnor U13271 (N_13271,N_12345,N_12182);
xor U13272 (N_13272,N_12864,N_12209);
nand U13273 (N_13273,N_12666,N_12063);
and U13274 (N_13274,N_12909,N_12946);
xnor U13275 (N_13275,N_12230,N_12065);
or U13276 (N_13276,N_12950,N_12507);
nor U13277 (N_13277,N_12173,N_12994);
and U13278 (N_13278,N_12414,N_12029);
nand U13279 (N_13279,N_12768,N_12834);
nor U13280 (N_13280,N_12050,N_12824);
and U13281 (N_13281,N_12835,N_12934);
nand U13282 (N_13282,N_12344,N_12267);
nor U13283 (N_13283,N_12704,N_12970);
and U13284 (N_13284,N_12262,N_12609);
nand U13285 (N_13285,N_12175,N_12897);
and U13286 (N_13286,N_12696,N_12874);
nand U13287 (N_13287,N_12638,N_12006);
xor U13288 (N_13288,N_12531,N_12680);
nand U13289 (N_13289,N_12115,N_12549);
or U13290 (N_13290,N_12795,N_12842);
and U13291 (N_13291,N_12089,N_12872);
nor U13292 (N_13292,N_12876,N_12090);
xnor U13293 (N_13293,N_12714,N_12304);
nand U13294 (N_13294,N_12792,N_12567);
or U13295 (N_13295,N_12797,N_12046);
or U13296 (N_13296,N_12165,N_12590);
nor U13297 (N_13297,N_12222,N_12737);
or U13298 (N_13298,N_12902,N_12936);
or U13299 (N_13299,N_12983,N_12878);
nand U13300 (N_13300,N_12013,N_12025);
or U13301 (N_13301,N_12350,N_12660);
or U13302 (N_13302,N_12381,N_12195);
nand U13303 (N_13303,N_12593,N_12958);
and U13304 (N_13304,N_12575,N_12543);
or U13305 (N_13305,N_12608,N_12047);
nor U13306 (N_13306,N_12133,N_12433);
xor U13307 (N_13307,N_12179,N_12402);
nor U13308 (N_13308,N_12405,N_12986);
nor U13309 (N_13309,N_12287,N_12802);
nor U13310 (N_13310,N_12846,N_12921);
nor U13311 (N_13311,N_12782,N_12853);
nor U13312 (N_13312,N_12084,N_12486);
xor U13313 (N_13313,N_12935,N_12309);
nor U13314 (N_13314,N_12663,N_12191);
xor U13315 (N_13315,N_12127,N_12582);
and U13316 (N_13316,N_12848,N_12905);
nand U13317 (N_13317,N_12202,N_12024);
or U13318 (N_13318,N_12784,N_12277);
xnor U13319 (N_13319,N_12681,N_12941);
nor U13320 (N_13320,N_12091,N_12944);
and U13321 (N_13321,N_12746,N_12576);
xor U13322 (N_13322,N_12401,N_12500);
xnor U13323 (N_13323,N_12081,N_12563);
xnor U13324 (N_13324,N_12470,N_12723);
nand U13325 (N_13325,N_12915,N_12379);
or U13326 (N_13326,N_12413,N_12993);
xnor U13327 (N_13327,N_12557,N_12419);
nor U13328 (N_13328,N_12270,N_12977);
or U13329 (N_13329,N_12096,N_12542);
and U13330 (N_13330,N_12984,N_12033);
nand U13331 (N_13331,N_12343,N_12026);
and U13332 (N_13332,N_12450,N_12541);
xnor U13333 (N_13333,N_12743,N_12957);
nand U13334 (N_13334,N_12034,N_12204);
nor U13335 (N_13335,N_12854,N_12395);
nand U13336 (N_13336,N_12995,N_12726);
nor U13337 (N_13337,N_12756,N_12464);
or U13338 (N_13338,N_12533,N_12221);
nand U13339 (N_13339,N_12424,N_12049);
or U13340 (N_13340,N_12295,N_12913);
or U13341 (N_13341,N_12683,N_12528);
nor U13342 (N_13342,N_12882,N_12250);
nand U13343 (N_13343,N_12103,N_12788);
nand U13344 (N_13344,N_12211,N_12366);
and U13345 (N_13345,N_12796,N_12248);
and U13346 (N_13346,N_12130,N_12719);
nand U13347 (N_13347,N_12220,N_12138);
nand U13348 (N_13348,N_12341,N_12943);
nand U13349 (N_13349,N_12094,N_12459);
or U13350 (N_13350,N_12742,N_12786);
or U13351 (N_13351,N_12186,N_12054);
nand U13352 (N_13352,N_12580,N_12727);
or U13353 (N_13353,N_12900,N_12111);
or U13354 (N_13354,N_12851,N_12451);
xor U13355 (N_13355,N_12042,N_12904);
xnor U13356 (N_13356,N_12868,N_12973);
and U13357 (N_13357,N_12391,N_12066);
nor U13358 (N_13358,N_12991,N_12870);
xnor U13359 (N_13359,N_12241,N_12364);
nand U13360 (N_13360,N_12462,N_12713);
xnor U13361 (N_13361,N_12461,N_12783);
nor U13362 (N_13362,N_12161,N_12170);
nand U13363 (N_13363,N_12678,N_12174);
xor U13364 (N_13364,N_12444,N_12135);
nor U13365 (N_13365,N_12763,N_12585);
nor U13366 (N_13366,N_12885,N_12011);
and U13367 (N_13367,N_12807,N_12843);
xnor U13368 (N_13368,N_12212,N_12712);
and U13369 (N_13369,N_12574,N_12388);
xor U13370 (N_13370,N_12612,N_12554);
or U13371 (N_13371,N_12059,N_12314);
or U13372 (N_13372,N_12396,N_12306);
and U13373 (N_13373,N_12562,N_12446);
or U13374 (N_13374,N_12342,N_12707);
xnor U13375 (N_13375,N_12881,N_12406);
and U13376 (N_13376,N_12674,N_12208);
nor U13377 (N_13377,N_12069,N_12398);
xnor U13378 (N_13378,N_12238,N_12100);
or U13379 (N_13379,N_12320,N_12569);
and U13380 (N_13380,N_12118,N_12256);
nor U13381 (N_13381,N_12159,N_12588);
and U13382 (N_13382,N_12020,N_12352);
xor U13383 (N_13383,N_12190,N_12073);
xor U13384 (N_13384,N_12275,N_12751);
xnor U13385 (N_13385,N_12652,N_12695);
and U13386 (N_13386,N_12057,N_12579);
nor U13387 (N_13387,N_12658,N_12811);
or U13388 (N_13388,N_12534,N_12099);
nand U13389 (N_13389,N_12027,N_12167);
nor U13390 (N_13390,N_12914,N_12429);
xor U13391 (N_13391,N_12601,N_12621);
or U13392 (N_13392,N_12926,N_12561);
nand U13393 (N_13393,N_12082,N_12269);
nor U13394 (N_13394,N_12480,N_12693);
nor U13395 (N_13395,N_12725,N_12798);
or U13396 (N_13396,N_12587,N_12884);
xor U13397 (N_13397,N_12323,N_12374);
xnor U13398 (N_13398,N_12933,N_12105);
or U13399 (N_13399,N_12310,N_12261);
or U13400 (N_13400,N_12758,N_12515);
and U13401 (N_13401,N_12426,N_12407);
nor U13402 (N_13402,N_12007,N_12482);
nor U13403 (N_13403,N_12650,N_12239);
nand U13404 (N_13404,N_12833,N_12338);
xnor U13405 (N_13405,N_12164,N_12427);
and U13406 (N_13406,N_12491,N_12136);
xnor U13407 (N_13407,N_12362,N_12908);
and U13408 (N_13408,N_12665,N_12803);
nand U13409 (N_13409,N_12817,N_12778);
nor U13410 (N_13410,N_12801,N_12297);
or U13411 (N_13411,N_12635,N_12308);
or U13412 (N_13412,N_12787,N_12358);
nand U13413 (N_13413,N_12948,N_12888);
or U13414 (N_13414,N_12039,N_12747);
nor U13415 (N_13415,N_12456,N_12018);
xor U13416 (N_13416,N_12923,N_12141);
nand U13417 (N_13417,N_12112,N_12224);
xor U13418 (N_13418,N_12152,N_12307);
xor U13419 (N_13419,N_12040,N_12602);
nand U13420 (N_13420,N_12272,N_12113);
xnor U13421 (N_13421,N_12960,N_12988);
and U13422 (N_13422,N_12898,N_12210);
nor U13423 (N_13423,N_12128,N_12361);
nand U13424 (N_13424,N_12385,N_12037);
and U13425 (N_13425,N_12499,N_12428);
or U13426 (N_13426,N_12197,N_12809);
and U13427 (N_13427,N_12969,N_12439);
nor U13428 (N_13428,N_12850,N_12484);
nor U13429 (N_13429,N_12283,N_12776);
nor U13430 (N_13430,N_12060,N_12276);
nor U13431 (N_13431,N_12137,N_12740);
nand U13432 (N_13432,N_12279,N_12822);
xnor U13433 (N_13433,N_12110,N_12611);
nor U13434 (N_13434,N_12653,N_12584);
nand U13435 (N_13435,N_12974,N_12085);
nand U13436 (N_13436,N_12002,N_12375);
xor U13437 (N_13437,N_12473,N_12148);
or U13438 (N_13438,N_12157,N_12411);
and U13439 (N_13439,N_12016,N_12689);
and U13440 (N_13440,N_12671,N_12041);
nor U13441 (N_13441,N_12030,N_12976);
nor U13442 (N_13442,N_12386,N_12964);
and U13443 (N_13443,N_12645,N_12716);
nand U13444 (N_13444,N_12775,N_12839);
and U13445 (N_13445,N_12998,N_12012);
nand U13446 (N_13446,N_12201,N_12759);
xor U13447 (N_13447,N_12129,N_12317);
nand U13448 (N_13448,N_12530,N_12032);
and U13449 (N_13449,N_12438,N_12931);
nand U13450 (N_13450,N_12684,N_12753);
xor U13451 (N_13451,N_12125,N_12075);
nand U13452 (N_13452,N_12363,N_12278);
nor U13453 (N_13453,N_12437,N_12185);
and U13454 (N_13454,N_12236,N_12291);
nor U13455 (N_13455,N_12302,N_12501);
xnor U13456 (N_13456,N_12953,N_12733);
xor U13457 (N_13457,N_12546,N_12856);
nand U13458 (N_13458,N_12570,N_12045);
xnor U13459 (N_13459,N_12617,N_12351);
and U13460 (N_13460,N_12599,N_12153);
nor U13461 (N_13461,N_12818,N_12454);
nor U13462 (N_13462,N_12589,N_12648);
nand U13463 (N_13463,N_12477,N_12321);
nand U13464 (N_13464,N_12836,N_12061);
or U13465 (N_13465,N_12871,N_12326);
and U13466 (N_13466,N_12423,N_12489);
nor U13467 (N_13467,N_12855,N_12793);
nand U13468 (N_13468,N_12654,N_12086);
and U13469 (N_13469,N_12487,N_12831);
nor U13470 (N_13470,N_12056,N_12813);
nand U13471 (N_13471,N_12478,N_12455);
and U13472 (N_13472,N_12384,N_12647);
nand U13473 (N_13473,N_12468,N_12772);
nor U13474 (N_13474,N_12717,N_12301);
nand U13475 (N_13475,N_12538,N_12072);
nand U13476 (N_13476,N_12971,N_12339);
nand U13477 (N_13477,N_12106,N_12686);
xor U13478 (N_13478,N_12698,N_12242);
nor U13479 (N_13479,N_12804,N_12353);
or U13480 (N_13480,N_12764,N_12458);
nand U13481 (N_13481,N_12067,N_12422);
nand U13482 (N_13482,N_12337,N_12789);
xor U13483 (N_13483,N_12215,N_12873);
nand U13484 (N_13484,N_12010,N_12975);
nand U13485 (N_13485,N_12600,N_12187);
nor U13486 (N_13486,N_12688,N_12810);
xnor U13487 (N_13487,N_12123,N_12022);
and U13488 (N_13488,N_12399,N_12620);
and U13489 (N_13489,N_12325,N_12271);
nand U13490 (N_13490,N_12154,N_12028);
xor U13491 (N_13491,N_12290,N_12207);
xnor U13492 (N_13492,N_12249,N_12595);
or U13493 (N_13493,N_12102,N_12107);
xor U13494 (N_13494,N_12336,N_12180);
or U13495 (N_13495,N_12649,N_12728);
and U13496 (N_13496,N_12051,N_12244);
and U13497 (N_13497,N_12639,N_12571);
xnor U13498 (N_13498,N_12521,N_12636);
nor U13499 (N_13499,N_12518,N_12911);
and U13500 (N_13500,N_12643,N_12965);
nand U13501 (N_13501,N_12047,N_12669);
xnor U13502 (N_13502,N_12360,N_12181);
nand U13503 (N_13503,N_12069,N_12407);
and U13504 (N_13504,N_12976,N_12367);
xnor U13505 (N_13505,N_12392,N_12590);
nor U13506 (N_13506,N_12576,N_12100);
and U13507 (N_13507,N_12938,N_12806);
nand U13508 (N_13508,N_12262,N_12309);
xnor U13509 (N_13509,N_12244,N_12321);
and U13510 (N_13510,N_12030,N_12357);
xnor U13511 (N_13511,N_12303,N_12136);
nand U13512 (N_13512,N_12696,N_12653);
nand U13513 (N_13513,N_12553,N_12113);
nand U13514 (N_13514,N_12016,N_12609);
nand U13515 (N_13515,N_12289,N_12769);
nor U13516 (N_13516,N_12226,N_12964);
or U13517 (N_13517,N_12996,N_12853);
nand U13518 (N_13518,N_12067,N_12650);
or U13519 (N_13519,N_12277,N_12857);
or U13520 (N_13520,N_12276,N_12048);
or U13521 (N_13521,N_12797,N_12372);
nor U13522 (N_13522,N_12461,N_12173);
and U13523 (N_13523,N_12621,N_12768);
nand U13524 (N_13524,N_12535,N_12991);
nand U13525 (N_13525,N_12642,N_12323);
and U13526 (N_13526,N_12712,N_12742);
nor U13527 (N_13527,N_12021,N_12282);
and U13528 (N_13528,N_12271,N_12962);
xnor U13529 (N_13529,N_12304,N_12488);
xor U13530 (N_13530,N_12941,N_12371);
xor U13531 (N_13531,N_12657,N_12679);
nand U13532 (N_13532,N_12244,N_12086);
or U13533 (N_13533,N_12079,N_12050);
xor U13534 (N_13534,N_12844,N_12465);
and U13535 (N_13535,N_12358,N_12813);
and U13536 (N_13536,N_12939,N_12796);
nor U13537 (N_13537,N_12890,N_12232);
xnor U13538 (N_13538,N_12838,N_12058);
xnor U13539 (N_13539,N_12773,N_12096);
xor U13540 (N_13540,N_12954,N_12610);
nand U13541 (N_13541,N_12481,N_12836);
or U13542 (N_13542,N_12659,N_12122);
nor U13543 (N_13543,N_12592,N_12685);
and U13544 (N_13544,N_12434,N_12651);
or U13545 (N_13545,N_12427,N_12053);
or U13546 (N_13546,N_12865,N_12184);
and U13547 (N_13547,N_12815,N_12401);
xor U13548 (N_13548,N_12072,N_12415);
or U13549 (N_13549,N_12127,N_12675);
nor U13550 (N_13550,N_12644,N_12285);
xnor U13551 (N_13551,N_12466,N_12693);
nor U13552 (N_13552,N_12460,N_12929);
xor U13553 (N_13553,N_12598,N_12344);
xnor U13554 (N_13554,N_12892,N_12127);
or U13555 (N_13555,N_12012,N_12569);
nor U13556 (N_13556,N_12385,N_12394);
or U13557 (N_13557,N_12957,N_12424);
or U13558 (N_13558,N_12354,N_12975);
nand U13559 (N_13559,N_12080,N_12496);
and U13560 (N_13560,N_12688,N_12377);
nand U13561 (N_13561,N_12816,N_12588);
nand U13562 (N_13562,N_12188,N_12054);
and U13563 (N_13563,N_12475,N_12476);
xor U13564 (N_13564,N_12275,N_12916);
nand U13565 (N_13565,N_12727,N_12735);
or U13566 (N_13566,N_12088,N_12859);
nor U13567 (N_13567,N_12084,N_12078);
xnor U13568 (N_13568,N_12975,N_12884);
or U13569 (N_13569,N_12964,N_12069);
nand U13570 (N_13570,N_12340,N_12578);
nor U13571 (N_13571,N_12603,N_12148);
nand U13572 (N_13572,N_12491,N_12433);
xnor U13573 (N_13573,N_12905,N_12011);
nor U13574 (N_13574,N_12122,N_12181);
nand U13575 (N_13575,N_12503,N_12125);
and U13576 (N_13576,N_12921,N_12259);
or U13577 (N_13577,N_12287,N_12087);
xor U13578 (N_13578,N_12255,N_12312);
xnor U13579 (N_13579,N_12815,N_12855);
nand U13580 (N_13580,N_12845,N_12758);
or U13581 (N_13581,N_12133,N_12753);
nand U13582 (N_13582,N_12293,N_12467);
and U13583 (N_13583,N_12177,N_12570);
xnor U13584 (N_13584,N_12037,N_12211);
xnor U13585 (N_13585,N_12964,N_12584);
or U13586 (N_13586,N_12571,N_12403);
xor U13587 (N_13587,N_12992,N_12505);
nand U13588 (N_13588,N_12119,N_12949);
or U13589 (N_13589,N_12324,N_12445);
and U13590 (N_13590,N_12845,N_12458);
xnor U13591 (N_13591,N_12614,N_12625);
nor U13592 (N_13592,N_12627,N_12510);
or U13593 (N_13593,N_12964,N_12982);
and U13594 (N_13594,N_12751,N_12774);
nor U13595 (N_13595,N_12651,N_12649);
and U13596 (N_13596,N_12803,N_12946);
and U13597 (N_13597,N_12225,N_12141);
and U13598 (N_13598,N_12298,N_12856);
nand U13599 (N_13599,N_12754,N_12352);
nor U13600 (N_13600,N_12054,N_12472);
nand U13601 (N_13601,N_12053,N_12836);
or U13602 (N_13602,N_12521,N_12019);
nor U13603 (N_13603,N_12880,N_12941);
xor U13604 (N_13604,N_12235,N_12083);
and U13605 (N_13605,N_12523,N_12117);
and U13606 (N_13606,N_12297,N_12060);
xor U13607 (N_13607,N_12592,N_12891);
nor U13608 (N_13608,N_12865,N_12428);
or U13609 (N_13609,N_12348,N_12079);
nor U13610 (N_13610,N_12955,N_12705);
or U13611 (N_13611,N_12493,N_12591);
nor U13612 (N_13612,N_12767,N_12150);
and U13613 (N_13613,N_12271,N_12544);
or U13614 (N_13614,N_12438,N_12869);
nand U13615 (N_13615,N_12757,N_12738);
nand U13616 (N_13616,N_12203,N_12506);
or U13617 (N_13617,N_12479,N_12894);
and U13618 (N_13618,N_12364,N_12612);
nand U13619 (N_13619,N_12926,N_12885);
and U13620 (N_13620,N_12577,N_12217);
and U13621 (N_13621,N_12980,N_12968);
nand U13622 (N_13622,N_12182,N_12636);
or U13623 (N_13623,N_12726,N_12171);
or U13624 (N_13624,N_12001,N_12906);
xor U13625 (N_13625,N_12097,N_12914);
nor U13626 (N_13626,N_12596,N_12327);
xor U13627 (N_13627,N_12913,N_12398);
nor U13628 (N_13628,N_12199,N_12605);
or U13629 (N_13629,N_12541,N_12830);
nor U13630 (N_13630,N_12866,N_12506);
and U13631 (N_13631,N_12946,N_12301);
nand U13632 (N_13632,N_12516,N_12975);
nor U13633 (N_13633,N_12310,N_12720);
and U13634 (N_13634,N_12558,N_12117);
or U13635 (N_13635,N_12866,N_12121);
xnor U13636 (N_13636,N_12347,N_12190);
nor U13637 (N_13637,N_12361,N_12494);
or U13638 (N_13638,N_12788,N_12598);
xnor U13639 (N_13639,N_12458,N_12838);
nor U13640 (N_13640,N_12065,N_12487);
and U13641 (N_13641,N_12459,N_12196);
or U13642 (N_13642,N_12914,N_12795);
or U13643 (N_13643,N_12329,N_12264);
nand U13644 (N_13644,N_12709,N_12972);
nand U13645 (N_13645,N_12854,N_12118);
and U13646 (N_13646,N_12674,N_12929);
nor U13647 (N_13647,N_12981,N_12075);
and U13648 (N_13648,N_12608,N_12170);
nor U13649 (N_13649,N_12074,N_12265);
xor U13650 (N_13650,N_12317,N_12689);
nand U13651 (N_13651,N_12238,N_12602);
or U13652 (N_13652,N_12322,N_12043);
xor U13653 (N_13653,N_12470,N_12774);
or U13654 (N_13654,N_12501,N_12799);
nand U13655 (N_13655,N_12424,N_12563);
or U13656 (N_13656,N_12364,N_12222);
xor U13657 (N_13657,N_12106,N_12469);
nor U13658 (N_13658,N_12812,N_12816);
xor U13659 (N_13659,N_12312,N_12377);
nand U13660 (N_13660,N_12176,N_12873);
xor U13661 (N_13661,N_12565,N_12990);
or U13662 (N_13662,N_12004,N_12916);
or U13663 (N_13663,N_12420,N_12895);
xnor U13664 (N_13664,N_12135,N_12026);
nand U13665 (N_13665,N_12163,N_12453);
xor U13666 (N_13666,N_12336,N_12926);
and U13667 (N_13667,N_12511,N_12313);
and U13668 (N_13668,N_12077,N_12992);
or U13669 (N_13669,N_12743,N_12072);
and U13670 (N_13670,N_12516,N_12050);
nand U13671 (N_13671,N_12569,N_12586);
xnor U13672 (N_13672,N_12936,N_12376);
or U13673 (N_13673,N_12298,N_12349);
or U13674 (N_13674,N_12506,N_12164);
or U13675 (N_13675,N_12707,N_12547);
or U13676 (N_13676,N_12075,N_12666);
or U13677 (N_13677,N_12258,N_12445);
or U13678 (N_13678,N_12210,N_12453);
xor U13679 (N_13679,N_12439,N_12728);
nor U13680 (N_13680,N_12616,N_12309);
and U13681 (N_13681,N_12247,N_12587);
or U13682 (N_13682,N_12574,N_12139);
nand U13683 (N_13683,N_12646,N_12834);
xnor U13684 (N_13684,N_12370,N_12577);
and U13685 (N_13685,N_12244,N_12805);
nor U13686 (N_13686,N_12193,N_12340);
nand U13687 (N_13687,N_12923,N_12482);
nor U13688 (N_13688,N_12341,N_12821);
xnor U13689 (N_13689,N_12159,N_12257);
and U13690 (N_13690,N_12291,N_12986);
nand U13691 (N_13691,N_12040,N_12107);
nand U13692 (N_13692,N_12648,N_12965);
and U13693 (N_13693,N_12085,N_12292);
xnor U13694 (N_13694,N_12613,N_12653);
nand U13695 (N_13695,N_12224,N_12416);
and U13696 (N_13696,N_12550,N_12821);
or U13697 (N_13697,N_12068,N_12588);
or U13698 (N_13698,N_12175,N_12308);
or U13699 (N_13699,N_12554,N_12863);
nor U13700 (N_13700,N_12476,N_12997);
xnor U13701 (N_13701,N_12988,N_12340);
nor U13702 (N_13702,N_12941,N_12088);
xnor U13703 (N_13703,N_12997,N_12840);
and U13704 (N_13704,N_12989,N_12929);
xor U13705 (N_13705,N_12321,N_12334);
nand U13706 (N_13706,N_12019,N_12495);
xor U13707 (N_13707,N_12496,N_12145);
nor U13708 (N_13708,N_12101,N_12847);
nand U13709 (N_13709,N_12301,N_12860);
nor U13710 (N_13710,N_12383,N_12717);
and U13711 (N_13711,N_12563,N_12979);
nor U13712 (N_13712,N_12658,N_12210);
and U13713 (N_13713,N_12897,N_12737);
and U13714 (N_13714,N_12381,N_12221);
nand U13715 (N_13715,N_12686,N_12013);
or U13716 (N_13716,N_12065,N_12866);
xnor U13717 (N_13717,N_12407,N_12024);
or U13718 (N_13718,N_12303,N_12954);
and U13719 (N_13719,N_12540,N_12762);
nor U13720 (N_13720,N_12554,N_12261);
nand U13721 (N_13721,N_12680,N_12523);
xnor U13722 (N_13722,N_12620,N_12157);
and U13723 (N_13723,N_12159,N_12437);
nor U13724 (N_13724,N_12221,N_12879);
xor U13725 (N_13725,N_12384,N_12938);
xnor U13726 (N_13726,N_12036,N_12712);
nor U13727 (N_13727,N_12746,N_12531);
nor U13728 (N_13728,N_12191,N_12835);
and U13729 (N_13729,N_12226,N_12473);
nor U13730 (N_13730,N_12586,N_12101);
xor U13731 (N_13731,N_12016,N_12282);
nand U13732 (N_13732,N_12595,N_12978);
xnor U13733 (N_13733,N_12120,N_12116);
nand U13734 (N_13734,N_12461,N_12635);
xnor U13735 (N_13735,N_12963,N_12513);
nand U13736 (N_13736,N_12885,N_12107);
nand U13737 (N_13737,N_12336,N_12133);
nand U13738 (N_13738,N_12034,N_12839);
or U13739 (N_13739,N_12814,N_12265);
xor U13740 (N_13740,N_12844,N_12845);
or U13741 (N_13741,N_12050,N_12828);
xnor U13742 (N_13742,N_12449,N_12161);
and U13743 (N_13743,N_12647,N_12827);
nor U13744 (N_13744,N_12539,N_12574);
xnor U13745 (N_13745,N_12265,N_12897);
nor U13746 (N_13746,N_12325,N_12784);
and U13747 (N_13747,N_12217,N_12442);
nor U13748 (N_13748,N_12282,N_12558);
xor U13749 (N_13749,N_12662,N_12995);
nor U13750 (N_13750,N_12049,N_12111);
nor U13751 (N_13751,N_12064,N_12656);
xor U13752 (N_13752,N_12871,N_12434);
nor U13753 (N_13753,N_12079,N_12795);
xor U13754 (N_13754,N_12917,N_12747);
or U13755 (N_13755,N_12927,N_12120);
xor U13756 (N_13756,N_12094,N_12331);
or U13757 (N_13757,N_12258,N_12839);
and U13758 (N_13758,N_12629,N_12210);
and U13759 (N_13759,N_12790,N_12606);
nor U13760 (N_13760,N_12710,N_12465);
nand U13761 (N_13761,N_12087,N_12231);
and U13762 (N_13762,N_12340,N_12861);
nor U13763 (N_13763,N_12035,N_12506);
or U13764 (N_13764,N_12931,N_12570);
and U13765 (N_13765,N_12978,N_12942);
nand U13766 (N_13766,N_12093,N_12018);
xnor U13767 (N_13767,N_12352,N_12912);
and U13768 (N_13768,N_12641,N_12667);
nand U13769 (N_13769,N_12949,N_12381);
nor U13770 (N_13770,N_12853,N_12162);
or U13771 (N_13771,N_12304,N_12835);
or U13772 (N_13772,N_12759,N_12181);
nand U13773 (N_13773,N_12051,N_12667);
nor U13774 (N_13774,N_12186,N_12816);
or U13775 (N_13775,N_12912,N_12670);
and U13776 (N_13776,N_12457,N_12291);
xor U13777 (N_13777,N_12267,N_12778);
xnor U13778 (N_13778,N_12444,N_12611);
xor U13779 (N_13779,N_12811,N_12415);
nand U13780 (N_13780,N_12335,N_12348);
nand U13781 (N_13781,N_12315,N_12926);
nor U13782 (N_13782,N_12486,N_12303);
or U13783 (N_13783,N_12926,N_12239);
xor U13784 (N_13784,N_12864,N_12525);
and U13785 (N_13785,N_12545,N_12713);
nand U13786 (N_13786,N_12283,N_12372);
xnor U13787 (N_13787,N_12933,N_12905);
xor U13788 (N_13788,N_12589,N_12847);
nand U13789 (N_13789,N_12320,N_12718);
and U13790 (N_13790,N_12894,N_12078);
or U13791 (N_13791,N_12017,N_12081);
nand U13792 (N_13792,N_12269,N_12605);
xnor U13793 (N_13793,N_12887,N_12018);
and U13794 (N_13794,N_12066,N_12099);
or U13795 (N_13795,N_12867,N_12654);
nor U13796 (N_13796,N_12772,N_12729);
xnor U13797 (N_13797,N_12684,N_12316);
or U13798 (N_13798,N_12494,N_12644);
xnor U13799 (N_13799,N_12195,N_12021);
nor U13800 (N_13800,N_12163,N_12234);
nor U13801 (N_13801,N_12784,N_12247);
or U13802 (N_13802,N_12542,N_12373);
nor U13803 (N_13803,N_12675,N_12557);
nor U13804 (N_13804,N_12185,N_12862);
xor U13805 (N_13805,N_12369,N_12455);
nor U13806 (N_13806,N_12614,N_12150);
xnor U13807 (N_13807,N_12477,N_12139);
and U13808 (N_13808,N_12350,N_12414);
nor U13809 (N_13809,N_12232,N_12563);
nor U13810 (N_13810,N_12163,N_12089);
or U13811 (N_13811,N_12702,N_12893);
nand U13812 (N_13812,N_12978,N_12702);
or U13813 (N_13813,N_12294,N_12431);
xnor U13814 (N_13814,N_12086,N_12401);
or U13815 (N_13815,N_12324,N_12543);
nand U13816 (N_13816,N_12566,N_12039);
xnor U13817 (N_13817,N_12647,N_12691);
nor U13818 (N_13818,N_12458,N_12724);
nand U13819 (N_13819,N_12834,N_12949);
xor U13820 (N_13820,N_12779,N_12554);
nand U13821 (N_13821,N_12608,N_12931);
or U13822 (N_13822,N_12920,N_12247);
xnor U13823 (N_13823,N_12059,N_12317);
xor U13824 (N_13824,N_12314,N_12762);
xnor U13825 (N_13825,N_12675,N_12954);
and U13826 (N_13826,N_12493,N_12660);
nor U13827 (N_13827,N_12254,N_12776);
nand U13828 (N_13828,N_12254,N_12954);
nand U13829 (N_13829,N_12389,N_12850);
xnor U13830 (N_13830,N_12656,N_12722);
or U13831 (N_13831,N_12049,N_12377);
nor U13832 (N_13832,N_12167,N_12227);
nor U13833 (N_13833,N_12229,N_12634);
xnor U13834 (N_13834,N_12114,N_12058);
xnor U13835 (N_13835,N_12680,N_12136);
or U13836 (N_13836,N_12663,N_12080);
and U13837 (N_13837,N_12832,N_12525);
xnor U13838 (N_13838,N_12293,N_12340);
or U13839 (N_13839,N_12831,N_12467);
nand U13840 (N_13840,N_12597,N_12588);
nor U13841 (N_13841,N_12349,N_12002);
or U13842 (N_13842,N_12401,N_12855);
nor U13843 (N_13843,N_12438,N_12652);
nand U13844 (N_13844,N_12475,N_12759);
nand U13845 (N_13845,N_12057,N_12570);
xnor U13846 (N_13846,N_12607,N_12394);
xor U13847 (N_13847,N_12206,N_12957);
xnor U13848 (N_13848,N_12988,N_12266);
or U13849 (N_13849,N_12628,N_12209);
nor U13850 (N_13850,N_12507,N_12067);
xnor U13851 (N_13851,N_12570,N_12980);
or U13852 (N_13852,N_12898,N_12851);
nor U13853 (N_13853,N_12346,N_12792);
nand U13854 (N_13854,N_12561,N_12372);
or U13855 (N_13855,N_12251,N_12977);
and U13856 (N_13856,N_12245,N_12385);
and U13857 (N_13857,N_12119,N_12705);
nor U13858 (N_13858,N_12822,N_12458);
and U13859 (N_13859,N_12933,N_12417);
nor U13860 (N_13860,N_12702,N_12452);
nand U13861 (N_13861,N_12353,N_12227);
nor U13862 (N_13862,N_12010,N_12599);
nor U13863 (N_13863,N_12057,N_12440);
nand U13864 (N_13864,N_12622,N_12215);
and U13865 (N_13865,N_12202,N_12337);
xnor U13866 (N_13866,N_12986,N_12579);
and U13867 (N_13867,N_12568,N_12059);
xnor U13868 (N_13868,N_12222,N_12903);
nor U13869 (N_13869,N_12056,N_12904);
nand U13870 (N_13870,N_12564,N_12672);
xor U13871 (N_13871,N_12673,N_12746);
nor U13872 (N_13872,N_12386,N_12123);
nor U13873 (N_13873,N_12688,N_12359);
nor U13874 (N_13874,N_12743,N_12399);
nor U13875 (N_13875,N_12891,N_12346);
nor U13876 (N_13876,N_12893,N_12846);
nand U13877 (N_13877,N_12318,N_12140);
or U13878 (N_13878,N_12740,N_12655);
nand U13879 (N_13879,N_12105,N_12538);
or U13880 (N_13880,N_12783,N_12248);
nand U13881 (N_13881,N_12265,N_12192);
nor U13882 (N_13882,N_12990,N_12240);
or U13883 (N_13883,N_12380,N_12670);
or U13884 (N_13884,N_12931,N_12493);
nand U13885 (N_13885,N_12525,N_12413);
nand U13886 (N_13886,N_12655,N_12335);
nand U13887 (N_13887,N_12223,N_12051);
nor U13888 (N_13888,N_12632,N_12957);
nor U13889 (N_13889,N_12235,N_12056);
or U13890 (N_13890,N_12550,N_12889);
xor U13891 (N_13891,N_12350,N_12788);
nor U13892 (N_13892,N_12767,N_12831);
or U13893 (N_13893,N_12388,N_12772);
nand U13894 (N_13894,N_12287,N_12117);
nor U13895 (N_13895,N_12988,N_12028);
nand U13896 (N_13896,N_12350,N_12134);
or U13897 (N_13897,N_12213,N_12110);
xnor U13898 (N_13898,N_12355,N_12207);
and U13899 (N_13899,N_12540,N_12714);
nor U13900 (N_13900,N_12533,N_12477);
or U13901 (N_13901,N_12240,N_12567);
xnor U13902 (N_13902,N_12367,N_12821);
or U13903 (N_13903,N_12505,N_12061);
nand U13904 (N_13904,N_12308,N_12531);
xnor U13905 (N_13905,N_12169,N_12036);
and U13906 (N_13906,N_12770,N_12734);
nor U13907 (N_13907,N_12827,N_12346);
nand U13908 (N_13908,N_12838,N_12234);
nand U13909 (N_13909,N_12077,N_12791);
nor U13910 (N_13910,N_12794,N_12671);
and U13911 (N_13911,N_12345,N_12303);
nand U13912 (N_13912,N_12855,N_12772);
or U13913 (N_13913,N_12623,N_12329);
xnor U13914 (N_13914,N_12705,N_12137);
or U13915 (N_13915,N_12132,N_12910);
and U13916 (N_13916,N_12099,N_12125);
nor U13917 (N_13917,N_12162,N_12387);
nor U13918 (N_13918,N_12556,N_12909);
nand U13919 (N_13919,N_12387,N_12946);
nand U13920 (N_13920,N_12279,N_12103);
xor U13921 (N_13921,N_12226,N_12530);
nor U13922 (N_13922,N_12449,N_12972);
xnor U13923 (N_13923,N_12112,N_12116);
xor U13924 (N_13924,N_12587,N_12314);
and U13925 (N_13925,N_12174,N_12049);
nor U13926 (N_13926,N_12359,N_12325);
nand U13927 (N_13927,N_12344,N_12708);
nand U13928 (N_13928,N_12333,N_12304);
and U13929 (N_13929,N_12006,N_12153);
xnor U13930 (N_13930,N_12403,N_12974);
xnor U13931 (N_13931,N_12474,N_12773);
nor U13932 (N_13932,N_12582,N_12456);
or U13933 (N_13933,N_12107,N_12938);
nand U13934 (N_13934,N_12362,N_12890);
xor U13935 (N_13935,N_12739,N_12626);
xor U13936 (N_13936,N_12476,N_12530);
nand U13937 (N_13937,N_12466,N_12629);
or U13938 (N_13938,N_12482,N_12831);
and U13939 (N_13939,N_12217,N_12142);
or U13940 (N_13940,N_12865,N_12253);
and U13941 (N_13941,N_12407,N_12478);
or U13942 (N_13942,N_12624,N_12507);
xor U13943 (N_13943,N_12329,N_12432);
or U13944 (N_13944,N_12176,N_12948);
xor U13945 (N_13945,N_12048,N_12323);
or U13946 (N_13946,N_12028,N_12832);
xnor U13947 (N_13947,N_12506,N_12239);
nand U13948 (N_13948,N_12034,N_12270);
nand U13949 (N_13949,N_12751,N_12450);
nor U13950 (N_13950,N_12364,N_12279);
xor U13951 (N_13951,N_12735,N_12441);
xor U13952 (N_13952,N_12689,N_12133);
and U13953 (N_13953,N_12885,N_12137);
nand U13954 (N_13954,N_12508,N_12817);
or U13955 (N_13955,N_12698,N_12966);
nor U13956 (N_13956,N_12196,N_12066);
xor U13957 (N_13957,N_12100,N_12270);
xnor U13958 (N_13958,N_12952,N_12976);
nor U13959 (N_13959,N_12622,N_12996);
or U13960 (N_13960,N_12790,N_12035);
and U13961 (N_13961,N_12709,N_12501);
or U13962 (N_13962,N_12524,N_12952);
or U13963 (N_13963,N_12997,N_12080);
xnor U13964 (N_13964,N_12363,N_12939);
and U13965 (N_13965,N_12909,N_12292);
or U13966 (N_13966,N_12318,N_12940);
or U13967 (N_13967,N_12216,N_12132);
nand U13968 (N_13968,N_12585,N_12280);
nand U13969 (N_13969,N_12326,N_12002);
nor U13970 (N_13970,N_12136,N_12542);
nand U13971 (N_13971,N_12459,N_12241);
or U13972 (N_13972,N_12491,N_12917);
and U13973 (N_13973,N_12989,N_12758);
or U13974 (N_13974,N_12219,N_12047);
and U13975 (N_13975,N_12984,N_12286);
nand U13976 (N_13976,N_12129,N_12984);
or U13977 (N_13977,N_12309,N_12876);
and U13978 (N_13978,N_12083,N_12005);
nor U13979 (N_13979,N_12624,N_12610);
nor U13980 (N_13980,N_12874,N_12026);
and U13981 (N_13981,N_12547,N_12467);
nand U13982 (N_13982,N_12289,N_12272);
xnor U13983 (N_13983,N_12851,N_12135);
or U13984 (N_13984,N_12803,N_12631);
xnor U13985 (N_13985,N_12740,N_12060);
and U13986 (N_13986,N_12128,N_12449);
and U13987 (N_13987,N_12166,N_12564);
or U13988 (N_13988,N_12539,N_12307);
xor U13989 (N_13989,N_12934,N_12528);
or U13990 (N_13990,N_12776,N_12522);
xor U13991 (N_13991,N_12609,N_12321);
or U13992 (N_13992,N_12176,N_12001);
or U13993 (N_13993,N_12621,N_12525);
or U13994 (N_13994,N_12320,N_12419);
nor U13995 (N_13995,N_12233,N_12674);
nor U13996 (N_13996,N_12169,N_12092);
xor U13997 (N_13997,N_12812,N_12526);
nand U13998 (N_13998,N_12605,N_12903);
and U13999 (N_13999,N_12163,N_12963);
or U14000 (N_14000,N_13441,N_13571);
nand U14001 (N_14001,N_13399,N_13889);
xnor U14002 (N_14002,N_13683,N_13372);
and U14003 (N_14003,N_13418,N_13915);
and U14004 (N_14004,N_13885,N_13522);
xnor U14005 (N_14005,N_13264,N_13628);
xnor U14006 (N_14006,N_13447,N_13704);
xor U14007 (N_14007,N_13845,N_13805);
and U14008 (N_14008,N_13289,N_13942);
xnor U14009 (N_14009,N_13682,N_13717);
nor U14010 (N_14010,N_13030,N_13993);
nor U14011 (N_14011,N_13755,N_13856);
xor U14012 (N_14012,N_13220,N_13147);
xnor U14013 (N_14013,N_13413,N_13462);
and U14014 (N_14014,N_13892,N_13047);
nor U14015 (N_14015,N_13467,N_13839);
or U14016 (N_14016,N_13108,N_13017);
and U14017 (N_14017,N_13419,N_13451);
xnor U14018 (N_14018,N_13888,N_13050);
and U14019 (N_14019,N_13563,N_13238);
and U14020 (N_14020,N_13354,N_13662);
or U14021 (N_14021,N_13958,N_13392);
xor U14022 (N_14022,N_13574,N_13280);
or U14023 (N_14023,N_13626,N_13529);
nand U14024 (N_14024,N_13216,N_13226);
nor U14025 (N_14025,N_13935,N_13016);
xnor U14026 (N_14026,N_13429,N_13635);
xor U14027 (N_14027,N_13715,N_13336);
and U14028 (N_14028,N_13273,N_13292);
xnor U14029 (N_14029,N_13351,N_13981);
and U14030 (N_14030,N_13896,N_13149);
and U14031 (N_14031,N_13294,N_13933);
and U14032 (N_14032,N_13903,N_13437);
nor U14033 (N_14033,N_13514,N_13559);
xor U14034 (N_14034,N_13056,N_13601);
nand U14035 (N_14035,N_13787,N_13008);
nor U14036 (N_14036,N_13802,N_13980);
nor U14037 (N_14037,N_13155,N_13389);
xnor U14038 (N_14038,N_13127,N_13257);
xor U14039 (N_14039,N_13078,N_13159);
nand U14040 (N_14040,N_13509,N_13209);
or U14041 (N_14041,N_13863,N_13846);
nor U14042 (N_14042,N_13893,N_13024);
nand U14043 (N_14043,N_13594,N_13849);
or U14044 (N_14044,N_13205,N_13577);
nor U14045 (N_14045,N_13157,N_13886);
and U14046 (N_14046,N_13227,N_13585);
nand U14047 (N_14047,N_13565,N_13525);
nor U14048 (N_14048,N_13552,N_13458);
nor U14049 (N_14049,N_13681,N_13171);
nand U14050 (N_14050,N_13262,N_13048);
xor U14051 (N_14051,N_13440,N_13907);
and U14052 (N_14052,N_13511,N_13781);
xnor U14053 (N_14053,N_13150,N_13766);
nand U14054 (N_14054,N_13368,N_13790);
and U14055 (N_14055,N_13290,N_13617);
and U14056 (N_14056,N_13712,N_13535);
and U14057 (N_14057,N_13070,N_13986);
and U14058 (N_14058,N_13870,N_13096);
and U14059 (N_14059,N_13597,N_13541);
or U14060 (N_14060,N_13723,N_13497);
nor U14061 (N_14061,N_13539,N_13039);
and U14062 (N_14062,N_13409,N_13533);
nor U14063 (N_14063,N_13148,N_13374);
and U14064 (N_14064,N_13680,N_13639);
or U14065 (N_14065,N_13385,N_13302);
nor U14066 (N_14066,N_13198,N_13143);
or U14067 (N_14067,N_13170,N_13854);
xor U14068 (N_14068,N_13791,N_13794);
and U14069 (N_14069,N_13929,N_13875);
or U14070 (N_14070,N_13486,N_13627);
and U14071 (N_14071,N_13334,N_13081);
xnor U14072 (N_14072,N_13003,N_13813);
nand U14073 (N_14073,N_13065,N_13855);
xor U14074 (N_14074,N_13260,N_13901);
and U14075 (N_14075,N_13167,N_13999);
and U14076 (N_14076,N_13689,N_13518);
and U14077 (N_14077,N_13809,N_13828);
and U14078 (N_14078,N_13006,N_13954);
nor U14079 (N_14079,N_13645,N_13801);
nand U14080 (N_14080,N_13820,N_13025);
nand U14081 (N_14081,N_13621,N_13156);
or U14082 (N_14082,N_13353,N_13387);
xor U14083 (N_14083,N_13974,N_13350);
and U14084 (N_14084,N_13201,N_13277);
or U14085 (N_14085,N_13530,N_13701);
or U14086 (N_14086,N_13270,N_13027);
or U14087 (N_14087,N_13707,N_13811);
nand U14088 (N_14088,N_13076,N_13971);
nand U14089 (N_14089,N_13948,N_13221);
nand U14090 (N_14090,N_13588,N_13745);
nor U14091 (N_14091,N_13864,N_13412);
nor U14092 (N_14092,N_13589,N_13946);
xnor U14093 (N_14093,N_13659,N_13778);
nand U14094 (N_14094,N_13873,N_13567);
nor U14095 (N_14095,N_13632,N_13152);
xor U14096 (N_14096,N_13636,N_13910);
or U14097 (N_14097,N_13840,N_13424);
xnor U14098 (N_14098,N_13814,N_13806);
xnor U14099 (N_14099,N_13106,N_13861);
xor U14100 (N_14100,N_13261,N_13105);
or U14101 (N_14101,N_13450,N_13477);
or U14102 (N_14102,N_13568,N_13322);
nor U14103 (N_14103,N_13022,N_13416);
xor U14104 (N_14104,N_13191,N_13400);
and U14105 (N_14105,N_13987,N_13528);
or U14106 (N_14106,N_13242,N_13734);
or U14107 (N_14107,N_13034,N_13950);
and U14108 (N_14108,N_13582,N_13190);
and U14109 (N_14109,N_13454,N_13376);
and U14110 (N_14110,N_13203,N_13579);
and U14111 (N_14111,N_13083,N_13713);
xnor U14112 (N_14112,N_13132,N_13179);
or U14113 (N_14113,N_13668,N_13009);
nor U14114 (N_14114,N_13938,N_13222);
or U14115 (N_14115,N_13783,N_13857);
or U14116 (N_14116,N_13442,N_13307);
nand U14117 (N_14117,N_13874,N_13556);
nor U14118 (N_14118,N_13599,N_13544);
and U14119 (N_14119,N_13268,N_13188);
nand U14120 (N_14120,N_13275,N_13004);
or U14121 (N_14121,N_13972,N_13433);
nand U14122 (N_14122,N_13575,N_13869);
nand U14123 (N_14123,N_13561,N_13310);
and U14124 (N_14124,N_13797,N_13320);
xor U14125 (N_14125,N_13118,N_13134);
nand U14126 (N_14126,N_13973,N_13510);
nor U14127 (N_14127,N_13474,N_13905);
xor U14128 (N_14128,N_13943,N_13452);
or U14129 (N_14129,N_13557,N_13103);
or U14130 (N_14130,N_13285,N_13671);
nor U14131 (N_14131,N_13696,N_13169);
nand U14132 (N_14132,N_13629,N_13168);
xnor U14133 (N_14133,N_13194,N_13042);
and U14134 (N_14134,N_13084,N_13064);
nor U14135 (N_14135,N_13494,N_13041);
nand U14136 (N_14136,N_13153,N_13521);
and U14137 (N_14137,N_13546,N_13463);
nand U14138 (N_14138,N_13286,N_13737);
or U14139 (N_14139,N_13775,N_13061);
xnor U14140 (N_14140,N_13945,N_13199);
xnor U14141 (N_14141,N_13381,N_13982);
nand U14142 (N_14142,N_13291,N_13918);
and U14143 (N_14143,N_13578,N_13214);
nand U14144 (N_14144,N_13736,N_13821);
xnor U14145 (N_14145,N_13773,N_13506);
nand U14146 (N_14146,N_13101,N_13512);
or U14147 (N_14147,N_13730,N_13665);
or U14148 (N_14148,N_13975,N_13448);
or U14149 (N_14149,N_13742,N_13465);
and U14150 (N_14150,N_13097,N_13142);
nand U14151 (N_14151,N_13023,N_13965);
or U14152 (N_14152,N_13332,N_13555);
xnor U14153 (N_14153,N_13240,N_13998);
or U14154 (N_14154,N_13379,N_13165);
nand U14155 (N_14155,N_13688,N_13378);
nor U14156 (N_14156,N_13739,N_13388);
and U14157 (N_14157,N_13230,N_13002);
or U14158 (N_14158,N_13218,N_13053);
xnor U14159 (N_14159,N_13941,N_13908);
nor U14160 (N_14160,N_13031,N_13407);
nand U14161 (N_14161,N_13693,N_13259);
nor U14162 (N_14162,N_13189,N_13576);
xnor U14163 (N_14163,N_13995,N_13115);
nor U14164 (N_14164,N_13923,N_13658);
nand U14165 (N_14165,N_13455,N_13445);
xnor U14166 (N_14166,N_13095,N_13532);
or U14167 (N_14167,N_13326,N_13902);
nand U14168 (N_14168,N_13883,N_13345);
nand U14169 (N_14169,N_13210,N_13196);
and U14170 (N_14170,N_13069,N_13234);
nor U14171 (N_14171,N_13666,N_13059);
or U14172 (N_14172,N_13733,N_13035);
or U14173 (N_14173,N_13288,N_13066);
xnor U14174 (N_14174,N_13318,N_13862);
or U14175 (N_14175,N_13010,N_13241);
and U14176 (N_14176,N_13921,N_13427);
xor U14177 (N_14177,N_13197,N_13560);
or U14178 (N_14178,N_13865,N_13001);
nand U14179 (N_14179,N_13648,N_13371);
nor U14180 (N_14180,N_13033,N_13835);
and U14181 (N_14181,N_13876,N_13204);
xnor U14182 (N_14182,N_13804,N_13303);
xnor U14183 (N_14183,N_13939,N_13894);
nand U14184 (N_14184,N_13356,N_13123);
and U14185 (N_14185,N_13164,N_13866);
nor U14186 (N_14186,N_13706,N_13361);
and U14187 (N_14187,N_13542,N_13130);
or U14188 (N_14188,N_13485,N_13674);
xnor U14189 (N_14189,N_13848,N_13761);
and U14190 (N_14190,N_13301,N_13306);
and U14191 (N_14191,N_13788,N_13075);
xor U14192 (N_14192,N_13128,N_13604);
or U14193 (N_14193,N_13135,N_13898);
and U14194 (N_14194,N_13235,N_13367);
or U14195 (N_14195,N_13384,N_13679);
nand U14196 (N_14196,N_13192,N_13670);
nor U14197 (N_14197,N_13151,N_13847);
nor U14198 (N_14198,N_13049,N_13746);
or U14199 (N_14199,N_13484,N_13082);
or U14200 (N_14200,N_13364,N_13686);
xor U14201 (N_14201,N_13110,N_13114);
xnor U14202 (N_14202,N_13776,N_13882);
and U14203 (N_14203,N_13058,N_13583);
and U14204 (N_14204,N_13838,N_13046);
xnor U14205 (N_14205,N_13104,N_13178);
xnor U14206 (N_14206,N_13481,N_13175);
or U14207 (N_14207,N_13710,N_13055);
xor U14208 (N_14208,N_13258,N_13697);
nand U14209 (N_14209,N_13432,N_13774);
nor U14210 (N_14210,N_13355,N_13767);
and U14211 (N_14211,N_13314,N_13077);
nand U14212 (N_14212,N_13482,N_13436);
xor U14213 (N_14213,N_13834,N_13523);
nand U14214 (N_14214,N_13906,N_13616);
and U14215 (N_14215,N_13393,N_13415);
or U14216 (N_14216,N_13446,N_13607);
nor U14217 (N_14217,N_13623,N_13187);
nor U14218 (N_14218,N_13630,N_13186);
nor U14219 (N_14219,N_13824,N_13703);
or U14220 (N_14220,N_13284,N_13045);
xor U14221 (N_14221,N_13961,N_13471);
and U14222 (N_14222,N_13928,N_13342);
or U14223 (N_14223,N_13282,N_13011);
or U14224 (N_14224,N_13656,N_13468);
xor U14225 (N_14225,N_13655,N_13653);
nand U14226 (N_14226,N_13229,N_13687);
or U14227 (N_14227,N_13837,N_13983);
nor U14228 (N_14228,N_13743,N_13019);
nand U14229 (N_14229,N_13373,N_13453);
and U14230 (N_14230,N_13633,N_13920);
nand U14231 (N_14231,N_13182,N_13072);
nand U14232 (N_14232,N_13914,N_13496);
or U14233 (N_14233,N_13762,N_13036);
nand U14234 (N_14234,N_13478,N_13324);
nor U14235 (N_14235,N_13581,N_13278);
or U14236 (N_14236,N_13493,N_13732);
or U14237 (N_14237,N_13858,N_13836);
nand U14238 (N_14238,N_13642,N_13449);
nor U14239 (N_14239,N_13185,N_13719);
nand U14240 (N_14240,N_13224,N_13113);
xor U14241 (N_14241,N_13705,N_13490);
nor U14242 (N_14242,N_13989,N_13333);
nor U14243 (N_14243,N_13722,N_13428);
nor U14244 (N_14244,N_13460,N_13803);
nor U14245 (N_14245,N_13536,N_13138);
or U14246 (N_14246,N_13233,N_13540);
xor U14247 (N_14247,N_13338,N_13466);
xor U14248 (N_14248,N_13608,N_13872);
and U14249 (N_14249,N_13405,N_13505);
nand U14250 (N_14250,N_13348,N_13649);
nor U14251 (N_14251,N_13700,N_13699);
and U14252 (N_14252,N_13266,N_13363);
nor U14253 (N_14253,N_13420,N_13650);
nand U14254 (N_14254,N_13744,N_13718);
nor U14255 (N_14255,N_13508,N_13231);
xnor U14256 (N_14256,N_13228,N_13800);
xor U14257 (N_14257,N_13756,N_13963);
and U14258 (N_14258,N_13044,N_13144);
nor U14259 (N_14259,N_13771,N_13988);
xor U14260 (N_14260,N_13362,N_13764);
or U14261 (N_14261,N_13232,N_13779);
or U14262 (N_14262,N_13513,N_13817);
nor U14263 (N_14263,N_13283,N_13877);
and U14264 (N_14264,N_13469,N_13960);
nand U14265 (N_14265,N_13099,N_13161);
nor U14266 (N_14266,N_13622,N_13654);
or U14267 (N_14267,N_13319,N_13037);
xnor U14268 (N_14268,N_13660,N_13964);
nand U14269 (N_14269,N_13396,N_13976);
or U14270 (N_14270,N_13352,N_13038);
xnor U14271 (N_14271,N_13272,N_13695);
and U14272 (N_14272,N_13526,N_13758);
and U14273 (N_14273,N_13184,N_13634);
or U14274 (N_14274,N_13211,N_13422);
xor U14275 (N_14275,N_13909,N_13538);
and U14276 (N_14276,N_13212,N_13459);
and U14277 (N_14277,N_13977,N_13215);
nor U14278 (N_14278,N_13491,N_13884);
xor U14279 (N_14279,N_13815,N_13631);
or U14280 (N_14280,N_13014,N_13602);
nand U14281 (N_14281,N_13299,N_13305);
nor U14282 (N_14282,N_13431,N_13068);
nand U14283 (N_14283,N_13217,N_13444);
and U14284 (N_14284,N_13207,N_13638);
and U14285 (N_14285,N_13590,N_13109);
nor U14286 (N_14286,N_13676,N_13456);
xor U14287 (N_14287,N_13430,N_13018);
and U14288 (N_14288,N_13461,N_13370);
nor U14289 (N_14289,N_13154,N_13625);
or U14290 (N_14290,N_13652,N_13054);
xnor U14291 (N_14291,N_13600,N_13959);
or U14292 (N_14292,N_13021,N_13895);
and U14293 (N_14293,N_13740,N_13669);
nand U14294 (N_14294,N_13380,N_13279);
or U14295 (N_14295,N_13253,N_13052);
or U14296 (N_14296,N_13093,N_13074);
and U14297 (N_14297,N_13812,N_13741);
nand U14298 (N_14298,N_13472,N_13359);
or U14299 (N_14299,N_13537,N_13944);
nor U14300 (N_14300,N_13615,N_13966);
or U14301 (N_14301,N_13166,N_13871);
or U14302 (N_14302,N_13911,N_13947);
nor U14303 (N_14303,N_13738,N_13750);
nor U14304 (N_14304,N_13426,N_13819);
xnor U14305 (N_14305,N_13757,N_13916);
nand U14306 (N_14306,N_13488,N_13661);
and U14307 (N_14307,N_13562,N_13726);
nand U14308 (N_14308,N_13735,N_13133);
or U14309 (N_14309,N_13867,N_13271);
xnor U14310 (N_14310,N_13969,N_13040);
and U14311 (N_14311,N_13953,N_13564);
nor U14312 (N_14312,N_13470,N_13090);
nor U14313 (N_14313,N_13624,N_13618);
nor U14314 (N_14314,N_13489,N_13598);
xnor U14315 (N_14315,N_13256,N_13434);
xor U14316 (N_14316,N_13487,N_13709);
or U14317 (N_14317,N_13495,N_13769);
nor U14318 (N_14318,N_13934,N_13749);
nand U14319 (N_14319,N_13408,N_13287);
nor U14320 (N_14320,N_13213,N_13527);
or U14321 (N_14321,N_13254,N_13690);
or U14322 (N_14322,N_13312,N_13347);
nor U14323 (N_14323,N_13116,N_13646);
nor U14324 (N_14324,N_13702,N_13644);
nand U14325 (N_14325,N_13851,N_13094);
nor U14326 (N_14326,N_13970,N_13425);
and U14327 (N_14327,N_13507,N_13637);
or U14328 (N_14328,N_13247,N_13913);
or U14329 (N_14329,N_13401,N_13088);
or U14330 (N_14330,N_13293,N_13558);
xnor U14331 (N_14331,N_13841,N_13267);
nand U14332 (N_14332,N_13772,N_13193);
xnor U14333 (N_14333,N_13464,N_13949);
and U14334 (N_14334,N_13691,N_13789);
xor U14335 (N_14335,N_13091,N_13092);
and U14336 (N_14336,N_13675,N_13295);
nor U14337 (N_14337,N_13765,N_13780);
or U14338 (N_14338,N_13316,N_13032);
and U14339 (N_14339,N_13798,N_13968);
nor U14340 (N_14340,N_13202,N_13760);
or U14341 (N_14341,N_13503,N_13410);
or U14342 (N_14342,N_13952,N_13071);
xor U14343 (N_14343,N_13519,N_13844);
or U14344 (N_14344,N_13079,N_13026);
xor U14345 (N_14345,N_13647,N_13515);
or U14346 (N_14346,N_13793,N_13304);
nor U14347 (N_14347,N_13028,N_13296);
nand U14348 (N_14348,N_13818,N_13940);
nand U14349 (N_14349,N_13122,N_13610);
and U14350 (N_14350,N_13724,N_13891);
and U14351 (N_14351,N_13163,N_13951);
nand U14352 (N_14352,N_13102,N_13657);
nand U14353 (N_14353,N_13534,N_13225);
nand U14354 (N_14354,N_13043,N_13850);
nor U14355 (N_14355,N_13501,N_13878);
nor U14356 (N_14356,N_13421,N_13395);
and U14357 (N_14357,N_13341,N_13897);
and U14358 (N_14358,N_13176,N_13181);
nor U14359 (N_14359,N_13605,N_13587);
nand U14360 (N_14360,N_13816,N_13978);
xor U14361 (N_14361,N_13580,N_13208);
nand U14362 (N_14362,N_13782,N_13754);
and U14363 (N_14363,N_13435,N_13842);
nor U14364 (N_14364,N_13339,N_13728);
or U14365 (N_14365,N_13140,N_13369);
or U14366 (N_14366,N_13711,N_13829);
xor U14367 (N_14367,N_13331,N_13553);
or U14368 (N_14368,N_13007,N_13125);
or U14369 (N_14369,N_13573,N_13263);
nand U14370 (N_14370,N_13985,N_13708);
or U14371 (N_14371,N_13141,N_13309);
xnor U14372 (N_14372,N_13930,N_13725);
nand U14373 (N_14373,N_13015,N_13139);
nand U14374 (N_14374,N_13759,N_13593);
xnor U14375 (N_14375,N_13276,N_13927);
xor U14376 (N_14376,N_13000,N_13752);
nand U14377 (N_14377,N_13062,N_13868);
and U14378 (N_14378,N_13281,N_13584);
or U14379 (N_14379,N_13543,N_13398);
xnor U14380 (N_14380,N_13063,N_13606);
nor U14381 (N_14381,N_13195,N_13795);
and U14382 (N_14382,N_13881,N_13912);
xnor U14383 (N_14383,N_13620,N_13830);
nand U14384 (N_14384,N_13479,N_13344);
and U14385 (N_14385,N_13126,N_13298);
nor U14386 (N_14386,N_13173,N_13520);
nor U14387 (N_14387,N_13329,N_13569);
nand U14388 (N_14388,N_13531,N_13770);
and U14389 (N_14389,N_13498,N_13545);
nor U14390 (N_14390,N_13366,N_13890);
or U14391 (N_14391,N_13483,N_13162);
xor U14392 (N_14392,N_13475,N_13112);
and U14393 (N_14393,N_13786,N_13614);
and U14394 (N_14394,N_13252,N_13547);
xnor U14395 (N_14395,N_13146,N_13925);
nor U14396 (N_14396,N_13524,N_13439);
xor U14397 (N_14397,N_13360,N_13183);
or U14398 (N_14398,N_13349,N_13924);
or U14399 (N_14399,N_13394,N_13994);
nand U14400 (N_14400,N_13404,N_13651);
nor U14401 (N_14401,N_13346,N_13124);
nand U14402 (N_14402,N_13997,N_13119);
and U14403 (N_14403,N_13922,N_13566);
xnor U14404 (N_14404,N_13714,N_13586);
and U14405 (N_14405,N_13411,N_13784);
nand U14406 (N_14406,N_13777,N_13956);
nor U14407 (N_14407,N_13554,N_13200);
nand U14408 (N_14408,N_13219,N_13992);
xnor U14409 (N_14409,N_13751,N_13438);
nand U14410 (N_14410,N_13067,N_13297);
nor U14411 (N_14411,N_13249,N_13832);
nand U14412 (N_14412,N_13810,N_13315);
xnor U14413 (N_14413,N_13936,N_13685);
xnor U14414 (N_14414,N_13255,N_13492);
and U14415 (N_14415,N_13603,N_13129);
xor U14416 (N_14416,N_13158,N_13323);
xnor U14417 (N_14417,N_13317,N_13570);
nor U14418 (N_14418,N_13926,N_13340);
or U14419 (N_14419,N_13859,N_13414);
nor U14420 (N_14420,N_13619,N_13808);
and U14421 (N_14421,N_13382,N_13990);
xnor U14422 (N_14422,N_13747,N_13962);
nand U14423 (N_14423,N_13500,N_13612);
and U14424 (N_14424,N_13677,N_13269);
or U14425 (N_14425,N_13698,N_13753);
or U14426 (N_14426,N_13517,N_13796);
and U14427 (N_14427,N_13731,N_13476);
or U14428 (N_14428,N_13337,N_13641);
or U14429 (N_14429,N_13057,N_13423);
nand U14430 (N_14430,N_13991,N_13357);
nor U14431 (N_14431,N_13223,N_13406);
nand U14432 (N_14432,N_13822,N_13852);
and U14433 (N_14433,N_13785,N_13716);
and U14434 (N_14434,N_13720,N_13879);
xnor U14435 (N_14435,N_13365,N_13321);
or U14436 (N_14436,N_13694,N_13473);
xnor U14437 (N_14437,N_13311,N_13826);
nor U14438 (N_14438,N_13937,N_13174);
nor U14439 (N_14439,N_13145,N_13051);
or U14440 (N_14440,N_13206,N_13480);
and U14441 (N_14441,N_13085,N_13328);
nand U14442 (N_14442,N_13799,N_13265);
or U14443 (N_14443,N_13919,N_13087);
or U14444 (N_14444,N_13107,N_13086);
xnor U14445 (N_14445,N_13012,N_13548);
and U14446 (N_14446,N_13343,N_13136);
and U14447 (N_14447,N_13377,N_13640);
nor U14448 (N_14448,N_13692,N_13609);
nand U14449 (N_14449,N_13443,N_13239);
nand U14450 (N_14450,N_13899,N_13613);
and U14451 (N_14451,N_13792,N_13073);
and U14452 (N_14452,N_13243,N_13248);
or U14453 (N_14453,N_13313,N_13768);
nor U14454 (N_14454,N_13502,N_13663);
nor U14455 (N_14455,N_13403,N_13131);
xnor U14456 (N_14456,N_13833,N_13020);
and U14457 (N_14457,N_13823,N_13236);
or U14458 (N_14458,N_13013,N_13967);
xor U14459 (N_14459,N_13550,N_13391);
or U14460 (N_14460,N_13572,N_13664);
nand U14461 (N_14461,N_13121,N_13727);
and U14462 (N_14462,N_13996,N_13120);
or U14463 (N_14463,N_13827,N_13729);
nand U14464 (N_14464,N_13386,N_13375);
nand U14465 (N_14465,N_13029,N_13327);
and U14466 (N_14466,N_13807,N_13900);
xor U14467 (N_14467,N_13250,N_13005);
or U14468 (N_14468,N_13672,N_13499);
or U14469 (N_14469,N_13244,N_13117);
and U14470 (N_14470,N_13504,N_13955);
nand U14471 (N_14471,N_13611,N_13308);
xnor U14472 (N_14472,N_13957,N_13595);
nand U14473 (N_14473,N_13932,N_13358);
xor U14474 (N_14474,N_13325,N_13853);
nor U14475 (N_14475,N_13831,N_13643);
and U14476 (N_14476,N_13060,N_13904);
xnor U14477 (N_14477,N_13330,N_13237);
nor U14478 (N_14478,N_13089,N_13667);
or U14479 (N_14479,N_13111,N_13843);
and U14480 (N_14480,N_13591,N_13390);
nor U14481 (N_14481,N_13300,N_13100);
or U14482 (N_14482,N_13457,N_13397);
and U14483 (N_14483,N_13917,N_13274);
and U14484 (N_14484,N_13673,N_13684);
nand U14485 (N_14485,N_13979,N_13748);
and U14486 (N_14486,N_13383,N_13763);
or U14487 (N_14487,N_13180,N_13172);
or U14488 (N_14488,N_13402,N_13551);
and U14489 (N_14489,N_13335,N_13137);
or U14490 (N_14490,N_13177,N_13984);
and U14491 (N_14491,N_13098,N_13245);
and U14492 (N_14492,N_13080,N_13678);
and U14493 (N_14493,N_13860,N_13880);
or U14494 (N_14494,N_13516,N_13417);
and U14495 (N_14495,N_13825,N_13592);
or U14496 (N_14496,N_13246,N_13549);
nand U14497 (N_14497,N_13596,N_13931);
nand U14498 (N_14498,N_13887,N_13160);
nand U14499 (N_14499,N_13721,N_13251);
nand U14500 (N_14500,N_13390,N_13223);
or U14501 (N_14501,N_13846,N_13829);
nand U14502 (N_14502,N_13520,N_13800);
nand U14503 (N_14503,N_13752,N_13619);
or U14504 (N_14504,N_13903,N_13236);
or U14505 (N_14505,N_13536,N_13854);
and U14506 (N_14506,N_13753,N_13583);
nor U14507 (N_14507,N_13128,N_13818);
xnor U14508 (N_14508,N_13200,N_13540);
or U14509 (N_14509,N_13229,N_13752);
nand U14510 (N_14510,N_13868,N_13011);
nor U14511 (N_14511,N_13919,N_13207);
and U14512 (N_14512,N_13741,N_13562);
xnor U14513 (N_14513,N_13244,N_13261);
xor U14514 (N_14514,N_13149,N_13330);
and U14515 (N_14515,N_13569,N_13443);
or U14516 (N_14516,N_13427,N_13766);
and U14517 (N_14517,N_13845,N_13681);
and U14518 (N_14518,N_13370,N_13792);
nand U14519 (N_14519,N_13523,N_13222);
xnor U14520 (N_14520,N_13881,N_13128);
nand U14521 (N_14521,N_13325,N_13905);
or U14522 (N_14522,N_13672,N_13486);
xnor U14523 (N_14523,N_13133,N_13746);
nor U14524 (N_14524,N_13407,N_13546);
nor U14525 (N_14525,N_13487,N_13454);
nand U14526 (N_14526,N_13420,N_13599);
nor U14527 (N_14527,N_13396,N_13157);
nor U14528 (N_14528,N_13344,N_13111);
nand U14529 (N_14529,N_13056,N_13160);
xor U14530 (N_14530,N_13804,N_13135);
nand U14531 (N_14531,N_13324,N_13462);
nand U14532 (N_14532,N_13049,N_13917);
and U14533 (N_14533,N_13731,N_13370);
and U14534 (N_14534,N_13552,N_13625);
or U14535 (N_14535,N_13810,N_13747);
or U14536 (N_14536,N_13265,N_13076);
nor U14537 (N_14537,N_13348,N_13367);
and U14538 (N_14538,N_13527,N_13014);
or U14539 (N_14539,N_13791,N_13634);
and U14540 (N_14540,N_13396,N_13433);
nand U14541 (N_14541,N_13597,N_13302);
nand U14542 (N_14542,N_13426,N_13614);
xor U14543 (N_14543,N_13328,N_13174);
and U14544 (N_14544,N_13070,N_13956);
nand U14545 (N_14545,N_13433,N_13379);
and U14546 (N_14546,N_13980,N_13184);
and U14547 (N_14547,N_13274,N_13028);
nor U14548 (N_14548,N_13669,N_13939);
and U14549 (N_14549,N_13218,N_13104);
or U14550 (N_14550,N_13578,N_13312);
or U14551 (N_14551,N_13562,N_13054);
or U14552 (N_14552,N_13346,N_13507);
and U14553 (N_14553,N_13028,N_13525);
xnor U14554 (N_14554,N_13439,N_13574);
and U14555 (N_14555,N_13088,N_13334);
xnor U14556 (N_14556,N_13817,N_13941);
xnor U14557 (N_14557,N_13173,N_13020);
xor U14558 (N_14558,N_13020,N_13895);
xnor U14559 (N_14559,N_13013,N_13362);
and U14560 (N_14560,N_13853,N_13792);
nor U14561 (N_14561,N_13018,N_13413);
or U14562 (N_14562,N_13360,N_13284);
or U14563 (N_14563,N_13816,N_13025);
nor U14564 (N_14564,N_13928,N_13329);
xnor U14565 (N_14565,N_13491,N_13215);
xnor U14566 (N_14566,N_13876,N_13235);
nand U14567 (N_14567,N_13424,N_13405);
nand U14568 (N_14568,N_13036,N_13345);
nor U14569 (N_14569,N_13983,N_13713);
and U14570 (N_14570,N_13674,N_13426);
nand U14571 (N_14571,N_13852,N_13747);
or U14572 (N_14572,N_13808,N_13657);
or U14573 (N_14573,N_13283,N_13017);
xnor U14574 (N_14574,N_13968,N_13944);
and U14575 (N_14575,N_13859,N_13710);
or U14576 (N_14576,N_13818,N_13056);
nor U14577 (N_14577,N_13040,N_13031);
and U14578 (N_14578,N_13067,N_13375);
nand U14579 (N_14579,N_13563,N_13068);
nand U14580 (N_14580,N_13331,N_13386);
nand U14581 (N_14581,N_13551,N_13016);
or U14582 (N_14582,N_13188,N_13611);
xor U14583 (N_14583,N_13522,N_13651);
nand U14584 (N_14584,N_13608,N_13554);
and U14585 (N_14585,N_13174,N_13825);
xnor U14586 (N_14586,N_13252,N_13756);
or U14587 (N_14587,N_13191,N_13591);
and U14588 (N_14588,N_13324,N_13042);
or U14589 (N_14589,N_13974,N_13878);
nand U14590 (N_14590,N_13263,N_13129);
or U14591 (N_14591,N_13604,N_13420);
nor U14592 (N_14592,N_13779,N_13451);
or U14593 (N_14593,N_13138,N_13788);
nand U14594 (N_14594,N_13949,N_13328);
xnor U14595 (N_14595,N_13656,N_13027);
nor U14596 (N_14596,N_13244,N_13815);
nor U14597 (N_14597,N_13390,N_13933);
or U14598 (N_14598,N_13288,N_13485);
or U14599 (N_14599,N_13123,N_13922);
and U14600 (N_14600,N_13527,N_13852);
xor U14601 (N_14601,N_13260,N_13365);
and U14602 (N_14602,N_13168,N_13336);
xor U14603 (N_14603,N_13237,N_13115);
and U14604 (N_14604,N_13823,N_13594);
nor U14605 (N_14605,N_13739,N_13343);
nor U14606 (N_14606,N_13593,N_13584);
and U14607 (N_14607,N_13433,N_13512);
and U14608 (N_14608,N_13337,N_13970);
and U14609 (N_14609,N_13494,N_13442);
or U14610 (N_14610,N_13058,N_13745);
or U14611 (N_14611,N_13177,N_13837);
xnor U14612 (N_14612,N_13464,N_13033);
nor U14613 (N_14613,N_13374,N_13758);
and U14614 (N_14614,N_13213,N_13745);
nand U14615 (N_14615,N_13709,N_13842);
nand U14616 (N_14616,N_13458,N_13155);
nor U14617 (N_14617,N_13074,N_13738);
xnor U14618 (N_14618,N_13133,N_13074);
or U14619 (N_14619,N_13856,N_13519);
nand U14620 (N_14620,N_13244,N_13510);
nand U14621 (N_14621,N_13110,N_13651);
nand U14622 (N_14622,N_13337,N_13386);
and U14623 (N_14623,N_13663,N_13568);
or U14624 (N_14624,N_13340,N_13697);
nand U14625 (N_14625,N_13180,N_13107);
or U14626 (N_14626,N_13677,N_13515);
or U14627 (N_14627,N_13641,N_13560);
and U14628 (N_14628,N_13081,N_13054);
and U14629 (N_14629,N_13907,N_13590);
xor U14630 (N_14630,N_13551,N_13294);
nor U14631 (N_14631,N_13927,N_13947);
xor U14632 (N_14632,N_13588,N_13473);
xnor U14633 (N_14633,N_13584,N_13112);
nand U14634 (N_14634,N_13901,N_13693);
or U14635 (N_14635,N_13903,N_13252);
and U14636 (N_14636,N_13631,N_13808);
and U14637 (N_14637,N_13651,N_13465);
and U14638 (N_14638,N_13455,N_13465);
xnor U14639 (N_14639,N_13669,N_13018);
nand U14640 (N_14640,N_13818,N_13148);
xor U14641 (N_14641,N_13834,N_13727);
and U14642 (N_14642,N_13212,N_13516);
xnor U14643 (N_14643,N_13704,N_13300);
and U14644 (N_14644,N_13218,N_13630);
xor U14645 (N_14645,N_13965,N_13696);
xor U14646 (N_14646,N_13486,N_13859);
or U14647 (N_14647,N_13348,N_13280);
nand U14648 (N_14648,N_13922,N_13990);
nor U14649 (N_14649,N_13439,N_13949);
or U14650 (N_14650,N_13934,N_13640);
xnor U14651 (N_14651,N_13378,N_13491);
and U14652 (N_14652,N_13908,N_13656);
or U14653 (N_14653,N_13026,N_13085);
nand U14654 (N_14654,N_13089,N_13387);
and U14655 (N_14655,N_13514,N_13842);
or U14656 (N_14656,N_13171,N_13760);
and U14657 (N_14657,N_13698,N_13091);
or U14658 (N_14658,N_13029,N_13779);
xnor U14659 (N_14659,N_13581,N_13863);
xor U14660 (N_14660,N_13468,N_13398);
nor U14661 (N_14661,N_13966,N_13752);
and U14662 (N_14662,N_13400,N_13915);
nor U14663 (N_14663,N_13207,N_13282);
and U14664 (N_14664,N_13624,N_13535);
xnor U14665 (N_14665,N_13160,N_13335);
nand U14666 (N_14666,N_13899,N_13047);
and U14667 (N_14667,N_13951,N_13605);
nand U14668 (N_14668,N_13756,N_13106);
and U14669 (N_14669,N_13129,N_13775);
and U14670 (N_14670,N_13232,N_13623);
nand U14671 (N_14671,N_13105,N_13687);
xor U14672 (N_14672,N_13866,N_13629);
or U14673 (N_14673,N_13958,N_13587);
and U14674 (N_14674,N_13066,N_13263);
nand U14675 (N_14675,N_13317,N_13125);
nor U14676 (N_14676,N_13072,N_13783);
nand U14677 (N_14677,N_13054,N_13060);
and U14678 (N_14678,N_13375,N_13546);
xor U14679 (N_14679,N_13651,N_13001);
and U14680 (N_14680,N_13535,N_13370);
nor U14681 (N_14681,N_13718,N_13201);
and U14682 (N_14682,N_13247,N_13551);
or U14683 (N_14683,N_13596,N_13136);
and U14684 (N_14684,N_13236,N_13524);
xor U14685 (N_14685,N_13086,N_13080);
nand U14686 (N_14686,N_13591,N_13086);
nor U14687 (N_14687,N_13354,N_13649);
nand U14688 (N_14688,N_13273,N_13867);
nand U14689 (N_14689,N_13524,N_13183);
nor U14690 (N_14690,N_13417,N_13894);
or U14691 (N_14691,N_13452,N_13174);
nand U14692 (N_14692,N_13391,N_13030);
or U14693 (N_14693,N_13938,N_13865);
nand U14694 (N_14694,N_13858,N_13047);
xor U14695 (N_14695,N_13886,N_13988);
nand U14696 (N_14696,N_13088,N_13521);
nor U14697 (N_14697,N_13070,N_13023);
or U14698 (N_14698,N_13569,N_13205);
or U14699 (N_14699,N_13328,N_13780);
and U14700 (N_14700,N_13991,N_13034);
nand U14701 (N_14701,N_13707,N_13227);
nor U14702 (N_14702,N_13083,N_13489);
or U14703 (N_14703,N_13690,N_13386);
and U14704 (N_14704,N_13701,N_13669);
nor U14705 (N_14705,N_13820,N_13117);
and U14706 (N_14706,N_13049,N_13579);
or U14707 (N_14707,N_13627,N_13483);
or U14708 (N_14708,N_13282,N_13368);
nor U14709 (N_14709,N_13047,N_13330);
nor U14710 (N_14710,N_13825,N_13154);
xor U14711 (N_14711,N_13797,N_13381);
and U14712 (N_14712,N_13455,N_13724);
and U14713 (N_14713,N_13032,N_13064);
and U14714 (N_14714,N_13501,N_13398);
xnor U14715 (N_14715,N_13563,N_13780);
nand U14716 (N_14716,N_13637,N_13124);
and U14717 (N_14717,N_13517,N_13418);
and U14718 (N_14718,N_13934,N_13025);
xor U14719 (N_14719,N_13588,N_13822);
and U14720 (N_14720,N_13553,N_13243);
nand U14721 (N_14721,N_13925,N_13102);
nand U14722 (N_14722,N_13237,N_13532);
and U14723 (N_14723,N_13590,N_13630);
nor U14724 (N_14724,N_13131,N_13039);
or U14725 (N_14725,N_13855,N_13002);
and U14726 (N_14726,N_13469,N_13178);
xnor U14727 (N_14727,N_13724,N_13964);
and U14728 (N_14728,N_13990,N_13628);
xor U14729 (N_14729,N_13239,N_13872);
nand U14730 (N_14730,N_13897,N_13128);
and U14731 (N_14731,N_13979,N_13697);
and U14732 (N_14732,N_13011,N_13664);
nand U14733 (N_14733,N_13493,N_13702);
nand U14734 (N_14734,N_13865,N_13602);
xnor U14735 (N_14735,N_13982,N_13731);
or U14736 (N_14736,N_13814,N_13600);
nor U14737 (N_14737,N_13772,N_13493);
and U14738 (N_14738,N_13527,N_13118);
nand U14739 (N_14739,N_13358,N_13536);
or U14740 (N_14740,N_13163,N_13958);
or U14741 (N_14741,N_13037,N_13468);
xnor U14742 (N_14742,N_13153,N_13968);
and U14743 (N_14743,N_13162,N_13707);
or U14744 (N_14744,N_13933,N_13635);
and U14745 (N_14745,N_13794,N_13171);
and U14746 (N_14746,N_13598,N_13780);
and U14747 (N_14747,N_13604,N_13213);
nand U14748 (N_14748,N_13193,N_13528);
nor U14749 (N_14749,N_13273,N_13993);
nand U14750 (N_14750,N_13445,N_13199);
or U14751 (N_14751,N_13866,N_13566);
nand U14752 (N_14752,N_13611,N_13589);
nand U14753 (N_14753,N_13787,N_13465);
nor U14754 (N_14754,N_13095,N_13546);
and U14755 (N_14755,N_13890,N_13751);
or U14756 (N_14756,N_13249,N_13561);
xnor U14757 (N_14757,N_13107,N_13914);
or U14758 (N_14758,N_13451,N_13618);
xor U14759 (N_14759,N_13097,N_13861);
or U14760 (N_14760,N_13106,N_13971);
nand U14761 (N_14761,N_13669,N_13073);
xnor U14762 (N_14762,N_13422,N_13470);
and U14763 (N_14763,N_13527,N_13799);
and U14764 (N_14764,N_13130,N_13766);
nor U14765 (N_14765,N_13913,N_13182);
nand U14766 (N_14766,N_13075,N_13147);
or U14767 (N_14767,N_13738,N_13355);
and U14768 (N_14768,N_13754,N_13743);
and U14769 (N_14769,N_13572,N_13054);
nor U14770 (N_14770,N_13289,N_13741);
or U14771 (N_14771,N_13096,N_13949);
nand U14772 (N_14772,N_13157,N_13306);
xnor U14773 (N_14773,N_13359,N_13300);
and U14774 (N_14774,N_13465,N_13901);
or U14775 (N_14775,N_13272,N_13154);
nor U14776 (N_14776,N_13667,N_13248);
and U14777 (N_14777,N_13553,N_13592);
or U14778 (N_14778,N_13020,N_13898);
or U14779 (N_14779,N_13008,N_13363);
nor U14780 (N_14780,N_13299,N_13035);
nor U14781 (N_14781,N_13454,N_13004);
nor U14782 (N_14782,N_13135,N_13409);
nand U14783 (N_14783,N_13661,N_13296);
and U14784 (N_14784,N_13267,N_13113);
nand U14785 (N_14785,N_13154,N_13467);
and U14786 (N_14786,N_13396,N_13439);
nor U14787 (N_14787,N_13838,N_13645);
xor U14788 (N_14788,N_13872,N_13801);
and U14789 (N_14789,N_13551,N_13884);
xor U14790 (N_14790,N_13609,N_13732);
nor U14791 (N_14791,N_13306,N_13055);
and U14792 (N_14792,N_13269,N_13854);
or U14793 (N_14793,N_13923,N_13579);
and U14794 (N_14794,N_13762,N_13813);
nor U14795 (N_14795,N_13287,N_13087);
or U14796 (N_14796,N_13776,N_13098);
nor U14797 (N_14797,N_13762,N_13081);
and U14798 (N_14798,N_13088,N_13666);
or U14799 (N_14799,N_13267,N_13578);
nand U14800 (N_14800,N_13604,N_13296);
xnor U14801 (N_14801,N_13051,N_13359);
xor U14802 (N_14802,N_13803,N_13671);
nand U14803 (N_14803,N_13806,N_13839);
and U14804 (N_14804,N_13120,N_13587);
xnor U14805 (N_14805,N_13250,N_13882);
nand U14806 (N_14806,N_13303,N_13494);
xnor U14807 (N_14807,N_13480,N_13083);
and U14808 (N_14808,N_13836,N_13125);
nor U14809 (N_14809,N_13061,N_13546);
or U14810 (N_14810,N_13682,N_13568);
nand U14811 (N_14811,N_13317,N_13397);
and U14812 (N_14812,N_13933,N_13638);
nor U14813 (N_14813,N_13441,N_13847);
nor U14814 (N_14814,N_13598,N_13218);
nor U14815 (N_14815,N_13353,N_13384);
xnor U14816 (N_14816,N_13389,N_13584);
or U14817 (N_14817,N_13965,N_13377);
or U14818 (N_14818,N_13299,N_13394);
and U14819 (N_14819,N_13720,N_13686);
nor U14820 (N_14820,N_13218,N_13874);
nand U14821 (N_14821,N_13293,N_13325);
and U14822 (N_14822,N_13312,N_13818);
nand U14823 (N_14823,N_13454,N_13247);
or U14824 (N_14824,N_13079,N_13378);
and U14825 (N_14825,N_13716,N_13805);
or U14826 (N_14826,N_13456,N_13121);
and U14827 (N_14827,N_13502,N_13651);
nand U14828 (N_14828,N_13335,N_13190);
nand U14829 (N_14829,N_13783,N_13347);
xor U14830 (N_14830,N_13532,N_13273);
xor U14831 (N_14831,N_13976,N_13736);
or U14832 (N_14832,N_13632,N_13638);
nand U14833 (N_14833,N_13909,N_13665);
or U14834 (N_14834,N_13486,N_13773);
or U14835 (N_14835,N_13576,N_13808);
and U14836 (N_14836,N_13830,N_13057);
nand U14837 (N_14837,N_13239,N_13983);
xnor U14838 (N_14838,N_13499,N_13345);
nor U14839 (N_14839,N_13716,N_13573);
and U14840 (N_14840,N_13231,N_13230);
nand U14841 (N_14841,N_13596,N_13521);
nor U14842 (N_14842,N_13802,N_13775);
or U14843 (N_14843,N_13365,N_13664);
xnor U14844 (N_14844,N_13943,N_13648);
or U14845 (N_14845,N_13397,N_13991);
and U14846 (N_14846,N_13019,N_13869);
and U14847 (N_14847,N_13711,N_13401);
and U14848 (N_14848,N_13598,N_13266);
and U14849 (N_14849,N_13773,N_13844);
and U14850 (N_14850,N_13671,N_13175);
or U14851 (N_14851,N_13726,N_13779);
and U14852 (N_14852,N_13007,N_13804);
xor U14853 (N_14853,N_13768,N_13125);
and U14854 (N_14854,N_13417,N_13256);
and U14855 (N_14855,N_13305,N_13812);
and U14856 (N_14856,N_13041,N_13395);
nand U14857 (N_14857,N_13525,N_13693);
and U14858 (N_14858,N_13890,N_13123);
xnor U14859 (N_14859,N_13236,N_13622);
and U14860 (N_14860,N_13947,N_13848);
and U14861 (N_14861,N_13322,N_13154);
and U14862 (N_14862,N_13405,N_13939);
nor U14863 (N_14863,N_13369,N_13185);
nor U14864 (N_14864,N_13590,N_13391);
nor U14865 (N_14865,N_13851,N_13129);
nor U14866 (N_14866,N_13132,N_13421);
or U14867 (N_14867,N_13080,N_13661);
nor U14868 (N_14868,N_13828,N_13870);
and U14869 (N_14869,N_13678,N_13082);
or U14870 (N_14870,N_13948,N_13656);
or U14871 (N_14871,N_13240,N_13268);
and U14872 (N_14872,N_13859,N_13676);
or U14873 (N_14873,N_13625,N_13196);
nand U14874 (N_14874,N_13488,N_13008);
and U14875 (N_14875,N_13843,N_13228);
nor U14876 (N_14876,N_13365,N_13790);
xor U14877 (N_14877,N_13065,N_13665);
nor U14878 (N_14878,N_13009,N_13464);
nor U14879 (N_14879,N_13356,N_13984);
xnor U14880 (N_14880,N_13397,N_13405);
or U14881 (N_14881,N_13665,N_13255);
nor U14882 (N_14882,N_13072,N_13689);
xor U14883 (N_14883,N_13575,N_13303);
xnor U14884 (N_14884,N_13217,N_13582);
and U14885 (N_14885,N_13823,N_13951);
nor U14886 (N_14886,N_13159,N_13141);
nor U14887 (N_14887,N_13431,N_13171);
and U14888 (N_14888,N_13713,N_13584);
or U14889 (N_14889,N_13061,N_13877);
xnor U14890 (N_14890,N_13984,N_13677);
or U14891 (N_14891,N_13063,N_13767);
and U14892 (N_14892,N_13473,N_13533);
or U14893 (N_14893,N_13917,N_13023);
or U14894 (N_14894,N_13562,N_13686);
nand U14895 (N_14895,N_13973,N_13775);
and U14896 (N_14896,N_13777,N_13639);
or U14897 (N_14897,N_13285,N_13930);
or U14898 (N_14898,N_13365,N_13597);
or U14899 (N_14899,N_13341,N_13733);
nand U14900 (N_14900,N_13287,N_13765);
nand U14901 (N_14901,N_13226,N_13325);
xor U14902 (N_14902,N_13009,N_13444);
nand U14903 (N_14903,N_13920,N_13672);
or U14904 (N_14904,N_13691,N_13011);
nand U14905 (N_14905,N_13804,N_13346);
nor U14906 (N_14906,N_13746,N_13640);
and U14907 (N_14907,N_13166,N_13738);
and U14908 (N_14908,N_13739,N_13344);
nand U14909 (N_14909,N_13951,N_13534);
or U14910 (N_14910,N_13281,N_13798);
or U14911 (N_14911,N_13441,N_13825);
or U14912 (N_14912,N_13730,N_13848);
xor U14913 (N_14913,N_13195,N_13357);
and U14914 (N_14914,N_13361,N_13015);
or U14915 (N_14915,N_13196,N_13588);
xnor U14916 (N_14916,N_13167,N_13077);
nor U14917 (N_14917,N_13131,N_13051);
or U14918 (N_14918,N_13283,N_13235);
nand U14919 (N_14919,N_13413,N_13919);
or U14920 (N_14920,N_13765,N_13323);
nor U14921 (N_14921,N_13887,N_13775);
nor U14922 (N_14922,N_13218,N_13683);
nand U14923 (N_14923,N_13262,N_13324);
and U14924 (N_14924,N_13603,N_13684);
or U14925 (N_14925,N_13756,N_13575);
xnor U14926 (N_14926,N_13172,N_13087);
nand U14927 (N_14927,N_13779,N_13807);
nor U14928 (N_14928,N_13596,N_13258);
and U14929 (N_14929,N_13387,N_13153);
and U14930 (N_14930,N_13614,N_13888);
nor U14931 (N_14931,N_13604,N_13471);
and U14932 (N_14932,N_13478,N_13116);
or U14933 (N_14933,N_13778,N_13231);
xor U14934 (N_14934,N_13146,N_13942);
or U14935 (N_14935,N_13425,N_13625);
or U14936 (N_14936,N_13504,N_13869);
or U14937 (N_14937,N_13319,N_13619);
xnor U14938 (N_14938,N_13783,N_13623);
xnor U14939 (N_14939,N_13043,N_13788);
or U14940 (N_14940,N_13751,N_13208);
or U14941 (N_14941,N_13014,N_13020);
xnor U14942 (N_14942,N_13708,N_13888);
and U14943 (N_14943,N_13734,N_13419);
nor U14944 (N_14944,N_13532,N_13004);
and U14945 (N_14945,N_13520,N_13784);
xor U14946 (N_14946,N_13685,N_13392);
xor U14947 (N_14947,N_13891,N_13573);
xor U14948 (N_14948,N_13933,N_13562);
nand U14949 (N_14949,N_13114,N_13640);
or U14950 (N_14950,N_13793,N_13871);
and U14951 (N_14951,N_13920,N_13895);
and U14952 (N_14952,N_13709,N_13459);
nor U14953 (N_14953,N_13130,N_13587);
nand U14954 (N_14954,N_13895,N_13647);
and U14955 (N_14955,N_13278,N_13379);
or U14956 (N_14956,N_13737,N_13228);
nand U14957 (N_14957,N_13157,N_13555);
nor U14958 (N_14958,N_13387,N_13260);
nand U14959 (N_14959,N_13849,N_13938);
xor U14960 (N_14960,N_13669,N_13374);
nand U14961 (N_14961,N_13112,N_13680);
nor U14962 (N_14962,N_13787,N_13196);
and U14963 (N_14963,N_13119,N_13852);
nand U14964 (N_14964,N_13915,N_13809);
or U14965 (N_14965,N_13214,N_13964);
nand U14966 (N_14966,N_13820,N_13566);
nand U14967 (N_14967,N_13719,N_13163);
xor U14968 (N_14968,N_13492,N_13871);
xnor U14969 (N_14969,N_13251,N_13180);
xor U14970 (N_14970,N_13191,N_13175);
nand U14971 (N_14971,N_13898,N_13714);
nor U14972 (N_14972,N_13212,N_13298);
nor U14973 (N_14973,N_13009,N_13073);
and U14974 (N_14974,N_13262,N_13257);
xnor U14975 (N_14975,N_13164,N_13342);
or U14976 (N_14976,N_13170,N_13500);
or U14977 (N_14977,N_13513,N_13325);
nand U14978 (N_14978,N_13365,N_13835);
xor U14979 (N_14979,N_13630,N_13919);
and U14980 (N_14980,N_13839,N_13556);
or U14981 (N_14981,N_13888,N_13900);
and U14982 (N_14982,N_13486,N_13302);
and U14983 (N_14983,N_13764,N_13508);
and U14984 (N_14984,N_13698,N_13461);
nand U14985 (N_14985,N_13487,N_13871);
and U14986 (N_14986,N_13068,N_13089);
and U14987 (N_14987,N_13263,N_13789);
or U14988 (N_14988,N_13200,N_13978);
and U14989 (N_14989,N_13370,N_13069);
or U14990 (N_14990,N_13591,N_13077);
xor U14991 (N_14991,N_13662,N_13425);
nand U14992 (N_14992,N_13409,N_13250);
nand U14993 (N_14993,N_13673,N_13913);
xor U14994 (N_14994,N_13418,N_13020);
nand U14995 (N_14995,N_13763,N_13585);
xor U14996 (N_14996,N_13371,N_13610);
nand U14997 (N_14997,N_13139,N_13778);
and U14998 (N_14998,N_13749,N_13010);
nand U14999 (N_14999,N_13567,N_13727);
nor U15000 (N_15000,N_14463,N_14048);
or U15001 (N_15001,N_14883,N_14067);
or U15002 (N_15002,N_14809,N_14217);
xnor U15003 (N_15003,N_14008,N_14066);
and U15004 (N_15004,N_14962,N_14475);
nand U15005 (N_15005,N_14150,N_14636);
and U15006 (N_15006,N_14671,N_14766);
and U15007 (N_15007,N_14509,N_14247);
and U15008 (N_15008,N_14496,N_14355);
nor U15009 (N_15009,N_14141,N_14874);
xor U15010 (N_15010,N_14910,N_14451);
xor U15011 (N_15011,N_14428,N_14801);
nand U15012 (N_15012,N_14591,N_14711);
nor U15013 (N_15013,N_14612,N_14578);
nor U15014 (N_15014,N_14977,N_14710);
and U15015 (N_15015,N_14957,N_14269);
or U15016 (N_15016,N_14631,N_14569);
or U15017 (N_15017,N_14527,N_14658);
nor U15018 (N_15018,N_14167,N_14897);
or U15019 (N_15019,N_14972,N_14516);
nand U15020 (N_15020,N_14641,N_14727);
nor U15021 (N_15021,N_14948,N_14429);
and U15022 (N_15022,N_14168,N_14003);
and U15023 (N_15023,N_14486,N_14885);
nand U15024 (N_15024,N_14361,N_14354);
nand U15025 (N_15025,N_14925,N_14776);
nand U15026 (N_15026,N_14949,N_14637);
and U15027 (N_15027,N_14223,N_14615);
nor U15028 (N_15028,N_14552,N_14338);
xnor U15029 (N_15029,N_14876,N_14845);
xnor U15030 (N_15030,N_14622,N_14916);
nand U15031 (N_15031,N_14878,N_14126);
and U15032 (N_15032,N_14287,N_14781);
nor U15033 (N_15033,N_14915,N_14240);
xor U15034 (N_15034,N_14239,N_14387);
xnor U15035 (N_15035,N_14382,N_14100);
or U15036 (N_15036,N_14911,N_14785);
nand U15037 (N_15037,N_14861,N_14263);
and U15038 (N_15038,N_14480,N_14027);
nor U15039 (N_15039,N_14488,N_14155);
xnor U15040 (N_15040,N_14937,N_14335);
xnor U15041 (N_15041,N_14576,N_14495);
nand U15042 (N_15042,N_14314,N_14884);
or U15043 (N_15043,N_14396,N_14774);
xnor U15044 (N_15044,N_14905,N_14867);
nand U15045 (N_15045,N_14248,N_14843);
or U15046 (N_15046,N_14912,N_14819);
nor U15047 (N_15047,N_14933,N_14605);
and U15048 (N_15048,N_14865,N_14717);
and U15049 (N_15049,N_14097,N_14812);
and U15050 (N_15050,N_14246,N_14792);
or U15051 (N_15051,N_14392,N_14662);
or U15052 (N_15052,N_14198,N_14947);
or U15053 (N_15053,N_14805,N_14713);
xnor U15054 (N_15054,N_14857,N_14091);
nor U15055 (N_15055,N_14836,N_14318);
nor U15056 (N_15056,N_14252,N_14186);
xor U15057 (N_15057,N_14046,N_14336);
or U15058 (N_15058,N_14934,N_14259);
xnor U15059 (N_15059,N_14062,N_14136);
xor U15060 (N_15060,N_14148,N_14123);
xnor U15061 (N_15061,N_14329,N_14011);
nor U15062 (N_15062,N_14784,N_14006);
nor U15063 (N_15063,N_14386,N_14726);
and U15064 (N_15064,N_14230,N_14670);
or U15065 (N_15065,N_14852,N_14850);
and U15066 (N_15066,N_14096,N_14546);
nand U15067 (N_15067,N_14431,N_14600);
nand U15068 (N_15068,N_14903,N_14295);
nand U15069 (N_15069,N_14040,N_14459);
nand U15070 (N_15070,N_14364,N_14704);
nand U15071 (N_15071,N_14748,N_14778);
nor U15072 (N_15072,N_14729,N_14777);
and U15073 (N_15073,N_14630,N_14417);
nor U15074 (N_15074,N_14927,N_14731);
xnor U15075 (N_15075,N_14233,N_14004);
or U15076 (N_15076,N_14742,N_14242);
nand U15077 (N_15077,N_14427,N_14754);
or U15078 (N_15078,N_14807,N_14455);
nand U15079 (N_15079,N_14112,N_14362);
xnor U15080 (N_15080,N_14825,N_14026);
nor U15081 (N_15081,N_14675,N_14913);
nand U15082 (N_15082,N_14154,N_14465);
or U15083 (N_15083,N_14530,N_14732);
nor U15084 (N_15084,N_14288,N_14199);
nand U15085 (N_15085,N_14250,N_14697);
or U15086 (N_15086,N_14373,N_14452);
and U15087 (N_15087,N_14353,N_14558);
nand U15088 (N_15088,N_14178,N_14529);
and U15089 (N_15089,N_14325,N_14579);
nand U15090 (N_15090,N_14478,N_14402);
or U15091 (N_15091,N_14256,N_14620);
nor U15092 (N_15092,N_14661,N_14705);
nand U15093 (N_15093,N_14950,N_14310);
nor U15094 (N_15094,N_14871,N_14009);
and U15095 (N_15095,N_14038,N_14724);
or U15096 (N_15096,N_14660,N_14984);
or U15097 (N_15097,N_14739,N_14593);
nor U15098 (N_15098,N_14350,N_14497);
nor U15099 (N_15099,N_14179,N_14680);
xor U15100 (N_15100,N_14113,N_14177);
or U15101 (N_15101,N_14589,N_14623);
xnor U15102 (N_15102,N_14237,N_14370);
or U15103 (N_15103,N_14152,N_14059);
xnor U15104 (N_15104,N_14821,N_14592);
nand U15105 (N_15105,N_14110,N_14270);
and U15106 (N_15106,N_14088,N_14289);
nand U15107 (N_15107,N_14514,N_14831);
and U15108 (N_15108,N_14952,N_14360);
nor U15109 (N_15109,N_14818,N_14251);
nor U15110 (N_15110,N_14042,N_14944);
or U15111 (N_15111,N_14565,N_14235);
nand U15112 (N_15112,N_14290,N_14209);
nand U15113 (N_15113,N_14722,N_14941);
and U15114 (N_15114,N_14121,N_14886);
nand U15115 (N_15115,N_14770,N_14526);
and U15116 (N_15116,N_14519,N_14545);
or U15117 (N_15117,N_14830,N_14063);
or U15118 (N_15118,N_14967,N_14868);
xnor U15119 (N_15119,N_14734,N_14752);
nor U15120 (N_15120,N_14855,N_14448);
and U15121 (N_15121,N_14371,N_14975);
nand U15122 (N_15122,N_14312,N_14320);
nand U15123 (N_15123,N_14982,N_14332);
nor U15124 (N_15124,N_14388,N_14577);
nor U15125 (N_15125,N_14932,N_14838);
or U15126 (N_15126,N_14438,N_14378);
nand U15127 (N_15127,N_14130,N_14163);
nand U15128 (N_15128,N_14033,N_14433);
xor U15129 (N_15129,N_14823,N_14306);
nand U15130 (N_15130,N_14049,N_14837);
and U15131 (N_15131,N_14512,N_14385);
and U15132 (N_15132,N_14134,N_14586);
xor U15133 (N_15133,N_14212,N_14566);
and U15134 (N_15134,N_14682,N_14559);
and U15135 (N_15135,N_14077,N_14162);
xnor U15136 (N_15136,N_14669,N_14173);
and U15137 (N_15137,N_14331,N_14880);
nor U15138 (N_15138,N_14634,N_14638);
and U15139 (N_15139,N_14639,N_14946);
and U15140 (N_15140,N_14347,N_14549);
or U15141 (N_15141,N_14583,N_14501);
xor U15142 (N_15142,N_14323,N_14460);
and U15143 (N_15143,N_14943,N_14745);
nor U15144 (N_15144,N_14833,N_14738);
nand U15145 (N_15145,N_14829,N_14089);
nor U15146 (N_15146,N_14842,N_14648);
and U15147 (N_15147,N_14442,N_14909);
nand U15148 (N_15148,N_14135,N_14513);
nor U15149 (N_15149,N_14069,N_14646);
xor U15150 (N_15150,N_14346,N_14317);
and U15151 (N_15151,N_14899,N_14220);
nand U15152 (N_15152,N_14339,N_14053);
or U15153 (N_15153,N_14344,N_14137);
nand U15154 (N_15154,N_14120,N_14720);
or U15155 (N_15155,N_14574,N_14917);
or U15156 (N_15156,N_14476,N_14951);
nand U15157 (N_15157,N_14298,N_14227);
xnor U15158 (N_15158,N_14036,N_14430);
and U15159 (N_15159,N_14504,N_14032);
nor U15160 (N_15160,N_14083,N_14188);
or U15161 (N_15161,N_14733,N_14743);
nor U15162 (N_15162,N_14606,N_14019);
nor U15163 (N_15163,N_14283,N_14305);
and U15164 (N_15164,N_14226,N_14201);
or U15165 (N_15165,N_14443,N_14065);
and U15166 (N_15166,N_14681,N_14816);
and U15167 (N_15167,N_14249,N_14893);
or U15168 (N_15168,N_14060,N_14002);
and U15169 (N_15169,N_14603,N_14128);
and U15170 (N_15170,N_14616,N_14632);
and U15171 (N_15171,N_14494,N_14324);
nand U15172 (N_15172,N_14158,N_14853);
nor U15173 (N_15173,N_14303,N_14342);
and U15174 (N_15174,N_14507,N_14587);
or U15175 (N_15175,N_14166,N_14222);
or U15176 (N_15176,N_14232,N_14528);
xnor U15177 (N_15177,N_14098,N_14993);
and U15178 (N_15178,N_14118,N_14117);
nor U15179 (N_15179,N_14755,N_14095);
xnor U15180 (N_15180,N_14462,N_14555);
and U15181 (N_15181,N_14231,N_14444);
nor U15182 (N_15182,N_14047,N_14081);
nor U15183 (N_15183,N_14441,N_14372);
xnor U15184 (N_15184,N_14763,N_14079);
nand U15185 (N_15185,N_14769,N_14300);
nor U15186 (N_15186,N_14706,N_14862);
or U15187 (N_15187,N_14034,N_14064);
nand U15188 (N_15188,N_14969,N_14481);
nand U15189 (N_15189,N_14258,N_14426);
xor U15190 (N_15190,N_14976,N_14928);
nand U15191 (N_15191,N_14692,N_14960);
or U15192 (N_15192,N_14881,N_14073);
xnor U15193 (N_15193,N_14992,N_14472);
and U15194 (N_15194,N_14918,N_14490);
nor U15195 (N_15195,N_14619,N_14759);
or U15196 (N_15196,N_14958,N_14534);
nor U15197 (N_15197,N_14389,N_14806);
or U15198 (N_15198,N_14010,N_14174);
nor U15199 (N_15199,N_14533,N_14169);
nand U15200 (N_15200,N_14058,N_14543);
or U15201 (N_15201,N_14018,N_14892);
nand U15202 (N_15202,N_14890,N_14072);
xnor U15203 (N_15203,N_14985,N_14684);
or U15204 (N_15204,N_14326,N_14815);
nand U15205 (N_15205,N_14989,N_14075);
nand U15206 (N_15206,N_14687,N_14275);
and U15207 (N_15207,N_14464,N_14959);
nor U15208 (N_15208,N_14521,N_14557);
xnor U15209 (N_15209,N_14030,N_14416);
nor U15210 (N_15210,N_14103,N_14847);
xnor U15211 (N_15211,N_14735,N_14930);
nor U15212 (N_15212,N_14409,N_14707);
nand U15213 (N_15213,N_14453,N_14919);
nand U15214 (N_15214,N_14856,N_14202);
or U15215 (N_15215,N_14377,N_14802);
nand U15216 (N_15216,N_14359,N_14206);
or U15217 (N_15217,N_14293,N_14111);
xnor U15218 (N_15218,N_14786,N_14550);
nor U15219 (N_15219,N_14257,N_14278);
or U15220 (N_15220,N_14413,N_14834);
xor U15221 (N_15221,N_14243,N_14765);
nand U15222 (N_15222,N_14824,N_14470);
nand U15223 (N_15223,N_14037,N_14974);
or U15224 (N_15224,N_14085,N_14654);
nand U15225 (N_15225,N_14477,N_14092);
and U15226 (N_15226,N_14554,N_14466);
nand U15227 (N_15227,N_14689,N_14594);
and U15228 (N_15228,N_14425,N_14160);
and U15229 (N_15229,N_14125,N_14194);
nand U15230 (N_15230,N_14891,N_14045);
or U15231 (N_15231,N_14285,N_14983);
or U15232 (N_15232,N_14510,N_14653);
nor U15233 (N_15233,N_14189,N_14832);
xnor U15234 (N_15234,N_14780,N_14375);
nand U15235 (N_15235,N_14645,N_14716);
nor U15236 (N_15236,N_14449,N_14624);
and U15237 (N_15237,N_14633,N_14151);
nand U15238 (N_15238,N_14800,N_14467);
or U15239 (N_15239,N_14261,N_14115);
xnor U15240 (N_15240,N_14422,N_14907);
or U15241 (N_15241,N_14536,N_14159);
nand U15242 (N_15242,N_14888,N_14568);
and U15243 (N_15243,N_14419,N_14381);
or U15244 (N_15244,N_14082,N_14399);
and U15245 (N_15245,N_14954,N_14817);
xor U15246 (N_15246,N_14228,N_14695);
nor U15247 (N_15247,N_14175,N_14216);
xor U15248 (N_15248,N_14268,N_14170);
or U15249 (N_15249,N_14181,N_14445);
nand U15250 (N_15250,N_14562,N_14408);
or U15251 (N_15251,N_14914,N_14213);
nor U15252 (N_15252,N_14119,N_14548);
nand U15253 (N_15253,N_14628,N_14254);
and U15254 (N_15254,N_14608,N_14221);
nor U15255 (N_15255,N_14980,N_14978);
and U15256 (N_15256,N_14182,N_14901);
nor U15257 (N_15257,N_14651,N_14436);
nor U15258 (N_15258,N_14281,N_14635);
nand U15259 (N_15259,N_14798,N_14998);
nor U15260 (N_15260,N_14099,N_14407);
or U15261 (N_15261,N_14921,N_14652);
and U15262 (N_15262,N_14761,N_14005);
xor U15263 (N_15263,N_14677,N_14374);
nand U15264 (N_15264,N_14393,N_14538);
or U15265 (N_15265,N_14524,N_14647);
and U15266 (N_15266,N_14506,N_14939);
nor U15267 (N_15267,N_14650,N_14328);
and U15268 (N_15268,N_14986,N_14043);
nand U15269 (N_15269,N_14076,N_14403);
nand U15270 (N_15270,N_14563,N_14573);
xnor U15271 (N_15271,N_14351,N_14601);
xor U15272 (N_15272,N_14851,N_14762);
xor U15273 (N_15273,N_14035,N_14410);
nand U15274 (N_15274,N_14297,N_14284);
nand U15275 (N_15275,N_14703,N_14185);
nor U15276 (N_15276,N_14023,N_14340);
and U15277 (N_15277,N_14165,N_14797);
xnor U15278 (N_15278,N_14094,N_14561);
xor U15279 (N_15279,N_14074,N_14813);
and U15280 (N_15280,N_14788,N_14904);
xor U15281 (N_15281,N_14013,N_14757);
xor U15282 (N_15282,N_14691,N_14145);
nor U15283 (N_15283,N_14302,N_14966);
nor U15284 (N_15284,N_14531,N_14143);
or U15285 (N_15285,N_14725,N_14255);
nand U15286 (N_15286,N_14187,N_14588);
or U15287 (N_15287,N_14979,N_14981);
xnor U15288 (N_15288,N_14747,N_14610);
and U15289 (N_15289,N_14101,N_14668);
or U15290 (N_15290,N_14124,N_14811);
or U15291 (N_15291,N_14491,N_14301);
xnor U15292 (N_15292,N_14663,N_14995);
or U15293 (N_15293,N_14087,N_14746);
or U15294 (N_15294,N_14511,N_14022);
and U15295 (N_15295,N_14363,N_14398);
and U15296 (N_15296,N_14487,N_14183);
xnor U15297 (N_15297,N_14349,N_14078);
or U15298 (N_15298,N_14493,N_14712);
nor U15299 (N_15299,N_14207,N_14860);
xor U15300 (N_15300,N_14728,N_14469);
xnor U15301 (N_15301,N_14142,N_14191);
nor U15302 (N_15302,N_14029,N_14196);
xnor U15303 (N_15303,N_14582,N_14820);
or U15304 (N_15304,N_14280,N_14996);
xor U15305 (N_15305,N_14131,N_14471);
and U15306 (N_15306,N_14054,N_14211);
nand U15307 (N_15307,N_14515,N_14322);
xor U15308 (N_15308,N_14474,N_14840);
nand U15309 (N_15309,N_14334,N_14107);
nor U15310 (N_15310,N_14935,N_14241);
or U15311 (N_15311,N_14454,N_14773);
xor U15312 (N_15312,N_14693,N_14315);
nor U15313 (N_15313,N_14758,N_14750);
nor U15314 (N_15314,N_14938,N_14642);
nand U15315 (N_15315,N_14849,N_14420);
xnor U15316 (N_15316,N_14676,N_14764);
or U15317 (N_15317,N_14313,N_14597);
xnor U15318 (N_15318,N_14994,N_14024);
xnor U15319 (N_15319,N_14584,N_14551);
xnor U15320 (N_15320,N_14139,N_14873);
xnor U15321 (N_15321,N_14744,N_14896);
nor U15322 (N_15322,N_14936,N_14379);
or U15323 (N_15323,N_14879,N_14180);
xor U15324 (N_15324,N_14990,N_14685);
xor U15325 (N_15325,N_14266,N_14264);
nand U15326 (N_15326,N_14376,N_14140);
or U15327 (N_15327,N_14595,N_14276);
nand U15328 (N_15328,N_14015,N_14737);
and U15329 (N_15329,N_14394,N_14423);
or U15330 (N_15330,N_14391,N_14138);
or U15331 (N_15331,N_14395,N_14204);
xor U15332 (N_15332,N_14133,N_14795);
and U15333 (N_15333,N_14749,N_14790);
nor U15334 (N_15334,N_14869,N_14014);
nand U15335 (N_15335,N_14380,N_14304);
or U15336 (N_15336,N_14665,N_14614);
xnor U15337 (N_15337,N_14730,N_14644);
nor U15338 (N_15338,N_14157,N_14193);
nand U15339 (N_15339,N_14659,N_14017);
nand U15340 (N_15340,N_14782,N_14768);
and U15341 (N_15341,N_14236,N_14457);
nor U15342 (N_15342,N_14352,N_14225);
nor U15343 (N_15343,N_14841,N_14068);
xor U15344 (N_15344,N_14090,N_14424);
xor U15345 (N_15345,N_14721,N_14702);
and U15346 (N_15346,N_14215,N_14564);
xor U15347 (N_15347,N_14719,N_14116);
and U15348 (N_15348,N_14963,N_14343);
nor U15349 (N_15349,N_14508,N_14229);
nand U15350 (N_15350,N_14277,N_14894);
and U15351 (N_15351,N_14200,N_14520);
nand U15352 (N_15352,N_14699,N_14205);
and U15353 (N_15353,N_14356,N_14238);
xor U15354 (N_15354,N_14787,N_14522);
nand U15355 (N_15355,N_14771,N_14964);
or U15356 (N_15356,N_14105,N_14794);
nor U15357 (N_15357,N_14596,N_14643);
or U15358 (N_15358,N_14122,N_14922);
nand U15359 (N_15359,N_14369,N_14330);
nor U15360 (N_15360,N_14626,N_14826);
and U15361 (N_15361,N_14299,N_14144);
xor U15362 (N_15362,N_14482,N_14505);
and U15363 (N_15363,N_14146,N_14108);
or U15364 (N_15364,N_14450,N_14708);
nor U15365 (N_15365,N_14827,N_14655);
xnor U15366 (N_15366,N_14560,N_14412);
nor U15367 (N_15367,N_14197,N_14253);
nor U15368 (N_15368,N_14106,N_14273);
or U15369 (N_15369,N_14499,N_14000);
nor U15370 (N_15370,N_14208,N_14822);
xor U15371 (N_15371,N_14102,N_14674);
xnor U15372 (N_15372,N_14164,N_14859);
nand U15373 (N_15373,N_14908,N_14945);
xnor U15374 (N_15374,N_14940,N_14052);
nor U15375 (N_15375,N_14999,N_14629);
xnor U15376 (N_15376,N_14598,N_14244);
nor U15377 (N_15377,N_14171,N_14321);
and U15378 (N_15378,N_14673,N_14988);
nand U15379 (N_15379,N_14846,N_14664);
or U15380 (N_15380,N_14542,N_14070);
and U15381 (N_15381,N_14924,N_14400);
xnor U15382 (N_15382,N_14872,N_14666);
nor U15383 (N_15383,N_14814,N_14541);
and U15384 (N_15384,N_14698,N_14153);
nand U15385 (N_15385,N_14955,N_14736);
xnor U15386 (N_15386,N_14599,N_14532);
and U15387 (N_15387,N_14751,N_14055);
xnor U15388 (N_15388,N_14319,N_14683);
or U15389 (N_15389,N_14411,N_14585);
nor U15390 (N_15390,N_14617,N_14882);
nand U15391 (N_15391,N_14556,N_14953);
and U15392 (N_15392,N_14265,N_14741);
nor U15393 (N_15393,N_14149,N_14923);
nand U15394 (N_15394,N_14877,N_14390);
nand U15395 (N_15395,N_14518,N_14437);
nor U15396 (N_15396,N_14456,N_14753);
or U15397 (N_15397,N_14001,N_14678);
xor U15398 (N_15398,N_14084,N_14621);
and U15399 (N_15399,N_14272,N_14071);
and U15400 (N_15400,N_14970,N_14640);
and U15401 (N_15401,N_14649,N_14050);
xor U15402 (N_15402,N_14041,N_14929);
xnor U15403 (N_15403,N_14129,N_14895);
or U15404 (N_15404,N_14114,N_14291);
and U15405 (N_15405,N_14889,N_14657);
nor U15406 (N_15406,N_14061,N_14973);
nand U15407 (N_15407,N_14971,N_14544);
and U15408 (N_15408,N_14618,N_14828);
or U15409 (N_15409,N_14613,N_14580);
or U15410 (N_15410,N_14961,N_14808);
or U15411 (N_15411,N_14161,N_14432);
or U15412 (N_15412,N_14709,N_14447);
xnor U15413 (N_15413,N_14367,N_14540);
nor U15414 (N_15414,N_14537,N_14492);
xor U15415 (N_15415,N_14421,N_14345);
nor U15416 (N_15416,N_14686,N_14926);
nand U15417 (N_15417,N_14931,N_14234);
nand U15418 (N_15418,N_14775,N_14575);
and U15419 (N_15419,N_14415,N_14348);
and U15420 (N_15420,N_14920,N_14218);
or U15421 (N_15421,N_14357,N_14854);
nor U15422 (N_15422,N_14740,N_14906);
nand U15423 (N_15423,N_14311,N_14461);
nor U15424 (N_15424,N_14274,N_14523);
nand U15425 (N_15425,N_14296,N_14397);
nand U15426 (N_15426,N_14844,N_14016);
and U15427 (N_15427,N_14696,N_14760);
or U15428 (N_15428,N_14767,N_14479);
or U15429 (N_15429,N_14690,N_14987);
nor U15430 (N_15430,N_14245,N_14127);
nor U15431 (N_15431,N_14309,N_14271);
nand U15432 (N_15432,N_14021,N_14203);
xnor U15433 (N_15433,N_14864,N_14679);
xnor U15434 (N_15434,N_14571,N_14500);
xnor U15435 (N_15435,N_14366,N_14219);
nand U15436 (N_15436,N_14570,N_14965);
or U15437 (N_15437,N_14418,N_14991);
or U15438 (N_15438,N_14887,N_14404);
and U15439 (N_15439,N_14789,N_14547);
nor U15440 (N_15440,N_14866,N_14956);
or U15441 (N_15441,N_14484,N_14756);
or U15442 (N_15442,N_14525,N_14405);
nand U15443 (N_15443,N_14810,N_14384);
nor U15444 (N_15444,N_14093,N_14609);
xnor U15445 (N_15445,N_14104,N_14156);
or U15446 (N_15446,N_14875,N_14132);
nand U15447 (N_15447,N_14383,N_14718);
xnor U15448 (N_15448,N_14485,N_14406);
xnor U15449 (N_15449,N_14656,N_14553);
and U15450 (N_15450,N_14667,N_14799);
or U15451 (N_15451,N_14688,N_14715);
nand U15452 (N_15452,N_14056,N_14031);
xor U15453 (N_15453,N_14517,N_14368);
and U15454 (N_15454,N_14192,N_14473);
xnor U15455 (N_15455,N_14458,N_14468);
and U15456 (N_15456,N_14316,N_14292);
and U15457 (N_15457,N_14333,N_14604);
or U15458 (N_15458,N_14898,N_14414);
or U15459 (N_15459,N_14701,N_14870);
and U15460 (N_15460,N_14307,N_14435);
and U15461 (N_15461,N_14900,N_14308);
nor U15462 (N_15462,N_14365,N_14007);
nor U15463 (N_15463,N_14434,N_14086);
xor U15464 (N_15464,N_14147,N_14341);
and U15465 (N_15465,N_14858,N_14942);
nand U15466 (N_15466,N_14224,N_14080);
and U15467 (N_15467,N_14439,N_14627);
and U15468 (N_15468,N_14779,N_14803);
and U15469 (N_15469,N_14997,N_14195);
or U15470 (N_15470,N_14286,N_14539);
and U15471 (N_15471,N_14176,N_14210);
nor U15472 (N_15472,N_14723,N_14793);
nand U15473 (N_15473,N_14489,N_14611);
xnor U15474 (N_15474,N_14863,N_14968);
nand U15475 (N_15475,N_14184,N_14502);
nor U15476 (N_15476,N_14572,N_14012);
and U15477 (N_15477,N_14057,N_14498);
xnor U15478 (N_15478,N_14327,N_14051);
or U15479 (N_15479,N_14279,N_14440);
xnor U15480 (N_15480,N_14791,N_14700);
or U15481 (N_15481,N_14028,N_14190);
xor U15482 (N_15482,N_14020,N_14039);
nand U15483 (N_15483,N_14602,N_14044);
xnor U15484 (N_15484,N_14109,N_14590);
nor U15485 (N_15485,N_14567,N_14446);
nor U15486 (N_15486,N_14262,N_14214);
nor U15487 (N_15487,N_14839,N_14672);
and U15488 (N_15488,N_14294,N_14401);
or U15489 (N_15489,N_14902,N_14772);
nand U15490 (N_15490,N_14694,N_14535);
nand U15491 (N_15491,N_14607,N_14625);
and U15492 (N_15492,N_14172,N_14796);
and U15493 (N_15493,N_14848,N_14358);
and U15494 (N_15494,N_14804,N_14503);
or U15495 (N_15495,N_14025,N_14835);
nor U15496 (N_15496,N_14337,N_14581);
nor U15497 (N_15497,N_14483,N_14267);
nor U15498 (N_15498,N_14260,N_14282);
and U15499 (N_15499,N_14783,N_14714);
xor U15500 (N_15500,N_14641,N_14920);
nand U15501 (N_15501,N_14057,N_14420);
or U15502 (N_15502,N_14038,N_14106);
nand U15503 (N_15503,N_14018,N_14009);
nand U15504 (N_15504,N_14927,N_14554);
or U15505 (N_15505,N_14953,N_14897);
nor U15506 (N_15506,N_14437,N_14662);
xnor U15507 (N_15507,N_14381,N_14616);
xnor U15508 (N_15508,N_14610,N_14953);
xnor U15509 (N_15509,N_14759,N_14486);
or U15510 (N_15510,N_14380,N_14077);
nand U15511 (N_15511,N_14465,N_14789);
and U15512 (N_15512,N_14830,N_14780);
or U15513 (N_15513,N_14519,N_14361);
and U15514 (N_15514,N_14933,N_14831);
and U15515 (N_15515,N_14711,N_14978);
nor U15516 (N_15516,N_14054,N_14736);
xnor U15517 (N_15517,N_14333,N_14680);
xor U15518 (N_15518,N_14907,N_14632);
xnor U15519 (N_15519,N_14495,N_14777);
or U15520 (N_15520,N_14123,N_14156);
and U15521 (N_15521,N_14957,N_14038);
and U15522 (N_15522,N_14245,N_14653);
xor U15523 (N_15523,N_14648,N_14051);
nand U15524 (N_15524,N_14478,N_14944);
nor U15525 (N_15525,N_14835,N_14448);
nor U15526 (N_15526,N_14475,N_14016);
or U15527 (N_15527,N_14641,N_14007);
and U15528 (N_15528,N_14659,N_14077);
xor U15529 (N_15529,N_14011,N_14388);
nand U15530 (N_15530,N_14673,N_14587);
nand U15531 (N_15531,N_14969,N_14838);
nor U15532 (N_15532,N_14260,N_14675);
nor U15533 (N_15533,N_14796,N_14279);
or U15534 (N_15534,N_14847,N_14204);
and U15535 (N_15535,N_14361,N_14839);
or U15536 (N_15536,N_14189,N_14984);
nand U15537 (N_15537,N_14574,N_14655);
or U15538 (N_15538,N_14354,N_14452);
xnor U15539 (N_15539,N_14079,N_14251);
or U15540 (N_15540,N_14734,N_14156);
nor U15541 (N_15541,N_14325,N_14072);
or U15542 (N_15542,N_14819,N_14036);
and U15543 (N_15543,N_14782,N_14891);
or U15544 (N_15544,N_14498,N_14868);
and U15545 (N_15545,N_14200,N_14068);
xor U15546 (N_15546,N_14590,N_14646);
xnor U15547 (N_15547,N_14662,N_14527);
or U15548 (N_15548,N_14870,N_14358);
and U15549 (N_15549,N_14821,N_14904);
nand U15550 (N_15550,N_14960,N_14778);
xnor U15551 (N_15551,N_14244,N_14039);
or U15552 (N_15552,N_14196,N_14201);
or U15553 (N_15553,N_14744,N_14163);
and U15554 (N_15554,N_14190,N_14376);
nand U15555 (N_15555,N_14097,N_14419);
xor U15556 (N_15556,N_14677,N_14315);
xnor U15557 (N_15557,N_14738,N_14633);
and U15558 (N_15558,N_14233,N_14187);
or U15559 (N_15559,N_14971,N_14755);
nor U15560 (N_15560,N_14209,N_14246);
xnor U15561 (N_15561,N_14522,N_14674);
and U15562 (N_15562,N_14481,N_14851);
or U15563 (N_15563,N_14111,N_14663);
and U15564 (N_15564,N_14218,N_14811);
nor U15565 (N_15565,N_14448,N_14850);
and U15566 (N_15566,N_14628,N_14194);
xnor U15567 (N_15567,N_14641,N_14286);
and U15568 (N_15568,N_14886,N_14551);
nor U15569 (N_15569,N_14302,N_14925);
xor U15570 (N_15570,N_14044,N_14297);
and U15571 (N_15571,N_14629,N_14657);
nand U15572 (N_15572,N_14863,N_14126);
or U15573 (N_15573,N_14313,N_14082);
nor U15574 (N_15574,N_14429,N_14291);
xnor U15575 (N_15575,N_14580,N_14625);
nor U15576 (N_15576,N_14755,N_14128);
or U15577 (N_15577,N_14566,N_14466);
nand U15578 (N_15578,N_14520,N_14416);
xnor U15579 (N_15579,N_14928,N_14084);
or U15580 (N_15580,N_14050,N_14471);
nand U15581 (N_15581,N_14528,N_14669);
nor U15582 (N_15582,N_14473,N_14244);
and U15583 (N_15583,N_14893,N_14343);
nor U15584 (N_15584,N_14115,N_14372);
nand U15585 (N_15585,N_14365,N_14852);
or U15586 (N_15586,N_14676,N_14720);
xnor U15587 (N_15587,N_14938,N_14809);
or U15588 (N_15588,N_14353,N_14399);
or U15589 (N_15589,N_14377,N_14579);
nor U15590 (N_15590,N_14299,N_14669);
or U15591 (N_15591,N_14801,N_14609);
and U15592 (N_15592,N_14625,N_14708);
or U15593 (N_15593,N_14111,N_14400);
nor U15594 (N_15594,N_14828,N_14431);
or U15595 (N_15595,N_14741,N_14536);
nand U15596 (N_15596,N_14772,N_14694);
xor U15597 (N_15597,N_14793,N_14208);
nor U15598 (N_15598,N_14867,N_14292);
or U15599 (N_15599,N_14817,N_14443);
or U15600 (N_15600,N_14327,N_14014);
or U15601 (N_15601,N_14191,N_14774);
xnor U15602 (N_15602,N_14377,N_14784);
or U15603 (N_15603,N_14666,N_14814);
nor U15604 (N_15604,N_14435,N_14824);
xnor U15605 (N_15605,N_14524,N_14207);
or U15606 (N_15606,N_14103,N_14891);
nor U15607 (N_15607,N_14484,N_14357);
and U15608 (N_15608,N_14501,N_14228);
or U15609 (N_15609,N_14567,N_14712);
xor U15610 (N_15610,N_14612,N_14994);
and U15611 (N_15611,N_14189,N_14058);
nand U15612 (N_15612,N_14674,N_14082);
and U15613 (N_15613,N_14839,N_14849);
nand U15614 (N_15614,N_14957,N_14134);
or U15615 (N_15615,N_14058,N_14208);
xor U15616 (N_15616,N_14106,N_14926);
nor U15617 (N_15617,N_14510,N_14103);
xnor U15618 (N_15618,N_14000,N_14832);
nor U15619 (N_15619,N_14880,N_14292);
or U15620 (N_15620,N_14456,N_14497);
or U15621 (N_15621,N_14718,N_14375);
nand U15622 (N_15622,N_14585,N_14492);
xor U15623 (N_15623,N_14760,N_14117);
and U15624 (N_15624,N_14182,N_14857);
nand U15625 (N_15625,N_14837,N_14249);
nor U15626 (N_15626,N_14815,N_14047);
or U15627 (N_15627,N_14139,N_14158);
or U15628 (N_15628,N_14432,N_14582);
xor U15629 (N_15629,N_14530,N_14891);
and U15630 (N_15630,N_14714,N_14352);
nand U15631 (N_15631,N_14249,N_14215);
nand U15632 (N_15632,N_14761,N_14408);
or U15633 (N_15633,N_14548,N_14100);
and U15634 (N_15634,N_14855,N_14563);
xnor U15635 (N_15635,N_14991,N_14823);
nand U15636 (N_15636,N_14677,N_14349);
or U15637 (N_15637,N_14900,N_14365);
and U15638 (N_15638,N_14690,N_14682);
xnor U15639 (N_15639,N_14185,N_14504);
or U15640 (N_15640,N_14445,N_14757);
or U15641 (N_15641,N_14645,N_14504);
xnor U15642 (N_15642,N_14294,N_14246);
and U15643 (N_15643,N_14715,N_14530);
and U15644 (N_15644,N_14812,N_14820);
and U15645 (N_15645,N_14579,N_14831);
nand U15646 (N_15646,N_14422,N_14064);
or U15647 (N_15647,N_14599,N_14622);
nand U15648 (N_15648,N_14091,N_14711);
or U15649 (N_15649,N_14575,N_14750);
nor U15650 (N_15650,N_14986,N_14454);
xnor U15651 (N_15651,N_14620,N_14614);
nand U15652 (N_15652,N_14705,N_14289);
or U15653 (N_15653,N_14071,N_14548);
or U15654 (N_15654,N_14497,N_14529);
nor U15655 (N_15655,N_14604,N_14265);
or U15656 (N_15656,N_14015,N_14183);
nor U15657 (N_15657,N_14103,N_14098);
nand U15658 (N_15658,N_14728,N_14751);
xor U15659 (N_15659,N_14746,N_14256);
nand U15660 (N_15660,N_14381,N_14720);
nand U15661 (N_15661,N_14380,N_14341);
xor U15662 (N_15662,N_14843,N_14207);
nand U15663 (N_15663,N_14006,N_14866);
xnor U15664 (N_15664,N_14119,N_14986);
nand U15665 (N_15665,N_14157,N_14152);
xnor U15666 (N_15666,N_14237,N_14423);
or U15667 (N_15667,N_14426,N_14517);
nand U15668 (N_15668,N_14351,N_14625);
xor U15669 (N_15669,N_14712,N_14814);
and U15670 (N_15670,N_14718,N_14142);
xnor U15671 (N_15671,N_14865,N_14353);
nand U15672 (N_15672,N_14125,N_14388);
nand U15673 (N_15673,N_14586,N_14493);
and U15674 (N_15674,N_14523,N_14322);
xor U15675 (N_15675,N_14232,N_14995);
or U15676 (N_15676,N_14307,N_14052);
xnor U15677 (N_15677,N_14933,N_14131);
or U15678 (N_15678,N_14042,N_14787);
and U15679 (N_15679,N_14623,N_14683);
nand U15680 (N_15680,N_14682,N_14132);
or U15681 (N_15681,N_14676,N_14058);
or U15682 (N_15682,N_14966,N_14866);
and U15683 (N_15683,N_14856,N_14500);
xor U15684 (N_15684,N_14953,N_14969);
and U15685 (N_15685,N_14423,N_14493);
nor U15686 (N_15686,N_14985,N_14181);
xor U15687 (N_15687,N_14562,N_14810);
nor U15688 (N_15688,N_14588,N_14368);
nor U15689 (N_15689,N_14353,N_14337);
or U15690 (N_15690,N_14195,N_14230);
xnor U15691 (N_15691,N_14183,N_14047);
and U15692 (N_15692,N_14098,N_14304);
nor U15693 (N_15693,N_14484,N_14282);
or U15694 (N_15694,N_14941,N_14297);
xor U15695 (N_15695,N_14396,N_14076);
and U15696 (N_15696,N_14614,N_14222);
nor U15697 (N_15697,N_14233,N_14640);
nor U15698 (N_15698,N_14448,N_14635);
nor U15699 (N_15699,N_14695,N_14262);
or U15700 (N_15700,N_14880,N_14936);
nor U15701 (N_15701,N_14174,N_14052);
or U15702 (N_15702,N_14904,N_14976);
nor U15703 (N_15703,N_14337,N_14115);
nor U15704 (N_15704,N_14587,N_14624);
and U15705 (N_15705,N_14058,N_14352);
xor U15706 (N_15706,N_14384,N_14778);
and U15707 (N_15707,N_14453,N_14479);
nand U15708 (N_15708,N_14666,N_14771);
nand U15709 (N_15709,N_14881,N_14095);
or U15710 (N_15710,N_14623,N_14808);
and U15711 (N_15711,N_14097,N_14221);
and U15712 (N_15712,N_14194,N_14852);
nand U15713 (N_15713,N_14837,N_14706);
nand U15714 (N_15714,N_14296,N_14713);
nor U15715 (N_15715,N_14104,N_14175);
nand U15716 (N_15716,N_14657,N_14048);
xnor U15717 (N_15717,N_14020,N_14803);
and U15718 (N_15718,N_14909,N_14250);
xnor U15719 (N_15719,N_14248,N_14056);
xor U15720 (N_15720,N_14860,N_14442);
xor U15721 (N_15721,N_14119,N_14404);
and U15722 (N_15722,N_14396,N_14504);
xor U15723 (N_15723,N_14295,N_14614);
nor U15724 (N_15724,N_14409,N_14359);
and U15725 (N_15725,N_14386,N_14252);
xnor U15726 (N_15726,N_14003,N_14407);
and U15727 (N_15727,N_14975,N_14608);
nand U15728 (N_15728,N_14502,N_14426);
xnor U15729 (N_15729,N_14609,N_14909);
xor U15730 (N_15730,N_14810,N_14163);
and U15731 (N_15731,N_14599,N_14256);
nor U15732 (N_15732,N_14092,N_14778);
or U15733 (N_15733,N_14484,N_14832);
and U15734 (N_15734,N_14621,N_14894);
and U15735 (N_15735,N_14599,N_14566);
nand U15736 (N_15736,N_14493,N_14565);
nor U15737 (N_15737,N_14529,N_14493);
or U15738 (N_15738,N_14238,N_14267);
nor U15739 (N_15739,N_14956,N_14421);
nor U15740 (N_15740,N_14429,N_14830);
or U15741 (N_15741,N_14879,N_14603);
nand U15742 (N_15742,N_14965,N_14078);
and U15743 (N_15743,N_14955,N_14049);
nand U15744 (N_15744,N_14750,N_14701);
and U15745 (N_15745,N_14314,N_14239);
nand U15746 (N_15746,N_14961,N_14921);
xnor U15747 (N_15747,N_14840,N_14114);
xnor U15748 (N_15748,N_14214,N_14946);
or U15749 (N_15749,N_14108,N_14309);
or U15750 (N_15750,N_14642,N_14026);
and U15751 (N_15751,N_14276,N_14374);
or U15752 (N_15752,N_14325,N_14539);
and U15753 (N_15753,N_14275,N_14595);
nor U15754 (N_15754,N_14839,N_14691);
xor U15755 (N_15755,N_14175,N_14983);
xnor U15756 (N_15756,N_14665,N_14649);
xnor U15757 (N_15757,N_14511,N_14112);
and U15758 (N_15758,N_14166,N_14128);
nand U15759 (N_15759,N_14453,N_14113);
and U15760 (N_15760,N_14079,N_14541);
or U15761 (N_15761,N_14471,N_14853);
nor U15762 (N_15762,N_14378,N_14502);
nand U15763 (N_15763,N_14726,N_14890);
nand U15764 (N_15764,N_14657,N_14118);
xnor U15765 (N_15765,N_14262,N_14480);
nand U15766 (N_15766,N_14982,N_14261);
xnor U15767 (N_15767,N_14508,N_14641);
and U15768 (N_15768,N_14441,N_14481);
or U15769 (N_15769,N_14598,N_14948);
xor U15770 (N_15770,N_14727,N_14262);
xor U15771 (N_15771,N_14121,N_14572);
nand U15772 (N_15772,N_14444,N_14710);
and U15773 (N_15773,N_14585,N_14379);
and U15774 (N_15774,N_14047,N_14870);
xnor U15775 (N_15775,N_14354,N_14524);
or U15776 (N_15776,N_14005,N_14990);
xnor U15777 (N_15777,N_14819,N_14124);
or U15778 (N_15778,N_14498,N_14553);
and U15779 (N_15779,N_14335,N_14805);
nor U15780 (N_15780,N_14104,N_14457);
or U15781 (N_15781,N_14629,N_14125);
and U15782 (N_15782,N_14970,N_14866);
xor U15783 (N_15783,N_14968,N_14347);
nor U15784 (N_15784,N_14319,N_14118);
xor U15785 (N_15785,N_14988,N_14152);
nand U15786 (N_15786,N_14722,N_14094);
and U15787 (N_15787,N_14570,N_14581);
and U15788 (N_15788,N_14534,N_14684);
and U15789 (N_15789,N_14693,N_14911);
or U15790 (N_15790,N_14078,N_14375);
and U15791 (N_15791,N_14768,N_14340);
nand U15792 (N_15792,N_14167,N_14900);
xnor U15793 (N_15793,N_14261,N_14995);
nand U15794 (N_15794,N_14050,N_14612);
and U15795 (N_15795,N_14649,N_14011);
xor U15796 (N_15796,N_14714,N_14090);
nand U15797 (N_15797,N_14370,N_14502);
xnor U15798 (N_15798,N_14733,N_14845);
xor U15799 (N_15799,N_14845,N_14517);
nand U15800 (N_15800,N_14339,N_14076);
nand U15801 (N_15801,N_14665,N_14871);
nor U15802 (N_15802,N_14767,N_14635);
xor U15803 (N_15803,N_14699,N_14510);
nand U15804 (N_15804,N_14543,N_14714);
xor U15805 (N_15805,N_14371,N_14063);
nor U15806 (N_15806,N_14764,N_14249);
and U15807 (N_15807,N_14228,N_14796);
nor U15808 (N_15808,N_14336,N_14725);
and U15809 (N_15809,N_14388,N_14556);
xnor U15810 (N_15810,N_14647,N_14109);
nor U15811 (N_15811,N_14909,N_14345);
xor U15812 (N_15812,N_14606,N_14315);
nand U15813 (N_15813,N_14200,N_14610);
nor U15814 (N_15814,N_14086,N_14675);
xor U15815 (N_15815,N_14445,N_14995);
nand U15816 (N_15816,N_14134,N_14605);
nand U15817 (N_15817,N_14624,N_14181);
and U15818 (N_15818,N_14542,N_14048);
and U15819 (N_15819,N_14896,N_14713);
xnor U15820 (N_15820,N_14153,N_14391);
and U15821 (N_15821,N_14696,N_14065);
nor U15822 (N_15822,N_14826,N_14043);
nand U15823 (N_15823,N_14548,N_14021);
nor U15824 (N_15824,N_14030,N_14397);
nand U15825 (N_15825,N_14707,N_14543);
nand U15826 (N_15826,N_14201,N_14184);
nor U15827 (N_15827,N_14057,N_14447);
and U15828 (N_15828,N_14699,N_14693);
nor U15829 (N_15829,N_14306,N_14110);
nor U15830 (N_15830,N_14447,N_14066);
nand U15831 (N_15831,N_14796,N_14597);
and U15832 (N_15832,N_14643,N_14850);
nand U15833 (N_15833,N_14557,N_14037);
nor U15834 (N_15834,N_14476,N_14831);
or U15835 (N_15835,N_14384,N_14964);
xnor U15836 (N_15836,N_14312,N_14590);
xor U15837 (N_15837,N_14550,N_14540);
or U15838 (N_15838,N_14889,N_14437);
nor U15839 (N_15839,N_14399,N_14408);
xnor U15840 (N_15840,N_14281,N_14415);
and U15841 (N_15841,N_14320,N_14617);
or U15842 (N_15842,N_14553,N_14235);
xor U15843 (N_15843,N_14523,N_14784);
nor U15844 (N_15844,N_14846,N_14390);
xnor U15845 (N_15845,N_14754,N_14451);
xnor U15846 (N_15846,N_14665,N_14737);
and U15847 (N_15847,N_14388,N_14105);
nor U15848 (N_15848,N_14172,N_14121);
or U15849 (N_15849,N_14313,N_14774);
and U15850 (N_15850,N_14766,N_14663);
and U15851 (N_15851,N_14693,N_14904);
nor U15852 (N_15852,N_14714,N_14472);
and U15853 (N_15853,N_14159,N_14509);
xnor U15854 (N_15854,N_14401,N_14503);
xor U15855 (N_15855,N_14299,N_14346);
nand U15856 (N_15856,N_14784,N_14246);
nand U15857 (N_15857,N_14090,N_14176);
and U15858 (N_15858,N_14302,N_14669);
or U15859 (N_15859,N_14330,N_14869);
and U15860 (N_15860,N_14282,N_14486);
and U15861 (N_15861,N_14948,N_14664);
xor U15862 (N_15862,N_14043,N_14195);
nor U15863 (N_15863,N_14706,N_14411);
nor U15864 (N_15864,N_14428,N_14282);
nor U15865 (N_15865,N_14849,N_14891);
nand U15866 (N_15866,N_14097,N_14397);
or U15867 (N_15867,N_14709,N_14242);
xnor U15868 (N_15868,N_14625,N_14791);
and U15869 (N_15869,N_14795,N_14902);
nand U15870 (N_15870,N_14805,N_14230);
and U15871 (N_15871,N_14637,N_14335);
nor U15872 (N_15872,N_14001,N_14029);
nand U15873 (N_15873,N_14624,N_14120);
nand U15874 (N_15874,N_14664,N_14399);
nand U15875 (N_15875,N_14228,N_14262);
xnor U15876 (N_15876,N_14497,N_14525);
or U15877 (N_15877,N_14070,N_14499);
nand U15878 (N_15878,N_14700,N_14569);
nor U15879 (N_15879,N_14985,N_14913);
nand U15880 (N_15880,N_14185,N_14563);
xor U15881 (N_15881,N_14201,N_14227);
nor U15882 (N_15882,N_14334,N_14391);
xnor U15883 (N_15883,N_14694,N_14835);
xnor U15884 (N_15884,N_14583,N_14944);
nor U15885 (N_15885,N_14251,N_14276);
and U15886 (N_15886,N_14873,N_14461);
nor U15887 (N_15887,N_14200,N_14878);
xor U15888 (N_15888,N_14316,N_14364);
nor U15889 (N_15889,N_14547,N_14725);
nor U15890 (N_15890,N_14669,N_14028);
nor U15891 (N_15891,N_14439,N_14854);
and U15892 (N_15892,N_14717,N_14954);
and U15893 (N_15893,N_14780,N_14568);
or U15894 (N_15894,N_14347,N_14265);
or U15895 (N_15895,N_14871,N_14057);
or U15896 (N_15896,N_14992,N_14508);
nor U15897 (N_15897,N_14380,N_14611);
or U15898 (N_15898,N_14841,N_14502);
and U15899 (N_15899,N_14179,N_14193);
and U15900 (N_15900,N_14513,N_14199);
nor U15901 (N_15901,N_14819,N_14706);
xnor U15902 (N_15902,N_14383,N_14906);
or U15903 (N_15903,N_14479,N_14971);
or U15904 (N_15904,N_14708,N_14255);
or U15905 (N_15905,N_14835,N_14221);
nor U15906 (N_15906,N_14478,N_14915);
xnor U15907 (N_15907,N_14426,N_14055);
nand U15908 (N_15908,N_14861,N_14594);
or U15909 (N_15909,N_14011,N_14900);
and U15910 (N_15910,N_14078,N_14937);
and U15911 (N_15911,N_14130,N_14284);
and U15912 (N_15912,N_14292,N_14787);
nand U15913 (N_15913,N_14216,N_14546);
nor U15914 (N_15914,N_14414,N_14462);
nand U15915 (N_15915,N_14056,N_14819);
nor U15916 (N_15916,N_14451,N_14578);
nor U15917 (N_15917,N_14731,N_14589);
nand U15918 (N_15918,N_14598,N_14235);
and U15919 (N_15919,N_14672,N_14683);
or U15920 (N_15920,N_14059,N_14110);
nor U15921 (N_15921,N_14769,N_14469);
nand U15922 (N_15922,N_14134,N_14070);
and U15923 (N_15923,N_14195,N_14951);
or U15924 (N_15924,N_14083,N_14116);
nor U15925 (N_15925,N_14262,N_14539);
or U15926 (N_15926,N_14674,N_14373);
nor U15927 (N_15927,N_14979,N_14947);
nand U15928 (N_15928,N_14626,N_14507);
or U15929 (N_15929,N_14572,N_14373);
or U15930 (N_15930,N_14770,N_14088);
nand U15931 (N_15931,N_14795,N_14056);
xor U15932 (N_15932,N_14882,N_14360);
nand U15933 (N_15933,N_14977,N_14887);
or U15934 (N_15934,N_14728,N_14851);
and U15935 (N_15935,N_14487,N_14081);
nor U15936 (N_15936,N_14147,N_14504);
nor U15937 (N_15937,N_14065,N_14561);
xnor U15938 (N_15938,N_14964,N_14224);
or U15939 (N_15939,N_14289,N_14019);
nand U15940 (N_15940,N_14566,N_14791);
nand U15941 (N_15941,N_14743,N_14870);
xnor U15942 (N_15942,N_14888,N_14546);
or U15943 (N_15943,N_14048,N_14866);
nand U15944 (N_15944,N_14249,N_14167);
and U15945 (N_15945,N_14124,N_14519);
and U15946 (N_15946,N_14220,N_14429);
nand U15947 (N_15947,N_14824,N_14915);
xnor U15948 (N_15948,N_14024,N_14165);
nand U15949 (N_15949,N_14334,N_14413);
nand U15950 (N_15950,N_14517,N_14566);
nand U15951 (N_15951,N_14754,N_14282);
or U15952 (N_15952,N_14453,N_14648);
and U15953 (N_15953,N_14359,N_14300);
xnor U15954 (N_15954,N_14957,N_14817);
xor U15955 (N_15955,N_14938,N_14479);
or U15956 (N_15956,N_14874,N_14457);
or U15957 (N_15957,N_14642,N_14273);
nor U15958 (N_15958,N_14826,N_14324);
and U15959 (N_15959,N_14551,N_14737);
and U15960 (N_15960,N_14580,N_14685);
and U15961 (N_15961,N_14860,N_14610);
nor U15962 (N_15962,N_14847,N_14194);
or U15963 (N_15963,N_14115,N_14769);
and U15964 (N_15964,N_14341,N_14718);
and U15965 (N_15965,N_14303,N_14669);
xor U15966 (N_15966,N_14325,N_14081);
and U15967 (N_15967,N_14163,N_14098);
nand U15968 (N_15968,N_14851,N_14904);
xnor U15969 (N_15969,N_14674,N_14221);
and U15970 (N_15970,N_14278,N_14369);
and U15971 (N_15971,N_14224,N_14211);
or U15972 (N_15972,N_14225,N_14170);
xnor U15973 (N_15973,N_14499,N_14167);
nand U15974 (N_15974,N_14104,N_14580);
and U15975 (N_15975,N_14272,N_14130);
xor U15976 (N_15976,N_14675,N_14295);
or U15977 (N_15977,N_14654,N_14211);
and U15978 (N_15978,N_14394,N_14846);
nand U15979 (N_15979,N_14124,N_14354);
and U15980 (N_15980,N_14597,N_14959);
and U15981 (N_15981,N_14030,N_14840);
nand U15982 (N_15982,N_14181,N_14150);
nor U15983 (N_15983,N_14292,N_14249);
nor U15984 (N_15984,N_14310,N_14002);
or U15985 (N_15985,N_14052,N_14535);
and U15986 (N_15986,N_14094,N_14378);
or U15987 (N_15987,N_14118,N_14641);
nor U15988 (N_15988,N_14177,N_14643);
and U15989 (N_15989,N_14756,N_14509);
or U15990 (N_15990,N_14631,N_14381);
or U15991 (N_15991,N_14999,N_14621);
xor U15992 (N_15992,N_14926,N_14237);
or U15993 (N_15993,N_14490,N_14189);
or U15994 (N_15994,N_14532,N_14230);
or U15995 (N_15995,N_14471,N_14979);
xor U15996 (N_15996,N_14038,N_14817);
nand U15997 (N_15997,N_14315,N_14309);
or U15998 (N_15998,N_14639,N_14551);
or U15999 (N_15999,N_14123,N_14840);
and U16000 (N_16000,N_15984,N_15616);
or U16001 (N_16001,N_15046,N_15287);
nand U16002 (N_16002,N_15332,N_15681);
xor U16003 (N_16003,N_15222,N_15406);
nand U16004 (N_16004,N_15131,N_15313);
and U16005 (N_16005,N_15949,N_15037);
xor U16006 (N_16006,N_15108,N_15490);
nor U16007 (N_16007,N_15031,N_15898);
xor U16008 (N_16008,N_15404,N_15291);
nor U16009 (N_16009,N_15712,N_15646);
and U16010 (N_16010,N_15192,N_15893);
and U16011 (N_16011,N_15821,N_15415);
nor U16012 (N_16012,N_15755,N_15320);
nor U16013 (N_16013,N_15897,N_15628);
and U16014 (N_16014,N_15247,N_15564);
nand U16015 (N_16015,N_15118,N_15938);
or U16016 (N_16016,N_15358,N_15825);
xnor U16017 (N_16017,N_15075,N_15253);
or U16018 (N_16018,N_15030,N_15283);
nand U16019 (N_16019,N_15085,N_15877);
xor U16020 (N_16020,N_15610,N_15019);
xnor U16021 (N_16021,N_15289,N_15492);
nand U16022 (N_16022,N_15272,N_15922);
nand U16023 (N_16023,N_15117,N_15235);
xor U16024 (N_16024,N_15400,N_15625);
nor U16025 (N_16025,N_15782,N_15779);
xor U16026 (N_16026,N_15401,N_15070);
nand U16027 (N_16027,N_15660,N_15423);
or U16028 (N_16028,N_15630,N_15336);
or U16029 (N_16029,N_15501,N_15387);
or U16030 (N_16030,N_15953,N_15138);
nor U16031 (N_16031,N_15568,N_15839);
or U16032 (N_16032,N_15013,N_15134);
xor U16033 (N_16033,N_15209,N_15381);
or U16034 (N_16034,N_15029,N_15202);
xor U16035 (N_16035,N_15523,N_15986);
nor U16036 (N_16036,N_15964,N_15872);
nor U16037 (N_16037,N_15757,N_15484);
nor U16038 (N_16038,N_15974,N_15471);
nand U16039 (N_16039,N_15275,N_15833);
or U16040 (N_16040,N_15746,N_15337);
xnor U16041 (N_16041,N_15081,N_15560);
xnor U16042 (N_16042,N_15944,N_15852);
and U16043 (N_16043,N_15120,N_15677);
and U16044 (N_16044,N_15596,N_15014);
or U16045 (N_16045,N_15851,N_15142);
xnor U16046 (N_16046,N_15507,N_15215);
xnor U16047 (N_16047,N_15078,N_15301);
nor U16048 (N_16048,N_15856,N_15694);
nor U16049 (N_16049,N_15152,N_15583);
or U16050 (N_16050,N_15547,N_15655);
nand U16051 (N_16051,N_15649,N_15816);
xnor U16052 (N_16052,N_15060,N_15840);
and U16053 (N_16053,N_15052,N_15614);
xor U16054 (N_16054,N_15556,N_15334);
or U16055 (N_16055,N_15578,N_15505);
nor U16056 (N_16056,N_15742,N_15548);
nand U16057 (N_16057,N_15510,N_15359);
xor U16058 (N_16058,N_15457,N_15148);
nor U16059 (N_16059,N_15519,N_15563);
nor U16060 (N_16060,N_15561,N_15486);
or U16061 (N_16061,N_15074,N_15585);
xnor U16062 (N_16062,N_15865,N_15262);
and U16063 (N_16063,N_15092,N_15431);
xnor U16064 (N_16064,N_15213,N_15061);
xor U16065 (N_16065,N_15318,N_15673);
xor U16066 (N_16066,N_15443,N_15419);
or U16067 (N_16067,N_15808,N_15341);
nor U16068 (N_16068,N_15229,N_15708);
and U16069 (N_16069,N_15954,N_15239);
or U16070 (N_16070,N_15914,N_15803);
or U16071 (N_16071,N_15530,N_15996);
or U16072 (N_16072,N_15164,N_15819);
nand U16073 (N_16073,N_15424,N_15298);
nor U16074 (N_16074,N_15151,N_15991);
nor U16075 (N_16075,N_15770,N_15979);
nand U16076 (N_16076,N_15611,N_15663);
or U16077 (N_16077,N_15998,N_15043);
xor U16078 (N_16078,N_15088,N_15993);
nor U16079 (N_16079,N_15084,N_15985);
xnor U16080 (N_16080,N_15176,N_15141);
xnor U16081 (N_16081,N_15284,N_15943);
or U16082 (N_16082,N_15942,N_15714);
or U16083 (N_16083,N_15073,N_15269);
or U16084 (N_16084,N_15378,N_15474);
nand U16085 (N_16085,N_15144,N_15196);
or U16086 (N_16086,N_15410,N_15379);
xnor U16087 (N_16087,N_15089,N_15934);
xor U16088 (N_16088,N_15086,N_15408);
and U16089 (N_16089,N_15753,N_15296);
and U16090 (N_16090,N_15890,N_15704);
nor U16091 (N_16091,N_15157,N_15537);
or U16092 (N_16092,N_15465,N_15445);
xnor U16093 (N_16093,N_15399,N_15987);
xor U16094 (N_16094,N_15216,N_15180);
nand U16095 (N_16095,N_15121,N_15822);
nor U16096 (N_16096,N_15983,N_15003);
and U16097 (N_16097,N_15715,N_15606);
xnor U16098 (N_16098,N_15487,N_15231);
or U16099 (N_16099,N_15861,N_15766);
nor U16100 (N_16100,N_15475,N_15367);
xnor U16101 (N_16101,N_15693,N_15736);
xor U16102 (N_16102,N_15842,N_15689);
nor U16103 (N_16103,N_15347,N_15158);
nand U16104 (N_16104,N_15321,N_15838);
nand U16105 (N_16105,N_15754,N_15631);
and U16106 (N_16106,N_15188,N_15805);
nor U16107 (N_16107,N_15096,N_15559);
and U16108 (N_16108,N_15153,N_15896);
and U16109 (N_16109,N_15648,N_15163);
or U16110 (N_16110,N_15047,N_15807);
nor U16111 (N_16111,N_15421,N_15299);
or U16112 (N_16112,N_15133,N_15446);
nor U16113 (N_16113,N_15207,N_15128);
nor U16114 (N_16114,N_15385,N_15988);
nor U16115 (N_16115,N_15271,N_15187);
xnor U16116 (N_16116,N_15834,N_15869);
xnor U16117 (N_16117,N_15267,N_15069);
xor U16118 (N_16118,N_15867,N_15665);
xnor U16119 (N_16119,N_15668,N_15363);
xnor U16120 (N_16120,N_15442,N_15100);
and U16121 (N_16121,N_15224,N_15413);
or U16122 (N_16122,N_15077,N_15717);
and U16123 (N_16123,N_15126,N_15639);
and U16124 (N_16124,N_15016,N_15422);
or U16125 (N_16125,N_15217,N_15544);
or U16126 (N_16126,N_15863,N_15461);
and U16127 (N_16127,N_15554,N_15600);
nor U16128 (N_16128,N_15058,N_15438);
xnor U16129 (N_16129,N_15466,N_15258);
nand U16130 (N_16130,N_15909,N_15420);
and U16131 (N_16131,N_15377,N_15645);
nor U16132 (N_16132,N_15109,N_15590);
nor U16133 (N_16133,N_15039,N_15124);
and U16134 (N_16134,N_15908,N_15850);
and U16135 (N_16135,N_15875,N_15778);
nand U16136 (N_16136,N_15342,N_15254);
nand U16137 (N_16137,N_15620,N_15957);
xor U16138 (N_16138,N_15618,N_15835);
nand U16139 (N_16139,N_15509,N_15601);
or U16140 (N_16140,N_15023,N_15784);
and U16141 (N_16141,N_15558,N_15726);
xnor U16142 (N_16142,N_15703,N_15418);
nor U16143 (N_16143,N_15171,N_15670);
and U16144 (N_16144,N_15116,N_15436);
or U16145 (N_16145,N_15889,N_15885);
and U16146 (N_16146,N_15674,N_15278);
or U16147 (N_16147,N_15388,N_15727);
nor U16148 (N_16148,N_15178,N_15122);
xnor U16149 (N_16149,N_15064,N_15427);
nor U16150 (N_16150,N_15059,N_15405);
or U16151 (N_16151,N_15761,N_15691);
xor U16152 (N_16152,N_15550,N_15573);
or U16153 (N_16153,N_15302,N_15886);
or U16154 (N_16154,N_15608,N_15973);
and U16155 (N_16155,N_15728,N_15783);
and U16156 (N_16156,N_15053,N_15204);
nor U16157 (N_16157,N_15932,N_15903);
or U16158 (N_16158,N_15435,N_15488);
and U16159 (N_16159,N_15551,N_15522);
and U16160 (N_16160,N_15054,N_15102);
or U16161 (N_16161,N_15006,N_15305);
and U16162 (N_16162,N_15534,N_15552);
xor U16163 (N_16163,N_15426,N_15532);
nor U16164 (N_16164,N_15723,N_15653);
or U16165 (N_16165,N_15165,N_15351);
xnor U16166 (N_16166,N_15591,N_15658);
or U16167 (N_16167,N_15543,N_15276);
nor U16168 (N_16168,N_15915,N_15758);
or U16169 (N_16169,N_15651,N_15966);
nor U16170 (N_16170,N_15542,N_15925);
or U16171 (N_16171,N_15732,N_15748);
xor U16172 (N_16172,N_15469,N_15846);
nand U16173 (N_16173,N_15156,N_15963);
and U16174 (N_16174,N_15724,N_15273);
xor U16175 (N_16175,N_15429,N_15586);
nor U16176 (N_16176,N_15540,N_15478);
and U16177 (N_16177,N_15999,N_15393);
nand U16178 (N_16178,N_15190,N_15076);
and U16179 (N_16179,N_15967,N_15049);
and U16180 (N_16180,N_15259,N_15232);
and U16181 (N_16181,N_15604,N_15355);
nand U16182 (N_16182,N_15011,N_15268);
xnor U16183 (N_16183,N_15227,N_15323);
nand U16184 (N_16184,N_15022,N_15184);
and U16185 (N_16185,N_15666,N_15062);
nor U16186 (N_16186,N_15900,N_15883);
or U16187 (N_16187,N_15297,N_15961);
nor U16188 (N_16188,N_15773,N_15091);
nor U16189 (N_16189,N_15671,N_15437);
nor U16190 (N_16190,N_15769,N_15464);
or U16191 (N_16191,N_15661,N_15536);
nor U16192 (N_16192,N_15672,N_15786);
and U16193 (N_16193,N_15485,N_15647);
xor U16194 (N_16194,N_15170,N_15503);
nand U16195 (N_16195,N_15211,N_15495);
and U16196 (N_16196,N_15995,N_15114);
nand U16197 (N_16197,N_15292,N_15637);
nor U16198 (N_16198,N_15099,N_15506);
nor U16199 (N_16199,N_15981,N_15051);
nand U16200 (N_16200,N_15139,N_15855);
xnor U16201 (N_16201,N_15787,N_15449);
nor U16202 (N_16202,N_15680,N_15010);
nand U16203 (N_16203,N_15389,N_15894);
nor U16204 (N_16204,N_15252,N_15266);
or U16205 (N_16205,N_15725,N_15652);
and U16206 (N_16206,N_15945,N_15454);
xnor U16207 (N_16207,N_15132,N_15771);
xnor U16208 (N_16208,N_15310,N_15592);
or U16209 (N_16209,N_15166,N_15792);
nor U16210 (N_16210,N_15913,N_15172);
and U16211 (N_16211,N_15038,N_15360);
nand U16212 (N_16212,N_15160,N_15324);
or U16213 (N_16213,N_15033,N_15095);
and U16214 (N_16214,N_15588,N_15005);
nand U16215 (N_16215,N_15990,N_15582);
and U16216 (N_16216,N_15517,N_15179);
or U16217 (N_16217,N_15857,N_15854);
or U16218 (N_16218,N_15345,N_15312);
nor U16219 (N_16219,N_15391,N_15416);
nand U16220 (N_16220,N_15080,N_15626);
nand U16221 (N_16221,N_15828,N_15493);
nor U16222 (N_16222,N_15191,N_15907);
nand U16223 (N_16223,N_15975,N_15417);
nand U16224 (N_16224,N_15710,N_15526);
and U16225 (N_16225,N_15675,N_15001);
and U16226 (N_16226,N_15892,N_15669);
xor U16227 (N_16227,N_15304,N_15899);
xnor U16228 (N_16228,N_15498,N_15879);
nor U16229 (N_16229,N_15220,N_15319);
nor U16230 (N_16230,N_15214,N_15125);
nand U16231 (N_16231,N_15829,N_15881);
and U16232 (N_16232,N_15960,N_15226);
xnor U16233 (N_16233,N_15760,N_15901);
xnor U16234 (N_16234,N_15830,N_15237);
nor U16235 (N_16235,N_15386,N_15512);
and U16236 (N_16236,N_15477,N_15546);
nor U16237 (N_16237,N_15799,N_15845);
or U16238 (N_16238,N_15657,N_15994);
and U16239 (N_16239,N_15315,N_15968);
or U16240 (N_16240,N_15251,N_15448);
nor U16241 (N_16241,N_15848,N_15333);
nor U16242 (N_16242,N_15339,N_15440);
xnor U16243 (N_16243,N_15826,N_15814);
nand U16244 (N_16244,N_15679,N_15707);
xor U16245 (N_16245,N_15836,N_15776);
nor U16246 (N_16246,N_15844,N_15823);
nand U16247 (N_16247,N_15820,N_15200);
and U16248 (N_16248,N_15238,N_15884);
nand U16249 (N_16249,N_15240,N_15467);
nand U16250 (N_16250,N_15402,N_15831);
nand U16251 (N_16251,N_15941,N_15135);
or U16252 (N_16252,N_15571,N_15183);
or U16253 (N_16253,N_15127,N_15853);
nor U16254 (N_16254,N_15504,N_15702);
nor U16255 (N_16255,N_15162,N_15462);
and U16256 (N_16256,N_15765,N_15722);
or U16257 (N_16257,N_15939,N_15041);
xor U16258 (N_16258,N_15595,N_15093);
nor U16259 (N_16259,N_15260,N_15294);
nand U16260 (N_16260,N_15325,N_15699);
xor U16261 (N_16261,N_15380,N_15789);
and U16262 (N_16262,N_15577,N_15687);
nor U16263 (N_16263,N_15083,N_15300);
xnor U16264 (N_16264,N_15317,N_15434);
nor U16265 (N_16265,N_15514,N_15057);
nor U16266 (N_16266,N_15017,N_15228);
or U16267 (N_16267,N_15734,N_15000);
and U16268 (N_16268,N_15136,N_15303);
xnor U16269 (N_16269,N_15549,N_15221);
nor U16270 (N_16270,N_15911,N_15664);
or U16271 (N_16271,N_15801,N_15972);
nand U16272 (N_16272,N_15456,N_15891);
nor U16273 (N_16273,N_15264,N_15072);
or U16274 (N_16274,N_15982,N_15824);
or U16275 (N_16275,N_15015,N_15977);
and U16276 (N_16276,N_15640,N_15969);
nand U16277 (N_16277,N_15905,N_15432);
or U16278 (N_16278,N_15937,N_15201);
or U16279 (N_16279,N_15094,N_15212);
nor U16280 (N_16280,N_15644,N_15929);
and U16281 (N_16281,N_15567,N_15729);
nor U16282 (N_16282,N_15980,N_15871);
nand U16283 (N_16283,N_15880,N_15481);
nor U16284 (N_16284,N_15575,N_15101);
or U16285 (N_16285,N_15453,N_15926);
and U16286 (N_16286,N_15818,N_15887);
or U16287 (N_16287,N_15731,N_15739);
nand U16288 (N_16288,N_15344,N_15263);
or U16289 (N_16289,N_15622,N_15407);
xor U16290 (N_16290,N_15112,N_15804);
nand U16291 (N_16291,N_15690,N_15565);
xnor U16292 (N_16292,N_15793,N_15612);
nand U16293 (N_16293,N_15502,N_15027);
xor U16294 (N_16294,N_15107,N_15806);
nor U16295 (N_16295,N_15350,N_15809);
nor U16296 (N_16296,N_15018,N_15356);
or U16297 (N_16297,N_15810,N_15130);
or U16298 (N_16298,N_15912,N_15918);
nand U16299 (N_16299,N_15656,N_15572);
nor U16300 (N_16300,N_15225,N_15813);
and U16301 (N_16301,N_15230,N_15695);
nand U16302 (N_16302,N_15700,N_15615);
or U16303 (N_16303,N_15527,N_15412);
or U16304 (N_16304,N_15002,N_15357);
and U16305 (N_16305,N_15555,N_15397);
or U16306 (N_16306,N_15959,N_15322);
xnor U16307 (N_16307,N_15256,N_15638);
xnor U16308 (N_16308,N_15798,N_15489);
or U16309 (N_16309,N_15243,N_15286);
nand U16310 (N_16310,N_15439,N_15249);
or U16311 (N_16311,N_15459,N_15335);
or U16312 (N_16312,N_15643,N_15511);
nand U16313 (N_16313,N_15667,N_15827);
nor U16314 (N_16314,N_15686,N_15795);
nand U16315 (N_16315,N_15989,N_15012);
nand U16316 (N_16316,N_15716,N_15082);
xor U16317 (N_16317,N_15295,N_15390);
nand U16318 (N_16318,N_15352,N_15428);
nand U16319 (N_16319,N_15071,N_15433);
nand U16320 (N_16320,N_15520,N_15587);
nand U16321 (N_16321,N_15398,N_15696);
nor U16322 (N_16322,N_15521,N_15451);
nor U16323 (N_16323,N_15468,N_15065);
and U16324 (N_16324,N_15346,N_15870);
nand U16325 (N_16325,N_15594,N_15569);
xnor U16326 (N_16326,N_15790,N_15343);
nor U16327 (N_16327,N_15103,N_15182);
nor U16328 (N_16328,N_15067,N_15832);
or U16329 (N_16329,N_15045,N_15177);
nor U16330 (N_16330,N_15970,N_15603);
nand U16331 (N_16331,N_15692,N_15508);
nor U16332 (N_16332,N_15154,N_15411);
nand U16333 (N_16333,N_15307,N_15623);
and U16334 (N_16334,N_15785,N_15106);
or U16335 (N_16335,N_15167,N_15374);
nand U16336 (N_16336,N_15992,N_15328);
nor U16337 (N_16337,N_15329,N_15584);
or U16338 (N_16338,N_15425,N_15713);
nor U16339 (N_16339,N_15115,N_15617);
xor U16340 (N_16340,N_15876,N_15528);
nand U16341 (N_16341,N_15414,N_15524);
or U16342 (N_16342,N_15007,N_15950);
or U16343 (N_16343,N_15441,N_15483);
and U16344 (N_16344,N_15479,N_15137);
or U16345 (N_16345,N_15173,N_15340);
xnor U16346 (N_16346,N_15396,N_15598);
nand U16347 (N_16347,N_15035,N_15282);
and U16348 (N_16348,N_15032,N_15161);
and U16349 (N_16349,N_15633,N_15123);
xor U16350 (N_16350,N_15460,N_15208);
or U16351 (N_16351,N_15193,N_15175);
or U16352 (N_16352,N_15535,N_15409);
and U16353 (N_16353,N_15104,N_15372);
nand U16354 (N_16354,N_15186,N_15662);
nand U16355 (N_16355,N_15740,N_15730);
xnor U16356 (N_16356,N_15197,N_15858);
nand U16357 (N_16357,N_15920,N_15314);
xnor U16358 (N_16358,N_15233,N_15762);
nand U16359 (N_16359,N_15525,N_15910);
nand U16360 (N_16360,N_15494,N_15055);
nor U16361 (N_16361,N_15921,N_15709);
or U16362 (N_16362,N_15364,N_15491);
xnor U16363 (N_16363,N_15234,N_15366);
nand U16364 (N_16364,N_15923,N_15248);
or U16365 (N_16365,N_15290,N_15772);
nor U16366 (N_16366,N_15581,N_15203);
nor U16367 (N_16367,N_15634,N_15931);
or U16368 (N_16368,N_15750,N_15194);
nand U16369 (N_16369,N_15744,N_15129);
and U16370 (N_16370,N_15815,N_15198);
or U16371 (N_16371,N_15353,N_15553);
nor U16372 (N_16372,N_15745,N_15326);
nor U16373 (N_16373,N_15562,N_15538);
and U16374 (N_16374,N_15629,N_15794);
nand U16375 (N_16375,N_15895,N_15650);
and U16376 (N_16376,N_15997,N_15579);
xnor U16377 (N_16377,N_15864,N_15048);
or U16378 (N_16378,N_15497,N_15020);
and U16379 (N_16379,N_15607,N_15916);
or U16380 (N_16380,N_15371,N_15403);
nor U16381 (N_16381,N_15362,N_15955);
xnor U16382 (N_16382,N_15641,N_15306);
nor U16383 (N_16383,N_15447,N_15775);
xor U16384 (N_16384,N_15539,N_15159);
nand U16385 (N_16385,N_15008,N_15878);
nor U16386 (N_16386,N_15948,N_15338);
or U16387 (N_16387,N_15255,N_15150);
nand U16388 (N_16388,N_15309,N_15705);
nor U16389 (N_16389,N_15837,N_15654);
and U16390 (N_16390,N_15028,N_15580);
nand U16391 (N_16391,N_15919,N_15902);
xor U16392 (N_16392,N_15882,N_15682);
xnor U16393 (N_16393,N_15843,N_15529);
nor U16394 (N_16394,N_15155,N_15458);
nor U16395 (N_16395,N_15743,N_15450);
nand U16396 (N_16396,N_15956,N_15242);
nor U16397 (N_16397,N_15365,N_15802);
nand U16398 (N_16398,N_15145,N_15683);
and U16399 (N_16399,N_15361,N_15697);
nand U16400 (N_16400,N_15024,N_15257);
nor U16401 (N_16401,N_15597,N_15500);
and U16402 (N_16402,N_15330,N_15764);
xor U16403 (N_16403,N_15463,N_15797);
nand U16404 (N_16404,N_15951,N_15791);
or U16405 (N_16405,N_15383,N_15605);
or U16406 (N_16406,N_15349,N_15288);
nand U16407 (N_16407,N_15749,N_15574);
and U16408 (N_16408,N_15195,N_15777);
nor U16409 (N_16409,N_15004,N_15781);
and U16410 (N_16410,N_15499,N_15685);
xor U16411 (N_16411,N_15050,N_15040);
xnor U16412 (N_16412,N_15621,N_15531);
and U16413 (N_16413,N_15636,N_15533);
nor U16414 (N_16414,N_15025,N_15368);
nand U16415 (N_16415,N_15370,N_15245);
and U16416 (N_16416,N_15684,N_15143);
and U16417 (N_16417,N_15244,N_15168);
and U16418 (N_16418,N_15721,N_15455);
nor U16419 (N_16419,N_15706,N_15146);
and U16420 (N_16420,N_15090,N_15261);
nand U16421 (N_16421,N_15720,N_15009);
or U16422 (N_16422,N_15473,N_15768);
and U16423 (N_16423,N_15281,N_15589);
and U16424 (N_16424,N_15904,N_15788);
nor U16425 (N_16425,N_15241,N_15265);
nor U16426 (N_16426,N_15873,N_15952);
or U16427 (N_16427,N_15718,N_15635);
nand U16428 (N_16428,N_15541,N_15609);
and U16429 (N_16429,N_15936,N_15888);
nand U16430 (N_16430,N_15056,N_15678);
nand U16431 (N_16431,N_15759,N_15280);
and U16432 (N_16432,N_15701,N_15774);
xor U16433 (N_16433,N_15223,N_15933);
nor U16434 (N_16434,N_15140,N_15277);
nor U16435 (N_16435,N_15392,N_15866);
nand U16436 (N_16436,N_15735,N_15516);
and U16437 (N_16437,N_15210,N_15097);
or U16438 (N_16438,N_15868,N_15874);
xnor U16439 (N_16439,N_15218,N_15026);
and U16440 (N_16440,N_15927,N_15613);
or U16441 (N_16441,N_15105,N_15557);
xor U16442 (N_16442,N_15110,N_15373);
nand U16443 (N_16443,N_15236,N_15113);
nor U16444 (N_16444,N_15219,N_15978);
and U16445 (N_16445,N_15811,N_15079);
nor U16446 (N_16446,N_15308,N_15752);
nor U16447 (N_16447,N_15928,N_15602);
nor U16448 (N_16448,N_15737,N_15659);
xnor U16449 (N_16449,N_15246,N_15513);
or U16450 (N_16450,N_15375,N_15741);
and U16451 (N_16451,N_15627,N_15738);
nand U16452 (N_16452,N_15756,N_15250);
and U16453 (N_16453,N_15619,N_15369);
and U16454 (N_16454,N_15149,N_15935);
and U16455 (N_16455,N_15817,N_15747);
xor U16456 (N_16456,N_15593,N_15394);
or U16457 (N_16457,N_15476,N_15711);
and U16458 (N_16458,N_15917,N_15098);
or U16459 (N_16459,N_15036,N_15293);
xor U16460 (N_16460,N_15068,N_15698);
nand U16461 (N_16461,N_15632,N_15111);
nand U16462 (N_16462,N_15472,N_15570);
nor U16463 (N_16463,N_15395,N_15311);
and U16464 (N_16464,N_15545,N_15841);
nand U16465 (N_16465,N_15812,N_15947);
xnor U16466 (N_16466,N_15185,N_15780);
and U16467 (N_16467,N_15976,N_15063);
nand U16468 (N_16468,N_15452,N_15958);
xnor U16469 (N_16469,N_15354,N_15279);
nand U16470 (N_16470,N_15962,N_15021);
and U16471 (N_16471,N_15496,N_15206);
nand U16472 (N_16472,N_15862,N_15719);
and U16473 (N_16473,N_15767,N_15119);
or U16474 (N_16474,N_15382,N_15930);
xor U16475 (N_16475,N_15566,N_15480);
xor U16476 (N_16476,N_15965,N_15518);
and U16477 (N_16477,N_15205,N_15482);
and U16478 (N_16478,N_15924,N_15384);
and U16479 (N_16479,N_15331,N_15376);
and U16480 (N_16480,N_15430,N_15971);
nand U16481 (N_16481,N_15599,N_15189);
nand U16482 (N_16482,N_15847,N_15270);
xnor U16483 (N_16483,N_15444,N_15327);
and U16484 (N_16484,N_15181,N_15169);
nor U16485 (N_16485,N_15087,N_15066);
xnor U16486 (N_16486,N_15624,N_15147);
nand U16487 (N_16487,N_15796,N_15174);
nor U16488 (N_16488,N_15470,N_15940);
and U16489 (N_16489,N_15906,N_15316);
and U16490 (N_16490,N_15285,N_15751);
or U16491 (N_16491,N_15763,N_15199);
nor U16492 (N_16492,N_15576,N_15688);
xor U16493 (N_16493,N_15676,N_15800);
xor U16494 (N_16494,N_15042,N_15044);
or U16495 (N_16495,N_15274,N_15860);
or U16496 (N_16496,N_15849,N_15348);
or U16497 (N_16497,N_15733,N_15515);
xnor U16498 (N_16498,N_15034,N_15946);
xnor U16499 (N_16499,N_15859,N_15642);
nor U16500 (N_16500,N_15098,N_15133);
nand U16501 (N_16501,N_15866,N_15960);
or U16502 (N_16502,N_15141,N_15812);
and U16503 (N_16503,N_15224,N_15495);
xor U16504 (N_16504,N_15509,N_15903);
and U16505 (N_16505,N_15320,N_15067);
nand U16506 (N_16506,N_15628,N_15686);
nand U16507 (N_16507,N_15658,N_15612);
and U16508 (N_16508,N_15425,N_15850);
or U16509 (N_16509,N_15130,N_15230);
or U16510 (N_16510,N_15573,N_15615);
and U16511 (N_16511,N_15950,N_15311);
and U16512 (N_16512,N_15447,N_15359);
or U16513 (N_16513,N_15113,N_15165);
or U16514 (N_16514,N_15836,N_15931);
and U16515 (N_16515,N_15043,N_15007);
xor U16516 (N_16516,N_15301,N_15139);
nor U16517 (N_16517,N_15177,N_15244);
xnor U16518 (N_16518,N_15150,N_15476);
or U16519 (N_16519,N_15778,N_15898);
or U16520 (N_16520,N_15551,N_15682);
or U16521 (N_16521,N_15235,N_15148);
xor U16522 (N_16522,N_15161,N_15502);
or U16523 (N_16523,N_15383,N_15806);
nand U16524 (N_16524,N_15476,N_15739);
xnor U16525 (N_16525,N_15193,N_15794);
or U16526 (N_16526,N_15955,N_15215);
or U16527 (N_16527,N_15449,N_15700);
or U16528 (N_16528,N_15531,N_15347);
nand U16529 (N_16529,N_15894,N_15950);
nor U16530 (N_16530,N_15889,N_15181);
nand U16531 (N_16531,N_15451,N_15321);
or U16532 (N_16532,N_15095,N_15778);
nand U16533 (N_16533,N_15324,N_15272);
nand U16534 (N_16534,N_15208,N_15490);
nand U16535 (N_16535,N_15180,N_15748);
and U16536 (N_16536,N_15909,N_15139);
nor U16537 (N_16537,N_15577,N_15167);
and U16538 (N_16538,N_15308,N_15192);
or U16539 (N_16539,N_15175,N_15253);
nor U16540 (N_16540,N_15319,N_15711);
and U16541 (N_16541,N_15556,N_15395);
nand U16542 (N_16542,N_15551,N_15011);
or U16543 (N_16543,N_15489,N_15893);
xnor U16544 (N_16544,N_15417,N_15238);
xnor U16545 (N_16545,N_15477,N_15757);
xnor U16546 (N_16546,N_15038,N_15342);
or U16547 (N_16547,N_15607,N_15821);
or U16548 (N_16548,N_15349,N_15617);
xor U16549 (N_16549,N_15438,N_15466);
or U16550 (N_16550,N_15944,N_15299);
nor U16551 (N_16551,N_15014,N_15246);
xor U16552 (N_16552,N_15924,N_15793);
and U16553 (N_16553,N_15222,N_15468);
and U16554 (N_16554,N_15644,N_15005);
or U16555 (N_16555,N_15800,N_15951);
or U16556 (N_16556,N_15144,N_15142);
nand U16557 (N_16557,N_15971,N_15752);
nor U16558 (N_16558,N_15402,N_15809);
xnor U16559 (N_16559,N_15113,N_15465);
xor U16560 (N_16560,N_15920,N_15250);
or U16561 (N_16561,N_15206,N_15859);
and U16562 (N_16562,N_15934,N_15760);
or U16563 (N_16563,N_15322,N_15839);
nor U16564 (N_16564,N_15835,N_15937);
nand U16565 (N_16565,N_15816,N_15173);
or U16566 (N_16566,N_15109,N_15442);
nand U16567 (N_16567,N_15063,N_15081);
or U16568 (N_16568,N_15226,N_15667);
nor U16569 (N_16569,N_15069,N_15422);
nand U16570 (N_16570,N_15346,N_15517);
and U16571 (N_16571,N_15075,N_15641);
and U16572 (N_16572,N_15495,N_15994);
nand U16573 (N_16573,N_15322,N_15695);
nand U16574 (N_16574,N_15250,N_15234);
or U16575 (N_16575,N_15797,N_15436);
nor U16576 (N_16576,N_15470,N_15082);
and U16577 (N_16577,N_15588,N_15830);
and U16578 (N_16578,N_15320,N_15980);
nor U16579 (N_16579,N_15182,N_15593);
and U16580 (N_16580,N_15353,N_15493);
nor U16581 (N_16581,N_15211,N_15405);
and U16582 (N_16582,N_15322,N_15031);
nand U16583 (N_16583,N_15811,N_15379);
nor U16584 (N_16584,N_15372,N_15272);
xor U16585 (N_16585,N_15381,N_15805);
or U16586 (N_16586,N_15869,N_15799);
or U16587 (N_16587,N_15120,N_15388);
nor U16588 (N_16588,N_15047,N_15495);
xor U16589 (N_16589,N_15079,N_15464);
and U16590 (N_16590,N_15627,N_15692);
xor U16591 (N_16591,N_15609,N_15825);
xor U16592 (N_16592,N_15789,N_15701);
or U16593 (N_16593,N_15175,N_15909);
or U16594 (N_16594,N_15544,N_15637);
xor U16595 (N_16595,N_15208,N_15069);
or U16596 (N_16596,N_15034,N_15360);
and U16597 (N_16597,N_15285,N_15194);
nor U16598 (N_16598,N_15743,N_15043);
nor U16599 (N_16599,N_15097,N_15972);
xnor U16600 (N_16600,N_15676,N_15227);
nand U16601 (N_16601,N_15024,N_15250);
or U16602 (N_16602,N_15938,N_15675);
and U16603 (N_16603,N_15542,N_15136);
or U16604 (N_16604,N_15369,N_15878);
xnor U16605 (N_16605,N_15291,N_15046);
or U16606 (N_16606,N_15203,N_15228);
and U16607 (N_16607,N_15896,N_15221);
xor U16608 (N_16608,N_15225,N_15206);
xnor U16609 (N_16609,N_15822,N_15110);
or U16610 (N_16610,N_15988,N_15334);
nor U16611 (N_16611,N_15640,N_15939);
nand U16612 (N_16612,N_15608,N_15213);
xnor U16613 (N_16613,N_15045,N_15231);
or U16614 (N_16614,N_15645,N_15786);
xor U16615 (N_16615,N_15509,N_15496);
nor U16616 (N_16616,N_15943,N_15729);
or U16617 (N_16617,N_15137,N_15787);
nor U16618 (N_16618,N_15526,N_15270);
nor U16619 (N_16619,N_15809,N_15927);
nand U16620 (N_16620,N_15177,N_15148);
nor U16621 (N_16621,N_15635,N_15746);
xnor U16622 (N_16622,N_15668,N_15490);
nand U16623 (N_16623,N_15893,N_15537);
nor U16624 (N_16624,N_15824,N_15057);
xnor U16625 (N_16625,N_15861,N_15763);
nand U16626 (N_16626,N_15860,N_15596);
nand U16627 (N_16627,N_15218,N_15543);
nor U16628 (N_16628,N_15606,N_15234);
and U16629 (N_16629,N_15175,N_15517);
nor U16630 (N_16630,N_15483,N_15392);
nand U16631 (N_16631,N_15937,N_15692);
xnor U16632 (N_16632,N_15981,N_15316);
xnor U16633 (N_16633,N_15794,N_15388);
nand U16634 (N_16634,N_15079,N_15933);
nor U16635 (N_16635,N_15925,N_15708);
xnor U16636 (N_16636,N_15548,N_15525);
nor U16637 (N_16637,N_15840,N_15376);
or U16638 (N_16638,N_15555,N_15240);
nand U16639 (N_16639,N_15249,N_15154);
xor U16640 (N_16640,N_15674,N_15808);
or U16641 (N_16641,N_15004,N_15733);
or U16642 (N_16642,N_15713,N_15628);
nand U16643 (N_16643,N_15804,N_15670);
nor U16644 (N_16644,N_15397,N_15169);
xor U16645 (N_16645,N_15341,N_15121);
xor U16646 (N_16646,N_15333,N_15965);
xor U16647 (N_16647,N_15722,N_15046);
nand U16648 (N_16648,N_15907,N_15324);
nand U16649 (N_16649,N_15281,N_15393);
and U16650 (N_16650,N_15185,N_15615);
nand U16651 (N_16651,N_15582,N_15731);
nor U16652 (N_16652,N_15841,N_15656);
or U16653 (N_16653,N_15726,N_15239);
nor U16654 (N_16654,N_15676,N_15805);
nand U16655 (N_16655,N_15936,N_15656);
nor U16656 (N_16656,N_15646,N_15088);
xnor U16657 (N_16657,N_15970,N_15252);
nand U16658 (N_16658,N_15261,N_15392);
nand U16659 (N_16659,N_15282,N_15818);
xor U16660 (N_16660,N_15729,N_15112);
or U16661 (N_16661,N_15129,N_15589);
or U16662 (N_16662,N_15175,N_15060);
xor U16663 (N_16663,N_15743,N_15837);
nor U16664 (N_16664,N_15456,N_15801);
or U16665 (N_16665,N_15316,N_15838);
or U16666 (N_16666,N_15657,N_15120);
nand U16667 (N_16667,N_15601,N_15980);
nand U16668 (N_16668,N_15424,N_15342);
nand U16669 (N_16669,N_15126,N_15513);
and U16670 (N_16670,N_15657,N_15692);
and U16671 (N_16671,N_15687,N_15923);
xnor U16672 (N_16672,N_15702,N_15793);
nor U16673 (N_16673,N_15092,N_15854);
or U16674 (N_16674,N_15391,N_15161);
xnor U16675 (N_16675,N_15198,N_15317);
or U16676 (N_16676,N_15766,N_15980);
xnor U16677 (N_16677,N_15468,N_15092);
or U16678 (N_16678,N_15528,N_15853);
nand U16679 (N_16679,N_15412,N_15644);
xnor U16680 (N_16680,N_15501,N_15385);
or U16681 (N_16681,N_15172,N_15889);
nand U16682 (N_16682,N_15321,N_15735);
nor U16683 (N_16683,N_15642,N_15094);
or U16684 (N_16684,N_15582,N_15785);
or U16685 (N_16685,N_15383,N_15337);
xor U16686 (N_16686,N_15330,N_15289);
and U16687 (N_16687,N_15875,N_15759);
xor U16688 (N_16688,N_15695,N_15398);
nand U16689 (N_16689,N_15258,N_15764);
xnor U16690 (N_16690,N_15807,N_15500);
nor U16691 (N_16691,N_15585,N_15463);
and U16692 (N_16692,N_15326,N_15780);
or U16693 (N_16693,N_15656,N_15577);
nor U16694 (N_16694,N_15745,N_15790);
and U16695 (N_16695,N_15250,N_15006);
or U16696 (N_16696,N_15194,N_15019);
nand U16697 (N_16697,N_15289,N_15822);
nand U16698 (N_16698,N_15327,N_15473);
xor U16699 (N_16699,N_15386,N_15625);
or U16700 (N_16700,N_15941,N_15500);
nand U16701 (N_16701,N_15393,N_15006);
and U16702 (N_16702,N_15016,N_15499);
and U16703 (N_16703,N_15711,N_15942);
nand U16704 (N_16704,N_15353,N_15338);
and U16705 (N_16705,N_15298,N_15880);
xor U16706 (N_16706,N_15463,N_15501);
nand U16707 (N_16707,N_15381,N_15859);
and U16708 (N_16708,N_15208,N_15659);
nand U16709 (N_16709,N_15205,N_15562);
xor U16710 (N_16710,N_15815,N_15701);
nor U16711 (N_16711,N_15542,N_15900);
nor U16712 (N_16712,N_15631,N_15743);
and U16713 (N_16713,N_15501,N_15373);
xor U16714 (N_16714,N_15693,N_15026);
nand U16715 (N_16715,N_15326,N_15914);
nand U16716 (N_16716,N_15552,N_15106);
xor U16717 (N_16717,N_15704,N_15883);
nand U16718 (N_16718,N_15992,N_15420);
nor U16719 (N_16719,N_15046,N_15501);
nand U16720 (N_16720,N_15605,N_15461);
and U16721 (N_16721,N_15406,N_15856);
or U16722 (N_16722,N_15338,N_15870);
or U16723 (N_16723,N_15105,N_15248);
and U16724 (N_16724,N_15370,N_15571);
xnor U16725 (N_16725,N_15041,N_15645);
or U16726 (N_16726,N_15333,N_15824);
and U16727 (N_16727,N_15781,N_15074);
and U16728 (N_16728,N_15672,N_15716);
or U16729 (N_16729,N_15099,N_15657);
nor U16730 (N_16730,N_15655,N_15251);
or U16731 (N_16731,N_15103,N_15083);
xnor U16732 (N_16732,N_15254,N_15015);
xnor U16733 (N_16733,N_15490,N_15686);
and U16734 (N_16734,N_15944,N_15372);
xor U16735 (N_16735,N_15900,N_15331);
nand U16736 (N_16736,N_15023,N_15615);
and U16737 (N_16737,N_15987,N_15297);
nor U16738 (N_16738,N_15547,N_15055);
nor U16739 (N_16739,N_15275,N_15515);
nor U16740 (N_16740,N_15115,N_15239);
nor U16741 (N_16741,N_15534,N_15277);
xnor U16742 (N_16742,N_15079,N_15785);
or U16743 (N_16743,N_15479,N_15510);
nand U16744 (N_16744,N_15670,N_15387);
xnor U16745 (N_16745,N_15466,N_15659);
xor U16746 (N_16746,N_15599,N_15125);
and U16747 (N_16747,N_15707,N_15178);
or U16748 (N_16748,N_15314,N_15438);
nand U16749 (N_16749,N_15303,N_15163);
and U16750 (N_16750,N_15169,N_15029);
or U16751 (N_16751,N_15179,N_15941);
and U16752 (N_16752,N_15869,N_15321);
xor U16753 (N_16753,N_15783,N_15841);
xnor U16754 (N_16754,N_15284,N_15805);
and U16755 (N_16755,N_15338,N_15078);
nand U16756 (N_16756,N_15608,N_15554);
or U16757 (N_16757,N_15999,N_15027);
and U16758 (N_16758,N_15902,N_15258);
nor U16759 (N_16759,N_15812,N_15356);
nand U16760 (N_16760,N_15578,N_15385);
xnor U16761 (N_16761,N_15518,N_15230);
nand U16762 (N_16762,N_15560,N_15268);
xor U16763 (N_16763,N_15428,N_15414);
or U16764 (N_16764,N_15963,N_15283);
xnor U16765 (N_16765,N_15208,N_15782);
xnor U16766 (N_16766,N_15141,N_15119);
xnor U16767 (N_16767,N_15496,N_15918);
or U16768 (N_16768,N_15644,N_15749);
nand U16769 (N_16769,N_15600,N_15511);
and U16770 (N_16770,N_15458,N_15572);
nand U16771 (N_16771,N_15545,N_15509);
nand U16772 (N_16772,N_15030,N_15759);
or U16773 (N_16773,N_15823,N_15324);
and U16774 (N_16774,N_15095,N_15677);
nor U16775 (N_16775,N_15553,N_15292);
xnor U16776 (N_16776,N_15443,N_15015);
nand U16777 (N_16777,N_15236,N_15341);
xor U16778 (N_16778,N_15144,N_15770);
nor U16779 (N_16779,N_15466,N_15980);
nor U16780 (N_16780,N_15467,N_15105);
and U16781 (N_16781,N_15250,N_15907);
xor U16782 (N_16782,N_15247,N_15092);
xnor U16783 (N_16783,N_15698,N_15997);
nor U16784 (N_16784,N_15503,N_15790);
or U16785 (N_16785,N_15369,N_15777);
nand U16786 (N_16786,N_15023,N_15229);
xnor U16787 (N_16787,N_15149,N_15991);
xor U16788 (N_16788,N_15507,N_15500);
nor U16789 (N_16789,N_15269,N_15090);
nand U16790 (N_16790,N_15660,N_15308);
or U16791 (N_16791,N_15707,N_15177);
xnor U16792 (N_16792,N_15941,N_15327);
nor U16793 (N_16793,N_15771,N_15088);
or U16794 (N_16794,N_15223,N_15620);
and U16795 (N_16795,N_15506,N_15048);
or U16796 (N_16796,N_15577,N_15055);
nor U16797 (N_16797,N_15632,N_15479);
nor U16798 (N_16798,N_15688,N_15254);
nor U16799 (N_16799,N_15080,N_15543);
nand U16800 (N_16800,N_15149,N_15114);
or U16801 (N_16801,N_15907,N_15177);
nand U16802 (N_16802,N_15200,N_15895);
nand U16803 (N_16803,N_15418,N_15443);
nor U16804 (N_16804,N_15324,N_15680);
or U16805 (N_16805,N_15333,N_15947);
xnor U16806 (N_16806,N_15590,N_15864);
nand U16807 (N_16807,N_15322,N_15344);
xor U16808 (N_16808,N_15560,N_15951);
xor U16809 (N_16809,N_15679,N_15376);
and U16810 (N_16810,N_15715,N_15664);
nand U16811 (N_16811,N_15798,N_15274);
or U16812 (N_16812,N_15984,N_15653);
or U16813 (N_16813,N_15334,N_15101);
xor U16814 (N_16814,N_15356,N_15906);
nor U16815 (N_16815,N_15648,N_15488);
xor U16816 (N_16816,N_15011,N_15260);
or U16817 (N_16817,N_15662,N_15236);
xor U16818 (N_16818,N_15824,N_15619);
nor U16819 (N_16819,N_15470,N_15182);
xor U16820 (N_16820,N_15685,N_15959);
nor U16821 (N_16821,N_15659,N_15657);
and U16822 (N_16822,N_15623,N_15299);
and U16823 (N_16823,N_15852,N_15229);
nor U16824 (N_16824,N_15708,N_15453);
and U16825 (N_16825,N_15471,N_15540);
or U16826 (N_16826,N_15738,N_15366);
nor U16827 (N_16827,N_15716,N_15617);
nor U16828 (N_16828,N_15730,N_15756);
and U16829 (N_16829,N_15473,N_15698);
nor U16830 (N_16830,N_15688,N_15335);
nand U16831 (N_16831,N_15410,N_15947);
xnor U16832 (N_16832,N_15620,N_15422);
and U16833 (N_16833,N_15136,N_15528);
or U16834 (N_16834,N_15255,N_15952);
or U16835 (N_16835,N_15345,N_15440);
or U16836 (N_16836,N_15876,N_15284);
xor U16837 (N_16837,N_15684,N_15905);
or U16838 (N_16838,N_15606,N_15863);
nand U16839 (N_16839,N_15331,N_15162);
xnor U16840 (N_16840,N_15861,N_15335);
xor U16841 (N_16841,N_15115,N_15842);
nand U16842 (N_16842,N_15731,N_15829);
or U16843 (N_16843,N_15790,N_15926);
nand U16844 (N_16844,N_15351,N_15299);
nand U16845 (N_16845,N_15531,N_15199);
or U16846 (N_16846,N_15252,N_15740);
or U16847 (N_16847,N_15214,N_15931);
and U16848 (N_16848,N_15818,N_15001);
xor U16849 (N_16849,N_15782,N_15050);
or U16850 (N_16850,N_15822,N_15713);
xnor U16851 (N_16851,N_15049,N_15168);
or U16852 (N_16852,N_15067,N_15494);
xnor U16853 (N_16853,N_15235,N_15584);
nor U16854 (N_16854,N_15844,N_15105);
xnor U16855 (N_16855,N_15827,N_15867);
xnor U16856 (N_16856,N_15139,N_15601);
and U16857 (N_16857,N_15954,N_15265);
nor U16858 (N_16858,N_15044,N_15220);
xor U16859 (N_16859,N_15947,N_15534);
xnor U16860 (N_16860,N_15899,N_15051);
nor U16861 (N_16861,N_15005,N_15333);
nand U16862 (N_16862,N_15837,N_15744);
and U16863 (N_16863,N_15278,N_15101);
nand U16864 (N_16864,N_15882,N_15929);
nor U16865 (N_16865,N_15475,N_15834);
or U16866 (N_16866,N_15945,N_15224);
nor U16867 (N_16867,N_15874,N_15475);
nand U16868 (N_16868,N_15603,N_15093);
and U16869 (N_16869,N_15418,N_15203);
nand U16870 (N_16870,N_15476,N_15664);
or U16871 (N_16871,N_15364,N_15794);
nor U16872 (N_16872,N_15694,N_15557);
or U16873 (N_16873,N_15726,N_15121);
xnor U16874 (N_16874,N_15232,N_15725);
or U16875 (N_16875,N_15559,N_15892);
xnor U16876 (N_16876,N_15911,N_15388);
and U16877 (N_16877,N_15805,N_15232);
or U16878 (N_16878,N_15286,N_15152);
nand U16879 (N_16879,N_15599,N_15555);
xnor U16880 (N_16880,N_15451,N_15477);
xnor U16881 (N_16881,N_15629,N_15468);
nand U16882 (N_16882,N_15675,N_15094);
xnor U16883 (N_16883,N_15262,N_15503);
or U16884 (N_16884,N_15043,N_15702);
xnor U16885 (N_16885,N_15837,N_15512);
and U16886 (N_16886,N_15792,N_15737);
nor U16887 (N_16887,N_15910,N_15631);
xor U16888 (N_16888,N_15194,N_15071);
xor U16889 (N_16889,N_15051,N_15882);
or U16890 (N_16890,N_15273,N_15448);
and U16891 (N_16891,N_15899,N_15790);
nor U16892 (N_16892,N_15320,N_15448);
xnor U16893 (N_16893,N_15158,N_15214);
xor U16894 (N_16894,N_15198,N_15359);
and U16895 (N_16895,N_15851,N_15649);
nor U16896 (N_16896,N_15059,N_15024);
nor U16897 (N_16897,N_15282,N_15971);
and U16898 (N_16898,N_15658,N_15802);
xnor U16899 (N_16899,N_15658,N_15256);
and U16900 (N_16900,N_15288,N_15512);
nand U16901 (N_16901,N_15689,N_15699);
or U16902 (N_16902,N_15472,N_15856);
and U16903 (N_16903,N_15659,N_15993);
xor U16904 (N_16904,N_15906,N_15749);
nor U16905 (N_16905,N_15618,N_15135);
or U16906 (N_16906,N_15416,N_15023);
nand U16907 (N_16907,N_15174,N_15618);
and U16908 (N_16908,N_15976,N_15121);
nand U16909 (N_16909,N_15847,N_15900);
or U16910 (N_16910,N_15183,N_15958);
nand U16911 (N_16911,N_15843,N_15986);
and U16912 (N_16912,N_15892,N_15560);
and U16913 (N_16913,N_15402,N_15167);
or U16914 (N_16914,N_15666,N_15845);
nand U16915 (N_16915,N_15440,N_15168);
nor U16916 (N_16916,N_15222,N_15863);
xnor U16917 (N_16917,N_15579,N_15595);
and U16918 (N_16918,N_15929,N_15767);
and U16919 (N_16919,N_15220,N_15734);
and U16920 (N_16920,N_15691,N_15357);
nand U16921 (N_16921,N_15357,N_15540);
nor U16922 (N_16922,N_15594,N_15498);
and U16923 (N_16923,N_15160,N_15320);
or U16924 (N_16924,N_15274,N_15774);
nand U16925 (N_16925,N_15405,N_15063);
nand U16926 (N_16926,N_15654,N_15278);
or U16927 (N_16927,N_15658,N_15039);
nor U16928 (N_16928,N_15263,N_15522);
and U16929 (N_16929,N_15789,N_15181);
nand U16930 (N_16930,N_15020,N_15285);
or U16931 (N_16931,N_15446,N_15860);
or U16932 (N_16932,N_15949,N_15897);
and U16933 (N_16933,N_15461,N_15260);
or U16934 (N_16934,N_15319,N_15325);
xor U16935 (N_16935,N_15208,N_15128);
nand U16936 (N_16936,N_15923,N_15524);
xnor U16937 (N_16937,N_15542,N_15943);
xor U16938 (N_16938,N_15123,N_15041);
and U16939 (N_16939,N_15246,N_15448);
nor U16940 (N_16940,N_15831,N_15421);
nand U16941 (N_16941,N_15916,N_15667);
nand U16942 (N_16942,N_15347,N_15957);
or U16943 (N_16943,N_15496,N_15992);
or U16944 (N_16944,N_15742,N_15133);
or U16945 (N_16945,N_15131,N_15237);
or U16946 (N_16946,N_15438,N_15656);
xor U16947 (N_16947,N_15574,N_15506);
xor U16948 (N_16948,N_15716,N_15819);
nor U16949 (N_16949,N_15788,N_15300);
or U16950 (N_16950,N_15770,N_15923);
and U16951 (N_16951,N_15659,N_15717);
or U16952 (N_16952,N_15312,N_15497);
nand U16953 (N_16953,N_15684,N_15593);
or U16954 (N_16954,N_15020,N_15931);
nand U16955 (N_16955,N_15204,N_15123);
nand U16956 (N_16956,N_15662,N_15807);
and U16957 (N_16957,N_15744,N_15902);
nor U16958 (N_16958,N_15016,N_15964);
and U16959 (N_16959,N_15416,N_15396);
xor U16960 (N_16960,N_15669,N_15767);
and U16961 (N_16961,N_15376,N_15999);
nand U16962 (N_16962,N_15605,N_15500);
and U16963 (N_16963,N_15289,N_15095);
or U16964 (N_16964,N_15049,N_15830);
xnor U16965 (N_16965,N_15748,N_15558);
xor U16966 (N_16966,N_15192,N_15144);
xor U16967 (N_16967,N_15278,N_15094);
and U16968 (N_16968,N_15366,N_15519);
xnor U16969 (N_16969,N_15414,N_15961);
nand U16970 (N_16970,N_15722,N_15223);
and U16971 (N_16971,N_15617,N_15873);
nor U16972 (N_16972,N_15816,N_15944);
or U16973 (N_16973,N_15883,N_15051);
xor U16974 (N_16974,N_15461,N_15896);
or U16975 (N_16975,N_15495,N_15296);
nor U16976 (N_16976,N_15964,N_15694);
and U16977 (N_16977,N_15759,N_15913);
nand U16978 (N_16978,N_15988,N_15586);
and U16979 (N_16979,N_15202,N_15522);
xnor U16980 (N_16980,N_15243,N_15218);
or U16981 (N_16981,N_15597,N_15820);
xnor U16982 (N_16982,N_15375,N_15009);
xnor U16983 (N_16983,N_15576,N_15484);
and U16984 (N_16984,N_15616,N_15672);
nor U16985 (N_16985,N_15384,N_15874);
and U16986 (N_16986,N_15083,N_15261);
xnor U16987 (N_16987,N_15068,N_15416);
nor U16988 (N_16988,N_15455,N_15284);
or U16989 (N_16989,N_15883,N_15824);
nand U16990 (N_16990,N_15304,N_15002);
and U16991 (N_16991,N_15737,N_15225);
nor U16992 (N_16992,N_15703,N_15251);
nor U16993 (N_16993,N_15880,N_15973);
nor U16994 (N_16994,N_15854,N_15883);
nor U16995 (N_16995,N_15341,N_15415);
nand U16996 (N_16996,N_15255,N_15814);
nor U16997 (N_16997,N_15904,N_15800);
nand U16998 (N_16998,N_15109,N_15649);
nand U16999 (N_16999,N_15683,N_15532);
and U17000 (N_17000,N_16932,N_16136);
or U17001 (N_17001,N_16059,N_16393);
or U17002 (N_17002,N_16614,N_16230);
nor U17003 (N_17003,N_16904,N_16713);
xor U17004 (N_17004,N_16867,N_16953);
or U17005 (N_17005,N_16769,N_16518);
nand U17006 (N_17006,N_16607,N_16359);
or U17007 (N_17007,N_16716,N_16263);
and U17008 (N_17008,N_16666,N_16862);
xnor U17009 (N_17009,N_16679,N_16421);
nor U17010 (N_17010,N_16451,N_16299);
or U17011 (N_17011,N_16731,N_16377);
nand U17012 (N_17012,N_16815,N_16826);
xor U17013 (N_17013,N_16523,N_16423);
or U17014 (N_17014,N_16215,N_16336);
and U17015 (N_17015,N_16751,N_16290);
xnor U17016 (N_17016,N_16705,N_16467);
or U17017 (N_17017,N_16793,N_16834);
and U17018 (N_17018,N_16908,N_16387);
nand U17019 (N_17019,N_16099,N_16554);
nand U17020 (N_17020,N_16999,N_16756);
nor U17021 (N_17021,N_16732,N_16311);
nand U17022 (N_17022,N_16181,N_16695);
and U17023 (N_17023,N_16086,N_16573);
nand U17024 (N_17024,N_16665,N_16762);
nand U17025 (N_17025,N_16042,N_16191);
nor U17026 (N_17026,N_16422,N_16744);
nor U17027 (N_17027,N_16753,N_16588);
or U17028 (N_17028,N_16582,N_16894);
nand U17029 (N_17029,N_16839,N_16209);
or U17030 (N_17030,N_16205,N_16077);
nor U17031 (N_17031,N_16802,N_16707);
nand U17032 (N_17032,N_16322,N_16273);
and U17033 (N_17033,N_16124,N_16015);
nand U17034 (N_17034,N_16537,N_16982);
or U17035 (N_17035,N_16658,N_16696);
nor U17036 (N_17036,N_16197,N_16417);
and U17037 (N_17037,N_16628,N_16211);
or U17038 (N_17038,N_16176,N_16613);
and U17039 (N_17039,N_16175,N_16975);
nand U17040 (N_17040,N_16725,N_16631);
nand U17041 (N_17041,N_16689,N_16328);
or U17042 (N_17042,N_16061,N_16901);
nor U17043 (N_17043,N_16801,N_16062);
xnor U17044 (N_17044,N_16830,N_16533);
and U17045 (N_17045,N_16313,N_16693);
nand U17046 (N_17046,N_16357,N_16065);
and U17047 (N_17047,N_16361,N_16105);
or U17048 (N_17048,N_16638,N_16045);
nor U17049 (N_17049,N_16775,N_16318);
or U17050 (N_17050,N_16850,N_16781);
or U17051 (N_17051,N_16216,N_16097);
xnor U17052 (N_17052,N_16228,N_16545);
or U17053 (N_17053,N_16761,N_16231);
nand U17054 (N_17054,N_16708,N_16212);
xor U17055 (N_17055,N_16568,N_16429);
nand U17056 (N_17056,N_16122,N_16486);
xnor U17057 (N_17057,N_16066,N_16021);
or U17058 (N_17058,N_16164,N_16046);
nor U17059 (N_17059,N_16390,N_16369);
xor U17060 (N_17060,N_16297,N_16427);
and U17061 (N_17061,N_16902,N_16684);
nand U17062 (N_17062,N_16567,N_16748);
nand U17063 (N_17063,N_16505,N_16360);
nor U17064 (N_17064,N_16782,N_16170);
or U17065 (N_17065,N_16399,N_16965);
xnor U17066 (N_17066,N_16171,N_16247);
nor U17067 (N_17067,N_16749,N_16504);
nand U17068 (N_17068,N_16434,N_16818);
xor U17069 (N_17069,N_16629,N_16340);
nand U17070 (N_17070,N_16321,N_16489);
xor U17071 (N_17071,N_16715,N_16188);
nand U17072 (N_17072,N_16616,N_16411);
nand U17073 (N_17073,N_16030,N_16962);
nand U17074 (N_17074,N_16510,N_16825);
xor U17075 (N_17075,N_16788,N_16052);
or U17076 (N_17076,N_16553,N_16719);
nor U17077 (N_17077,N_16722,N_16883);
or U17078 (N_17078,N_16098,N_16544);
nor U17079 (N_17079,N_16245,N_16827);
nand U17080 (N_17080,N_16298,N_16797);
xor U17081 (N_17081,N_16271,N_16840);
and U17082 (N_17082,N_16226,N_16376);
xnor U17083 (N_17083,N_16539,N_16010);
nor U17084 (N_17084,N_16771,N_16139);
or U17085 (N_17085,N_16773,N_16893);
or U17086 (N_17086,N_16661,N_16535);
xor U17087 (N_17087,N_16796,N_16326);
nand U17088 (N_17088,N_16534,N_16577);
nor U17089 (N_17089,N_16630,N_16286);
nand U17090 (N_17090,N_16499,N_16846);
nand U17091 (N_17091,N_16724,N_16559);
or U17092 (N_17092,N_16528,N_16746);
xor U17093 (N_17093,N_16625,N_16940);
nor U17094 (N_17094,N_16084,N_16005);
nand U17095 (N_17095,N_16853,N_16453);
nor U17096 (N_17096,N_16847,N_16512);
xor U17097 (N_17097,N_16088,N_16640);
xor U17098 (N_17098,N_16955,N_16865);
nand U17099 (N_17099,N_16547,N_16706);
nor U17100 (N_17100,N_16881,N_16593);
and U17101 (N_17101,N_16020,N_16141);
nor U17102 (N_17102,N_16174,N_16668);
or U17103 (N_17103,N_16524,N_16208);
and U17104 (N_17104,N_16758,N_16153);
and U17105 (N_17105,N_16096,N_16248);
and U17106 (N_17106,N_16019,N_16312);
or U17107 (N_17107,N_16754,N_16498);
or U17108 (N_17108,N_16458,N_16239);
nand U17109 (N_17109,N_16293,N_16024);
or U17110 (N_17110,N_16092,N_16119);
and U17111 (N_17111,N_16283,N_16919);
and U17112 (N_17112,N_16161,N_16323);
or U17113 (N_17113,N_16605,N_16770);
nor U17114 (N_17114,N_16222,N_16718);
nor U17115 (N_17115,N_16995,N_16849);
and U17116 (N_17116,N_16664,N_16246);
xnor U17117 (N_17117,N_16506,N_16575);
or U17118 (N_17118,N_16536,N_16876);
and U17119 (N_17119,N_16712,N_16039);
and U17120 (N_17120,N_16911,N_16514);
nand U17121 (N_17121,N_16483,N_16494);
nand U17122 (N_17122,N_16241,N_16670);
nand U17123 (N_17123,N_16845,N_16626);
nor U17124 (N_17124,N_16115,N_16728);
or U17125 (N_17125,N_16768,N_16617);
xor U17126 (N_17126,N_16651,N_16282);
nor U17127 (N_17127,N_16385,N_16492);
and U17128 (N_17128,N_16193,N_16497);
xnor U17129 (N_17129,N_16841,N_16765);
xnor U17130 (N_17130,N_16063,N_16159);
and U17131 (N_17131,N_16150,N_16319);
nand U17132 (N_17132,N_16950,N_16674);
nand U17133 (N_17133,N_16366,N_16147);
or U17134 (N_17134,N_16831,N_16898);
or U17135 (N_17135,N_16623,N_16268);
xor U17136 (N_17136,N_16990,N_16420);
and U17137 (N_17137,N_16527,N_16978);
xor U17138 (N_17138,N_16168,N_16333);
nand U17139 (N_17139,N_16866,N_16406);
or U17140 (N_17140,N_16743,N_16291);
xnor U17141 (N_17141,N_16274,N_16048);
nor U17142 (N_17142,N_16714,N_16407);
xor U17143 (N_17143,N_16662,N_16763);
xnor U17144 (N_17144,N_16659,N_16493);
nor U17145 (N_17145,N_16267,N_16158);
and U17146 (N_17146,N_16060,N_16799);
or U17147 (N_17147,N_16214,N_16936);
nand U17148 (N_17148,N_16229,N_16704);
xnor U17149 (N_17149,N_16075,N_16073);
nand U17150 (N_17150,N_16634,N_16103);
and U17151 (N_17151,N_16516,N_16221);
or U17152 (N_17152,N_16008,N_16766);
xor U17153 (N_17153,N_16424,N_16178);
xor U17154 (N_17154,N_16252,N_16832);
nand U17155 (N_17155,N_16302,N_16167);
xor U17156 (N_17156,N_16249,N_16350);
or U17157 (N_17157,N_16857,N_16145);
xnor U17158 (N_17158,N_16317,N_16113);
and U17159 (N_17159,N_16757,N_16811);
and U17160 (N_17160,N_16445,N_16315);
xor U17161 (N_17161,N_16121,N_16984);
and U17162 (N_17162,N_16805,N_16808);
or U17163 (N_17163,N_16438,N_16899);
xor U17164 (N_17164,N_16471,N_16993);
nor U17165 (N_17165,N_16220,N_16963);
or U17166 (N_17166,N_16179,N_16924);
nand U17167 (N_17167,N_16058,N_16259);
nor U17168 (N_17168,N_16070,N_16927);
and U17169 (N_17169,N_16806,N_16152);
nor U17170 (N_17170,N_16278,N_16495);
and U17171 (N_17171,N_16690,N_16325);
xor U17172 (N_17172,N_16777,N_16403);
xor U17173 (N_17173,N_16683,N_16117);
xnor U17174 (N_17174,N_16412,N_16233);
nor U17175 (N_17175,N_16597,N_16076);
and U17176 (N_17176,N_16198,N_16740);
nand U17177 (N_17177,N_16977,N_16384);
and U17178 (N_17178,N_16525,N_16300);
nor U17179 (N_17179,N_16223,N_16087);
nor U17180 (N_17180,N_16346,N_16882);
and U17181 (N_17181,N_16352,N_16371);
xnor U17182 (N_17182,N_16444,N_16501);
or U17183 (N_17183,N_16314,N_16676);
and U17184 (N_17184,N_16907,N_16921);
or U17185 (N_17185,N_16697,N_16373);
or U17186 (N_17186,N_16870,N_16143);
nor U17187 (N_17187,N_16917,N_16730);
nand U17188 (N_17188,N_16602,N_16860);
or U17189 (N_17189,N_16966,N_16054);
xnor U17190 (N_17190,N_16354,N_16204);
and U17191 (N_17191,N_16381,N_16854);
nand U17192 (N_17192,N_16723,N_16603);
xnor U17193 (N_17193,N_16726,N_16289);
or U17194 (N_17194,N_16186,N_16093);
or U17195 (N_17195,N_16800,N_16388);
nor U17196 (N_17196,N_16935,N_16426);
nand U17197 (N_17197,N_16165,N_16006);
nor U17198 (N_17198,N_16303,N_16433);
xor U17199 (N_17199,N_16102,N_16736);
and U17200 (N_17200,N_16824,N_16491);
or U17201 (N_17201,N_16686,N_16435);
nor U17202 (N_17202,N_16851,N_16108);
nand U17203 (N_17203,N_16116,N_16192);
xor U17204 (N_17204,N_16415,N_16945);
xor U17205 (N_17205,N_16878,N_16584);
and U17206 (N_17206,N_16244,N_16969);
or U17207 (N_17207,N_16028,N_16219);
or U17208 (N_17208,N_16050,N_16379);
and U17209 (N_17209,N_16069,N_16237);
nor U17210 (N_17210,N_16146,N_16017);
xor U17211 (N_17211,N_16803,N_16540);
nand U17212 (N_17212,N_16639,N_16998);
and U17213 (N_17213,N_16563,N_16861);
and U17214 (N_17214,N_16589,N_16368);
xnor U17215 (N_17215,N_16138,N_16473);
xor U17216 (N_17216,N_16864,N_16657);
and U17217 (N_17217,N_16155,N_16632);
or U17218 (N_17218,N_16700,N_16428);
and U17219 (N_17219,N_16583,N_16624);
and U17220 (N_17220,N_16701,N_16997);
or U17221 (N_17221,N_16913,N_16745);
nand U17222 (N_17222,N_16305,N_16968);
nor U17223 (N_17223,N_16942,N_16081);
xor U17224 (N_17224,N_16787,N_16372);
nand U17225 (N_17225,N_16600,N_16018);
nor U17226 (N_17226,N_16261,N_16419);
nand U17227 (N_17227,N_16660,N_16462);
xnor U17228 (N_17228,N_16272,N_16142);
nor U17229 (N_17229,N_16418,N_16546);
or U17230 (N_17230,N_16673,N_16238);
xor U17231 (N_17231,N_16580,N_16441);
nor U17232 (N_17232,N_16025,N_16067);
and U17233 (N_17233,N_16364,N_16110);
nor U17234 (N_17234,N_16530,N_16646);
nand U17235 (N_17235,N_16111,N_16329);
xor U17236 (N_17236,N_16177,N_16100);
nor U17237 (N_17237,N_16790,N_16585);
or U17238 (N_17238,N_16083,N_16079);
xnor U17239 (N_17239,N_16739,N_16031);
nand U17240 (N_17240,N_16408,N_16842);
or U17241 (N_17241,N_16256,N_16255);
nand U17242 (N_17242,N_16389,N_16721);
xor U17243 (N_17243,N_16644,N_16780);
nor U17244 (N_17244,N_16710,N_16513);
nor U17245 (N_17245,N_16040,N_16874);
or U17246 (N_17246,N_16078,N_16737);
xor U17247 (N_17247,N_16443,N_16468);
and U17248 (N_17248,N_16502,N_16447);
nor U17249 (N_17249,N_16033,N_16351);
and U17250 (N_17250,N_16785,N_16488);
and U17251 (N_17251,N_16571,N_16759);
or U17252 (N_17252,N_16621,N_16341);
nor U17253 (N_17253,N_16541,N_16203);
xnor U17254 (N_17254,N_16812,N_16948);
and U17255 (N_17255,N_16064,N_16413);
nor U17256 (N_17256,N_16049,N_16859);
nand U17257 (N_17257,N_16285,N_16500);
xor U17258 (N_17258,N_16980,N_16206);
xnor U17259 (N_17259,N_16126,N_16635);
nand U17260 (N_17260,N_16596,N_16843);
nor U17261 (N_17261,N_16038,N_16292);
and U17262 (N_17262,N_16735,N_16118);
nand U17263 (N_17263,N_16051,N_16671);
and U17264 (N_17264,N_16410,N_16699);
and U17265 (N_17265,N_16128,N_16449);
nor U17266 (N_17266,N_16946,N_16560);
nand U17267 (N_17267,N_16234,N_16154);
or U17268 (N_17268,N_16041,N_16558);
xor U17269 (N_17269,N_16933,N_16988);
and U17270 (N_17270,N_16717,N_16307);
nand U17271 (N_17271,N_16356,N_16809);
xnor U17272 (N_17272,N_16983,N_16264);
or U17273 (N_17273,N_16002,N_16074);
xor U17274 (N_17274,N_16798,N_16452);
xnor U17275 (N_17275,N_16729,N_16938);
nor U17276 (N_17276,N_16856,N_16095);
and U17277 (N_17277,N_16464,N_16822);
or U17278 (N_17278,N_16401,N_16649);
or U17279 (N_17279,N_16184,N_16457);
or U17280 (N_17280,N_16565,N_16681);
and U17281 (N_17281,N_16912,N_16875);
xnor U17282 (N_17282,N_16133,N_16833);
nand U17283 (N_17283,N_16162,N_16416);
and U17284 (N_17284,N_16375,N_16543);
and U17285 (N_17285,N_16370,N_16331);
xor U17286 (N_17286,N_16561,N_16251);
nor U17287 (N_17287,N_16578,N_16232);
nor U17288 (N_17288,N_16555,N_16182);
or U17289 (N_17289,N_16643,N_16531);
nand U17290 (N_17290,N_16804,N_16581);
nand U17291 (N_17291,N_16572,N_16956);
xor U17292 (N_17292,N_16470,N_16606);
and U17293 (N_17293,N_16398,N_16755);
xor U17294 (N_17294,N_16014,N_16277);
nand U17295 (N_17295,N_16210,N_16709);
xor U17296 (N_17296,N_16916,N_16240);
and U17297 (N_17297,N_16217,N_16873);
and U17298 (N_17298,N_16994,N_16342);
and U17299 (N_17299,N_16374,N_16144);
and U17300 (N_17300,N_16973,N_16194);
xnor U17301 (N_17301,N_16478,N_16301);
or U17302 (N_17302,N_16125,N_16521);
xnor U17303 (N_17303,N_16654,N_16227);
nand U17304 (N_17304,N_16253,N_16642);
or U17305 (N_17305,N_16914,N_16837);
or U17306 (N_17306,N_16094,N_16480);
or U17307 (N_17307,N_16574,N_16542);
nor U17308 (N_17308,N_16280,N_16918);
nor U17309 (N_17309,N_16767,N_16947);
and U17310 (N_17310,N_16915,N_16810);
nor U17311 (N_17311,N_16877,N_16734);
nand U17312 (N_17312,N_16466,N_16905);
nand U17313 (N_17313,N_16669,N_16934);
nor U17314 (N_17314,N_16667,N_16258);
nand U17315 (N_17315,N_16482,N_16974);
and U17316 (N_17316,N_16814,N_16254);
or U17317 (N_17317,N_16627,N_16207);
nor U17318 (N_17318,N_16347,N_16633);
nor U17319 (N_17319,N_16131,N_16134);
or U17320 (N_17320,N_16169,N_16149);
or U17321 (N_17321,N_16257,N_16243);
xor U17322 (N_17322,N_16475,N_16446);
or U17323 (N_17323,N_16455,N_16636);
nor U17324 (N_17324,N_16053,N_16454);
nor U17325 (N_17325,N_16871,N_16711);
xor U17326 (N_17326,N_16106,N_16309);
and U17327 (N_17327,N_16620,N_16476);
nor U17328 (N_17328,N_16027,N_16242);
and U17329 (N_17329,N_16450,N_16348);
xor U17330 (N_17330,N_16836,N_16549);
xor U17331 (N_17331,N_16479,N_16703);
and U17332 (N_17332,N_16764,N_16202);
or U17333 (N_17333,N_16355,N_16647);
xor U17334 (N_17334,N_16784,N_16090);
nor U17335 (N_17335,N_16880,N_16199);
nand U17336 (N_17336,N_16160,N_16702);
xnor U17337 (N_17337,N_16594,N_16404);
or U17338 (N_17338,N_16358,N_16349);
nand U17339 (N_17339,N_16532,N_16156);
and U17340 (N_17340,N_16405,N_16114);
nand U17341 (N_17341,N_16490,N_16035);
nor U17342 (N_17342,N_16989,N_16391);
and U17343 (N_17343,N_16085,N_16971);
nor U17344 (N_17344,N_16012,N_16382);
or U17345 (N_17345,N_16986,N_16485);
xnor U17346 (N_17346,N_16637,N_16195);
xnor U17347 (N_17347,N_16296,N_16733);
nor U17348 (N_17348,N_16747,N_16858);
nor U17349 (N_17349,N_16477,N_16201);
and U17350 (N_17350,N_16439,N_16465);
nor U17351 (N_17351,N_16519,N_16047);
xor U17352 (N_17352,N_16397,N_16320);
or U17353 (N_17353,N_16432,N_16895);
xnor U17354 (N_17354,N_16440,N_16392);
or U17355 (N_17355,N_16992,N_16872);
nor U17356 (N_17356,N_16520,N_16592);
or U17357 (N_17357,N_16991,N_16402);
and U17358 (N_17358,N_16619,N_16650);
xnor U17359 (N_17359,N_16180,N_16869);
or U17360 (N_17360,N_16648,N_16187);
nor U17361 (N_17361,N_16148,N_16250);
nor U17362 (N_17362,N_16786,N_16691);
xnor U17363 (N_17363,N_16260,N_16007);
or U17364 (N_17364,N_16172,N_16557);
or U17365 (N_17365,N_16225,N_16795);
xnor U17366 (N_17366,N_16928,N_16071);
xnor U17367 (N_17367,N_16678,N_16601);
nand U17368 (N_17368,N_16101,N_16294);
or U17369 (N_17369,N_16910,N_16823);
nand U17370 (N_17370,N_16332,N_16414);
nor U17371 (N_17371,N_16848,N_16698);
nand U17372 (N_17372,N_16813,N_16409);
or U17373 (N_17373,N_16284,N_16779);
nor U17374 (N_17374,N_16548,N_16163);
or U17375 (N_17375,N_16615,N_16609);
and U17376 (N_17376,N_16562,N_16107);
nand U17377 (N_17377,N_16967,N_16276);
nand U17378 (N_17378,N_16213,N_16001);
or U17379 (N_17379,N_16011,N_16951);
nor U17380 (N_17380,N_16906,N_16949);
nand U17381 (N_17381,N_16436,N_16886);
and U17382 (N_17382,N_16807,N_16032);
nor U17383 (N_17383,N_16460,N_16653);
nand U17384 (N_17384,N_16599,N_16330);
or U17385 (N_17385,N_16996,N_16132);
and U17386 (N_17386,N_16396,N_16400);
and U17387 (N_17387,N_16929,N_16044);
or U17388 (N_17388,N_16269,N_16463);
xor U17389 (N_17389,N_16752,N_16891);
nor U17390 (N_17390,N_16569,N_16022);
nand U17391 (N_17391,N_16009,N_16386);
or U17392 (N_17392,N_16920,N_16970);
or U17393 (N_17393,N_16496,N_16509);
or U17394 (N_17394,N_16655,N_16383);
or U17395 (N_17395,N_16288,N_16004);
nand U17396 (N_17396,N_16335,N_16394);
nand U17397 (N_17397,N_16774,N_16926);
nand U17398 (N_17398,N_16964,N_16590);
nand U17399 (N_17399,N_16218,N_16838);
and U17400 (N_17400,N_16281,N_16692);
xor U17401 (N_17401,N_16448,N_16566);
nor U17402 (N_17402,N_16080,N_16741);
xnor U17403 (N_17403,N_16685,N_16091);
nand U17404 (N_17404,N_16611,N_16173);
nor U17405 (N_17405,N_16235,N_16591);
nor U17406 (N_17406,N_16508,N_16943);
and U17407 (N_17407,N_16043,N_16958);
xnor U17408 (N_17408,N_16484,N_16961);
or U17409 (N_17409,N_16675,N_16890);
xnor U17410 (N_17410,N_16855,N_16036);
nor U17411 (N_17411,N_16430,N_16016);
nor U17412 (N_17412,N_16622,N_16189);
and U17413 (N_17413,N_16987,N_16835);
nand U17414 (N_17414,N_16129,N_16380);
nor U17415 (N_17415,N_16897,N_16789);
nor U17416 (N_17416,N_16265,N_16262);
or U17417 (N_17417,N_16353,N_16889);
xor U17418 (N_17418,N_16551,N_16343);
nor U17419 (N_17419,N_16295,N_16750);
or U17420 (N_17420,N_16941,N_16337);
or U17421 (N_17421,N_16395,N_16688);
nor U17422 (N_17422,N_16344,N_16816);
and U17423 (N_17423,N_16304,N_16960);
nand U17424 (N_17424,N_16552,N_16275);
nor U17425 (N_17425,N_16641,N_16474);
and U17426 (N_17426,N_16868,N_16287);
xor U17427 (N_17427,N_16576,N_16892);
and U17428 (N_17428,N_16887,N_16055);
nand U17429 (N_17429,N_16538,N_16185);
xor U17430 (N_17430,N_16109,N_16112);
or U17431 (N_17431,N_16306,N_16363);
nand U17432 (N_17432,N_16579,N_16930);
nand U17433 (N_17433,N_16123,N_16431);
and U17434 (N_17434,N_16308,N_16598);
or U17435 (N_17435,N_16760,N_16135);
nand U17436 (N_17436,N_16863,N_16196);
nor U17437 (N_17437,N_16517,N_16672);
nor U17438 (N_17438,N_16663,N_16820);
or U17439 (N_17439,N_16957,N_16610);
nand U17440 (N_17440,N_16056,N_16338);
nand U17441 (N_17441,N_16236,N_16618);
and U17442 (N_17442,N_16923,N_16529);
nor U17443 (N_17443,N_16190,N_16003);
nor U17444 (N_17444,N_16270,N_16680);
and U17445 (N_17445,N_16324,N_16979);
xnor U17446 (N_17446,N_16556,N_16166);
and U17447 (N_17447,N_16200,N_16738);
xor U17448 (N_17448,N_16057,N_16279);
nor U17449 (N_17449,N_16487,N_16526);
nor U17450 (N_17450,N_16976,N_16727);
xnor U17451 (N_17451,N_16939,N_16652);
and U17452 (N_17452,N_16687,N_16682);
xor U17453 (N_17453,N_16792,N_16612);
and U17454 (N_17454,N_16183,N_16776);
nand U17455 (N_17455,N_16137,N_16425);
nand U17456 (N_17456,N_16645,N_16000);
nor U17457 (N_17457,N_16985,N_16817);
or U17458 (N_17458,N_16608,N_16791);
or U17459 (N_17459,N_16034,N_16586);
or U17460 (N_17460,N_16456,N_16345);
xnor U17461 (N_17461,N_16511,N_16507);
or U17462 (N_17462,N_16925,N_16140);
and U17463 (N_17463,N_16461,N_16224);
or U17464 (N_17464,N_16922,N_16900);
xnor U17465 (N_17465,N_16127,N_16515);
nor U17466 (N_17466,N_16829,N_16157);
and U17467 (N_17467,N_16952,N_16972);
nand U17468 (N_17468,N_16896,N_16082);
nand U17469 (N_17469,N_16819,N_16954);
nand U17470 (N_17470,N_16742,N_16604);
or U17471 (N_17471,N_16334,N_16130);
xnor U17472 (N_17472,N_16378,N_16772);
nand U17473 (N_17473,N_16909,N_16469);
xor U17474 (N_17474,N_16023,N_16937);
nor U17475 (N_17475,N_16885,N_16794);
nor U17476 (N_17476,N_16037,N_16821);
nand U17477 (N_17477,N_16852,N_16089);
nand U17478 (N_17478,N_16437,N_16472);
and U17479 (N_17479,N_16503,N_16959);
and U17480 (N_17480,N_16778,N_16367);
xor U17481 (N_17481,N_16522,N_16564);
or U17482 (N_17482,N_16903,N_16339);
or U17483 (N_17483,N_16151,N_16888);
xnor U17484 (N_17484,N_16362,N_16587);
nand U17485 (N_17485,N_16266,N_16327);
and U17486 (N_17486,N_16828,N_16595);
xnor U17487 (N_17487,N_16029,N_16120);
nor U17488 (N_17488,N_16677,N_16694);
xnor U17489 (N_17489,N_16981,N_16068);
and U17490 (N_17490,N_16310,N_16072);
and U17491 (N_17491,N_16026,N_16365);
or U17492 (N_17492,N_16844,N_16013);
nand U17493 (N_17493,N_16104,N_16944);
and U17494 (N_17494,N_16459,N_16550);
or U17495 (N_17495,N_16931,N_16884);
nor U17496 (N_17496,N_16481,N_16316);
or U17497 (N_17497,N_16720,N_16570);
nand U17498 (N_17498,N_16442,N_16879);
or U17499 (N_17499,N_16656,N_16783);
xnor U17500 (N_17500,N_16566,N_16428);
nor U17501 (N_17501,N_16037,N_16316);
xor U17502 (N_17502,N_16430,N_16082);
nand U17503 (N_17503,N_16114,N_16251);
nor U17504 (N_17504,N_16500,N_16936);
nand U17505 (N_17505,N_16274,N_16053);
and U17506 (N_17506,N_16206,N_16009);
and U17507 (N_17507,N_16599,N_16328);
and U17508 (N_17508,N_16307,N_16984);
nor U17509 (N_17509,N_16487,N_16555);
or U17510 (N_17510,N_16111,N_16094);
nor U17511 (N_17511,N_16533,N_16847);
or U17512 (N_17512,N_16787,N_16625);
nand U17513 (N_17513,N_16897,N_16223);
xor U17514 (N_17514,N_16431,N_16918);
or U17515 (N_17515,N_16839,N_16781);
and U17516 (N_17516,N_16000,N_16633);
xnor U17517 (N_17517,N_16892,N_16882);
or U17518 (N_17518,N_16483,N_16056);
nand U17519 (N_17519,N_16034,N_16668);
nor U17520 (N_17520,N_16311,N_16604);
and U17521 (N_17521,N_16703,N_16142);
nor U17522 (N_17522,N_16872,N_16142);
or U17523 (N_17523,N_16741,N_16290);
or U17524 (N_17524,N_16643,N_16732);
nand U17525 (N_17525,N_16482,N_16427);
or U17526 (N_17526,N_16188,N_16909);
nor U17527 (N_17527,N_16066,N_16812);
xnor U17528 (N_17528,N_16120,N_16919);
nor U17529 (N_17529,N_16658,N_16555);
nand U17530 (N_17530,N_16417,N_16806);
nand U17531 (N_17531,N_16455,N_16897);
nand U17532 (N_17532,N_16198,N_16113);
and U17533 (N_17533,N_16859,N_16866);
nor U17534 (N_17534,N_16728,N_16929);
nor U17535 (N_17535,N_16001,N_16309);
nand U17536 (N_17536,N_16745,N_16006);
nor U17537 (N_17537,N_16290,N_16027);
nor U17538 (N_17538,N_16503,N_16601);
or U17539 (N_17539,N_16927,N_16186);
or U17540 (N_17540,N_16211,N_16154);
and U17541 (N_17541,N_16178,N_16479);
or U17542 (N_17542,N_16644,N_16887);
xnor U17543 (N_17543,N_16128,N_16798);
nor U17544 (N_17544,N_16383,N_16702);
or U17545 (N_17545,N_16658,N_16650);
nor U17546 (N_17546,N_16499,N_16096);
or U17547 (N_17547,N_16610,N_16195);
nor U17548 (N_17548,N_16471,N_16923);
nor U17549 (N_17549,N_16877,N_16489);
nand U17550 (N_17550,N_16371,N_16688);
xnor U17551 (N_17551,N_16189,N_16143);
xor U17552 (N_17552,N_16697,N_16631);
and U17553 (N_17553,N_16610,N_16692);
xor U17554 (N_17554,N_16747,N_16572);
nor U17555 (N_17555,N_16442,N_16321);
or U17556 (N_17556,N_16837,N_16299);
nand U17557 (N_17557,N_16214,N_16410);
and U17558 (N_17558,N_16337,N_16037);
or U17559 (N_17559,N_16567,N_16674);
nand U17560 (N_17560,N_16316,N_16039);
nand U17561 (N_17561,N_16793,N_16263);
and U17562 (N_17562,N_16296,N_16349);
xor U17563 (N_17563,N_16484,N_16688);
xor U17564 (N_17564,N_16786,N_16189);
nor U17565 (N_17565,N_16087,N_16531);
nand U17566 (N_17566,N_16606,N_16566);
xor U17567 (N_17567,N_16368,N_16892);
nor U17568 (N_17568,N_16170,N_16889);
xnor U17569 (N_17569,N_16097,N_16051);
and U17570 (N_17570,N_16997,N_16850);
and U17571 (N_17571,N_16536,N_16341);
nor U17572 (N_17572,N_16455,N_16420);
xor U17573 (N_17573,N_16227,N_16854);
xor U17574 (N_17574,N_16728,N_16688);
xnor U17575 (N_17575,N_16215,N_16916);
nand U17576 (N_17576,N_16740,N_16345);
xor U17577 (N_17577,N_16564,N_16687);
nor U17578 (N_17578,N_16648,N_16392);
xnor U17579 (N_17579,N_16697,N_16953);
and U17580 (N_17580,N_16559,N_16649);
and U17581 (N_17581,N_16008,N_16300);
nand U17582 (N_17582,N_16686,N_16235);
nand U17583 (N_17583,N_16844,N_16696);
and U17584 (N_17584,N_16817,N_16562);
or U17585 (N_17585,N_16111,N_16174);
xor U17586 (N_17586,N_16052,N_16301);
or U17587 (N_17587,N_16844,N_16137);
xor U17588 (N_17588,N_16585,N_16702);
nand U17589 (N_17589,N_16073,N_16237);
nand U17590 (N_17590,N_16476,N_16978);
nor U17591 (N_17591,N_16825,N_16277);
and U17592 (N_17592,N_16287,N_16750);
or U17593 (N_17593,N_16494,N_16455);
nor U17594 (N_17594,N_16433,N_16048);
and U17595 (N_17595,N_16037,N_16941);
or U17596 (N_17596,N_16937,N_16585);
or U17597 (N_17597,N_16310,N_16661);
nor U17598 (N_17598,N_16808,N_16206);
and U17599 (N_17599,N_16593,N_16195);
nand U17600 (N_17600,N_16590,N_16334);
nor U17601 (N_17601,N_16266,N_16557);
or U17602 (N_17602,N_16549,N_16181);
or U17603 (N_17603,N_16901,N_16563);
nor U17604 (N_17604,N_16943,N_16583);
or U17605 (N_17605,N_16476,N_16835);
nand U17606 (N_17606,N_16183,N_16471);
and U17607 (N_17607,N_16156,N_16216);
nor U17608 (N_17608,N_16469,N_16562);
or U17609 (N_17609,N_16541,N_16643);
nand U17610 (N_17610,N_16777,N_16085);
nor U17611 (N_17611,N_16693,N_16852);
nand U17612 (N_17612,N_16189,N_16252);
xor U17613 (N_17613,N_16294,N_16741);
and U17614 (N_17614,N_16212,N_16206);
nand U17615 (N_17615,N_16949,N_16971);
nor U17616 (N_17616,N_16654,N_16347);
and U17617 (N_17617,N_16485,N_16993);
and U17618 (N_17618,N_16176,N_16337);
xor U17619 (N_17619,N_16390,N_16522);
nand U17620 (N_17620,N_16901,N_16854);
xnor U17621 (N_17621,N_16497,N_16877);
and U17622 (N_17622,N_16032,N_16248);
nor U17623 (N_17623,N_16264,N_16011);
nand U17624 (N_17624,N_16687,N_16052);
nand U17625 (N_17625,N_16367,N_16483);
nor U17626 (N_17626,N_16433,N_16948);
nand U17627 (N_17627,N_16223,N_16420);
xor U17628 (N_17628,N_16894,N_16756);
xor U17629 (N_17629,N_16830,N_16757);
nand U17630 (N_17630,N_16934,N_16164);
xnor U17631 (N_17631,N_16522,N_16643);
and U17632 (N_17632,N_16791,N_16508);
nor U17633 (N_17633,N_16071,N_16113);
nand U17634 (N_17634,N_16044,N_16048);
xnor U17635 (N_17635,N_16573,N_16716);
or U17636 (N_17636,N_16103,N_16757);
or U17637 (N_17637,N_16682,N_16286);
xor U17638 (N_17638,N_16174,N_16450);
or U17639 (N_17639,N_16583,N_16994);
xnor U17640 (N_17640,N_16057,N_16879);
nor U17641 (N_17641,N_16996,N_16098);
or U17642 (N_17642,N_16400,N_16242);
or U17643 (N_17643,N_16453,N_16548);
xor U17644 (N_17644,N_16108,N_16360);
nor U17645 (N_17645,N_16153,N_16359);
nand U17646 (N_17646,N_16734,N_16085);
or U17647 (N_17647,N_16017,N_16072);
nand U17648 (N_17648,N_16521,N_16661);
nand U17649 (N_17649,N_16281,N_16130);
xor U17650 (N_17650,N_16112,N_16964);
and U17651 (N_17651,N_16457,N_16093);
xor U17652 (N_17652,N_16618,N_16768);
xnor U17653 (N_17653,N_16707,N_16464);
nor U17654 (N_17654,N_16413,N_16357);
xor U17655 (N_17655,N_16297,N_16722);
and U17656 (N_17656,N_16885,N_16992);
or U17657 (N_17657,N_16939,N_16934);
xnor U17658 (N_17658,N_16969,N_16637);
nor U17659 (N_17659,N_16148,N_16699);
and U17660 (N_17660,N_16996,N_16963);
and U17661 (N_17661,N_16668,N_16287);
nor U17662 (N_17662,N_16938,N_16913);
nor U17663 (N_17663,N_16365,N_16100);
nand U17664 (N_17664,N_16171,N_16407);
and U17665 (N_17665,N_16155,N_16475);
nand U17666 (N_17666,N_16916,N_16467);
and U17667 (N_17667,N_16929,N_16450);
and U17668 (N_17668,N_16869,N_16447);
nor U17669 (N_17669,N_16314,N_16261);
nor U17670 (N_17670,N_16322,N_16584);
xor U17671 (N_17671,N_16416,N_16508);
or U17672 (N_17672,N_16674,N_16174);
xnor U17673 (N_17673,N_16206,N_16165);
or U17674 (N_17674,N_16853,N_16141);
and U17675 (N_17675,N_16919,N_16284);
nand U17676 (N_17676,N_16227,N_16412);
nand U17677 (N_17677,N_16310,N_16082);
nand U17678 (N_17678,N_16761,N_16919);
nor U17679 (N_17679,N_16441,N_16547);
nand U17680 (N_17680,N_16782,N_16593);
nand U17681 (N_17681,N_16842,N_16640);
or U17682 (N_17682,N_16512,N_16518);
nand U17683 (N_17683,N_16183,N_16717);
or U17684 (N_17684,N_16655,N_16592);
xor U17685 (N_17685,N_16926,N_16411);
xor U17686 (N_17686,N_16989,N_16223);
xnor U17687 (N_17687,N_16651,N_16778);
xor U17688 (N_17688,N_16610,N_16539);
and U17689 (N_17689,N_16348,N_16746);
nand U17690 (N_17690,N_16702,N_16947);
and U17691 (N_17691,N_16040,N_16607);
and U17692 (N_17692,N_16970,N_16895);
and U17693 (N_17693,N_16289,N_16383);
nor U17694 (N_17694,N_16729,N_16206);
and U17695 (N_17695,N_16357,N_16229);
and U17696 (N_17696,N_16476,N_16137);
and U17697 (N_17697,N_16263,N_16217);
or U17698 (N_17698,N_16662,N_16898);
nand U17699 (N_17699,N_16110,N_16476);
or U17700 (N_17700,N_16806,N_16163);
xor U17701 (N_17701,N_16880,N_16743);
and U17702 (N_17702,N_16341,N_16728);
xor U17703 (N_17703,N_16792,N_16478);
and U17704 (N_17704,N_16531,N_16924);
or U17705 (N_17705,N_16757,N_16398);
or U17706 (N_17706,N_16983,N_16954);
and U17707 (N_17707,N_16119,N_16198);
xnor U17708 (N_17708,N_16930,N_16381);
nor U17709 (N_17709,N_16662,N_16515);
and U17710 (N_17710,N_16189,N_16881);
xor U17711 (N_17711,N_16895,N_16252);
nand U17712 (N_17712,N_16358,N_16809);
nor U17713 (N_17713,N_16709,N_16966);
nand U17714 (N_17714,N_16634,N_16238);
nor U17715 (N_17715,N_16829,N_16246);
xor U17716 (N_17716,N_16229,N_16745);
xnor U17717 (N_17717,N_16757,N_16806);
nor U17718 (N_17718,N_16577,N_16388);
nor U17719 (N_17719,N_16723,N_16213);
nand U17720 (N_17720,N_16192,N_16755);
or U17721 (N_17721,N_16038,N_16110);
or U17722 (N_17722,N_16629,N_16846);
nor U17723 (N_17723,N_16570,N_16518);
nor U17724 (N_17724,N_16983,N_16365);
nor U17725 (N_17725,N_16703,N_16516);
and U17726 (N_17726,N_16331,N_16136);
and U17727 (N_17727,N_16728,N_16046);
and U17728 (N_17728,N_16542,N_16620);
xnor U17729 (N_17729,N_16233,N_16559);
xnor U17730 (N_17730,N_16455,N_16347);
nor U17731 (N_17731,N_16408,N_16713);
nand U17732 (N_17732,N_16353,N_16424);
nand U17733 (N_17733,N_16443,N_16844);
or U17734 (N_17734,N_16526,N_16131);
and U17735 (N_17735,N_16592,N_16051);
and U17736 (N_17736,N_16385,N_16103);
and U17737 (N_17737,N_16951,N_16650);
nor U17738 (N_17738,N_16450,N_16485);
nor U17739 (N_17739,N_16355,N_16890);
or U17740 (N_17740,N_16565,N_16043);
nand U17741 (N_17741,N_16416,N_16914);
nor U17742 (N_17742,N_16081,N_16085);
nand U17743 (N_17743,N_16366,N_16713);
and U17744 (N_17744,N_16728,N_16378);
or U17745 (N_17745,N_16100,N_16477);
nand U17746 (N_17746,N_16525,N_16576);
nor U17747 (N_17747,N_16019,N_16549);
nor U17748 (N_17748,N_16561,N_16813);
nor U17749 (N_17749,N_16616,N_16357);
nor U17750 (N_17750,N_16754,N_16714);
and U17751 (N_17751,N_16151,N_16290);
or U17752 (N_17752,N_16149,N_16445);
nand U17753 (N_17753,N_16334,N_16054);
xor U17754 (N_17754,N_16947,N_16817);
and U17755 (N_17755,N_16407,N_16332);
nand U17756 (N_17756,N_16214,N_16883);
nand U17757 (N_17757,N_16103,N_16296);
xnor U17758 (N_17758,N_16671,N_16394);
xnor U17759 (N_17759,N_16448,N_16044);
or U17760 (N_17760,N_16754,N_16355);
nor U17761 (N_17761,N_16724,N_16191);
xnor U17762 (N_17762,N_16966,N_16348);
and U17763 (N_17763,N_16918,N_16702);
xnor U17764 (N_17764,N_16111,N_16960);
xnor U17765 (N_17765,N_16671,N_16976);
and U17766 (N_17766,N_16837,N_16152);
and U17767 (N_17767,N_16438,N_16788);
nor U17768 (N_17768,N_16934,N_16579);
xnor U17769 (N_17769,N_16184,N_16514);
nand U17770 (N_17770,N_16501,N_16991);
and U17771 (N_17771,N_16793,N_16507);
nand U17772 (N_17772,N_16992,N_16379);
nand U17773 (N_17773,N_16490,N_16766);
or U17774 (N_17774,N_16853,N_16056);
nand U17775 (N_17775,N_16425,N_16341);
nor U17776 (N_17776,N_16918,N_16035);
xor U17777 (N_17777,N_16959,N_16619);
or U17778 (N_17778,N_16959,N_16573);
or U17779 (N_17779,N_16017,N_16416);
xor U17780 (N_17780,N_16017,N_16084);
or U17781 (N_17781,N_16868,N_16527);
and U17782 (N_17782,N_16133,N_16841);
nor U17783 (N_17783,N_16648,N_16831);
or U17784 (N_17784,N_16234,N_16548);
nand U17785 (N_17785,N_16011,N_16750);
and U17786 (N_17786,N_16548,N_16578);
or U17787 (N_17787,N_16717,N_16874);
and U17788 (N_17788,N_16385,N_16637);
nor U17789 (N_17789,N_16916,N_16704);
nor U17790 (N_17790,N_16914,N_16391);
xor U17791 (N_17791,N_16679,N_16530);
nor U17792 (N_17792,N_16123,N_16780);
nor U17793 (N_17793,N_16670,N_16973);
or U17794 (N_17794,N_16568,N_16244);
xor U17795 (N_17795,N_16619,N_16452);
and U17796 (N_17796,N_16005,N_16304);
or U17797 (N_17797,N_16796,N_16456);
nand U17798 (N_17798,N_16790,N_16533);
nor U17799 (N_17799,N_16305,N_16689);
xor U17800 (N_17800,N_16313,N_16946);
nand U17801 (N_17801,N_16015,N_16737);
or U17802 (N_17802,N_16719,N_16125);
nand U17803 (N_17803,N_16426,N_16388);
nand U17804 (N_17804,N_16050,N_16840);
xor U17805 (N_17805,N_16080,N_16736);
and U17806 (N_17806,N_16447,N_16057);
xor U17807 (N_17807,N_16447,N_16243);
xnor U17808 (N_17808,N_16639,N_16679);
and U17809 (N_17809,N_16489,N_16201);
xor U17810 (N_17810,N_16393,N_16533);
and U17811 (N_17811,N_16522,N_16959);
or U17812 (N_17812,N_16468,N_16422);
nand U17813 (N_17813,N_16464,N_16269);
and U17814 (N_17814,N_16083,N_16243);
xnor U17815 (N_17815,N_16362,N_16589);
and U17816 (N_17816,N_16950,N_16691);
or U17817 (N_17817,N_16250,N_16168);
nand U17818 (N_17818,N_16430,N_16098);
or U17819 (N_17819,N_16816,N_16252);
nor U17820 (N_17820,N_16446,N_16871);
xnor U17821 (N_17821,N_16146,N_16576);
or U17822 (N_17822,N_16659,N_16021);
xnor U17823 (N_17823,N_16322,N_16723);
and U17824 (N_17824,N_16990,N_16835);
nand U17825 (N_17825,N_16576,N_16845);
xor U17826 (N_17826,N_16781,N_16246);
nor U17827 (N_17827,N_16062,N_16710);
xnor U17828 (N_17828,N_16513,N_16335);
nand U17829 (N_17829,N_16451,N_16323);
nand U17830 (N_17830,N_16282,N_16196);
nand U17831 (N_17831,N_16003,N_16273);
xor U17832 (N_17832,N_16760,N_16175);
xnor U17833 (N_17833,N_16250,N_16843);
xor U17834 (N_17834,N_16139,N_16458);
or U17835 (N_17835,N_16028,N_16741);
or U17836 (N_17836,N_16424,N_16535);
and U17837 (N_17837,N_16842,N_16369);
nand U17838 (N_17838,N_16047,N_16964);
and U17839 (N_17839,N_16537,N_16452);
and U17840 (N_17840,N_16570,N_16826);
nor U17841 (N_17841,N_16336,N_16740);
nor U17842 (N_17842,N_16823,N_16788);
and U17843 (N_17843,N_16187,N_16969);
or U17844 (N_17844,N_16279,N_16184);
xor U17845 (N_17845,N_16857,N_16343);
xnor U17846 (N_17846,N_16089,N_16539);
nor U17847 (N_17847,N_16370,N_16213);
or U17848 (N_17848,N_16001,N_16459);
nand U17849 (N_17849,N_16161,N_16847);
or U17850 (N_17850,N_16747,N_16574);
nand U17851 (N_17851,N_16832,N_16716);
nor U17852 (N_17852,N_16189,N_16419);
nor U17853 (N_17853,N_16689,N_16763);
xnor U17854 (N_17854,N_16368,N_16900);
and U17855 (N_17855,N_16976,N_16472);
or U17856 (N_17856,N_16306,N_16044);
nor U17857 (N_17857,N_16613,N_16594);
nor U17858 (N_17858,N_16189,N_16711);
and U17859 (N_17859,N_16415,N_16635);
or U17860 (N_17860,N_16668,N_16687);
xnor U17861 (N_17861,N_16401,N_16744);
nand U17862 (N_17862,N_16195,N_16117);
xor U17863 (N_17863,N_16141,N_16574);
xnor U17864 (N_17864,N_16429,N_16312);
xnor U17865 (N_17865,N_16559,N_16420);
nand U17866 (N_17866,N_16957,N_16825);
or U17867 (N_17867,N_16330,N_16871);
and U17868 (N_17868,N_16036,N_16726);
xnor U17869 (N_17869,N_16628,N_16270);
or U17870 (N_17870,N_16267,N_16855);
and U17871 (N_17871,N_16822,N_16435);
or U17872 (N_17872,N_16094,N_16809);
xnor U17873 (N_17873,N_16566,N_16023);
and U17874 (N_17874,N_16543,N_16434);
nor U17875 (N_17875,N_16620,N_16888);
nand U17876 (N_17876,N_16162,N_16656);
and U17877 (N_17877,N_16579,N_16041);
and U17878 (N_17878,N_16674,N_16634);
nand U17879 (N_17879,N_16024,N_16068);
nor U17880 (N_17880,N_16231,N_16749);
or U17881 (N_17881,N_16396,N_16894);
nor U17882 (N_17882,N_16717,N_16131);
nand U17883 (N_17883,N_16505,N_16001);
and U17884 (N_17884,N_16922,N_16801);
or U17885 (N_17885,N_16338,N_16698);
nor U17886 (N_17886,N_16916,N_16027);
or U17887 (N_17887,N_16884,N_16672);
or U17888 (N_17888,N_16820,N_16110);
nor U17889 (N_17889,N_16359,N_16092);
xnor U17890 (N_17890,N_16253,N_16179);
and U17891 (N_17891,N_16364,N_16932);
nor U17892 (N_17892,N_16181,N_16426);
xor U17893 (N_17893,N_16709,N_16142);
nand U17894 (N_17894,N_16885,N_16787);
and U17895 (N_17895,N_16686,N_16646);
nor U17896 (N_17896,N_16927,N_16108);
and U17897 (N_17897,N_16499,N_16073);
and U17898 (N_17898,N_16041,N_16456);
xor U17899 (N_17899,N_16717,N_16600);
or U17900 (N_17900,N_16795,N_16680);
or U17901 (N_17901,N_16596,N_16401);
xor U17902 (N_17902,N_16583,N_16747);
and U17903 (N_17903,N_16293,N_16980);
nor U17904 (N_17904,N_16113,N_16779);
and U17905 (N_17905,N_16747,N_16340);
xnor U17906 (N_17906,N_16578,N_16573);
nand U17907 (N_17907,N_16324,N_16872);
nor U17908 (N_17908,N_16552,N_16161);
xnor U17909 (N_17909,N_16901,N_16330);
xnor U17910 (N_17910,N_16568,N_16670);
nor U17911 (N_17911,N_16357,N_16309);
and U17912 (N_17912,N_16606,N_16928);
or U17913 (N_17913,N_16130,N_16469);
or U17914 (N_17914,N_16525,N_16869);
and U17915 (N_17915,N_16293,N_16857);
nor U17916 (N_17916,N_16230,N_16553);
and U17917 (N_17917,N_16512,N_16879);
nand U17918 (N_17918,N_16403,N_16324);
or U17919 (N_17919,N_16919,N_16377);
xor U17920 (N_17920,N_16574,N_16244);
nand U17921 (N_17921,N_16775,N_16451);
nor U17922 (N_17922,N_16135,N_16198);
xnor U17923 (N_17923,N_16727,N_16699);
xor U17924 (N_17924,N_16970,N_16598);
or U17925 (N_17925,N_16436,N_16263);
and U17926 (N_17926,N_16875,N_16386);
and U17927 (N_17927,N_16554,N_16382);
nor U17928 (N_17928,N_16220,N_16333);
nor U17929 (N_17929,N_16353,N_16425);
and U17930 (N_17930,N_16699,N_16224);
and U17931 (N_17931,N_16444,N_16641);
xnor U17932 (N_17932,N_16843,N_16529);
or U17933 (N_17933,N_16509,N_16106);
nand U17934 (N_17934,N_16959,N_16795);
xnor U17935 (N_17935,N_16719,N_16181);
and U17936 (N_17936,N_16909,N_16371);
and U17937 (N_17937,N_16625,N_16655);
nand U17938 (N_17938,N_16552,N_16932);
or U17939 (N_17939,N_16153,N_16449);
nand U17940 (N_17940,N_16228,N_16544);
or U17941 (N_17941,N_16614,N_16388);
or U17942 (N_17942,N_16299,N_16911);
nor U17943 (N_17943,N_16226,N_16338);
nand U17944 (N_17944,N_16302,N_16882);
xnor U17945 (N_17945,N_16138,N_16536);
or U17946 (N_17946,N_16657,N_16587);
and U17947 (N_17947,N_16123,N_16181);
xor U17948 (N_17948,N_16182,N_16208);
nand U17949 (N_17949,N_16888,N_16680);
xor U17950 (N_17950,N_16275,N_16808);
nand U17951 (N_17951,N_16824,N_16105);
xnor U17952 (N_17952,N_16831,N_16409);
or U17953 (N_17953,N_16268,N_16384);
nor U17954 (N_17954,N_16240,N_16239);
nand U17955 (N_17955,N_16682,N_16497);
and U17956 (N_17956,N_16717,N_16598);
and U17957 (N_17957,N_16261,N_16810);
or U17958 (N_17958,N_16754,N_16789);
xor U17959 (N_17959,N_16964,N_16637);
nand U17960 (N_17960,N_16911,N_16265);
xor U17961 (N_17961,N_16962,N_16944);
and U17962 (N_17962,N_16685,N_16112);
xnor U17963 (N_17963,N_16712,N_16332);
and U17964 (N_17964,N_16046,N_16401);
and U17965 (N_17965,N_16828,N_16803);
nor U17966 (N_17966,N_16552,N_16362);
xor U17967 (N_17967,N_16276,N_16504);
or U17968 (N_17968,N_16383,N_16608);
nor U17969 (N_17969,N_16426,N_16465);
xor U17970 (N_17970,N_16339,N_16344);
and U17971 (N_17971,N_16745,N_16164);
or U17972 (N_17972,N_16870,N_16409);
nor U17973 (N_17973,N_16758,N_16986);
xor U17974 (N_17974,N_16070,N_16563);
and U17975 (N_17975,N_16864,N_16757);
nor U17976 (N_17976,N_16589,N_16026);
nand U17977 (N_17977,N_16604,N_16370);
xnor U17978 (N_17978,N_16413,N_16550);
nor U17979 (N_17979,N_16266,N_16355);
nor U17980 (N_17980,N_16014,N_16213);
nor U17981 (N_17981,N_16882,N_16058);
nor U17982 (N_17982,N_16990,N_16869);
xnor U17983 (N_17983,N_16453,N_16412);
nor U17984 (N_17984,N_16347,N_16855);
nand U17985 (N_17985,N_16102,N_16688);
and U17986 (N_17986,N_16458,N_16859);
nand U17987 (N_17987,N_16745,N_16891);
nand U17988 (N_17988,N_16342,N_16227);
nor U17989 (N_17989,N_16683,N_16329);
nand U17990 (N_17990,N_16641,N_16186);
nand U17991 (N_17991,N_16824,N_16847);
and U17992 (N_17992,N_16547,N_16744);
nand U17993 (N_17993,N_16650,N_16605);
nor U17994 (N_17994,N_16266,N_16111);
and U17995 (N_17995,N_16986,N_16364);
nor U17996 (N_17996,N_16357,N_16906);
and U17997 (N_17997,N_16573,N_16032);
nand U17998 (N_17998,N_16021,N_16867);
xnor U17999 (N_17999,N_16943,N_16060);
xor U18000 (N_18000,N_17593,N_17592);
xnor U18001 (N_18001,N_17737,N_17029);
or U18002 (N_18002,N_17343,N_17287);
nor U18003 (N_18003,N_17021,N_17251);
nor U18004 (N_18004,N_17570,N_17858);
xor U18005 (N_18005,N_17361,N_17863);
nor U18006 (N_18006,N_17012,N_17900);
nor U18007 (N_18007,N_17846,N_17149);
or U18008 (N_18008,N_17991,N_17365);
or U18009 (N_18009,N_17183,N_17467);
and U18010 (N_18010,N_17627,N_17696);
xor U18011 (N_18011,N_17448,N_17958);
xor U18012 (N_18012,N_17832,N_17612);
nand U18013 (N_18013,N_17165,N_17314);
nor U18014 (N_18014,N_17647,N_17117);
xnor U18015 (N_18015,N_17542,N_17291);
or U18016 (N_18016,N_17013,N_17651);
nand U18017 (N_18017,N_17884,N_17182);
nor U18018 (N_18018,N_17233,N_17814);
nor U18019 (N_18019,N_17600,N_17833);
or U18020 (N_18020,N_17126,N_17247);
and U18021 (N_18021,N_17636,N_17803);
or U18022 (N_18022,N_17129,N_17604);
and U18023 (N_18023,N_17450,N_17209);
and U18024 (N_18024,N_17667,N_17691);
nand U18025 (N_18025,N_17288,N_17828);
and U18026 (N_18026,N_17175,N_17700);
or U18027 (N_18027,N_17329,N_17577);
and U18028 (N_18028,N_17402,N_17718);
or U18029 (N_18029,N_17285,N_17510);
and U18030 (N_18030,N_17644,N_17809);
nor U18031 (N_18031,N_17387,N_17940);
or U18032 (N_18032,N_17692,N_17683);
and U18033 (N_18033,N_17608,N_17877);
or U18034 (N_18034,N_17018,N_17461);
xor U18035 (N_18035,N_17420,N_17249);
or U18036 (N_18036,N_17847,N_17466);
nor U18037 (N_18037,N_17825,N_17163);
nand U18038 (N_18038,N_17802,N_17389);
or U18039 (N_18039,N_17215,N_17845);
nor U18040 (N_18040,N_17630,N_17731);
xnor U18041 (N_18041,N_17048,N_17468);
xnor U18042 (N_18042,N_17722,N_17319);
or U18043 (N_18043,N_17295,N_17167);
nor U18044 (N_18044,N_17200,N_17758);
nand U18045 (N_18045,N_17978,N_17443);
and U18046 (N_18046,N_17697,N_17554);
and U18047 (N_18047,N_17095,N_17837);
or U18048 (N_18048,N_17304,N_17996);
nor U18049 (N_18049,N_17224,N_17426);
or U18050 (N_18050,N_17144,N_17223);
and U18051 (N_18051,N_17123,N_17548);
nand U18052 (N_18052,N_17926,N_17742);
and U18053 (N_18053,N_17830,N_17528);
nand U18054 (N_18054,N_17891,N_17116);
xor U18055 (N_18055,N_17629,N_17072);
and U18056 (N_18056,N_17925,N_17949);
nand U18057 (N_18057,N_17106,N_17975);
xnor U18058 (N_18058,N_17128,N_17646);
nand U18059 (N_18059,N_17195,N_17869);
xor U18060 (N_18060,N_17815,N_17901);
nor U18061 (N_18061,N_17866,N_17055);
nand U18062 (N_18062,N_17039,N_17614);
nor U18063 (N_18063,N_17179,N_17566);
or U18064 (N_18064,N_17171,N_17112);
or U18065 (N_18065,N_17166,N_17313);
and U18066 (N_18066,N_17007,N_17610);
or U18067 (N_18067,N_17491,N_17935);
or U18068 (N_18068,N_17439,N_17801);
nor U18069 (N_18069,N_17005,N_17555);
xor U18070 (N_18070,N_17934,N_17516);
nor U18071 (N_18071,N_17457,N_17244);
nand U18072 (N_18072,N_17198,N_17827);
or U18073 (N_18073,N_17156,N_17130);
nor U18074 (N_18074,N_17841,N_17921);
nor U18075 (N_18075,N_17367,N_17709);
nor U18076 (N_18076,N_17945,N_17536);
and U18077 (N_18077,N_17643,N_17404);
and U18078 (N_18078,N_17196,N_17181);
and U18079 (N_18079,N_17693,N_17660);
nand U18080 (N_18080,N_17435,N_17706);
nor U18081 (N_18081,N_17980,N_17352);
or U18082 (N_18082,N_17458,N_17518);
nor U18083 (N_18083,N_17716,N_17492);
nor U18084 (N_18084,N_17486,N_17987);
xnor U18085 (N_18085,N_17812,N_17872);
nor U18086 (N_18086,N_17037,N_17221);
and U18087 (N_18087,N_17628,N_17730);
or U18088 (N_18088,N_17414,N_17050);
nand U18089 (N_18089,N_17799,N_17559);
and U18090 (N_18090,N_17409,N_17369);
nand U18091 (N_18091,N_17937,N_17587);
nand U18092 (N_18092,N_17246,N_17260);
or U18093 (N_18093,N_17360,N_17893);
and U18094 (N_18094,N_17044,N_17908);
xor U18095 (N_18095,N_17724,N_17805);
or U18096 (N_18096,N_17065,N_17774);
nand U18097 (N_18097,N_17519,N_17652);
or U18098 (N_18098,N_17054,N_17359);
xnor U18099 (N_18099,N_17423,N_17685);
nand U18100 (N_18100,N_17346,N_17194);
and U18101 (N_18101,N_17914,N_17002);
and U18102 (N_18102,N_17428,N_17719);
nand U18103 (N_18103,N_17840,N_17431);
or U18104 (N_18104,N_17063,N_17019);
nand U18105 (N_18105,N_17804,N_17944);
xnor U18106 (N_18106,N_17954,N_17541);
and U18107 (N_18107,N_17424,N_17333);
nand U18108 (N_18108,N_17659,N_17292);
nor U18109 (N_18109,N_17392,N_17595);
or U18110 (N_18110,N_17087,N_17806);
xor U18111 (N_18111,N_17969,N_17856);
or U18112 (N_18112,N_17357,N_17043);
nor U18113 (N_18113,N_17870,N_17701);
xnor U18114 (N_18114,N_17715,N_17464);
and U18115 (N_18115,N_17663,N_17584);
and U18116 (N_18116,N_17120,N_17642);
and U18117 (N_18117,N_17897,N_17421);
and U18118 (N_18118,N_17682,N_17430);
xor U18119 (N_18119,N_17537,N_17680);
nand U18120 (N_18120,N_17698,N_17711);
xor U18121 (N_18121,N_17101,N_17222);
nor U18122 (N_18122,N_17650,N_17531);
xor U18123 (N_18123,N_17155,N_17429);
nor U18124 (N_18124,N_17535,N_17192);
xnor U18125 (N_18125,N_17476,N_17992);
xor U18126 (N_18126,N_17579,N_17546);
xor U18127 (N_18127,N_17558,N_17294);
xnor U18128 (N_18128,N_17765,N_17966);
xor U18129 (N_18129,N_17315,N_17411);
or U18130 (N_18130,N_17245,N_17883);
or U18131 (N_18131,N_17781,N_17523);
xnor U18132 (N_18132,N_17093,N_17318);
and U18133 (N_18133,N_17271,N_17049);
or U18134 (N_18134,N_17511,N_17859);
or U18135 (N_18135,N_17576,N_17817);
and U18136 (N_18136,N_17382,N_17638);
nand U18137 (N_18137,N_17842,N_17772);
nand U18138 (N_18138,N_17808,N_17968);
xnor U18139 (N_18139,N_17740,N_17658);
nor U18140 (N_18140,N_17308,N_17977);
xnor U18141 (N_18141,N_17438,N_17427);
nor U18142 (N_18142,N_17540,N_17899);
nor U18143 (N_18143,N_17979,N_17248);
nor U18144 (N_18144,N_17026,N_17796);
and U18145 (N_18145,N_17059,N_17092);
xnor U18146 (N_18146,N_17826,N_17052);
and U18147 (N_18147,N_17316,N_17490);
nor U18148 (N_18148,N_17342,N_17205);
nand U18149 (N_18149,N_17985,N_17906);
xnor U18150 (N_18150,N_17177,N_17415);
xor U18151 (N_18151,N_17227,N_17533);
and U18152 (N_18152,N_17383,N_17390);
xnor U18153 (N_18153,N_17960,N_17241);
nor U18154 (N_18154,N_17494,N_17606);
xnor U18155 (N_18155,N_17391,N_17916);
nor U18156 (N_18156,N_17732,N_17907);
xor U18157 (N_18157,N_17851,N_17797);
and U18158 (N_18158,N_17634,N_17407);
nor U18159 (N_18159,N_17376,N_17143);
or U18160 (N_18160,N_17347,N_17560);
xnor U18161 (N_18161,N_17720,N_17855);
nor U18162 (N_18162,N_17964,N_17211);
or U18163 (N_18163,N_17372,N_17097);
xnor U18164 (N_18164,N_17405,N_17904);
and U18165 (N_18165,N_17734,N_17524);
nand U18166 (N_18166,N_17505,N_17232);
nor U18167 (N_18167,N_17930,N_17728);
or U18168 (N_18168,N_17004,N_17578);
xnor U18169 (N_18169,N_17556,N_17860);
nor U18170 (N_18170,N_17497,N_17836);
xnor U18171 (N_18171,N_17514,N_17989);
nor U18172 (N_18172,N_17483,N_17867);
xnor U18173 (N_18173,N_17823,N_17296);
xor U18174 (N_18174,N_17947,N_17838);
and U18175 (N_18175,N_17437,N_17290);
or U18176 (N_18176,N_17127,N_17366);
and U18177 (N_18177,N_17334,N_17010);
nand U18178 (N_18178,N_17626,N_17780);
or U18179 (N_18179,N_17707,N_17413);
nor U18180 (N_18180,N_17521,N_17950);
and U18181 (N_18181,N_17132,N_17034);
nand U18182 (N_18182,N_17114,N_17140);
and U18183 (N_18183,N_17498,N_17076);
and U18184 (N_18184,N_17588,N_17278);
nand U18185 (N_18185,N_17264,N_17023);
xor U18186 (N_18186,N_17027,N_17375);
and U18187 (N_18187,N_17527,N_17480);
or U18188 (N_18188,N_17180,N_17664);
or U18189 (N_18189,N_17136,N_17613);
nand U18190 (N_18190,N_17024,N_17670);
xnor U18191 (N_18191,N_17206,N_17263);
nor U18192 (N_18192,N_17311,N_17714);
or U18193 (N_18193,N_17882,N_17911);
nand U18194 (N_18194,N_17539,N_17293);
and U18195 (N_18195,N_17621,N_17253);
nor U18196 (N_18196,N_17761,N_17948);
or U18197 (N_18197,N_17990,N_17506);
nand U18198 (N_18198,N_17124,N_17214);
nand U18199 (N_18199,N_17553,N_17096);
and U18200 (N_18200,N_17225,N_17862);
or U18201 (N_18201,N_17432,N_17008);
nand U18202 (N_18202,N_17125,N_17905);
and U18203 (N_18203,N_17150,N_17635);
xor U18204 (N_18204,N_17082,N_17605);
xor U18205 (N_18205,N_17547,N_17673);
or U18206 (N_18206,N_17928,N_17080);
nor U18207 (N_18207,N_17003,N_17993);
xor U18208 (N_18208,N_17850,N_17481);
xnor U18209 (N_18209,N_17028,N_17186);
or U18210 (N_18210,N_17035,N_17220);
nand U18211 (N_18211,N_17060,N_17751);
nand U18212 (N_18212,N_17786,N_17148);
and U18213 (N_18213,N_17077,N_17695);
xnor U18214 (N_18214,N_17199,N_17561);
or U18215 (N_18215,N_17289,N_17190);
nor U18216 (N_18216,N_17831,N_17640);
xnor U18217 (N_18217,N_17079,N_17267);
and U18218 (N_18218,N_17040,N_17704);
xor U18219 (N_18219,N_17623,N_17662);
nor U18220 (N_18220,N_17756,N_17754);
nand U18221 (N_18221,N_17477,N_17009);
and U18222 (N_18222,N_17504,N_17164);
and U18223 (N_18223,N_17385,N_17403);
or U18224 (N_18224,N_17237,N_17834);
and U18225 (N_18225,N_17456,N_17378);
nand U18226 (N_18226,N_17967,N_17508);
and U18227 (N_18227,N_17568,N_17653);
xnor U18228 (N_18228,N_17912,N_17299);
nor U18229 (N_18229,N_17469,N_17145);
nand U18230 (N_18230,N_17699,N_17956);
xor U18231 (N_18231,N_17522,N_17580);
nor U18232 (N_18232,N_17401,N_17572);
nand U18233 (N_18233,N_17564,N_17777);
or U18234 (N_18234,N_17793,N_17417);
and U18235 (N_18235,N_17589,N_17368);
xnor U18236 (N_18236,N_17999,N_17871);
nand U18237 (N_18237,N_17460,N_17813);
nor U18238 (N_18238,N_17800,N_17567);
xor U18239 (N_18239,N_17513,N_17455);
and U18240 (N_18240,N_17345,N_17938);
xor U18241 (N_18241,N_17810,N_17876);
xor U18242 (N_18242,N_17064,N_17303);
or U18243 (N_18243,N_17771,N_17344);
xnor U18244 (N_18244,N_17534,N_17529);
nand U18245 (N_18245,N_17686,N_17672);
xor U18246 (N_18246,N_17549,N_17807);
nor U18247 (N_18247,N_17231,N_17203);
or U18248 (N_18248,N_17103,N_17723);
nor U18249 (N_18249,N_17852,N_17955);
and U18250 (N_18250,N_17084,N_17773);
nand U18251 (N_18251,N_17500,N_17440);
nand U18252 (N_18252,N_17000,N_17759);
or U18253 (N_18253,N_17787,N_17573);
xnor U18254 (N_18254,N_17743,N_17351);
nand U18255 (N_18255,N_17708,N_17767);
or U18256 (N_18256,N_17769,N_17675);
or U18257 (N_18257,N_17962,N_17462);
nand U18258 (N_18258,N_17109,N_17075);
or U18259 (N_18259,N_17482,N_17277);
nand U18260 (N_18260,N_17370,N_17433);
xor U18261 (N_18261,N_17425,N_17972);
nor U18262 (N_18262,N_17998,N_17868);
and U18263 (N_18263,N_17137,N_17768);
nand U18264 (N_18264,N_17835,N_17110);
xor U18265 (N_18265,N_17274,N_17412);
or U18266 (N_18266,N_17001,N_17472);
xor U18267 (N_18267,N_17281,N_17317);
nand U18268 (N_18268,N_17113,N_17622);
xor U18269 (N_18269,N_17543,N_17353);
nor U18270 (N_18270,N_17894,N_17961);
and U18271 (N_18271,N_17762,N_17509);
and U18272 (N_18272,N_17590,N_17265);
nor U18273 (N_18273,N_17441,N_17408);
and U18274 (N_18274,N_17074,N_17208);
and U18275 (N_18275,N_17121,N_17268);
and U18276 (N_18276,N_17364,N_17615);
xor U18277 (N_18277,N_17550,N_17393);
xor U18278 (N_18278,N_17666,N_17158);
and U18279 (N_18279,N_17187,N_17406);
xnor U18280 (N_18280,N_17301,N_17920);
nand U18281 (N_18281,N_17434,N_17735);
nand U18282 (N_18282,N_17104,N_17350);
or U18283 (N_18283,N_17887,N_17058);
xnor U18284 (N_18284,N_17300,N_17388);
nor U18285 (N_18285,N_17485,N_17377);
or U18286 (N_18286,N_17286,N_17645);
nor U18287 (N_18287,N_17684,N_17445);
nand U18288 (N_18288,N_17085,N_17396);
and U18289 (N_18289,N_17229,N_17849);
nor U18290 (N_18290,N_17363,N_17162);
and U18291 (N_18291,N_17824,N_17976);
and U18292 (N_18292,N_17349,N_17380);
nand U18293 (N_18293,N_17465,N_17478);
or U18294 (N_18294,N_17325,N_17878);
and U18295 (N_18295,N_17282,N_17599);
nand U18296 (N_18296,N_17874,N_17655);
nor U18297 (N_18297,N_17459,N_17083);
and U18298 (N_18298,N_17302,N_17499);
xnor U18299 (N_18299,N_17184,N_17896);
xor U18300 (N_18300,N_17532,N_17710);
xor U18301 (N_18301,N_17782,N_17086);
or U18302 (N_18302,N_17262,N_17853);
nor U18303 (N_18303,N_17020,N_17603);
xnor U18304 (N_18304,N_17811,N_17471);
and U18305 (N_18305,N_17631,N_17170);
and U18306 (N_18306,N_17067,N_17503);
nand U18307 (N_18307,N_17705,N_17596);
nand U18308 (N_18308,N_17160,N_17254);
xnor U18309 (N_18309,N_17111,N_17910);
and U18310 (N_18310,N_17520,N_17875);
nor U18311 (N_18311,N_17918,N_17108);
or U18312 (N_18312,N_17261,N_17749);
and U18313 (N_18313,N_17105,N_17168);
nor U18314 (N_18314,N_17755,N_17942);
nor U18315 (N_18315,N_17197,N_17270);
nor U18316 (N_18316,N_17562,N_17217);
nor U18317 (N_18317,N_17854,N_17792);
or U18318 (N_18318,N_17679,N_17131);
nand U18319 (N_18319,N_17014,N_17931);
xor U18320 (N_18320,N_17202,N_17974);
nand U18321 (N_18321,N_17178,N_17135);
or U18322 (N_18322,N_17620,N_17051);
or U18323 (N_18323,N_17422,N_17753);
nand U18324 (N_18324,N_17641,N_17436);
nor U18325 (N_18325,N_17848,N_17046);
nor U18326 (N_18326,N_17933,N_17530);
or U18327 (N_18327,N_17310,N_17927);
xor U18328 (N_18328,N_17922,N_17169);
nor U18329 (N_18329,N_17864,N_17747);
and U18330 (N_18330,N_17212,N_17218);
nand U18331 (N_18331,N_17795,N_17517);
nor U18332 (N_18332,N_17453,N_17057);
or U18333 (N_18333,N_17507,N_17098);
xnor U18334 (N_18334,N_17726,N_17449);
or U18335 (N_18335,N_17791,N_17818);
nand U18336 (N_18336,N_17141,N_17022);
xnor U18337 (N_18337,N_17915,N_17242);
or U18338 (N_18338,N_17873,N_17677);
xnor U18339 (N_18339,N_17902,N_17502);
nor U18340 (N_18340,N_17031,N_17844);
nor U18341 (N_18341,N_17495,N_17280);
and U18342 (N_18342,N_17757,N_17235);
nor U18343 (N_18343,N_17102,N_17965);
and U18344 (N_18344,N_17624,N_17829);
xor U18345 (N_18345,N_17172,N_17207);
xnor U18346 (N_18346,N_17702,N_17821);
nor U18347 (N_18347,N_17088,N_17690);
nor U18348 (N_18348,N_17094,N_17358);
xnor U18349 (N_18349,N_17474,N_17888);
xor U18350 (N_18350,N_17775,N_17038);
and U18351 (N_18351,N_17475,N_17115);
nor U18352 (N_18352,N_17748,N_17997);
or U18353 (N_18353,N_17939,N_17678);
nand U18354 (N_18354,N_17419,N_17721);
nor U18355 (N_18355,N_17011,N_17591);
nand U18356 (N_18356,N_17146,N_17488);
xor U18357 (N_18357,N_17886,N_17784);
xnor U18358 (N_18358,N_17323,N_17913);
nor U18359 (N_18359,N_17397,N_17321);
nor U18360 (N_18360,N_17654,N_17879);
and U18361 (N_18361,N_17881,N_17618);
nand U18362 (N_18362,N_17671,N_17783);
nand U18363 (N_18363,N_17307,N_17006);
nor U18364 (N_18364,N_17236,N_17332);
and U18365 (N_18365,N_17741,N_17442);
nand U18366 (N_18366,N_17750,N_17661);
or U18367 (N_18367,N_17305,N_17416);
nor U18368 (N_18368,N_17946,N_17609);
and U18369 (N_18369,N_17032,N_17272);
xor U18370 (N_18370,N_17790,N_17681);
xnor U18371 (N_18371,N_17496,N_17250);
and U18372 (N_18372,N_17586,N_17033);
and U18373 (N_18373,N_17725,N_17030);
xor U18374 (N_18374,N_17982,N_17766);
nor U18375 (N_18375,N_17061,N_17258);
nor U18376 (N_18376,N_17276,N_17070);
and U18377 (N_18377,N_17736,N_17138);
or U18378 (N_18378,N_17694,N_17484);
or U18379 (N_18379,N_17569,N_17374);
and U18380 (N_18380,N_17400,N_17326);
or U18381 (N_18381,N_17788,N_17703);
nor U18382 (N_18382,N_17252,N_17355);
nand U18383 (N_18383,N_17598,N_17986);
xnor U18384 (N_18384,N_17571,N_17994);
or U18385 (N_18385,N_17036,N_17760);
nor U18386 (N_18386,N_17119,N_17099);
nand U18387 (N_18387,N_17228,N_17118);
and U18388 (N_18388,N_17776,N_17189);
nand U18389 (N_18389,N_17889,N_17712);
and U18390 (N_18390,N_17373,N_17957);
xor U18391 (N_18391,N_17959,N_17238);
or U18392 (N_18392,N_17885,N_17487);
and U18393 (N_18393,N_17895,N_17234);
or U18394 (N_18394,N_17473,N_17384);
xor U18395 (N_18395,N_17582,N_17257);
and U18396 (N_18396,N_17341,N_17557);
xor U18397 (N_18397,N_17924,N_17327);
or U18398 (N_18398,N_17575,N_17335);
nor U18399 (N_18399,N_17193,N_17770);
and U18400 (N_18400,N_17594,N_17066);
xor U18401 (N_18401,N_17279,N_17454);
or U18402 (N_18402,N_17995,N_17356);
and U18403 (N_18403,N_17213,N_17607);
nor U18404 (N_18404,N_17953,N_17139);
xnor U18405 (N_18405,N_17324,N_17399);
nand U18406 (N_18406,N_17340,N_17665);
xnor U18407 (N_18407,N_17988,N_17015);
nand U18408 (N_18408,N_17493,N_17574);
and U18409 (N_18409,N_17919,N_17689);
nor U18410 (N_18410,N_17619,N_17047);
and U18411 (N_18411,N_17648,N_17284);
and U18412 (N_18412,N_17107,N_17071);
nor U18413 (N_18413,N_17379,N_17880);
xnor U18414 (N_18414,N_17243,N_17789);
and U18415 (N_18415,N_17744,N_17738);
nand U18416 (N_18416,N_17226,N_17688);
or U18417 (N_18417,N_17045,N_17339);
nor U18418 (N_18418,N_17746,N_17625);
or U18419 (N_18419,N_17822,N_17134);
nand U18420 (N_18420,N_17779,N_17597);
nor U18421 (N_18421,N_17336,N_17585);
nand U18422 (N_18422,N_17053,N_17544);
xor U18423 (N_18423,N_17210,N_17565);
and U18424 (N_18424,N_17159,N_17923);
or U18425 (N_18425,N_17929,N_17410);
and U18426 (N_18426,N_17551,N_17941);
nor U18427 (N_18427,N_17298,N_17312);
and U18428 (N_18428,N_17444,N_17328);
or U18429 (N_18429,N_17963,N_17563);
or U18430 (N_18430,N_17078,N_17983);
nor U18431 (N_18431,N_17151,N_17525);
or U18432 (N_18432,N_17616,N_17451);
nand U18433 (N_18433,N_17632,N_17639);
nand U18434 (N_18434,N_17637,N_17778);
nand U18435 (N_18435,N_17297,N_17185);
or U18436 (N_18436,N_17337,N_17331);
nor U18437 (N_18437,N_17256,N_17479);
xor U18438 (N_18438,N_17676,N_17191);
or U18439 (N_18439,N_17068,N_17239);
and U18440 (N_18440,N_17843,N_17042);
xnor U18441 (N_18441,N_17794,N_17552);
and U18442 (N_18442,N_17240,N_17970);
xnor U18443 (N_18443,N_17489,N_17752);
xnor U18444 (N_18444,N_17656,N_17739);
nor U18445 (N_18445,N_17362,N_17330);
or U18446 (N_18446,N_17745,N_17157);
nand U18447 (N_18447,N_17538,N_17090);
xor U18448 (N_18448,N_17386,N_17657);
xor U18449 (N_18449,N_17371,N_17674);
xnor U18450 (N_18450,N_17819,N_17259);
xnor U18451 (N_18451,N_17016,N_17602);
and U18452 (N_18452,N_17216,N_17152);
and U18453 (N_18453,N_17898,N_17091);
and U18454 (N_18454,N_17501,N_17201);
xnor U18455 (N_18455,N_17951,N_17943);
nand U18456 (N_18456,N_17173,N_17581);
xnor U18457 (N_18457,N_17729,N_17122);
and U18458 (N_18458,N_17269,N_17649);
or U18459 (N_18459,N_17447,N_17266);
xnor U18460 (N_18460,N_17764,N_17633);
xnor U18461 (N_18461,N_17348,N_17394);
and U18462 (N_18462,N_17526,N_17446);
or U18463 (N_18463,N_17320,N_17418);
nand U18464 (N_18464,N_17717,N_17981);
nor U18465 (N_18465,N_17611,N_17176);
nand U18466 (N_18466,N_17865,N_17973);
xor U18467 (N_18467,N_17069,N_17230);
or U18468 (N_18468,N_17154,N_17909);
and U18469 (N_18469,N_17153,N_17395);
nor U18470 (N_18470,N_17452,N_17669);
or U18471 (N_18471,N_17255,N_17275);
nor U18472 (N_18472,N_17617,N_17041);
nor U18473 (N_18473,N_17984,N_17583);
nor U18474 (N_18474,N_17381,N_17073);
and U18475 (N_18475,N_17798,N_17890);
nand U18476 (N_18476,N_17161,N_17785);
nand U18477 (N_18477,N_17816,N_17515);
nor U18478 (N_18478,N_17219,N_17273);
xnor U18479 (N_18479,N_17545,N_17903);
or U18480 (N_18480,N_17763,N_17174);
xnor U18481 (N_18481,N_17971,N_17056);
nor U18482 (N_18482,N_17283,N_17062);
nor U18483 (N_18483,N_17089,N_17306);
nor U18484 (N_18484,N_17025,N_17727);
or U18485 (N_18485,N_17512,N_17713);
or U18486 (N_18486,N_17952,N_17733);
nand U18487 (N_18487,N_17398,N_17017);
and U18488 (N_18488,N_17839,N_17188);
or U18489 (N_18489,N_17601,N_17892);
nand U18490 (N_18490,N_17861,N_17932);
and U18491 (N_18491,N_17463,N_17857);
and U18492 (N_18492,N_17470,N_17081);
xnor U18493 (N_18493,N_17338,N_17309);
nand U18494 (N_18494,N_17917,N_17100);
and U18495 (N_18495,N_17354,N_17204);
nand U18496 (N_18496,N_17147,N_17668);
or U18497 (N_18497,N_17142,N_17322);
and U18498 (N_18498,N_17687,N_17936);
nor U18499 (N_18499,N_17820,N_17133);
xnor U18500 (N_18500,N_17752,N_17724);
or U18501 (N_18501,N_17721,N_17916);
xor U18502 (N_18502,N_17018,N_17660);
nand U18503 (N_18503,N_17911,N_17136);
xnor U18504 (N_18504,N_17739,N_17610);
nor U18505 (N_18505,N_17194,N_17574);
or U18506 (N_18506,N_17236,N_17923);
and U18507 (N_18507,N_17466,N_17753);
and U18508 (N_18508,N_17943,N_17759);
or U18509 (N_18509,N_17524,N_17391);
nor U18510 (N_18510,N_17048,N_17687);
xnor U18511 (N_18511,N_17347,N_17723);
or U18512 (N_18512,N_17232,N_17152);
xor U18513 (N_18513,N_17173,N_17867);
xor U18514 (N_18514,N_17705,N_17164);
nor U18515 (N_18515,N_17853,N_17940);
nor U18516 (N_18516,N_17404,N_17739);
or U18517 (N_18517,N_17201,N_17061);
nor U18518 (N_18518,N_17886,N_17845);
and U18519 (N_18519,N_17700,N_17796);
xor U18520 (N_18520,N_17607,N_17265);
nor U18521 (N_18521,N_17376,N_17385);
nor U18522 (N_18522,N_17022,N_17122);
nor U18523 (N_18523,N_17579,N_17718);
nor U18524 (N_18524,N_17602,N_17264);
nand U18525 (N_18525,N_17925,N_17679);
and U18526 (N_18526,N_17011,N_17744);
or U18527 (N_18527,N_17832,N_17937);
nand U18528 (N_18528,N_17784,N_17763);
nand U18529 (N_18529,N_17471,N_17352);
nor U18530 (N_18530,N_17958,N_17826);
nand U18531 (N_18531,N_17136,N_17669);
nor U18532 (N_18532,N_17214,N_17092);
nand U18533 (N_18533,N_17498,N_17163);
nor U18534 (N_18534,N_17813,N_17248);
xor U18535 (N_18535,N_17208,N_17867);
nor U18536 (N_18536,N_17079,N_17863);
and U18537 (N_18537,N_17238,N_17068);
or U18538 (N_18538,N_17381,N_17678);
nand U18539 (N_18539,N_17376,N_17657);
xor U18540 (N_18540,N_17927,N_17138);
and U18541 (N_18541,N_17022,N_17444);
nand U18542 (N_18542,N_17704,N_17288);
or U18543 (N_18543,N_17959,N_17434);
or U18544 (N_18544,N_17254,N_17111);
nor U18545 (N_18545,N_17698,N_17838);
xnor U18546 (N_18546,N_17564,N_17504);
or U18547 (N_18547,N_17977,N_17998);
nor U18548 (N_18548,N_17453,N_17968);
nand U18549 (N_18549,N_17703,N_17713);
and U18550 (N_18550,N_17485,N_17675);
xnor U18551 (N_18551,N_17603,N_17864);
nand U18552 (N_18552,N_17837,N_17171);
nand U18553 (N_18553,N_17171,N_17129);
nand U18554 (N_18554,N_17485,N_17076);
xor U18555 (N_18555,N_17511,N_17527);
nor U18556 (N_18556,N_17598,N_17397);
and U18557 (N_18557,N_17309,N_17420);
nor U18558 (N_18558,N_17329,N_17937);
and U18559 (N_18559,N_17369,N_17585);
nor U18560 (N_18560,N_17391,N_17878);
nor U18561 (N_18561,N_17711,N_17521);
nor U18562 (N_18562,N_17127,N_17040);
and U18563 (N_18563,N_17450,N_17554);
nor U18564 (N_18564,N_17964,N_17360);
and U18565 (N_18565,N_17805,N_17359);
and U18566 (N_18566,N_17632,N_17181);
nand U18567 (N_18567,N_17466,N_17170);
and U18568 (N_18568,N_17075,N_17050);
nor U18569 (N_18569,N_17915,N_17622);
nand U18570 (N_18570,N_17457,N_17898);
nand U18571 (N_18571,N_17917,N_17865);
xor U18572 (N_18572,N_17932,N_17566);
nand U18573 (N_18573,N_17894,N_17668);
nor U18574 (N_18574,N_17851,N_17454);
nor U18575 (N_18575,N_17356,N_17614);
nand U18576 (N_18576,N_17577,N_17291);
or U18577 (N_18577,N_17117,N_17967);
and U18578 (N_18578,N_17093,N_17604);
nand U18579 (N_18579,N_17510,N_17406);
or U18580 (N_18580,N_17232,N_17992);
and U18581 (N_18581,N_17606,N_17400);
or U18582 (N_18582,N_17318,N_17109);
or U18583 (N_18583,N_17831,N_17391);
or U18584 (N_18584,N_17806,N_17071);
nor U18585 (N_18585,N_17054,N_17561);
or U18586 (N_18586,N_17010,N_17189);
and U18587 (N_18587,N_17474,N_17397);
nor U18588 (N_18588,N_17497,N_17298);
and U18589 (N_18589,N_17736,N_17219);
nand U18590 (N_18590,N_17800,N_17835);
nand U18591 (N_18591,N_17312,N_17937);
or U18592 (N_18592,N_17265,N_17166);
nand U18593 (N_18593,N_17147,N_17250);
nor U18594 (N_18594,N_17023,N_17772);
or U18595 (N_18595,N_17496,N_17950);
nand U18596 (N_18596,N_17596,N_17443);
nand U18597 (N_18597,N_17786,N_17078);
or U18598 (N_18598,N_17517,N_17650);
or U18599 (N_18599,N_17653,N_17139);
xor U18600 (N_18600,N_17699,N_17444);
xnor U18601 (N_18601,N_17119,N_17896);
and U18602 (N_18602,N_17202,N_17870);
nor U18603 (N_18603,N_17935,N_17209);
or U18604 (N_18604,N_17333,N_17240);
nor U18605 (N_18605,N_17793,N_17759);
xnor U18606 (N_18606,N_17430,N_17503);
and U18607 (N_18607,N_17277,N_17833);
or U18608 (N_18608,N_17269,N_17981);
nor U18609 (N_18609,N_17963,N_17172);
and U18610 (N_18610,N_17359,N_17217);
nand U18611 (N_18611,N_17075,N_17130);
nand U18612 (N_18612,N_17014,N_17337);
nand U18613 (N_18613,N_17125,N_17286);
and U18614 (N_18614,N_17081,N_17076);
nand U18615 (N_18615,N_17901,N_17045);
nand U18616 (N_18616,N_17378,N_17839);
nand U18617 (N_18617,N_17889,N_17385);
and U18618 (N_18618,N_17578,N_17589);
xnor U18619 (N_18619,N_17113,N_17274);
nand U18620 (N_18620,N_17891,N_17800);
or U18621 (N_18621,N_17345,N_17948);
xor U18622 (N_18622,N_17452,N_17353);
nand U18623 (N_18623,N_17669,N_17569);
nor U18624 (N_18624,N_17357,N_17476);
and U18625 (N_18625,N_17638,N_17312);
nand U18626 (N_18626,N_17052,N_17843);
nor U18627 (N_18627,N_17931,N_17460);
and U18628 (N_18628,N_17878,N_17446);
or U18629 (N_18629,N_17844,N_17003);
xnor U18630 (N_18630,N_17516,N_17218);
or U18631 (N_18631,N_17283,N_17402);
nand U18632 (N_18632,N_17786,N_17403);
and U18633 (N_18633,N_17928,N_17472);
nor U18634 (N_18634,N_17170,N_17939);
xnor U18635 (N_18635,N_17158,N_17370);
or U18636 (N_18636,N_17972,N_17802);
xor U18637 (N_18637,N_17144,N_17009);
nand U18638 (N_18638,N_17819,N_17403);
xnor U18639 (N_18639,N_17678,N_17712);
nor U18640 (N_18640,N_17480,N_17969);
xor U18641 (N_18641,N_17663,N_17418);
nand U18642 (N_18642,N_17306,N_17416);
nand U18643 (N_18643,N_17642,N_17012);
nor U18644 (N_18644,N_17995,N_17910);
and U18645 (N_18645,N_17200,N_17450);
nand U18646 (N_18646,N_17082,N_17392);
nor U18647 (N_18647,N_17396,N_17715);
or U18648 (N_18648,N_17387,N_17667);
nand U18649 (N_18649,N_17826,N_17284);
nor U18650 (N_18650,N_17813,N_17670);
or U18651 (N_18651,N_17501,N_17683);
and U18652 (N_18652,N_17865,N_17710);
and U18653 (N_18653,N_17182,N_17362);
or U18654 (N_18654,N_17307,N_17170);
xor U18655 (N_18655,N_17160,N_17749);
xnor U18656 (N_18656,N_17904,N_17525);
xnor U18657 (N_18657,N_17011,N_17720);
nor U18658 (N_18658,N_17381,N_17892);
nor U18659 (N_18659,N_17891,N_17061);
nor U18660 (N_18660,N_17129,N_17192);
or U18661 (N_18661,N_17303,N_17123);
or U18662 (N_18662,N_17392,N_17574);
xnor U18663 (N_18663,N_17374,N_17112);
nand U18664 (N_18664,N_17779,N_17013);
nand U18665 (N_18665,N_17567,N_17438);
nand U18666 (N_18666,N_17950,N_17816);
and U18667 (N_18667,N_17049,N_17192);
nand U18668 (N_18668,N_17179,N_17627);
or U18669 (N_18669,N_17314,N_17796);
and U18670 (N_18670,N_17125,N_17258);
or U18671 (N_18671,N_17780,N_17815);
and U18672 (N_18672,N_17508,N_17203);
nor U18673 (N_18673,N_17882,N_17749);
xnor U18674 (N_18674,N_17819,N_17299);
and U18675 (N_18675,N_17557,N_17339);
nand U18676 (N_18676,N_17932,N_17927);
and U18677 (N_18677,N_17307,N_17925);
xnor U18678 (N_18678,N_17457,N_17161);
and U18679 (N_18679,N_17900,N_17807);
xor U18680 (N_18680,N_17754,N_17469);
nor U18681 (N_18681,N_17782,N_17959);
nor U18682 (N_18682,N_17135,N_17377);
or U18683 (N_18683,N_17641,N_17941);
or U18684 (N_18684,N_17507,N_17750);
or U18685 (N_18685,N_17180,N_17692);
xnor U18686 (N_18686,N_17944,N_17435);
and U18687 (N_18687,N_17860,N_17527);
xnor U18688 (N_18688,N_17837,N_17184);
nor U18689 (N_18689,N_17225,N_17075);
xor U18690 (N_18690,N_17242,N_17404);
and U18691 (N_18691,N_17304,N_17707);
and U18692 (N_18692,N_17320,N_17188);
or U18693 (N_18693,N_17822,N_17414);
and U18694 (N_18694,N_17526,N_17692);
nand U18695 (N_18695,N_17729,N_17104);
nor U18696 (N_18696,N_17594,N_17680);
nor U18697 (N_18697,N_17855,N_17231);
nand U18698 (N_18698,N_17455,N_17631);
and U18699 (N_18699,N_17071,N_17371);
xnor U18700 (N_18700,N_17474,N_17821);
and U18701 (N_18701,N_17528,N_17657);
nor U18702 (N_18702,N_17941,N_17347);
nor U18703 (N_18703,N_17145,N_17273);
and U18704 (N_18704,N_17213,N_17127);
xor U18705 (N_18705,N_17721,N_17076);
nor U18706 (N_18706,N_17211,N_17117);
nor U18707 (N_18707,N_17580,N_17571);
nor U18708 (N_18708,N_17321,N_17289);
and U18709 (N_18709,N_17150,N_17433);
and U18710 (N_18710,N_17607,N_17015);
xnor U18711 (N_18711,N_17292,N_17540);
or U18712 (N_18712,N_17027,N_17881);
xor U18713 (N_18713,N_17042,N_17249);
xor U18714 (N_18714,N_17487,N_17151);
nor U18715 (N_18715,N_17948,N_17248);
xnor U18716 (N_18716,N_17896,N_17965);
or U18717 (N_18717,N_17346,N_17516);
nor U18718 (N_18718,N_17191,N_17113);
xor U18719 (N_18719,N_17414,N_17606);
xor U18720 (N_18720,N_17641,N_17133);
xor U18721 (N_18721,N_17725,N_17263);
nor U18722 (N_18722,N_17697,N_17300);
nand U18723 (N_18723,N_17613,N_17907);
xnor U18724 (N_18724,N_17727,N_17179);
nor U18725 (N_18725,N_17988,N_17288);
or U18726 (N_18726,N_17583,N_17820);
xnor U18727 (N_18727,N_17710,N_17885);
xor U18728 (N_18728,N_17849,N_17351);
nor U18729 (N_18729,N_17616,N_17191);
and U18730 (N_18730,N_17955,N_17871);
or U18731 (N_18731,N_17691,N_17750);
and U18732 (N_18732,N_17539,N_17665);
nor U18733 (N_18733,N_17138,N_17882);
nor U18734 (N_18734,N_17194,N_17714);
or U18735 (N_18735,N_17347,N_17694);
or U18736 (N_18736,N_17989,N_17761);
nand U18737 (N_18737,N_17644,N_17325);
xor U18738 (N_18738,N_17434,N_17220);
nor U18739 (N_18739,N_17266,N_17421);
and U18740 (N_18740,N_17676,N_17391);
xor U18741 (N_18741,N_17682,N_17376);
and U18742 (N_18742,N_17033,N_17313);
and U18743 (N_18743,N_17547,N_17035);
and U18744 (N_18744,N_17620,N_17288);
nor U18745 (N_18745,N_17945,N_17151);
nand U18746 (N_18746,N_17597,N_17764);
nor U18747 (N_18747,N_17484,N_17105);
or U18748 (N_18748,N_17868,N_17129);
or U18749 (N_18749,N_17101,N_17377);
nor U18750 (N_18750,N_17258,N_17497);
xnor U18751 (N_18751,N_17978,N_17528);
nand U18752 (N_18752,N_17322,N_17251);
nor U18753 (N_18753,N_17338,N_17868);
nor U18754 (N_18754,N_17553,N_17504);
or U18755 (N_18755,N_17881,N_17762);
or U18756 (N_18756,N_17532,N_17693);
xnor U18757 (N_18757,N_17623,N_17552);
and U18758 (N_18758,N_17927,N_17205);
nand U18759 (N_18759,N_17503,N_17201);
nand U18760 (N_18760,N_17081,N_17080);
nand U18761 (N_18761,N_17496,N_17755);
xnor U18762 (N_18762,N_17377,N_17127);
or U18763 (N_18763,N_17638,N_17781);
and U18764 (N_18764,N_17467,N_17148);
or U18765 (N_18765,N_17688,N_17933);
and U18766 (N_18766,N_17387,N_17097);
nand U18767 (N_18767,N_17920,N_17499);
and U18768 (N_18768,N_17416,N_17133);
and U18769 (N_18769,N_17344,N_17765);
xor U18770 (N_18770,N_17420,N_17831);
xor U18771 (N_18771,N_17885,N_17850);
nor U18772 (N_18772,N_17160,N_17332);
or U18773 (N_18773,N_17748,N_17441);
or U18774 (N_18774,N_17487,N_17053);
nand U18775 (N_18775,N_17523,N_17564);
nand U18776 (N_18776,N_17645,N_17163);
nand U18777 (N_18777,N_17981,N_17163);
xnor U18778 (N_18778,N_17114,N_17130);
nand U18779 (N_18779,N_17544,N_17632);
nor U18780 (N_18780,N_17343,N_17149);
nand U18781 (N_18781,N_17788,N_17894);
and U18782 (N_18782,N_17867,N_17163);
nor U18783 (N_18783,N_17634,N_17131);
xnor U18784 (N_18784,N_17414,N_17906);
nand U18785 (N_18785,N_17562,N_17308);
nand U18786 (N_18786,N_17249,N_17129);
xnor U18787 (N_18787,N_17936,N_17489);
or U18788 (N_18788,N_17111,N_17469);
nand U18789 (N_18789,N_17848,N_17156);
xnor U18790 (N_18790,N_17702,N_17884);
xnor U18791 (N_18791,N_17243,N_17002);
nor U18792 (N_18792,N_17677,N_17208);
nand U18793 (N_18793,N_17544,N_17183);
nand U18794 (N_18794,N_17334,N_17525);
xor U18795 (N_18795,N_17904,N_17346);
and U18796 (N_18796,N_17862,N_17255);
xnor U18797 (N_18797,N_17123,N_17358);
nor U18798 (N_18798,N_17608,N_17587);
xor U18799 (N_18799,N_17199,N_17856);
nand U18800 (N_18800,N_17330,N_17429);
xor U18801 (N_18801,N_17530,N_17068);
xnor U18802 (N_18802,N_17978,N_17549);
xnor U18803 (N_18803,N_17136,N_17637);
nand U18804 (N_18804,N_17808,N_17979);
or U18805 (N_18805,N_17281,N_17889);
and U18806 (N_18806,N_17080,N_17975);
or U18807 (N_18807,N_17968,N_17598);
or U18808 (N_18808,N_17531,N_17832);
and U18809 (N_18809,N_17597,N_17792);
or U18810 (N_18810,N_17705,N_17794);
or U18811 (N_18811,N_17302,N_17684);
or U18812 (N_18812,N_17758,N_17869);
and U18813 (N_18813,N_17437,N_17805);
nor U18814 (N_18814,N_17412,N_17909);
nor U18815 (N_18815,N_17123,N_17977);
nand U18816 (N_18816,N_17837,N_17140);
and U18817 (N_18817,N_17244,N_17148);
nand U18818 (N_18818,N_17690,N_17350);
and U18819 (N_18819,N_17277,N_17473);
and U18820 (N_18820,N_17048,N_17982);
nand U18821 (N_18821,N_17279,N_17285);
nand U18822 (N_18822,N_17995,N_17914);
and U18823 (N_18823,N_17734,N_17463);
or U18824 (N_18824,N_17775,N_17271);
xnor U18825 (N_18825,N_17060,N_17582);
or U18826 (N_18826,N_17355,N_17561);
nand U18827 (N_18827,N_17616,N_17638);
nor U18828 (N_18828,N_17564,N_17370);
nor U18829 (N_18829,N_17927,N_17458);
xor U18830 (N_18830,N_17848,N_17975);
nor U18831 (N_18831,N_17388,N_17672);
nand U18832 (N_18832,N_17308,N_17019);
nor U18833 (N_18833,N_17594,N_17411);
and U18834 (N_18834,N_17524,N_17533);
xor U18835 (N_18835,N_17005,N_17683);
or U18836 (N_18836,N_17030,N_17085);
and U18837 (N_18837,N_17200,N_17745);
or U18838 (N_18838,N_17130,N_17956);
nand U18839 (N_18839,N_17519,N_17405);
nand U18840 (N_18840,N_17638,N_17967);
nor U18841 (N_18841,N_17444,N_17817);
and U18842 (N_18842,N_17314,N_17480);
and U18843 (N_18843,N_17424,N_17968);
nand U18844 (N_18844,N_17043,N_17234);
nand U18845 (N_18845,N_17603,N_17542);
nand U18846 (N_18846,N_17428,N_17193);
xor U18847 (N_18847,N_17649,N_17256);
nand U18848 (N_18848,N_17760,N_17951);
or U18849 (N_18849,N_17953,N_17116);
or U18850 (N_18850,N_17372,N_17096);
and U18851 (N_18851,N_17634,N_17839);
and U18852 (N_18852,N_17640,N_17136);
and U18853 (N_18853,N_17978,N_17704);
or U18854 (N_18854,N_17375,N_17895);
xnor U18855 (N_18855,N_17826,N_17407);
nand U18856 (N_18856,N_17917,N_17500);
nand U18857 (N_18857,N_17027,N_17400);
nor U18858 (N_18858,N_17841,N_17277);
xor U18859 (N_18859,N_17578,N_17990);
nand U18860 (N_18860,N_17693,N_17580);
or U18861 (N_18861,N_17753,N_17431);
xnor U18862 (N_18862,N_17679,N_17328);
xnor U18863 (N_18863,N_17614,N_17407);
and U18864 (N_18864,N_17990,N_17859);
nand U18865 (N_18865,N_17453,N_17529);
nor U18866 (N_18866,N_17104,N_17757);
and U18867 (N_18867,N_17231,N_17018);
nand U18868 (N_18868,N_17364,N_17780);
xor U18869 (N_18869,N_17606,N_17220);
xnor U18870 (N_18870,N_17063,N_17348);
or U18871 (N_18871,N_17564,N_17517);
nand U18872 (N_18872,N_17591,N_17421);
xnor U18873 (N_18873,N_17451,N_17135);
nand U18874 (N_18874,N_17361,N_17112);
nand U18875 (N_18875,N_17626,N_17521);
xnor U18876 (N_18876,N_17301,N_17035);
xnor U18877 (N_18877,N_17628,N_17283);
nand U18878 (N_18878,N_17220,N_17136);
nand U18879 (N_18879,N_17180,N_17987);
nor U18880 (N_18880,N_17037,N_17430);
or U18881 (N_18881,N_17907,N_17452);
xor U18882 (N_18882,N_17367,N_17515);
or U18883 (N_18883,N_17827,N_17361);
nor U18884 (N_18884,N_17395,N_17130);
nand U18885 (N_18885,N_17721,N_17653);
and U18886 (N_18886,N_17478,N_17163);
or U18887 (N_18887,N_17121,N_17202);
nor U18888 (N_18888,N_17895,N_17969);
nand U18889 (N_18889,N_17803,N_17864);
or U18890 (N_18890,N_17872,N_17881);
or U18891 (N_18891,N_17219,N_17758);
and U18892 (N_18892,N_17633,N_17052);
nand U18893 (N_18893,N_17941,N_17386);
and U18894 (N_18894,N_17915,N_17152);
nand U18895 (N_18895,N_17824,N_17631);
nor U18896 (N_18896,N_17532,N_17826);
and U18897 (N_18897,N_17498,N_17499);
nand U18898 (N_18898,N_17927,N_17440);
and U18899 (N_18899,N_17332,N_17952);
nor U18900 (N_18900,N_17277,N_17142);
or U18901 (N_18901,N_17705,N_17027);
or U18902 (N_18902,N_17995,N_17869);
xor U18903 (N_18903,N_17831,N_17156);
or U18904 (N_18904,N_17325,N_17376);
xor U18905 (N_18905,N_17939,N_17044);
xor U18906 (N_18906,N_17253,N_17742);
nor U18907 (N_18907,N_17467,N_17143);
xnor U18908 (N_18908,N_17028,N_17655);
and U18909 (N_18909,N_17482,N_17242);
nand U18910 (N_18910,N_17903,N_17198);
xor U18911 (N_18911,N_17084,N_17797);
nand U18912 (N_18912,N_17501,N_17113);
or U18913 (N_18913,N_17763,N_17927);
nor U18914 (N_18914,N_17014,N_17148);
nor U18915 (N_18915,N_17552,N_17498);
or U18916 (N_18916,N_17914,N_17631);
or U18917 (N_18917,N_17191,N_17453);
and U18918 (N_18918,N_17596,N_17471);
nand U18919 (N_18919,N_17893,N_17156);
nand U18920 (N_18920,N_17545,N_17214);
and U18921 (N_18921,N_17083,N_17557);
or U18922 (N_18922,N_17961,N_17866);
or U18923 (N_18923,N_17615,N_17955);
nand U18924 (N_18924,N_17089,N_17353);
nand U18925 (N_18925,N_17076,N_17200);
xnor U18926 (N_18926,N_17363,N_17967);
xnor U18927 (N_18927,N_17802,N_17209);
or U18928 (N_18928,N_17785,N_17068);
or U18929 (N_18929,N_17520,N_17874);
nor U18930 (N_18930,N_17284,N_17853);
nor U18931 (N_18931,N_17021,N_17555);
nor U18932 (N_18932,N_17662,N_17235);
nand U18933 (N_18933,N_17437,N_17262);
and U18934 (N_18934,N_17701,N_17020);
nand U18935 (N_18935,N_17114,N_17808);
or U18936 (N_18936,N_17653,N_17688);
or U18937 (N_18937,N_17562,N_17945);
nor U18938 (N_18938,N_17728,N_17800);
or U18939 (N_18939,N_17911,N_17348);
and U18940 (N_18940,N_17506,N_17440);
nand U18941 (N_18941,N_17005,N_17855);
and U18942 (N_18942,N_17085,N_17911);
nor U18943 (N_18943,N_17749,N_17135);
nor U18944 (N_18944,N_17609,N_17695);
and U18945 (N_18945,N_17895,N_17825);
nand U18946 (N_18946,N_17686,N_17996);
xor U18947 (N_18947,N_17117,N_17143);
and U18948 (N_18948,N_17634,N_17722);
or U18949 (N_18949,N_17649,N_17519);
nor U18950 (N_18950,N_17302,N_17754);
nor U18951 (N_18951,N_17843,N_17305);
nor U18952 (N_18952,N_17202,N_17292);
nand U18953 (N_18953,N_17640,N_17455);
or U18954 (N_18954,N_17505,N_17819);
nor U18955 (N_18955,N_17956,N_17468);
or U18956 (N_18956,N_17592,N_17435);
nor U18957 (N_18957,N_17779,N_17257);
nor U18958 (N_18958,N_17697,N_17721);
or U18959 (N_18959,N_17374,N_17775);
nor U18960 (N_18960,N_17376,N_17713);
and U18961 (N_18961,N_17951,N_17296);
and U18962 (N_18962,N_17185,N_17412);
nor U18963 (N_18963,N_17829,N_17471);
or U18964 (N_18964,N_17677,N_17930);
nand U18965 (N_18965,N_17315,N_17189);
and U18966 (N_18966,N_17184,N_17116);
xnor U18967 (N_18967,N_17139,N_17688);
nor U18968 (N_18968,N_17107,N_17041);
nor U18969 (N_18969,N_17213,N_17247);
or U18970 (N_18970,N_17643,N_17215);
xnor U18971 (N_18971,N_17443,N_17271);
or U18972 (N_18972,N_17121,N_17531);
xnor U18973 (N_18973,N_17887,N_17925);
xor U18974 (N_18974,N_17743,N_17012);
nor U18975 (N_18975,N_17024,N_17421);
and U18976 (N_18976,N_17097,N_17776);
xnor U18977 (N_18977,N_17923,N_17422);
xor U18978 (N_18978,N_17489,N_17623);
nor U18979 (N_18979,N_17049,N_17072);
xnor U18980 (N_18980,N_17169,N_17364);
xnor U18981 (N_18981,N_17242,N_17170);
nand U18982 (N_18982,N_17877,N_17442);
and U18983 (N_18983,N_17717,N_17643);
or U18984 (N_18984,N_17770,N_17936);
nand U18985 (N_18985,N_17443,N_17157);
and U18986 (N_18986,N_17244,N_17968);
nand U18987 (N_18987,N_17730,N_17096);
xor U18988 (N_18988,N_17003,N_17809);
and U18989 (N_18989,N_17046,N_17661);
nand U18990 (N_18990,N_17859,N_17740);
xnor U18991 (N_18991,N_17203,N_17958);
and U18992 (N_18992,N_17538,N_17833);
or U18993 (N_18993,N_17877,N_17210);
and U18994 (N_18994,N_17328,N_17487);
and U18995 (N_18995,N_17665,N_17721);
nand U18996 (N_18996,N_17426,N_17041);
or U18997 (N_18997,N_17460,N_17464);
nand U18998 (N_18998,N_17629,N_17280);
or U18999 (N_18999,N_17745,N_17643);
and U19000 (N_19000,N_18137,N_18420);
xor U19001 (N_19001,N_18063,N_18117);
xnor U19002 (N_19002,N_18536,N_18730);
or U19003 (N_19003,N_18393,N_18700);
xor U19004 (N_19004,N_18029,N_18292);
and U19005 (N_19005,N_18083,N_18235);
xnor U19006 (N_19006,N_18004,N_18696);
xor U19007 (N_19007,N_18825,N_18974);
and U19008 (N_19008,N_18555,N_18866);
nand U19009 (N_19009,N_18633,N_18512);
nand U19010 (N_19010,N_18734,N_18355);
and U19011 (N_19011,N_18240,N_18964);
nand U19012 (N_19012,N_18546,N_18402);
or U19013 (N_19013,N_18897,N_18035);
and U19014 (N_19014,N_18168,N_18685);
xnor U19015 (N_19015,N_18702,N_18229);
xnor U19016 (N_19016,N_18557,N_18281);
nand U19017 (N_19017,N_18710,N_18648);
nand U19018 (N_19018,N_18698,N_18791);
xnor U19019 (N_19019,N_18826,N_18580);
or U19020 (N_19020,N_18357,N_18829);
nor U19021 (N_19021,N_18712,N_18170);
or U19022 (N_19022,N_18875,N_18819);
nor U19023 (N_19023,N_18216,N_18255);
xnor U19024 (N_19024,N_18461,N_18543);
xor U19025 (N_19025,N_18395,N_18842);
xnor U19026 (N_19026,N_18720,N_18232);
and U19027 (N_19027,N_18195,N_18894);
and U19028 (N_19028,N_18850,N_18244);
nand U19029 (N_19029,N_18697,N_18873);
xnor U19030 (N_19030,N_18532,N_18618);
nand U19031 (N_19031,N_18781,N_18883);
nand U19032 (N_19032,N_18413,N_18201);
and U19033 (N_19033,N_18946,N_18885);
and U19034 (N_19034,N_18677,N_18230);
and U19035 (N_19035,N_18537,N_18373);
nor U19036 (N_19036,N_18878,N_18774);
xnor U19037 (N_19037,N_18835,N_18972);
nand U19038 (N_19038,N_18877,N_18694);
xnor U19039 (N_19039,N_18469,N_18488);
xor U19040 (N_19040,N_18550,N_18114);
or U19041 (N_19041,N_18726,N_18669);
nor U19042 (N_19042,N_18573,N_18160);
and U19043 (N_19043,N_18100,N_18764);
xnor U19044 (N_19044,N_18706,N_18064);
and U19045 (N_19045,N_18735,N_18305);
xnor U19046 (N_19046,N_18300,N_18310);
or U19047 (N_19047,N_18672,N_18338);
xor U19048 (N_19048,N_18335,N_18797);
nor U19049 (N_19049,N_18467,N_18369);
nand U19050 (N_19050,N_18453,N_18777);
xnor U19051 (N_19051,N_18585,N_18602);
and U19052 (N_19052,N_18813,N_18445);
nor U19053 (N_19053,N_18705,N_18760);
or U19054 (N_19054,N_18802,N_18960);
nand U19055 (N_19055,N_18852,N_18379);
xnor U19056 (N_19056,N_18771,N_18458);
nor U19057 (N_19057,N_18107,N_18922);
or U19058 (N_19058,N_18495,N_18994);
nand U19059 (N_19059,N_18456,N_18525);
or U19060 (N_19060,N_18879,N_18851);
nor U19061 (N_19061,N_18646,N_18856);
or U19062 (N_19062,N_18892,N_18208);
nand U19063 (N_19063,N_18221,N_18403);
nor U19064 (N_19064,N_18586,N_18249);
and U19065 (N_19065,N_18020,N_18548);
xor U19066 (N_19066,N_18328,N_18342);
and U19067 (N_19067,N_18803,N_18671);
or U19068 (N_19068,N_18653,N_18845);
and U19069 (N_19069,N_18670,N_18361);
and U19070 (N_19070,N_18407,N_18619);
xor U19071 (N_19071,N_18794,N_18806);
xnor U19072 (N_19072,N_18059,N_18718);
and U19073 (N_19073,N_18193,N_18278);
nand U19074 (N_19074,N_18389,N_18578);
nand U19075 (N_19075,N_18975,N_18641);
nor U19076 (N_19076,N_18891,N_18131);
nand U19077 (N_19077,N_18674,N_18742);
xnor U19078 (N_19078,N_18971,N_18088);
xor U19079 (N_19079,N_18763,N_18606);
nor U19080 (N_19080,N_18583,N_18282);
xor U19081 (N_19081,N_18723,N_18448);
nor U19082 (N_19082,N_18030,N_18787);
and U19083 (N_19083,N_18053,N_18459);
nand U19084 (N_19084,N_18007,N_18758);
and U19085 (N_19085,N_18317,N_18765);
and U19086 (N_19086,N_18098,N_18783);
nand U19087 (N_19087,N_18424,N_18079);
nor U19088 (N_19088,N_18324,N_18350);
or U19089 (N_19089,N_18935,N_18238);
xnor U19090 (N_19090,N_18211,N_18397);
nor U19091 (N_19091,N_18092,N_18487);
nand U19092 (N_19092,N_18754,N_18937);
xnor U19093 (N_19093,N_18655,N_18219);
or U19094 (N_19094,N_18479,N_18101);
nor U19095 (N_19095,N_18486,N_18051);
and U19096 (N_19096,N_18509,N_18880);
nor U19097 (N_19097,N_18108,N_18480);
or U19098 (N_19098,N_18233,N_18534);
nor U19099 (N_19099,N_18273,N_18854);
or U19100 (N_19100,N_18270,N_18628);
nor U19101 (N_19101,N_18419,N_18881);
nor U19102 (N_19102,N_18620,N_18508);
and U19103 (N_19103,N_18034,N_18465);
xor U19104 (N_19104,N_18337,N_18242);
or U19105 (N_19105,N_18567,N_18582);
and U19106 (N_19106,N_18860,N_18267);
nor U19107 (N_19107,N_18776,N_18942);
or U19108 (N_19108,N_18675,N_18316);
nand U19109 (N_19109,N_18524,N_18996);
xnor U19110 (N_19110,N_18128,N_18770);
nand U19111 (N_19111,N_18401,N_18442);
xnor U19112 (N_19112,N_18556,N_18868);
or U19113 (N_19113,N_18591,N_18970);
and U19114 (N_19114,N_18903,N_18625);
and U19115 (N_19115,N_18916,N_18070);
nand U19116 (N_19116,N_18416,N_18306);
nand U19117 (N_19117,N_18999,N_18659);
xnor U19118 (N_19118,N_18045,N_18033);
xnor U19119 (N_19119,N_18717,N_18356);
or U19120 (N_19120,N_18275,N_18535);
nor U19121 (N_19121,N_18027,N_18804);
and U19122 (N_19122,N_18731,N_18336);
xnor U19123 (N_19123,N_18381,N_18222);
and U19124 (N_19124,N_18719,N_18099);
and U19125 (N_19125,N_18500,N_18944);
nand U19126 (N_19126,N_18017,N_18779);
nor U19127 (N_19127,N_18398,N_18388);
nor U19128 (N_19128,N_18786,N_18150);
nor U19129 (N_19129,N_18657,N_18940);
and U19130 (N_19130,N_18713,N_18664);
and U19131 (N_19131,N_18189,N_18977);
nand U19132 (N_19132,N_18539,N_18434);
nand U19133 (N_19133,N_18417,N_18740);
nor U19134 (N_19134,N_18118,N_18483);
nand U19135 (N_19135,N_18234,N_18068);
and U19136 (N_19136,N_18060,N_18482);
and U19137 (N_19137,N_18872,N_18252);
xnor U19138 (N_19138,N_18624,N_18969);
nand U19139 (N_19139,N_18334,N_18440);
or U19140 (N_19140,N_18400,N_18149);
and U19141 (N_19141,N_18236,N_18656);
and U19142 (N_19142,N_18135,N_18176);
and U19143 (N_19143,N_18514,N_18154);
and U19144 (N_19144,N_18595,N_18733);
or U19145 (N_19145,N_18805,N_18186);
or U19146 (N_19146,N_18295,N_18410);
or U19147 (N_19147,N_18206,N_18956);
nor U19148 (N_19148,N_18124,N_18767);
xor U19149 (N_19149,N_18741,N_18490);
nand U19150 (N_19150,N_18976,N_18002);
nor U19151 (N_19151,N_18253,N_18784);
and U19152 (N_19152,N_18287,N_18732);
xnor U19153 (N_19153,N_18950,N_18649);
nand U19154 (N_19154,N_18086,N_18093);
nor U19155 (N_19155,N_18811,N_18988);
nor U19156 (N_19156,N_18485,N_18260);
or U19157 (N_19157,N_18676,N_18914);
or U19158 (N_19158,N_18966,N_18297);
xor U19159 (N_19159,N_18807,N_18691);
or U19160 (N_19160,N_18863,N_18775);
and U19161 (N_19161,N_18184,N_18681);
nor U19162 (N_19162,N_18016,N_18254);
xnor U19163 (N_19163,N_18392,N_18921);
nand U19164 (N_19164,N_18640,N_18967);
or U19165 (N_19165,N_18542,N_18056);
xnor U19166 (N_19166,N_18869,N_18147);
or U19167 (N_19167,N_18477,N_18202);
and U19168 (N_19168,N_18432,N_18443);
nand U19169 (N_19169,N_18982,N_18609);
xnor U19170 (N_19170,N_18951,N_18096);
and U19171 (N_19171,N_18311,N_18642);
xor U19172 (N_19172,N_18048,N_18431);
or U19173 (N_19173,N_18217,N_18279);
nor U19174 (N_19174,N_18464,N_18259);
or U19175 (N_19175,N_18846,N_18614);
and U19176 (N_19176,N_18598,N_18044);
and U19177 (N_19177,N_18849,N_18130);
xnor U19178 (N_19178,N_18204,N_18715);
or U19179 (N_19179,N_18721,N_18836);
or U19180 (N_19180,N_18547,N_18936);
nor U19181 (N_19181,N_18121,N_18394);
nand U19182 (N_19182,N_18899,N_18828);
or U19183 (N_19183,N_18747,N_18180);
xnor U19184 (N_19184,N_18041,N_18841);
and U19185 (N_19185,N_18028,N_18298);
nor U19186 (N_19186,N_18887,N_18608);
nor U19187 (N_19187,N_18954,N_18945);
nor U19188 (N_19188,N_18075,N_18798);
and U19189 (N_19189,N_18927,N_18523);
and U19190 (N_19190,N_18102,N_18521);
or U19191 (N_19191,N_18010,N_18612);
xor U19192 (N_19192,N_18153,N_18889);
nand U19193 (N_19193,N_18895,N_18658);
nand U19194 (N_19194,N_18319,N_18519);
nand U19195 (N_19195,N_18171,N_18687);
nand U19196 (N_19196,N_18009,N_18005);
and U19197 (N_19197,N_18104,N_18055);
nand U19198 (N_19198,N_18579,N_18145);
and U19199 (N_19199,N_18241,N_18593);
nor U19200 (N_19200,N_18981,N_18581);
or U19201 (N_19201,N_18187,N_18663);
nand U19202 (N_19202,N_18882,N_18917);
or U19203 (N_19203,N_18631,N_18227);
nor U19204 (N_19204,N_18066,N_18165);
nor U19205 (N_19205,N_18404,N_18761);
xnor U19206 (N_19206,N_18426,N_18815);
xnor U19207 (N_19207,N_18177,N_18478);
nand U19208 (N_19208,N_18062,N_18264);
nand U19209 (N_19209,N_18637,N_18412);
or U19210 (N_19210,N_18090,N_18644);
xnor U19211 (N_19211,N_18638,N_18837);
xnor U19212 (N_19212,N_18327,N_18576);
nor U19213 (N_19213,N_18665,N_18751);
nor U19214 (N_19214,N_18320,N_18588);
nor U19215 (N_19215,N_18499,N_18908);
and U19216 (N_19216,N_18617,N_18296);
nand U19217 (N_19217,N_18584,N_18294);
nor U19218 (N_19218,N_18823,N_18973);
nand U19219 (N_19219,N_18043,N_18134);
nand U19220 (N_19220,N_18695,N_18623);
and U19221 (N_19221,N_18666,N_18364);
and U19222 (N_19222,N_18630,N_18615);
nand U19223 (N_19223,N_18923,N_18192);
xnor U19224 (N_19224,N_18693,N_18955);
or U19225 (N_19225,N_18446,N_18024);
and U19226 (N_19226,N_18780,N_18587);
and U19227 (N_19227,N_18680,N_18449);
or U19228 (N_19228,N_18329,N_18261);
xor U19229 (N_19229,N_18475,N_18948);
and U19230 (N_19230,N_18330,N_18228);
xor U19231 (N_19231,N_18910,N_18549);
or U19232 (N_19232,N_18569,N_18447);
and U19233 (N_19233,N_18616,N_18961);
and U19234 (N_19234,N_18427,N_18853);
or U19235 (N_19235,N_18941,N_18714);
or U19236 (N_19236,N_18590,N_18900);
and U19237 (N_19237,N_18888,N_18057);
xnor U19238 (N_19238,N_18142,N_18571);
or U19239 (N_19239,N_18513,N_18605);
or U19240 (N_19240,N_18037,N_18861);
and U19241 (N_19241,N_18909,N_18943);
nand U19242 (N_19242,N_18621,N_18289);
nand U19243 (N_19243,N_18358,N_18089);
and U19244 (N_19244,N_18349,N_18678);
nand U19245 (N_19245,N_18643,N_18023);
and U19246 (N_19246,N_18708,N_18790);
and U19247 (N_19247,N_18864,N_18816);
xnor U19248 (N_19248,N_18772,N_18049);
and U19249 (N_19249,N_18172,N_18552);
and U19250 (N_19250,N_18778,N_18709);
xor U19251 (N_19251,N_18871,N_18928);
nand U19252 (N_19252,N_18737,N_18762);
nand U19253 (N_19253,N_18686,N_18566);
xor U19254 (N_19254,N_18155,N_18144);
nor U19255 (N_19255,N_18210,N_18876);
xnor U19256 (N_19256,N_18843,N_18231);
xnor U19257 (N_19257,N_18162,N_18148);
xor U19258 (N_19258,N_18391,N_18188);
or U19259 (N_19259,N_18827,N_18913);
xor U19260 (N_19260,N_18462,N_18736);
nor U19261 (N_19261,N_18354,N_18239);
xnor U19262 (N_19262,N_18346,N_18199);
xnor U19263 (N_19263,N_18245,N_18690);
and U19264 (N_19264,N_18194,N_18484);
nand U19265 (N_19265,N_18901,N_18015);
and U19266 (N_19266,N_18538,N_18930);
xnor U19267 (N_19267,N_18243,N_18505);
nand U19268 (N_19268,N_18476,N_18998);
and U19269 (N_19269,N_18314,N_18990);
and U19270 (N_19270,N_18912,N_18414);
xor U19271 (N_19271,N_18668,N_18387);
or U19272 (N_19272,N_18191,N_18283);
nand U19273 (N_19273,N_18560,N_18793);
xor U19274 (N_19274,N_18257,N_18380);
nand U19275 (N_19275,N_18838,N_18931);
or U19276 (N_19276,N_18529,N_18722);
xor U19277 (N_19277,N_18247,N_18115);
xor U19278 (N_19278,N_18592,N_18012);
and U19279 (N_19279,N_18652,N_18660);
and U19280 (N_19280,N_18237,N_18284);
nor U19281 (N_19281,N_18570,N_18596);
and U19282 (N_19282,N_18366,N_18333);
nand U19283 (N_19283,N_18109,N_18473);
nor U19284 (N_19284,N_18506,N_18603);
xor U19285 (N_19285,N_18810,N_18429);
or U19286 (N_19286,N_18692,N_18067);
xor U19287 (N_19287,N_18220,N_18526);
nand U19288 (N_19288,N_18163,N_18455);
nor U19289 (N_19289,N_18345,N_18745);
nand U19290 (N_19290,N_18906,N_18274);
or U19291 (N_19291,N_18785,N_18157);
or U19292 (N_19292,N_18285,N_18989);
and U19293 (N_19293,N_18510,N_18036);
xor U19294 (N_19294,N_18707,N_18197);
nand U19295 (N_19295,N_18038,N_18520);
xor U19296 (N_19296,N_18701,N_18753);
nand U19297 (N_19297,N_18371,N_18095);
or U19298 (N_19298,N_18933,N_18992);
nor U19299 (N_19299,N_18212,N_18926);
nor U19300 (N_19300,N_18341,N_18046);
and U19301 (N_19301,N_18450,N_18859);
xnor U19302 (N_19302,N_18611,N_18207);
and U19303 (N_19303,N_18932,N_18302);
and U19304 (N_19304,N_18175,N_18301);
or U19305 (N_19305,N_18516,N_18463);
nor U19306 (N_19306,N_18136,N_18303);
nand U19307 (N_19307,N_18980,N_18504);
nor U19308 (N_19308,N_18559,N_18047);
xnor U19309 (N_19309,N_18597,N_18052);
or U19310 (N_19310,N_18498,N_18138);
and U19311 (N_19311,N_18026,N_18452);
and U19312 (N_19312,N_18326,N_18323);
nor U19313 (N_19313,N_18688,N_18439);
and U19314 (N_19314,N_18166,N_18246);
nor U19315 (N_19315,N_18411,N_18437);
or U19316 (N_19316,N_18639,N_18127);
nor U19317 (N_19317,N_18689,N_18082);
nand U19318 (N_19318,N_18087,N_18929);
xor U19319 (N_19319,N_18801,N_18517);
xnor U19320 (N_19320,N_18312,N_18058);
xor U19321 (N_19321,N_18152,N_18120);
nand U19322 (N_19322,N_18789,N_18321);
nor U19323 (N_19323,N_18818,N_18293);
xnor U19324 (N_19324,N_18902,N_18962);
xnor U19325 (N_19325,N_18265,N_18375);
or U19326 (N_19326,N_18531,N_18018);
and U19327 (N_19327,N_18367,N_18000);
nand U19328 (N_19328,N_18073,N_18919);
or U19329 (N_19329,N_18169,N_18574);
xnor U19330 (N_19330,N_18116,N_18792);
xor U19331 (N_19331,N_18179,N_18558);
xor U19332 (N_19332,N_18938,N_18986);
and U19333 (N_19333,N_18979,N_18214);
and U19334 (N_19334,N_18554,N_18481);
and U19335 (N_19335,N_18799,N_18178);
or U19336 (N_19336,N_18377,N_18949);
nor U19337 (N_19337,N_18870,N_18290);
nand U19338 (N_19338,N_18629,N_18418);
xor U19339 (N_19339,N_18812,N_18288);
or U19340 (N_19340,N_18915,N_18182);
nor U19341 (N_19341,N_18286,N_18527);
or U19342 (N_19342,N_18991,N_18308);
nand U19343 (N_19343,N_18081,N_18339);
nor U19344 (N_19344,N_18541,N_18359);
xnor U19345 (N_19345,N_18577,N_18496);
or U19346 (N_19346,N_18146,N_18258);
and U19347 (N_19347,N_18858,N_18280);
xnor U19348 (N_19348,N_18352,N_18025);
xnor U19349 (N_19349,N_18890,N_18080);
nand U19350 (N_19350,N_18351,N_18076);
xnor U19351 (N_19351,N_18224,N_18756);
xnor U19352 (N_19352,N_18291,N_18362);
or U19353 (N_19353,N_18183,N_18441);
or U19354 (N_19354,N_18905,N_18304);
xnor U19355 (N_19355,N_18983,N_18271);
nor U19356 (N_19356,N_18679,N_18752);
nor U19357 (N_19357,N_18167,N_18987);
xnor U19358 (N_19358,N_18491,N_18112);
nand U19359 (N_19359,N_18601,N_18132);
nand U19360 (N_19360,N_18728,N_18645);
or U19361 (N_19361,N_18494,N_18934);
and U19362 (N_19362,N_18021,N_18911);
and U19363 (N_19363,N_18406,N_18110);
nand U19364 (N_19364,N_18551,N_18563);
and U19365 (N_19365,N_18173,N_18968);
or U19366 (N_19366,N_18014,N_18769);
and U19367 (N_19367,N_18632,N_18604);
xor U19368 (N_19368,N_18839,N_18077);
nand U19369 (N_19369,N_18126,N_18435);
or U19370 (N_19370,N_18530,N_18382);
nand U19371 (N_19371,N_18907,N_18262);
nand U19372 (N_19372,N_18074,N_18003);
or U19373 (N_19373,N_18796,N_18097);
xor U19374 (N_19374,N_18190,N_18139);
xor U19375 (N_19375,N_18372,N_18553);
xor U19376 (N_19376,N_18867,N_18203);
or U19377 (N_19377,N_18111,N_18113);
nor U19378 (N_19378,N_18383,N_18276);
and U19379 (N_19379,N_18322,N_18425);
nand U19380 (N_19380,N_18344,N_18353);
or U19381 (N_19381,N_18269,N_18423);
and U19382 (N_19382,N_18782,N_18433);
nor U19383 (N_19383,N_18831,N_18198);
nand U19384 (N_19384,N_18896,N_18143);
xor U19385 (N_19385,N_18748,N_18122);
or U19386 (N_19386,N_18613,N_18457);
nand U19387 (N_19387,N_18474,N_18370);
nand U19388 (N_19388,N_18408,N_18006);
and U19389 (N_19389,N_18847,N_18773);
or U19390 (N_19390,N_18011,N_18865);
or U19391 (N_19391,N_18348,N_18125);
or U19392 (N_19392,N_18958,N_18684);
nor U19393 (N_19393,N_18133,N_18422);
or U19394 (N_19394,N_18492,N_18040);
and U19395 (N_19395,N_18699,N_18716);
and U19396 (N_19396,N_18185,N_18788);
xnor U19397 (N_19397,N_18468,N_18140);
or U19398 (N_19398,N_18156,N_18898);
and U19399 (N_19399,N_18739,N_18251);
or U19400 (N_19400,N_18200,N_18711);
or U19401 (N_19401,N_18084,N_18589);
and U19402 (N_19402,N_18844,N_18743);
or U19403 (N_19403,N_18634,N_18451);
xnor U19404 (N_19404,N_18545,N_18091);
or U19405 (N_19405,N_18503,N_18196);
or U19406 (N_19406,N_18331,N_18065);
nor U19407 (N_19407,N_18054,N_18824);
or U19408 (N_19408,N_18757,N_18385);
nor U19409 (N_19409,N_18248,N_18997);
and U19410 (N_19410,N_18848,N_18834);
xor U19411 (N_19411,N_18572,N_18667);
and U19412 (N_19412,N_18094,N_18340);
or U19413 (N_19413,N_18515,N_18360);
and U19414 (N_19414,N_18993,N_18151);
and U19415 (N_19415,N_18855,N_18309);
or U19416 (N_19416,N_18650,N_18141);
nor U19417 (N_19417,N_18072,N_18744);
nor U19418 (N_19418,N_18978,N_18862);
nor U19419 (N_19419,N_18444,N_18755);
nor U19420 (N_19420,N_18378,N_18959);
or U19421 (N_19421,N_18925,N_18493);
or U19422 (N_19422,N_18750,N_18682);
or U19423 (N_19423,N_18662,N_18085);
or U19424 (N_19424,N_18884,N_18313);
nand U19425 (N_19425,N_18363,N_18218);
or U19426 (N_19426,N_18738,N_18874);
or U19427 (N_19427,N_18471,N_18315);
nand U19428 (N_19428,N_18409,N_18518);
or U19429 (N_19429,N_18307,N_18749);
or U19430 (N_19430,N_18857,N_18565);
nand U19431 (N_19431,N_18820,N_18042);
xnor U19432 (N_19432,N_18032,N_18561);
and U19433 (N_19433,N_18918,N_18399);
xnor U19434 (N_19434,N_18533,N_18390);
nor U19435 (N_19435,N_18318,N_18268);
nand U19436 (N_19436,N_18953,N_18325);
and U19437 (N_19437,N_18647,N_18904);
or U19438 (N_19438,N_18626,N_18161);
or U19439 (N_19439,N_18600,N_18472);
and U19440 (N_19440,N_18939,N_18635);
nor U19441 (N_19441,N_18250,N_18725);
xor U19442 (N_19442,N_18947,N_18421);
xor U19443 (N_19443,N_18522,N_18544);
nor U19444 (N_19444,N_18454,N_18636);
nand U19445 (N_19445,N_18223,N_18466);
nor U19446 (N_19446,N_18768,N_18528);
nor U19447 (N_19447,N_18501,N_18105);
and U19448 (N_19448,N_18575,N_18272);
nor U19449 (N_19449,N_18511,N_18808);
and U19450 (N_19450,N_18022,N_18562);
or U19451 (N_19451,N_18415,N_18123);
and U19452 (N_19452,N_18164,N_18830);
and U19453 (N_19453,N_18800,N_18119);
or U19454 (N_19454,N_18683,N_18226);
or U19455 (N_19455,N_18594,N_18368);
or U19456 (N_19456,N_18001,N_18277);
nor U19457 (N_19457,N_18832,N_18893);
or U19458 (N_19458,N_18822,N_18766);
xor U19459 (N_19459,N_18704,N_18985);
xnor U19460 (N_19460,N_18965,N_18205);
xor U19461 (N_19461,N_18957,N_18489);
or U19462 (N_19462,N_18507,N_18727);
nor U19463 (N_19463,N_18061,N_18031);
or U19464 (N_19464,N_18209,N_18266);
xnor U19465 (N_19465,N_18814,N_18984);
or U19466 (N_19466,N_18396,N_18069);
and U19467 (N_19467,N_18365,N_18746);
xor U19468 (N_19468,N_18158,N_18129);
xnor U19469 (N_19469,N_18174,N_18256);
nor U19470 (N_19470,N_18817,N_18920);
nand U19471 (N_19471,N_18343,N_18995);
nor U19472 (N_19472,N_18430,N_18386);
nand U19473 (N_19473,N_18833,N_18622);
or U19474 (N_19474,N_18039,N_18008);
or U19475 (N_19475,N_18374,N_18263);
nor U19476 (N_19476,N_18729,N_18013);
or U19477 (N_19477,N_18564,N_18071);
and U19478 (N_19478,N_18599,N_18703);
or U19479 (N_19479,N_18050,N_18332);
or U19480 (N_19480,N_18840,N_18299);
nand U19481 (N_19481,N_18502,N_18106);
xor U19482 (N_19482,N_18809,N_18460);
nand U19483 (N_19483,N_18159,N_18497);
xor U19484 (N_19484,N_18952,N_18568);
or U19485 (N_19485,N_18924,N_18795);
or U19486 (N_19486,N_18347,N_18078);
nor U19487 (N_19487,N_18213,N_18376);
or U19488 (N_19488,N_18759,N_18215);
nand U19489 (N_19489,N_18103,N_18724);
or U19490 (N_19490,N_18661,N_18405);
or U19491 (N_19491,N_18181,N_18540);
nor U19492 (N_19492,N_18886,N_18627);
and U19493 (N_19493,N_18651,N_18438);
or U19494 (N_19494,N_18470,N_18019);
or U19495 (N_19495,N_18610,N_18673);
xnor U19496 (N_19496,N_18821,N_18428);
or U19497 (N_19497,N_18384,N_18436);
nand U19498 (N_19498,N_18963,N_18607);
nand U19499 (N_19499,N_18225,N_18654);
nor U19500 (N_19500,N_18199,N_18808);
and U19501 (N_19501,N_18012,N_18676);
nand U19502 (N_19502,N_18526,N_18702);
nand U19503 (N_19503,N_18354,N_18563);
nor U19504 (N_19504,N_18266,N_18125);
nand U19505 (N_19505,N_18214,N_18090);
xnor U19506 (N_19506,N_18945,N_18470);
or U19507 (N_19507,N_18226,N_18636);
and U19508 (N_19508,N_18845,N_18275);
nor U19509 (N_19509,N_18373,N_18497);
xor U19510 (N_19510,N_18976,N_18909);
and U19511 (N_19511,N_18573,N_18806);
nor U19512 (N_19512,N_18848,N_18791);
nand U19513 (N_19513,N_18147,N_18741);
or U19514 (N_19514,N_18855,N_18293);
nand U19515 (N_19515,N_18038,N_18547);
nor U19516 (N_19516,N_18953,N_18383);
nand U19517 (N_19517,N_18276,N_18697);
nand U19518 (N_19518,N_18349,N_18528);
nor U19519 (N_19519,N_18241,N_18809);
nand U19520 (N_19520,N_18397,N_18310);
and U19521 (N_19521,N_18765,N_18164);
and U19522 (N_19522,N_18165,N_18942);
xor U19523 (N_19523,N_18789,N_18722);
and U19524 (N_19524,N_18850,N_18359);
nor U19525 (N_19525,N_18707,N_18753);
xnor U19526 (N_19526,N_18835,N_18630);
xnor U19527 (N_19527,N_18780,N_18506);
nand U19528 (N_19528,N_18001,N_18353);
or U19529 (N_19529,N_18679,N_18008);
xor U19530 (N_19530,N_18689,N_18281);
nor U19531 (N_19531,N_18865,N_18841);
nor U19532 (N_19532,N_18691,N_18675);
xor U19533 (N_19533,N_18125,N_18788);
nand U19534 (N_19534,N_18864,N_18813);
or U19535 (N_19535,N_18128,N_18143);
or U19536 (N_19536,N_18051,N_18435);
xnor U19537 (N_19537,N_18590,N_18874);
nor U19538 (N_19538,N_18858,N_18852);
nand U19539 (N_19539,N_18772,N_18727);
or U19540 (N_19540,N_18680,N_18428);
nand U19541 (N_19541,N_18739,N_18651);
xor U19542 (N_19542,N_18608,N_18215);
or U19543 (N_19543,N_18710,N_18104);
nor U19544 (N_19544,N_18146,N_18648);
and U19545 (N_19545,N_18253,N_18313);
or U19546 (N_19546,N_18534,N_18396);
nor U19547 (N_19547,N_18919,N_18322);
xnor U19548 (N_19548,N_18690,N_18239);
and U19549 (N_19549,N_18311,N_18359);
or U19550 (N_19550,N_18071,N_18693);
nand U19551 (N_19551,N_18472,N_18380);
and U19552 (N_19552,N_18543,N_18805);
and U19553 (N_19553,N_18365,N_18416);
nor U19554 (N_19554,N_18599,N_18057);
nor U19555 (N_19555,N_18507,N_18891);
or U19556 (N_19556,N_18125,N_18582);
xor U19557 (N_19557,N_18693,N_18082);
nor U19558 (N_19558,N_18333,N_18439);
xnor U19559 (N_19559,N_18410,N_18405);
nand U19560 (N_19560,N_18946,N_18683);
xor U19561 (N_19561,N_18901,N_18938);
xor U19562 (N_19562,N_18295,N_18710);
xnor U19563 (N_19563,N_18688,N_18445);
and U19564 (N_19564,N_18940,N_18379);
xnor U19565 (N_19565,N_18883,N_18439);
nor U19566 (N_19566,N_18530,N_18522);
and U19567 (N_19567,N_18371,N_18561);
nor U19568 (N_19568,N_18570,N_18600);
nor U19569 (N_19569,N_18201,N_18958);
or U19570 (N_19570,N_18560,N_18007);
nand U19571 (N_19571,N_18314,N_18256);
xnor U19572 (N_19572,N_18121,N_18246);
nand U19573 (N_19573,N_18326,N_18824);
or U19574 (N_19574,N_18797,N_18171);
or U19575 (N_19575,N_18149,N_18786);
xor U19576 (N_19576,N_18016,N_18297);
and U19577 (N_19577,N_18006,N_18365);
nor U19578 (N_19578,N_18842,N_18595);
and U19579 (N_19579,N_18916,N_18874);
nand U19580 (N_19580,N_18839,N_18384);
or U19581 (N_19581,N_18277,N_18701);
or U19582 (N_19582,N_18466,N_18933);
or U19583 (N_19583,N_18431,N_18634);
and U19584 (N_19584,N_18690,N_18025);
or U19585 (N_19585,N_18936,N_18194);
or U19586 (N_19586,N_18183,N_18538);
nand U19587 (N_19587,N_18206,N_18680);
or U19588 (N_19588,N_18259,N_18959);
nor U19589 (N_19589,N_18256,N_18916);
xor U19590 (N_19590,N_18955,N_18858);
nand U19591 (N_19591,N_18209,N_18548);
or U19592 (N_19592,N_18343,N_18133);
and U19593 (N_19593,N_18203,N_18233);
and U19594 (N_19594,N_18872,N_18401);
xor U19595 (N_19595,N_18832,N_18810);
and U19596 (N_19596,N_18953,N_18852);
or U19597 (N_19597,N_18370,N_18566);
nand U19598 (N_19598,N_18236,N_18823);
and U19599 (N_19599,N_18928,N_18328);
nor U19600 (N_19600,N_18277,N_18311);
or U19601 (N_19601,N_18515,N_18084);
xnor U19602 (N_19602,N_18055,N_18655);
and U19603 (N_19603,N_18209,N_18124);
and U19604 (N_19604,N_18947,N_18833);
or U19605 (N_19605,N_18723,N_18760);
nor U19606 (N_19606,N_18373,N_18740);
and U19607 (N_19607,N_18784,N_18966);
nor U19608 (N_19608,N_18872,N_18961);
and U19609 (N_19609,N_18898,N_18000);
or U19610 (N_19610,N_18554,N_18798);
or U19611 (N_19611,N_18338,N_18538);
xor U19612 (N_19612,N_18316,N_18622);
xnor U19613 (N_19613,N_18705,N_18505);
or U19614 (N_19614,N_18906,N_18878);
xor U19615 (N_19615,N_18059,N_18574);
xnor U19616 (N_19616,N_18304,N_18456);
or U19617 (N_19617,N_18233,N_18028);
nor U19618 (N_19618,N_18560,N_18470);
and U19619 (N_19619,N_18579,N_18697);
nor U19620 (N_19620,N_18583,N_18029);
nor U19621 (N_19621,N_18370,N_18967);
nor U19622 (N_19622,N_18766,N_18543);
nor U19623 (N_19623,N_18881,N_18716);
nor U19624 (N_19624,N_18882,N_18849);
xnor U19625 (N_19625,N_18613,N_18434);
xor U19626 (N_19626,N_18663,N_18836);
nand U19627 (N_19627,N_18015,N_18513);
and U19628 (N_19628,N_18132,N_18686);
nand U19629 (N_19629,N_18845,N_18620);
xor U19630 (N_19630,N_18204,N_18037);
xnor U19631 (N_19631,N_18011,N_18834);
xor U19632 (N_19632,N_18542,N_18246);
or U19633 (N_19633,N_18520,N_18434);
and U19634 (N_19634,N_18745,N_18013);
and U19635 (N_19635,N_18166,N_18702);
xor U19636 (N_19636,N_18778,N_18612);
and U19637 (N_19637,N_18103,N_18424);
nand U19638 (N_19638,N_18043,N_18627);
nand U19639 (N_19639,N_18275,N_18416);
xor U19640 (N_19640,N_18144,N_18143);
nor U19641 (N_19641,N_18877,N_18928);
nand U19642 (N_19642,N_18468,N_18330);
xor U19643 (N_19643,N_18966,N_18740);
xnor U19644 (N_19644,N_18585,N_18476);
and U19645 (N_19645,N_18796,N_18491);
or U19646 (N_19646,N_18227,N_18216);
xnor U19647 (N_19647,N_18547,N_18096);
nor U19648 (N_19648,N_18196,N_18447);
and U19649 (N_19649,N_18990,N_18190);
nand U19650 (N_19650,N_18998,N_18996);
or U19651 (N_19651,N_18230,N_18382);
and U19652 (N_19652,N_18194,N_18020);
and U19653 (N_19653,N_18366,N_18464);
xor U19654 (N_19654,N_18747,N_18861);
nor U19655 (N_19655,N_18036,N_18878);
nor U19656 (N_19656,N_18128,N_18663);
nor U19657 (N_19657,N_18726,N_18274);
nand U19658 (N_19658,N_18512,N_18413);
or U19659 (N_19659,N_18044,N_18903);
xor U19660 (N_19660,N_18591,N_18415);
and U19661 (N_19661,N_18419,N_18546);
and U19662 (N_19662,N_18133,N_18557);
nand U19663 (N_19663,N_18976,N_18700);
and U19664 (N_19664,N_18266,N_18846);
nand U19665 (N_19665,N_18894,N_18676);
nand U19666 (N_19666,N_18860,N_18376);
nor U19667 (N_19667,N_18937,N_18132);
and U19668 (N_19668,N_18521,N_18564);
and U19669 (N_19669,N_18537,N_18764);
nor U19670 (N_19670,N_18884,N_18228);
nand U19671 (N_19671,N_18263,N_18325);
or U19672 (N_19672,N_18822,N_18624);
and U19673 (N_19673,N_18276,N_18711);
nor U19674 (N_19674,N_18496,N_18289);
nand U19675 (N_19675,N_18017,N_18629);
nor U19676 (N_19676,N_18313,N_18777);
and U19677 (N_19677,N_18999,N_18148);
nand U19678 (N_19678,N_18292,N_18850);
xnor U19679 (N_19679,N_18180,N_18809);
and U19680 (N_19680,N_18393,N_18745);
nand U19681 (N_19681,N_18415,N_18598);
nand U19682 (N_19682,N_18275,N_18828);
nand U19683 (N_19683,N_18299,N_18855);
nand U19684 (N_19684,N_18714,N_18206);
nand U19685 (N_19685,N_18148,N_18644);
or U19686 (N_19686,N_18878,N_18069);
and U19687 (N_19687,N_18064,N_18125);
xor U19688 (N_19688,N_18297,N_18300);
nor U19689 (N_19689,N_18324,N_18777);
xnor U19690 (N_19690,N_18520,N_18159);
or U19691 (N_19691,N_18046,N_18107);
nand U19692 (N_19692,N_18696,N_18561);
and U19693 (N_19693,N_18301,N_18418);
xnor U19694 (N_19694,N_18961,N_18016);
and U19695 (N_19695,N_18885,N_18525);
xnor U19696 (N_19696,N_18849,N_18648);
and U19697 (N_19697,N_18199,N_18803);
nand U19698 (N_19698,N_18358,N_18345);
xnor U19699 (N_19699,N_18502,N_18885);
nand U19700 (N_19700,N_18594,N_18553);
nand U19701 (N_19701,N_18744,N_18137);
and U19702 (N_19702,N_18905,N_18127);
and U19703 (N_19703,N_18743,N_18946);
and U19704 (N_19704,N_18785,N_18061);
and U19705 (N_19705,N_18035,N_18609);
nor U19706 (N_19706,N_18589,N_18377);
and U19707 (N_19707,N_18193,N_18041);
nor U19708 (N_19708,N_18545,N_18778);
xnor U19709 (N_19709,N_18002,N_18234);
nand U19710 (N_19710,N_18991,N_18313);
nor U19711 (N_19711,N_18137,N_18757);
nand U19712 (N_19712,N_18645,N_18383);
xor U19713 (N_19713,N_18780,N_18315);
and U19714 (N_19714,N_18382,N_18396);
nor U19715 (N_19715,N_18485,N_18987);
nor U19716 (N_19716,N_18148,N_18114);
xor U19717 (N_19717,N_18165,N_18442);
xor U19718 (N_19718,N_18072,N_18134);
and U19719 (N_19719,N_18591,N_18021);
xnor U19720 (N_19720,N_18330,N_18932);
nand U19721 (N_19721,N_18356,N_18704);
nand U19722 (N_19722,N_18922,N_18994);
nor U19723 (N_19723,N_18702,N_18597);
and U19724 (N_19724,N_18413,N_18601);
and U19725 (N_19725,N_18129,N_18186);
xnor U19726 (N_19726,N_18378,N_18555);
nand U19727 (N_19727,N_18922,N_18040);
and U19728 (N_19728,N_18593,N_18419);
or U19729 (N_19729,N_18599,N_18586);
nand U19730 (N_19730,N_18942,N_18689);
and U19731 (N_19731,N_18155,N_18271);
nor U19732 (N_19732,N_18966,N_18752);
and U19733 (N_19733,N_18682,N_18533);
or U19734 (N_19734,N_18884,N_18869);
and U19735 (N_19735,N_18467,N_18649);
xnor U19736 (N_19736,N_18658,N_18346);
and U19737 (N_19737,N_18252,N_18131);
or U19738 (N_19738,N_18971,N_18227);
nor U19739 (N_19739,N_18227,N_18177);
and U19740 (N_19740,N_18939,N_18499);
or U19741 (N_19741,N_18221,N_18896);
nand U19742 (N_19742,N_18558,N_18853);
or U19743 (N_19743,N_18861,N_18386);
nand U19744 (N_19744,N_18415,N_18008);
or U19745 (N_19745,N_18610,N_18086);
xnor U19746 (N_19746,N_18103,N_18446);
nor U19747 (N_19747,N_18021,N_18117);
and U19748 (N_19748,N_18602,N_18672);
and U19749 (N_19749,N_18490,N_18020);
nor U19750 (N_19750,N_18248,N_18242);
or U19751 (N_19751,N_18299,N_18094);
nand U19752 (N_19752,N_18566,N_18794);
or U19753 (N_19753,N_18542,N_18042);
nor U19754 (N_19754,N_18209,N_18121);
xnor U19755 (N_19755,N_18588,N_18187);
xnor U19756 (N_19756,N_18079,N_18658);
nand U19757 (N_19757,N_18286,N_18113);
nor U19758 (N_19758,N_18131,N_18818);
nor U19759 (N_19759,N_18565,N_18581);
nand U19760 (N_19760,N_18423,N_18628);
xnor U19761 (N_19761,N_18025,N_18770);
nor U19762 (N_19762,N_18372,N_18094);
nor U19763 (N_19763,N_18147,N_18744);
and U19764 (N_19764,N_18295,N_18762);
nand U19765 (N_19765,N_18311,N_18149);
nand U19766 (N_19766,N_18929,N_18805);
or U19767 (N_19767,N_18822,N_18471);
xor U19768 (N_19768,N_18282,N_18681);
or U19769 (N_19769,N_18657,N_18313);
nand U19770 (N_19770,N_18020,N_18236);
or U19771 (N_19771,N_18824,N_18669);
xor U19772 (N_19772,N_18828,N_18149);
nand U19773 (N_19773,N_18523,N_18059);
and U19774 (N_19774,N_18053,N_18694);
nor U19775 (N_19775,N_18401,N_18078);
xnor U19776 (N_19776,N_18509,N_18431);
nor U19777 (N_19777,N_18183,N_18270);
xor U19778 (N_19778,N_18477,N_18610);
and U19779 (N_19779,N_18961,N_18137);
xor U19780 (N_19780,N_18945,N_18108);
nor U19781 (N_19781,N_18285,N_18136);
and U19782 (N_19782,N_18345,N_18227);
and U19783 (N_19783,N_18975,N_18245);
nand U19784 (N_19784,N_18187,N_18239);
and U19785 (N_19785,N_18287,N_18873);
xor U19786 (N_19786,N_18181,N_18756);
nand U19787 (N_19787,N_18991,N_18760);
or U19788 (N_19788,N_18589,N_18528);
and U19789 (N_19789,N_18225,N_18908);
xnor U19790 (N_19790,N_18930,N_18355);
or U19791 (N_19791,N_18066,N_18508);
nand U19792 (N_19792,N_18899,N_18770);
nor U19793 (N_19793,N_18742,N_18259);
and U19794 (N_19794,N_18910,N_18540);
and U19795 (N_19795,N_18386,N_18749);
or U19796 (N_19796,N_18216,N_18321);
or U19797 (N_19797,N_18139,N_18813);
nand U19798 (N_19798,N_18854,N_18454);
and U19799 (N_19799,N_18948,N_18593);
xor U19800 (N_19800,N_18598,N_18266);
or U19801 (N_19801,N_18271,N_18451);
or U19802 (N_19802,N_18812,N_18187);
nand U19803 (N_19803,N_18738,N_18103);
xnor U19804 (N_19804,N_18822,N_18262);
or U19805 (N_19805,N_18697,N_18739);
nor U19806 (N_19806,N_18348,N_18352);
or U19807 (N_19807,N_18585,N_18867);
or U19808 (N_19808,N_18011,N_18314);
xor U19809 (N_19809,N_18399,N_18298);
nor U19810 (N_19810,N_18651,N_18773);
xor U19811 (N_19811,N_18832,N_18189);
nand U19812 (N_19812,N_18478,N_18872);
xor U19813 (N_19813,N_18607,N_18554);
nand U19814 (N_19814,N_18462,N_18153);
nor U19815 (N_19815,N_18528,N_18076);
nor U19816 (N_19816,N_18183,N_18525);
nand U19817 (N_19817,N_18537,N_18845);
or U19818 (N_19818,N_18321,N_18576);
nor U19819 (N_19819,N_18673,N_18573);
xnor U19820 (N_19820,N_18536,N_18888);
xor U19821 (N_19821,N_18510,N_18738);
nor U19822 (N_19822,N_18678,N_18858);
or U19823 (N_19823,N_18828,N_18736);
and U19824 (N_19824,N_18402,N_18063);
xnor U19825 (N_19825,N_18719,N_18455);
or U19826 (N_19826,N_18641,N_18565);
or U19827 (N_19827,N_18869,N_18909);
nand U19828 (N_19828,N_18611,N_18676);
or U19829 (N_19829,N_18645,N_18578);
nor U19830 (N_19830,N_18951,N_18470);
nand U19831 (N_19831,N_18711,N_18205);
nor U19832 (N_19832,N_18664,N_18414);
nor U19833 (N_19833,N_18606,N_18444);
and U19834 (N_19834,N_18955,N_18768);
nand U19835 (N_19835,N_18173,N_18695);
or U19836 (N_19836,N_18231,N_18350);
nand U19837 (N_19837,N_18611,N_18571);
nor U19838 (N_19838,N_18703,N_18089);
nor U19839 (N_19839,N_18369,N_18148);
nor U19840 (N_19840,N_18779,N_18904);
nor U19841 (N_19841,N_18985,N_18485);
nand U19842 (N_19842,N_18414,N_18853);
nor U19843 (N_19843,N_18072,N_18917);
or U19844 (N_19844,N_18293,N_18713);
nor U19845 (N_19845,N_18376,N_18249);
xor U19846 (N_19846,N_18584,N_18444);
or U19847 (N_19847,N_18026,N_18255);
xnor U19848 (N_19848,N_18777,N_18842);
nand U19849 (N_19849,N_18861,N_18553);
nand U19850 (N_19850,N_18553,N_18204);
or U19851 (N_19851,N_18447,N_18258);
and U19852 (N_19852,N_18031,N_18474);
nand U19853 (N_19853,N_18593,N_18549);
nand U19854 (N_19854,N_18475,N_18009);
or U19855 (N_19855,N_18013,N_18951);
and U19856 (N_19856,N_18980,N_18929);
nand U19857 (N_19857,N_18760,N_18169);
nor U19858 (N_19858,N_18354,N_18053);
and U19859 (N_19859,N_18655,N_18532);
or U19860 (N_19860,N_18889,N_18582);
nand U19861 (N_19861,N_18388,N_18185);
or U19862 (N_19862,N_18720,N_18473);
nand U19863 (N_19863,N_18106,N_18007);
and U19864 (N_19864,N_18599,N_18757);
nor U19865 (N_19865,N_18899,N_18166);
xnor U19866 (N_19866,N_18776,N_18784);
nand U19867 (N_19867,N_18137,N_18367);
nand U19868 (N_19868,N_18611,N_18386);
and U19869 (N_19869,N_18987,N_18581);
and U19870 (N_19870,N_18533,N_18197);
nand U19871 (N_19871,N_18546,N_18236);
nor U19872 (N_19872,N_18141,N_18140);
and U19873 (N_19873,N_18864,N_18448);
nor U19874 (N_19874,N_18137,N_18580);
xnor U19875 (N_19875,N_18368,N_18138);
nor U19876 (N_19876,N_18900,N_18406);
and U19877 (N_19877,N_18799,N_18454);
or U19878 (N_19878,N_18367,N_18239);
nand U19879 (N_19879,N_18319,N_18343);
xnor U19880 (N_19880,N_18917,N_18091);
xor U19881 (N_19881,N_18437,N_18112);
nor U19882 (N_19882,N_18025,N_18940);
and U19883 (N_19883,N_18345,N_18403);
nor U19884 (N_19884,N_18641,N_18542);
or U19885 (N_19885,N_18256,N_18188);
nor U19886 (N_19886,N_18637,N_18471);
nand U19887 (N_19887,N_18335,N_18728);
or U19888 (N_19888,N_18975,N_18147);
nor U19889 (N_19889,N_18913,N_18219);
nand U19890 (N_19890,N_18142,N_18442);
nand U19891 (N_19891,N_18302,N_18131);
or U19892 (N_19892,N_18901,N_18089);
and U19893 (N_19893,N_18536,N_18658);
xor U19894 (N_19894,N_18167,N_18396);
or U19895 (N_19895,N_18430,N_18001);
and U19896 (N_19896,N_18913,N_18385);
nor U19897 (N_19897,N_18146,N_18987);
and U19898 (N_19898,N_18022,N_18697);
xnor U19899 (N_19899,N_18628,N_18140);
xor U19900 (N_19900,N_18186,N_18380);
nor U19901 (N_19901,N_18877,N_18527);
xor U19902 (N_19902,N_18349,N_18154);
and U19903 (N_19903,N_18482,N_18673);
or U19904 (N_19904,N_18690,N_18188);
xor U19905 (N_19905,N_18581,N_18127);
or U19906 (N_19906,N_18412,N_18239);
nor U19907 (N_19907,N_18091,N_18180);
or U19908 (N_19908,N_18158,N_18343);
nand U19909 (N_19909,N_18520,N_18752);
xor U19910 (N_19910,N_18104,N_18827);
or U19911 (N_19911,N_18003,N_18802);
and U19912 (N_19912,N_18868,N_18215);
xnor U19913 (N_19913,N_18933,N_18448);
and U19914 (N_19914,N_18779,N_18988);
xor U19915 (N_19915,N_18233,N_18361);
nor U19916 (N_19916,N_18593,N_18925);
or U19917 (N_19917,N_18427,N_18064);
or U19918 (N_19918,N_18523,N_18708);
and U19919 (N_19919,N_18549,N_18370);
and U19920 (N_19920,N_18336,N_18547);
or U19921 (N_19921,N_18822,N_18113);
xor U19922 (N_19922,N_18456,N_18901);
nor U19923 (N_19923,N_18972,N_18175);
or U19924 (N_19924,N_18994,N_18730);
xnor U19925 (N_19925,N_18625,N_18398);
and U19926 (N_19926,N_18573,N_18204);
or U19927 (N_19927,N_18535,N_18908);
xnor U19928 (N_19928,N_18026,N_18251);
nand U19929 (N_19929,N_18527,N_18935);
nor U19930 (N_19930,N_18563,N_18763);
xnor U19931 (N_19931,N_18961,N_18723);
xnor U19932 (N_19932,N_18704,N_18880);
nand U19933 (N_19933,N_18365,N_18620);
or U19934 (N_19934,N_18194,N_18351);
xor U19935 (N_19935,N_18378,N_18818);
and U19936 (N_19936,N_18255,N_18673);
nand U19937 (N_19937,N_18040,N_18941);
or U19938 (N_19938,N_18688,N_18464);
or U19939 (N_19939,N_18273,N_18172);
xnor U19940 (N_19940,N_18249,N_18100);
and U19941 (N_19941,N_18645,N_18947);
or U19942 (N_19942,N_18993,N_18426);
and U19943 (N_19943,N_18321,N_18855);
nand U19944 (N_19944,N_18656,N_18248);
and U19945 (N_19945,N_18936,N_18233);
xor U19946 (N_19946,N_18656,N_18310);
xnor U19947 (N_19947,N_18529,N_18371);
or U19948 (N_19948,N_18630,N_18235);
and U19949 (N_19949,N_18285,N_18535);
nor U19950 (N_19950,N_18220,N_18541);
or U19951 (N_19951,N_18264,N_18555);
and U19952 (N_19952,N_18016,N_18534);
nor U19953 (N_19953,N_18179,N_18393);
nand U19954 (N_19954,N_18872,N_18935);
and U19955 (N_19955,N_18922,N_18722);
xor U19956 (N_19956,N_18199,N_18669);
and U19957 (N_19957,N_18041,N_18363);
or U19958 (N_19958,N_18587,N_18390);
or U19959 (N_19959,N_18104,N_18814);
nand U19960 (N_19960,N_18317,N_18046);
nor U19961 (N_19961,N_18395,N_18607);
or U19962 (N_19962,N_18484,N_18354);
nand U19963 (N_19963,N_18153,N_18106);
or U19964 (N_19964,N_18877,N_18312);
xnor U19965 (N_19965,N_18929,N_18233);
and U19966 (N_19966,N_18208,N_18080);
or U19967 (N_19967,N_18370,N_18851);
or U19968 (N_19968,N_18159,N_18229);
xor U19969 (N_19969,N_18337,N_18915);
and U19970 (N_19970,N_18155,N_18781);
and U19971 (N_19971,N_18060,N_18099);
nor U19972 (N_19972,N_18914,N_18828);
and U19973 (N_19973,N_18288,N_18413);
nand U19974 (N_19974,N_18226,N_18583);
and U19975 (N_19975,N_18981,N_18211);
xor U19976 (N_19976,N_18977,N_18353);
or U19977 (N_19977,N_18514,N_18785);
and U19978 (N_19978,N_18755,N_18067);
and U19979 (N_19979,N_18026,N_18926);
xor U19980 (N_19980,N_18048,N_18835);
or U19981 (N_19981,N_18120,N_18538);
xnor U19982 (N_19982,N_18101,N_18710);
and U19983 (N_19983,N_18788,N_18896);
nor U19984 (N_19984,N_18832,N_18503);
nand U19985 (N_19985,N_18055,N_18947);
nor U19986 (N_19986,N_18232,N_18218);
nor U19987 (N_19987,N_18895,N_18934);
nor U19988 (N_19988,N_18713,N_18346);
and U19989 (N_19989,N_18213,N_18711);
nor U19990 (N_19990,N_18390,N_18469);
and U19991 (N_19991,N_18812,N_18456);
xor U19992 (N_19992,N_18525,N_18642);
nand U19993 (N_19993,N_18780,N_18779);
or U19994 (N_19994,N_18637,N_18212);
xnor U19995 (N_19995,N_18070,N_18833);
nor U19996 (N_19996,N_18123,N_18443);
and U19997 (N_19997,N_18949,N_18636);
xnor U19998 (N_19998,N_18415,N_18778);
xor U19999 (N_19999,N_18540,N_18442);
nor U20000 (N_20000,N_19386,N_19622);
xor U20001 (N_20001,N_19178,N_19542);
and U20002 (N_20002,N_19826,N_19526);
nor U20003 (N_20003,N_19568,N_19229);
xnor U20004 (N_20004,N_19165,N_19806);
nand U20005 (N_20005,N_19121,N_19192);
xor U20006 (N_20006,N_19434,N_19637);
or U20007 (N_20007,N_19939,N_19673);
nand U20008 (N_20008,N_19864,N_19799);
or U20009 (N_20009,N_19522,N_19848);
nor U20010 (N_20010,N_19881,N_19527);
nor U20011 (N_20011,N_19075,N_19055);
nand U20012 (N_20012,N_19683,N_19795);
xnor U20013 (N_20013,N_19454,N_19796);
nand U20014 (N_20014,N_19014,N_19923);
xor U20015 (N_20015,N_19747,N_19624);
nor U20016 (N_20016,N_19094,N_19347);
xnor U20017 (N_20017,N_19890,N_19515);
xnor U20018 (N_20018,N_19834,N_19874);
xor U20019 (N_20019,N_19538,N_19373);
nand U20020 (N_20020,N_19761,N_19958);
and U20021 (N_20021,N_19493,N_19584);
nor U20022 (N_20022,N_19311,N_19812);
nor U20023 (N_20023,N_19539,N_19644);
nor U20024 (N_20024,N_19452,N_19701);
xnor U20025 (N_20025,N_19294,N_19798);
or U20026 (N_20026,N_19019,N_19955);
xor U20027 (N_20027,N_19163,N_19477);
xnor U20028 (N_20028,N_19088,N_19141);
and U20029 (N_20029,N_19885,N_19704);
and U20030 (N_20030,N_19700,N_19167);
or U20031 (N_20031,N_19720,N_19916);
xor U20032 (N_20032,N_19763,N_19419);
xor U20033 (N_20033,N_19020,N_19979);
nand U20034 (N_20034,N_19004,N_19145);
or U20035 (N_20035,N_19389,N_19310);
nor U20036 (N_20036,N_19387,N_19569);
nand U20037 (N_20037,N_19820,N_19684);
and U20038 (N_20038,N_19614,N_19651);
and U20039 (N_20039,N_19572,N_19974);
and U20040 (N_20040,N_19366,N_19458);
or U20041 (N_20041,N_19697,N_19549);
nor U20042 (N_20042,N_19717,N_19532);
xor U20043 (N_20043,N_19368,N_19432);
nor U20044 (N_20044,N_19585,N_19575);
nor U20045 (N_20045,N_19792,N_19730);
nor U20046 (N_20046,N_19833,N_19374);
or U20047 (N_20047,N_19171,N_19241);
and U20048 (N_20048,N_19453,N_19956);
or U20049 (N_20049,N_19027,N_19408);
and U20050 (N_20050,N_19922,N_19361);
or U20051 (N_20051,N_19587,N_19272);
xnor U20052 (N_20052,N_19971,N_19814);
and U20053 (N_20053,N_19010,N_19647);
xor U20054 (N_20054,N_19774,N_19384);
nor U20055 (N_20055,N_19724,N_19096);
xor U20056 (N_20056,N_19865,N_19540);
nand U20057 (N_20057,N_19355,N_19503);
xnor U20058 (N_20058,N_19816,N_19337);
and U20059 (N_20059,N_19136,N_19559);
xor U20060 (N_20060,N_19489,N_19589);
xnor U20061 (N_20061,N_19506,N_19359);
or U20062 (N_20062,N_19160,N_19153);
or U20063 (N_20063,N_19997,N_19467);
nor U20064 (N_20064,N_19079,N_19068);
nand U20065 (N_20065,N_19067,N_19742);
nor U20066 (N_20066,N_19581,N_19312);
nor U20067 (N_20067,N_19764,N_19656);
xnor U20068 (N_20068,N_19660,N_19738);
and U20069 (N_20069,N_19775,N_19450);
xnor U20070 (N_20070,N_19256,N_19557);
nor U20071 (N_20071,N_19334,N_19894);
xnor U20072 (N_20072,N_19106,N_19155);
xor U20073 (N_20073,N_19957,N_19169);
or U20074 (N_20074,N_19586,N_19054);
nand U20075 (N_20075,N_19904,N_19174);
nand U20076 (N_20076,N_19983,N_19843);
xnor U20077 (N_20077,N_19635,N_19433);
and U20078 (N_20078,N_19789,N_19487);
or U20079 (N_20079,N_19238,N_19950);
and U20080 (N_20080,N_19024,N_19367);
and U20081 (N_20081,N_19222,N_19070);
nand U20082 (N_20082,N_19511,N_19606);
xnor U20083 (N_20083,N_19759,N_19550);
xnor U20084 (N_20084,N_19715,N_19228);
or U20085 (N_20085,N_19329,N_19492);
and U20086 (N_20086,N_19046,N_19401);
and U20087 (N_20087,N_19811,N_19154);
xnor U20088 (N_20088,N_19109,N_19849);
nor U20089 (N_20089,N_19645,N_19803);
or U20090 (N_20090,N_19464,N_19360);
nand U20091 (N_20091,N_19444,N_19854);
nor U20092 (N_20092,N_19250,N_19605);
or U20093 (N_20093,N_19535,N_19425);
nand U20094 (N_20094,N_19966,N_19986);
nand U20095 (N_20095,N_19852,N_19164);
and U20096 (N_20096,N_19883,N_19502);
xor U20097 (N_20097,N_19262,N_19188);
and U20098 (N_20098,N_19151,N_19322);
and U20099 (N_20099,N_19889,N_19828);
or U20100 (N_20100,N_19092,N_19264);
xor U20101 (N_20101,N_19420,N_19223);
or U20102 (N_20102,N_19655,N_19343);
nand U20103 (N_20103,N_19767,N_19779);
xnor U20104 (N_20104,N_19518,N_19085);
or U20105 (N_20105,N_19421,N_19847);
xor U20106 (N_20106,N_19607,N_19975);
nand U20107 (N_20107,N_19059,N_19516);
xnor U20108 (N_20108,N_19571,N_19807);
or U20109 (N_20109,N_19486,N_19842);
nor U20110 (N_20110,N_19582,N_19591);
and U20111 (N_20111,N_19306,N_19261);
or U20112 (N_20112,N_19166,N_19388);
xor U20113 (N_20113,N_19888,N_19623);
and U20114 (N_20114,N_19157,N_19415);
or U20115 (N_20115,N_19325,N_19275);
and U20116 (N_20116,N_19824,N_19056);
and U20117 (N_20117,N_19112,N_19081);
xor U20118 (N_20118,N_19615,N_19616);
or U20119 (N_20119,N_19898,N_19414);
or U20120 (N_20120,N_19937,N_19265);
nand U20121 (N_20121,N_19128,N_19926);
nor U20122 (N_20122,N_19702,N_19047);
nand U20123 (N_20123,N_19267,N_19077);
and U20124 (N_20124,N_19841,N_19760);
xor U20125 (N_20125,N_19741,N_19175);
and U20126 (N_20126,N_19138,N_19321);
xor U20127 (N_20127,N_19039,N_19028);
xor U20128 (N_20128,N_19711,N_19208);
or U20129 (N_20129,N_19314,N_19235);
nand U20130 (N_20130,N_19765,N_19696);
and U20131 (N_20131,N_19447,N_19289);
xnor U20132 (N_20132,N_19441,N_19773);
xnor U20133 (N_20133,N_19925,N_19122);
nand U20134 (N_20134,N_19546,N_19993);
and U20135 (N_20135,N_19198,N_19206);
nor U20136 (N_20136,N_19282,N_19844);
or U20137 (N_20137,N_19439,N_19135);
nand U20138 (N_20138,N_19992,N_19876);
xnor U20139 (N_20139,N_19687,N_19427);
or U20140 (N_20140,N_19065,N_19544);
nor U20141 (N_20141,N_19234,N_19195);
nand U20142 (N_20142,N_19423,N_19574);
nand U20143 (N_20143,N_19269,N_19335);
or U20144 (N_20144,N_19001,N_19132);
nor U20145 (N_20145,N_19479,N_19147);
xor U20146 (N_20146,N_19686,N_19525);
and U20147 (N_20147,N_19497,N_19358);
xnor U20148 (N_20148,N_19236,N_19921);
and U20149 (N_20149,N_19541,N_19665);
or U20150 (N_20150,N_19281,N_19612);
and U20151 (N_20151,N_19588,N_19209);
xor U20152 (N_20152,N_19891,N_19125);
or U20153 (N_20153,N_19573,N_19168);
xnor U20154 (N_20154,N_19719,N_19110);
nand U20155 (N_20155,N_19514,N_19910);
or U20156 (N_20156,N_19033,N_19899);
and U20157 (N_20157,N_19652,N_19064);
xor U20158 (N_20158,N_19330,N_19076);
xor U20159 (N_20159,N_19363,N_19815);
nor U20160 (N_20160,N_19397,N_19357);
and U20161 (N_20161,N_19045,N_19158);
nand U20162 (N_20162,N_19661,N_19703);
or U20163 (N_20163,N_19181,N_19346);
and U20164 (N_20164,N_19246,N_19405);
nand U20165 (N_20165,N_19838,N_19602);
or U20166 (N_20166,N_19317,N_19817);
xor U20167 (N_20167,N_19823,N_19618);
xor U20168 (N_20168,N_19193,N_19431);
and U20169 (N_20169,N_19049,N_19553);
xor U20170 (N_20170,N_19633,N_19886);
and U20171 (N_20171,N_19219,N_19286);
xnor U20172 (N_20172,N_19469,N_19103);
or U20173 (N_20173,N_19291,N_19907);
xnor U20174 (N_20174,N_19689,N_19669);
xor U20175 (N_20175,N_19555,N_19259);
nor U20176 (N_20176,N_19710,N_19478);
nand U20177 (N_20177,N_19830,N_19919);
nor U20178 (N_20178,N_19908,N_19170);
nor U20179 (N_20179,N_19436,N_19914);
nor U20180 (N_20180,N_19935,N_19255);
nor U20181 (N_20181,N_19215,N_19508);
nand U20182 (N_20182,N_19396,N_19271);
xor U20183 (N_20183,N_19105,N_19426);
nor U20184 (N_20184,N_19475,N_19101);
nand U20185 (N_20185,N_19999,N_19877);
xnor U20186 (N_20186,N_19802,N_19107);
nand U20187 (N_20187,N_19768,N_19007);
xnor U20188 (N_20188,N_19179,N_19733);
nand U20189 (N_20189,N_19845,N_19734);
nand U20190 (N_20190,N_19777,N_19912);
and U20191 (N_20191,N_19032,N_19752);
or U20192 (N_20192,N_19012,N_19731);
or U20193 (N_20193,N_19531,N_19352);
xnor U20194 (N_20194,N_19998,N_19184);
and U20195 (N_20195,N_19579,N_19629);
or U20196 (N_20196,N_19987,N_19932);
nand U20197 (N_20197,N_19643,N_19859);
nand U20198 (N_20198,N_19491,N_19091);
or U20199 (N_20199,N_19757,N_19082);
or U20200 (N_20200,N_19592,N_19943);
and U20201 (N_20201,N_19976,N_19340);
nor U20202 (N_20202,N_19245,N_19481);
xor U20203 (N_20203,N_19520,N_19430);
or U20204 (N_20204,N_19762,N_19496);
nor U20205 (N_20205,N_19356,N_19626);
or U20206 (N_20206,N_19878,N_19484);
or U20207 (N_20207,N_19946,N_19459);
nand U20208 (N_20208,N_19945,N_19089);
or U20209 (N_20209,N_19625,N_19131);
nand U20210 (N_20210,N_19350,N_19949);
nor U20211 (N_20211,N_19378,N_19861);
nand U20212 (N_20212,N_19455,N_19102);
nor U20213 (N_20213,N_19097,N_19872);
xnor U20214 (N_20214,N_19302,N_19688);
and U20215 (N_20215,N_19456,N_19810);
xnor U20216 (N_20216,N_19124,N_19410);
and U20217 (N_20217,N_19940,N_19021);
or U20218 (N_20218,N_19982,N_19737);
xor U20219 (N_20219,N_19393,N_19226);
xor U20220 (N_20220,N_19276,N_19536);
and U20221 (N_20221,N_19977,N_19036);
nor U20222 (N_20222,N_19610,N_19349);
and U20223 (N_20223,N_19895,N_19778);
xor U20224 (N_20224,N_19855,N_19692);
and U20225 (N_20225,N_19951,N_19658);
xnor U20226 (N_20226,N_19679,N_19353);
nand U20227 (N_20227,N_19280,N_19451);
nor U20228 (N_20228,N_19634,N_19190);
and U20229 (N_20229,N_19108,N_19394);
and U20230 (N_20230,N_19090,N_19504);
or U20231 (N_20231,N_19879,N_19413);
or U20232 (N_20232,N_19776,N_19718);
or U20233 (N_20233,N_19461,N_19002);
and U20234 (N_20234,N_19237,N_19490);
xnor U20235 (N_20235,N_19784,N_19560);
nor U20236 (N_20236,N_19695,N_19954);
xnor U20237 (N_20237,N_19244,N_19025);
and U20238 (N_20238,N_19331,N_19488);
nor U20239 (N_20239,N_19893,N_19037);
nand U20240 (N_20240,N_19130,N_19978);
and U20241 (N_20241,N_19911,N_19274);
or U20242 (N_20242,N_19266,N_19632);
nand U20243 (N_20243,N_19476,N_19827);
nor U20244 (N_20244,N_19008,N_19751);
xor U20245 (N_20245,N_19172,N_19822);
nor U20246 (N_20246,N_19220,N_19973);
nor U20247 (N_20247,N_19189,N_19918);
and U20248 (N_20248,N_19463,N_19985);
or U20249 (N_20249,N_19023,N_19562);
nand U20250 (N_20250,N_19084,N_19788);
or U20251 (N_20251,N_19071,N_19224);
xnor U20252 (N_20252,N_19248,N_19214);
xnor U20253 (N_20253,N_19176,N_19725);
nand U20254 (N_20254,N_19797,N_19466);
or U20255 (N_20255,N_19551,N_19369);
and U20256 (N_20256,N_19654,N_19407);
nor U20257 (N_20257,N_19137,N_19676);
xor U20258 (N_20258,N_19595,N_19293);
xnor U20259 (N_20259,N_19204,N_19866);
xnor U20260 (N_20260,N_19364,N_19308);
xnor U20261 (N_20261,N_19853,N_19257);
and U20262 (N_20262,N_19743,N_19500);
or U20263 (N_20263,N_19341,N_19249);
nand U20264 (N_20264,N_19446,N_19197);
and U20265 (N_20265,N_19996,N_19869);
nor U20266 (N_20266,N_19967,N_19095);
nand U20267 (N_20267,N_19561,N_19111);
and U20268 (N_20268,N_19263,N_19545);
and U20269 (N_20269,N_19548,N_19682);
nand U20270 (N_20270,N_19416,N_19667);
or U20271 (N_20271,N_19113,N_19013);
nor U20272 (N_20272,N_19287,N_19638);
nand U20273 (N_20273,N_19969,N_19846);
xor U20274 (N_20274,N_19348,N_19242);
and U20275 (N_20275,N_19793,N_19860);
xor U20276 (N_20276,N_19944,N_19370);
xnor U20277 (N_20277,N_19603,N_19554);
nor U20278 (N_20278,N_19058,N_19417);
nor U20279 (N_20279,N_19318,N_19230);
or U20280 (N_20280,N_19690,N_19604);
nand U20281 (N_20281,N_19297,N_19781);
nand U20282 (N_20282,N_19061,N_19116);
and U20283 (N_20283,N_19512,N_19173);
nand U20284 (N_20284,N_19800,N_19597);
and U20285 (N_20285,N_19722,N_19565);
xor U20286 (N_20286,N_19677,N_19713);
nand U20287 (N_20287,N_19593,N_19323);
and U20288 (N_20288,N_19161,N_19791);
nand U20289 (N_20289,N_19099,N_19611);
or U20290 (N_20290,N_19344,N_19460);
and U20291 (N_20291,N_19933,N_19284);
nand U20292 (N_20292,N_19309,N_19529);
xor U20293 (N_20293,N_19143,N_19411);
and U20294 (N_20294,N_19285,N_19739);
nand U20295 (N_20295,N_19941,N_19851);
nand U20296 (N_20296,N_19041,N_19558);
nand U20297 (N_20297,N_19495,N_19523);
nor U20298 (N_20298,N_19474,N_19884);
nor U20299 (N_20299,N_19114,N_19783);
and U20300 (N_20300,N_19863,N_19207);
nand U20301 (N_20301,N_19896,N_19786);
or U20302 (N_20302,N_19485,N_19505);
nor U20303 (N_20303,N_19972,N_19498);
and U20304 (N_20304,N_19887,N_19753);
or U20305 (N_20305,N_19148,N_19104);
xor U20306 (N_20306,N_19552,N_19543);
or U20307 (N_20307,N_19707,N_19399);
and U20308 (N_20308,N_19670,N_19300);
nor U20309 (N_20309,N_19354,N_19243);
nor U20310 (N_20310,N_19857,N_19875);
nand U20311 (N_20311,N_19794,N_19578);
xnor U20312 (N_20312,N_19005,N_19048);
nand U20313 (N_20313,N_19156,N_19936);
xnor U20314 (N_20314,N_19011,N_19438);
xor U20315 (N_20315,N_19333,N_19712);
nand U20316 (N_20316,N_19319,N_19913);
nor U20317 (N_20317,N_19398,N_19429);
or U20318 (N_20318,N_19424,N_19534);
nand U20319 (N_20319,N_19442,N_19903);
xor U20320 (N_20320,N_19115,N_19959);
nand U20321 (N_20321,N_19517,N_19640);
nor U20322 (N_20322,N_19462,N_19406);
nand U20323 (N_20323,N_19342,N_19970);
and U20324 (N_20324,N_19570,N_19443);
or U20325 (N_20325,N_19862,N_19187);
nor U20326 (N_20326,N_19301,N_19034);
xnor U20327 (N_20327,N_19721,N_19043);
xnor U20328 (N_20328,N_19726,N_19307);
and U20329 (N_20329,N_19596,N_19418);
nor U20330 (N_20330,N_19251,N_19126);
or U20331 (N_20331,N_19252,N_19038);
nand U20332 (N_20332,N_19196,N_19227);
or U20333 (N_20333,N_19290,N_19057);
nand U20334 (N_20334,N_19052,N_19239);
nor U20335 (N_20335,N_19808,N_19375);
and U20336 (N_20336,N_19445,N_19305);
nand U20337 (N_20337,N_19989,N_19362);
or U20338 (N_20338,N_19772,N_19729);
and U20339 (N_20339,N_19609,N_19785);
nand U20340 (N_20340,N_19093,N_19631);
or U20341 (N_20341,N_19339,N_19769);
xor U20342 (N_20342,N_19328,N_19755);
or U20343 (N_20343,N_19233,N_19580);
nand U20344 (N_20344,N_19031,N_19299);
xor U20345 (N_20345,N_19938,N_19758);
nor U20346 (N_20346,N_19062,N_19288);
and U20347 (N_20347,N_19390,N_19766);
xor U20348 (N_20348,N_19867,N_19017);
and U20349 (N_20349,N_19296,N_19240);
and U20350 (N_20350,N_19650,N_19980);
or U20351 (N_20351,N_19199,N_19030);
nor U20352 (N_20352,N_19412,N_19620);
and U20353 (N_20353,N_19152,N_19901);
nand U20354 (N_20354,N_19920,N_19134);
nor U20355 (N_20355,N_19371,N_19142);
xor U20356 (N_20356,N_19457,N_19471);
or U20357 (N_20357,N_19313,N_19519);
nor U20358 (N_20358,N_19952,N_19391);
xnor U20359 (N_20359,N_19801,N_19927);
xnor U20360 (N_20360,N_19599,N_19917);
nand U20361 (N_20361,N_19825,N_19277);
nor U20362 (N_20362,N_19210,N_19501);
or U20363 (N_20363,N_19608,N_19381);
nor U20364 (N_20364,N_19962,N_19931);
or U20365 (N_20365,N_19900,N_19440);
nand U20366 (N_20366,N_19392,N_19351);
nand U20367 (N_20367,N_19377,N_19934);
nand U20368 (N_20368,N_19016,N_19691);
xnor U20369 (N_20369,N_19947,N_19448);
nor U20370 (N_20370,N_19693,N_19871);
nand U20371 (N_20371,N_19991,N_19182);
nand U20372 (N_20372,N_19694,N_19217);
nor U20373 (N_20373,N_19409,N_19988);
or U20374 (N_20374,N_19530,N_19636);
nor U20375 (N_20375,N_19735,N_19402);
xnor U20376 (N_20376,N_19080,N_19732);
or U20377 (N_20377,N_19345,N_19205);
xnor U20378 (N_20378,N_19681,N_19746);
nor U20379 (N_20379,N_19483,N_19221);
xnor U20380 (N_20380,N_19663,N_19678);
or U20381 (N_20381,N_19521,N_19225);
nor U20382 (N_20382,N_19231,N_19327);
and U20383 (N_20383,N_19211,N_19180);
or U20384 (N_20384,N_19577,N_19022);
or U20385 (N_20385,N_19664,N_19659);
and U20386 (N_20386,N_19837,N_19074);
nor U20387 (N_20387,N_19494,N_19365);
nor U20388 (N_20388,N_19547,N_19063);
xor U20389 (N_20389,N_19098,N_19123);
nand U20390 (N_20390,N_19805,N_19050);
nand U20391 (N_20391,N_19648,N_19379);
xnor U20392 (N_20392,N_19600,N_19716);
xnor U20393 (N_20393,N_19882,N_19736);
nand U20394 (N_20394,N_19771,N_19902);
xor U20395 (N_20395,N_19965,N_19006);
xnor U20396 (N_20396,N_19437,N_19254);
nand U20397 (N_20397,N_19268,N_19086);
xor U20398 (N_20398,N_19470,N_19000);
nor U20399 (N_20399,N_19556,N_19200);
nor U20400 (N_20400,N_19953,N_19782);
and U20401 (N_20401,N_19909,N_19203);
or U20402 (N_20402,N_19380,N_19995);
xor U20403 (N_20403,N_19332,N_19942);
xor U20404 (N_20404,N_19133,N_19566);
nor U20405 (N_20405,N_19315,N_19928);
and U20406 (N_20406,N_19303,N_19699);
nand U20407 (N_20407,N_19621,N_19706);
xor U20408 (N_20408,N_19260,N_19856);
nand U20409 (N_20409,N_19750,N_19078);
and U20410 (N_20410,N_19748,N_19641);
xor U20411 (N_20411,N_19594,N_19044);
nor U20412 (N_20412,N_19279,N_19482);
and U20413 (N_20413,N_19619,N_19672);
and U20414 (N_20414,N_19723,N_19385);
and U20415 (N_20415,N_19499,N_19120);
nand U20416 (N_20416,N_19709,N_19924);
or U20417 (N_20417,N_19666,N_19868);
nor U20418 (N_20418,N_19821,N_19029);
nor U20419 (N_20419,N_19372,N_19507);
nor U20420 (N_20420,N_19326,N_19510);
or U20421 (N_20421,N_19382,N_19671);
or U20422 (N_20422,N_19149,N_19292);
or U20423 (N_20423,N_19528,N_19298);
xor U20424 (N_20424,N_19770,N_19858);
xor U20425 (N_20425,N_19336,N_19929);
nor U20426 (N_20426,N_19087,N_19185);
or U20427 (N_20427,N_19590,N_19533);
nor U20428 (N_20428,N_19480,N_19583);
nand U20429 (N_20429,N_19316,N_19472);
xnor U20430 (N_20430,N_19627,N_19674);
nand U20431 (N_20431,N_19278,N_19146);
xor U20432 (N_20432,N_19740,N_19513);
xnor U20433 (N_20433,N_19015,N_19119);
nor U20434 (N_20434,N_19617,N_19435);
or U20435 (N_20435,N_19127,N_19283);
xnor U20436 (N_20436,N_19873,N_19051);
nor U20437 (N_20437,N_19839,N_19930);
or U20438 (N_20438,N_19780,N_19657);
nand U20439 (N_20439,N_19026,N_19850);
nor U20440 (N_20440,N_19727,N_19749);
and U20441 (N_20441,N_19139,N_19646);
nand U20442 (N_20442,N_19790,N_19129);
nor U20443 (N_20443,N_19567,N_19018);
or U20444 (N_20444,N_19668,N_19509);
and U20445 (N_20445,N_19338,N_19073);
nand U20446 (N_20446,N_19201,N_19639);
and U20447 (N_20447,N_19598,N_19270);
and U20448 (N_20448,N_19675,N_19897);
nor U20449 (N_20449,N_19072,N_19613);
nor U20450 (N_20450,N_19981,N_19804);
and U20451 (N_20451,N_19449,N_19662);
xnor U20452 (N_20452,N_19060,N_19144);
nand U20453 (N_20453,N_19009,N_19628);
nand U20454 (N_20454,N_19832,N_19320);
or U20455 (N_20455,N_19601,N_19653);
or U20456 (N_20456,N_19906,N_19159);
or U20457 (N_20457,N_19100,N_19213);
or U20458 (N_20458,N_19003,N_19984);
xor U20459 (N_20459,N_19880,N_19216);
nor U20460 (N_20460,N_19150,N_19870);
nor U20461 (N_20461,N_19035,N_19708);
nor U20462 (N_20462,N_19705,N_19642);
xor U20463 (N_20463,N_19040,N_19756);
nand U20464 (N_20464,N_19422,N_19787);
nor U20465 (N_20465,N_19232,N_19468);
nor U20466 (N_20466,N_19813,N_19273);
xor U20467 (N_20467,N_19819,N_19376);
or U20468 (N_20468,N_19186,N_19698);
xor U20469 (N_20469,N_19994,N_19714);
nand U20470 (N_20470,N_19576,N_19258);
nand U20471 (N_20471,N_19162,N_19053);
xor U20472 (N_20472,N_19836,N_19754);
xnor U20473 (N_20473,N_19960,N_19042);
nor U20474 (N_20474,N_19465,N_19963);
xnor U20475 (N_20475,N_19630,N_19745);
or U20476 (N_20476,N_19829,N_19247);
nand U20477 (N_20477,N_19403,N_19191);
xor U20478 (N_20478,N_19649,N_19905);
and U20479 (N_20479,N_19948,N_19680);
or U20480 (N_20480,N_19961,N_19183);
and U20481 (N_20481,N_19066,N_19383);
xnor U20482 (N_20482,N_19964,N_19395);
nor U20483 (N_20483,N_19473,N_19744);
xnor U20484 (N_20484,N_19563,N_19892);
and U20485 (N_20485,N_19140,N_19295);
nand U20486 (N_20486,N_19537,N_19835);
nor U20487 (N_20487,N_19118,N_19524);
nor U20488 (N_20488,N_19117,N_19069);
or U20489 (N_20489,N_19968,N_19915);
and U20490 (N_20490,N_19324,N_19400);
and U20491 (N_20491,N_19428,N_19194);
or U20492 (N_20492,N_19728,N_19404);
nor U20493 (N_20493,N_19218,N_19990);
xnor U20494 (N_20494,N_19304,N_19685);
nor U20495 (N_20495,N_19564,N_19818);
xnor U20496 (N_20496,N_19177,N_19212);
or U20497 (N_20497,N_19831,N_19253);
nor U20498 (N_20498,N_19809,N_19083);
nand U20499 (N_20499,N_19202,N_19840);
nor U20500 (N_20500,N_19567,N_19829);
and U20501 (N_20501,N_19292,N_19864);
xnor U20502 (N_20502,N_19066,N_19878);
or U20503 (N_20503,N_19668,N_19940);
or U20504 (N_20504,N_19137,N_19850);
nor U20505 (N_20505,N_19441,N_19421);
or U20506 (N_20506,N_19219,N_19883);
nor U20507 (N_20507,N_19681,N_19503);
xnor U20508 (N_20508,N_19517,N_19692);
and U20509 (N_20509,N_19273,N_19626);
nor U20510 (N_20510,N_19943,N_19330);
nand U20511 (N_20511,N_19215,N_19864);
nand U20512 (N_20512,N_19862,N_19541);
or U20513 (N_20513,N_19334,N_19313);
nand U20514 (N_20514,N_19149,N_19761);
nand U20515 (N_20515,N_19246,N_19863);
or U20516 (N_20516,N_19167,N_19035);
or U20517 (N_20517,N_19097,N_19963);
nor U20518 (N_20518,N_19609,N_19483);
nor U20519 (N_20519,N_19887,N_19990);
or U20520 (N_20520,N_19740,N_19504);
xor U20521 (N_20521,N_19357,N_19083);
and U20522 (N_20522,N_19656,N_19729);
nor U20523 (N_20523,N_19849,N_19429);
and U20524 (N_20524,N_19239,N_19250);
xnor U20525 (N_20525,N_19952,N_19898);
nor U20526 (N_20526,N_19982,N_19182);
nand U20527 (N_20527,N_19197,N_19582);
nand U20528 (N_20528,N_19613,N_19905);
and U20529 (N_20529,N_19331,N_19685);
nor U20530 (N_20530,N_19580,N_19577);
or U20531 (N_20531,N_19535,N_19716);
xor U20532 (N_20532,N_19648,N_19220);
or U20533 (N_20533,N_19188,N_19756);
xnor U20534 (N_20534,N_19463,N_19129);
xnor U20535 (N_20535,N_19927,N_19840);
and U20536 (N_20536,N_19039,N_19993);
or U20537 (N_20537,N_19744,N_19404);
or U20538 (N_20538,N_19336,N_19848);
or U20539 (N_20539,N_19113,N_19730);
xor U20540 (N_20540,N_19308,N_19560);
nand U20541 (N_20541,N_19718,N_19495);
nand U20542 (N_20542,N_19577,N_19209);
nor U20543 (N_20543,N_19188,N_19192);
nand U20544 (N_20544,N_19416,N_19214);
and U20545 (N_20545,N_19386,N_19028);
nor U20546 (N_20546,N_19182,N_19799);
xor U20547 (N_20547,N_19346,N_19531);
xor U20548 (N_20548,N_19165,N_19905);
nor U20549 (N_20549,N_19613,N_19878);
nor U20550 (N_20550,N_19325,N_19340);
and U20551 (N_20551,N_19702,N_19715);
xnor U20552 (N_20552,N_19437,N_19432);
and U20553 (N_20553,N_19335,N_19087);
nand U20554 (N_20554,N_19064,N_19015);
and U20555 (N_20555,N_19713,N_19400);
and U20556 (N_20556,N_19000,N_19903);
nor U20557 (N_20557,N_19321,N_19910);
nor U20558 (N_20558,N_19669,N_19857);
nand U20559 (N_20559,N_19220,N_19632);
xnor U20560 (N_20560,N_19360,N_19714);
nor U20561 (N_20561,N_19928,N_19974);
xnor U20562 (N_20562,N_19737,N_19588);
nor U20563 (N_20563,N_19889,N_19905);
xnor U20564 (N_20564,N_19443,N_19161);
nand U20565 (N_20565,N_19540,N_19442);
and U20566 (N_20566,N_19951,N_19597);
and U20567 (N_20567,N_19427,N_19907);
xor U20568 (N_20568,N_19514,N_19855);
xnor U20569 (N_20569,N_19394,N_19581);
nand U20570 (N_20570,N_19644,N_19054);
nor U20571 (N_20571,N_19205,N_19853);
xor U20572 (N_20572,N_19099,N_19177);
nand U20573 (N_20573,N_19280,N_19875);
or U20574 (N_20574,N_19888,N_19569);
or U20575 (N_20575,N_19433,N_19655);
nand U20576 (N_20576,N_19371,N_19033);
nand U20577 (N_20577,N_19590,N_19901);
and U20578 (N_20578,N_19806,N_19138);
nor U20579 (N_20579,N_19002,N_19075);
nor U20580 (N_20580,N_19297,N_19992);
or U20581 (N_20581,N_19190,N_19060);
and U20582 (N_20582,N_19286,N_19007);
nor U20583 (N_20583,N_19721,N_19871);
nor U20584 (N_20584,N_19975,N_19140);
nor U20585 (N_20585,N_19651,N_19667);
and U20586 (N_20586,N_19003,N_19945);
xor U20587 (N_20587,N_19035,N_19592);
xor U20588 (N_20588,N_19565,N_19454);
xnor U20589 (N_20589,N_19754,N_19742);
or U20590 (N_20590,N_19883,N_19460);
or U20591 (N_20591,N_19473,N_19372);
xor U20592 (N_20592,N_19708,N_19469);
nor U20593 (N_20593,N_19717,N_19250);
xnor U20594 (N_20594,N_19523,N_19831);
nand U20595 (N_20595,N_19051,N_19675);
nand U20596 (N_20596,N_19677,N_19735);
nor U20597 (N_20597,N_19353,N_19699);
or U20598 (N_20598,N_19768,N_19401);
or U20599 (N_20599,N_19038,N_19926);
or U20600 (N_20600,N_19286,N_19953);
and U20601 (N_20601,N_19318,N_19583);
nor U20602 (N_20602,N_19806,N_19399);
xor U20603 (N_20603,N_19531,N_19187);
or U20604 (N_20604,N_19195,N_19496);
nor U20605 (N_20605,N_19620,N_19315);
nor U20606 (N_20606,N_19993,N_19910);
and U20607 (N_20607,N_19405,N_19864);
xnor U20608 (N_20608,N_19700,N_19518);
or U20609 (N_20609,N_19224,N_19179);
and U20610 (N_20610,N_19470,N_19280);
or U20611 (N_20611,N_19730,N_19810);
nand U20612 (N_20612,N_19723,N_19188);
xnor U20613 (N_20613,N_19262,N_19211);
and U20614 (N_20614,N_19764,N_19639);
nor U20615 (N_20615,N_19847,N_19456);
nand U20616 (N_20616,N_19801,N_19961);
nand U20617 (N_20617,N_19420,N_19885);
nand U20618 (N_20618,N_19734,N_19804);
nor U20619 (N_20619,N_19889,N_19540);
xor U20620 (N_20620,N_19291,N_19801);
and U20621 (N_20621,N_19071,N_19609);
and U20622 (N_20622,N_19291,N_19713);
or U20623 (N_20623,N_19787,N_19550);
nand U20624 (N_20624,N_19997,N_19446);
nand U20625 (N_20625,N_19688,N_19243);
nor U20626 (N_20626,N_19155,N_19830);
nor U20627 (N_20627,N_19295,N_19806);
nor U20628 (N_20628,N_19935,N_19421);
nor U20629 (N_20629,N_19926,N_19125);
xnor U20630 (N_20630,N_19582,N_19609);
nand U20631 (N_20631,N_19955,N_19839);
or U20632 (N_20632,N_19087,N_19508);
or U20633 (N_20633,N_19858,N_19953);
and U20634 (N_20634,N_19795,N_19672);
or U20635 (N_20635,N_19736,N_19538);
nor U20636 (N_20636,N_19210,N_19073);
or U20637 (N_20637,N_19456,N_19845);
and U20638 (N_20638,N_19437,N_19970);
and U20639 (N_20639,N_19765,N_19392);
nand U20640 (N_20640,N_19983,N_19930);
or U20641 (N_20641,N_19334,N_19669);
and U20642 (N_20642,N_19239,N_19989);
and U20643 (N_20643,N_19255,N_19268);
xnor U20644 (N_20644,N_19400,N_19976);
or U20645 (N_20645,N_19251,N_19245);
and U20646 (N_20646,N_19986,N_19364);
and U20647 (N_20647,N_19505,N_19453);
xnor U20648 (N_20648,N_19723,N_19294);
nor U20649 (N_20649,N_19938,N_19965);
nand U20650 (N_20650,N_19427,N_19103);
nor U20651 (N_20651,N_19579,N_19852);
nor U20652 (N_20652,N_19569,N_19891);
or U20653 (N_20653,N_19582,N_19426);
xnor U20654 (N_20654,N_19268,N_19584);
and U20655 (N_20655,N_19890,N_19654);
or U20656 (N_20656,N_19212,N_19851);
or U20657 (N_20657,N_19955,N_19403);
nor U20658 (N_20658,N_19701,N_19954);
or U20659 (N_20659,N_19690,N_19350);
nand U20660 (N_20660,N_19920,N_19560);
and U20661 (N_20661,N_19113,N_19217);
and U20662 (N_20662,N_19099,N_19337);
and U20663 (N_20663,N_19883,N_19922);
xor U20664 (N_20664,N_19215,N_19662);
nor U20665 (N_20665,N_19364,N_19156);
and U20666 (N_20666,N_19253,N_19682);
xnor U20667 (N_20667,N_19731,N_19872);
xnor U20668 (N_20668,N_19757,N_19451);
xnor U20669 (N_20669,N_19199,N_19371);
nor U20670 (N_20670,N_19741,N_19203);
or U20671 (N_20671,N_19553,N_19192);
xor U20672 (N_20672,N_19041,N_19514);
and U20673 (N_20673,N_19440,N_19752);
nor U20674 (N_20674,N_19705,N_19701);
and U20675 (N_20675,N_19297,N_19043);
and U20676 (N_20676,N_19500,N_19606);
and U20677 (N_20677,N_19866,N_19864);
xnor U20678 (N_20678,N_19574,N_19147);
nor U20679 (N_20679,N_19833,N_19266);
nor U20680 (N_20680,N_19826,N_19603);
nor U20681 (N_20681,N_19172,N_19544);
or U20682 (N_20682,N_19743,N_19262);
or U20683 (N_20683,N_19349,N_19935);
nor U20684 (N_20684,N_19502,N_19505);
nor U20685 (N_20685,N_19552,N_19928);
nor U20686 (N_20686,N_19069,N_19460);
nor U20687 (N_20687,N_19757,N_19806);
nor U20688 (N_20688,N_19169,N_19939);
nand U20689 (N_20689,N_19983,N_19329);
or U20690 (N_20690,N_19050,N_19580);
and U20691 (N_20691,N_19353,N_19971);
nor U20692 (N_20692,N_19465,N_19361);
nand U20693 (N_20693,N_19563,N_19821);
nand U20694 (N_20694,N_19416,N_19476);
xor U20695 (N_20695,N_19942,N_19664);
or U20696 (N_20696,N_19204,N_19438);
and U20697 (N_20697,N_19072,N_19839);
nor U20698 (N_20698,N_19523,N_19974);
nor U20699 (N_20699,N_19791,N_19201);
nand U20700 (N_20700,N_19424,N_19448);
and U20701 (N_20701,N_19842,N_19821);
nor U20702 (N_20702,N_19545,N_19278);
or U20703 (N_20703,N_19424,N_19512);
nand U20704 (N_20704,N_19511,N_19668);
or U20705 (N_20705,N_19608,N_19170);
or U20706 (N_20706,N_19059,N_19838);
xor U20707 (N_20707,N_19141,N_19161);
or U20708 (N_20708,N_19032,N_19315);
and U20709 (N_20709,N_19174,N_19238);
or U20710 (N_20710,N_19746,N_19456);
nand U20711 (N_20711,N_19798,N_19070);
xor U20712 (N_20712,N_19036,N_19855);
xor U20713 (N_20713,N_19411,N_19465);
xor U20714 (N_20714,N_19476,N_19614);
and U20715 (N_20715,N_19052,N_19193);
or U20716 (N_20716,N_19674,N_19605);
and U20717 (N_20717,N_19559,N_19284);
xnor U20718 (N_20718,N_19355,N_19013);
xnor U20719 (N_20719,N_19583,N_19135);
nand U20720 (N_20720,N_19312,N_19909);
and U20721 (N_20721,N_19595,N_19825);
xnor U20722 (N_20722,N_19788,N_19889);
and U20723 (N_20723,N_19145,N_19836);
nand U20724 (N_20724,N_19546,N_19056);
nor U20725 (N_20725,N_19318,N_19748);
nor U20726 (N_20726,N_19267,N_19973);
and U20727 (N_20727,N_19005,N_19748);
and U20728 (N_20728,N_19876,N_19387);
nand U20729 (N_20729,N_19513,N_19519);
xnor U20730 (N_20730,N_19775,N_19330);
xor U20731 (N_20731,N_19843,N_19095);
and U20732 (N_20732,N_19341,N_19820);
xnor U20733 (N_20733,N_19780,N_19404);
and U20734 (N_20734,N_19074,N_19471);
or U20735 (N_20735,N_19966,N_19301);
and U20736 (N_20736,N_19689,N_19297);
and U20737 (N_20737,N_19920,N_19108);
and U20738 (N_20738,N_19147,N_19962);
nor U20739 (N_20739,N_19192,N_19333);
nor U20740 (N_20740,N_19955,N_19370);
or U20741 (N_20741,N_19308,N_19054);
nand U20742 (N_20742,N_19453,N_19708);
xnor U20743 (N_20743,N_19167,N_19387);
or U20744 (N_20744,N_19588,N_19912);
and U20745 (N_20745,N_19506,N_19985);
nor U20746 (N_20746,N_19848,N_19282);
and U20747 (N_20747,N_19059,N_19382);
nand U20748 (N_20748,N_19915,N_19392);
nor U20749 (N_20749,N_19183,N_19046);
xnor U20750 (N_20750,N_19379,N_19786);
nand U20751 (N_20751,N_19049,N_19886);
nor U20752 (N_20752,N_19188,N_19900);
and U20753 (N_20753,N_19827,N_19393);
xnor U20754 (N_20754,N_19486,N_19160);
or U20755 (N_20755,N_19210,N_19269);
nand U20756 (N_20756,N_19188,N_19402);
xnor U20757 (N_20757,N_19689,N_19843);
nor U20758 (N_20758,N_19131,N_19442);
or U20759 (N_20759,N_19369,N_19229);
xor U20760 (N_20760,N_19365,N_19475);
xnor U20761 (N_20761,N_19121,N_19325);
xor U20762 (N_20762,N_19389,N_19890);
nor U20763 (N_20763,N_19709,N_19544);
or U20764 (N_20764,N_19167,N_19650);
xnor U20765 (N_20765,N_19463,N_19416);
xor U20766 (N_20766,N_19348,N_19950);
xor U20767 (N_20767,N_19358,N_19942);
xor U20768 (N_20768,N_19272,N_19133);
xnor U20769 (N_20769,N_19101,N_19097);
nand U20770 (N_20770,N_19483,N_19500);
or U20771 (N_20771,N_19031,N_19573);
nand U20772 (N_20772,N_19354,N_19272);
nor U20773 (N_20773,N_19047,N_19340);
and U20774 (N_20774,N_19075,N_19636);
nand U20775 (N_20775,N_19206,N_19418);
xnor U20776 (N_20776,N_19749,N_19018);
and U20777 (N_20777,N_19713,N_19565);
nor U20778 (N_20778,N_19964,N_19020);
xnor U20779 (N_20779,N_19345,N_19514);
xor U20780 (N_20780,N_19036,N_19156);
nand U20781 (N_20781,N_19769,N_19623);
and U20782 (N_20782,N_19873,N_19482);
or U20783 (N_20783,N_19155,N_19568);
nor U20784 (N_20784,N_19727,N_19816);
and U20785 (N_20785,N_19261,N_19247);
or U20786 (N_20786,N_19994,N_19717);
or U20787 (N_20787,N_19802,N_19288);
xor U20788 (N_20788,N_19655,N_19462);
xnor U20789 (N_20789,N_19989,N_19157);
xor U20790 (N_20790,N_19464,N_19871);
or U20791 (N_20791,N_19445,N_19055);
nand U20792 (N_20792,N_19793,N_19605);
nor U20793 (N_20793,N_19180,N_19246);
nand U20794 (N_20794,N_19250,N_19329);
nor U20795 (N_20795,N_19520,N_19748);
xnor U20796 (N_20796,N_19351,N_19594);
xnor U20797 (N_20797,N_19383,N_19886);
xor U20798 (N_20798,N_19825,N_19152);
nor U20799 (N_20799,N_19086,N_19793);
and U20800 (N_20800,N_19936,N_19767);
and U20801 (N_20801,N_19442,N_19689);
nor U20802 (N_20802,N_19037,N_19973);
nor U20803 (N_20803,N_19047,N_19581);
and U20804 (N_20804,N_19230,N_19204);
or U20805 (N_20805,N_19696,N_19027);
nand U20806 (N_20806,N_19368,N_19887);
nand U20807 (N_20807,N_19165,N_19445);
nand U20808 (N_20808,N_19580,N_19878);
nand U20809 (N_20809,N_19006,N_19641);
nand U20810 (N_20810,N_19731,N_19787);
and U20811 (N_20811,N_19279,N_19602);
or U20812 (N_20812,N_19206,N_19636);
nor U20813 (N_20813,N_19454,N_19074);
or U20814 (N_20814,N_19877,N_19556);
and U20815 (N_20815,N_19424,N_19868);
xor U20816 (N_20816,N_19146,N_19904);
and U20817 (N_20817,N_19793,N_19376);
or U20818 (N_20818,N_19174,N_19824);
nor U20819 (N_20819,N_19336,N_19091);
nor U20820 (N_20820,N_19838,N_19675);
xor U20821 (N_20821,N_19089,N_19651);
and U20822 (N_20822,N_19566,N_19081);
or U20823 (N_20823,N_19757,N_19892);
or U20824 (N_20824,N_19637,N_19605);
or U20825 (N_20825,N_19362,N_19203);
nor U20826 (N_20826,N_19527,N_19930);
nand U20827 (N_20827,N_19061,N_19911);
nor U20828 (N_20828,N_19541,N_19314);
nand U20829 (N_20829,N_19816,N_19981);
nand U20830 (N_20830,N_19447,N_19756);
nor U20831 (N_20831,N_19403,N_19914);
nand U20832 (N_20832,N_19909,N_19464);
and U20833 (N_20833,N_19813,N_19412);
xor U20834 (N_20834,N_19041,N_19992);
nand U20835 (N_20835,N_19310,N_19140);
xnor U20836 (N_20836,N_19412,N_19685);
nand U20837 (N_20837,N_19473,N_19760);
xnor U20838 (N_20838,N_19878,N_19746);
nor U20839 (N_20839,N_19567,N_19145);
and U20840 (N_20840,N_19495,N_19931);
or U20841 (N_20841,N_19242,N_19070);
or U20842 (N_20842,N_19211,N_19024);
xor U20843 (N_20843,N_19571,N_19755);
and U20844 (N_20844,N_19960,N_19843);
nor U20845 (N_20845,N_19895,N_19314);
nor U20846 (N_20846,N_19825,N_19719);
or U20847 (N_20847,N_19692,N_19981);
nand U20848 (N_20848,N_19147,N_19089);
and U20849 (N_20849,N_19263,N_19783);
nand U20850 (N_20850,N_19366,N_19115);
and U20851 (N_20851,N_19267,N_19547);
and U20852 (N_20852,N_19065,N_19214);
nand U20853 (N_20853,N_19311,N_19245);
and U20854 (N_20854,N_19334,N_19622);
or U20855 (N_20855,N_19358,N_19628);
xor U20856 (N_20856,N_19096,N_19042);
nand U20857 (N_20857,N_19579,N_19096);
or U20858 (N_20858,N_19104,N_19662);
nand U20859 (N_20859,N_19842,N_19000);
or U20860 (N_20860,N_19760,N_19845);
nand U20861 (N_20861,N_19936,N_19495);
and U20862 (N_20862,N_19657,N_19036);
nand U20863 (N_20863,N_19017,N_19673);
nor U20864 (N_20864,N_19509,N_19084);
nor U20865 (N_20865,N_19226,N_19321);
and U20866 (N_20866,N_19547,N_19825);
or U20867 (N_20867,N_19637,N_19479);
or U20868 (N_20868,N_19218,N_19391);
or U20869 (N_20869,N_19789,N_19892);
or U20870 (N_20870,N_19670,N_19219);
and U20871 (N_20871,N_19918,N_19603);
nand U20872 (N_20872,N_19586,N_19011);
and U20873 (N_20873,N_19753,N_19561);
and U20874 (N_20874,N_19170,N_19027);
nor U20875 (N_20875,N_19703,N_19761);
xor U20876 (N_20876,N_19299,N_19049);
or U20877 (N_20877,N_19804,N_19534);
nor U20878 (N_20878,N_19457,N_19997);
or U20879 (N_20879,N_19727,N_19934);
nand U20880 (N_20880,N_19722,N_19571);
nand U20881 (N_20881,N_19364,N_19731);
or U20882 (N_20882,N_19958,N_19130);
xor U20883 (N_20883,N_19340,N_19216);
nor U20884 (N_20884,N_19477,N_19804);
nand U20885 (N_20885,N_19596,N_19109);
or U20886 (N_20886,N_19822,N_19903);
xnor U20887 (N_20887,N_19669,N_19306);
nand U20888 (N_20888,N_19520,N_19523);
or U20889 (N_20889,N_19790,N_19639);
nand U20890 (N_20890,N_19289,N_19976);
xnor U20891 (N_20891,N_19403,N_19727);
xnor U20892 (N_20892,N_19937,N_19961);
or U20893 (N_20893,N_19932,N_19321);
nor U20894 (N_20894,N_19120,N_19406);
or U20895 (N_20895,N_19751,N_19347);
nand U20896 (N_20896,N_19646,N_19073);
nor U20897 (N_20897,N_19261,N_19986);
nor U20898 (N_20898,N_19534,N_19106);
or U20899 (N_20899,N_19683,N_19081);
nor U20900 (N_20900,N_19863,N_19714);
nor U20901 (N_20901,N_19905,N_19184);
or U20902 (N_20902,N_19758,N_19561);
nand U20903 (N_20903,N_19868,N_19955);
xor U20904 (N_20904,N_19352,N_19839);
nor U20905 (N_20905,N_19286,N_19518);
or U20906 (N_20906,N_19748,N_19624);
nor U20907 (N_20907,N_19382,N_19943);
and U20908 (N_20908,N_19673,N_19039);
and U20909 (N_20909,N_19397,N_19769);
nor U20910 (N_20910,N_19623,N_19723);
xor U20911 (N_20911,N_19707,N_19679);
or U20912 (N_20912,N_19984,N_19951);
and U20913 (N_20913,N_19123,N_19282);
or U20914 (N_20914,N_19632,N_19670);
xnor U20915 (N_20915,N_19051,N_19577);
or U20916 (N_20916,N_19158,N_19762);
or U20917 (N_20917,N_19935,N_19741);
or U20918 (N_20918,N_19904,N_19827);
and U20919 (N_20919,N_19161,N_19316);
nor U20920 (N_20920,N_19853,N_19111);
and U20921 (N_20921,N_19047,N_19683);
or U20922 (N_20922,N_19741,N_19551);
nand U20923 (N_20923,N_19143,N_19329);
xor U20924 (N_20924,N_19615,N_19783);
nor U20925 (N_20925,N_19368,N_19414);
or U20926 (N_20926,N_19662,N_19268);
nand U20927 (N_20927,N_19563,N_19323);
and U20928 (N_20928,N_19044,N_19176);
nand U20929 (N_20929,N_19641,N_19250);
xnor U20930 (N_20930,N_19564,N_19068);
or U20931 (N_20931,N_19985,N_19317);
xor U20932 (N_20932,N_19598,N_19845);
nor U20933 (N_20933,N_19220,N_19855);
nor U20934 (N_20934,N_19566,N_19680);
nand U20935 (N_20935,N_19821,N_19525);
nand U20936 (N_20936,N_19011,N_19921);
or U20937 (N_20937,N_19741,N_19886);
nand U20938 (N_20938,N_19415,N_19418);
xor U20939 (N_20939,N_19421,N_19516);
and U20940 (N_20940,N_19112,N_19879);
nor U20941 (N_20941,N_19739,N_19895);
and U20942 (N_20942,N_19093,N_19865);
nor U20943 (N_20943,N_19374,N_19145);
and U20944 (N_20944,N_19055,N_19469);
and U20945 (N_20945,N_19681,N_19027);
nand U20946 (N_20946,N_19931,N_19887);
xnor U20947 (N_20947,N_19978,N_19797);
nor U20948 (N_20948,N_19769,N_19820);
and U20949 (N_20949,N_19933,N_19798);
or U20950 (N_20950,N_19053,N_19557);
and U20951 (N_20951,N_19911,N_19958);
or U20952 (N_20952,N_19059,N_19429);
nand U20953 (N_20953,N_19997,N_19711);
xor U20954 (N_20954,N_19120,N_19461);
or U20955 (N_20955,N_19717,N_19351);
nor U20956 (N_20956,N_19195,N_19313);
and U20957 (N_20957,N_19878,N_19309);
nand U20958 (N_20958,N_19302,N_19678);
and U20959 (N_20959,N_19646,N_19189);
nor U20960 (N_20960,N_19420,N_19564);
nor U20961 (N_20961,N_19752,N_19146);
nand U20962 (N_20962,N_19730,N_19547);
nor U20963 (N_20963,N_19196,N_19281);
nand U20964 (N_20964,N_19757,N_19216);
nand U20965 (N_20965,N_19890,N_19138);
nand U20966 (N_20966,N_19702,N_19372);
xnor U20967 (N_20967,N_19568,N_19606);
nor U20968 (N_20968,N_19014,N_19807);
and U20969 (N_20969,N_19411,N_19214);
and U20970 (N_20970,N_19672,N_19596);
nor U20971 (N_20971,N_19216,N_19429);
nor U20972 (N_20972,N_19271,N_19569);
nor U20973 (N_20973,N_19783,N_19010);
and U20974 (N_20974,N_19345,N_19537);
and U20975 (N_20975,N_19495,N_19649);
and U20976 (N_20976,N_19860,N_19685);
and U20977 (N_20977,N_19727,N_19931);
or U20978 (N_20978,N_19230,N_19668);
nand U20979 (N_20979,N_19577,N_19148);
xnor U20980 (N_20980,N_19055,N_19919);
nand U20981 (N_20981,N_19628,N_19743);
xor U20982 (N_20982,N_19999,N_19279);
or U20983 (N_20983,N_19399,N_19442);
nor U20984 (N_20984,N_19272,N_19832);
nand U20985 (N_20985,N_19836,N_19114);
xnor U20986 (N_20986,N_19687,N_19568);
nor U20987 (N_20987,N_19547,N_19446);
or U20988 (N_20988,N_19410,N_19966);
xor U20989 (N_20989,N_19046,N_19524);
and U20990 (N_20990,N_19319,N_19343);
or U20991 (N_20991,N_19313,N_19027);
xor U20992 (N_20992,N_19419,N_19075);
nor U20993 (N_20993,N_19029,N_19500);
and U20994 (N_20994,N_19712,N_19580);
nand U20995 (N_20995,N_19098,N_19777);
nand U20996 (N_20996,N_19816,N_19283);
nor U20997 (N_20997,N_19759,N_19476);
nand U20998 (N_20998,N_19178,N_19190);
and U20999 (N_20999,N_19907,N_19814);
nand U21000 (N_21000,N_20223,N_20685);
nand U21001 (N_21001,N_20792,N_20087);
nand U21002 (N_21002,N_20882,N_20316);
and U21003 (N_21003,N_20907,N_20432);
and U21004 (N_21004,N_20412,N_20005);
and U21005 (N_21005,N_20219,N_20177);
xnor U21006 (N_21006,N_20894,N_20895);
nor U21007 (N_21007,N_20926,N_20850);
and U21008 (N_21008,N_20269,N_20286);
and U21009 (N_21009,N_20035,N_20231);
nor U21010 (N_21010,N_20298,N_20478);
xor U21011 (N_21011,N_20575,N_20550);
xnor U21012 (N_21012,N_20862,N_20527);
nand U21013 (N_21013,N_20119,N_20936);
or U21014 (N_21014,N_20167,N_20910);
nor U21015 (N_21015,N_20331,N_20008);
and U21016 (N_21016,N_20111,N_20442);
xor U21017 (N_21017,N_20144,N_20509);
nor U21018 (N_21018,N_20308,N_20507);
nand U21019 (N_21019,N_20612,N_20299);
nand U21020 (N_21020,N_20236,N_20967);
nand U21021 (N_21021,N_20040,N_20013);
xnor U21022 (N_21022,N_20654,N_20991);
or U21023 (N_21023,N_20402,N_20597);
nor U21024 (N_21024,N_20630,N_20650);
xnor U21025 (N_21025,N_20257,N_20004);
or U21026 (N_21026,N_20747,N_20871);
and U21027 (N_21027,N_20136,N_20033);
nand U21028 (N_21028,N_20373,N_20572);
and U21029 (N_21029,N_20647,N_20904);
xor U21030 (N_21030,N_20184,N_20954);
and U21031 (N_21031,N_20890,N_20424);
xnor U21032 (N_21032,N_20985,N_20578);
xnor U21033 (N_21033,N_20073,N_20157);
nand U21034 (N_21034,N_20672,N_20729);
nand U21035 (N_21035,N_20237,N_20543);
or U21036 (N_21036,N_20878,N_20334);
nand U21037 (N_21037,N_20381,N_20680);
nand U21038 (N_21038,N_20275,N_20888);
xnor U21039 (N_21039,N_20526,N_20185);
and U21040 (N_21040,N_20302,N_20753);
or U21041 (N_21041,N_20273,N_20559);
nand U21042 (N_21042,N_20263,N_20925);
nand U21043 (N_21043,N_20815,N_20287);
xnor U21044 (N_21044,N_20928,N_20706);
nand U21045 (N_21045,N_20554,N_20030);
and U21046 (N_21046,N_20682,N_20834);
nor U21047 (N_21047,N_20999,N_20305);
nand U21048 (N_21048,N_20588,N_20245);
xor U21049 (N_21049,N_20677,N_20240);
and U21050 (N_21050,N_20494,N_20060);
nand U21051 (N_21051,N_20425,N_20534);
or U21052 (N_21052,N_20149,N_20312);
or U21053 (N_21053,N_20718,N_20842);
nand U21054 (N_21054,N_20746,N_20439);
xnor U21055 (N_21055,N_20311,N_20964);
nor U21056 (N_21056,N_20020,N_20464);
nand U21057 (N_21057,N_20244,N_20376);
nor U21058 (N_21058,N_20480,N_20186);
xor U21059 (N_21059,N_20931,N_20912);
or U21060 (N_21060,N_20134,N_20486);
xnor U21061 (N_21061,N_20835,N_20600);
nand U21062 (N_21062,N_20864,N_20128);
nand U21063 (N_21063,N_20582,N_20504);
nand U21064 (N_21064,N_20730,N_20972);
xnor U21065 (N_21065,N_20467,N_20566);
nand U21066 (N_21066,N_20561,N_20495);
xnor U21067 (N_21067,N_20084,N_20556);
xor U21068 (N_21068,N_20352,N_20713);
or U21069 (N_21069,N_20262,N_20632);
or U21070 (N_21070,N_20328,N_20569);
xor U21071 (N_21071,N_20103,N_20209);
nand U21072 (N_21072,N_20121,N_20044);
and U21073 (N_21073,N_20843,N_20962);
and U21074 (N_21074,N_20268,N_20333);
nand U21075 (N_21075,N_20868,N_20330);
and U21076 (N_21076,N_20293,N_20071);
xor U21077 (N_21077,N_20295,N_20978);
nand U21078 (N_21078,N_20857,N_20806);
nand U21079 (N_21079,N_20518,N_20047);
or U21080 (N_21080,N_20711,N_20960);
and U21081 (N_21081,N_20933,N_20377);
nor U21082 (N_21082,N_20454,N_20015);
nand U21083 (N_21083,N_20175,N_20590);
or U21084 (N_21084,N_20816,N_20292);
and U21085 (N_21085,N_20796,N_20836);
or U21086 (N_21086,N_20459,N_20000);
nand U21087 (N_21087,N_20318,N_20341);
nor U21088 (N_21088,N_20965,N_20327);
nor U21089 (N_21089,N_20165,N_20877);
and U21090 (N_21090,N_20276,N_20876);
or U21091 (N_21091,N_20143,N_20421);
or U21092 (N_21092,N_20752,N_20045);
and U21093 (N_21093,N_20351,N_20409);
nand U21094 (N_21094,N_20780,N_20675);
and U21095 (N_21095,N_20542,N_20379);
or U21096 (N_21096,N_20174,N_20118);
or U21097 (N_21097,N_20885,N_20468);
and U21098 (N_21098,N_20131,N_20354);
or U21099 (N_21099,N_20445,N_20350);
and U21100 (N_21100,N_20538,N_20717);
nor U21101 (N_21101,N_20761,N_20707);
xnor U21102 (N_21102,N_20763,N_20493);
and U21103 (N_21103,N_20473,N_20902);
or U21104 (N_21104,N_20019,N_20749);
nor U21105 (N_21105,N_20031,N_20636);
nand U21106 (N_21106,N_20499,N_20633);
xor U21107 (N_21107,N_20986,N_20858);
or U21108 (N_21108,N_20502,N_20036);
nand U21109 (N_21109,N_20724,N_20935);
xnor U21110 (N_21110,N_20610,N_20026);
xnor U21111 (N_21111,N_20346,N_20148);
nor U21112 (N_21112,N_20197,N_20152);
and U21113 (N_21113,N_20889,N_20697);
or U21114 (N_21114,N_20827,N_20670);
nand U21115 (N_21115,N_20759,N_20553);
nand U21116 (N_21116,N_20129,N_20058);
xor U21117 (N_21117,N_20039,N_20475);
and U21118 (N_21118,N_20782,N_20199);
nand U21119 (N_21119,N_20260,N_20874);
and U21120 (N_21120,N_20684,N_20604);
xnor U21121 (N_21121,N_20043,N_20090);
and U21122 (N_21122,N_20080,N_20410);
and U21123 (N_21123,N_20279,N_20731);
nor U21124 (N_21124,N_20694,N_20700);
and U21125 (N_21125,N_20422,N_20229);
and U21126 (N_21126,N_20998,N_20809);
nor U21127 (N_21127,N_20360,N_20411);
xnor U21128 (N_21128,N_20772,N_20142);
or U21129 (N_21129,N_20021,N_20726);
xor U21130 (N_21130,N_20062,N_20066);
xnor U21131 (N_21131,N_20951,N_20251);
xor U21132 (N_21132,N_20042,N_20905);
nand U21133 (N_21133,N_20117,N_20278);
nor U21134 (N_21134,N_20304,N_20640);
or U21135 (N_21135,N_20793,N_20235);
nor U21136 (N_21136,N_20139,N_20628);
and U21137 (N_21137,N_20108,N_20290);
xor U21138 (N_21138,N_20703,N_20748);
nor U21139 (N_21139,N_20329,N_20055);
and U21140 (N_21140,N_20022,N_20539);
or U21141 (N_21141,N_20392,N_20068);
xor U21142 (N_21142,N_20384,N_20714);
and U21143 (N_21143,N_20133,N_20923);
nor U21144 (N_21144,N_20363,N_20938);
nand U21145 (N_21145,N_20820,N_20064);
or U21146 (N_21146,N_20389,N_20678);
and U21147 (N_21147,N_20007,N_20088);
nor U21148 (N_21148,N_20297,N_20823);
nand U21149 (N_21149,N_20147,N_20406);
nand U21150 (N_21150,N_20140,N_20973);
xnor U21151 (N_21151,N_20181,N_20396);
nor U21152 (N_21152,N_20104,N_20638);
or U21153 (N_21153,N_20949,N_20370);
nor U21154 (N_21154,N_20228,N_20288);
or U21155 (N_21155,N_20547,N_20603);
and U21156 (N_21156,N_20217,N_20623);
nor U21157 (N_21157,N_20997,N_20848);
nor U21158 (N_21158,N_20880,N_20657);
xnor U21159 (N_21159,N_20621,N_20110);
or U21160 (N_21160,N_20735,N_20191);
nor U21161 (N_21161,N_20977,N_20272);
xnor U21162 (N_21162,N_20161,N_20570);
nand U21163 (N_21163,N_20479,N_20941);
xnor U21164 (N_21164,N_20616,N_20881);
nor U21165 (N_21165,N_20914,N_20562);
nand U21166 (N_21166,N_20664,N_20595);
or U21167 (N_21167,N_20461,N_20852);
nand U21168 (N_21168,N_20799,N_20125);
and U21169 (N_21169,N_20057,N_20294);
nand U21170 (N_21170,N_20845,N_20601);
or U21171 (N_21171,N_20641,N_20206);
nor U21172 (N_21172,N_20488,N_20750);
nand U21173 (N_21173,N_20227,N_20025);
or U21174 (N_21174,N_20375,N_20489);
nor U21175 (N_21175,N_20577,N_20916);
and U21176 (N_21176,N_20520,N_20808);
xor U21177 (N_21177,N_20401,N_20795);
nor U21178 (N_21178,N_20082,N_20383);
and U21179 (N_21179,N_20307,N_20500);
nor U21180 (N_21180,N_20844,N_20497);
and U21181 (N_21181,N_20803,N_20230);
xnor U21182 (N_21182,N_20911,N_20146);
nand U21183 (N_21183,N_20573,N_20754);
xnor U21184 (N_21184,N_20899,N_20180);
nand U21185 (N_21185,N_20611,N_20691);
nand U21186 (N_21186,N_20172,N_20221);
nor U21187 (N_21187,N_20705,N_20183);
nand U21188 (N_21188,N_20557,N_20982);
xnor U21189 (N_21189,N_20704,N_20618);
xor U21190 (N_21190,N_20154,N_20281);
nand U21191 (N_21191,N_20443,N_20742);
nand U21192 (N_21192,N_20313,N_20980);
nand U21193 (N_21193,N_20171,N_20825);
nand U21194 (N_21194,N_20107,N_20721);
nor U21195 (N_21195,N_20741,N_20810);
nand U21196 (N_21196,N_20574,N_20458);
nor U21197 (N_21197,N_20204,N_20284);
nor U21198 (N_21198,N_20248,N_20947);
or U21199 (N_21199,N_20884,N_20169);
nor U21200 (N_21200,N_20599,N_20336);
or U21201 (N_21201,N_20849,N_20851);
nand U21202 (N_21202,N_20176,N_20247);
nand U21203 (N_21203,N_20188,N_20395);
nor U21204 (N_21204,N_20723,N_20265);
nand U21205 (N_21205,N_20001,N_20854);
and U21206 (N_21206,N_20743,N_20920);
or U21207 (N_21207,N_20764,N_20563);
and U21208 (N_21208,N_20788,N_20699);
and U21209 (N_21209,N_20434,N_20783);
xnor U21210 (N_21210,N_20692,N_20813);
and U21211 (N_21211,N_20267,N_20061);
nand U21212 (N_21212,N_20010,N_20866);
nor U21213 (N_21213,N_20417,N_20405);
nand U21214 (N_21214,N_20974,N_20833);
nand U21215 (N_21215,N_20163,N_20745);
and U21216 (N_21216,N_20074,N_20734);
nand U21217 (N_21217,N_20988,N_20164);
and U21218 (N_21218,N_20637,N_20626);
xnor U21219 (N_21219,N_20246,N_20676);
or U21220 (N_21220,N_20644,N_20335);
nor U21221 (N_21221,N_20800,N_20506);
nand U21222 (N_21222,N_20853,N_20971);
nor U21223 (N_21223,N_20940,N_20598);
or U21224 (N_21224,N_20444,N_20112);
and U21225 (N_21225,N_20322,N_20791);
and U21226 (N_21226,N_20870,N_20846);
nand U21227 (N_21227,N_20744,N_20314);
or U21228 (N_21228,N_20673,N_20252);
nand U21229 (N_21229,N_20887,N_20465);
nor U21230 (N_21230,N_20138,N_20091);
nor U21231 (N_21231,N_20525,N_20811);
nor U21232 (N_21232,N_20725,N_20403);
and U21233 (N_21233,N_20285,N_20807);
xor U21234 (N_21234,N_20583,N_20652);
xor U21235 (N_21235,N_20576,N_20875);
and U21236 (N_21236,N_20116,N_20660);
and U21237 (N_21237,N_20189,N_20303);
and U21238 (N_21238,N_20266,N_20173);
and U21239 (N_21239,N_20708,N_20918);
or U21240 (N_21240,N_20786,N_20115);
nand U21241 (N_21241,N_20153,N_20737);
and U21242 (N_21242,N_20837,N_20602);
xor U21243 (N_21243,N_20581,N_20089);
and U21244 (N_21244,N_20016,N_20215);
or U21245 (N_21245,N_20102,N_20767);
xnor U21246 (N_21246,N_20032,N_20201);
and U21247 (N_21247,N_20420,N_20552);
and U21248 (N_21248,N_20913,N_20380);
xor U21249 (N_21249,N_20873,N_20413);
nor U21250 (N_21250,N_20289,N_20642);
nand U21251 (N_21251,N_20211,N_20757);
xnor U21252 (N_21252,N_20399,N_20930);
nand U21253 (N_21253,N_20254,N_20233);
or U21254 (N_21254,N_20781,N_20270);
nand U21255 (N_21255,N_20716,N_20255);
nor U21256 (N_21256,N_20300,N_20242);
and U21257 (N_21257,N_20106,N_20041);
and U21258 (N_21258,N_20798,N_20948);
xnor U21259 (N_21259,N_20415,N_20407);
or U21260 (N_21260,N_20447,N_20605);
and U21261 (N_21261,N_20879,N_20961);
and U21262 (N_21262,N_20586,N_20661);
nand U21263 (N_21263,N_20096,N_20225);
xor U21264 (N_21264,N_20984,N_20338);
nand U21265 (N_21265,N_20987,N_20368);
and U21266 (N_21266,N_20469,N_20006);
xor U21267 (N_21267,N_20277,N_20306);
nand U21268 (N_21268,N_20388,N_20950);
xor U21269 (N_21269,N_20579,N_20785);
nand U21270 (N_21270,N_20200,N_20009);
nand U21271 (N_21271,N_20264,N_20756);
nor U21272 (N_21272,N_20929,N_20733);
or U21273 (N_21273,N_20135,N_20466);
nand U21274 (N_21274,N_20414,N_20514);
and U21275 (N_21275,N_20470,N_20541);
xnor U21276 (N_21276,N_20448,N_20531);
nand U21277 (N_21277,N_20883,N_20766);
or U21278 (N_21278,N_20840,N_20720);
nor U21279 (N_21279,N_20155,N_20450);
nor U21280 (N_21280,N_20571,N_20474);
or U21281 (N_21281,N_20784,N_20830);
or U21282 (N_21282,N_20968,N_20822);
nand U21283 (N_21283,N_20770,N_20337);
nor U21284 (N_21284,N_20683,N_20615);
or U21285 (N_21285,N_20937,N_20841);
and U21286 (N_21286,N_20151,N_20361);
and U21287 (N_21287,N_20100,N_20635);
or U21288 (N_21288,N_20908,N_20995);
nand U21289 (N_21289,N_20012,N_20340);
nor U21290 (N_21290,N_20378,N_20053);
nor U21291 (N_21291,N_20498,N_20606);
nor U21292 (N_21292,N_20086,N_20769);
or U21293 (N_21293,N_20787,N_20324);
and U21294 (N_21294,N_20491,N_20867);
nor U21295 (N_21295,N_20709,N_20326);
and U21296 (N_21296,N_20034,N_20693);
nand U21297 (N_21297,N_20449,N_20668);
and U21298 (N_21298,N_20777,N_20418);
nor U21299 (N_21299,N_20046,N_20301);
or U21300 (N_21300,N_20567,N_20762);
or U21301 (N_21301,N_20958,N_20438);
nor U21302 (N_21302,N_20076,N_20536);
and U21303 (N_21303,N_20460,N_20924);
and U21304 (N_21304,N_20521,N_20014);
or U21305 (N_21305,N_20123,N_20054);
and U21306 (N_21306,N_20203,N_20390);
and U21307 (N_21307,N_20695,N_20214);
xnor U21308 (N_21308,N_20942,N_20440);
nor U21309 (N_21309,N_20321,N_20701);
nor U21310 (N_21310,N_20508,N_20093);
nor U21311 (N_21311,N_20946,N_20037);
nor U21312 (N_21312,N_20622,N_20528);
or U21313 (N_21313,N_20667,N_20487);
and U21314 (N_21314,N_20476,N_20775);
nor U21315 (N_21315,N_20249,N_20639);
or U21316 (N_21316,N_20210,N_20385);
and U21317 (N_21317,N_20627,N_20715);
or U21318 (N_21318,N_20532,N_20095);
xor U21319 (N_21319,N_20921,N_20819);
and U21320 (N_21320,N_20092,N_20317);
and U21321 (N_21321,N_20537,N_20397);
xor U21322 (N_21322,N_20944,N_20271);
nor U21323 (N_21323,N_20592,N_20482);
xor U21324 (N_21324,N_20625,N_20256);
or U21325 (N_21325,N_20357,N_20158);
xnor U21326 (N_21326,N_20838,N_20778);
or U21327 (N_21327,N_20202,N_20990);
nor U21328 (N_21328,N_20099,N_20310);
xor U21329 (N_21329,N_20490,N_20085);
nand U21330 (N_21330,N_20132,N_20220);
and U21331 (N_21331,N_20366,N_20259);
and U21332 (N_21332,N_20141,N_20856);
nor U21333 (N_21333,N_20441,N_20195);
and U21334 (N_21334,N_20540,N_20817);
and U21335 (N_21335,N_20686,N_20137);
nand U21336 (N_21336,N_20634,N_20859);
or U21337 (N_21337,N_20789,N_20956);
xor U21338 (N_21338,N_20011,N_20651);
and U21339 (N_21339,N_20319,N_20484);
or U21340 (N_21340,N_20959,N_20483);
and U21341 (N_21341,N_20915,N_20981);
nor U21342 (N_21342,N_20159,N_20828);
xnor U21343 (N_21343,N_20179,N_20624);
nor U21344 (N_21344,N_20059,N_20513);
and U21345 (N_21345,N_20027,N_20872);
nor U21346 (N_21346,N_20127,N_20387);
nand U21347 (N_21347,N_20560,N_20182);
and U21348 (N_21348,N_20665,N_20280);
nand U21349 (N_21349,N_20736,N_20679);
or U21350 (N_21350,N_20712,N_20234);
or U21351 (N_21351,N_20453,N_20122);
nor U21352 (N_21352,N_20893,N_20187);
xor U21353 (N_21353,N_20239,N_20213);
or U21354 (N_21354,N_20613,N_20649);
xnor U21355 (N_21355,N_20617,N_20205);
or U21356 (N_21356,N_20689,N_20069);
nor U21357 (N_21357,N_20955,N_20922);
xnor U21358 (N_21358,N_20477,N_20332);
and U21359 (N_21359,N_20511,N_20456);
and U21360 (N_21360,N_20768,N_20629);
xnor U21361 (N_21361,N_20347,N_20758);
nor U21362 (N_21362,N_20452,N_20932);
and U21363 (N_21363,N_20070,N_20218);
or U21364 (N_21364,N_20208,N_20802);
nand U21365 (N_21365,N_20056,N_20992);
or U21366 (N_21366,N_20078,N_20253);
xor U21367 (N_21367,N_20821,N_20261);
nor U21368 (N_21368,N_20976,N_20391);
and U21369 (N_21369,N_20865,N_20897);
or U21370 (N_21370,N_20994,N_20212);
and U21371 (N_21371,N_20790,N_20934);
or U21372 (N_21372,N_20050,N_20886);
and U21373 (N_21373,N_20162,N_20529);
nor U21374 (N_21374,N_20320,N_20427);
nor U21375 (N_21375,N_20274,N_20224);
nand U21376 (N_21376,N_20462,N_20696);
nor U21377 (N_21377,N_20619,N_20232);
nand U21378 (N_21378,N_20728,N_20243);
and U21379 (N_21379,N_20408,N_20359);
or U21380 (N_21380,N_20656,N_20655);
nor U21381 (N_21381,N_20049,N_20751);
or U21382 (N_21382,N_20426,N_20342);
nor U21383 (N_21383,N_20945,N_20433);
or U21384 (N_21384,N_20190,N_20416);
and U21385 (N_21385,N_20607,N_20832);
and U21386 (N_21386,N_20906,N_20194);
nand U21387 (N_21387,N_20356,N_20993);
nor U21388 (N_21388,N_20609,N_20524);
nand U21389 (N_21389,N_20943,N_20472);
or U21390 (N_21390,N_20596,N_20437);
nor U21391 (N_21391,N_20681,N_20957);
and U21392 (N_21392,N_20648,N_20903);
and U21393 (N_21393,N_20028,N_20283);
or U21394 (N_21394,N_20564,N_20038);
or U21395 (N_21395,N_20367,N_20471);
nand U21396 (N_21396,N_20797,N_20966);
nand U21397 (N_21397,N_20178,N_20952);
and U21398 (N_21398,N_20812,N_20855);
and U21399 (N_21399,N_20386,N_20503);
xnor U21400 (N_21400,N_20098,N_20512);
nand U21401 (N_21401,N_20382,N_20501);
nor U21402 (N_21402,N_20463,N_20863);
nor U21403 (N_21403,N_20740,N_20549);
xor U21404 (N_21404,N_20017,N_20404);
nor U21405 (N_21405,N_20774,N_20097);
nor U21406 (N_21406,N_20343,N_20002);
nand U21407 (N_21407,N_20101,N_20496);
xor U21408 (N_21408,N_20738,N_20126);
nor U21409 (N_21409,N_20643,N_20156);
nand U21410 (N_21410,N_20687,N_20801);
nand U21411 (N_21411,N_20900,N_20722);
and U21412 (N_21412,N_20969,N_20063);
xor U21413 (N_21413,N_20568,N_20374);
or U21414 (N_21414,N_20429,N_20358);
nor U21415 (N_21415,N_20614,N_20051);
nand U21416 (N_21416,N_20548,N_20258);
nor U21417 (N_21417,N_20939,N_20546);
nand U21418 (N_21418,N_20369,N_20565);
xor U21419 (N_21419,N_20094,N_20818);
or U21420 (N_21420,N_20024,N_20674);
nor U21421 (N_21421,N_20349,N_20898);
nor U21422 (N_21422,N_20831,N_20241);
xor U21423 (N_21423,N_20710,N_20166);
nand U21424 (N_21424,N_20533,N_20989);
and U21425 (N_21425,N_20065,N_20584);
or U21426 (N_21426,N_20523,N_20207);
xor U21427 (N_21427,N_20170,N_20591);
nand U21428 (N_21428,N_20419,N_20355);
nor U21429 (N_21429,N_20431,N_20891);
nor U21430 (N_21430,N_20394,N_20535);
and U21431 (N_21431,N_20216,N_20052);
xnor U21432 (N_21432,N_20446,N_20522);
nand U21433 (N_21433,N_20516,N_20398);
nand U21434 (N_21434,N_20530,N_20919);
or U21435 (N_21435,N_20423,N_20645);
nor U21436 (N_21436,N_20755,N_20291);
nor U21437 (N_21437,N_20435,N_20124);
nand U21438 (N_21438,N_20023,N_20455);
and U21439 (N_21439,N_20688,N_20168);
or U21440 (N_21440,N_20839,N_20739);
and U21441 (N_21441,N_20296,N_20003);
or U21442 (N_21442,N_20492,N_20400);
nor U21443 (N_21443,N_20805,N_20339);
and U21444 (N_21444,N_20771,N_20282);
nor U21445 (N_21445,N_20659,N_20804);
xnor U21446 (N_21446,N_20160,N_20824);
and U21447 (N_21447,N_20826,N_20896);
and U21448 (N_21448,N_20558,N_20620);
xnor U21449 (N_21449,N_20669,N_20372);
or U21450 (N_21450,N_20083,N_20365);
xnor U21451 (N_21451,N_20732,N_20515);
nor U21452 (N_21452,N_20593,N_20067);
xor U21453 (N_21453,N_20315,N_20018);
and U21454 (N_21454,N_20430,N_20075);
xnor U21455 (N_21455,N_20861,N_20585);
and U21456 (N_21456,N_20238,N_20779);
nand U21457 (N_21457,N_20829,N_20587);
nand U21458 (N_21458,N_20196,N_20589);
nand U21459 (N_21459,N_20979,N_20983);
nor U21460 (N_21460,N_20927,N_20760);
xor U21461 (N_21461,N_20963,N_20077);
and U21462 (N_21462,N_20109,N_20663);
nand U21463 (N_21463,N_20451,N_20727);
nor U21464 (N_21464,N_20371,N_20653);
or U21465 (N_21465,N_20481,N_20544);
and U21466 (N_21466,N_20662,N_20702);
nand U21467 (N_21467,N_20505,N_20608);
nor U21468 (N_21468,N_20250,N_20580);
and U21469 (N_21469,N_20198,N_20226);
nand U21470 (N_21470,N_20666,N_20393);
nor U21471 (N_21471,N_20970,N_20120);
xor U21472 (N_21472,N_20517,N_20345);
xnor U21473 (N_21473,N_20860,N_20631);
nor U21474 (N_21474,N_20953,N_20690);
nor U21475 (N_21475,N_20362,N_20658);
nand U21476 (N_21476,N_20072,N_20079);
xor U21477 (N_21477,N_20551,N_20814);
nand U21478 (N_21478,N_20555,N_20917);
xnor U21479 (N_21479,N_20594,N_20436);
nor U21480 (N_21480,N_20794,N_20671);
or U21481 (N_21481,N_20353,N_20869);
and U21482 (N_21482,N_20646,N_20909);
nor U21483 (N_21483,N_20428,N_20048);
nand U21484 (N_21484,N_20975,N_20996);
or U21485 (N_21485,N_20776,N_20485);
nand U21486 (N_21486,N_20364,N_20081);
nand U21487 (N_21487,N_20457,N_20348);
nor U21488 (N_21488,N_20150,N_20114);
nand U21489 (N_21489,N_20309,N_20892);
or U21490 (N_21490,N_20847,N_20113);
nor U21491 (N_21491,N_20222,N_20323);
and U21492 (N_21492,N_20325,N_20719);
and U21493 (N_21493,N_20765,N_20510);
nor U21494 (N_21494,N_20519,N_20105);
and U21495 (N_21495,N_20029,N_20901);
nor U21496 (N_21496,N_20192,N_20130);
and U21497 (N_21497,N_20145,N_20698);
and U21498 (N_21498,N_20193,N_20545);
and U21499 (N_21499,N_20344,N_20773);
or U21500 (N_21500,N_20505,N_20534);
or U21501 (N_21501,N_20000,N_20764);
or U21502 (N_21502,N_20904,N_20355);
or U21503 (N_21503,N_20852,N_20421);
nor U21504 (N_21504,N_20653,N_20806);
nor U21505 (N_21505,N_20498,N_20653);
or U21506 (N_21506,N_20339,N_20636);
or U21507 (N_21507,N_20597,N_20031);
nand U21508 (N_21508,N_20557,N_20192);
or U21509 (N_21509,N_20810,N_20785);
and U21510 (N_21510,N_20383,N_20473);
or U21511 (N_21511,N_20521,N_20140);
xor U21512 (N_21512,N_20402,N_20167);
nand U21513 (N_21513,N_20335,N_20750);
and U21514 (N_21514,N_20635,N_20040);
nor U21515 (N_21515,N_20811,N_20301);
and U21516 (N_21516,N_20997,N_20751);
and U21517 (N_21517,N_20881,N_20807);
nand U21518 (N_21518,N_20770,N_20222);
and U21519 (N_21519,N_20246,N_20644);
or U21520 (N_21520,N_20316,N_20000);
xor U21521 (N_21521,N_20184,N_20560);
and U21522 (N_21522,N_20421,N_20096);
or U21523 (N_21523,N_20618,N_20871);
nand U21524 (N_21524,N_20056,N_20113);
or U21525 (N_21525,N_20760,N_20634);
nand U21526 (N_21526,N_20287,N_20294);
and U21527 (N_21527,N_20593,N_20693);
xor U21528 (N_21528,N_20061,N_20841);
or U21529 (N_21529,N_20658,N_20305);
and U21530 (N_21530,N_20635,N_20921);
nor U21531 (N_21531,N_20393,N_20986);
or U21532 (N_21532,N_20321,N_20239);
xor U21533 (N_21533,N_20190,N_20732);
or U21534 (N_21534,N_20024,N_20197);
nand U21535 (N_21535,N_20791,N_20142);
xor U21536 (N_21536,N_20357,N_20855);
xnor U21537 (N_21537,N_20361,N_20380);
or U21538 (N_21538,N_20225,N_20849);
nand U21539 (N_21539,N_20198,N_20493);
and U21540 (N_21540,N_20531,N_20871);
xnor U21541 (N_21541,N_20224,N_20058);
or U21542 (N_21542,N_20647,N_20219);
and U21543 (N_21543,N_20036,N_20170);
nor U21544 (N_21544,N_20309,N_20923);
or U21545 (N_21545,N_20809,N_20463);
or U21546 (N_21546,N_20440,N_20342);
or U21547 (N_21547,N_20550,N_20252);
nor U21548 (N_21548,N_20441,N_20229);
nor U21549 (N_21549,N_20534,N_20019);
xor U21550 (N_21550,N_20765,N_20737);
and U21551 (N_21551,N_20681,N_20602);
xnor U21552 (N_21552,N_20799,N_20981);
or U21553 (N_21553,N_20086,N_20874);
nor U21554 (N_21554,N_20437,N_20143);
and U21555 (N_21555,N_20518,N_20190);
nand U21556 (N_21556,N_20036,N_20482);
or U21557 (N_21557,N_20437,N_20058);
nand U21558 (N_21558,N_20630,N_20048);
nand U21559 (N_21559,N_20117,N_20987);
or U21560 (N_21560,N_20359,N_20960);
or U21561 (N_21561,N_20258,N_20979);
and U21562 (N_21562,N_20170,N_20909);
nand U21563 (N_21563,N_20539,N_20376);
nor U21564 (N_21564,N_20725,N_20548);
xnor U21565 (N_21565,N_20543,N_20160);
and U21566 (N_21566,N_20582,N_20175);
or U21567 (N_21567,N_20269,N_20380);
or U21568 (N_21568,N_20056,N_20415);
xor U21569 (N_21569,N_20302,N_20005);
nand U21570 (N_21570,N_20037,N_20977);
nor U21571 (N_21571,N_20659,N_20833);
nor U21572 (N_21572,N_20064,N_20496);
nand U21573 (N_21573,N_20250,N_20310);
nand U21574 (N_21574,N_20870,N_20701);
or U21575 (N_21575,N_20613,N_20269);
nand U21576 (N_21576,N_20833,N_20031);
or U21577 (N_21577,N_20346,N_20455);
nor U21578 (N_21578,N_20728,N_20557);
xor U21579 (N_21579,N_20374,N_20737);
nor U21580 (N_21580,N_20853,N_20329);
or U21581 (N_21581,N_20715,N_20859);
nand U21582 (N_21582,N_20279,N_20941);
nor U21583 (N_21583,N_20469,N_20748);
or U21584 (N_21584,N_20427,N_20387);
xnor U21585 (N_21585,N_20895,N_20007);
and U21586 (N_21586,N_20844,N_20227);
or U21587 (N_21587,N_20948,N_20556);
and U21588 (N_21588,N_20332,N_20007);
nor U21589 (N_21589,N_20776,N_20244);
xor U21590 (N_21590,N_20403,N_20707);
and U21591 (N_21591,N_20208,N_20680);
nor U21592 (N_21592,N_20672,N_20822);
xnor U21593 (N_21593,N_20226,N_20141);
xor U21594 (N_21594,N_20718,N_20554);
or U21595 (N_21595,N_20335,N_20614);
and U21596 (N_21596,N_20082,N_20754);
and U21597 (N_21597,N_20482,N_20775);
nand U21598 (N_21598,N_20462,N_20421);
nand U21599 (N_21599,N_20787,N_20703);
nor U21600 (N_21600,N_20941,N_20231);
and U21601 (N_21601,N_20961,N_20627);
and U21602 (N_21602,N_20476,N_20338);
or U21603 (N_21603,N_20222,N_20138);
or U21604 (N_21604,N_20045,N_20371);
nor U21605 (N_21605,N_20387,N_20679);
nand U21606 (N_21606,N_20190,N_20906);
and U21607 (N_21607,N_20694,N_20195);
xor U21608 (N_21608,N_20684,N_20934);
xnor U21609 (N_21609,N_20789,N_20008);
xor U21610 (N_21610,N_20832,N_20187);
and U21611 (N_21611,N_20693,N_20103);
or U21612 (N_21612,N_20213,N_20544);
nand U21613 (N_21613,N_20795,N_20996);
and U21614 (N_21614,N_20520,N_20286);
xor U21615 (N_21615,N_20127,N_20818);
or U21616 (N_21616,N_20814,N_20818);
nor U21617 (N_21617,N_20754,N_20119);
xor U21618 (N_21618,N_20004,N_20726);
xor U21619 (N_21619,N_20508,N_20754);
and U21620 (N_21620,N_20464,N_20983);
and U21621 (N_21621,N_20274,N_20188);
nand U21622 (N_21622,N_20826,N_20780);
nor U21623 (N_21623,N_20222,N_20598);
and U21624 (N_21624,N_20951,N_20005);
nand U21625 (N_21625,N_20845,N_20640);
xor U21626 (N_21626,N_20909,N_20991);
xnor U21627 (N_21627,N_20992,N_20946);
and U21628 (N_21628,N_20841,N_20075);
xnor U21629 (N_21629,N_20273,N_20248);
and U21630 (N_21630,N_20195,N_20162);
or U21631 (N_21631,N_20484,N_20638);
xor U21632 (N_21632,N_20368,N_20667);
or U21633 (N_21633,N_20663,N_20479);
and U21634 (N_21634,N_20398,N_20570);
nand U21635 (N_21635,N_20132,N_20473);
and U21636 (N_21636,N_20354,N_20404);
nor U21637 (N_21637,N_20132,N_20502);
and U21638 (N_21638,N_20308,N_20095);
nand U21639 (N_21639,N_20657,N_20669);
or U21640 (N_21640,N_20861,N_20452);
nand U21641 (N_21641,N_20908,N_20061);
nand U21642 (N_21642,N_20860,N_20103);
xor U21643 (N_21643,N_20707,N_20030);
nand U21644 (N_21644,N_20414,N_20886);
nor U21645 (N_21645,N_20501,N_20945);
or U21646 (N_21646,N_20564,N_20709);
xnor U21647 (N_21647,N_20391,N_20597);
nor U21648 (N_21648,N_20914,N_20601);
and U21649 (N_21649,N_20009,N_20561);
xnor U21650 (N_21650,N_20452,N_20244);
nor U21651 (N_21651,N_20748,N_20518);
xor U21652 (N_21652,N_20566,N_20950);
and U21653 (N_21653,N_20008,N_20692);
nor U21654 (N_21654,N_20907,N_20211);
or U21655 (N_21655,N_20577,N_20225);
nand U21656 (N_21656,N_20169,N_20277);
and U21657 (N_21657,N_20452,N_20745);
nand U21658 (N_21658,N_20794,N_20922);
xor U21659 (N_21659,N_20576,N_20598);
and U21660 (N_21660,N_20434,N_20054);
xnor U21661 (N_21661,N_20003,N_20065);
nor U21662 (N_21662,N_20720,N_20522);
nor U21663 (N_21663,N_20711,N_20103);
nor U21664 (N_21664,N_20688,N_20769);
and U21665 (N_21665,N_20154,N_20186);
nor U21666 (N_21666,N_20135,N_20334);
or U21667 (N_21667,N_20256,N_20984);
nor U21668 (N_21668,N_20796,N_20019);
xor U21669 (N_21669,N_20845,N_20533);
nor U21670 (N_21670,N_20155,N_20782);
and U21671 (N_21671,N_20070,N_20637);
or U21672 (N_21672,N_20132,N_20655);
nand U21673 (N_21673,N_20107,N_20574);
xor U21674 (N_21674,N_20002,N_20933);
and U21675 (N_21675,N_20847,N_20318);
nor U21676 (N_21676,N_20709,N_20340);
and U21677 (N_21677,N_20440,N_20674);
nor U21678 (N_21678,N_20160,N_20722);
or U21679 (N_21679,N_20442,N_20796);
nor U21680 (N_21680,N_20201,N_20373);
nand U21681 (N_21681,N_20393,N_20293);
nand U21682 (N_21682,N_20863,N_20196);
nand U21683 (N_21683,N_20392,N_20871);
nand U21684 (N_21684,N_20788,N_20647);
nand U21685 (N_21685,N_20162,N_20775);
nand U21686 (N_21686,N_20516,N_20237);
nand U21687 (N_21687,N_20686,N_20272);
nor U21688 (N_21688,N_20975,N_20816);
and U21689 (N_21689,N_20221,N_20767);
nor U21690 (N_21690,N_20023,N_20561);
and U21691 (N_21691,N_20937,N_20912);
xnor U21692 (N_21692,N_20848,N_20039);
xor U21693 (N_21693,N_20080,N_20655);
nand U21694 (N_21694,N_20670,N_20431);
nand U21695 (N_21695,N_20498,N_20650);
nand U21696 (N_21696,N_20185,N_20432);
nand U21697 (N_21697,N_20049,N_20438);
xor U21698 (N_21698,N_20370,N_20996);
nand U21699 (N_21699,N_20164,N_20286);
nand U21700 (N_21700,N_20440,N_20117);
nor U21701 (N_21701,N_20446,N_20544);
nor U21702 (N_21702,N_20306,N_20389);
and U21703 (N_21703,N_20788,N_20081);
nor U21704 (N_21704,N_20086,N_20922);
xnor U21705 (N_21705,N_20798,N_20257);
xnor U21706 (N_21706,N_20733,N_20049);
xnor U21707 (N_21707,N_20318,N_20678);
and U21708 (N_21708,N_20504,N_20770);
nand U21709 (N_21709,N_20533,N_20140);
nor U21710 (N_21710,N_20740,N_20555);
nand U21711 (N_21711,N_20773,N_20733);
xnor U21712 (N_21712,N_20304,N_20506);
nor U21713 (N_21713,N_20265,N_20883);
xor U21714 (N_21714,N_20131,N_20379);
nand U21715 (N_21715,N_20017,N_20747);
or U21716 (N_21716,N_20321,N_20912);
xnor U21717 (N_21717,N_20016,N_20675);
nor U21718 (N_21718,N_20256,N_20464);
or U21719 (N_21719,N_20729,N_20995);
xor U21720 (N_21720,N_20605,N_20566);
nor U21721 (N_21721,N_20130,N_20555);
nand U21722 (N_21722,N_20927,N_20951);
nor U21723 (N_21723,N_20263,N_20968);
nand U21724 (N_21724,N_20406,N_20397);
and U21725 (N_21725,N_20106,N_20385);
nor U21726 (N_21726,N_20140,N_20760);
or U21727 (N_21727,N_20593,N_20156);
or U21728 (N_21728,N_20883,N_20055);
nand U21729 (N_21729,N_20065,N_20484);
xor U21730 (N_21730,N_20251,N_20400);
nand U21731 (N_21731,N_20934,N_20678);
or U21732 (N_21732,N_20418,N_20497);
or U21733 (N_21733,N_20477,N_20336);
and U21734 (N_21734,N_20674,N_20358);
xor U21735 (N_21735,N_20274,N_20635);
or U21736 (N_21736,N_20359,N_20872);
nor U21737 (N_21737,N_20291,N_20729);
and U21738 (N_21738,N_20042,N_20145);
xnor U21739 (N_21739,N_20640,N_20714);
xnor U21740 (N_21740,N_20411,N_20462);
and U21741 (N_21741,N_20034,N_20503);
xnor U21742 (N_21742,N_20984,N_20138);
xor U21743 (N_21743,N_20358,N_20265);
nor U21744 (N_21744,N_20178,N_20447);
nand U21745 (N_21745,N_20492,N_20378);
and U21746 (N_21746,N_20623,N_20313);
xor U21747 (N_21747,N_20678,N_20569);
nand U21748 (N_21748,N_20955,N_20340);
xor U21749 (N_21749,N_20535,N_20668);
and U21750 (N_21750,N_20043,N_20851);
xnor U21751 (N_21751,N_20955,N_20239);
nor U21752 (N_21752,N_20020,N_20575);
xnor U21753 (N_21753,N_20167,N_20589);
or U21754 (N_21754,N_20761,N_20307);
or U21755 (N_21755,N_20171,N_20362);
or U21756 (N_21756,N_20861,N_20359);
or U21757 (N_21757,N_20761,N_20738);
xor U21758 (N_21758,N_20323,N_20111);
xnor U21759 (N_21759,N_20318,N_20754);
nand U21760 (N_21760,N_20694,N_20342);
xor U21761 (N_21761,N_20063,N_20639);
and U21762 (N_21762,N_20567,N_20372);
nand U21763 (N_21763,N_20061,N_20356);
nand U21764 (N_21764,N_20383,N_20436);
nand U21765 (N_21765,N_20405,N_20483);
nand U21766 (N_21766,N_20537,N_20447);
and U21767 (N_21767,N_20480,N_20761);
nor U21768 (N_21768,N_20128,N_20605);
xnor U21769 (N_21769,N_20289,N_20118);
nor U21770 (N_21770,N_20662,N_20616);
nor U21771 (N_21771,N_20148,N_20410);
or U21772 (N_21772,N_20540,N_20959);
and U21773 (N_21773,N_20711,N_20227);
and U21774 (N_21774,N_20524,N_20666);
nor U21775 (N_21775,N_20982,N_20540);
or U21776 (N_21776,N_20942,N_20963);
and U21777 (N_21777,N_20028,N_20831);
nor U21778 (N_21778,N_20434,N_20622);
xnor U21779 (N_21779,N_20819,N_20432);
or U21780 (N_21780,N_20341,N_20387);
nand U21781 (N_21781,N_20541,N_20055);
and U21782 (N_21782,N_20131,N_20410);
or U21783 (N_21783,N_20934,N_20364);
and U21784 (N_21784,N_20739,N_20730);
and U21785 (N_21785,N_20660,N_20591);
nand U21786 (N_21786,N_20428,N_20193);
nand U21787 (N_21787,N_20539,N_20154);
nand U21788 (N_21788,N_20336,N_20551);
or U21789 (N_21789,N_20859,N_20975);
xnor U21790 (N_21790,N_20199,N_20331);
nand U21791 (N_21791,N_20686,N_20719);
nand U21792 (N_21792,N_20852,N_20727);
xnor U21793 (N_21793,N_20847,N_20008);
and U21794 (N_21794,N_20430,N_20500);
nand U21795 (N_21795,N_20733,N_20077);
and U21796 (N_21796,N_20994,N_20746);
and U21797 (N_21797,N_20430,N_20284);
xnor U21798 (N_21798,N_20080,N_20796);
nand U21799 (N_21799,N_20637,N_20892);
nand U21800 (N_21800,N_20932,N_20880);
nor U21801 (N_21801,N_20985,N_20656);
and U21802 (N_21802,N_20855,N_20140);
and U21803 (N_21803,N_20004,N_20375);
and U21804 (N_21804,N_20585,N_20165);
or U21805 (N_21805,N_20509,N_20052);
and U21806 (N_21806,N_20518,N_20221);
nand U21807 (N_21807,N_20843,N_20494);
nand U21808 (N_21808,N_20680,N_20164);
nor U21809 (N_21809,N_20378,N_20719);
and U21810 (N_21810,N_20094,N_20679);
nor U21811 (N_21811,N_20258,N_20831);
xor U21812 (N_21812,N_20581,N_20913);
nor U21813 (N_21813,N_20926,N_20198);
xor U21814 (N_21814,N_20140,N_20431);
nor U21815 (N_21815,N_20620,N_20955);
nor U21816 (N_21816,N_20175,N_20928);
xor U21817 (N_21817,N_20380,N_20600);
nand U21818 (N_21818,N_20073,N_20831);
nor U21819 (N_21819,N_20373,N_20352);
nand U21820 (N_21820,N_20933,N_20160);
xnor U21821 (N_21821,N_20443,N_20226);
and U21822 (N_21822,N_20160,N_20643);
nand U21823 (N_21823,N_20309,N_20082);
nand U21824 (N_21824,N_20057,N_20224);
nor U21825 (N_21825,N_20685,N_20483);
and U21826 (N_21826,N_20916,N_20877);
and U21827 (N_21827,N_20847,N_20526);
nand U21828 (N_21828,N_20478,N_20058);
or U21829 (N_21829,N_20538,N_20901);
or U21830 (N_21830,N_20165,N_20397);
xnor U21831 (N_21831,N_20642,N_20449);
xnor U21832 (N_21832,N_20588,N_20314);
nand U21833 (N_21833,N_20703,N_20025);
xor U21834 (N_21834,N_20696,N_20666);
nand U21835 (N_21835,N_20183,N_20568);
nand U21836 (N_21836,N_20234,N_20107);
and U21837 (N_21837,N_20057,N_20327);
nand U21838 (N_21838,N_20096,N_20478);
nand U21839 (N_21839,N_20260,N_20195);
and U21840 (N_21840,N_20940,N_20318);
xor U21841 (N_21841,N_20827,N_20260);
and U21842 (N_21842,N_20380,N_20604);
and U21843 (N_21843,N_20587,N_20306);
or U21844 (N_21844,N_20487,N_20526);
or U21845 (N_21845,N_20109,N_20050);
nand U21846 (N_21846,N_20524,N_20619);
and U21847 (N_21847,N_20124,N_20448);
nand U21848 (N_21848,N_20003,N_20255);
and U21849 (N_21849,N_20655,N_20930);
and U21850 (N_21850,N_20913,N_20250);
nor U21851 (N_21851,N_20588,N_20232);
nor U21852 (N_21852,N_20067,N_20703);
nor U21853 (N_21853,N_20386,N_20732);
xnor U21854 (N_21854,N_20339,N_20162);
nand U21855 (N_21855,N_20983,N_20744);
nand U21856 (N_21856,N_20456,N_20998);
and U21857 (N_21857,N_20364,N_20953);
and U21858 (N_21858,N_20288,N_20524);
nor U21859 (N_21859,N_20163,N_20457);
and U21860 (N_21860,N_20472,N_20065);
nor U21861 (N_21861,N_20541,N_20675);
xor U21862 (N_21862,N_20846,N_20682);
and U21863 (N_21863,N_20928,N_20680);
or U21864 (N_21864,N_20970,N_20598);
nor U21865 (N_21865,N_20193,N_20874);
or U21866 (N_21866,N_20964,N_20417);
nor U21867 (N_21867,N_20856,N_20619);
and U21868 (N_21868,N_20714,N_20742);
xnor U21869 (N_21869,N_20733,N_20446);
and U21870 (N_21870,N_20440,N_20248);
xor U21871 (N_21871,N_20050,N_20368);
xor U21872 (N_21872,N_20211,N_20377);
nor U21873 (N_21873,N_20237,N_20575);
nor U21874 (N_21874,N_20287,N_20010);
nor U21875 (N_21875,N_20467,N_20190);
and U21876 (N_21876,N_20493,N_20829);
xnor U21877 (N_21877,N_20816,N_20630);
nand U21878 (N_21878,N_20610,N_20543);
and U21879 (N_21879,N_20509,N_20304);
and U21880 (N_21880,N_20442,N_20762);
nand U21881 (N_21881,N_20223,N_20309);
or U21882 (N_21882,N_20432,N_20004);
nand U21883 (N_21883,N_20972,N_20063);
nor U21884 (N_21884,N_20581,N_20772);
xor U21885 (N_21885,N_20685,N_20506);
nand U21886 (N_21886,N_20211,N_20303);
nand U21887 (N_21887,N_20399,N_20683);
nand U21888 (N_21888,N_20123,N_20330);
and U21889 (N_21889,N_20623,N_20180);
and U21890 (N_21890,N_20352,N_20585);
xnor U21891 (N_21891,N_20404,N_20550);
xnor U21892 (N_21892,N_20131,N_20479);
xor U21893 (N_21893,N_20463,N_20590);
nor U21894 (N_21894,N_20792,N_20941);
and U21895 (N_21895,N_20494,N_20275);
nor U21896 (N_21896,N_20260,N_20325);
or U21897 (N_21897,N_20046,N_20967);
nor U21898 (N_21898,N_20140,N_20802);
nor U21899 (N_21899,N_20824,N_20390);
xnor U21900 (N_21900,N_20795,N_20820);
or U21901 (N_21901,N_20627,N_20613);
xor U21902 (N_21902,N_20915,N_20330);
nand U21903 (N_21903,N_20291,N_20336);
or U21904 (N_21904,N_20127,N_20506);
nor U21905 (N_21905,N_20007,N_20802);
and U21906 (N_21906,N_20147,N_20264);
xor U21907 (N_21907,N_20573,N_20710);
nor U21908 (N_21908,N_20186,N_20600);
nor U21909 (N_21909,N_20943,N_20283);
nor U21910 (N_21910,N_20989,N_20011);
or U21911 (N_21911,N_20796,N_20296);
or U21912 (N_21912,N_20849,N_20485);
and U21913 (N_21913,N_20596,N_20586);
nor U21914 (N_21914,N_20385,N_20058);
xor U21915 (N_21915,N_20864,N_20791);
or U21916 (N_21916,N_20433,N_20810);
xnor U21917 (N_21917,N_20557,N_20599);
nor U21918 (N_21918,N_20668,N_20806);
nand U21919 (N_21919,N_20503,N_20498);
or U21920 (N_21920,N_20031,N_20002);
nand U21921 (N_21921,N_20907,N_20731);
nor U21922 (N_21922,N_20256,N_20713);
nor U21923 (N_21923,N_20606,N_20511);
nand U21924 (N_21924,N_20582,N_20585);
or U21925 (N_21925,N_20170,N_20837);
or U21926 (N_21926,N_20109,N_20146);
nor U21927 (N_21927,N_20131,N_20680);
nor U21928 (N_21928,N_20048,N_20252);
or U21929 (N_21929,N_20880,N_20212);
and U21930 (N_21930,N_20520,N_20317);
and U21931 (N_21931,N_20525,N_20195);
nand U21932 (N_21932,N_20532,N_20150);
or U21933 (N_21933,N_20357,N_20199);
xor U21934 (N_21934,N_20176,N_20978);
nor U21935 (N_21935,N_20499,N_20154);
nand U21936 (N_21936,N_20795,N_20436);
nor U21937 (N_21937,N_20189,N_20499);
nand U21938 (N_21938,N_20260,N_20018);
xor U21939 (N_21939,N_20130,N_20662);
nand U21940 (N_21940,N_20949,N_20127);
or U21941 (N_21941,N_20846,N_20978);
or U21942 (N_21942,N_20490,N_20557);
nor U21943 (N_21943,N_20157,N_20826);
nor U21944 (N_21944,N_20292,N_20778);
nand U21945 (N_21945,N_20438,N_20462);
or U21946 (N_21946,N_20789,N_20627);
or U21947 (N_21947,N_20843,N_20880);
xnor U21948 (N_21948,N_20139,N_20589);
and U21949 (N_21949,N_20008,N_20925);
or U21950 (N_21950,N_20146,N_20481);
or U21951 (N_21951,N_20628,N_20591);
nand U21952 (N_21952,N_20309,N_20251);
and U21953 (N_21953,N_20614,N_20564);
nor U21954 (N_21954,N_20772,N_20964);
or U21955 (N_21955,N_20844,N_20395);
or U21956 (N_21956,N_20100,N_20465);
or U21957 (N_21957,N_20995,N_20036);
or U21958 (N_21958,N_20167,N_20085);
xnor U21959 (N_21959,N_20119,N_20927);
xnor U21960 (N_21960,N_20448,N_20132);
nor U21961 (N_21961,N_20330,N_20896);
nor U21962 (N_21962,N_20076,N_20947);
and U21963 (N_21963,N_20869,N_20103);
nand U21964 (N_21964,N_20140,N_20005);
nor U21965 (N_21965,N_20334,N_20837);
or U21966 (N_21966,N_20781,N_20038);
xnor U21967 (N_21967,N_20372,N_20720);
xnor U21968 (N_21968,N_20902,N_20949);
or U21969 (N_21969,N_20774,N_20059);
and U21970 (N_21970,N_20417,N_20032);
nor U21971 (N_21971,N_20010,N_20662);
and U21972 (N_21972,N_20172,N_20997);
nand U21973 (N_21973,N_20485,N_20528);
nor U21974 (N_21974,N_20116,N_20192);
nand U21975 (N_21975,N_20770,N_20508);
or U21976 (N_21976,N_20909,N_20534);
xnor U21977 (N_21977,N_20282,N_20065);
and U21978 (N_21978,N_20947,N_20498);
or U21979 (N_21979,N_20360,N_20966);
and U21980 (N_21980,N_20142,N_20301);
or U21981 (N_21981,N_20556,N_20963);
nor U21982 (N_21982,N_20936,N_20754);
nor U21983 (N_21983,N_20109,N_20210);
or U21984 (N_21984,N_20678,N_20009);
nor U21985 (N_21985,N_20713,N_20835);
nor U21986 (N_21986,N_20733,N_20539);
xnor U21987 (N_21987,N_20260,N_20746);
and U21988 (N_21988,N_20364,N_20112);
or U21989 (N_21989,N_20745,N_20923);
or U21990 (N_21990,N_20125,N_20237);
nand U21991 (N_21991,N_20658,N_20738);
or U21992 (N_21992,N_20452,N_20477);
nand U21993 (N_21993,N_20721,N_20473);
and U21994 (N_21994,N_20688,N_20648);
nand U21995 (N_21995,N_20505,N_20492);
or U21996 (N_21996,N_20448,N_20922);
or U21997 (N_21997,N_20425,N_20021);
or U21998 (N_21998,N_20724,N_20742);
nor U21999 (N_21999,N_20248,N_20317);
nand U22000 (N_22000,N_21211,N_21731);
and U22001 (N_22001,N_21702,N_21274);
nand U22002 (N_22002,N_21691,N_21002);
nand U22003 (N_22003,N_21737,N_21989);
nor U22004 (N_22004,N_21385,N_21161);
nor U22005 (N_22005,N_21828,N_21463);
and U22006 (N_22006,N_21452,N_21009);
nand U22007 (N_22007,N_21352,N_21842);
nor U22008 (N_22008,N_21992,N_21778);
xnor U22009 (N_22009,N_21602,N_21435);
and U22010 (N_22010,N_21649,N_21964);
or U22011 (N_22011,N_21894,N_21865);
nor U22012 (N_22012,N_21845,N_21835);
and U22013 (N_22013,N_21292,N_21119);
xnor U22014 (N_22014,N_21394,N_21508);
xnor U22015 (N_22015,N_21575,N_21182);
xor U22016 (N_22016,N_21882,N_21809);
and U22017 (N_22017,N_21539,N_21640);
and U22018 (N_22018,N_21355,N_21822);
and U22019 (N_22019,N_21062,N_21242);
nand U22020 (N_22020,N_21429,N_21227);
or U22021 (N_22021,N_21192,N_21499);
and U22022 (N_22022,N_21748,N_21843);
or U22023 (N_22023,N_21913,N_21909);
nand U22024 (N_22024,N_21545,N_21785);
nor U22025 (N_22025,N_21636,N_21250);
nor U22026 (N_22026,N_21346,N_21848);
nand U22027 (N_22027,N_21921,N_21807);
nand U22028 (N_22028,N_21726,N_21271);
nand U22029 (N_22029,N_21144,N_21003);
or U22030 (N_22030,N_21634,N_21162);
or U22031 (N_22031,N_21333,N_21998);
nor U22032 (N_22032,N_21163,N_21598);
nand U22033 (N_22033,N_21076,N_21485);
xnor U22034 (N_22034,N_21444,N_21969);
or U22035 (N_22035,N_21628,N_21241);
nor U22036 (N_22036,N_21120,N_21465);
and U22037 (N_22037,N_21732,N_21703);
nor U22038 (N_22038,N_21551,N_21688);
xor U22039 (N_22039,N_21072,N_21048);
nor U22040 (N_22040,N_21685,N_21949);
and U22041 (N_22041,N_21010,N_21087);
or U22042 (N_22042,N_21814,N_21191);
xor U22043 (N_22043,N_21523,N_21514);
nand U22044 (N_22044,N_21993,N_21826);
and U22045 (N_22045,N_21586,N_21771);
and U22046 (N_22046,N_21942,N_21692);
xnor U22047 (N_22047,N_21125,N_21859);
xor U22048 (N_22048,N_21321,N_21915);
nor U22049 (N_22049,N_21733,N_21312);
nand U22050 (N_22050,N_21900,N_21681);
nor U22051 (N_22051,N_21366,N_21092);
xor U22052 (N_22052,N_21089,N_21779);
xor U22053 (N_22053,N_21388,N_21565);
or U22054 (N_22054,N_21730,N_21212);
nand U22055 (N_22055,N_21777,N_21378);
nand U22056 (N_22056,N_21864,N_21559);
and U22057 (N_22057,N_21699,N_21364);
nor U22058 (N_22058,N_21108,N_21044);
xor U22059 (N_22059,N_21739,N_21392);
xor U22060 (N_22060,N_21275,N_21439);
nor U22061 (N_22061,N_21967,N_21888);
or U22062 (N_22062,N_21999,N_21493);
xor U22063 (N_22063,N_21898,N_21314);
or U22064 (N_22064,N_21566,N_21356);
and U22065 (N_22065,N_21955,N_21338);
nor U22066 (N_22066,N_21045,N_21047);
xnor U22067 (N_22067,N_21549,N_21766);
xnor U22068 (N_22068,N_21375,N_21976);
nor U22069 (N_22069,N_21391,N_21489);
or U22070 (N_22070,N_21324,N_21299);
or U22071 (N_22071,N_21742,N_21284);
xor U22072 (N_22072,N_21122,N_21660);
or U22073 (N_22073,N_21341,N_21094);
nand U22074 (N_22074,N_21610,N_21664);
and U22075 (N_22075,N_21446,N_21963);
nand U22076 (N_22076,N_21339,N_21676);
and U22077 (N_22077,N_21533,N_21831);
xor U22078 (N_22078,N_21247,N_21906);
nor U22079 (N_22079,N_21836,N_21400);
nor U22080 (N_22080,N_21436,N_21269);
nor U22081 (N_22081,N_21884,N_21220);
or U22082 (N_22082,N_21960,N_21368);
or U22083 (N_22083,N_21725,N_21957);
nand U22084 (N_22084,N_21103,N_21051);
and U22085 (N_22085,N_21153,N_21406);
and U22086 (N_22086,N_21187,N_21719);
nor U22087 (N_22087,N_21695,N_21986);
xnor U22088 (N_22088,N_21698,N_21880);
and U22089 (N_22089,N_21427,N_21421);
or U22090 (N_22090,N_21804,N_21905);
and U22091 (N_22091,N_21077,N_21308);
or U22092 (N_22092,N_21152,N_21000);
nand U22093 (N_22093,N_21277,N_21146);
nor U22094 (N_22094,N_21659,N_21530);
nand U22095 (N_22095,N_21064,N_21883);
and U22096 (N_22096,N_21040,N_21617);
or U22097 (N_22097,N_21768,N_21343);
and U22098 (N_22098,N_21154,N_21196);
or U22099 (N_22099,N_21399,N_21136);
nand U22100 (N_22100,N_21148,N_21524);
nor U22101 (N_22101,N_21395,N_21600);
and U22102 (N_22102,N_21408,N_21879);
or U22103 (N_22103,N_21177,N_21653);
xor U22104 (N_22104,N_21933,N_21684);
or U22105 (N_22105,N_21244,N_21816);
nor U22106 (N_22106,N_21607,N_21491);
nand U22107 (N_22107,N_21510,N_21556);
or U22108 (N_22108,N_21757,N_21431);
and U22109 (N_22109,N_21052,N_21025);
nor U22110 (N_22110,N_21801,N_21516);
or U22111 (N_22111,N_21226,N_21774);
nand U22112 (N_22112,N_21389,N_21145);
nand U22113 (N_22113,N_21380,N_21994);
or U22114 (N_22114,N_21576,N_21724);
or U22115 (N_22115,N_21522,N_21716);
nor U22116 (N_22116,N_21800,N_21334);
nor U22117 (N_22117,N_21150,N_21765);
xor U22118 (N_22118,N_21283,N_21759);
xor U22119 (N_22119,N_21167,N_21903);
or U22120 (N_22120,N_21796,N_21932);
or U22121 (N_22121,N_21371,N_21206);
and U22122 (N_22122,N_21142,N_21416);
and U22123 (N_22123,N_21892,N_21423);
or U22124 (N_22124,N_21643,N_21294);
or U22125 (N_22125,N_21877,N_21129);
xnor U22126 (N_22126,N_21024,N_21233);
xor U22127 (N_22127,N_21750,N_21793);
and U22128 (N_22128,N_21770,N_21488);
nor U22129 (N_22129,N_21840,N_21507);
xnor U22130 (N_22130,N_21131,N_21946);
and U22131 (N_22131,N_21708,N_21310);
nand U22132 (N_22132,N_21683,N_21678);
xor U22133 (N_22133,N_21173,N_21953);
nand U22134 (N_22134,N_21198,N_21056);
nand U22135 (N_22135,N_21783,N_21934);
xor U22136 (N_22136,N_21803,N_21020);
and U22137 (N_22137,N_21365,N_21904);
xnor U22138 (N_22138,N_21453,N_21004);
and U22139 (N_22139,N_21574,N_21581);
or U22140 (N_22140,N_21971,N_21528);
nor U22141 (N_22141,N_21571,N_21289);
or U22142 (N_22142,N_21509,N_21464);
and U22143 (N_22143,N_21591,N_21350);
nor U22144 (N_22144,N_21631,N_21318);
or U22145 (N_22145,N_21572,N_21332);
or U22146 (N_22146,N_21214,N_21582);
xnor U22147 (N_22147,N_21862,N_21068);
or U22148 (N_22148,N_21995,N_21797);
or U22149 (N_22149,N_21105,N_21029);
and U22150 (N_22150,N_21095,N_21078);
or U22151 (N_22151,N_21147,N_21336);
xor U22152 (N_22152,N_21449,N_21734);
nor U22153 (N_22153,N_21140,N_21867);
xnor U22154 (N_22154,N_21369,N_21937);
xnor U22155 (N_22155,N_21128,N_21956);
and U22156 (N_22156,N_21217,N_21966);
and U22157 (N_22157,N_21311,N_21305);
nor U22158 (N_22158,N_21601,N_21171);
xor U22159 (N_22159,N_21260,N_21419);
xnor U22160 (N_22160,N_21561,N_21032);
nor U22161 (N_22161,N_21023,N_21744);
nor U22162 (N_22162,N_21176,N_21902);
or U22163 (N_22163,N_21091,N_21172);
xnor U22164 (N_22164,N_21268,N_21330);
and U22165 (N_22165,N_21208,N_21001);
nor U22166 (N_22166,N_21914,N_21013);
or U22167 (N_22167,N_21614,N_21819);
nand U22168 (N_22168,N_21603,N_21353);
nand U22169 (N_22169,N_21362,N_21053);
nor U22170 (N_22170,N_21098,N_21124);
and U22171 (N_22171,N_21856,N_21972);
and U22172 (N_22172,N_21700,N_21276);
and U22173 (N_22173,N_21460,N_21457);
nor U22174 (N_22174,N_21074,N_21169);
nor U22175 (N_22175,N_21409,N_21039);
and U22176 (N_22176,N_21787,N_21805);
or U22177 (N_22177,N_21237,N_21199);
or U22178 (N_22178,N_21070,N_21526);
and U22179 (N_22179,N_21773,N_21629);
and U22180 (N_22180,N_21808,N_21492);
and U22181 (N_22181,N_21997,N_21912);
nand U22182 (N_22182,N_21181,N_21302);
xnor U22183 (N_22183,N_21065,N_21673);
nand U22184 (N_22184,N_21417,N_21531);
and U22185 (N_22185,N_21016,N_21962);
or U22186 (N_22186,N_21265,N_21975);
or U22187 (N_22187,N_21827,N_21296);
nand U22188 (N_22188,N_21207,N_21515);
nand U22189 (N_22189,N_21935,N_21623);
xnor U22190 (N_22190,N_21769,N_21030);
nand U22191 (N_22191,N_21981,N_21535);
and U22192 (N_22192,N_21511,N_21958);
xor U22193 (N_22193,N_21081,N_21890);
nor U22194 (N_22194,N_21301,N_21382);
nor U22195 (N_22195,N_21871,N_21767);
and U22196 (N_22196,N_21714,N_21841);
nor U22197 (N_22197,N_21459,N_21627);
and U22198 (N_22198,N_21749,N_21041);
nor U22199 (N_22199,N_21213,N_21677);
xor U22200 (N_22200,N_21430,N_21322);
nor U22201 (N_22201,N_21857,N_21420);
nor U22202 (N_22202,N_21323,N_21650);
or U22203 (N_22203,N_21616,N_21210);
or U22204 (N_22204,N_21319,N_21927);
nand U22205 (N_22205,N_21263,N_21126);
and U22206 (N_22206,N_21763,N_21735);
nand U22207 (N_22207,N_21118,N_21224);
nor U22208 (N_22208,N_21891,N_21548);
nand U22209 (N_22209,N_21589,N_21498);
xnor U22210 (N_22210,N_21156,N_21985);
or U22211 (N_22211,N_21878,N_21058);
nand U22212 (N_22212,N_21990,N_21258);
or U22213 (N_22213,N_21109,N_21069);
xnor U22214 (N_22214,N_21645,N_21007);
nor U22215 (N_22215,N_21943,N_21253);
xor U22216 (N_22216,N_21597,N_21799);
and U22217 (N_22217,N_21837,N_21448);
xnor U22218 (N_22218,N_21850,N_21741);
xnor U22219 (N_22219,N_21520,N_21722);
nor U22220 (N_22220,N_21893,N_21205);
nand U22221 (N_22221,N_21709,N_21428);
and U22222 (N_22222,N_21854,N_21647);
and U22223 (N_22223,N_21049,N_21811);
xnor U22224 (N_22224,N_21521,N_21021);
xor U22225 (N_22225,N_21386,N_21916);
nand U22226 (N_22226,N_21736,N_21036);
xor U22227 (N_22227,N_21656,N_21063);
or U22228 (N_22228,N_21588,N_21760);
nand U22229 (N_22229,N_21578,N_21690);
and U22230 (N_22230,N_21279,N_21505);
nand U22231 (N_22231,N_21746,N_21151);
nand U22232 (N_22232,N_21222,N_21849);
xor U22233 (N_22233,N_21495,N_21223);
and U22234 (N_22234,N_21978,N_21675);
nand U22235 (N_22235,N_21789,N_21954);
and U22236 (N_22236,N_21562,N_21861);
nand U22237 (N_22237,N_21357,N_21221);
xor U22238 (N_22238,N_21812,N_21335);
nor U22239 (N_22239,N_21328,N_21924);
and U22240 (N_22240,N_21107,N_21740);
nand U22241 (N_22241,N_21537,N_21345);
nor U22242 (N_22242,N_21689,N_21249);
nor U22243 (N_22243,N_21866,N_21494);
and U22244 (N_22244,N_21821,N_21829);
and U22245 (N_22245,N_21824,N_21729);
or U22246 (N_22246,N_21133,N_21300);
nor U22247 (N_22247,N_21547,N_21846);
or U22248 (N_22248,N_21433,N_21544);
nand U22249 (N_22249,N_21863,N_21974);
and U22250 (N_22250,N_21424,N_21868);
nand U22251 (N_22251,N_21473,N_21928);
nor U22252 (N_22252,N_21286,N_21686);
nor U22253 (N_22253,N_21102,N_21360);
or U22254 (N_22254,N_21847,N_21178);
and U22255 (N_22255,N_21679,N_21784);
and U22256 (N_22256,N_21006,N_21504);
nand U22257 (N_22257,N_21349,N_21374);
and U22258 (N_22258,N_21272,N_21813);
and U22259 (N_22259,N_21232,N_21104);
nand U22260 (N_22260,N_21633,N_21996);
nand U22261 (N_22261,N_21758,N_21099);
nand U22262 (N_22262,N_21306,N_21968);
xor U22263 (N_22263,N_21980,N_21037);
or U22264 (N_22264,N_21327,N_21550);
xnor U22265 (N_22265,N_21390,N_21005);
or U22266 (N_22266,N_21480,N_21387);
and U22267 (N_22267,N_21209,N_21532);
nand U22268 (N_22268,N_21644,N_21938);
or U22269 (N_22269,N_21573,N_21881);
nor U22270 (N_22270,N_21101,N_21027);
or U22271 (N_22271,N_21426,N_21071);
xor U22272 (N_22272,N_21606,N_21625);
nor U22273 (N_22273,N_21184,N_21825);
nor U22274 (N_22274,N_21609,N_21639);
nand U22275 (N_22275,N_21347,N_21202);
nand U22276 (N_22276,N_21682,N_21696);
or U22277 (N_22277,N_21988,N_21422);
xnor U22278 (N_22278,N_21959,N_21899);
nand U22279 (N_22279,N_21764,N_21256);
xor U22280 (N_22280,N_21243,N_21743);
and U22281 (N_22281,N_21671,N_21484);
or U22282 (N_22282,N_21950,N_21790);
and U22283 (N_22283,N_21035,N_21130);
and U22284 (N_22284,N_21093,N_21874);
nand U22285 (N_22285,N_21907,N_21604);
and U22286 (N_22286,N_21665,N_21834);
or U22287 (N_22287,N_21666,N_21513);
and U22288 (N_22288,N_21127,N_21315);
xor U22289 (N_22289,N_21662,N_21090);
nand U22290 (N_22290,N_21012,N_21100);
and U22291 (N_22291,N_21646,N_21466);
nor U22292 (N_22292,N_21376,N_21501);
nor U22293 (N_22293,N_21175,N_21663);
xnor U22294 (N_22294,N_21482,N_21694);
or U22295 (N_22295,N_21782,N_21940);
or U22296 (N_22296,N_21383,N_21414);
or U22297 (N_22297,N_21479,N_21710);
nor U22298 (N_22298,N_21919,N_21525);
nand U22299 (N_22299,N_21246,N_21641);
or U22300 (N_22300,N_21621,N_21096);
xnor U22301 (N_22301,N_21290,N_21925);
or U22302 (N_22302,N_21658,N_21059);
nand U22303 (N_22303,N_21541,N_21158);
nand U22304 (N_22304,N_21066,N_21450);
and U22305 (N_22305,N_21931,N_21164);
and U22306 (N_22306,N_21858,N_21454);
and U22307 (N_22307,N_21885,N_21538);
xnor U22308 (N_22308,N_21280,N_21185);
and U22309 (N_22309,N_21188,N_21711);
nand U22310 (N_22310,N_21546,N_21611);
nand U22311 (N_22311,N_21470,N_21159);
xor U22312 (N_22312,N_21132,N_21674);
nor U22313 (N_22313,N_21379,N_21193);
or U22314 (N_22314,N_21624,N_21613);
nor U22315 (N_22315,N_21234,N_21403);
or U22316 (N_22316,N_21195,N_21751);
nor U22317 (N_22317,N_21011,N_21342);
or U22318 (N_22318,N_21791,N_21288);
xor U22319 (N_22319,N_21259,N_21780);
nor U22320 (N_22320,N_21086,N_21626);
nor U22321 (N_22321,N_21632,N_21612);
or U22322 (N_22322,N_21088,N_21451);
nor U22323 (N_22323,N_21855,N_21445);
nor U22324 (N_22324,N_21372,N_21084);
nor U22325 (N_22325,N_21496,N_21442);
or U22326 (N_22326,N_21872,N_21254);
and U22327 (N_22327,N_21552,N_21745);
or U22328 (N_22328,N_21017,N_21034);
nor U22329 (N_22329,N_21031,N_21652);
or U22330 (N_22330,N_21543,N_21952);
and U22331 (N_22331,N_21381,N_21326);
and U22332 (N_22332,N_21500,N_21723);
and U22333 (N_22333,N_21046,N_21018);
xor U22334 (N_22334,N_21363,N_21707);
or U22335 (N_22335,N_21190,N_21638);
or U22336 (N_22336,N_21786,N_21307);
or U22337 (N_22337,N_21057,N_21218);
or U22338 (N_22338,N_21948,N_21183);
and U22339 (N_22339,N_21317,N_21287);
xor U22340 (N_22340,N_21293,N_21402);
nor U22341 (N_22341,N_21236,N_21168);
xor U22342 (N_22342,N_21987,N_21415);
or U22343 (N_22343,N_21082,N_21079);
or U22344 (N_22344,N_21615,N_21478);
and U22345 (N_22345,N_21553,N_21973);
and U22346 (N_22346,N_21486,N_21762);
nor U22347 (N_22347,N_21635,N_21303);
or U22348 (N_22348,N_21245,N_21519);
xor U22349 (N_22349,N_21873,N_21920);
nor U22350 (N_22350,N_21738,N_21897);
or U22351 (N_22351,N_21019,N_21060);
and U22352 (N_22352,N_21475,N_21802);
nand U22353 (N_22353,N_21367,N_21425);
nor U22354 (N_22354,N_21396,N_21728);
and U22355 (N_22355,N_21945,N_21584);
nor U22356 (N_22356,N_21983,N_21410);
or U22357 (N_22357,N_21359,N_21895);
and U22358 (N_22358,N_21490,N_21917);
nand U22359 (N_22359,N_21687,N_21637);
and U22360 (N_22360,N_21908,N_21197);
xor U22361 (N_22361,N_21441,N_21536);
xnor U22362 (N_22362,N_21139,N_21563);
nand U22363 (N_22363,N_21577,N_21080);
xnor U22364 (N_22364,N_21851,N_21067);
and U22365 (N_22365,N_21155,N_21413);
nor U22366 (N_22366,N_21618,N_21304);
nor U22367 (N_22367,N_21896,N_21619);
nor U22368 (N_22368,N_21160,N_21593);
and U22369 (N_22369,N_21720,N_21529);
xor U22370 (N_22370,N_21404,N_21592);
nor U22371 (N_22371,N_21886,N_21697);
or U22372 (N_22372,N_21203,N_21469);
nor U22373 (N_22373,N_21929,N_21149);
or U22374 (N_22374,N_21337,N_21930);
nand U22375 (N_22375,N_21014,N_21590);
nor U22376 (N_22376,N_21527,N_21412);
xor U22377 (N_22377,N_21398,N_21718);
and U22378 (N_22378,N_21278,N_21216);
nand U22379 (N_22379,N_21033,N_21818);
or U22380 (N_22380,N_21170,N_21141);
nor U22381 (N_22381,N_21434,N_21028);
or U22382 (N_22382,N_21860,N_21557);
nor U22383 (N_22383,N_21788,N_21648);
nor U22384 (N_22384,N_21461,N_21794);
or U22385 (N_22385,N_21248,N_21201);
nor U22386 (N_22386,N_21965,N_21462);
and U22387 (N_22387,N_21455,N_21143);
nor U22388 (N_22388,N_21225,N_21984);
xor U22389 (N_22389,N_21137,N_21889);
and U22390 (N_22390,N_21923,N_21951);
or U22391 (N_22391,N_21166,N_21472);
xnor U22392 (N_22392,N_21114,N_21407);
or U22393 (N_22393,N_21839,N_21651);
xor U22394 (N_22394,N_21110,N_21106);
and U22395 (N_22395,N_21443,N_21186);
xnor U22396 (N_22396,N_21112,N_21961);
nor U22397 (N_22397,N_21157,N_21630);
nor U22398 (N_22398,N_21316,N_21135);
nand U22399 (N_22399,N_21540,N_21438);
or U22400 (N_22400,N_21926,N_21165);
nor U22401 (N_22401,N_21910,N_21111);
or U22402 (N_22402,N_21798,N_21776);
nand U22403 (N_22403,N_21097,N_21121);
or U22404 (N_22404,N_21668,N_21752);
nor U22405 (N_22405,N_21116,N_21747);
and U22406 (N_22406,N_21781,N_21228);
nand U22407 (N_22407,N_21054,N_21437);
nor U22408 (N_22408,N_21497,N_21117);
or U22409 (N_22409,N_21123,N_21255);
xor U22410 (N_22410,N_21432,N_21918);
and U22411 (N_22411,N_21705,N_21555);
or U22412 (N_22412,N_21832,N_21477);
and U22413 (N_22413,N_21594,N_21174);
nand U22414 (N_22414,N_21727,N_21568);
nor U22415 (N_22415,N_21792,N_21570);
or U22416 (N_22416,N_21073,N_21672);
and U22417 (N_22417,N_21876,N_21701);
nor U22418 (N_22418,N_21230,N_21580);
xor U22419 (N_22419,N_21761,N_21456);
xnor U22420 (N_22420,N_21313,N_21401);
nor U22421 (N_22421,N_21340,N_21043);
xnor U22422 (N_22422,N_21585,N_21823);
xor U22423 (N_22423,N_21042,N_21179);
or U22424 (N_22424,N_21870,N_21713);
or U22425 (N_22425,N_21329,N_21518);
nor U22426 (N_22426,N_21471,N_21844);
and U22427 (N_22427,N_21936,N_21564);
or U22428 (N_22428,N_21204,N_21838);
xor U22429 (N_22429,N_21754,N_21583);
or U22430 (N_22430,N_21229,N_21622);
or U22431 (N_22431,N_21815,N_21215);
xnor U22432 (N_22432,N_21756,N_21194);
or U22433 (N_22433,N_21817,N_21180);
nor U22434 (N_22434,N_21252,N_21820);
nor U22435 (N_22435,N_21373,N_21055);
xnor U22436 (N_22436,N_21596,N_21721);
and U22437 (N_22437,N_21560,N_21772);
nor U22438 (N_22438,N_21483,N_21704);
nor U22439 (N_22439,N_21506,N_21015);
xor U22440 (N_22440,N_21579,N_21503);
nand U22441 (N_22441,N_21026,N_21599);
and U22442 (N_22442,N_21325,N_21270);
nand U22443 (N_22443,N_21982,N_21251);
nand U22444 (N_22444,N_21657,N_21405);
xor U22445 (N_22445,N_21567,N_21189);
and U22446 (N_22446,N_21200,N_21775);
nand U22447 (N_22447,N_21083,N_21085);
and U22448 (N_22448,N_21458,N_21348);
or U22449 (N_22449,N_21554,N_21361);
nor U22450 (N_22450,N_21358,N_21654);
xor U22451 (N_22451,N_21810,N_21901);
nand U22452 (N_22452,N_21911,N_21642);
nand U22453 (N_22453,N_21680,N_21309);
xor U22454 (N_22454,N_21693,N_21354);
nand U22455 (N_22455,N_21257,N_21712);
nor U22456 (N_22456,N_21344,N_21806);
or U22457 (N_22457,N_21468,N_21605);
or U22458 (N_22458,N_21285,N_21869);
nand U22459 (N_22459,N_21397,N_21411);
nand U22460 (N_22460,N_21266,N_21273);
nand U22461 (N_22461,N_21587,N_21608);
nor U22462 (N_22462,N_21517,N_21655);
nand U22463 (N_22463,N_21370,N_21331);
or U22464 (N_22464,N_21295,N_21534);
and U22465 (N_22465,N_21853,N_21852);
nand U22466 (N_22466,N_21941,N_21467);
and U22467 (N_22467,N_21661,N_21239);
or U22468 (N_22468,N_21418,N_21231);
xor U22469 (N_22469,N_21384,N_21219);
nor U22470 (N_22470,N_21447,N_21542);
nor U22471 (N_22471,N_21922,N_21706);
and U22472 (N_22472,N_21944,N_21050);
xor U22473 (N_22473,N_21669,N_21134);
nor U22474 (N_22474,N_21569,N_21970);
or U22475 (N_22475,N_21830,N_21875);
nor U22476 (N_22476,N_21393,N_21620);
and U22477 (N_22477,N_21240,N_21440);
xor U22478 (N_22478,N_21487,N_21795);
or U22479 (N_22479,N_21595,N_21282);
nor U22480 (N_22480,N_21502,N_21320);
or U22481 (N_22481,N_21038,N_21267);
nor U22482 (N_22482,N_21075,N_21717);
or U22483 (N_22483,N_21351,N_21008);
and U22484 (N_22484,N_21755,N_21670);
or U22485 (N_22485,N_21474,N_21261);
or U22486 (N_22486,N_21753,N_21977);
or U22487 (N_22487,N_21947,N_21476);
or U22488 (N_22488,N_21235,N_21939);
nor U22489 (N_22489,N_21238,N_21481);
nand U22490 (N_22490,N_21833,N_21297);
or U22491 (N_22491,N_21022,N_21115);
and U22492 (N_22492,N_21264,N_21291);
or U22493 (N_22493,N_21887,N_21138);
xor U22494 (N_22494,N_21377,N_21262);
xor U22495 (N_22495,N_21298,N_21113);
xor U22496 (N_22496,N_21558,N_21667);
and U22497 (N_22497,N_21991,N_21979);
xnor U22498 (N_22498,N_21715,N_21061);
nand U22499 (N_22499,N_21512,N_21281);
nand U22500 (N_22500,N_21934,N_21946);
xnor U22501 (N_22501,N_21986,N_21765);
nor U22502 (N_22502,N_21888,N_21603);
or U22503 (N_22503,N_21893,N_21777);
or U22504 (N_22504,N_21635,N_21079);
and U22505 (N_22505,N_21012,N_21528);
xor U22506 (N_22506,N_21069,N_21915);
xnor U22507 (N_22507,N_21019,N_21958);
xnor U22508 (N_22508,N_21671,N_21287);
xnor U22509 (N_22509,N_21684,N_21500);
nor U22510 (N_22510,N_21912,N_21206);
and U22511 (N_22511,N_21836,N_21487);
xor U22512 (N_22512,N_21975,N_21224);
or U22513 (N_22513,N_21873,N_21001);
or U22514 (N_22514,N_21636,N_21241);
nor U22515 (N_22515,N_21723,N_21275);
nand U22516 (N_22516,N_21910,N_21949);
and U22517 (N_22517,N_21931,N_21809);
and U22518 (N_22518,N_21272,N_21723);
nor U22519 (N_22519,N_21960,N_21066);
nand U22520 (N_22520,N_21361,N_21515);
nand U22521 (N_22521,N_21616,N_21375);
or U22522 (N_22522,N_21339,N_21883);
or U22523 (N_22523,N_21718,N_21481);
nand U22524 (N_22524,N_21294,N_21630);
nor U22525 (N_22525,N_21849,N_21118);
nor U22526 (N_22526,N_21302,N_21917);
nand U22527 (N_22527,N_21270,N_21486);
nor U22528 (N_22528,N_21455,N_21661);
xnor U22529 (N_22529,N_21896,N_21453);
nor U22530 (N_22530,N_21667,N_21825);
nor U22531 (N_22531,N_21055,N_21663);
or U22532 (N_22532,N_21635,N_21512);
xor U22533 (N_22533,N_21795,N_21027);
nand U22534 (N_22534,N_21338,N_21176);
or U22535 (N_22535,N_21051,N_21242);
or U22536 (N_22536,N_21224,N_21472);
or U22537 (N_22537,N_21469,N_21368);
xor U22538 (N_22538,N_21356,N_21739);
or U22539 (N_22539,N_21852,N_21193);
and U22540 (N_22540,N_21314,N_21436);
nor U22541 (N_22541,N_21447,N_21686);
nor U22542 (N_22542,N_21684,N_21755);
nor U22543 (N_22543,N_21298,N_21584);
xnor U22544 (N_22544,N_21345,N_21417);
nor U22545 (N_22545,N_21905,N_21582);
and U22546 (N_22546,N_21897,N_21330);
or U22547 (N_22547,N_21138,N_21617);
and U22548 (N_22548,N_21243,N_21828);
xor U22549 (N_22549,N_21092,N_21742);
and U22550 (N_22550,N_21833,N_21011);
nand U22551 (N_22551,N_21364,N_21260);
nand U22552 (N_22552,N_21780,N_21603);
and U22553 (N_22553,N_21580,N_21242);
and U22554 (N_22554,N_21658,N_21066);
nand U22555 (N_22555,N_21140,N_21402);
nand U22556 (N_22556,N_21703,N_21133);
xor U22557 (N_22557,N_21086,N_21371);
nand U22558 (N_22558,N_21026,N_21310);
or U22559 (N_22559,N_21668,N_21783);
nand U22560 (N_22560,N_21909,N_21282);
nor U22561 (N_22561,N_21829,N_21375);
and U22562 (N_22562,N_21241,N_21102);
and U22563 (N_22563,N_21909,N_21260);
nor U22564 (N_22564,N_21792,N_21264);
and U22565 (N_22565,N_21049,N_21721);
nand U22566 (N_22566,N_21167,N_21844);
or U22567 (N_22567,N_21911,N_21516);
or U22568 (N_22568,N_21565,N_21755);
and U22569 (N_22569,N_21624,N_21916);
and U22570 (N_22570,N_21766,N_21722);
nand U22571 (N_22571,N_21277,N_21466);
or U22572 (N_22572,N_21143,N_21062);
or U22573 (N_22573,N_21309,N_21605);
xor U22574 (N_22574,N_21605,N_21945);
nand U22575 (N_22575,N_21822,N_21719);
xnor U22576 (N_22576,N_21367,N_21922);
nor U22577 (N_22577,N_21950,N_21981);
nand U22578 (N_22578,N_21116,N_21845);
nand U22579 (N_22579,N_21125,N_21586);
xor U22580 (N_22580,N_21836,N_21618);
xor U22581 (N_22581,N_21684,N_21035);
or U22582 (N_22582,N_21066,N_21372);
nor U22583 (N_22583,N_21295,N_21513);
or U22584 (N_22584,N_21625,N_21791);
xor U22585 (N_22585,N_21615,N_21370);
nor U22586 (N_22586,N_21027,N_21369);
and U22587 (N_22587,N_21334,N_21518);
or U22588 (N_22588,N_21756,N_21415);
xor U22589 (N_22589,N_21997,N_21274);
nor U22590 (N_22590,N_21073,N_21219);
or U22591 (N_22591,N_21553,N_21136);
nor U22592 (N_22592,N_21231,N_21581);
or U22593 (N_22593,N_21296,N_21579);
and U22594 (N_22594,N_21442,N_21335);
or U22595 (N_22595,N_21071,N_21900);
nand U22596 (N_22596,N_21427,N_21247);
or U22597 (N_22597,N_21540,N_21469);
nand U22598 (N_22598,N_21307,N_21426);
or U22599 (N_22599,N_21262,N_21364);
and U22600 (N_22600,N_21110,N_21282);
nor U22601 (N_22601,N_21139,N_21025);
nand U22602 (N_22602,N_21475,N_21604);
xnor U22603 (N_22603,N_21252,N_21163);
nor U22604 (N_22604,N_21459,N_21185);
or U22605 (N_22605,N_21917,N_21171);
and U22606 (N_22606,N_21538,N_21347);
nand U22607 (N_22607,N_21335,N_21423);
and U22608 (N_22608,N_21577,N_21891);
nor U22609 (N_22609,N_21144,N_21040);
nand U22610 (N_22610,N_21098,N_21357);
xor U22611 (N_22611,N_21680,N_21706);
xnor U22612 (N_22612,N_21204,N_21140);
nand U22613 (N_22613,N_21273,N_21989);
xor U22614 (N_22614,N_21691,N_21628);
and U22615 (N_22615,N_21951,N_21619);
and U22616 (N_22616,N_21294,N_21932);
xnor U22617 (N_22617,N_21434,N_21240);
nand U22618 (N_22618,N_21558,N_21174);
or U22619 (N_22619,N_21598,N_21106);
nand U22620 (N_22620,N_21082,N_21268);
xor U22621 (N_22621,N_21805,N_21343);
xnor U22622 (N_22622,N_21592,N_21844);
and U22623 (N_22623,N_21991,N_21484);
or U22624 (N_22624,N_21335,N_21781);
xor U22625 (N_22625,N_21211,N_21142);
nand U22626 (N_22626,N_21494,N_21750);
or U22627 (N_22627,N_21228,N_21848);
or U22628 (N_22628,N_21888,N_21464);
nand U22629 (N_22629,N_21419,N_21203);
nand U22630 (N_22630,N_21036,N_21103);
xor U22631 (N_22631,N_21051,N_21286);
and U22632 (N_22632,N_21653,N_21911);
nor U22633 (N_22633,N_21258,N_21798);
xnor U22634 (N_22634,N_21927,N_21012);
xnor U22635 (N_22635,N_21192,N_21812);
or U22636 (N_22636,N_21984,N_21506);
nand U22637 (N_22637,N_21154,N_21293);
nor U22638 (N_22638,N_21561,N_21390);
nand U22639 (N_22639,N_21425,N_21056);
nand U22640 (N_22640,N_21226,N_21965);
and U22641 (N_22641,N_21365,N_21456);
and U22642 (N_22642,N_21670,N_21442);
xnor U22643 (N_22643,N_21111,N_21430);
nand U22644 (N_22644,N_21826,N_21049);
nor U22645 (N_22645,N_21385,N_21103);
xor U22646 (N_22646,N_21920,N_21200);
nand U22647 (N_22647,N_21755,N_21115);
and U22648 (N_22648,N_21184,N_21020);
and U22649 (N_22649,N_21359,N_21116);
xor U22650 (N_22650,N_21951,N_21114);
or U22651 (N_22651,N_21701,N_21392);
xor U22652 (N_22652,N_21959,N_21206);
nand U22653 (N_22653,N_21179,N_21599);
nand U22654 (N_22654,N_21008,N_21722);
and U22655 (N_22655,N_21893,N_21153);
xor U22656 (N_22656,N_21326,N_21222);
nor U22657 (N_22657,N_21723,N_21594);
nor U22658 (N_22658,N_21194,N_21257);
xor U22659 (N_22659,N_21412,N_21296);
xor U22660 (N_22660,N_21272,N_21487);
nand U22661 (N_22661,N_21338,N_21554);
and U22662 (N_22662,N_21286,N_21296);
xor U22663 (N_22663,N_21682,N_21839);
xnor U22664 (N_22664,N_21329,N_21986);
xnor U22665 (N_22665,N_21217,N_21670);
and U22666 (N_22666,N_21744,N_21233);
nand U22667 (N_22667,N_21003,N_21773);
or U22668 (N_22668,N_21875,N_21337);
nand U22669 (N_22669,N_21701,N_21017);
nand U22670 (N_22670,N_21340,N_21624);
or U22671 (N_22671,N_21052,N_21308);
nor U22672 (N_22672,N_21641,N_21552);
nand U22673 (N_22673,N_21713,N_21402);
xor U22674 (N_22674,N_21637,N_21077);
nand U22675 (N_22675,N_21613,N_21712);
xnor U22676 (N_22676,N_21041,N_21191);
and U22677 (N_22677,N_21084,N_21036);
and U22678 (N_22678,N_21489,N_21916);
xnor U22679 (N_22679,N_21022,N_21661);
nand U22680 (N_22680,N_21236,N_21272);
nor U22681 (N_22681,N_21346,N_21351);
or U22682 (N_22682,N_21188,N_21741);
and U22683 (N_22683,N_21713,N_21832);
xor U22684 (N_22684,N_21420,N_21414);
nor U22685 (N_22685,N_21538,N_21255);
xnor U22686 (N_22686,N_21506,N_21113);
nor U22687 (N_22687,N_21676,N_21822);
xnor U22688 (N_22688,N_21168,N_21993);
or U22689 (N_22689,N_21722,N_21829);
and U22690 (N_22690,N_21684,N_21485);
and U22691 (N_22691,N_21259,N_21866);
xnor U22692 (N_22692,N_21350,N_21113);
nand U22693 (N_22693,N_21669,N_21154);
and U22694 (N_22694,N_21002,N_21924);
nor U22695 (N_22695,N_21693,N_21394);
nand U22696 (N_22696,N_21150,N_21344);
nand U22697 (N_22697,N_21391,N_21434);
and U22698 (N_22698,N_21134,N_21402);
xnor U22699 (N_22699,N_21514,N_21412);
xnor U22700 (N_22700,N_21492,N_21452);
nor U22701 (N_22701,N_21547,N_21404);
nor U22702 (N_22702,N_21370,N_21374);
nand U22703 (N_22703,N_21879,N_21322);
or U22704 (N_22704,N_21677,N_21786);
nor U22705 (N_22705,N_21270,N_21833);
xor U22706 (N_22706,N_21246,N_21939);
and U22707 (N_22707,N_21480,N_21473);
nand U22708 (N_22708,N_21388,N_21016);
nor U22709 (N_22709,N_21327,N_21162);
and U22710 (N_22710,N_21754,N_21076);
or U22711 (N_22711,N_21653,N_21225);
nor U22712 (N_22712,N_21189,N_21109);
xor U22713 (N_22713,N_21510,N_21559);
nand U22714 (N_22714,N_21143,N_21186);
xor U22715 (N_22715,N_21692,N_21971);
or U22716 (N_22716,N_21491,N_21699);
nor U22717 (N_22717,N_21761,N_21859);
or U22718 (N_22718,N_21639,N_21604);
nand U22719 (N_22719,N_21655,N_21037);
nor U22720 (N_22720,N_21562,N_21209);
nand U22721 (N_22721,N_21044,N_21510);
xnor U22722 (N_22722,N_21245,N_21544);
and U22723 (N_22723,N_21977,N_21075);
nand U22724 (N_22724,N_21988,N_21190);
nor U22725 (N_22725,N_21669,N_21624);
nand U22726 (N_22726,N_21502,N_21416);
or U22727 (N_22727,N_21271,N_21134);
xor U22728 (N_22728,N_21478,N_21518);
xor U22729 (N_22729,N_21882,N_21233);
and U22730 (N_22730,N_21614,N_21528);
nand U22731 (N_22731,N_21250,N_21085);
or U22732 (N_22732,N_21895,N_21524);
nand U22733 (N_22733,N_21433,N_21055);
xor U22734 (N_22734,N_21723,N_21822);
nand U22735 (N_22735,N_21696,N_21514);
nor U22736 (N_22736,N_21841,N_21747);
or U22737 (N_22737,N_21785,N_21366);
xnor U22738 (N_22738,N_21256,N_21845);
nand U22739 (N_22739,N_21583,N_21080);
xnor U22740 (N_22740,N_21150,N_21650);
or U22741 (N_22741,N_21048,N_21928);
nand U22742 (N_22742,N_21580,N_21328);
and U22743 (N_22743,N_21891,N_21994);
or U22744 (N_22744,N_21935,N_21106);
or U22745 (N_22745,N_21329,N_21809);
nor U22746 (N_22746,N_21213,N_21404);
or U22747 (N_22747,N_21796,N_21243);
or U22748 (N_22748,N_21953,N_21344);
nand U22749 (N_22749,N_21534,N_21868);
xor U22750 (N_22750,N_21394,N_21038);
nor U22751 (N_22751,N_21324,N_21534);
nand U22752 (N_22752,N_21862,N_21111);
or U22753 (N_22753,N_21607,N_21856);
xnor U22754 (N_22754,N_21906,N_21776);
xnor U22755 (N_22755,N_21753,N_21897);
nor U22756 (N_22756,N_21492,N_21607);
xor U22757 (N_22757,N_21347,N_21275);
and U22758 (N_22758,N_21060,N_21959);
nand U22759 (N_22759,N_21733,N_21791);
nand U22760 (N_22760,N_21630,N_21016);
and U22761 (N_22761,N_21781,N_21492);
and U22762 (N_22762,N_21946,N_21711);
and U22763 (N_22763,N_21917,N_21721);
nor U22764 (N_22764,N_21312,N_21573);
or U22765 (N_22765,N_21001,N_21428);
nor U22766 (N_22766,N_21482,N_21998);
or U22767 (N_22767,N_21369,N_21711);
or U22768 (N_22768,N_21054,N_21523);
nor U22769 (N_22769,N_21147,N_21902);
nand U22770 (N_22770,N_21592,N_21031);
nor U22771 (N_22771,N_21577,N_21145);
nor U22772 (N_22772,N_21755,N_21434);
or U22773 (N_22773,N_21285,N_21697);
or U22774 (N_22774,N_21241,N_21284);
and U22775 (N_22775,N_21781,N_21005);
xnor U22776 (N_22776,N_21252,N_21492);
nor U22777 (N_22777,N_21128,N_21157);
or U22778 (N_22778,N_21901,N_21518);
nor U22779 (N_22779,N_21121,N_21347);
xor U22780 (N_22780,N_21465,N_21047);
or U22781 (N_22781,N_21258,N_21428);
nor U22782 (N_22782,N_21276,N_21253);
xor U22783 (N_22783,N_21660,N_21288);
nand U22784 (N_22784,N_21204,N_21331);
xnor U22785 (N_22785,N_21657,N_21425);
or U22786 (N_22786,N_21737,N_21038);
nand U22787 (N_22787,N_21392,N_21240);
and U22788 (N_22788,N_21604,N_21436);
nor U22789 (N_22789,N_21669,N_21114);
or U22790 (N_22790,N_21136,N_21151);
xnor U22791 (N_22791,N_21231,N_21224);
and U22792 (N_22792,N_21359,N_21486);
nand U22793 (N_22793,N_21948,N_21736);
nor U22794 (N_22794,N_21897,N_21197);
nand U22795 (N_22795,N_21329,N_21063);
or U22796 (N_22796,N_21864,N_21908);
nor U22797 (N_22797,N_21789,N_21899);
nand U22798 (N_22798,N_21559,N_21018);
xor U22799 (N_22799,N_21478,N_21792);
nor U22800 (N_22800,N_21868,N_21623);
nor U22801 (N_22801,N_21754,N_21825);
xnor U22802 (N_22802,N_21080,N_21861);
or U22803 (N_22803,N_21190,N_21497);
nand U22804 (N_22804,N_21407,N_21640);
xor U22805 (N_22805,N_21034,N_21300);
xnor U22806 (N_22806,N_21468,N_21260);
nand U22807 (N_22807,N_21392,N_21649);
or U22808 (N_22808,N_21617,N_21657);
nand U22809 (N_22809,N_21982,N_21546);
xor U22810 (N_22810,N_21441,N_21810);
nor U22811 (N_22811,N_21214,N_21530);
nor U22812 (N_22812,N_21432,N_21032);
xor U22813 (N_22813,N_21201,N_21506);
xor U22814 (N_22814,N_21813,N_21301);
and U22815 (N_22815,N_21835,N_21926);
nand U22816 (N_22816,N_21052,N_21191);
xor U22817 (N_22817,N_21124,N_21667);
or U22818 (N_22818,N_21964,N_21759);
nand U22819 (N_22819,N_21137,N_21818);
or U22820 (N_22820,N_21495,N_21111);
or U22821 (N_22821,N_21545,N_21782);
xnor U22822 (N_22822,N_21985,N_21379);
or U22823 (N_22823,N_21740,N_21691);
or U22824 (N_22824,N_21671,N_21463);
or U22825 (N_22825,N_21851,N_21010);
nor U22826 (N_22826,N_21949,N_21384);
and U22827 (N_22827,N_21081,N_21440);
nor U22828 (N_22828,N_21945,N_21194);
and U22829 (N_22829,N_21771,N_21468);
nand U22830 (N_22830,N_21927,N_21021);
and U22831 (N_22831,N_21643,N_21017);
nand U22832 (N_22832,N_21601,N_21245);
and U22833 (N_22833,N_21195,N_21614);
xor U22834 (N_22834,N_21519,N_21686);
or U22835 (N_22835,N_21375,N_21069);
or U22836 (N_22836,N_21077,N_21437);
xor U22837 (N_22837,N_21596,N_21191);
xor U22838 (N_22838,N_21113,N_21725);
nand U22839 (N_22839,N_21488,N_21209);
xnor U22840 (N_22840,N_21497,N_21559);
nor U22841 (N_22841,N_21183,N_21010);
nor U22842 (N_22842,N_21527,N_21232);
and U22843 (N_22843,N_21542,N_21730);
nand U22844 (N_22844,N_21777,N_21694);
xor U22845 (N_22845,N_21208,N_21062);
xnor U22846 (N_22846,N_21749,N_21156);
xor U22847 (N_22847,N_21237,N_21472);
xor U22848 (N_22848,N_21192,N_21799);
nand U22849 (N_22849,N_21300,N_21735);
nor U22850 (N_22850,N_21607,N_21752);
nand U22851 (N_22851,N_21582,N_21813);
nand U22852 (N_22852,N_21387,N_21818);
and U22853 (N_22853,N_21706,N_21119);
nor U22854 (N_22854,N_21257,N_21719);
or U22855 (N_22855,N_21711,N_21900);
nand U22856 (N_22856,N_21118,N_21601);
xnor U22857 (N_22857,N_21554,N_21090);
and U22858 (N_22858,N_21680,N_21848);
xnor U22859 (N_22859,N_21375,N_21010);
and U22860 (N_22860,N_21026,N_21142);
and U22861 (N_22861,N_21231,N_21096);
nand U22862 (N_22862,N_21581,N_21928);
nand U22863 (N_22863,N_21819,N_21932);
and U22864 (N_22864,N_21451,N_21521);
or U22865 (N_22865,N_21820,N_21935);
nand U22866 (N_22866,N_21292,N_21903);
and U22867 (N_22867,N_21613,N_21930);
nand U22868 (N_22868,N_21215,N_21280);
or U22869 (N_22869,N_21513,N_21053);
nand U22870 (N_22870,N_21309,N_21916);
or U22871 (N_22871,N_21787,N_21669);
xor U22872 (N_22872,N_21471,N_21970);
and U22873 (N_22873,N_21393,N_21403);
xor U22874 (N_22874,N_21127,N_21602);
nor U22875 (N_22875,N_21561,N_21387);
xnor U22876 (N_22876,N_21894,N_21788);
nand U22877 (N_22877,N_21148,N_21294);
and U22878 (N_22878,N_21004,N_21068);
and U22879 (N_22879,N_21450,N_21872);
and U22880 (N_22880,N_21658,N_21389);
nand U22881 (N_22881,N_21743,N_21282);
or U22882 (N_22882,N_21259,N_21757);
and U22883 (N_22883,N_21319,N_21982);
nand U22884 (N_22884,N_21514,N_21614);
or U22885 (N_22885,N_21907,N_21352);
and U22886 (N_22886,N_21477,N_21566);
or U22887 (N_22887,N_21032,N_21641);
or U22888 (N_22888,N_21857,N_21000);
and U22889 (N_22889,N_21307,N_21977);
nand U22890 (N_22890,N_21494,N_21017);
or U22891 (N_22891,N_21219,N_21388);
or U22892 (N_22892,N_21516,N_21985);
nand U22893 (N_22893,N_21376,N_21118);
nand U22894 (N_22894,N_21089,N_21903);
xnor U22895 (N_22895,N_21380,N_21187);
xnor U22896 (N_22896,N_21496,N_21265);
nand U22897 (N_22897,N_21926,N_21047);
or U22898 (N_22898,N_21030,N_21354);
xor U22899 (N_22899,N_21633,N_21465);
nand U22900 (N_22900,N_21758,N_21045);
nand U22901 (N_22901,N_21056,N_21474);
and U22902 (N_22902,N_21928,N_21939);
nand U22903 (N_22903,N_21115,N_21275);
nor U22904 (N_22904,N_21974,N_21787);
nor U22905 (N_22905,N_21187,N_21619);
and U22906 (N_22906,N_21392,N_21740);
or U22907 (N_22907,N_21162,N_21936);
and U22908 (N_22908,N_21884,N_21465);
nor U22909 (N_22909,N_21514,N_21488);
nor U22910 (N_22910,N_21908,N_21265);
and U22911 (N_22911,N_21877,N_21249);
nand U22912 (N_22912,N_21184,N_21892);
xor U22913 (N_22913,N_21700,N_21788);
nor U22914 (N_22914,N_21398,N_21004);
nand U22915 (N_22915,N_21829,N_21607);
nor U22916 (N_22916,N_21141,N_21916);
or U22917 (N_22917,N_21970,N_21812);
nor U22918 (N_22918,N_21757,N_21604);
xor U22919 (N_22919,N_21882,N_21553);
or U22920 (N_22920,N_21848,N_21904);
nor U22921 (N_22921,N_21449,N_21336);
nor U22922 (N_22922,N_21388,N_21921);
and U22923 (N_22923,N_21522,N_21706);
or U22924 (N_22924,N_21712,N_21569);
nand U22925 (N_22925,N_21682,N_21415);
nor U22926 (N_22926,N_21915,N_21602);
nand U22927 (N_22927,N_21260,N_21246);
nand U22928 (N_22928,N_21018,N_21141);
nor U22929 (N_22929,N_21903,N_21443);
and U22930 (N_22930,N_21735,N_21390);
or U22931 (N_22931,N_21586,N_21899);
and U22932 (N_22932,N_21248,N_21087);
and U22933 (N_22933,N_21634,N_21577);
nand U22934 (N_22934,N_21378,N_21314);
or U22935 (N_22935,N_21223,N_21124);
and U22936 (N_22936,N_21037,N_21441);
xnor U22937 (N_22937,N_21761,N_21007);
or U22938 (N_22938,N_21673,N_21310);
or U22939 (N_22939,N_21701,N_21364);
xnor U22940 (N_22940,N_21608,N_21130);
and U22941 (N_22941,N_21048,N_21654);
or U22942 (N_22942,N_21214,N_21235);
nand U22943 (N_22943,N_21725,N_21633);
nor U22944 (N_22944,N_21458,N_21616);
or U22945 (N_22945,N_21159,N_21075);
xor U22946 (N_22946,N_21425,N_21044);
or U22947 (N_22947,N_21013,N_21579);
nand U22948 (N_22948,N_21012,N_21377);
xor U22949 (N_22949,N_21717,N_21942);
nand U22950 (N_22950,N_21361,N_21478);
xnor U22951 (N_22951,N_21840,N_21244);
xor U22952 (N_22952,N_21755,N_21224);
and U22953 (N_22953,N_21306,N_21595);
nor U22954 (N_22954,N_21568,N_21182);
or U22955 (N_22955,N_21376,N_21387);
nand U22956 (N_22956,N_21028,N_21528);
nand U22957 (N_22957,N_21739,N_21414);
nand U22958 (N_22958,N_21797,N_21219);
nand U22959 (N_22959,N_21814,N_21793);
nor U22960 (N_22960,N_21587,N_21784);
xor U22961 (N_22961,N_21037,N_21499);
nor U22962 (N_22962,N_21049,N_21591);
or U22963 (N_22963,N_21168,N_21759);
nand U22964 (N_22964,N_21288,N_21365);
xor U22965 (N_22965,N_21666,N_21558);
or U22966 (N_22966,N_21535,N_21248);
and U22967 (N_22967,N_21219,N_21719);
nand U22968 (N_22968,N_21775,N_21927);
or U22969 (N_22969,N_21734,N_21716);
nand U22970 (N_22970,N_21225,N_21502);
or U22971 (N_22971,N_21821,N_21624);
xnor U22972 (N_22972,N_21133,N_21619);
nor U22973 (N_22973,N_21617,N_21289);
or U22974 (N_22974,N_21399,N_21357);
nor U22975 (N_22975,N_21899,N_21003);
and U22976 (N_22976,N_21678,N_21779);
or U22977 (N_22977,N_21485,N_21177);
xnor U22978 (N_22978,N_21391,N_21846);
nor U22979 (N_22979,N_21499,N_21141);
nand U22980 (N_22980,N_21060,N_21530);
nand U22981 (N_22981,N_21286,N_21381);
xnor U22982 (N_22982,N_21183,N_21968);
nand U22983 (N_22983,N_21780,N_21003);
and U22984 (N_22984,N_21000,N_21096);
xor U22985 (N_22985,N_21304,N_21276);
or U22986 (N_22986,N_21046,N_21808);
and U22987 (N_22987,N_21476,N_21602);
nor U22988 (N_22988,N_21059,N_21569);
nor U22989 (N_22989,N_21277,N_21454);
nor U22990 (N_22990,N_21525,N_21459);
xnor U22991 (N_22991,N_21243,N_21184);
or U22992 (N_22992,N_21636,N_21465);
and U22993 (N_22993,N_21633,N_21002);
nor U22994 (N_22994,N_21779,N_21760);
and U22995 (N_22995,N_21011,N_21466);
nor U22996 (N_22996,N_21893,N_21852);
and U22997 (N_22997,N_21902,N_21984);
or U22998 (N_22998,N_21068,N_21044);
nor U22999 (N_22999,N_21711,N_21593);
nor U23000 (N_23000,N_22695,N_22135);
nor U23001 (N_23001,N_22208,N_22255);
and U23002 (N_23002,N_22162,N_22715);
xnor U23003 (N_23003,N_22552,N_22098);
xnor U23004 (N_23004,N_22846,N_22259);
nor U23005 (N_23005,N_22563,N_22944);
and U23006 (N_23006,N_22906,N_22340);
nand U23007 (N_23007,N_22431,N_22395);
and U23008 (N_23008,N_22169,N_22678);
or U23009 (N_23009,N_22618,N_22869);
and U23010 (N_23010,N_22933,N_22280);
or U23011 (N_23011,N_22472,N_22610);
nor U23012 (N_23012,N_22133,N_22331);
and U23013 (N_23013,N_22424,N_22612);
or U23014 (N_23014,N_22912,N_22544);
or U23015 (N_23015,N_22288,N_22414);
nor U23016 (N_23016,N_22389,N_22591);
or U23017 (N_23017,N_22894,N_22951);
nor U23018 (N_23018,N_22700,N_22038);
xnor U23019 (N_23019,N_22959,N_22304);
and U23020 (N_23020,N_22290,N_22952);
nor U23021 (N_23021,N_22228,N_22823);
nor U23022 (N_23022,N_22198,N_22307);
nand U23023 (N_23023,N_22181,N_22673);
nand U23024 (N_23024,N_22390,N_22454);
and U23025 (N_23025,N_22024,N_22187);
and U23026 (N_23026,N_22252,N_22438);
nor U23027 (N_23027,N_22836,N_22412);
xor U23028 (N_23028,N_22811,N_22603);
xnor U23029 (N_23029,N_22097,N_22997);
or U23030 (N_23030,N_22049,N_22352);
and U23031 (N_23031,N_22175,N_22273);
or U23032 (N_23032,N_22157,N_22735);
nand U23033 (N_23033,N_22163,N_22191);
nor U23034 (N_23034,N_22817,N_22281);
and U23035 (N_23035,N_22372,N_22654);
or U23036 (N_23036,N_22860,N_22423);
nor U23037 (N_23037,N_22556,N_22201);
or U23038 (N_23038,N_22889,N_22911);
and U23039 (N_23039,N_22752,N_22853);
xnor U23040 (N_23040,N_22196,N_22266);
or U23041 (N_23041,N_22670,N_22029);
and U23042 (N_23042,N_22623,N_22689);
nor U23043 (N_23043,N_22643,N_22709);
or U23044 (N_23044,N_22599,N_22347);
nand U23045 (N_23045,N_22743,N_22158);
nand U23046 (N_23046,N_22718,N_22303);
xor U23047 (N_23047,N_22770,N_22286);
and U23048 (N_23048,N_22248,N_22453);
xnor U23049 (N_23049,N_22131,N_22102);
or U23050 (N_23050,N_22408,N_22047);
and U23051 (N_23051,N_22436,N_22510);
nand U23052 (N_23052,N_22236,N_22642);
and U23053 (N_23053,N_22921,N_22663);
xnor U23054 (N_23054,N_22729,N_22440);
or U23055 (N_23055,N_22891,N_22828);
or U23056 (N_23056,N_22607,N_22213);
or U23057 (N_23057,N_22584,N_22398);
nor U23058 (N_23058,N_22361,N_22675);
xor U23059 (N_23059,N_22815,N_22399);
nor U23060 (N_23060,N_22795,N_22018);
nor U23061 (N_23061,N_22940,N_22659);
xor U23062 (N_23062,N_22503,N_22983);
or U23063 (N_23063,N_22793,N_22798);
xnor U23064 (N_23064,N_22920,N_22238);
xnor U23065 (N_23065,N_22899,N_22230);
or U23066 (N_23066,N_22696,N_22277);
nor U23067 (N_23067,N_22148,N_22996);
xor U23068 (N_23068,N_22123,N_22426);
nand U23069 (N_23069,N_22545,N_22995);
and U23070 (N_23070,N_22596,N_22980);
or U23071 (N_23071,N_22884,N_22564);
or U23072 (N_23072,N_22876,N_22801);
nor U23073 (N_23073,N_22594,N_22573);
xor U23074 (N_23074,N_22922,N_22393);
and U23075 (N_23075,N_22989,N_22542);
nand U23076 (N_23076,N_22125,N_22759);
and U23077 (N_23077,N_22404,N_22726);
xor U23078 (N_23078,N_22085,N_22275);
nor U23079 (N_23079,N_22572,N_22524);
nand U23080 (N_23080,N_22760,N_22189);
or U23081 (N_23081,N_22958,N_22676);
nand U23082 (N_23082,N_22088,N_22879);
nor U23083 (N_23083,N_22566,N_22261);
or U23084 (N_23084,N_22720,N_22224);
nand U23085 (N_23085,N_22342,N_22174);
and U23086 (N_23086,N_22245,N_22704);
xor U23087 (N_23087,N_22755,N_22387);
or U23088 (N_23088,N_22656,N_22433);
xnor U23089 (N_23089,N_22851,N_22750);
and U23090 (N_23090,N_22568,N_22027);
xor U23091 (N_23091,N_22848,N_22621);
nor U23092 (N_23092,N_22341,N_22407);
and U23093 (N_23093,N_22325,N_22740);
xnor U23094 (N_23094,N_22481,N_22880);
nand U23095 (N_23095,N_22871,N_22712);
nand U23096 (N_23096,N_22890,N_22113);
nand U23097 (N_23097,N_22216,N_22114);
xor U23098 (N_23098,N_22075,N_22515);
and U23099 (N_23099,N_22167,N_22053);
xor U23100 (N_23100,N_22519,N_22804);
nand U23101 (N_23101,N_22953,N_22666);
or U23102 (N_23102,N_22600,N_22222);
and U23103 (N_23103,N_22355,N_22956);
nor U23104 (N_23104,N_22776,N_22816);
and U23105 (N_23105,N_22362,N_22727);
nand U23106 (N_23106,N_22437,N_22379);
or U23107 (N_23107,N_22762,N_22608);
nor U23108 (N_23108,N_22525,N_22268);
or U23109 (N_23109,N_22963,N_22471);
xor U23110 (N_23110,N_22716,N_22223);
nor U23111 (N_23111,N_22265,N_22246);
xnor U23112 (N_23112,N_22378,N_22107);
and U23113 (N_23113,N_22301,N_22410);
nor U23114 (N_23114,N_22929,N_22353);
nand U23115 (N_23115,N_22509,N_22072);
xnor U23116 (N_23116,N_22139,N_22893);
xor U23117 (N_23117,N_22930,N_22732);
xnor U23118 (N_23118,N_22419,N_22651);
nor U23119 (N_23119,N_22905,N_22791);
and U23120 (N_23120,N_22885,N_22578);
or U23121 (N_23121,N_22861,N_22206);
or U23122 (N_23122,N_22367,N_22212);
nand U23123 (N_23123,N_22442,N_22311);
and U23124 (N_23124,N_22234,N_22310);
nor U23125 (N_23125,N_22090,N_22766);
or U23126 (N_23126,N_22405,N_22664);
nand U23127 (N_23127,N_22910,N_22486);
nand U23128 (N_23128,N_22647,N_22232);
or U23129 (N_23129,N_22999,N_22067);
nor U23130 (N_23130,N_22706,N_22909);
or U23131 (N_23131,N_22333,N_22420);
nor U23132 (N_23132,N_22253,N_22830);
nand U23133 (N_23133,N_22579,N_22744);
xnor U23134 (N_23134,N_22011,N_22150);
or U23135 (N_23135,N_22692,N_22723);
nor U23136 (N_23136,N_22904,N_22479);
nor U23137 (N_23137,N_22315,N_22957);
nor U23138 (N_23138,N_22687,N_22660);
xor U23139 (N_23139,N_22104,N_22862);
and U23140 (N_23140,N_22639,N_22932);
or U23141 (N_23141,N_22827,N_22403);
and U23142 (N_23142,N_22192,N_22734);
and U23143 (N_23143,N_22597,N_22655);
or U23144 (N_23144,N_22915,N_22209);
or U23145 (N_23145,N_22271,N_22448);
nor U23146 (N_23146,N_22042,N_22942);
and U23147 (N_23147,N_22276,N_22863);
nand U23148 (N_23148,N_22330,N_22926);
and U23149 (N_23149,N_22938,N_22961);
or U23150 (N_23150,N_22172,N_22028);
or U23151 (N_23151,N_22121,N_22226);
nand U23152 (N_23152,N_22781,N_22745);
nor U23153 (N_23153,N_22470,N_22316);
nand U23154 (N_23154,N_22590,N_22918);
nand U23155 (N_23155,N_22358,N_22540);
and U23156 (N_23156,N_22825,N_22243);
and U23157 (N_23157,N_22892,N_22110);
or U23158 (N_23158,N_22914,N_22849);
nand U23159 (N_23159,N_22300,N_22244);
nor U23160 (N_23160,N_22523,N_22026);
nand U23161 (N_23161,N_22981,N_22327);
or U23162 (N_23162,N_22866,N_22284);
and U23163 (N_23163,N_22546,N_22834);
nor U23164 (N_23164,N_22400,N_22570);
nor U23165 (N_23165,N_22332,N_22161);
nand U23166 (N_23166,N_22577,N_22364);
and U23167 (N_23167,N_22051,N_22185);
or U23168 (N_23168,N_22459,N_22394);
nand U23169 (N_23169,N_22576,N_22155);
nand U23170 (N_23170,N_22071,N_22728);
or U23171 (N_23171,N_22747,N_22941);
nor U23172 (N_23172,N_22875,N_22007);
nor U23173 (N_23173,N_22679,N_22547);
nand U23174 (N_23174,N_22535,N_22699);
nor U23175 (N_23175,N_22883,N_22581);
nor U23176 (N_23176,N_22129,N_22124);
xor U23177 (N_23177,N_22320,N_22754);
xnor U23178 (N_23178,N_22377,N_22146);
nand U23179 (N_23179,N_22409,N_22344);
and U23180 (N_23180,N_22324,N_22778);
or U23181 (N_23181,N_22837,N_22193);
nand U23182 (N_23182,N_22595,N_22683);
nor U23183 (N_23183,N_22800,N_22978);
and U23184 (N_23184,N_22009,N_22421);
or U23185 (N_23185,N_22313,N_22166);
and U23186 (N_23186,N_22622,N_22505);
nor U23187 (N_23187,N_22388,N_22231);
nor U23188 (N_23188,N_22374,N_22701);
nor U23189 (N_23189,N_22203,N_22887);
or U23190 (N_23190,N_22021,N_22713);
and U23191 (N_23191,N_22466,N_22588);
xnor U23192 (N_23192,N_22336,N_22428);
nor U23193 (N_23193,N_22658,N_22988);
nand U23194 (N_23194,N_22457,N_22677);
or U23195 (N_23195,N_22548,N_22013);
or U23196 (N_23196,N_22636,N_22613);
or U23197 (N_23197,N_22907,N_22160);
xnor U23198 (N_23198,N_22298,N_22491);
nor U23199 (N_23199,N_22178,N_22725);
and U23200 (N_23200,N_22966,N_22583);
or U23201 (N_23201,N_22946,N_22063);
and U23202 (N_23202,N_22396,N_22217);
xor U23203 (N_23203,N_22173,N_22775);
and U23204 (N_23204,N_22625,N_22418);
xnor U23205 (N_23205,N_22434,N_22010);
nand U23206 (N_23206,N_22200,N_22627);
nor U23207 (N_23207,N_22258,N_22617);
nand U23208 (N_23208,N_22631,N_22368);
nor U23209 (N_23209,N_22257,N_22429);
nand U23210 (N_23210,N_22094,N_22263);
and U23211 (N_23211,N_22741,N_22194);
nand U23212 (N_23212,N_22845,N_22137);
or U23213 (N_23213,N_22052,N_22035);
xor U23214 (N_23214,N_22370,N_22142);
and U23215 (N_23215,N_22649,N_22074);
nand U23216 (N_23216,N_22215,N_22635);
xnor U23217 (N_23217,N_22787,N_22669);
nor U23218 (N_23218,N_22006,N_22425);
xor U23219 (N_23219,N_22780,N_22287);
nand U23220 (N_23220,N_22923,N_22349);
or U23221 (N_23221,N_22291,N_22012);
nor U23222 (N_23222,N_22960,N_22177);
nor U23223 (N_23223,N_22569,N_22348);
and U23224 (N_23224,N_22343,N_22821);
or U23225 (N_23225,N_22242,N_22841);
nor U23226 (N_23226,N_22492,N_22984);
nor U23227 (N_23227,N_22864,N_22705);
or U23228 (N_23228,N_22154,N_22506);
and U23229 (N_23229,N_22199,N_22587);
xor U23230 (N_23230,N_22903,N_22842);
nand U23231 (N_23231,N_22159,N_22707);
nor U23232 (N_23232,N_22784,N_22384);
and U23233 (N_23233,N_22068,N_22919);
or U23234 (N_23234,N_22814,N_22970);
xnor U23235 (N_23235,N_22087,N_22282);
and U23236 (N_23236,N_22939,N_22122);
nor U23237 (N_23237,N_22888,N_22771);
or U23238 (N_23238,N_22992,N_22176);
or U23239 (N_23239,N_22977,N_22065);
or U23240 (N_23240,N_22500,N_22308);
nand U23241 (N_23241,N_22764,N_22809);
nand U23242 (N_23242,N_22401,N_22708);
and U23243 (N_23243,N_22589,N_22501);
nor U23244 (N_23244,N_22822,N_22812);
xor U23245 (N_23245,N_22549,N_22886);
nand U23246 (N_23246,N_22334,N_22422);
nand U23247 (N_23247,N_22877,N_22688);
nand U23248 (N_23248,N_22338,N_22329);
nor U23249 (N_23249,N_22168,N_22974);
nand U23250 (N_23250,N_22789,N_22373);
nor U23251 (N_23251,N_22902,N_22668);
or U23252 (N_23252,N_22702,N_22947);
or U23253 (N_23253,N_22991,N_22628);
nand U23254 (N_23254,N_22824,N_22739);
or U23255 (N_23255,N_22672,N_22554);
nand U23256 (N_23256,N_22116,N_22296);
nor U23257 (N_23257,N_22844,N_22934);
xor U23258 (N_23258,N_22698,N_22153);
nor U23259 (N_23259,N_22742,N_22083);
and U23260 (N_23260,N_22015,N_22602);
nand U23261 (N_23261,N_22084,N_22852);
xnor U23262 (N_23262,N_22030,N_22593);
nand U23263 (N_23263,N_22514,N_22768);
xnor U23264 (N_23264,N_22604,N_22819);
nor U23265 (N_23265,N_22064,N_22897);
xnor U23266 (N_23266,N_22003,N_22773);
nor U23267 (N_23267,N_22369,N_22553);
nor U23268 (N_23268,N_22218,N_22359);
and U23269 (N_23269,N_22360,N_22896);
nor U23270 (N_23270,N_22838,N_22629);
and U23271 (N_23271,N_22054,N_22000);
xnor U23272 (N_23272,N_22684,N_22949);
nand U23273 (N_23273,N_22565,N_22445);
and U23274 (N_23274,N_22820,N_22070);
xor U23275 (N_23275,N_22490,N_22207);
or U23276 (N_23276,N_22620,N_22641);
and U23277 (N_23277,N_22449,N_22513);
xnor U23278 (N_23278,N_22335,N_22210);
nand U23279 (N_23279,N_22127,N_22312);
nand U23280 (N_23280,N_22522,N_22592);
and U23281 (N_23281,N_22898,N_22662);
nor U23282 (N_23282,N_22046,N_22017);
and U23283 (N_23283,N_22551,N_22417);
nand U23284 (N_23284,N_22019,N_22681);
and U23285 (N_23285,N_22475,N_22487);
xnor U23286 (N_23286,N_22204,N_22667);
nand U23287 (N_23287,N_22719,N_22488);
and U23288 (N_23288,N_22632,N_22240);
or U23289 (N_23289,N_22460,N_22044);
xnor U23290 (N_23290,N_22045,N_22859);
and U23291 (N_23291,N_22803,N_22972);
or U23292 (N_23292,N_22868,N_22916);
xor U23293 (N_23293,N_22994,N_22143);
and U23294 (N_23294,N_22250,N_22443);
nand U23295 (N_23295,N_22810,N_22925);
or U23296 (N_23296,N_22461,N_22652);
xor U23297 (N_23297,N_22722,N_22987);
nor U23298 (N_23298,N_22152,N_22794);
and U23299 (N_23299,N_22843,N_22126);
nand U23300 (N_23300,N_22508,N_22640);
or U23301 (N_23301,N_22467,N_22882);
and U23302 (N_23302,N_22924,N_22145);
nand U23303 (N_23303,N_22598,N_22808);
nor U23304 (N_23304,N_22717,N_22724);
and U23305 (N_23305,N_22661,N_22873);
nand U23306 (N_23306,N_22283,N_22802);
xor U23307 (N_23307,N_22202,N_22937);
and U23308 (N_23308,N_22078,N_22455);
nor U23309 (N_23309,N_22993,N_22415);
xnor U23310 (N_23310,N_22458,N_22381);
xor U23311 (N_23311,N_22239,N_22103);
nand U23312 (N_23312,N_22285,N_22171);
and U23313 (N_23313,N_22278,N_22541);
xnor U23314 (N_23314,N_22913,N_22432);
nand U23315 (N_23315,N_22339,N_22366);
nand U23316 (N_23316,N_22386,N_22101);
or U23317 (N_23317,N_22091,N_22350);
nand U23318 (N_23318,N_22697,N_22856);
nand U23319 (N_23319,N_22066,N_22512);
and U23320 (N_23320,N_22375,N_22763);
xnor U23321 (N_23321,N_22507,N_22140);
or U23322 (N_23322,N_22680,N_22337);
nand U23323 (N_23323,N_22518,N_22016);
nor U23324 (N_23324,N_22262,N_22558);
and U23325 (N_23325,N_22060,N_22156);
nand U23326 (N_23326,N_22219,N_22986);
xnor U23327 (N_23327,N_22528,N_22790);
xor U23328 (N_23328,N_22867,N_22758);
and U23329 (N_23329,N_22674,N_22685);
nand U23330 (N_23330,N_22797,N_22430);
and U23331 (N_23331,N_22005,N_22247);
or U23332 (N_23332,N_22965,N_22023);
nand U23333 (N_23333,N_22138,N_22998);
xor U23334 (N_23334,N_22482,N_22130);
xnor U23335 (N_23335,N_22108,N_22233);
xor U23336 (N_23336,N_22274,N_22235);
or U23337 (N_23337,N_22297,N_22948);
nand U23338 (N_23338,N_22733,N_22690);
xnor U23339 (N_23339,N_22955,N_22721);
or U23340 (N_23340,N_22456,N_22270);
and U23341 (N_23341,N_22112,N_22256);
and U23342 (N_23342,N_22575,N_22783);
nor U23343 (N_23343,N_22220,N_22008);
or U23344 (N_23344,N_22927,N_22550);
xor U23345 (N_23345,N_22227,N_22292);
or U23346 (N_23346,N_22241,N_22020);
nand U23347 (N_23347,N_22237,N_22062);
xor U23348 (N_23348,N_22582,N_22900);
xnor U23349 (N_23349,N_22533,N_22954);
or U23350 (N_23350,N_22637,N_22141);
nor U23351 (N_23351,N_22753,N_22567);
and U23352 (N_23352,N_22826,N_22840);
and U23353 (N_23353,N_22402,N_22186);
or U23354 (N_23354,N_22190,N_22749);
xnor U23355 (N_23355,N_22835,N_22985);
and U23356 (N_23356,N_22757,N_22653);
nor U23357 (N_23357,N_22973,N_22165);
xor U23358 (N_23358,N_22117,N_22805);
or U23359 (N_23359,N_22574,N_22267);
nand U23360 (N_23360,N_22936,N_22881);
nand U23361 (N_23361,N_22499,N_22543);
and U23362 (N_23362,N_22476,N_22463);
and U23363 (N_23363,N_22319,N_22391);
or U23364 (N_23364,N_22034,N_22626);
or U23365 (N_23365,N_22650,N_22188);
or U23366 (N_23366,N_22831,N_22183);
or U23367 (N_23367,N_22468,N_22609);
or U23368 (N_23368,N_22473,N_22562);
and U23369 (N_23369,N_22229,N_22782);
xnor U23370 (N_23370,N_22962,N_22971);
xor U23371 (N_23371,N_22179,N_22132);
xnor U23372 (N_23372,N_22439,N_22714);
and U23373 (N_23373,N_22872,N_22511);
nor U23374 (N_23374,N_22080,N_22096);
nand U23375 (N_23375,N_22295,N_22917);
and U23376 (N_23376,N_22093,N_22111);
or U23377 (N_23377,N_22082,N_22086);
nor U23378 (N_23378,N_22081,N_22813);
and U23379 (N_23379,N_22039,N_22738);
nor U23380 (N_23380,N_22731,N_22895);
and U23381 (N_23381,N_22099,N_22452);
and U23382 (N_23382,N_22799,N_22323);
and U23383 (N_23383,N_22833,N_22289);
nor U23384 (N_23384,N_22854,N_22785);
and U23385 (N_23385,N_22056,N_22170);
xnor U23386 (N_23386,N_22444,N_22119);
and U23387 (N_23387,N_22427,N_22365);
nand U23388 (N_23388,N_22571,N_22982);
nand U23389 (N_23389,N_22527,N_22326);
nor U23390 (N_23390,N_22560,N_22251);
or U23391 (N_23391,N_22314,N_22036);
and U23392 (N_23392,N_22025,N_22870);
and U23393 (N_23393,N_22967,N_22294);
xnor U23394 (N_23394,N_22069,N_22351);
xnor U23395 (N_23395,N_22057,N_22032);
or U23396 (N_23396,N_22788,N_22484);
nand U23397 (N_23397,N_22730,N_22345);
or U23398 (N_23398,N_22691,N_22526);
xnor U23399 (N_23399,N_22807,N_22502);
and U23400 (N_23400,N_22874,N_22976);
xnor U23401 (N_23401,N_22694,N_22441);
or U23402 (N_23402,N_22254,N_22968);
nand U23403 (N_23403,N_22149,N_22536);
xor U23404 (N_23404,N_22321,N_22392);
or U23405 (N_23405,N_22465,N_22109);
or U23406 (N_23406,N_22494,N_22769);
nor U23407 (N_23407,N_22648,N_22180);
nor U23408 (N_23408,N_22037,N_22638);
and U23409 (N_23409,N_22630,N_22601);
nor U23410 (N_23410,N_22464,N_22195);
nand U23411 (N_23411,N_22120,N_22964);
nand U23412 (N_23412,N_22774,N_22832);
nand U23413 (N_23413,N_22901,N_22004);
nand U23414 (N_23414,N_22945,N_22451);
and U23415 (N_23415,N_22031,N_22645);
xor U23416 (N_23416,N_22979,N_22634);
nor U23417 (N_23417,N_22520,N_22857);
and U23418 (N_23418,N_22328,N_22615);
and U23419 (N_23419,N_22624,N_22534);
or U23420 (N_23420,N_22309,N_22559);
xor U23421 (N_23421,N_22182,N_22606);
and U23422 (N_23422,N_22406,N_22498);
or U23423 (N_23423,N_22151,N_22865);
xnor U23424 (N_23424,N_22299,N_22605);
xor U23425 (N_23425,N_22002,N_22818);
or U23426 (N_23426,N_22839,N_22061);
and U23427 (N_23427,N_22646,N_22493);
or U23428 (N_23428,N_22073,N_22516);
or U23429 (N_23429,N_22530,N_22847);
or U23430 (N_23430,N_22211,N_22477);
nand U23431 (N_23431,N_22385,N_22371);
nor U23432 (N_23432,N_22413,N_22144);
nand U23433 (N_23433,N_22147,N_22703);
or U23434 (N_23434,N_22376,N_22480);
and U23435 (N_23435,N_22474,N_22450);
and U23436 (N_23436,N_22092,N_22197);
nand U23437 (N_23437,N_22040,N_22272);
and U23438 (N_23438,N_22264,N_22779);
or U23439 (N_23439,N_22225,N_22975);
or U23440 (N_23440,N_22356,N_22205);
xnor U23441 (N_23441,N_22682,N_22792);
or U23442 (N_23442,N_22858,N_22644);
xnor U23443 (N_23443,N_22496,N_22305);
or U23444 (N_23444,N_22935,N_22357);
nand U23445 (N_23445,N_22671,N_22665);
xnor U23446 (N_23446,N_22306,N_22633);
or U23447 (N_23447,N_22478,N_22495);
nor U23448 (N_23448,N_22416,N_22279);
xnor U23449 (N_23449,N_22184,N_22106);
or U23450 (N_23450,N_22055,N_22765);
or U23451 (N_23451,N_22557,N_22411);
nor U23452 (N_23452,N_22435,N_22751);
xnor U23453 (N_23453,N_22772,N_22611);
or U23454 (N_23454,N_22529,N_22969);
or U23455 (N_23455,N_22322,N_22829);
and U23456 (N_23456,N_22908,N_22076);
or U23457 (N_23457,N_22657,N_22517);
xor U23458 (N_23458,N_22950,N_22616);
and U23459 (N_23459,N_22767,N_22363);
or U23460 (N_23460,N_22521,N_22693);
xor U23461 (N_23461,N_22269,N_22058);
nand U23462 (N_23462,N_22033,N_22736);
xnor U23463 (N_23463,N_22317,N_22164);
nand U23464 (N_23464,N_22318,N_22043);
and U23465 (N_23465,N_22485,N_22531);
xnor U23466 (N_23466,N_22354,N_22489);
or U23467 (N_23467,N_22095,N_22050);
nor U23468 (N_23468,N_22447,N_22931);
nand U23469 (N_23469,N_22077,N_22796);
xor U23470 (N_23470,N_22555,N_22855);
nand U23471 (N_23471,N_22001,N_22756);
nand U23472 (N_23472,N_22504,N_22497);
nor U23473 (N_23473,N_22041,N_22786);
xnor U23474 (N_23474,N_22105,N_22059);
or U23475 (N_23475,N_22943,N_22538);
or U23476 (N_23476,N_22118,N_22383);
or U23477 (N_23477,N_22585,N_22079);
or U23478 (N_23478,N_22761,N_22878);
nand U23479 (N_23479,N_22532,N_22014);
nand U23480 (N_23480,N_22806,N_22134);
or U23481 (N_23481,N_22382,N_22580);
nor U23482 (N_23482,N_22048,N_22850);
nand U23483 (N_23483,N_22614,N_22221);
nor U23484 (N_23484,N_22380,N_22128);
and U23485 (N_23485,N_22462,N_22561);
or U23486 (N_23486,N_22686,N_22346);
nand U23487 (N_23487,N_22777,N_22710);
and U23488 (N_23488,N_22483,N_22711);
nor U23489 (N_23489,N_22746,N_22586);
or U23490 (N_23490,N_22737,N_22260);
xor U23491 (N_23491,N_22136,N_22539);
or U23492 (N_23492,N_22214,N_22293);
or U23493 (N_23493,N_22100,N_22115);
or U23494 (N_23494,N_22537,N_22089);
and U23495 (N_23495,N_22748,N_22619);
or U23496 (N_23496,N_22249,N_22469);
nand U23497 (N_23497,N_22302,N_22022);
xnor U23498 (N_23498,N_22397,N_22446);
xnor U23499 (N_23499,N_22928,N_22990);
nor U23500 (N_23500,N_22409,N_22121);
and U23501 (N_23501,N_22589,N_22459);
nor U23502 (N_23502,N_22952,N_22526);
nor U23503 (N_23503,N_22923,N_22883);
xnor U23504 (N_23504,N_22141,N_22170);
nand U23505 (N_23505,N_22141,N_22502);
nor U23506 (N_23506,N_22406,N_22328);
nand U23507 (N_23507,N_22411,N_22843);
or U23508 (N_23508,N_22313,N_22627);
xnor U23509 (N_23509,N_22699,N_22089);
xor U23510 (N_23510,N_22684,N_22377);
or U23511 (N_23511,N_22401,N_22112);
nand U23512 (N_23512,N_22601,N_22645);
or U23513 (N_23513,N_22316,N_22491);
nand U23514 (N_23514,N_22356,N_22704);
or U23515 (N_23515,N_22437,N_22597);
or U23516 (N_23516,N_22710,N_22794);
or U23517 (N_23517,N_22653,N_22983);
nand U23518 (N_23518,N_22605,N_22146);
or U23519 (N_23519,N_22336,N_22191);
and U23520 (N_23520,N_22137,N_22044);
or U23521 (N_23521,N_22714,N_22755);
nand U23522 (N_23522,N_22607,N_22930);
xnor U23523 (N_23523,N_22448,N_22122);
xor U23524 (N_23524,N_22240,N_22220);
or U23525 (N_23525,N_22200,N_22783);
nor U23526 (N_23526,N_22216,N_22934);
or U23527 (N_23527,N_22691,N_22945);
nor U23528 (N_23528,N_22376,N_22481);
nor U23529 (N_23529,N_22629,N_22655);
or U23530 (N_23530,N_22122,N_22584);
nand U23531 (N_23531,N_22629,N_22021);
and U23532 (N_23532,N_22928,N_22479);
nand U23533 (N_23533,N_22693,N_22698);
xnor U23534 (N_23534,N_22962,N_22360);
nor U23535 (N_23535,N_22634,N_22580);
or U23536 (N_23536,N_22342,N_22808);
or U23537 (N_23537,N_22828,N_22311);
or U23538 (N_23538,N_22935,N_22436);
nor U23539 (N_23539,N_22333,N_22764);
nor U23540 (N_23540,N_22367,N_22871);
or U23541 (N_23541,N_22558,N_22858);
nand U23542 (N_23542,N_22338,N_22550);
xnor U23543 (N_23543,N_22806,N_22878);
or U23544 (N_23544,N_22949,N_22417);
xor U23545 (N_23545,N_22707,N_22649);
xor U23546 (N_23546,N_22030,N_22851);
nor U23547 (N_23547,N_22503,N_22407);
nor U23548 (N_23548,N_22921,N_22881);
nand U23549 (N_23549,N_22199,N_22219);
or U23550 (N_23550,N_22299,N_22026);
nand U23551 (N_23551,N_22496,N_22975);
or U23552 (N_23552,N_22951,N_22253);
nand U23553 (N_23553,N_22016,N_22575);
nand U23554 (N_23554,N_22789,N_22707);
nor U23555 (N_23555,N_22237,N_22522);
xnor U23556 (N_23556,N_22341,N_22342);
or U23557 (N_23557,N_22005,N_22681);
and U23558 (N_23558,N_22838,N_22190);
and U23559 (N_23559,N_22973,N_22564);
nand U23560 (N_23560,N_22803,N_22990);
xor U23561 (N_23561,N_22284,N_22505);
xor U23562 (N_23562,N_22615,N_22270);
nand U23563 (N_23563,N_22150,N_22678);
nor U23564 (N_23564,N_22466,N_22572);
or U23565 (N_23565,N_22268,N_22864);
or U23566 (N_23566,N_22207,N_22761);
or U23567 (N_23567,N_22913,N_22206);
nand U23568 (N_23568,N_22926,N_22728);
xnor U23569 (N_23569,N_22114,N_22533);
nor U23570 (N_23570,N_22003,N_22293);
nand U23571 (N_23571,N_22081,N_22799);
xor U23572 (N_23572,N_22544,N_22259);
nand U23573 (N_23573,N_22341,N_22550);
and U23574 (N_23574,N_22479,N_22225);
nand U23575 (N_23575,N_22091,N_22107);
and U23576 (N_23576,N_22534,N_22455);
and U23577 (N_23577,N_22917,N_22241);
nor U23578 (N_23578,N_22629,N_22433);
nor U23579 (N_23579,N_22102,N_22224);
nand U23580 (N_23580,N_22345,N_22050);
or U23581 (N_23581,N_22667,N_22282);
nand U23582 (N_23582,N_22619,N_22084);
and U23583 (N_23583,N_22428,N_22554);
nor U23584 (N_23584,N_22871,N_22736);
xnor U23585 (N_23585,N_22768,N_22826);
xnor U23586 (N_23586,N_22563,N_22401);
xnor U23587 (N_23587,N_22151,N_22492);
nor U23588 (N_23588,N_22690,N_22314);
nor U23589 (N_23589,N_22892,N_22727);
nand U23590 (N_23590,N_22237,N_22806);
xnor U23591 (N_23591,N_22982,N_22541);
nand U23592 (N_23592,N_22616,N_22669);
xor U23593 (N_23593,N_22130,N_22117);
xor U23594 (N_23594,N_22758,N_22256);
or U23595 (N_23595,N_22260,N_22886);
or U23596 (N_23596,N_22605,N_22014);
nor U23597 (N_23597,N_22331,N_22336);
or U23598 (N_23598,N_22562,N_22731);
xnor U23599 (N_23599,N_22433,N_22354);
and U23600 (N_23600,N_22249,N_22854);
xor U23601 (N_23601,N_22062,N_22567);
or U23602 (N_23602,N_22983,N_22601);
and U23603 (N_23603,N_22914,N_22622);
or U23604 (N_23604,N_22693,N_22139);
or U23605 (N_23605,N_22349,N_22216);
or U23606 (N_23606,N_22545,N_22614);
and U23607 (N_23607,N_22186,N_22287);
and U23608 (N_23608,N_22364,N_22223);
or U23609 (N_23609,N_22750,N_22002);
nand U23610 (N_23610,N_22214,N_22274);
nand U23611 (N_23611,N_22069,N_22262);
nand U23612 (N_23612,N_22805,N_22162);
nor U23613 (N_23613,N_22407,N_22054);
xor U23614 (N_23614,N_22404,N_22496);
and U23615 (N_23615,N_22213,N_22137);
nor U23616 (N_23616,N_22182,N_22353);
and U23617 (N_23617,N_22885,N_22397);
and U23618 (N_23618,N_22770,N_22560);
xor U23619 (N_23619,N_22478,N_22084);
nor U23620 (N_23620,N_22136,N_22739);
or U23621 (N_23621,N_22438,N_22065);
or U23622 (N_23622,N_22119,N_22631);
xor U23623 (N_23623,N_22652,N_22789);
nor U23624 (N_23624,N_22708,N_22712);
or U23625 (N_23625,N_22768,N_22932);
nor U23626 (N_23626,N_22365,N_22605);
or U23627 (N_23627,N_22520,N_22239);
and U23628 (N_23628,N_22414,N_22903);
or U23629 (N_23629,N_22786,N_22398);
xnor U23630 (N_23630,N_22181,N_22410);
xor U23631 (N_23631,N_22535,N_22120);
and U23632 (N_23632,N_22883,N_22484);
or U23633 (N_23633,N_22891,N_22884);
and U23634 (N_23634,N_22080,N_22036);
or U23635 (N_23635,N_22852,N_22526);
and U23636 (N_23636,N_22864,N_22772);
or U23637 (N_23637,N_22568,N_22360);
xor U23638 (N_23638,N_22714,N_22214);
or U23639 (N_23639,N_22476,N_22353);
xnor U23640 (N_23640,N_22570,N_22216);
xor U23641 (N_23641,N_22976,N_22744);
or U23642 (N_23642,N_22625,N_22330);
or U23643 (N_23643,N_22365,N_22774);
nand U23644 (N_23644,N_22947,N_22685);
nor U23645 (N_23645,N_22998,N_22512);
nand U23646 (N_23646,N_22633,N_22833);
and U23647 (N_23647,N_22378,N_22093);
and U23648 (N_23648,N_22339,N_22324);
and U23649 (N_23649,N_22995,N_22868);
nand U23650 (N_23650,N_22183,N_22363);
xor U23651 (N_23651,N_22800,N_22507);
and U23652 (N_23652,N_22642,N_22002);
or U23653 (N_23653,N_22991,N_22990);
xor U23654 (N_23654,N_22046,N_22182);
or U23655 (N_23655,N_22778,N_22131);
nor U23656 (N_23656,N_22994,N_22762);
nor U23657 (N_23657,N_22366,N_22842);
nor U23658 (N_23658,N_22236,N_22107);
or U23659 (N_23659,N_22266,N_22275);
and U23660 (N_23660,N_22654,N_22027);
nor U23661 (N_23661,N_22896,N_22586);
nand U23662 (N_23662,N_22421,N_22916);
and U23663 (N_23663,N_22380,N_22482);
nand U23664 (N_23664,N_22542,N_22710);
nand U23665 (N_23665,N_22442,N_22587);
nor U23666 (N_23666,N_22556,N_22582);
nor U23667 (N_23667,N_22907,N_22058);
or U23668 (N_23668,N_22264,N_22409);
or U23669 (N_23669,N_22822,N_22178);
xor U23670 (N_23670,N_22071,N_22049);
nor U23671 (N_23671,N_22323,N_22350);
and U23672 (N_23672,N_22900,N_22237);
nor U23673 (N_23673,N_22378,N_22540);
or U23674 (N_23674,N_22958,N_22426);
or U23675 (N_23675,N_22475,N_22511);
or U23676 (N_23676,N_22570,N_22469);
or U23677 (N_23677,N_22753,N_22404);
nand U23678 (N_23678,N_22300,N_22535);
nor U23679 (N_23679,N_22007,N_22890);
nor U23680 (N_23680,N_22118,N_22168);
or U23681 (N_23681,N_22738,N_22368);
nor U23682 (N_23682,N_22256,N_22269);
or U23683 (N_23683,N_22849,N_22188);
nor U23684 (N_23684,N_22999,N_22524);
xnor U23685 (N_23685,N_22446,N_22277);
and U23686 (N_23686,N_22496,N_22761);
nor U23687 (N_23687,N_22887,N_22304);
and U23688 (N_23688,N_22287,N_22647);
nand U23689 (N_23689,N_22601,N_22499);
or U23690 (N_23690,N_22776,N_22625);
nor U23691 (N_23691,N_22786,N_22929);
or U23692 (N_23692,N_22931,N_22297);
nor U23693 (N_23693,N_22866,N_22943);
or U23694 (N_23694,N_22326,N_22122);
nor U23695 (N_23695,N_22315,N_22427);
and U23696 (N_23696,N_22715,N_22392);
nor U23697 (N_23697,N_22808,N_22077);
and U23698 (N_23698,N_22960,N_22837);
nand U23699 (N_23699,N_22775,N_22958);
xnor U23700 (N_23700,N_22309,N_22596);
nand U23701 (N_23701,N_22263,N_22939);
xnor U23702 (N_23702,N_22716,N_22677);
nor U23703 (N_23703,N_22175,N_22828);
nand U23704 (N_23704,N_22306,N_22595);
and U23705 (N_23705,N_22162,N_22014);
nor U23706 (N_23706,N_22065,N_22639);
nor U23707 (N_23707,N_22495,N_22750);
nor U23708 (N_23708,N_22633,N_22896);
nand U23709 (N_23709,N_22130,N_22494);
nor U23710 (N_23710,N_22668,N_22021);
xnor U23711 (N_23711,N_22579,N_22795);
xor U23712 (N_23712,N_22949,N_22254);
or U23713 (N_23713,N_22386,N_22973);
or U23714 (N_23714,N_22047,N_22452);
xnor U23715 (N_23715,N_22027,N_22174);
nor U23716 (N_23716,N_22069,N_22100);
nand U23717 (N_23717,N_22173,N_22452);
xor U23718 (N_23718,N_22840,N_22658);
xor U23719 (N_23719,N_22045,N_22143);
nor U23720 (N_23720,N_22317,N_22628);
nand U23721 (N_23721,N_22389,N_22410);
nor U23722 (N_23722,N_22154,N_22729);
nor U23723 (N_23723,N_22178,N_22400);
nand U23724 (N_23724,N_22316,N_22348);
and U23725 (N_23725,N_22935,N_22407);
xor U23726 (N_23726,N_22648,N_22079);
xor U23727 (N_23727,N_22430,N_22298);
nor U23728 (N_23728,N_22419,N_22123);
xor U23729 (N_23729,N_22084,N_22931);
nand U23730 (N_23730,N_22816,N_22961);
and U23731 (N_23731,N_22081,N_22794);
xor U23732 (N_23732,N_22968,N_22273);
and U23733 (N_23733,N_22429,N_22387);
xor U23734 (N_23734,N_22013,N_22726);
xor U23735 (N_23735,N_22605,N_22045);
xnor U23736 (N_23736,N_22645,N_22459);
and U23737 (N_23737,N_22997,N_22508);
nor U23738 (N_23738,N_22287,N_22078);
and U23739 (N_23739,N_22334,N_22941);
and U23740 (N_23740,N_22349,N_22878);
nor U23741 (N_23741,N_22015,N_22867);
and U23742 (N_23742,N_22149,N_22595);
nor U23743 (N_23743,N_22716,N_22235);
nand U23744 (N_23744,N_22758,N_22207);
nor U23745 (N_23745,N_22863,N_22289);
xor U23746 (N_23746,N_22277,N_22160);
nor U23747 (N_23747,N_22908,N_22140);
and U23748 (N_23748,N_22471,N_22794);
nor U23749 (N_23749,N_22671,N_22454);
xnor U23750 (N_23750,N_22959,N_22340);
xor U23751 (N_23751,N_22967,N_22053);
nand U23752 (N_23752,N_22884,N_22084);
or U23753 (N_23753,N_22766,N_22781);
xnor U23754 (N_23754,N_22483,N_22252);
nand U23755 (N_23755,N_22464,N_22789);
or U23756 (N_23756,N_22615,N_22799);
nand U23757 (N_23757,N_22929,N_22542);
or U23758 (N_23758,N_22467,N_22185);
nor U23759 (N_23759,N_22762,N_22004);
or U23760 (N_23760,N_22926,N_22883);
xor U23761 (N_23761,N_22085,N_22887);
and U23762 (N_23762,N_22602,N_22059);
nor U23763 (N_23763,N_22932,N_22091);
nand U23764 (N_23764,N_22829,N_22478);
and U23765 (N_23765,N_22462,N_22283);
nand U23766 (N_23766,N_22564,N_22220);
or U23767 (N_23767,N_22425,N_22770);
nor U23768 (N_23768,N_22979,N_22574);
and U23769 (N_23769,N_22026,N_22294);
nor U23770 (N_23770,N_22635,N_22738);
xnor U23771 (N_23771,N_22591,N_22060);
or U23772 (N_23772,N_22899,N_22094);
xor U23773 (N_23773,N_22583,N_22497);
xnor U23774 (N_23774,N_22779,N_22643);
xnor U23775 (N_23775,N_22174,N_22051);
nand U23776 (N_23776,N_22260,N_22053);
nor U23777 (N_23777,N_22118,N_22500);
xnor U23778 (N_23778,N_22320,N_22945);
or U23779 (N_23779,N_22005,N_22700);
xor U23780 (N_23780,N_22264,N_22171);
and U23781 (N_23781,N_22463,N_22489);
and U23782 (N_23782,N_22757,N_22438);
or U23783 (N_23783,N_22170,N_22780);
and U23784 (N_23784,N_22874,N_22581);
xor U23785 (N_23785,N_22761,N_22027);
nand U23786 (N_23786,N_22239,N_22797);
xnor U23787 (N_23787,N_22640,N_22843);
and U23788 (N_23788,N_22741,N_22052);
nand U23789 (N_23789,N_22279,N_22284);
and U23790 (N_23790,N_22981,N_22330);
or U23791 (N_23791,N_22278,N_22750);
nor U23792 (N_23792,N_22324,N_22543);
or U23793 (N_23793,N_22557,N_22963);
or U23794 (N_23794,N_22446,N_22324);
nor U23795 (N_23795,N_22772,N_22159);
nor U23796 (N_23796,N_22337,N_22202);
or U23797 (N_23797,N_22268,N_22756);
xnor U23798 (N_23798,N_22845,N_22410);
and U23799 (N_23799,N_22924,N_22502);
xnor U23800 (N_23800,N_22891,N_22676);
nand U23801 (N_23801,N_22274,N_22698);
xnor U23802 (N_23802,N_22755,N_22441);
or U23803 (N_23803,N_22941,N_22122);
nand U23804 (N_23804,N_22257,N_22239);
nor U23805 (N_23805,N_22995,N_22489);
nand U23806 (N_23806,N_22046,N_22913);
nand U23807 (N_23807,N_22416,N_22075);
and U23808 (N_23808,N_22261,N_22048);
or U23809 (N_23809,N_22843,N_22577);
xnor U23810 (N_23810,N_22654,N_22937);
or U23811 (N_23811,N_22073,N_22192);
nand U23812 (N_23812,N_22263,N_22736);
and U23813 (N_23813,N_22907,N_22148);
nand U23814 (N_23814,N_22885,N_22211);
nand U23815 (N_23815,N_22928,N_22815);
and U23816 (N_23816,N_22012,N_22898);
and U23817 (N_23817,N_22048,N_22106);
nand U23818 (N_23818,N_22817,N_22831);
or U23819 (N_23819,N_22899,N_22690);
nand U23820 (N_23820,N_22398,N_22763);
or U23821 (N_23821,N_22456,N_22371);
and U23822 (N_23822,N_22452,N_22376);
nand U23823 (N_23823,N_22422,N_22858);
nand U23824 (N_23824,N_22401,N_22969);
nand U23825 (N_23825,N_22940,N_22898);
or U23826 (N_23826,N_22368,N_22918);
xor U23827 (N_23827,N_22977,N_22422);
nand U23828 (N_23828,N_22778,N_22622);
or U23829 (N_23829,N_22162,N_22590);
nand U23830 (N_23830,N_22481,N_22099);
and U23831 (N_23831,N_22772,N_22394);
xnor U23832 (N_23832,N_22315,N_22252);
or U23833 (N_23833,N_22507,N_22134);
xor U23834 (N_23834,N_22562,N_22388);
nand U23835 (N_23835,N_22373,N_22290);
nand U23836 (N_23836,N_22192,N_22521);
nor U23837 (N_23837,N_22041,N_22154);
or U23838 (N_23838,N_22777,N_22896);
xor U23839 (N_23839,N_22315,N_22146);
nor U23840 (N_23840,N_22668,N_22297);
xnor U23841 (N_23841,N_22996,N_22021);
nand U23842 (N_23842,N_22622,N_22539);
xnor U23843 (N_23843,N_22798,N_22138);
nor U23844 (N_23844,N_22830,N_22033);
nand U23845 (N_23845,N_22417,N_22407);
xnor U23846 (N_23846,N_22061,N_22226);
nor U23847 (N_23847,N_22459,N_22477);
and U23848 (N_23848,N_22439,N_22644);
nor U23849 (N_23849,N_22635,N_22346);
nor U23850 (N_23850,N_22484,N_22858);
or U23851 (N_23851,N_22510,N_22651);
or U23852 (N_23852,N_22731,N_22899);
and U23853 (N_23853,N_22168,N_22363);
nor U23854 (N_23854,N_22239,N_22488);
or U23855 (N_23855,N_22084,N_22681);
nand U23856 (N_23856,N_22188,N_22191);
xnor U23857 (N_23857,N_22995,N_22243);
or U23858 (N_23858,N_22389,N_22096);
nor U23859 (N_23859,N_22360,N_22904);
or U23860 (N_23860,N_22217,N_22046);
and U23861 (N_23861,N_22156,N_22777);
or U23862 (N_23862,N_22371,N_22479);
nand U23863 (N_23863,N_22584,N_22401);
nand U23864 (N_23864,N_22292,N_22838);
or U23865 (N_23865,N_22211,N_22819);
nor U23866 (N_23866,N_22260,N_22443);
and U23867 (N_23867,N_22829,N_22920);
and U23868 (N_23868,N_22340,N_22839);
and U23869 (N_23869,N_22230,N_22017);
xor U23870 (N_23870,N_22675,N_22222);
nor U23871 (N_23871,N_22977,N_22996);
nand U23872 (N_23872,N_22265,N_22594);
nor U23873 (N_23873,N_22212,N_22588);
nor U23874 (N_23874,N_22742,N_22777);
xnor U23875 (N_23875,N_22334,N_22556);
nand U23876 (N_23876,N_22847,N_22868);
nand U23877 (N_23877,N_22008,N_22223);
or U23878 (N_23878,N_22085,N_22937);
and U23879 (N_23879,N_22092,N_22403);
nor U23880 (N_23880,N_22294,N_22177);
or U23881 (N_23881,N_22847,N_22925);
xnor U23882 (N_23882,N_22758,N_22566);
nor U23883 (N_23883,N_22888,N_22258);
xnor U23884 (N_23884,N_22693,N_22336);
xor U23885 (N_23885,N_22103,N_22997);
or U23886 (N_23886,N_22009,N_22784);
and U23887 (N_23887,N_22741,N_22998);
nand U23888 (N_23888,N_22290,N_22453);
and U23889 (N_23889,N_22469,N_22473);
nor U23890 (N_23890,N_22481,N_22710);
xor U23891 (N_23891,N_22022,N_22149);
or U23892 (N_23892,N_22396,N_22402);
xor U23893 (N_23893,N_22963,N_22236);
nand U23894 (N_23894,N_22901,N_22116);
nand U23895 (N_23895,N_22744,N_22473);
xor U23896 (N_23896,N_22508,N_22227);
nor U23897 (N_23897,N_22294,N_22260);
xnor U23898 (N_23898,N_22355,N_22791);
nor U23899 (N_23899,N_22792,N_22996);
and U23900 (N_23900,N_22197,N_22399);
nor U23901 (N_23901,N_22736,N_22615);
nor U23902 (N_23902,N_22847,N_22774);
nor U23903 (N_23903,N_22595,N_22130);
nor U23904 (N_23904,N_22216,N_22177);
nand U23905 (N_23905,N_22261,N_22193);
nand U23906 (N_23906,N_22681,N_22302);
and U23907 (N_23907,N_22130,N_22569);
nor U23908 (N_23908,N_22412,N_22489);
or U23909 (N_23909,N_22886,N_22236);
xnor U23910 (N_23910,N_22672,N_22977);
nand U23911 (N_23911,N_22211,N_22642);
and U23912 (N_23912,N_22842,N_22900);
and U23913 (N_23913,N_22797,N_22803);
nand U23914 (N_23914,N_22610,N_22044);
nor U23915 (N_23915,N_22757,N_22309);
xnor U23916 (N_23916,N_22509,N_22470);
xor U23917 (N_23917,N_22647,N_22656);
or U23918 (N_23918,N_22546,N_22283);
xor U23919 (N_23919,N_22973,N_22281);
or U23920 (N_23920,N_22849,N_22118);
nor U23921 (N_23921,N_22492,N_22623);
nand U23922 (N_23922,N_22193,N_22606);
nand U23923 (N_23923,N_22051,N_22010);
or U23924 (N_23924,N_22474,N_22091);
nand U23925 (N_23925,N_22167,N_22663);
or U23926 (N_23926,N_22592,N_22028);
or U23927 (N_23927,N_22015,N_22516);
nor U23928 (N_23928,N_22267,N_22166);
or U23929 (N_23929,N_22161,N_22780);
nand U23930 (N_23930,N_22056,N_22091);
nand U23931 (N_23931,N_22988,N_22043);
xnor U23932 (N_23932,N_22042,N_22562);
and U23933 (N_23933,N_22602,N_22349);
xnor U23934 (N_23934,N_22827,N_22256);
xnor U23935 (N_23935,N_22988,N_22679);
nand U23936 (N_23936,N_22263,N_22586);
xor U23937 (N_23937,N_22691,N_22209);
and U23938 (N_23938,N_22333,N_22739);
xor U23939 (N_23939,N_22818,N_22498);
or U23940 (N_23940,N_22404,N_22470);
nand U23941 (N_23941,N_22327,N_22731);
nor U23942 (N_23942,N_22434,N_22500);
xnor U23943 (N_23943,N_22614,N_22483);
nor U23944 (N_23944,N_22412,N_22419);
nor U23945 (N_23945,N_22146,N_22197);
xor U23946 (N_23946,N_22942,N_22806);
nand U23947 (N_23947,N_22587,N_22825);
nand U23948 (N_23948,N_22183,N_22032);
or U23949 (N_23949,N_22092,N_22180);
or U23950 (N_23950,N_22674,N_22351);
xnor U23951 (N_23951,N_22157,N_22915);
xor U23952 (N_23952,N_22459,N_22158);
xor U23953 (N_23953,N_22897,N_22748);
nor U23954 (N_23954,N_22909,N_22380);
nor U23955 (N_23955,N_22826,N_22862);
and U23956 (N_23956,N_22849,N_22233);
or U23957 (N_23957,N_22230,N_22935);
and U23958 (N_23958,N_22219,N_22027);
nand U23959 (N_23959,N_22087,N_22502);
xnor U23960 (N_23960,N_22828,N_22168);
and U23961 (N_23961,N_22146,N_22745);
nor U23962 (N_23962,N_22714,N_22508);
nor U23963 (N_23963,N_22112,N_22195);
nand U23964 (N_23964,N_22013,N_22580);
or U23965 (N_23965,N_22283,N_22300);
nand U23966 (N_23966,N_22008,N_22935);
or U23967 (N_23967,N_22983,N_22470);
xnor U23968 (N_23968,N_22657,N_22019);
or U23969 (N_23969,N_22101,N_22377);
xnor U23970 (N_23970,N_22286,N_22421);
nand U23971 (N_23971,N_22279,N_22658);
xnor U23972 (N_23972,N_22490,N_22836);
nor U23973 (N_23973,N_22668,N_22370);
xor U23974 (N_23974,N_22441,N_22549);
nor U23975 (N_23975,N_22053,N_22878);
and U23976 (N_23976,N_22409,N_22593);
nor U23977 (N_23977,N_22659,N_22032);
or U23978 (N_23978,N_22334,N_22043);
xnor U23979 (N_23979,N_22151,N_22352);
or U23980 (N_23980,N_22658,N_22819);
nand U23981 (N_23981,N_22157,N_22141);
or U23982 (N_23982,N_22772,N_22708);
and U23983 (N_23983,N_22006,N_22271);
nand U23984 (N_23984,N_22347,N_22405);
nand U23985 (N_23985,N_22916,N_22655);
nor U23986 (N_23986,N_22358,N_22890);
nor U23987 (N_23987,N_22668,N_22028);
or U23988 (N_23988,N_22899,N_22745);
nor U23989 (N_23989,N_22330,N_22582);
or U23990 (N_23990,N_22550,N_22191);
xor U23991 (N_23991,N_22644,N_22153);
and U23992 (N_23992,N_22781,N_22655);
or U23993 (N_23993,N_22428,N_22991);
and U23994 (N_23994,N_22275,N_22722);
xor U23995 (N_23995,N_22244,N_22084);
nand U23996 (N_23996,N_22651,N_22668);
xor U23997 (N_23997,N_22130,N_22554);
or U23998 (N_23998,N_22308,N_22635);
and U23999 (N_23999,N_22039,N_22058);
xor U24000 (N_24000,N_23783,N_23047);
nand U24001 (N_24001,N_23504,N_23440);
and U24002 (N_24002,N_23277,N_23165);
nor U24003 (N_24003,N_23311,N_23028);
nor U24004 (N_24004,N_23167,N_23644);
and U24005 (N_24005,N_23323,N_23891);
nand U24006 (N_24006,N_23658,N_23979);
or U24007 (N_24007,N_23705,N_23577);
or U24008 (N_24008,N_23627,N_23254);
and U24009 (N_24009,N_23915,N_23987);
and U24010 (N_24010,N_23051,N_23843);
nor U24011 (N_24011,N_23411,N_23893);
nor U24012 (N_24012,N_23838,N_23150);
xor U24013 (N_24013,N_23276,N_23333);
nor U24014 (N_24014,N_23287,N_23490);
xor U24015 (N_24015,N_23770,N_23675);
nor U24016 (N_24016,N_23849,N_23721);
nor U24017 (N_24017,N_23753,N_23942);
or U24018 (N_24018,N_23236,N_23886);
xnor U24019 (N_24019,N_23757,N_23813);
and U24020 (N_24020,N_23861,N_23765);
nand U24021 (N_24021,N_23230,N_23322);
nor U24022 (N_24022,N_23061,N_23380);
xor U24023 (N_24023,N_23889,N_23772);
nand U24024 (N_24024,N_23596,N_23518);
xor U24025 (N_24025,N_23102,N_23828);
and U24026 (N_24026,N_23928,N_23089);
and U24027 (N_24027,N_23584,N_23586);
nor U24028 (N_24028,N_23187,N_23592);
and U24029 (N_24029,N_23677,N_23630);
and U24030 (N_24030,N_23858,N_23736);
and U24031 (N_24031,N_23695,N_23662);
and U24032 (N_24032,N_23067,N_23030);
and U24033 (N_24033,N_23052,N_23247);
and U24034 (N_24034,N_23379,N_23807);
xor U24035 (N_24035,N_23732,N_23399);
nor U24036 (N_24036,N_23501,N_23599);
or U24037 (N_24037,N_23727,N_23650);
nor U24038 (N_24038,N_23910,N_23718);
nor U24039 (N_24039,N_23010,N_23980);
xnor U24040 (N_24040,N_23958,N_23710);
or U24041 (N_24041,N_23222,N_23069);
xnor U24042 (N_24042,N_23213,N_23057);
xnor U24043 (N_24043,N_23713,N_23835);
and U24044 (N_24044,N_23972,N_23652);
xnor U24045 (N_24045,N_23781,N_23962);
xor U24046 (N_24046,N_23066,N_23912);
nand U24047 (N_24047,N_23110,N_23758);
nor U24048 (N_24048,N_23378,N_23500);
nand U24049 (N_24049,N_23376,N_23320);
and U24050 (N_24050,N_23166,N_23448);
nor U24051 (N_24051,N_23146,N_23220);
and U24052 (N_24052,N_23356,N_23523);
nor U24053 (N_24053,N_23265,N_23648);
nor U24054 (N_24054,N_23443,N_23528);
xnor U24055 (N_24055,N_23111,N_23293);
xor U24056 (N_24056,N_23649,N_23453);
xnor U24057 (N_24057,N_23105,N_23846);
nor U24058 (N_24058,N_23328,N_23216);
and U24059 (N_24059,N_23346,N_23198);
or U24060 (N_24060,N_23688,N_23903);
nor U24061 (N_24061,N_23839,N_23696);
xor U24062 (N_24062,N_23050,N_23970);
xnor U24063 (N_24063,N_23270,N_23574);
nand U24064 (N_24064,N_23459,N_23869);
xor U24065 (N_24065,N_23179,N_23336);
and U24066 (N_24066,N_23551,N_23963);
or U24067 (N_24067,N_23879,N_23918);
nor U24068 (N_24068,N_23759,N_23444);
xnor U24069 (N_24069,N_23654,N_23473);
and U24070 (N_24070,N_23898,N_23545);
nor U24071 (N_24071,N_23482,N_23000);
or U24072 (N_24072,N_23730,N_23507);
xnor U24073 (N_24073,N_23331,N_23941);
nor U24074 (N_24074,N_23286,N_23782);
nor U24075 (N_24075,N_23132,N_23771);
nand U24076 (N_24076,N_23920,N_23284);
nor U24077 (N_24077,N_23170,N_23197);
nand U24078 (N_24078,N_23568,N_23318);
nor U24079 (N_24079,N_23703,N_23123);
and U24080 (N_24080,N_23349,N_23168);
and U24081 (N_24081,N_23304,N_23257);
nand U24082 (N_24082,N_23496,N_23935);
or U24083 (N_24083,N_23946,N_23321);
or U24084 (N_24084,N_23725,N_23564);
and U24085 (N_24085,N_23086,N_23316);
and U24086 (N_24086,N_23904,N_23780);
nand U24087 (N_24087,N_23635,N_23206);
xor U24088 (N_24088,N_23458,N_23288);
nor U24089 (N_24089,N_23077,N_23735);
or U24090 (N_24090,N_23296,N_23715);
or U24091 (N_24091,N_23505,N_23743);
nor U24092 (N_24092,N_23285,N_23412);
and U24093 (N_24093,N_23668,N_23629);
and U24094 (N_24094,N_23711,N_23364);
xnor U24095 (N_24095,N_23188,N_23508);
and U24096 (N_24096,N_23945,N_23452);
and U24097 (N_24097,N_23626,N_23267);
or U24098 (N_24098,N_23387,N_23693);
nand U24099 (N_24099,N_23674,N_23957);
xnor U24100 (N_24100,N_23651,N_23618);
xor U24101 (N_24101,N_23552,N_23090);
and U24102 (N_24102,N_23157,N_23262);
xor U24103 (N_24103,N_23205,N_23347);
nor U24104 (N_24104,N_23064,N_23038);
nor U24105 (N_24105,N_23366,N_23788);
xor U24106 (N_24106,N_23542,N_23513);
or U24107 (N_24107,N_23082,N_23881);
nand U24108 (N_24108,N_23249,N_23424);
nand U24109 (N_24109,N_23553,N_23454);
nand U24110 (N_24110,N_23532,N_23215);
nor U24111 (N_24111,N_23613,N_23789);
xor U24112 (N_24112,N_23708,N_23680);
or U24113 (N_24113,N_23075,N_23340);
nor U24114 (N_24114,N_23522,N_23547);
nand U24115 (N_24115,N_23182,N_23095);
and U24116 (N_24116,N_23685,N_23998);
xnor U24117 (N_24117,N_23238,N_23569);
nor U24118 (N_24118,N_23139,N_23255);
nand U24119 (N_24119,N_23756,N_23745);
or U24120 (N_24120,N_23830,N_23422);
or U24121 (N_24121,N_23009,N_23791);
nand U24122 (N_24122,N_23423,N_23925);
or U24123 (N_24123,N_23327,N_23271);
or U24124 (N_24124,N_23384,N_23540);
or U24125 (N_24125,N_23659,N_23707);
xnor U24126 (N_24126,N_23991,N_23520);
or U24127 (N_24127,N_23931,N_23389);
xor U24128 (N_24128,N_23589,N_23397);
nand U24129 (N_24129,N_23479,N_23723);
xor U24130 (N_24130,N_23619,N_23905);
and U24131 (N_24131,N_23381,N_23140);
and U24132 (N_24132,N_23524,N_23663);
xnor U24133 (N_24133,N_23733,N_23609);
nor U24134 (N_24134,N_23750,N_23135);
nand U24135 (N_24135,N_23803,N_23022);
nand U24136 (N_24136,N_23023,N_23731);
and U24137 (N_24137,N_23907,N_23204);
and U24138 (N_24138,N_23591,N_23895);
nor U24139 (N_24139,N_23472,N_23307);
xnor U24140 (N_24140,N_23128,N_23840);
or U24141 (N_24141,N_23162,N_23386);
or U24142 (N_24142,N_23950,N_23447);
xor U24143 (N_24143,N_23543,N_23984);
and U24144 (N_24144,N_23094,N_23431);
or U24145 (N_24145,N_23786,N_23734);
or U24146 (N_24146,N_23144,N_23722);
or U24147 (N_24147,N_23449,N_23093);
or U24148 (N_24148,N_23434,N_23059);
xnor U24149 (N_24149,N_23938,N_23768);
nand U24150 (N_24150,N_23926,N_23622);
or U24151 (N_24151,N_23706,N_23872);
nor U24152 (N_24152,N_23235,N_23761);
nor U24153 (N_24153,N_23279,N_23796);
xnor U24154 (N_24154,N_23005,N_23360);
or U24155 (N_24155,N_23201,N_23002);
or U24156 (N_24156,N_23309,N_23421);
nor U24157 (N_24157,N_23887,N_23043);
nor U24158 (N_24158,N_23940,N_23274);
nor U24159 (N_24159,N_23410,N_23814);
nor U24160 (N_24160,N_23329,N_23643);
xor U24161 (N_24161,N_23019,N_23882);
xor U24162 (N_24162,N_23959,N_23572);
and U24163 (N_24163,N_23171,N_23754);
nor U24164 (N_24164,N_23704,N_23185);
and U24165 (N_24165,N_23875,N_23610);
nor U24166 (N_24166,N_23014,N_23679);
nor U24167 (N_24167,N_23106,N_23724);
or U24168 (N_24168,N_23314,N_23499);
and U24169 (N_24169,N_23967,N_23809);
or U24170 (N_24170,N_23633,N_23510);
and U24171 (N_24171,N_23250,N_23006);
or U24172 (N_24172,N_23163,N_23189);
nand U24173 (N_24173,N_23107,N_23243);
nor U24174 (N_24174,N_23597,N_23888);
nor U24175 (N_24175,N_23948,N_23719);
and U24176 (N_24176,N_23874,N_23978);
nor U24177 (N_24177,N_23600,N_23739);
nand U24178 (N_24178,N_23933,N_23308);
xor U24179 (N_24179,N_23969,N_23624);
nor U24180 (N_24180,N_23485,N_23837);
nand U24181 (N_24181,N_23604,N_23492);
or U24182 (N_24182,N_23549,N_23511);
and U24183 (N_24183,N_23008,N_23438);
xor U24184 (N_24184,N_23916,N_23819);
xnor U24185 (N_24185,N_23169,N_23048);
or U24186 (N_24186,N_23605,N_23363);
nand U24187 (N_24187,N_23425,N_23611);
or U24188 (N_24188,N_23103,N_23478);
or U24189 (N_24189,N_23088,N_23203);
nor U24190 (N_24190,N_23108,N_23986);
xor U24191 (N_24191,N_23784,N_23195);
or U24192 (N_24192,N_23176,N_23324);
and U24193 (N_24193,N_23681,N_23159);
nand U24194 (N_24194,N_23359,N_23369);
or U24195 (N_24195,N_23896,N_23289);
xnor U24196 (N_24196,N_23880,N_23717);
or U24197 (N_24197,N_23673,N_23689);
xor U24198 (N_24198,N_23080,N_23660);
or U24199 (N_24199,N_23665,N_23079);
and U24200 (N_24200,N_23924,N_23385);
xor U24201 (N_24201,N_23766,N_23615);
nand U24202 (N_24202,N_23350,N_23691);
or U24203 (N_24203,N_23032,N_23798);
nand U24204 (N_24204,N_23684,N_23152);
xor U24205 (N_24205,N_23183,N_23831);
nor U24206 (N_24206,N_23078,N_23617);
and U24207 (N_24207,N_23191,N_23337);
and U24208 (N_24208,N_23332,N_23313);
nand U24209 (N_24209,N_23842,N_23178);
xor U24210 (N_24210,N_23398,N_23427);
nand U24211 (N_24211,N_23252,N_23908);
nand U24212 (N_24212,N_23502,N_23538);
and U24213 (N_24213,N_23012,N_23729);
xor U24214 (N_24214,N_23446,N_23746);
and U24215 (N_24215,N_23177,N_23436);
and U24216 (N_24216,N_23973,N_23535);
or U24217 (N_24217,N_23667,N_23760);
and U24218 (N_24218,N_23368,N_23836);
nor U24219 (N_24219,N_23455,N_23180);
nor U24220 (N_24220,N_23039,N_23468);
and U24221 (N_24221,N_23025,N_23046);
xor U24222 (N_24222,N_23352,N_23581);
xnor U24223 (N_24223,N_23870,N_23792);
or U24224 (N_24224,N_23683,N_23943);
and U24225 (N_24225,N_23263,N_23141);
or U24226 (N_24226,N_23070,N_23575);
and U24227 (N_24227,N_23890,N_23126);
or U24228 (N_24228,N_23442,N_23147);
nor U24229 (N_24229,N_23860,N_23130);
xor U24230 (N_24230,N_23698,N_23391);
nand U24231 (N_24231,N_23606,N_23430);
or U24232 (N_24232,N_23037,N_23388);
or U24233 (N_24233,N_23525,N_23560);
xnor U24234 (N_24234,N_23602,N_23697);
nor U24235 (N_24235,N_23212,N_23001);
nor U24236 (N_24236,N_23608,N_23237);
or U24237 (N_24237,N_23671,N_23233);
nand U24238 (N_24238,N_23228,N_23994);
or U24239 (N_24239,N_23866,N_23993);
and U24240 (N_24240,N_23873,N_23432);
or U24241 (N_24241,N_23937,N_23865);
nand U24242 (N_24242,N_23416,N_23637);
nor U24243 (N_24243,N_23377,N_23361);
nand U24244 (N_24244,N_23628,N_23480);
and U24245 (N_24245,N_23983,N_23864);
and U24246 (N_24246,N_23848,N_23699);
and U24247 (N_24247,N_23300,N_23148);
or U24248 (N_24248,N_23342,N_23640);
and U24249 (N_24249,N_23700,N_23127);
nor U24250 (N_24250,N_23588,N_23260);
xnor U24251 (N_24251,N_23947,N_23244);
nand U24252 (N_24252,N_23227,N_23669);
or U24253 (N_24253,N_23471,N_23137);
nor U24254 (N_24254,N_23242,N_23767);
nand U24255 (N_24255,N_23884,N_23952);
or U24256 (N_24256,N_23119,N_23283);
nor U24257 (N_24257,N_23015,N_23623);
and U24258 (N_24258,N_23985,N_23229);
nand U24259 (N_24259,N_23405,N_23390);
nand U24260 (N_24260,N_23939,N_23799);
or U24261 (N_24261,N_23445,N_23871);
or U24262 (N_24262,N_23488,N_23544);
xor U24263 (N_24263,N_23330,N_23465);
and U24264 (N_24264,N_23122,N_23497);
or U24265 (N_24265,N_23738,N_23409);
xnor U24266 (N_24266,N_23394,N_23690);
xor U24267 (N_24267,N_23367,N_23625);
xor U24268 (N_24268,N_23184,N_23607);
xnor U24269 (N_24269,N_23614,N_23678);
xor U24270 (N_24270,N_23661,N_23060);
nand U24271 (N_24271,N_23529,N_23464);
xor U24272 (N_24272,N_23795,N_23083);
and U24273 (N_24273,N_23018,N_23702);
and U24274 (N_24274,N_23219,N_23259);
or U24275 (N_24275,N_23856,N_23011);
xnor U24276 (N_24276,N_23955,N_23261);
or U24277 (N_24277,N_23256,N_23463);
nand U24278 (N_24278,N_23805,N_23295);
xor U24279 (N_24279,N_23777,N_23997);
and U24280 (N_24280,N_23292,N_23003);
nand U24281 (N_24281,N_23407,N_23797);
nand U24282 (N_24282,N_23917,N_23016);
or U24283 (N_24283,N_23563,N_23902);
or U24284 (N_24284,N_23100,N_23826);
xnor U24285 (N_24285,N_23966,N_23214);
or U24286 (N_24286,N_23121,N_23031);
or U24287 (N_24287,N_23832,N_23234);
nor U24288 (N_24288,N_23598,N_23202);
nand U24289 (N_24289,N_23282,N_23561);
nand U24290 (N_24290,N_23192,N_23981);
nand U24291 (N_24291,N_23857,N_23196);
or U24292 (N_24292,N_23557,N_23071);
or U24293 (N_24293,N_23800,N_23694);
nor U24294 (N_24294,N_23855,N_23631);
and U24295 (N_24295,N_23634,N_23310);
nand U24296 (N_24296,N_23160,N_23526);
xor U24297 (N_24297,N_23466,N_23158);
and U24298 (N_24298,N_23720,N_23303);
and U24299 (N_24299,N_23960,N_23325);
xnor U24300 (N_24300,N_23049,N_23541);
or U24301 (N_24301,N_23469,N_23117);
and U24302 (N_24302,N_23503,N_23420);
nor U24303 (N_24303,N_23317,N_23531);
nand U24304 (N_24304,N_23672,N_23053);
or U24305 (N_24305,N_23403,N_23024);
and U24306 (N_24306,N_23116,N_23539);
nor U24307 (N_24307,N_23656,N_23120);
and U24308 (N_24308,N_23280,N_23045);
nand U24309 (N_24309,N_23491,N_23036);
nor U24310 (N_24310,N_23516,N_23749);
xor U24311 (N_24311,N_23583,N_23686);
or U24312 (N_24312,N_23245,N_23467);
and U24313 (N_24313,N_23537,N_23982);
nor U24314 (N_24314,N_23240,N_23919);
and U24315 (N_24315,N_23246,N_23820);
xnor U24316 (N_24316,N_23714,N_23850);
and U24317 (N_24317,N_23954,N_23748);
and U24318 (N_24318,N_23451,N_23475);
or U24319 (N_24319,N_23867,N_23210);
and U24320 (N_24320,N_23995,N_23272);
nor U24321 (N_24321,N_23305,N_23514);
or U24322 (N_24322,N_23224,N_23087);
nand U24323 (N_24323,N_23226,N_23223);
nor U24324 (N_24324,N_23033,N_23486);
or U24325 (N_24325,N_23319,N_23877);
nand U24326 (N_24326,N_23081,N_23460);
and U24327 (N_24327,N_23527,N_23818);
xnor U24328 (N_24328,N_23999,N_23124);
xnor U24329 (N_24329,N_23426,N_23161);
xor U24330 (N_24330,N_23221,N_23172);
nand U24331 (N_24331,N_23382,N_23841);
nand U24332 (N_24332,N_23362,N_23670);
nor U24333 (N_24333,N_23450,N_23134);
nand U24334 (N_24334,N_23021,N_23042);
xnor U24335 (N_24335,N_23776,N_23258);
nand U24336 (N_24336,N_23193,N_23775);
nand U24337 (N_24337,N_23554,N_23175);
or U24338 (N_24338,N_23774,N_23393);
and U24339 (N_24339,N_23834,N_23054);
nand U24340 (N_24340,N_23573,N_23461);
or U24341 (N_24341,N_23944,N_23199);
or U24342 (N_24342,N_23582,N_23810);
nand U24343 (N_24343,N_23457,N_23477);
xor U24344 (N_24344,N_23275,N_23603);
nand U24345 (N_24345,N_23248,N_23439);
xnor U24346 (N_24346,N_23716,N_23664);
or U24347 (N_24347,N_23441,N_23335);
xor U24348 (N_24348,N_23534,N_23164);
or U24349 (N_24349,N_23264,N_23136);
nand U24350 (N_24350,N_23533,N_23822);
nand U24351 (N_24351,N_23231,N_23092);
or U24352 (N_24352,N_23207,N_23211);
nand U24353 (N_24353,N_23026,N_23326);
or U24354 (N_24354,N_23580,N_23989);
nand U24355 (N_24355,N_23437,N_23827);
and U24356 (N_24356,N_23041,N_23433);
xor U24357 (N_24357,N_23358,N_23996);
xnor U24358 (N_24358,N_23676,N_23181);
nand U24359 (N_24359,N_23883,N_23934);
or U24360 (N_24360,N_23932,N_23536);
nand U24361 (N_24361,N_23899,N_23816);
nor U24362 (N_24362,N_23370,N_23063);
xor U24363 (N_24363,N_23506,N_23641);
xnor U24364 (N_24364,N_23922,N_23741);
xor U24365 (N_24365,N_23435,N_23341);
nor U24366 (N_24366,N_23965,N_23892);
nor U24367 (N_24367,N_23585,N_23709);
nand U24368 (N_24368,N_23914,N_23339);
xnor U24369 (N_24369,N_23555,N_23666);
nand U24370 (N_24370,N_23862,N_23894);
nor U24371 (N_24371,N_23956,N_23620);
xor U24372 (N_24372,N_23515,N_23737);
xor U24373 (N_24373,N_23811,N_23638);
or U24374 (N_24374,N_23821,N_23149);
nor U24375 (N_24375,N_23779,N_23901);
nand U24376 (N_24376,N_23692,N_23801);
and U24377 (N_24377,N_23155,N_23371);
and U24378 (N_24378,N_23595,N_23927);
and U24379 (N_24379,N_23118,N_23773);
nand U24380 (N_24380,N_23101,N_23273);
nand U24381 (N_24381,N_23470,N_23373);
nor U24382 (N_24382,N_23129,N_23400);
xnor U24383 (N_24383,N_23383,N_23241);
xor U24384 (N_24384,N_23131,N_23936);
nand U24385 (N_24385,N_23639,N_23930);
xor U24386 (N_24386,N_23571,N_23351);
xor U24387 (N_24387,N_23406,N_23074);
xnor U24388 (N_24388,N_23530,N_23302);
nand U24389 (N_24389,N_23290,N_23949);
nor U24390 (N_24390,N_23402,N_23755);
and U24391 (N_24391,N_23790,N_23806);
nor U24392 (N_24392,N_23851,N_23298);
or U24393 (N_24393,N_23401,N_23594);
and U24394 (N_24394,N_23190,N_23853);
xor U24395 (N_24395,N_23209,N_23417);
or U24396 (N_24396,N_23493,N_23897);
or U24397 (N_24397,N_23239,N_23815);
and U24398 (N_24398,N_23113,N_23044);
or U24399 (N_24399,N_23808,N_23253);
and U24400 (N_24400,N_23096,N_23621);
or U24401 (N_24401,N_23115,N_23751);
and U24402 (N_24402,N_23072,N_23977);
or U24403 (N_24403,N_23601,N_23353);
nand U24404 (N_24404,N_23194,N_23173);
nor U24405 (N_24405,N_23007,N_23097);
xnor U24406 (N_24406,N_23909,N_23567);
nand U24407 (N_24407,N_23812,N_23975);
or U24408 (N_24408,N_23566,N_23374);
or U24409 (N_24409,N_23900,N_23268);
and U24410 (N_24410,N_23104,N_23845);
nor U24411 (N_24411,N_23740,N_23953);
nand U24412 (N_24412,N_23712,N_23348);
nand U24413 (N_24413,N_23186,N_23114);
nor U24414 (N_24414,N_23578,N_23065);
xnor U24415 (N_24415,N_23392,N_23653);
xor U24416 (N_24416,N_23225,N_23804);
xor U24417 (N_24417,N_23312,N_23546);
xor U24418 (N_24418,N_23297,N_23034);
nor U24419 (N_24419,N_23232,N_23429);
or U24420 (N_24420,N_23109,N_23084);
and U24421 (N_24421,N_23266,N_23579);
nand U24422 (N_24422,N_23971,N_23817);
xor U24423 (N_24423,N_23073,N_23301);
nand U24424 (N_24424,N_23404,N_23414);
nand U24425 (N_24425,N_23833,N_23876);
nor U24426 (N_24426,N_23787,N_23138);
and U24427 (N_24427,N_23612,N_23481);
nand U24428 (N_24428,N_23825,N_23415);
xnor U24429 (N_24429,N_23657,N_23512);
or U24430 (N_24430,N_23988,N_23112);
and U24431 (N_24431,N_23587,N_23418);
and U24432 (N_24432,N_23921,N_23847);
xnor U24433 (N_24433,N_23099,N_23153);
nand U24434 (N_24434,N_23055,N_23778);
or U24435 (N_24435,N_23728,N_23408);
nor U24436 (N_24436,N_23278,N_23474);
and U24437 (N_24437,N_23682,N_23854);
or U24438 (N_24438,N_23769,N_23154);
nor U24439 (N_24439,N_23911,N_23593);
nor U24440 (N_24440,N_23027,N_23085);
nand U24441 (N_24441,N_23004,N_23484);
nand U24442 (N_24442,N_23143,N_23785);
and U24443 (N_24443,N_23156,N_23646);
xnor U24444 (N_24444,N_23419,N_23040);
or U24445 (N_24445,N_23519,N_23558);
xor U24446 (N_24446,N_23726,N_23752);
and U24447 (N_24447,N_23636,N_23396);
nor U24448 (N_24448,N_23456,N_23823);
or U24449 (N_24449,N_23294,N_23334);
or U24450 (N_24450,N_23763,N_23035);
nand U24451 (N_24451,N_23961,N_23133);
and U24452 (N_24452,N_23562,N_23372);
nor U24453 (N_24453,N_23647,N_23565);
xor U24454 (N_24454,N_23550,N_23852);
nor U24455 (N_24455,N_23906,N_23489);
xor U24456 (N_24456,N_23345,N_23824);
xor U24457 (N_24457,N_23844,N_23576);
nand U24458 (N_24458,N_23992,N_23687);
nand U24459 (N_24459,N_23570,N_23747);
xnor U24460 (N_24460,N_23616,N_23125);
and U24461 (N_24461,N_23964,N_23794);
nor U24462 (N_24462,N_23645,N_23968);
nand U24463 (N_24463,N_23291,N_23338);
or U24464 (N_24464,N_23476,N_23357);
and U24465 (N_24465,N_23483,N_23174);
and U24466 (N_24466,N_23029,N_23375);
and U24467 (N_24467,N_23218,N_23642);
nand U24468 (N_24468,N_23487,N_23354);
xor U24469 (N_24469,N_23521,N_23517);
nor U24470 (N_24470,N_23868,N_23017);
and U24471 (N_24471,N_23913,N_23098);
and U24472 (N_24472,N_23655,N_23269);
xor U24473 (N_24473,N_23548,N_23142);
xor U24474 (N_24474,N_23923,N_23863);
nor U24475 (N_24475,N_23462,N_23701);
and U24476 (N_24476,N_23020,N_23974);
xnor U24477 (N_24477,N_23306,N_23764);
and U24478 (N_24478,N_23878,N_23281);
or U24479 (N_24479,N_23344,N_23056);
and U24480 (N_24480,N_23509,N_23299);
nand U24481 (N_24481,N_23744,N_23395);
or U24482 (N_24482,N_23802,N_23151);
and U24483 (N_24483,N_23076,N_23976);
nand U24484 (N_24484,N_23343,N_23951);
nor U24485 (N_24485,N_23885,N_23929);
xnor U24486 (N_24486,N_23428,N_23145);
xnor U24487 (N_24487,N_23590,N_23495);
xor U24488 (N_24488,N_23632,N_23251);
xor U24489 (N_24489,N_23091,N_23062);
and U24490 (N_24490,N_23315,N_23365);
xnor U24491 (N_24491,N_23058,N_23013);
nand U24492 (N_24492,N_23498,N_23413);
nand U24493 (N_24493,N_23793,N_23217);
or U24494 (N_24494,N_23200,N_23556);
nor U24495 (N_24495,N_23859,N_23208);
xnor U24496 (N_24496,N_23068,N_23559);
nor U24497 (N_24497,N_23829,N_23742);
nand U24498 (N_24498,N_23355,N_23494);
or U24499 (N_24499,N_23990,N_23762);
nand U24500 (N_24500,N_23817,N_23811);
nand U24501 (N_24501,N_23838,N_23241);
and U24502 (N_24502,N_23296,N_23000);
nand U24503 (N_24503,N_23411,N_23086);
nor U24504 (N_24504,N_23932,N_23060);
and U24505 (N_24505,N_23135,N_23033);
nand U24506 (N_24506,N_23811,N_23013);
nand U24507 (N_24507,N_23900,N_23716);
and U24508 (N_24508,N_23034,N_23115);
and U24509 (N_24509,N_23312,N_23531);
and U24510 (N_24510,N_23424,N_23202);
xnor U24511 (N_24511,N_23396,N_23709);
or U24512 (N_24512,N_23630,N_23567);
or U24513 (N_24513,N_23560,N_23248);
or U24514 (N_24514,N_23986,N_23004);
nor U24515 (N_24515,N_23298,N_23879);
and U24516 (N_24516,N_23757,N_23019);
and U24517 (N_24517,N_23300,N_23062);
or U24518 (N_24518,N_23044,N_23559);
nand U24519 (N_24519,N_23631,N_23129);
and U24520 (N_24520,N_23951,N_23940);
or U24521 (N_24521,N_23916,N_23496);
nor U24522 (N_24522,N_23962,N_23720);
nor U24523 (N_24523,N_23950,N_23542);
and U24524 (N_24524,N_23930,N_23616);
or U24525 (N_24525,N_23394,N_23045);
and U24526 (N_24526,N_23680,N_23010);
or U24527 (N_24527,N_23776,N_23803);
xor U24528 (N_24528,N_23819,N_23734);
and U24529 (N_24529,N_23672,N_23071);
nor U24530 (N_24530,N_23471,N_23642);
nor U24531 (N_24531,N_23521,N_23557);
xor U24532 (N_24532,N_23878,N_23206);
and U24533 (N_24533,N_23917,N_23440);
nor U24534 (N_24534,N_23195,N_23221);
or U24535 (N_24535,N_23065,N_23259);
nand U24536 (N_24536,N_23843,N_23008);
xor U24537 (N_24537,N_23782,N_23762);
nor U24538 (N_24538,N_23282,N_23457);
nor U24539 (N_24539,N_23899,N_23987);
and U24540 (N_24540,N_23254,N_23328);
xor U24541 (N_24541,N_23967,N_23024);
or U24542 (N_24542,N_23475,N_23524);
nor U24543 (N_24543,N_23532,N_23439);
or U24544 (N_24544,N_23718,N_23397);
xnor U24545 (N_24545,N_23185,N_23449);
nand U24546 (N_24546,N_23861,N_23887);
nor U24547 (N_24547,N_23667,N_23716);
nor U24548 (N_24548,N_23705,N_23430);
nand U24549 (N_24549,N_23282,N_23131);
and U24550 (N_24550,N_23155,N_23897);
xor U24551 (N_24551,N_23375,N_23337);
nand U24552 (N_24552,N_23770,N_23512);
or U24553 (N_24553,N_23645,N_23614);
nand U24554 (N_24554,N_23892,N_23700);
xor U24555 (N_24555,N_23279,N_23058);
xor U24556 (N_24556,N_23698,N_23156);
or U24557 (N_24557,N_23133,N_23064);
or U24558 (N_24558,N_23492,N_23100);
or U24559 (N_24559,N_23996,N_23869);
xor U24560 (N_24560,N_23491,N_23300);
nand U24561 (N_24561,N_23320,N_23254);
or U24562 (N_24562,N_23543,N_23678);
or U24563 (N_24563,N_23580,N_23727);
nand U24564 (N_24564,N_23878,N_23247);
or U24565 (N_24565,N_23172,N_23135);
nand U24566 (N_24566,N_23687,N_23376);
or U24567 (N_24567,N_23937,N_23462);
nor U24568 (N_24568,N_23502,N_23375);
nor U24569 (N_24569,N_23794,N_23795);
xor U24570 (N_24570,N_23263,N_23731);
or U24571 (N_24571,N_23890,N_23075);
nor U24572 (N_24572,N_23161,N_23638);
and U24573 (N_24573,N_23029,N_23325);
nand U24574 (N_24574,N_23750,N_23593);
nand U24575 (N_24575,N_23517,N_23542);
nand U24576 (N_24576,N_23989,N_23120);
xnor U24577 (N_24577,N_23133,N_23322);
nand U24578 (N_24578,N_23271,N_23389);
xor U24579 (N_24579,N_23581,N_23934);
and U24580 (N_24580,N_23085,N_23990);
xor U24581 (N_24581,N_23561,N_23776);
or U24582 (N_24582,N_23251,N_23769);
nand U24583 (N_24583,N_23230,N_23531);
nor U24584 (N_24584,N_23762,N_23725);
nand U24585 (N_24585,N_23323,N_23770);
and U24586 (N_24586,N_23678,N_23923);
nor U24587 (N_24587,N_23896,N_23751);
xor U24588 (N_24588,N_23455,N_23332);
and U24589 (N_24589,N_23550,N_23373);
or U24590 (N_24590,N_23067,N_23037);
xor U24591 (N_24591,N_23278,N_23627);
nor U24592 (N_24592,N_23018,N_23448);
nor U24593 (N_24593,N_23185,N_23196);
nor U24594 (N_24594,N_23934,N_23804);
and U24595 (N_24595,N_23842,N_23682);
nand U24596 (N_24596,N_23886,N_23124);
or U24597 (N_24597,N_23526,N_23257);
or U24598 (N_24598,N_23412,N_23153);
nor U24599 (N_24599,N_23667,N_23594);
nand U24600 (N_24600,N_23122,N_23395);
xnor U24601 (N_24601,N_23096,N_23709);
nor U24602 (N_24602,N_23031,N_23676);
or U24603 (N_24603,N_23751,N_23950);
nor U24604 (N_24604,N_23806,N_23539);
and U24605 (N_24605,N_23289,N_23155);
nor U24606 (N_24606,N_23520,N_23516);
nor U24607 (N_24607,N_23327,N_23973);
xor U24608 (N_24608,N_23865,N_23416);
and U24609 (N_24609,N_23180,N_23571);
or U24610 (N_24610,N_23426,N_23369);
xor U24611 (N_24611,N_23915,N_23048);
nand U24612 (N_24612,N_23098,N_23409);
and U24613 (N_24613,N_23310,N_23299);
or U24614 (N_24614,N_23167,N_23293);
nor U24615 (N_24615,N_23370,N_23181);
and U24616 (N_24616,N_23087,N_23388);
xor U24617 (N_24617,N_23047,N_23804);
nand U24618 (N_24618,N_23154,N_23072);
and U24619 (N_24619,N_23864,N_23386);
nor U24620 (N_24620,N_23908,N_23125);
nand U24621 (N_24621,N_23111,N_23340);
nor U24622 (N_24622,N_23128,N_23034);
nand U24623 (N_24623,N_23861,N_23715);
xnor U24624 (N_24624,N_23406,N_23342);
nand U24625 (N_24625,N_23627,N_23962);
nand U24626 (N_24626,N_23409,N_23683);
and U24627 (N_24627,N_23831,N_23129);
nand U24628 (N_24628,N_23219,N_23393);
or U24629 (N_24629,N_23483,N_23326);
xor U24630 (N_24630,N_23440,N_23316);
nand U24631 (N_24631,N_23646,N_23056);
nor U24632 (N_24632,N_23181,N_23299);
nor U24633 (N_24633,N_23158,N_23568);
xnor U24634 (N_24634,N_23154,N_23444);
nor U24635 (N_24635,N_23303,N_23748);
and U24636 (N_24636,N_23680,N_23657);
nand U24637 (N_24637,N_23403,N_23137);
or U24638 (N_24638,N_23314,N_23870);
xnor U24639 (N_24639,N_23611,N_23546);
xnor U24640 (N_24640,N_23292,N_23472);
xnor U24641 (N_24641,N_23873,N_23425);
or U24642 (N_24642,N_23590,N_23637);
or U24643 (N_24643,N_23311,N_23247);
and U24644 (N_24644,N_23745,N_23999);
or U24645 (N_24645,N_23088,N_23522);
or U24646 (N_24646,N_23299,N_23064);
xnor U24647 (N_24647,N_23505,N_23513);
xnor U24648 (N_24648,N_23442,N_23540);
and U24649 (N_24649,N_23107,N_23302);
and U24650 (N_24650,N_23231,N_23453);
or U24651 (N_24651,N_23338,N_23037);
and U24652 (N_24652,N_23900,N_23558);
or U24653 (N_24653,N_23253,N_23140);
nand U24654 (N_24654,N_23293,N_23779);
xnor U24655 (N_24655,N_23845,N_23562);
nor U24656 (N_24656,N_23294,N_23565);
nand U24657 (N_24657,N_23618,N_23832);
nor U24658 (N_24658,N_23584,N_23301);
or U24659 (N_24659,N_23604,N_23351);
nor U24660 (N_24660,N_23524,N_23828);
nand U24661 (N_24661,N_23684,N_23776);
or U24662 (N_24662,N_23723,N_23762);
or U24663 (N_24663,N_23204,N_23160);
nor U24664 (N_24664,N_23400,N_23317);
xnor U24665 (N_24665,N_23721,N_23373);
xnor U24666 (N_24666,N_23527,N_23476);
or U24667 (N_24667,N_23247,N_23376);
nand U24668 (N_24668,N_23950,N_23099);
and U24669 (N_24669,N_23660,N_23302);
nor U24670 (N_24670,N_23438,N_23155);
nor U24671 (N_24671,N_23861,N_23218);
nor U24672 (N_24672,N_23939,N_23349);
nor U24673 (N_24673,N_23931,N_23418);
nand U24674 (N_24674,N_23898,N_23083);
or U24675 (N_24675,N_23623,N_23265);
nand U24676 (N_24676,N_23091,N_23156);
nor U24677 (N_24677,N_23739,N_23723);
nor U24678 (N_24678,N_23146,N_23614);
xor U24679 (N_24679,N_23163,N_23073);
xnor U24680 (N_24680,N_23970,N_23414);
nor U24681 (N_24681,N_23425,N_23492);
or U24682 (N_24682,N_23946,N_23442);
nand U24683 (N_24683,N_23230,N_23080);
nand U24684 (N_24684,N_23467,N_23685);
nand U24685 (N_24685,N_23426,N_23450);
xnor U24686 (N_24686,N_23663,N_23842);
nand U24687 (N_24687,N_23739,N_23254);
and U24688 (N_24688,N_23379,N_23161);
or U24689 (N_24689,N_23520,N_23362);
or U24690 (N_24690,N_23466,N_23125);
and U24691 (N_24691,N_23817,N_23372);
nor U24692 (N_24692,N_23900,N_23223);
and U24693 (N_24693,N_23478,N_23455);
and U24694 (N_24694,N_23694,N_23579);
or U24695 (N_24695,N_23349,N_23996);
nand U24696 (N_24696,N_23972,N_23131);
nor U24697 (N_24697,N_23551,N_23033);
or U24698 (N_24698,N_23806,N_23393);
xnor U24699 (N_24699,N_23698,N_23301);
nor U24700 (N_24700,N_23040,N_23377);
nor U24701 (N_24701,N_23230,N_23516);
nand U24702 (N_24702,N_23606,N_23949);
xnor U24703 (N_24703,N_23999,N_23722);
nand U24704 (N_24704,N_23289,N_23114);
or U24705 (N_24705,N_23561,N_23005);
xnor U24706 (N_24706,N_23561,N_23137);
and U24707 (N_24707,N_23863,N_23608);
nand U24708 (N_24708,N_23584,N_23279);
nand U24709 (N_24709,N_23581,N_23828);
and U24710 (N_24710,N_23621,N_23960);
nor U24711 (N_24711,N_23342,N_23186);
nor U24712 (N_24712,N_23125,N_23640);
xnor U24713 (N_24713,N_23148,N_23918);
nand U24714 (N_24714,N_23074,N_23442);
xor U24715 (N_24715,N_23486,N_23272);
xnor U24716 (N_24716,N_23056,N_23473);
xor U24717 (N_24717,N_23922,N_23399);
nor U24718 (N_24718,N_23417,N_23553);
and U24719 (N_24719,N_23992,N_23739);
nand U24720 (N_24720,N_23444,N_23845);
xor U24721 (N_24721,N_23992,N_23079);
xor U24722 (N_24722,N_23960,N_23921);
nand U24723 (N_24723,N_23254,N_23230);
xor U24724 (N_24724,N_23523,N_23954);
and U24725 (N_24725,N_23059,N_23830);
or U24726 (N_24726,N_23935,N_23006);
and U24727 (N_24727,N_23676,N_23472);
and U24728 (N_24728,N_23367,N_23284);
or U24729 (N_24729,N_23033,N_23435);
nand U24730 (N_24730,N_23671,N_23059);
nor U24731 (N_24731,N_23044,N_23342);
and U24732 (N_24732,N_23132,N_23742);
xnor U24733 (N_24733,N_23825,N_23201);
or U24734 (N_24734,N_23532,N_23862);
nand U24735 (N_24735,N_23971,N_23419);
and U24736 (N_24736,N_23769,N_23688);
xnor U24737 (N_24737,N_23040,N_23792);
nand U24738 (N_24738,N_23869,N_23136);
nor U24739 (N_24739,N_23164,N_23250);
xor U24740 (N_24740,N_23743,N_23055);
nand U24741 (N_24741,N_23151,N_23658);
nand U24742 (N_24742,N_23596,N_23296);
and U24743 (N_24743,N_23435,N_23452);
and U24744 (N_24744,N_23617,N_23322);
nand U24745 (N_24745,N_23210,N_23280);
and U24746 (N_24746,N_23017,N_23923);
or U24747 (N_24747,N_23601,N_23441);
nand U24748 (N_24748,N_23158,N_23618);
nand U24749 (N_24749,N_23050,N_23437);
xnor U24750 (N_24750,N_23440,N_23354);
nor U24751 (N_24751,N_23649,N_23011);
nand U24752 (N_24752,N_23281,N_23301);
or U24753 (N_24753,N_23438,N_23544);
nor U24754 (N_24754,N_23307,N_23679);
nand U24755 (N_24755,N_23303,N_23011);
and U24756 (N_24756,N_23751,N_23337);
nand U24757 (N_24757,N_23876,N_23299);
xor U24758 (N_24758,N_23797,N_23331);
nor U24759 (N_24759,N_23916,N_23090);
nor U24760 (N_24760,N_23906,N_23838);
nand U24761 (N_24761,N_23009,N_23993);
nand U24762 (N_24762,N_23267,N_23208);
and U24763 (N_24763,N_23360,N_23961);
nor U24764 (N_24764,N_23396,N_23283);
nor U24765 (N_24765,N_23246,N_23227);
nand U24766 (N_24766,N_23993,N_23120);
or U24767 (N_24767,N_23067,N_23196);
nor U24768 (N_24768,N_23922,N_23618);
nand U24769 (N_24769,N_23359,N_23348);
and U24770 (N_24770,N_23850,N_23662);
or U24771 (N_24771,N_23960,N_23171);
or U24772 (N_24772,N_23774,N_23483);
nand U24773 (N_24773,N_23970,N_23376);
nor U24774 (N_24774,N_23406,N_23031);
nor U24775 (N_24775,N_23067,N_23793);
xor U24776 (N_24776,N_23781,N_23416);
or U24777 (N_24777,N_23171,N_23351);
and U24778 (N_24778,N_23362,N_23070);
nand U24779 (N_24779,N_23130,N_23284);
xor U24780 (N_24780,N_23283,N_23022);
or U24781 (N_24781,N_23677,N_23167);
nand U24782 (N_24782,N_23219,N_23842);
and U24783 (N_24783,N_23889,N_23549);
and U24784 (N_24784,N_23336,N_23062);
nor U24785 (N_24785,N_23893,N_23357);
and U24786 (N_24786,N_23115,N_23021);
xor U24787 (N_24787,N_23189,N_23398);
nand U24788 (N_24788,N_23882,N_23426);
nand U24789 (N_24789,N_23595,N_23718);
nor U24790 (N_24790,N_23189,N_23116);
nor U24791 (N_24791,N_23784,N_23027);
and U24792 (N_24792,N_23015,N_23774);
xnor U24793 (N_24793,N_23016,N_23467);
nand U24794 (N_24794,N_23911,N_23775);
nor U24795 (N_24795,N_23374,N_23666);
and U24796 (N_24796,N_23851,N_23079);
nor U24797 (N_24797,N_23930,N_23402);
xnor U24798 (N_24798,N_23331,N_23582);
nand U24799 (N_24799,N_23813,N_23938);
xor U24800 (N_24800,N_23918,N_23233);
and U24801 (N_24801,N_23987,N_23465);
nand U24802 (N_24802,N_23940,N_23839);
nor U24803 (N_24803,N_23722,N_23058);
or U24804 (N_24804,N_23435,N_23486);
or U24805 (N_24805,N_23187,N_23751);
nor U24806 (N_24806,N_23955,N_23491);
or U24807 (N_24807,N_23493,N_23930);
nor U24808 (N_24808,N_23362,N_23884);
or U24809 (N_24809,N_23411,N_23288);
nand U24810 (N_24810,N_23454,N_23363);
xnor U24811 (N_24811,N_23082,N_23261);
nand U24812 (N_24812,N_23421,N_23949);
nor U24813 (N_24813,N_23121,N_23194);
nand U24814 (N_24814,N_23253,N_23987);
xnor U24815 (N_24815,N_23512,N_23967);
xnor U24816 (N_24816,N_23191,N_23743);
xnor U24817 (N_24817,N_23637,N_23762);
or U24818 (N_24818,N_23563,N_23944);
or U24819 (N_24819,N_23940,N_23482);
xnor U24820 (N_24820,N_23922,N_23740);
nor U24821 (N_24821,N_23987,N_23988);
xnor U24822 (N_24822,N_23533,N_23351);
and U24823 (N_24823,N_23258,N_23441);
nor U24824 (N_24824,N_23482,N_23920);
xor U24825 (N_24825,N_23119,N_23858);
xor U24826 (N_24826,N_23979,N_23499);
nand U24827 (N_24827,N_23077,N_23128);
and U24828 (N_24828,N_23505,N_23088);
xnor U24829 (N_24829,N_23810,N_23335);
and U24830 (N_24830,N_23013,N_23054);
xnor U24831 (N_24831,N_23324,N_23607);
xor U24832 (N_24832,N_23239,N_23251);
xnor U24833 (N_24833,N_23565,N_23759);
nand U24834 (N_24834,N_23468,N_23259);
and U24835 (N_24835,N_23129,N_23149);
nand U24836 (N_24836,N_23828,N_23837);
and U24837 (N_24837,N_23866,N_23256);
and U24838 (N_24838,N_23369,N_23116);
and U24839 (N_24839,N_23422,N_23164);
and U24840 (N_24840,N_23908,N_23905);
xor U24841 (N_24841,N_23996,N_23968);
xnor U24842 (N_24842,N_23854,N_23574);
and U24843 (N_24843,N_23487,N_23197);
nor U24844 (N_24844,N_23884,N_23980);
nor U24845 (N_24845,N_23946,N_23665);
and U24846 (N_24846,N_23940,N_23846);
or U24847 (N_24847,N_23504,N_23515);
nand U24848 (N_24848,N_23054,N_23430);
or U24849 (N_24849,N_23235,N_23801);
and U24850 (N_24850,N_23223,N_23543);
and U24851 (N_24851,N_23307,N_23909);
xnor U24852 (N_24852,N_23908,N_23684);
nor U24853 (N_24853,N_23443,N_23738);
nand U24854 (N_24854,N_23246,N_23949);
nor U24855 (N_24855,N_23770,N_23404);
nor U24856 (N_24856,N_23408,N_23967);
nor U24857 (N_24857,N_23463,N_23987);
nor U24858 (N_24858,N_23494,N_23074);
xor U24859 (N_24859,N_23965,N_23064);
and U24860 (N_24860,N_23428,N_23263);
and U24861 (N_24861,N_23419,N_23551);
and U24862 (N_24862,N_23906,N_23385);
nor U24863 (N_24863,N_23863,N_23227);
nand U24864 (N_24864,N_23480,N_23418);
xor U24865 (N_24865,N_23140,N_23700);
or U24866 (N_24866,N_23564,N_23882);
nand U24867 (N_24867,N_23281,N_23395);
nor U24868 (N_24868,N_23464,N_23676);
and U24869 (N_24869,N_23483,N_23024);
xnor U24870 (N_24870,N_23980,N_23454);
xor U24871 (N_24871,N_23621,N_23010);
or U24872 (N_24872,N_23976,N_23347);
or U24873 (N_24873,N_23811,N_23223);
or U24874 (N_24874,N_23180,N_23668);
nor U24875 (N_24875,N_23718,N_23034);
xor U24876 (N_24876,N_23624,N_23384);
or U24877 (N_24877,N_23669,N_23833);
xnor U24878 (N_24878,N_23055,N_23439);
and U24879 (N_24879,N_23809,N_23342);
nor U24880 (N_24880,N_23305,N_23414);
nand U24881 (N_24881,N_23919,N_23224);
xor U24882 (N_24882,N_23119,N_23659);
and U24883 (N_24883,N_23924,N_23993);
and U24884 (N_24884,N_23007,N_23209);
xnor U24885 (N_24885,N_23676,N_23688);
and U24886 (N_24886,N_23899,N_23062);
and U24887 (N_24887,N_23953,N_23060);
nand U24888 (N_24888,N_23236,N_23955);
and U24889 (N_24889,N_23740,N_23076);
or U24890 (N_24890,N_23401,N_23703);
and U24891 (N_24891,N_23326,N_23695);
xnor U24892 (N_24892,N_23354,N_23776);
or U24893 (N_24893,N_23372,N_23950);
or U24894 (N_24894,N_23048,N_23887);
xor U24895 (N_24895,N_23068,N_23855);
nor U24896 (N_24896,N_23097,N_23476);
nand U24897 (N_24897,N_23187,N_23228);
xor U24898 (N_24898,N_23357,N_23372);
nor U24899 (N_24899,N_23222,N_23173);
nand U24900 (N_24900,N_23158,N_23713);
or U24901 (N_24901,N_23720,N_23885);
xor U24902 (N_24902,N_23463,N_23407);
xor U24903 (N_24903,N_23469,N_23048);
xnor U24904 (N_24904,N_23512,N_23805);
nor U24905 (N_24905,N_23496,N_23470);
and U24906 (N_24906,N_23331,N_23510);
nor U24907 (N_24907,N_23944,N_23006);
nand U24908 (N_24908,N_23325,N_23926);
or U24909 (N_24909,N_23939,N_23831);
nor U24910 (N_24910,N_23005,N_23595);
nand U24911 (N_24911,N_23411,N_23968);
and U24912 (N_24912,N_23346,N_23261);
and U24913 (N_24913,N_23156,N_23482);
and U24914 (N_24914,N_23960,N_23548);
nor U24915 (N_24915,N_23182,N_23768);
xor U24916 (N_24916,N_23584,N_23948);
nand U24917 (N_24917,N_23937,N_23959);
nand U24918 (N_24918,N_23643,N_23892);
or U24919 (N_24919,N_23500,N_23952);
nand U24920 (N_24920,N_23318,N_23090);
or U24921 (N_24921,N_23607,N_23219);
nor U24922 (N_24922,N_23107,N_23216);
or U24923 (N_24923,N_23213,N_23647);
xnor U24924 (N_24924,N_23357,N_23197);
xor U24925 (N_24925,N_23174,N_23110);
or U24926 (N_24926,N_23634,N_23038);
and U24927 (N_24927,N_23614,N_23112);
xor U24928 (N_24928,N_23930,N_23322);
nor U24929 (N_24929,N_23849,N_23830);
nor U24930 (N_24930,N_23295,N_23101);
or U24931 (N_24931,N_23686,N_23264);
or U24932 (N_24932,N_23756,N_23583);
and U24933 (N_24933,N_23344,N_23735);
xnor U24934 (N_24934,N_23330,N_23718);
nand U24935 (N_24935,N_23092,N_23046);
nor U24936 (N_24936,N_23758,N_23386);
nand U24937 (N_24937,N_23831,N_23644);
nor U24938 (N_24938,N_23842,N_23432);
or U24939 (N_24939,N_23886,N_23036);
xnor U24940 (N_24940,N_23617,N_23451);
and U24941 (N_24941,N_23854,N_23447);
nor U24942 (N_24942,N_23894,N_23403);
xnor U24943 (N_24943,N_23383,N_23922);
or U24944 (N_24944,N_23689,N_23725);
or U24945 (N_24945,N_23143,N_23776);
nand U24946 (N_24946,N_23390,N_23969);
nand U24947 (N_24947,N_23338,N_23121);
and U24948 (N_24948,N_23763,N_23097);
nor U24949 (N_24949,N_23460,N_23656);
or U24950 (N_24950,N_23832,N_23727);
nor U24951 (N_24951,N_23125,N_23551);
xnor U24952 (N_24952,N_23405,N_23423);
nor U24953 (N_24953,N_23706,N_23978);
nand U24954 (N_24954,N_23690,N_23076);
nor U24955 (N_24955,N_23669,N_23838);
nand U24956 (N_24956,N_23287,N_23805);
and U24957 (N_24957,N_23392,N_23561);
xnor U24958 (N_24958,N_23741,N_23379);
or U24959 (N_24959,N_23595,N_23936);
and U24960 (N_24960,N_23281,N_23377);
xnor U24961 (N_24961,N_23505,N_23512);
nor U24962 (N_24962,N_23806,N_23728);
xor U24963 (N_24963,N_23756,N_23630);
or U24964 (N_24964,N_23035,N_23758);
nand U24965 (N_24965,N_23683,N_23210);
and U24966 (N_24966,N_23268,N_23430);
xnor U24967 (N_24967,N_23440,N_23772);
and U24968 (N_24968,N_23360,N_23119);
and U24969 (N_24969,N_23108,N_23223);
and U24970 (N_24970,N_23754,N_23123);
and U24971 (N_24971,N_23963,N_23023);
nand U24972 (N_24972,N_23946,N_23980);
nor U24973 (N_24973,N_23806,N_23364);
xor U24974 (N_24974,N_23981,N_23625);
nor U24975 (N_24975,N_23851,N_23932);
and U24976 (N_24976,N_23786,N_23774);
nand U24977 (N_24977,N_23290,N_23606);
and U24978 (N_24978,N_23035,N_23294);
or U24979 (N_24979,N_23098,N_23624);
xor U24980 (N_24980,N_23644,N_23816);
nand U24981 (N_24981,N_23278,N_23201);
xnor U24982 (N_24982,N_23129,N_23877);
xor U24983 (N_24983,N_23394,N_23466);
nand U24984 (N_24984,N_23772,N_23775);
nand U24985 (N_24985,N_23433,N_23160);
and U24986 (N_24986,N_23788,N_23684);
nor U24987 (N_24987,N_23155,N_23975);
nand U24988 (N_24988,N_23634,N_23433);
xnor U24989 (N_24989,N_23228,N_23325);
and U24990 (N_24990,N_23955,N_23874);
xnor U24991 (N_24991,N_23392,N_23238);
nand U24992 (N_24992,N_23183,N_23460);
and U24993 (N_24993,N_23320,N_23496);
and U24994 (N_24994,N_23598,N_23693);
or U24995 (N_24995,N_23511,N_23707);
xnor U24996 (N_24996,N_23581,N_23360);
xnor U24997 (N_24997,N_23021,N_23340);
or U24998 (N_24998,N_23670,N_23813);
nor U24999 (N_24999,N_23038,N_23193);
nor U25000 (N_25000,N_24052,N_24427);
nor U25001 (N_25001,N_24182,N_24556);
xor U25002 (N_25002,N_24899,N_24012);
xor U25003 (N_25003,N_24832,N_24907);
and U25004 (N_25004,N_24931,N_24604);
nand U25005 (N_25005,N_24303,N_24664);
nand U25006 (N_25006,N_24080,N_24122);
nor U25007 (N_25007,N_24387,N_24500);
nand U25008 (N_25008,N_24239,N_24475);
nand U25009 (N_25009,N_24641,N_24712);
nand U25010 (N_25010,N_24623,N_24824);
nor U25011 (N_25011,N_24908,N_24237);
nor U25012 (N_25012,N_24968,N_24961);
nand U25013 (N_25013,N_24789,N_24002);
or U25014 (N_25014,N_24777,N_24981);
and U25015 (N_25015,N_24748,N_24661);
xor U25016 (N_25016,N_24693,N_24561);
or U25017 (N_25017,N_24138,N_24628);
xor U25018 (N_25018,N_24807,N_24761);
nor U25019 (N_25019,N_24440,N_24217);
or U25020 (N_25020,N_24861,N_24463);
xor U25021 (N_25021,N_24115,N_24081);
nor U25022 (N_25022,N_24046,N_24865);
xor U25023 (N_25023,N_24862,N_24855);
xor U25024 (N_25024,N_24021,N_24678);
or U25025 (N_25025,N_24649,N_24389);
nor U25026 (N_25026,N_24543,N_24309);
nand U25027 (N_25027,N_24786,N_24158);
or U25028 (N_25028,N_24477,N_24704);
nand U25029 (N_25029,N_24111,N_24375);
nor U25030 (N_25030,N_24569,N_24575);
xnor U25031 (N_25031,N_24214,N_24019);
nand U25032 (N_25032,N_24852,N_24950);
nor U25033 (N_25033,N_24103,N_24467);
nand U25034 (N_25034,N_24296,N_24620);
nor U25035 (N_25035,N_24334,N_24383);
nor U25036 (N_25036,N_24951,N_24105);
xnor U25037 (N_25037,N_24498,N_24281);
and U25038 (N_25038,N_24403,N_24711);
and U25039 (N_25039,N_24574,N_24354);
xor U25040 (N_25040,N_24897,N_24545);
and U25041 (N_25041,N_24532,N_24340);
and U25042 (N_25042,N_24109,N_24117);
xor U25043 (N_25043,N_24054,N_24790);
nand U25044 (N_25044,N_24558,N_24534);
and U25045 (N_25045,N_24251,N_24257);
xnor U25046 (N_25046,N_24429,N_24895);
nor U25047 (N_25047,N_24576,N_24982);
and U25048 (N_25048,N_24420,N_24579);
and U25049 (N_25049,N_24555,N_24888);
nand U25050 (N_25050,N_24552,N_24962);
and U25051 (N_25051,N_24922,N_24402);
or U25052 (N_25052,N_24470,N_24767);
xor U25053 (N_25053,N_24095,N_24644);
or U25054 (N_25054,N_24487,N_24528);
nor U25055 (N_25055,N_24921,N_24504);
xnor U25056 (N_25056,N_24956,N_24444);
nor U25057 (N_25057,N_24206,N_24356);
and U25058 (N_25058,N_24248,N_24010);
and U25059 (N_25059,N_24811,N_24934);
or U25060 (N_25060,N_24608,N_24377);
nor U25061 (N_25061,N_24850,N_24039);
nand U25062 (N_25062,N_24030,N_24026);
nand U25063 (N_25063,N_24565,N_24265);
xor U25064 (N_25064,N_24005,N_24755);
xnor U25065 (N_25065,N_24652,N_24568);
and U25066 (N_25066,N_24129,N_24462);
and U25067 (N_25067,N_24457,N_24174);
xnor U25068 (N_25068,N_24696,N_24107);
xnor U25069 (N_25069,N_24802,N_24959);
and U25070 (N_25070,N_24668,N_24379);
xnor U25071 (N_25071,N_24053,N_24726);
xor U25072 (N_25072,N_24345,N_24090);
or U25073 (N_25073,N_24706,N_24526);
and U25074 (N_25074,N_24267,N_24011);
xnor U25075 (N_25075,N_24683,N_24827);
nor U25076 (N_25076,N_24353,N_24796);
xor U25077 (N_25077,N_24488,N_24378);
nand U25078 (N_25078,N_24323,N_24141);
and U25079 (N_25079,N_24300,N_24215);
or U25080 (N_25080,N_24041,N_24537);
nor U25081 (N_25081,N_24876,N_24218);
nor U25082 (N_25082,N_24236,N_24370);
and U25083 (N_25083,N_24549,N_24229);
or U25084 (N_25084,N_24113,N_24671);
nor U25085 (N_25085,N_24814,N_24362);
or U25086 (N_25086,N_24737,N_24978);
or U25087 (N_25087,N_24770,N_24875);
xor U25088 (N_25088,N_24910,N_24725);
and U25089 (N_25089,N_24635,N_24909);
xor U25090 (N_25090,N_24104,N_24896);
xor U25091 (N_25091,N_24042,N_24878);
and U25092 (N_25092,N_24466,N_24607);
nor U25093 (N_25093,N_24305,N_24879);
or U25094 (N_25094,N_24242,N_24455);
xnor U25095 (N_25095,N_24792,N_24175);
or U25096 (N_25096,N_24201,N_24829);
nor U25097 (N_25097,N_24634,N_24401);
and U25098 (N_25098,N_24658,N_24369);
nand U25099 (N_25099,N_24847,N_24540);
nor U25100 (N_25100,N_24837,N_24139);
and U25101 (N_25101,N_24844,N_24009);
nor U25102 (N_25102,N_24840,N_24191);
nor U25103 (N_25103,N_24581,N_24295);
nand U25104 (N_25104,N_24784,N_24224);
xor U25105 (N_25105,N_24744,N_24253);
xor U25106 (N_25106,N_24904,N_24348);
and U25107 (N_25107,N_24318,N_24078);
xnor U25108 (N_25108,N_24096,N_24461);
nand U25109 (N_25109,N_24038,N_24456);
xor U25110 (N_25110,N_24361,N_24062);
and U25111 (N_25111,N_24343,N_24233);
and U25112 (N_25112,N_24559,N_24621);
xor U25113 (N_25113,N_24400,N_24991);
or U25114 (N_25114,N_24503,N_24302);
xor U25115 (N_25115,N_24252,N_24014);
nor U25116 (N_25116,N_24716,N_24371);
nand U25117 (N_25117,N_24849,N_24600);
nor U25118 (N_25118,N_24178,N_24690);
nand U25119 (N_25119,N_24100,N_24605);
nand U25120 (N_25120,N_24226,N_24294);
or U25121 (N_25121,N_24204,N_24816);
and U25122 (N_25122,N_24405,N_24809);
nor U25123 (N_25123,N_24173,N_24614);
or U25124 (N_25124,N_24842,N_24980);
nand U25125 (N_25125,N_24029,N_24593);
nand U25126 (N_25126,N_24927,N_24612);
or U25127 (N_25127,N_24374,N_24666);
xnor U25128 (N_25128,N_24828,N_24519);
or U25129 (N_25129,N_24358,N_24274);
xnor U25130 (N_25130,N_24602,N_24501);
nand U25131 (N_25131,N_24881,N_24264);
or U25132 (N_25132,N_24718,N_24486);
nand U25133 (N_25133,N_24198,N_24795);
xnor U25134 (N_25134,N_24164,N_24990);
and U25135 (N_25135,N_24151,N_24376);
xor U25136 (N_25136,N_24426,N_24815);
xor U25137 (N_25137,N_24186,N_24819);
nand U25138 (N_25138,N_24752,N_24924);
nand U25139 (N_25139,N_24863,N_24413);
nand U25140 (N_25140,N_24459,N_24538);
or U25141 (N_25141,N_24817,N_24774);
nand U25142 (N_25142,N_24258,N_24428);
or U25143 (N_25143,N_24473,N_24651);
xor U25144 (N_25144,N_24131,N_24072);
nor U25145 (N_25145,N_24476,N_24312);
xnor U25146 (N_25146,N_24443,N_24489);
xnor U25147 (N_25147,N_24411,N_24722);
or U25148 (N_25148,N_24800,N_24525);
and U25149 (N_25149,N_24342,N_24775);
and U25150 (N_25150,N_24025,N_24435);
or U25151 (N_25151,N_24393,N_24065);
nand U25152 (N_25152,N_24179,N_24381);
xnor U25153 (N_25153,N_24518,N_24143);
nor U25154 (N_25154,N_24165,N_24063);
nand U25155 (N_25155,N_24419,N_24527);
and U25156 (N_25156,N_24825,N_24149);
nand U25157 (N_25157,N_24893,N_24724);
or U25158 (N_25158,N_24040,N_24930);
nor U25159 (N_25159,N_24629,N_24000);
nand U25160 (N_25160,N_24169,N_24273);
nor U25161 (N_25161,N_24118,N_24860);
and U25162 (N_25162,N_24184,N_24536);
and U25163 (N_25163,N_24662,N_24275);
nand U25164 (N_25164,N_24452,N_24187);
or U25165 (N_25165,N_24570,N_24917);
or U25166 (N_25166,N_24957,N_24380);
xor U25167 (N_25167,N_24060,N_24099);
or U25168 (N_25168,N_24485,N_24915);
and U25169 (N_25169,N_24315,N_24680);
nand U25170 (N_25170,N_24263,N_24617);
nor U25171 (N_25171,N_24952,N_24747);
and U25172 (N_25172,N_24056,N_24886);
and U25173 (N_25173,N_24566,N_24513);
or U25174 (N_25174,N_24177,N_24373);
nor U25175 (N_25175,N_24967,N_24089);
nand U25176 (N_25176,N_24939,N_24554);
xor U25177 (N_25177,N_24582,N_24830);
nor U25178 (N_25178,N_24900,N_24512);
or U25179 (N_25179,N_24076,N_24707);
nor U25180 (N_25180,N_24431,N_24660);
xor U25181 (N_25181,N_24781,N_24140);
and U25182 (N_25182,N_24254,N_24762);
nor U25183 (N_25183,N_24928,N_24533);
nor U25184 (N_25184,N_24687,N_24208);
and U25185 (N_25185,N_24866,N_24289);
and U25186 (N_25186,N_24097,N_24497);
xor U25187 (N_25187,N_24667,N_24479);
nor U25188 (N_25188,N_24529,N_24654);
or U25189 (N_25189,N_24337,N_24517);
or U25190 (N_25190,N_24196,N_24839);
and U25191 (N_25191,N_24885,N_24259);
nand U25192 (N_25192,N_24494,N_24992);
nand U25193 (N_25193,N_24384,N_24856);
nor U25194 (N_25194,N_24130,N_24396);
or U25195 (N_25195,N_24898,N_24567);
nand U25196 (N_25196,N_24560,N_24889);
xnor U25197 (N_25197,N_24496,N_24086);
and U25198 (N_25198,N_24262,N_24495);
or U25199 (N_25199,N_24547,N_24066);
nor U25200 (N_25200,N_24162,N_24601);
xor U25201 (N_25201,N_24050,N_24764);
nor U25202 (N_25202,N_24047,N_24622);
xnor U25203 (N_25203,N_24867,N_24048);
xor U25204 (N_25204,N_24493,N_24616);
nand U25205 (N_25205,N_24759,N_24721);
xor U25206 (N_25206,N_24794,N_24720);
nor U25207 (N_25207,N_24698,N_24004);
nand U25208 (N_25208,N_24145,N_24133);
nand U25209 (N_25209,N_24768,N_24799);
and U25210 (N_25210,N_24787,N_24286);
or U25211 (N_25211,N_24003,N_24749);
nand U25212 (N_25212,N_24892,N_24619);
xor U25213 (N_25213,N_24914,N_24449);
and U25214 (N_25214,N_24806,N_24584);
and U25215 (N_25215,N_24542,N_24675);
xor U25216 (N_25216,N_24194,N_24701);
or U25217 (N_25217,N_24719,N_24125);
or U25218 (N_25218,N_24697,N_24299);
nand U25219 (N_25219,N_24677,N_24433);
and U25220 (N_25220,N_24778,N_24942);
xor U25221 (N_25221,N_24682,N_24171);
or U25222 (N_25222,N_24672,N_24448);
nor U25223 (N_25223,N_24170,N_24857);
and U25224 (N_25224,N_24211,N_24756);
nor U25225 (N_25225,N_24936,N_24727);
nand U25226 (N_25226,N_24395,N_24359);
nor U25227 (N_25227,N_24327,N_24142);
or U25228 (N_25228,N_24195,N_24835);
nor U25229 (N_25229,N_24788,N_24001);
nand U25230 (N_25230,N_24723,N_24058);
and U25231 (N_25231,N_24769,N_24679);
and U25232 (N_25232,N_24276,N_24188);
xnor U25233 (N_25233,N_24890,N_24713);
and U25234 (N_25234,N_24838,N_24779);
nor U25235 (N_25235,N_24851,N_24087);
and U25236 (N_25236,N_24606,N_24051);
and U25237 (N_25237,N_24074,N_24160);
nor U25238 (N_25238,N_24098,N_24699);
xnor U25239 (N_25239,N_24508,N_24548);
xor U25240 (N_25240,N_24321,N_24282);
xnor U25241 (N_25241,N_24422,N_24156);
or U25242 (N_25242,N_24804,N_24880);
nand U25243 (N_25243,N_24938,N_24415);
xnor U25244 (N_25244,N_24231,N_24708);
nor U25245 (N_25245,N_24669,N_24271);
xnor U25246 (N_25246,N_24083,N_24646);
nand U25247 (N_25247,N_24988,N_24243);
xnor U25248 (N_25248,N_24114,N_24335);
or U25249 (N_25249,N_24618,N_24925);
or U25250 (N_25250,N_24953,N_24571);
or U25251 (N_25251,N_24960,N_24193);
nor U25252 (N_25252,N_24831,N_24958);
nor U25253 (N_25253,N_24505,N_24238);
or U25254 (N_25254,N_24249,N_24205);
nand U25255 (N_25255,N_24624,N_24260);
nand U25256 (N_25256,N_24688,N_24673);
and U25257 (N_25257,N_24546,N_24995);
and U25258 (N_25258,N_24833,N_24034);
xnor U25259 (N_25259,N_24681,N_24771);
xor U25260 (N_25260,N_24210,N_24776);
nor U25261 (N_25261,N_24157,N_24611);
xor U25262 (N_25262,N_24805,N_24595);
nand U25263 (N_25263,N_24514,N_24288);
xor U25264 (N_25264,N_24082,N_24821);
or U25265 (N_25265,N_24094,N_24705);
and U25266 (N_25266,N_24324,N_24279);
nor U25267 (N_25267,N_24367,N_24750);
xor U25268 (N_25268,N_24557,N_24963);
or U25269 (N_25269,N_24167,N_24241);
and U25270 (N_25270,N_24023,N_24933);
nor U25271 (N_25271,N_24044,N_24481);
nand U25272 (N_25272,N_24108,N_24630);
nor U25273 (N_25273,N_24562,N_24906);
nand U25274 (N_25274,N_24740,N_24948);
and U25275 (N_25275,N_24310,N_24172);
and U25276 (N_25276,N_24333,N_24941);
nor U25277 (N_25277,N_24071,N_24027);
xor U25278 (N_25278,N_24035,N_24710);
xnor U25279 (N_25279,N_24385,N_24594);
nor U25280 (N_25280,N_24269,N_24181);
nor U25281 (N_25281,N_24454,N_24663);
nand U25282 (N_25282,N_24753,N_24643);
nor U25283 (N_25283,N_24355,N_24159);
or U25284 (N_25284,N_24969,N_24685);
nand U25285 (N_25285,N_24563,N_24996);
or U25286 (N_25286,N_24136,N_24372);
and U25287 (N_25287,N_24330,N_24882);
nor U25288 (N_25288,N_24067,N_24544);
and U25289 (N_25289,N_24993,N_24998);
nor U25290 (N_25290,N_24073,N_24316);
or U25291 (N_25291,N_24813,N_24013);
and U25292 (N_25292,N_24392,N_24591);
and U25293 (N_25293,N_24209,N_24222);
nor U25294 (N_25294,N_24820,N_24313);
xnor U25295 (N_25295,N_24092,N_24541);
and U25296 (N_25296,N_24293,N_24306);
and U25297 (N_25297,N_24287,N_24460);
or U25298 (N_25298,N_24192,N_24365);
nand U25299 (N_25299,N_24059,N_24070);
nor U25300 (N_25300,N_24798,N_24144);
or U25301 (N_25301,N_24609,N_24940);
and U25302 (N_25302,N_24451,N_24911);
nand U25303 (N_25303,N_24923,N_24414);
and U25304 (N_25304,N_24057,N_24797);
or U25305 (N_25305,N_24135,N_24423);
xor U25306 (N_25306,N_24386,N_24166);
and U25307 (N_25307,N_24255,N_24219);
or U25308 (N_25308,N_24979,N_24368);
nor U25309 (N_25309,N_24883,N_24007);
nand U25310 (N_25310,N_24946,N_24743);
or U25311 (N_25311,N_24736,N_24632);
nor U25312 (N_25312,N_24588,N_24290);
or U25313 (N_25313,N_24822,N_24535);
nor U25314 (N_25314,N_24846,N_24351);
and U25315 (N_25315,N_24434,N_24091);
nor U25316 (N_25316,N_24745,N_24746);
nand U25317 (N_25317,N_24116,N_24766);
nor U25318 (N_25318,N_24965,N_24596);
and U25319 (N_25319,N_24366,N_24382);
or U25320 (N_25320,N_24642,N_24410);
xor U25321 (N_25321,N_24702,N_24292);
and U25322 (N_25322,N_24971,N_24406);
or U25323 (N_25323,N_24877,N_24695);
xor U25324 (N_25324,N_24929,N_24152);
and U25325 (N_25325,N_24949,N_24905);
xnor U25326 (N_25326,N_24585,N_24437);
and U25327 (N_25327,N_24627,N_24036);
nor U25328 (N_25328,N_24424,N_24580);
xnor U25329 (N_25329,N_24586,N_24947);
xnor U25330 (N_25330,N_24553,N_24870);
nor U25331 (N_25331,N_24970,N_24008);
and U25332 (N_25332,N_24329,N_24220);
and U25333 (N_25333,N_24391,N_24572);
xor U25334 (N_25334,N_24350,N_24207);
and U25335 (N_25335,N_24101,N_24185);
nor U25336 (N_25336,N_24515,N_24810);
nor U25337 (N_25337,N_24626,N_24425);
and U25338 (N_25338,N_24499,N_24684);
nor U25339 (N_25339,N_24168,N_24730);
xnor U25340 (N_25340,N_24069,N_24943);
or U25341 (N_25341,N_24686,N_24738);
and U25342 (N_25342,N_24733,N_24509);
nor U25343 (N_25343,N_24016,N_24578);
or U25344 (N_25344,N_24480,N_24613);
nand U25345 (N_25345,N_24871,N_24232);
nand U25346 (N_25346,N_24598,N_24338);
and U25347 (N_25347,N_24216,N_24785);
or U25348 (N_25348,N_24818,N_24079);
nor U25349 (N_25349,N_24438,N_24700);
xor U25350 (N_25350,N_24028,N_24689);
or U25351 (N_25351,N_24364,N_24659);
nand U25352 (N_25352,N_24551,N_24439);
nor U25353 (N_25353,N_24280,N_24592);
xnor U25354 (N_25354,N_24577,N_24146);
or U25355 (N_25355,N_24319,N_24307);
and U25356 (N_25356,N_24045,N_24180);
nand U25357 (N_25357,N_24247,N_24843);
or U25358 (N_25358,N_24085,N_24388);
or U25359 (N_25359,N_24447,N_24587);
or U25360 (N_25360,N_24735,N_24913);
nand U25361 (N_25361,N_24037,N_24997);
xnor U25362 (N_25362,N_24801,N_24603);
and U25363 (N_25363,N_24360,N_24854);
and U25364 (N_25364,N_24270,N_24064);
xnor U25365 (N_25365,N_24638,N_24751);
xor U25366 (N_25366,N_24320,N_24148);
xnor U25367 (N_25367,N_24277,N_24521);
xor U25368 (N_25368,N_24783,N_24347);
nor U25369 (N_25369,N_24446,N_24502);
nor U25370 (N_25370,N_24346,N_24715);
xnor U25371 (N_25371,N_24154,N_24903);
nand U25372 (N_25372,N_24484,N_24197);
nand U25373 (N_25373,N_24363,N_24902);
and U25374 (N_25374,N_24161,N_24703);
and U25375 (N_25375,N_24511,N_24212);
or U25376 (N_25376,N_24823,N_24119);
nor U25377 (N_25377,N_24407,N_24339);
or U25378 (N_25378,N_24676,N_24006);
or U25379 (N_25379,N_24155,N_24328);
nor U25380 (N_25380,N_24412,N_24665);
and U25381 (N_25381,N_24564,N_24049);
or U25382 (N_25382,N_24966,N_24803);
nor U25383 (N_25383,N_24757,N_24937);
nand U25384 (N_25384,N_24227,N_24120);
or U25385 (N_25385,N_24134,N_24317);
xor U25386 (N_25386,N_24308,N_24015);
or U25387 (N_25387,N_24017,N_24834);
xor U25388 (N_25388,N_24772,N_24127);
and U25389 (N_25389,N_24311,N_24887);
and U25390 (N_25390,N_24826,N_24124);
xor U25391 (N_25391,N_24213,N_24977);
or U25392 (N_25392,N_24845,N_24973);
xor U25393 (N_25393,N_24599,N_24352);
and U25394 (N_25394,N_24331,N_24782);
nand U25395 (N_25395,N_24341,N_24478);
nand U25396 (N_25396,N_24482,N_24859);
nor U25397 (N_25397,N_24655,N_24297);
and U25398 (N_25398,N_24884,N_24935);
or U25399 (N_25399,N_24901,N_24983);
xnor U25400 (N_25400,N_24986,N_24397);
and U25401 (N_25401,N_24147,N_24490);
xnor U25402 (N_25402,N_24245,N_24674);
xnor U25403 (N_25403,N_24984,N_24873);
nor U25404 (N_25404,N_24024,N_24869);
nand U25405 (N_25405,N_24176,N_24336);
xor U25406 (N_25406,N_24625,N_24399);
or U25407 (N_25407,N_24106,N_24709);
or U25408 (N_25408,N_24610,N_24221);
xnor U25409 (N_25409,N_24657,N_24868);
and U25410 (N_25410,N_24717,N_24202);
and U25411 (N_25411,N_24033,N_24597);
xnor U25412 (N_25412,N_24442,N_24075);
xnor U25413 (N_25413,N_24483,N_24872);
nor U25414 (N_25414,N_24550,N_24266);
or U25415 (N_25415,N_24235,N_24110);
nand U25416 (N_25416,N_24228,N_24272);
or U25417 (N_25417,N_24421,N_24972);
nand U25418 (N_25418,N_24523,N_24453);
or U25419 (N_25419,N_24203,N_24123);
nor U25420 (N_25420,N_24780,N_24301);
and U25421 (N_25421,N_24430,N_24637);
nand U25422 (N_25422,N_24326,N_24077);
or U25423 (N_25423,N_24150,N_24763);
and U25424 (N_25424,N_24061,N_24506);
or U25425 (N_25425,N_24836,N_24390);
nor U25426 (N_25426,N_24731,N_24999);
xnor U25427 (N_25427,N_24223,N_24640);
or U25428 (N_25428,N_24692,N_24043);
and U25429 (N_25429,N_24357,N_24648);
and U25430 (N_25430,N_24298,N_24332);
nand U25431 (N_25431,N_24153,N_24464);
xor U25432 (N_25432,N_24520,N_24694);
xnor U25433 (N_25433,N_24760,N_24729);
nor U25434 (N_25434,N_24754,N_24994);
xnor U25435 (N_25435,N_24653,N_24284);
nor U25436 (N_25436,N_24132,N_24032);
or U25437 (N_25437,N_24250,N_24583);
nor U25438 (N_25438,N_24022,N_24573);
xnor U25439 (N_25439,N_24912,N_24864);
nor U25440 (N_25440,N_24732,N_24791);
nand U25441 (N_25441,N_24304,N_24920);
nor U25442 (N_25442,N_24808,N_24615);
xor U25443 (N_25443,N_24163,N_24137);
xor U25444 (N_25444,N_24975,N_24670);
xnor U25445 (N_25445,N_24894,N_24773);
and U25446 (N_25446,N_24278,N_24398);
nand U25447 (N_25447,N_24647,N_24200);
nand U25448 (N_25448,N_24758,N_24985);
nor U25449 (N_25449,N_24691,N_24516);
xor U25450 (N_25450,N_24018,N_24246);
nor U25451 (N_25451,N_24468,N_24944);
nand U25452 (N_25452,N_24987,N_24084);
and U25453 (N_25453,N_24055,N_24812);
and U25454 (N_25454,N_24793,N_24492);
or U25455 (N_25455,N_24349,N_24183);
or U25456 (N_25456,N_24853,N_24408);
and U25457 (N_25457,N_24955,N_24469);
nor U25458 (N_25458,N_24244,N_24126);
and U25459 (N_25459,N_24450,N_24068);
or U25460 (N_25460,N_24728,N_24394);
xnor U25461 (N_25461,N_24436,N_24954);
nor U25462 (N_25462,N_24261,N_24841);
xnor U25463 (N_25463,N_24765,N_24848);
nand U25464 (N_25464,N_24121,N_24418);
or U25465 (N_25465,N_24507,N_24441);
xor U25466 (N_25466,N_24639,N_24531);
nand U25467 (N_25467,N_24256,N_24633);
nand U25468 (N_25468,N_24020,N_24291);
xor U25469 (N_25469,N_24874,N_24471);
and U25470 (N_25470,N_24645,N_24522);
nor U25471 (N_25471,N_24976,N_24472);
xor U25472 (N_25472,N_24636,N_24240);
xnor U25473 (N_25473,N_24268,N_24590);
xnor U25474 (N_25474,N_24325,N_24714);
xnor U25475 (N_25475,N_24741,N_24589);
xnor U25476 (N_25476,N_24088,N_24524);
xnor U25477 (N_25477,N_24432,N_24491);
or U25478 (N_25478,N_24234,N_24650);
and U25479 (N_25479,N_24190,N_24409);
nor U25480 (N_25480,N_24112,N_24404);
nand U25481 (N_25481,N_24474,N_24656);
or U25482 (N_25482,N_24742,N_24458);
nor U25483 (N_25483,N_24932,N_24093);
nand U25484 (N_25484,N_24891,N_24989);
or U25485 (N_25485,N_24945,N_24919);
xnor U25486 (N_25486,N_24964,N_24285);
xor U25487 (N_25487,N_24631,N_24199);
nand U25488 (N_25488,N_24230,N_24916);
nand U25489 (N_25489,N_24225,N_24417);
and U25490 (N_25490,N_24283,N_24539);
or U25491 (N_25491,N_24416,N_24530);
xnor U25492 (N_25492,N_24322,N_24510);
nor U25493 (N_25493,N_24926,N_24445);
xor U25494 (N_25494,N_24314,N_24189);
xnor U25495 (N_25495,N_24344,N_24974);
nor U25496 (N_25496,N_24102,N_24734);
or U25497 (N_25497,N_24031,N_24465);
and U25498 (N_25498,N_24858,N_24918);
xnor U25499 (N_25499,N_24739,N_24128);
nand U25500 (N_25500,N_24823,N_24077);
or U25501 (N_25501,N_24090,N_24790);
and U25502 (N_25502,N_24250,N_24269);
nand U25503 (N_25503,N_24396,N_24138);
and U25504 (N_25504,N_24149,N_24302);
nand U25505 (N_25505,N_24384,N_24862);
xnor U25506 (N_25506,N_24937,N_24841);
or U25507 (N_25507,N_24763,N_24157);
and U25508 (N_25508,N_24859,N_24164);
nand U25509 (N_25509,N_24779,N_24009);
nor U25510 (N_25510,N_24684,N_24375);
nand U25511 (N_25511,N_24823,N_24032);
or U25512 (N_25512,N_24514,N_24572);
or U25513 (N_25513,N_24048,N_24915);
nand U25514 (N_25514,N_24626,N_24548);
nand U25515 (N_25515,N_24611,N_24805);
nor U25516 (N_25516,N_24689,N_24446);
or U25517 (N_25517,N_24807,N_24359);
nor U25518 (N_25518,N_24498,N_24698);
nand U25519 (N_25519,N_24102,N_24305);
nor U25520 (N_25520,N_24316,N_24499);
nor U25521 (N_25521,N_24448,N_24089);
nor U25522 (N_25522,N_24142,N_24413);
or U25523 (N_25523,N_24532,N_24824);
or U25524 (N_25524,N_24688,N_24297);
xor U25525 (N_25525,N_24381,N_24346);
and U25526 (N_25526,N_24187,N_24298);
or U25527 (N_25527,N_24133,N_24182);
or U25528 (N_25528,N_24304,N_24576);
nor U25529 (N_25529,N_24744,N_24718);
nor U25530 (N_25530,N_24029,N_24614);
and U25531 (N_25531,N_24548,N_24316);
or U25532 (N_25532,N_24588,N_24223);
nand U25533 (N_25533,N_24266,N_24479);
xor U25534 (N_25534,N_24709,N_24736);
or U25535 (N_25535,N_24673,N_24041);
nand U25536 (N_25536,N_24949,N_24941);
or U25537 (N_25537,N_24855,N_24533);
or U25538 (N_25538,N_24434,N_24277);
and U25539 (N_25539,N_24781,N_24065);
nor U25540 (N_25540,N_24467,N_24614);
and U25541 (N_25541,N_24200,N_24360);
nand U25542 (N_25542,N_24594,N_24398);
xnor U25543 (N_25543,N_24391,N_24842);
xnor U25544 (N_25544,N_24988,N_24662);
and U25545 (N_25545,N_24836,N_24425);
and U25546 (N_25546,N_24742,N_24807);
or U25547 (N_25547,N_24007,N_24245);
nor U25548 (N_25548,N_24938,N_24263);
nor U25549 (N_25549,N_24691,N_24074);
and U25550 (N_25550,N_24838,N_24148);
nand U25551 (N_25551,N_24906,N_24799);
or U25552 (N_25552,N_24918,N_24495);
and U25553 (N_25553,N_24952,N_24662);
nor U25554 (N_25554,N_24915,N_24770);
xor U25555 (N_25555,N_24693,N_24995);
or U25556 (N_25556,N_24851,N_24581);
and U25557 (N_25557,N_24366,N_24818);
nand U25558 (N_25558,N_24389,N_24784);
nand U25559 (N_25559,N_24996,N_24205);
or U25560 (N_25560,N_24535,N_24931);
or U25561 (N_25561,N_24119,N_24446);
and U25562 (N_25562,N_24428,N_24257);
nor U25563 (N_25563,N_24691,N_24947);
and U25564 (N_25564,N_24651,N_24622);
or U25565 (N_25565,N_24033,N_24667);
or U25566 (N_25566,N_24602,N_24902);
nor U25567 (N_25567,N_24562,N_24677);
nand U25568 (N_25568,N_24033,N_24196);
nor U25569 (N_25569,N_24921,N_24758);
nand U25570 (N_25570,N_24291,N_24225);
and U25571 (N_25571,N_24987,N_24371);
xnor U25572 (N_25572,N_24299,N_24698);
or U25573 (N_25573,N_24984,N_24222);
or U25574 (N_25574,N_24317,N_24398);
and U25575 (N_25575,N_24875,N_24029);
nor U25576 (N_25576,N_24616,N_24625);
nor U25577 (N_25577,N_24955,N_24380);
and U25578 (N_25578,N_24364,N_24699);
and U25579 (N_25579,N_24673,N_24018);
nand U25580 (N_25580,N_24160,N_24698);
or U25581 (N_25581,N_24544,N_24302);
or U25582 (N_25582,N_24715,N_24064);
nor U25583 (N_25583,N_24128,N_24191);
xnor U25584 (N_25584,N_24968,N_24545);
nor U25585 (N_25585,N_24519,N_24259);
or U25586 (N_25586,N_24895,N_24870);
and U25587 (N_25587,N_24905,N_24175);
or U25588 (N_25588,N_24542,N_24872);
nand U25589 (N_25589,N_24148,N_24195);
nor U25590 (N_25590,N_24283,N_24530);
nor U25591 (N_25591,N_24693,N_24459);
nand U25592 (N_25592,N_24004,N_24990);
or U25593 (N_25593,N_24782,N_24585);
nand U25594 (N_25594,N_24912,N_24009);
xnor U25595 (N_25595,N_24248,N_24489);
nand U25596 (N_25596,N_24426,N_24286);
xnor U25597 (N_25597,N_24367,N_24704);
nand U25598 (N_25598,N_24100,N_24420);
and U25599 (N_25599,N_24650,N_24699);
and U25600 (N_25600,N_24843,N_24537);
or U25601 (N_25601,N_24251,N_24669);
or U25602 (N_25602,N_24096,N_24113);
nand U25603 (N_25603,N_24112,N_24026);
nor U25604 (N_25604,N_24119,N_24156);
and U25605 (N_25605,N_24704,N_24423);
or U25606 (N_25606,N_24234,N_24631);
and U25607 (N_25607,N_24866,N_24905);
xnor U25608 (N_25608,N_24424,N_24862);
or U25609 (N_25609,N_24298,N_24929);
nand U25610 (N_25610,N_24638,N_24870);
or U25611 (N_25611,N_24566,N_24335);
and U25612 (N_25612,N_24039,N_24766);
nand U25613 (N_25613,N_24427,N_24638);
or U25614 (N_25614,N_24036,N_24643);
and U25615 (N_25615,N_24493,N_24411);
xnor U25616 (N_25616,N_24341,N_24360);
xor U25617 (N_25617,N_24652,N_24686);
or U25618 (N_25618,N_24840,N_24458);
nor U25619 (N_25619,N_24824,N_24752);
and U25620 (N_25620,N_24627,N_24709);
xor U25621 (N_25621,N_24285,N_24638);
nand U25622 (N_25622,N_24327,N_24891);
xor U25623 (N_25623,N_24248,N_24358);
xor U25624 (N_25624,N_24721,N_24745);
nand U25625 (N_25625,N_24449,N_24452);
and U25626 (N_25626,N_24559,N_24022);
or U25627 (N_25627,N_24047,N_24045);
nand U25628 (N_25628,N_24025,N_24288);
nor U25629 (N_25629,N_24940,N_24932);
nand U25630 (N_25630,N_24238,N_24167);
and U25631 (N_25631,N_24081,N_24579);
nand U25632 (N_25632,N_24478,N_24363);
nand U25633 (N_25633,N_24776,N_24704);
or U25634 (N_25634,N_24187,N_24131);
and U25635 (N_25635,N_24436,N_24707);
nand U25636 (N_25636,N_24816,N_24135);
nor U25637 (N_25637,N_24628,N_24070);
xor U25638 (N_25638,N_24436,N_24406);
and U25639 (N_25639,N_24713,N_24078);
xnor U25640 (N_25640,N_24788,N_24586);
nand U25641 (N_25641,N_24676,N_24686);
nor U25642 (N_25642,N_24875,N_24151);
and U25643 (N_25643,N_24904,N_24139);
and U25644 (N_25644,N_24925,N_24833);
nor U25645 (N_25645,N_24211,N_24384);
nand U25646 (N_25646,N_24331,N_24563);
xnor U25647 (N_25647,N_24496,N_24876);
xnor U25648 (N_25648,N_24688,N_24228);
and U25649 (N_25649,N_24489,N_24632);
nor U25650 (N_25650,N_24035,N_24241);
nand U25651 (N_25651,N_24524,N_24754);
or U25652 (N_25652,N_24220,N_24237);
nand U25653 (N_25653,N_24615,N_24064);
xnor U25654 (N_25654,N_24843,N_24086);
or U25655 (N_25655,N_24984,N_24116);
or U25656 (N_25656,N_24973,N_24963);
nor U25657 (N_25657,N_24208,N_24298);
or U25658 (N_25658,N_24307,N_24293);
and U25659 (N_25659,N_24029,N_24598);
nand U25660 (N_25660,N_24001,N_24366);
xnor U25661 (N_25661,N_24018,N_24185);
nor U25662 (N_25662,N_24474,N_24136);
nand U25663 (N_25663,N_24375,N_24269);
and U25664 (N_25664,N_24682,N_24529);
xor U25665 (N_25665,N_24430,N_24446);
nand U25666 (N_25666,N_24514,N_24891);
nand U25667 (N_25667,N_24331,N_24854);
and U25668 (N_25668,N_24374,N_24439);
nand U25669 (N_25669,N_24973,N_24561);
nand U25670 (N_25670,N_24489,N_24111);
and U25671 (N_25671,N_24967,N_24579);
nor U25672 (N_25672,N_24754,N_24165);
nor U25673 (N_25673,N_24145,N_24371);
nor U25674 (N_25674,N_24205,N_24892);
nand U25675 (N_25675,N_24517,N_24624);
nand U25676 (N_25676,N_24157,N_24304);
nand U25677 (N_25677,N_24953,N_24016);
and U25678 (N_25678,N_24317,N_24586);
or U25679 (N_25679,N_24776,N_24888);
and U25680 (N_25680,N_24607,N_24061);
nand U25681 (N_25681,N_24394,N_24675);
nand U25682 (N_25682,N_24736,N_24971);
xor U25683 (N_25683,N_24686,N_24682);
nor U25684 (N_25684,N_24655,N_24698);
or U25685 (N_25685,N_24445,N_24428);
nor U25686 (N_25686,N_24335,N_24324);
nor U25687 (N_25687,N_24866,N_24978);
xnor U25688 (N_25688,N_24611,N_24619);
or U25689 (N_25689,N_24304,N_24211);
and U25690 (N_25690,N_24715,N_24204);
xnor U25691 (N_25691,N_24472,N_24630);
or U25692 (N_25692,N_24988,N_24439);
nand U25693 (N_25693,N_24603,N_24945);
xor U25694 (N_25694,N_24039,N_24973);
or U25695 (N_25695,N_24760,N_24969);
and U25696 (N_25696,N_24170,N_24661);
xor U25697 (N_25697,N_24082,N_24263);
and U25698 (N_25698,N_24490,N_24522);
and U25699 (N_25699,N_24497,N_24508);
nand U25700 (N_25700,N_24591,N_24224);
or U25701 (N_25701,N_24183,N_24786);
and U25702 (N_25702,N_24047,N_24708);
nand U25703 (N_25703,N_24944,N_24147);
or U25704 (N_25704,N_24864,N_24424);
xor U25705 (N_25705,N_24802,N_24545);
xor U25706 (N_25706,N_24542,N_24943);
nor U25707 (N_25707,N_24606,N_24486);
nor U25708 (N_25708,N_24000,N_24380);
nand U25709 (N_25709,N_24314,N_24255);
nand U25710 (N_25710,N_24905,N_24154);
nand U25711 (N_25711,N_24939,N_24891);
nor U25712 (N_25712,N_24221,N_24325);
nand U25713 (N_25713,N_24871,N_24611);
xor U25714 (N_25714,N_24824,N_24075);
nor U25715 (N_25715,N_24233,N_24036);
nor U25716 (N_25716,N_24470,N_24010);
nand U25717 (N_25717,N_24749,N_24319);
and U25718 (N_25718,N_24274,N_24759);
xor U25719 (N_25719,N_24742,N_24895);
or U25720 (N_25720,N_24926,N_24385);
nand U25721 (N_25721,N_24531,N_24018);
or U25722 (N_25722,N_24290,N_24288);
and U25723 (N_25723,N_24445,N_24593);
and U25724 (N_25724,N_24336,N_24636);
xor U25725 (N_25725,N_24439,N_24697);
or U25726 (N_25726,N_24671,N_24785);
xor U25727 (N_25727,N_24562,N_24635);
or U25728 (N_25728,N_24734,N_24068);
nand U25729 (N_25729,N_24022,N_24632);
nor U25730 (N_25730,N_24190,N_24566);
nand U25731 (N_25731,N_24793,N_24588);
xnor U25732 (N_25732,N_24151,N_24835);
and U25733 (N_25733,N_24864,N_24742);
and U25734 (N_25734,N_24581,N_24084);
nand U25735 (N_25735,N_24670,N_24303);
xor U25736 (N_25736,N_24011,N_24613);
nand U25737 (N_25737,N_24287,N_24800);
nand U25738 (N_25738,N_24417,N_24832);
xnor U25739 (N_25739,N_24091,N_24472);
nand U25740 (N_25740,N_24487,N_24788);
nor U25741 (N_25741,N_24416,N_24852);
or U25742 (N_25742,N_24562,N_24951);
and U25743 (N_25743,N_24938,N_24469);
nor U25744 (N_25744,N_24095,N_24693);
and U25745 (N_25745,N_24596,N_24948);
or U25746 (N_25746,N_24217,N_24613);
nor U25747 (N_25747,N_24252,N_24690);
nor U25748 (N_25748,N_24810,N_24229);
nor U25749 (N_25749,N_24239,N_24909);
or U25750 (N_25750,N_24036,N_24676);
xor U25751 (N_25751,N_24448,N_24185);
xor U25752 (N_25752,N_24053,N_24318);
nand U25753 (N_25753,N_24766,N_24925);
nand U25754 (N_25754,N_24655,N_24027);
and U25755 (N_25755,N_24159,N_24633);
or U25756 (N_25756,N_24618,N_24914);
or U25757 (N_25757,N_24803,N_24733);
or U25758 (N_25758,N_24804,N_24727);
nand U25759 (N_25759,N_24906,N_24345);
xor U25760 (N_25760,N_24211,N_24759);
and U25761 (N_25761,N_24094,N_24862);
or U25762 (N_25762,N_24559,N_24443);
nor U25763 (N_25763,N_24420,N_24669);
or U25764 (N_25764,N_24530,N_24707);
nand U25765 (N_25765,N_24267,N_24684);
nor U25766 (N_25766,N_24025,N_24226);
nand U25767 (N_25767,N_24207,N_24645);
nor U25768 (N_25768,N_24962,N_24745);
or U25769 (N_25769,N_24026,N_24097);
xor U25770 (N_25770,N_24555,N_24212);
and U25771 (N_25771,N_24114,N_24826);
or U25772 (N_25772,N_24749,N_24614);
or U25773 (N_25773,N_24687,N_24065);
nand U25774 (N_25774,N_24970,N_24853);
xnor U25775 (N_25775,N_24457,N_24143);
and U25776 (N_25776,N_24126,N_24766);
or U25777 (N_25777,N_24383,N_24204);
or U25778 (N_25778,N_24162,N_24918);
nor U25779 (N_25779,N_24377,N_24392);
nand U25780 (N_25780,N_24303,N_24424);
nand U25781 (N_25781,N_24295,N_24507);
and U25782 (N_25782,N_24543,N_24852);
xnor U25783 (N_25783,N_24176,N_24702);
and U25784 (N_25784,N_24159,N_24385);
or U25785 (N_25785,N_24914,N_24943);
xnor U25786 (N_25786,N_24179,N_24662);
nand U25787 (N_25787,N_24296,N_24839);
or U25788 (N_25788,N_24535,N_24057);
or U25789 (N_25789,N_24847,N_24715);
and U25790 (N_25790,N_24685,N_24930);
and U25791 (N_25791,N_24335,N_24931);
nor U25792 (N_25792,N_24349,N_24926);
nand U25793 (N_25793,N_24487,N_24716);
nor U25794 (N_25794,N_24578,N_24411);
nand U25795 (N_25795,N_24114,N_24655);
or U25796 (N_25796,N_24010,N_24905);
xnor U25797 (N_25797,N_24569,N_24401);
nor U25798 (N_25798,N_24643,N_24578);
or U25799 (N_25799,N_24264,N_24941);
nor U25800 (N_25800,N_24023,N_24520);
or U25801 (N_25801,N_24552,N_24294);
xor U25802 (N_25802,N_24640,N_24302);
xor U25803 (N_25803,N_24819,N_24224);
nand U25804 (N_25804,N_24343,N_24161);
and U25805 (N_25805,N_24570,N_24273);
and U25806 (N_25806,N_24610,N_24426);
or U25807 (N_25807,N_24614,N_24855);
or U25808 (N_25808,N_24457,N_24192);
xor U25809 (N_25809,N_24801,N_24430);
nand U25810 (N_25810,N_24500,N_24056);
nor U25811 (N_25811,N_24039,N_24968);
nor U25812 (N_25812,N_24375,N_24417);
and U25813 (N_25813,N_24656,N_24924);
nand U25814 (N_25814,N_24319,N_24467);
nand U25815 (N_25815,N_24233,N_24136);
xor U25816 (N_25816,N_24297,N_24937);
or U25817 (N_25817,N_24561,N_24605);
xor U25818 (N_25818,N_24003,N_24952);
nand U25819 (N_25819,N_24423,N_24103);
xnor U25820 (N_25820,N_24922,N_24506);
and U25821 (N_25821,N_24441,N_24245);
nand U25822 (N_25822,N_24532,N_24073);
and U25823 (N_25823,N_24267,N_24633);
and U25824 (N_25824,N_24627,N_24195);
nand U25825 (N_25825,N_24649,N_24761);
nand U25826 (N_25826,N_24387,N_24030);
and U25827 (N_25827,N_24960,N_24143);
xnor U25828 (N_25828,N_24185,N_24415);
nand U25829 (N_25829,N_24889,N_24230);
or U25830 (N_25830,N_24464,N_24541);
and U25831 (N_25831,N_24811,N_24188);
nor U25832 (N_25832,N_24796,N_24434);
nand U25833 (N_25833,N_24189,N_24204);
nand U25834 (N_25834,N_24226,N_24393);
or U25835 (N_25835,N_24388,N_24146);
and U25836 (N_25836,N_24271,N_24780);
and U25837 (N_25837,N_24253,N_24666);
nand U25838 (N_25838,N_24789,N_24810);
xnor U25839 (N_25839,N_24854,N_24410);
and U25840 (N_25840,N_24004,N_24546);
and U25841 (N_25841,N_24394,N_24738);
nor U25842 (N_25842,N_24876,N_24327);
and U25843 (N_25843,N_24789,N_24279);
xor U25844 (N_25844,N_24756,N_24933);
or U25845 (N_25845,N_24080,N_24500);
and U25846 (N_25846,N_24807,N_24218);
nand U25847 (N_25847,N_24539,N_24631);
nor U25848 (N_25848,N_24857,N_24960);
nor U25849 (N_25849,N_24066,N_24534);
or U25850 (N_25850,N_24002,N_24885);
and U25851 (N_25851,N_24425,N_24195);
nor U25852 (N_25852,N_24470,N_24891);
nand U25853 (N_25853,N_24482,N_24116);
or U25854 (N_25854,N_24090,N_24441);
xnor U25855 (N_25855,N_24105,N_24524);
or U25856 (N_25856,N_24861,N_24910);
xor U25857 (N_25857,N_24461,N_24077);
nor U25858 (N_25858,N_24344,N_24779);
xnor U25859 (N_25859,N_24558,N_24872);
nand U25860 (N_25860,N_24600,N_24595);
or U25861 (N_25861,N_24233,N_24003);
nand U25862 (N_25862,N_24889,N_24265);
nor U25863 (N_25863,N_24339,N_24237);
nor U25864 (N_25864,N_24086,N_24396);
and U25865 (N_25865,N_24050,N_24436);
and U25866 (N_25866,N_24460,N_24096);
or U25867 (N_25867,N_24550,N_24519);
nand U25868 (N_25868,N_24507,N_24501);
nor U25869 (N_25869,N_24010,N_24262);
or U25870 (N_25870,N_24003,N_24596);
nand U25871 (N_25871,N_24710,N_24612);
nor U25872 (N_25872,N_24061,N_24209);
nor U25873 (N_25873,N_24492,N_24673);
nor U25874 (N_25874,N_24345,N_24263);
and U25875 (N_25875,N_24245,N_24268);
and U25876 (N_25876,N_24455,N_24471);
nor U25877 (N_25877,N_24174,N_24832);
xnor U25878 (N_25878,N_24834,N_24470);
nand U25879 (N_25879,N_24242,N_24329);
or U25880 (N_25880,N_24000,N_24715);
and U25881 (N_25881,N_24118,N_24333);
or U25882 (N_25882,N_24623,N_24604);
or U25883 (N_25883,N_24144,N_24258);
nor U25884 (N_25884,N_24079,N_24942);
or U25885 (N_25885,N_24893,N_24747);
nor U25886 (N_25886,N_24729,N_24769);
nor U25887 (N_25887,N_24712,N_24694);
or U25888 (N_25888,N_24649,N_24610);
or U25889 (N_25889,N_24159,N_24667);
or U25890 (N_25890,N_24839,N_24659);
nor U25891 (N_25891,N_24319,N_24543);
nor U25892 (N_25892,N_24770,N_24729);
or U25893 (N_25893,N_24982,N_24955);
or U25894 (N_25894,N_24279,N_24579);
or U25895 (N_25895,N_24101,N_24524);
nor U25896 (N_25896,N_24924,N_24585);
nor U25897 (N_25897,N_24273,N_24075);
xor U25898 (N_25898,N_24321,N_24074);
xnor U25899 (N_25899,N_24940,N_24535);
nand U25900 (N_25900,N_24771,N_24149);
nand U25901 (N_25901,N_24167,N_24038);
and U25902 (N_25902,N_24963,N_24247);
xor U25903 (N_25903,N_24143,N_24269);
or U25904 (N_25904,N_24480,N_24908);
or U25905 (N_25905,N_24273,N_24193);
or U25906 (N_25906,N_24705,N_24425);
nand U25907 (N_25907,N_24752,N_24028);
nand U25908 (N_25908,N_24615,N_24375);
or U25909 (N_25909,N_24897,N_24253);
or U25910 (N_25910,N_24449,N_24346);
and U25911 (N_25911,N_24200,N_24180);
nand U25912 (N_25912,N_24241,N_24121);
nand U25913 (N_25913,N_24696,N_24940);
or U25914 (N_25914,N_24970,N_24154);
xor U25915 (N_25915,N_24679,N_24589);
nor U25916 (N_25916,N_24666,N_24094);
and U25917 (N_25917,N_24904,N_24273);
or U25918 (N_25918,N_24037,N_24094);
nand U25919 (N_25919,N_24005,N_24971);
nand U25920 (N_25920,N_24443,N_24412);
or U25921 (N_25921,N_24533,N_24964);
or U25922 (N_25922,N_24324,N_24261);
and U25923 (N_25923,N_24840,N_24655);
nor U25924 (N_25924,N_24688,N_24078);
and U25925 (N_25925,N_24258,N_24212);
and U25926 (N_25926,N_24625,N_24546);
and U25927 (N_25927,N_24947,N_24474);
nor U25928 (N_25928,N_24307,N_24656);
nand U25929 (N_25929,N_24848,N_24412);
xor U25930 (N_25930,N_24645,N_24478);
nand U25931 (N_25931,N_24601,N_24690);
or U25932 (N_25932,N_24644,N_24360);
nand U25933 (N_25933,N_24793,N_24279);
xnor U25934 (N_25934,N_24358,N_24228);
nand U25935 (N_25935,N_24298,N_24035);
and U25936 (N_25936,N_24977,N_24126);
or U25937 (N_25937,N_24834,N_24123);
nand U25938 (N_25938,N_24160,N_24403);
and U25939 (N_25939,N_24657,N_24074);
nand U25940 (N_25940,N_24161,N_24845);
and U25941 (N_25941,N_24734,N_24765);
xor U25942 (N_25942,N_24911,N_24148);
nor U25943 (N_25943,N_24208,N_24069);
xnor U25944 (N_25944,N_24498,N_24326);
nor U25945 (N_25945,N_24418,N_24675);
or U25946 (N_25946,N_24711,N_24618);
and U25947 (N_25947,N_24337,N_24169);
or U25948 (N_25948,N_24453,N_24884);
or U25949 (N_25949,N_24534,N_24629);
xnor U25950 (N_25950,N_24332,N_24046);
xnor U25951 (N_25951,N_24433,N_24518);
nand U25952 (N_25952,N_24670,N_24173);
xnor U25953 (N_25953,N_24463,N_24479);
xor U25954 (N_25954,N_24796,N_24997);
xor U25955 (N_25955,N_24544,N_24210);
or U25956 (N_25956,N_24857,N_24054);
or U25957 (N_25957,N_24487,N_24991);
or U25958 (N_25958,N_24878,N_24658);
nand U25959 (N_25959,N_24595,N_24044);
and U25960 (N_25960,N_24420,N_24621);
or U25961 (N_25961,N_24706,N_24772);
and U25962 (N_25962,N_24900,N_24743);
xor U25963 (N_25963,N_24015,N_24703);
nor U25964 (N_25964,N_24439,N_24965);
or U25965 (N_25965,N_24134,N_24372);
or U25966 (N_25966,N_24072,N_24271);
nand U25967 (N_25967,N_24664,N_24919);
xnor U25968 (N_25968,N_24258,N_24252);
xnor U25969 (N_25969,N_24379,N_24072);
xor U25970 (N_25970,N_24423,N_24341);
and U25971 (N_25971,N_24687,N_24288);
nor U25972 (N_25972,N_24440,N_24572);
nand U25973 (N_25973,N_24022,N_24184);
xor U25974 (N_25974,N_24797,N_24583);
nor U25975 (N_25975,N_24256,N_24747);
and U25976 (N_25976,N_24485,N_24716);
xnor U25977 (N_25977,N_24972,N_24694);
nor U25978 (N_25978,N_24407,N_24583);
xnor U25979 (N_25979,N_24369,N_24480);
and U25980 (N_25980,N_24956,N_24723);
nand U25981 (N_25981,N_24422,N_24835);
and U25982 (N_25982,N_24830,N_24572);
and U25983 (N_25983,N_24593,N_24324);
nor U25984 (N_25984,N_24821,N_24520);
nand U25985 (N_25985,N_24582,N_24471);
nand U25986 (N_25986,N_24803,N_24374);
xnor U25987 (N_25987,N_24625,N_24492);
nor U25988 (N_25988,N_24150,N_24670);
xnor U25989 (N_25989,N_24381,N_24696);
xor U25990 (N_25990,N_24324,N_24235);
nor U25991 (N_25991,N_24081,N_24789);
or U25992 (N_25992,N_24336,N_24470);
nand U25993 (N_25993,N_24814,N_24381);
and U25994 (N_25994,N_24583,N_24360);
xnor U25995 (N_25995,N_24174,N_24042);
and U25996 (N_25996,N_24965,N_24717);
xnor U25997 (N_25997,N_24887,N_24595);
or U25998 (N_25998,N_24090,N_24630);
nand U25999 (N_25999,N_24815,N_24592);
and U26000 (N_26000,N_25903,N_25696);
nor U26001 (N_26001,N_25389,N_25534);
nand U26002 (N_26002,N_25437,N_25991);
nor U26003 (N_26003,N_25406,N_25070);
nand U26004 (N_26004,N_25046,N_25498);
and U26005 (N_26005,N_25178,N_25977);
nand U26006 (N_26006,N_25999,N_25659);
and U26007 (N_26007,N_25061,N_25203);
nand U26008 (N_26008,N_25719,N_25740);
xor U26009 (N_26009,N_25741,N_25876);
xnor U26010 (N_26010,N_25006,N_25086);
nand U26011 (N_26011,N_25867,N_25956);
nor U26012 (N_26012,N_25811,N_25017);
or U26013 (N_26013,N_25935,N_25943);
or U26014 (N_26014,N_25632,N_25299);
or U26015 (N_26015,N_25872,N_25553);
and U26016 (N_26016,N_25206,N_25924);
nor U26017 (N_26017,N_25704,N_25733);
and U26018 (N_26018,N_25367,N_25635);
and U26019 (N_26019,N_25947,N_25079);
xor U26020 (N_26020,N_25020,N_25929);
nor U26021 (N_26021,N_25010,N_25769);
nor U26022 (N_26022,N_25001,N_25892);
or U26023 (N_26023,N_25877,N_25096);
nor U26024 (N_26024,N_25965,N_25103);
xor U26025 (N_26025,N_25126,N_25717);
nand U26026 (N_26026,N_25312,N_25617);
xor U26027 (N_26027,N_25187,N_25400);
nor U26028 (N_26028,N_25621,N_25958);
xor U26029 (N_26029,N_25109,N_25906);
nand U26030 (N_26030,N_25328,N_25893);
or U26031 (N_26031,N_25597,N_25219);
nor U26032 (N_26032,N_25532,N_25468);
xnor U26033 (N_26033,N_25970,N_25535);
nor U26034 (N_26034,N_25923,N_25244);
xnor U26035 (N_26035,N_25317,N_25979);
or U26036 (N_26036,N_25194,N_25052);
and U26037 (N_26037,N_25922,N_25557);
or U26038 (N_26038,N_25916,N_25292);
nor U26039 (N_26039,N_25706,N_25209);
and U26040 (N_26040,N_25141,N_25624);
and U26041 (N_26041,N_25119,N_25786);
xnor U26042 (N_26042,N_25423,N_25134);
and U26043 (N_26043,N_25792,N_25607);
and U26044 (N_26044,N_25165,N_25365);
or U26045 (N_26045,N_25401,N_25510);
nor U26046 (N_26046,N_25580,N_25176);
nor U26047 (N_26047,N_25179,N_25403);
xnor U26048 (N_26048,N_25461,N_25730);
and U26049 (N_26049,N_25613,N_25930);
nor U26050 (N_26050,N_25612,N_25408);
xor U26051 (N_26051,N_25314,N_25253);
nor U26052 (N_26052,N_25186,N_25819);
xnor U26053 (N_26053,N_25752,N_25684);
and U26054 (N_26054,N_25793,N_25368);
nor U26055 (N_26055,N_25871,N_25963);
and U26056 (N_26056,N_25654,N_25810);
nor U26057 (N_26057,N_25080,N_25508);
or U26058 (N_26058,N_25236,N_25993);
xor U26059 (N_26059,N_25911,N_25854);
or U26060 (N_26060,N_25525,N_25962);
xnor U26061 (N_26061,N_25651,N_25297);
xnor U26062 (N_26062,N_25550,N_25638);
nand U26063 (N_26063,N_25715,N_25425);
nor U26064 (N_26064,N_25435,N_25390);
xnor U26065 (N_26065,N_25371,N_25265);
nor U26066 (N_26066,N_25216,N_25732);
or U26067 (N_26067,N_25776,N_25346);
nor U26068 (N_26068,N_25227,N_25658);
and U26069 (N_26069,N_25074,N_25538);
or U26070 (N_26070,N_25493,N_25116);
nand U26071 (N_26071,N_25221,N_25767);
and U26072 (N_26072,N_25479,N_25177);
or U26073 (N_26073,N_25279,N_25112);
nand U26074 (N_26074,N_25783,N_25688);
and U26075 (N_26075,N_25683,N_25814);
and U26076 (N_26076,N_25466,N_25207);
nand U26077 (N_26077,N_25832,N_25705);
nor U26078 (N_26078,N_25761,N_25238);
xor U26079 (N_26079,N_25222,N_25816);
nor U26080 (N_26080,N_25572,N_25024);
nand U26081 (N_26081,N_25589,N_25306);
or U26082 (N_26082,N_25931,N_25802);
or U26083 (N_26083,N_25100,N_25671);
and U26084 (N_26084,N_25462,N_25322);
xor U26085 (N_26085,N_25862,N_25066);
and U26086 (N_26086,N_25155,N_25307);
nor U26087 (N_26087,N_25590,N_25555);
xor U26088 (N_26088,N_25459,N_25012);
nand U26089 (N_26089,N_25541,N_25554);
xnor U26090 (N_26090,N_25797,N_25829);
and U26091 (N_26091,N_25057,N_25825);
nor U26092 (N_26092,N_25765,N_25353);
xnor U26093 (N_26093,N_25032,N_25240);
nor U26094 (N_26094,N_25626,N_25218);
nand U26095 (N_26095,N_25600,N_25151);
nand U26096 (N_26096,N_25455,N_25150);
nand U26097 (N_26097,N_25154,N_25350);
nand U26098 (N_26098,N_25491,N_25304);
or U26099 (N_26099,N_25475,N_25087);
or U26100 (N_26100,N_25526,N_25620);
nand U26101 (N_26101,N_25161,N_25137);
or U26102 (N_26102,N_25905,N_25095);
or U26103 (N_26103,N_25665,N_25714);
nor U26104 (N_26104,N_25038,N_25196);
nand U26105 (N_26105,N_25896,N_25851);
and U26106 (N_26106,N_25485,N_25125);
or U26107 (N_26107,N_25327,N_25047);
nand U26108 (N_26108,N_25500,N_25738);
xor U26109 (N_26109,N_25642,N_25961);
nand U26110 (N_26110,N_25439,N_25586);
xnor U26111 (N_26111,N_25633,N_25022);
nor U26112 (N_26112,N_25992,N_25914);
nor U26113 (N_26113,N_25595,N_25064);
xor U26114 (N_26114,N_25140,N_25364);
and U26115 (N_26115,N_25634,N_25679);
nand U26116 (N_26116,N_25477,N_25003);
and U26117 (N_26117,N_25989,N_25413);
or U26118 (N_26118,N_25859,N_25982);
and U26119 (N_26119,N_25676,N_25523);
xnor U26120 (N_26120,N_25894,N_25536);
nor U26121 (N_26121,N_25139,N_25252);
nand U26122 (N_26122,N_25019,N_25639);
nand U26123 (N_26123,N_25015,N_25418);
xnor U26124 (N_26124,N_25565,N_25849);
or U26125 (N_26125,N_25920,N_25381);
nor U26126 (N_26126,N_25083,N_25614);
xnor U26127 (N_26127,N_25185,N_25382);
or U26128 (N_26128,N_25640,N_25169);
or U26129 (N_26129,N_25972,N_25035);
nand U26130 (N_26130,N_25582,N_25104);
or U26131 (N_26131,N_25084,N_25742);
xnor U26132 (N_26132,N_25369,N_25444);
nand U26133 (N_26133,N_25611,N_25801);
nor U26134 (N_26134,N_25421,N_25530);
or U26135 (N_26135,N_25440,N_25649);
nor U26136 (N_26136,N_25197,N_25234);
nand U26137 (N_26137,N_25210,N_25443);
or U26138 (N_26138,N_25758,N_25743);
or U26139 (N_26139,N_25987,N_25942);
or U26140 (N_26140,N_25981,N_25148);
nor U26141 (N_26141,N_25745,N_25325);
nor U26142 (N_26142,N_25915,N_25492);
nor U26143 (N_26143,N_25152,N_25988);
nor U26144 (N_26144,N_25831,N_25330);
or U26145 (N_26145,N_25275,N_25108);
and U26146 (N_26146,N_25764,N_25564);
nand U26147 (N_26147,N_25997,N_25077);
or U26148 (N_26148,N_25636,N_25267);
and U26149 (N_26149,N_25242,N_25843);
or U26150 (N_26150,N_25653,N_25949);
nand U26151 (N_26151,N_25410,N_25718);
and U26152 (N_26152,N_25358,N_25448);
nand U26153 (N_26153,N_25841,N_25352);
or U26154 (N_26154,N_25546,N_25901);
or U26155 (N_26155,N_25030,N_25133);
xnor U26156 (N_26156,N_25575,N_25202);
or U26157 (N_26157,N_25127,N_25033);
nor U26158 (N_26158,N_25174,N_25781);
nand U26159 (N_26159,N_25506,N_25007);
nor U26160 (N_26160,N_25629,N_25789);
or U26161 (N_26161,N_25296,N_25168);
nand U26162 (N_26162,N_25496,N_25189);
nor U26163 (N_26163,N_25755,N_25147);
and U26164 (N_26164,N_25599,N_25505);
xor U26165 (N_26165,N_25584,N_25043);
or U26166 (N_26166,N_25908,N_25384);
xnor U26167 (N_26167,N_25039,N_25656);
xnor U26168 (N_26168,N_25310,N_25604);
xor U26169 (N_26169,N_25192,N_25858);
nand U26170 (N_26170,N_25092,N_25559);
nand U26171 (N_26171,N_25662,N_25374);
nand U26172 (N_26172,N_25644,N_25677);
nor U26173 (N_26173,N_25311,N_25701);
nand U26174 (N_26174,N_25837,N_25934);
nand U26175 (N_26175,N_25246,N_25652);
and U26176 (N_26176,N_25787,N_25980);
xnor U26177 (N_26177,N_25806,N_25808);
nand U26178 (N_26178,N_25848,N_25021);
xor U26179 (N_26179,N_25143,N_25592);
and U26180 (N_26180,N_25105,N_25868);
nand U26181 (N_26181,N_25135,N_25347);
xnor U26182 (N_26182,N_25875,N_25531);
or U26183 (N_26183,N_25616,N_25995);
or U26184 (N_26184,N_25295,N_25857);
xor U26185 (N_26185,N_25373,N_25902);
nor U26186 (N_26186,N_25458,N_25453);
nor U26187 (N_26187,N_25254,N_25520);
or U26188 (N_26188,N_25290,N_25243);
xor U26189 (N_26189,N_25158,N_25720);
nor U26190 (N_26190,N_25372,N_25724);
nand U26191 (N_26191,N_25261,N_25008);
and U26192 (N_26192,N_25514,N_25476);
or U26193 (N_26193,N_25250,N_25142);
and U26194 (N_26194,N_25521,N_25966);
xnor U26195 (N_26195,N_25433,N_25932);
or U26196 (N_26196,N_25434,N_25208);
nand U26197 (N_26197,N_25089,N_25130);
nand U26198 (N_26198,N_25537,N_25885);
xor U26199 (N_26199,N_25159,N_25248);
and U26200 (N_26200,N_25578,N_25097);
nor U26201 (N_26201,N_25771,N_25257);
or U26202 (N_26202,N_25345,N_25473);
nand U26203 (N_26203,N_25315,N_25303);
nand U26204 (N_26204,N_25274,N_25646);
nor U26205 (N_26205,N_25952,N_25588);
nor U26206 (N_26206,N_25669,N_25082);
xnor U26207 (N_26207,N_25772,N_25376);
xor U26208 (N_26208,N_25570,N_25175);
xnor U26209 (N_26209,N_25812,N_25280);
nand U26210 (N_26210,N_25391,N_25123);
nor U26211 (N_26211,N_25224,N_25115);
nor U26212 (N_26212,N_25497,N_25409);
xor U26213 (N_26213,N_25484,N_25971);
xor U26214 (N_26214,N_25018,N_25886);
nor U26215 (N_26215,N_25454,N_25517);
nor U26216 (N_26216,N_25360,N_25681);
xnor U26217 (N_26217,N_25320,N_25321);
nor U26218 (N_26218,N_25182,N_25533);
nor U26219 (N_26219,N_25263,N_25446);
xnor U26220 (N_26220,N_25556,N_25298);
nand U26221 (N_26221,N_25850,N_25566);
xor U26222 (N_26222,N_25957,N_25846);
xnor U26223 (N_26223,N_25258,N_25205);
nand U26224 (N_26224,N_25260,N_25648);
nor U26225 (N_26225,N_25287,N_25799);
xor U26226 (N_26226,N_25342,N_25983);
and U26227 (N_26227,N_25204,N_25445);
or U26228 (N_26228,N_25839,N_25073);
or U26229 (N_26229,N_25266,N_25004);
or U26230 (N_26230,N_25734,N_25309);
and U26231 (N_26231,N_25820,N_25936);
xnor U26232 (N_26232,N_25900,N_25464);
and U26233 (N_26233,N_25774,N_25005);
nand U26234 (N_26234,N_25044,N_25927);
nor U26235 (N_26235,N_25072,N_25488);
nand U26236 (N_26236,N_25552,N_25231);
nor U26237 (N_26237,N_25946,N_25838);
nor U26238 (N_26238,N_25377,N_25643);
nand U26239 (N_26239,N_25341,N_25667);
nor U26240 (N_26240,N_25507,N_25645);
xnor U26241 (N_26241,N_25269,N_25707);
and U26242 (N_26242,N_25913,N_25069);
and U26243 (N_26243,N_25235,N_25378);
and U26244 (N_26244,N_25756,N_25091);
nor U26245 (N_26245,N_25388,N_25528);
or U26246 (N_26246,N_25031,N_25598);
nand U26247 (N_26247,N_25319,N_25355);
nor U26248 (N_26248,N_25694,N_25145);
nand U26249 (N_26249,N_25777,N_25385);
or U26250 (N_26250,N_25994,N_25561);
nand U26251 (N_26251,N_25285,N_25288);
and U26252 (N_26252,N_25845,N_25291);
nand U26253 (N_26253,N_25809,N_25655);
and U26254 (N_26254,N_25065,N_25725);
nand U26255 (N_26255,N_25502,N_25703);
nand U26256 (N_26256,N_25869,N_25713);
or U26257 (N_26257,N_25770,N_25121);
nand U26258 (N_26258,N_25805,N_25996);
or U26259 (N_26259,N_25576,N_25283);
nor U26260 (N_26260,N_25751,N_25215);
and U26261 (N_26261,N_25630,N_25501);
nor U26262 (N_26262,N_25499,N_25230);
or U26263 (N_26263,N_25264,N_25563);
nor U26264 (N_26264,N_25474,N_25791);
xor U26265 (N_26265,N_25495,N_25313);
xor U26266 (N_26266,N_25359,N_25747);
nor U26267 (N_26267,N_25153,N_25217);
and U26268 (N_26268,N_25270,N_25339);
nor U26269 (N_26269,N_25504,N_25754);
nor U26270 (N_26270,N_25370,N_25471);
nor U26271 (N_26271,N_25700,N_25000);
and U26272 (N_26272,N_25099,N_25904);
and U26273 (N_26273,N_25860,N_25796);
and U26274 (N_26274,N_25071,N_25735);
or U26275 (N_26275,N_25807,N_25329);
and U26276 (N_26276,N_25657,N_25214);
xor U26277 (N_26277,N_25124,N_25262);
xor U26278 (N_26278,N_25239,N_25933);
and U26279 (N_26279,N_25702,N_25232);
xor U26280 (N_26280,N_25699,N_25027);
and U26281 (N_26281,N_25171,N_25647);
xor U26282 (N_26282,N_25835,N_25773);
nor U26283 (N_26283,N_25416,N_25737);
xnor U26284 (N_26284,N_25241,N_25025);
nor U26285 (N_26285,N_25058,N_25918);
or U26286 (N_26286,N_25910,N_25387);
nor U26287 (N_26287,N_25300,N_25467);
or U26288 (N_26288,N_25316,N_25011);
nand U26289 (N_26289,N_25690,N_25014);
nor U26290 (N_26290,N_25420,N_25427);
nor U26291 (N_26291,N_25394,N_25237);
or U26292 (N_26292,N_25511,N_25063);
xor U26293 (N_26293,N_25272,N_25571);
nor U26294 (N_26294,N_25088,N_25973);
or U26295 (N_26295,N_25487,N_25641);
nand U26296 (N_26296,N_25698,N_25509);
nand U26297 (N_26297,N_25053,N_25489);
or U26298 (N_26298,N_25967,N_25190);
nand U26299 (N_26299,N_25650,N_25748);
xor U26300 (N_26300,N_25276,N_25251);
or U26301 (N_26301,N_25693,N_25023);
and U26302 (N_26302,N_25986,N_25397);
nand U26303 (N_26303,N_25357,N_25048);
nand U26304 (N_26304,N_25193,N_25131);
or U26305 (N_26305,N_25567,N_25037);
nand U26306 (N_26306,N_25938,N_25824);
or U26307 (N_26307,N_25891,N_25460);
nand U26308 (N_26308,N_25138,N_25895);
or U26309 (N_26309,N_25395,N_25551);
nand U26310 (N_26310,N_25853,N_25823);
nor U26311 (N_26311,N_25587,N_25094);
and U26312 (N_26312,N_25919,N_25188);
nand U26313 (N_26313,N_25324,N_25211);
and U26314 (N_26314,N_25762,N_25054);
xnor U26315 (N_26315,N_25842,N_25928);
xor U26316 (N_26316,N_25463,N_25569);
or U26317 (N_26317,N_25163,N_25990);
nor U26318 (N_26318,N_25481,N_25465);
and U26319 (N_26319,N_25596,N_25132);
or U26320 (N_26320,N_25513,N_25674);
nor U26321 (N_26321,N_25539,N_25631);
nor U26322 (N_26322,N_25436,N_25579);
nor U26323 (N_26323,N_25430,N_25255);
and U26324 (N_26324,N_25195,N_25670);
nand U26325 (N_26325,N_25076,N_25954);
and U26326 (N_26326,N_25028,N_25804);
or U26327 (N_26327,N_25583,N_25785);
nand U26328 (N_26328,N_25009,N_25861);
or U26329 (N_26329,N_25759,N_25482);
xnor U26330 (N_26330,N_25338,N_25542);
nor U26331 (N_26331,N_25226,N_25380);
nand U26332 (N_26332,N_25167,N_25379);
nor U26333 (N_26333,N_25739,N_25917);
and U26334 (N_26334,N_25680,N_25974);
or U26335 (N_26335,N_25172,N_25697);
nor U26336 (N_26336,N_25308,N_25431);
nor U26337 (N_26337,N_25398,N_25518);
and U26338 (N_26338,N_25191,N_25623);
and U26339 (N_26339,N_25029,N_25627);
and U26340 (N_26340,N_25181,N_25815);
nand U26341 (N_26341,N_25950,N_25183);
or U26342 (N_26342,N_25289,N_25899);
xor U26343 (N_26343,N_25594,N_25136);
and U26344 (N_26344,N_25457,N_25666);
or U26345 (N_26345,N_25273,N_25162);
and U26346 (N_26346,N_25673,N_25780);
and U26347 (N_26347,N_25516,N_25603);
xor U26348 (N_26348,N_25784,N_25056);
and U26349 (N_26349,N_25062,N_25494);
and U26350 (N_26350,N_25736,N_25146);
and U26351 (N_26351,N_25075,N_25326);
or U26352 (N_26352,N_25618,N_25302);
and U26353 (N_26353,N_25349,N_25585);
nand U26354 (N_26354,N_25305,N_25548);
nand U26355 (N_26355,N_25955,N_25093);
or U26356 (N_26356,N_25549,N_25249);
nand U26357 (N_26357,N_25678,N_25716);
or U26358 (N_26358,N_25828,N_25881);
nor U26359 (N_26359,N_25711,N_25180);
and U26360 (N_26360,N_25944,N_25334);
nand U26361 (N_26361,N_25002,N_25422);
xor U26362 (N_26362,N_25301,N_25441);
nand U26363 (N_26363,N_25343,N_25726);
nand U26364 (N_26364,N_25813,N_25294);
and U26365 (N_26365,N_25055,N_25852);
or U26366 (N_26366,N_25951,N_25013);
and U26367 (N_26367,N_25577,N_25945);
nor U26368 (N_26368,N_25113,N_25386);
and U26369 (N_26369,N_25340,N_25512);
nor U26370 (N_26370,N_25562,N_25040);
xnor U26371 (N_26371,N_25429,N_25907);
nor U26372 (N_26372,N_25884,N_25268);
nand U26373 (N_26373,N_25602,N_25026);
or U26374 (N_26374,N_25964,N_25122);
nor U26375 (N_26375,N_25709,N_25689);
or U26376 (N_26376,N_25344,N_25247);
nor U26377 (N_26377,N_25478,N_25686);
and U26378 (N_26378,N_25201,N_25560);
and U26379 (N_26379,N_25515,N_25790);
nand U26380 (N_26380,N_25282,N_25503);
and U26381 (N_26381,N_25085,N_25415);
and U26382 (N_26382,N_25114,N_25608);
or U26383 (N_26383,N_25978,N_25794);
nand U26384 (N_26384,N_25129,N_25128);
nand U26385 (N_26385,N_25834,N_25890);
nand U26386 (N_26386,N_25050,N_25826);
or U26387 (N_26387,N_25685,N_25200);
nand U26388 (N_26388,N_25170,N_25428);
nand U26389 (N_26389,N_25847,N_25078);
xnor U26390 (N_26390,N_25591,N_25757);
and U26391 (N_26391,N_25975,N_25727);
nand U26392 (N_26392,N_25545,N_25225);
xor U26393 (N_26393,N_25863,N_25940);
and U26394 (N_26394,N_25354,N_25220);
xor U26395 (N_26395,N_25601,N_25414);
nor U26396 (N_26396,N_25160,N_25984);
nand U26397 (N_26397,N_25728,N_25278);
nand U26398 (N_26398,N_25897,N_25864);
nor U26399 (N_26399,N_25271,N_25404);
and U26400 (N_26400,N_25120,N_25438);
and U26401 (N_26401,N_25581,N_25909);
and U26402 (N_26402,N_25106,N_25332);
xnor U26403 (N_26403,N_25229,N_25912);
nor U26404 (N_26404,N_25941,N_25798);
and U26405 (N_26405,N_25879,N_25558);
xnor U26406 (N_26406,N_25959,N_25749);
or U26407 (N_26407,N_25800,N_25721);
and U26408 (N_26408,N_25760,N_25068);
nand U26409 (N_26409,N_25233,N_25383);
nor U26410 (N_26410,N_25985,N_25573);
nor U26411 (N_26411,N_25102,N_25118);
nor U26412 (N_26412,N_25331,N_25731);
and U26413 (N_26413,N_25953,N_25164);
and U26414 (N_26414,N_25111,N_25778);
nor U26415 (N_26415,N_25407,N_25782);
xor U26416 (N_26416,N_25323,N_25333);
and U26417 (N_26417,N_25199,N_25746);
nor U26418 (N_26418,N_25788,N_25042);
and U26419 (N_26419,N_25766,N_25873);
and U26420 (N_26420,N_25212,N_25779);
and U26421 (N_26421,N_25926,N_25149);
nor U26422 (N_26422,N_25744,N_25687);
nor U26423 (N_26423,N_25419,N_25016);
nand U26424 (N_26424,N_25432,N_25840);
xnor U26425 (N_26425,N_25543,N_25259);
nor U26426 (N_26426,N_25544,N_25540);
nand U26427 (N_26427,N_25098,N_25750);
or U26428 (N_26428,N_25049,N_25490);
nand U26429 (N_26429,N_25818,N_25472);
or U26430 (N_26430,N_25969,N_25483);
and U26431 (N_26431,N_25396,N_25664);
nor U26432 (N_26432,N_25405,N_25245);
and U26433 (N_26433,N_25609,N_25672);
and U26434 (N_26434,N_25878,N_25574);
nor U26435 (N_26435,N_25568,N_25480);
nand U26436 (N_26436,N_25855,N_25937);
or U26437 (N_26437,N_25411,N_25661);
nand U26438 (N_26438,N_25866,N_25695);
and U26439 (N_26439,N_25286,N_25803);
xor U26440 (N_26440,N_25622,N_25366);
nand U26441 (N_26441,N_25277,N_25045);
or U26442 (N_26442,N_25375,N_25844);
xor U26443 (N_26443,N_25392,N_25101);
or U26444 (N_26444,N_25469,N_25036);
nor U26445 (N_26445,N_25519,N_25865);
and U26446 (N_26446,N_25723,N_25921);
nor U26447 (N_26447,N_25522,N_25256);
nor U26448 (N_26448,N_25450,N_25668);
and U26449 (N_26449,N_25593,N_25691);
and U26450 (N_26450,N_25470,N_25775);
and U26451 (N_26451,N_25822,N_25402);
nor U26452 (N_26452,N_25060,N_25692);
nand U26453 (N_26453,N_25173,N_25817);
nor U26454 (N_26454,N_25090,N_25117);
nand U26455 (N_26455,N_25034,N_25361);
and U26456 (N_26456,N_25451,N_25281);
and U26457 (N_26457,N_25833,N_25663);
or U26458 (N_26458,N_25889,N_25293);
nor U26459 (N_26459,N_25335,N_25619);
nand U26460 (N_26460,N_25449,N_25628);
and U26461 (N_26461,N_25184,N_25874);
xor U26462 (N_26462,N_25753,N_25795);
nor U26463 (N_26463,N_25337,N_25393);
xor U26464 (N_26464,N_25960,N_25880);
and U26465 (N_26465,N_25948,N_25939);
xor U26466 (N_26466,N_25821,N_25998);
xor U26467 (N_26467,N_25486,N_25888);
and U26468 (N_26468,N_25051,N_25605);
nand U26469 (N_26469,N_25356,N_25336);
and U26470 (N_26470,N_25144,N_25363);
and U26471 (N_26471,N_25456,N_25198);
nor U26472 (N_26472,N_25156,N_25827);
or U26473 (N_26473,N_25527,N_25870);
and U26474 (N_26474,N_25660,N_25166);
xnor U26475 (N_26475,N_25318,N_25213);
nor U26476 (N_26476,N_25424,N_25615);
xnor U26477 (N_26477,N_25417,N_25524);
and U26478 (N_26478,N_25625,N_25768);
xnor U26479 (N_26479,N_25883,N_25348);
and U26480 (N_26480,N_25925,N_25081);
or U26481 (N_26481,N_25887,N_25107);
and U26482 (N_26482,N_25882,N_25399);
nor U26483 (N_26483,N_25610,N_25722);
and U26484 (N_26484,N_25708,N_25547);
and U26485 (N_26485,N_25452,N_25351);
xor U26486 (N_26486,N_25442,N_25447);
nor U26487 (N_26487,N_25606,N_25976);
nand U26488 (N_26488,N_25110,N_25712);
nand U26489 (N_26489,N_25675,N_25682);
nor U26490 (N_26490,N_25362,N_25898);
nand U26491 (N_26491,N_25830,N_25763);
and U26492 (N_26492,N_25412,N_25228);
and U26493 (N_26493,N_25041,N_25637);
or U26494 (N_26494,N_25284,N_25856);
nor U26495 (N_26495,N_25223,N_25710);
xnor U26496 (N_26496,N_25067,N_25426);
or U26497 (N_26497,N_25729,N_25059);
nand U26498 (N_26498,N_25529,N_25836);
nor U26499 (N_26499,N_25968,N_25157);
nand U26500 (N_26500,N_25963,N_25168);
and U26501 (N_26501,N_25163,N_25047);
nand U26502 (N_26502,N_25316,N_25547);
nor U26503 (N_26503,N_25877,N_25999);
nor U26504 (N_26504,N_25394,N_25123);
xnor U26505 (N_26505,N_25529,N_25381);
nor U26506 (N_26506,N_25540,N_25866);
nor U26507 (N_26507,N_25360,N_25168);
and U26508 (N_26508,N_25401,N_25315);
or U26509 (N_26509,N_25446,N_25225);
xnor U26510 (N_26510,N_25306,N_25232);
xor U26511 (N_26511,N_25200,N_25786);
nand U26512 (N_26512,N_25637,N_25517);
nor U26513 (N_26513,N_25817,N_25990);
xor U26514 (N_26514,N_25114,N_25457);
nand U26515 (N_26515,N_25016,N_25732);
or U26516 (N_26516,N_25131,N_25145);
xnor U26517 (N_26517,N_25736,N_25092);
or U26518 (N_26518,N_25770,N_25176);
and U26519 (N_26519,N_25014,N_25333);
xnor U26520 (N_26520,N_25481,N_25576);
xor U26521 (N_26521,N_25081,N_25307);
nor U26522 (N_26522,N_25182,N_25139);
xor U26523 (N_26523,N_25863,N_25590);
nor U26524 (N_26524,N_25457,N_25046);
or U26525 (N_26525,N_25203,N_25357);
xnor U26526 (N_26526,N_25128,N_25243);
nor U26527 (N_26527,N_25038,N_25187);
or U26528 (N_26528,N_25445,N_25378);
nand U26529 (N_26529,N_25139,N_25362);
nor U26530 (N_26530,N_25118,N_25714);
nor U26531 (N_26531,N_25449,N_25625);
nand U26532 (N_26532,N_25054,N_25697);
or U26533 (N_26533,N_25855,N_25744);
and U26534 (N_26534,N_25898,N_25077);
nand U26535 (N_26535,N_25510,N_25325);
or U26536 (N_26536,N_25156,N_25848);
or U26537 (N_26537,N_25156,N_25446);
xor U26538 (N_26538,N_25970,N_25282);
xnor U26539 (N_26539,N_25258,N_25103);
nand U26540 (N_26540,N_25515,N_25775);
nor U26541 (N_26541,N_25110,N_25172);
xor U26542 (N_26542,N_25408,N_25669);
or U26543 (N_26543,N_25339,N_25856);
or U26544 (N_26544,N_25901,N_25852);
or U26545 (N_26545,N_25822,N_25143);
nand U26546 (N_26546,N_25181,N_25191);
nor U26547 (N_26547,N_25490,N_25857);
nand U26548 (N_26548,N_25560,N_25564);
or U26549 (N_26549,N_25013,N_25025);
nand U26550 (N_26550,N_25659,N_25144);
nand U26551 (N_26551,N_25812,N_25760);
nor U26552 (N_26552,N_25833,N_25754);
or U26553 (N_26553,N_25686,N_25503);
nand U26554 (N_26554,N_25905,N_25523);
nor U26555 (N_26555,N_25351,N_25343);
nand U26556 (N_26556,N_25742,N_25743);
or U26557 (N_26557,N_25604,N_25817);
or U26558 (N_26558,N_25398,N_25993);
nand U26559 (N_26559,N_25907,N_25981);
or U26560 (N_26560,N_25361,N_25540);
nand U26561 (N_26561,N_25230,N_25718);
and U26562 (N_26562,N_25002,N_25914);
or U26563 (N_26563,N_25668,N_25180);
nor U26564 (N_26564,N_25205,N_25891);
xnor U26565 (N_26565,N_25830,N_25418);
or U26566 (N_26566,N_25731,N_25196);
xor U26567 (N_26567,N_25994,N_25123);
nor U26568 (N_26568,N_25221,N_25635);
nand U26569 (N_26569,N_25073,N_25490);
or U26570 (N_26570,N_25628,N_25147);
and U26571 (N_26571,N_25155,N_25562);
or U26572 (N_26572,N_25717,N_25924);
and U26573 (N_26573,N_25629,N_25995);
or U26574 (N_26574,N_25532,N_25016);
nor U26575 (N_26575,N_25096,N_25326);
and U26576 (N_26576,N_25710,N_25691);
nor U26577 (N_26577,N_25731,N_25327);
or U26578 (N_26578,N_25127,N_25323);
and U26579 (N_26579,N_25430,N_25349);
and U26580 (N_26580,N_25541,N_25283);
nor U26581 (N_26581,N_25886,N_25198);
and U26582 (N_26582,N_25140,N_25999);
or U26583 (N_26583,N_25075,N_25041);
nor U26584 (N_26584,N_25602,N_25533);
xnor U26585 (N_26585,N_25320,N_25815);
nand U26586 (N_26586,N_25636,N_25329);
nor U26587 (N_26587,N_25177,N_25979);
xnor U26588 (N_26588,N_25000,N_25046);
or U26589 (N_26589,N_25575,N_25680);
xor U26590 (N_26590,N_25369,N_25274);
xor U26591 (N_26591,N_25940,N_25230);
and U26592 (N_26592,N_25732,N_25593);
nor U26593 (N_26593,N_25976,N_25341);
or U26594 (N_26594,N_25719,N_25356);
or U26595 (N_26595,N_25127,N_25241);
or U26596 (N_26596,N_25739,N_25495);
or U26597 (N_26597,N_25008,N_25300);
or U26598 (N_26598,N_25757,N_25161);
nand U26599 (N_26599,N_25611,N_25530);
or U26600 (N_26600,N_25590,N_25952);
nor U26601 (N_26601,N_25772,N_25226);
nor U26602 (N_26602,N_25808,N_25881);
nand U26603 (N_26603,N_25932,N_25246);
nor U26604 (N_26604,N_25872,N_25124);
nand U26605 (N_26605,N_25540,N_25608);
and U26606 (N_26606,N_25146,N_25734);
xor U26607 (N_26607,N_25898,N_25254);
nand U26608 (N_26608,N_25485,N_25578);
nand U26609 (N_26609,N_25735,N_25504);
nor U26610 (N_26610,N_25782,N_25643);
or U26611 (N_26611,N_25717,N_25833);
or U26612 (N_26612,N_25746,N_25478);
and U26613 (N_26613,N_25785,N_25666);
nor U26614 (N_26614,N_25144,N_25117);
and U26615 (N_26615,N_25159,N_25866);
nand U26616 (N_26616,N_25465,N_25446);
and U26617 (N_26617,N_25402,N_25442);
nor U26618 (N_26618,N_25173,N_25036);
or U26619 (N_26619,N_25860,N_25940);
and U26620 (N_26620,N_25475,N_25556);
or U26621 (N_26621,N_25695,N_25204);
xor U26622 (N_26622,N_25964,N_25350);
xnor U26623 (N_26623,N_25259,N_25642);
and U26624 (N_26624,N_25283,N_25275);
xnor U26625 (N_26625,N_25961,N_25462);
nand U26626 (N_26626,N_25401,N_25865);
nand U26627 (N_26627,N_25167,N_25114);
and U26628 (N_26628,N_25415,N_25962);
and U26629 (N_26629,N_25269,N_25042);
nor U26630 (N_26630,N_25209,N_25634);
or U26631 (N_26631,N_25348,N_25230);
or U26632 (N_26632,N_25981,N_25700);
nor U26633 (N_26633,N_25604,N_25798);
xnor U26634 (N_26634,N_25387,N_25262);
nor U26635 (N_26635,N_25749,N_25460);
nor U26636 (N_26636,N_25285,N_25029);
nor U26637 (N_26637,N_25176,N_25983);
xnor U26638 (N_26638,N_25214,N_25710);
and U26639 (N_26639,N_25569,N_25524);
nor U26640 (N_26640,N_25591,N_25070);
or U26641 (N_26641,N_25401,N_25293);
xnor U26642 (N_26642,N_25544,N_25088);
nand U26643 (N_26643,N_25073,N_25659);
nand U26644 (N_26644,N_25485,N_25871);
nand U26645 (N_26645,N_25366,N_25676);
nand U26646 (N_26646,N_25545,N_25099);
or U26647 (N_26647,N_25427,N_25378);
xnor U26648 (N_26648,N_25977,N_25202);
and U26649 (N_26649,N_25693,N_25235);
nand U26650 (N_26650,N_25987,N_25122);
or U26651 (N_26651,N_25699,N_25820);
xnor U26652 (N_26652,N_25197,N_25390);
xor U26653 (N_26653,N_25666,N_25014);
or U26654 (N_26654,N_25637,N_25056);
nand U26655 (N_26655,N_25144,N_25307);
xnor U26656 (N_26656,N_25722,N_25860);
or U26657 (N_26657,N_25205,N_25388);
xnor U26658 (N_26658,N_25780,N_25796);
xnor U26659 (N_26659,N_25403,N_25895);
xor U26660 (N_26660,N_25695,N_25720);
nor U26661 (N_26661,N_25028,N_25556);
nor U26662 (N_26662,N_25471,N_25632);
nand U26663 (N_26663,N_25346,N_25298);
nor U26664 (N_26664,N_25812,N_25818);
or U26665 (N_26665,N_25258,N_25909);
xnor U26666 (N_26666,N_25535,N_25583);
nand U26667 (N_26667,N_25924,N_25880);
or U26668 (N_26668,N_25350,N_25011);
and U26669 (N_26669,N_25552,N_25276);
nand U26670 (N_26670,N_25661,N_25405);
nand U26671 (N_26671,N_25274,N_25327);
and U26672 (N_26672,N_25402,N_25730);
and U26673 (N_26673,N_25668,N_25036);
and U26674 (N_26674,N_25073,N_25656);
nor U26675 (N_26675,N_25240,N_25508);
and U26676 (N_26676,N_25873,N_25537);
xor U26677 (N_26677,N_25345,N_25284);
and U26678 (N_26678,N_25375,N_25168);
nor U26679 (N_26679,N_25474,N_25316);
nor U26680 (N_26680,N_25871,N_25261);
xnor U26681 (N_26681,N_25394,N_25965);
xor U26682 (N_26682,N_25047,N_25020);
nand U26683 (N_26683,N_25495,N_25050);
or U26684 (N_26684,N_25146,N_25056);
nor U26685 (N_26685,N_25072,N_25070);
nand U26686 (N_26686,N_25064,N_25483);
nand U26687 (N_26687,N_25080,N_25390);
or U26688 (N_26688,N_25913,N_25852);
and U26689 (N_26689,N_25614,N_25430);
xor U26690 (N_26690,N_25219,N_25802);
and U26691 (N_26691,N_25036,N_25128);
nand U26692 (N_26692,N_25129,N_25159);
or U26693 (N_26693,N_25668,N_25086);
xor U26694 (N_26694,N_25962,N_25482);
nand U26695 (N_26695,N_25763,N_25875);
xnor U26696 (N_26696,N_25090,N_25890);
or U26697 (N_26697,N_25910,N_25755);
nor U26698 (N_26698,N_25946,N_25844);
and U26699 (N_26699,N_25315,N_25240);
and U26700 (N_26700,N_25168,N_25310);
or U26701 (N_26701,N_25417,N_25519);
or U26702 (N_26702,N_25797,N_25158);
or U26703 (N_26703,N_25255,N_25122);
or U26704 (N_26704,N_25966,N_25825);
nor U26705 (N_26705,N_25702,N_25845);
or U26706 (N_26706,N_25170,N_25545);
nor U26707 (N_26707,N_25244,N_25850);
or U26708 (N_26708,N_25826,N_25652);
nand U26709 (N_26709,N_25873,N_25613);
or U26710 (N_26710,N_25033,N_25972);
nor U26711 (N_26711,N_25188,N_25012);
and U26712 (N_26712,N_25673,N_25677);
xor U26713 (N_26713,N_25829,N_25079);
and U26714 (N_26714,N_25570,N_25411);
nand U26715 (N_26715,N_25912,N_25413);
and U26716 (N_26716,N_25788,N_25179);
xnor U26717 (N_26717,N_25140,N_25066);
or U26718 (N_26718,N_25985,N_25207);
or U26719 (N_26719,N_25427,N_25514);
nand U26720 (N_26720,N_25629,N_25591);
and U26721 (N_26721,N_25253,N_25352);
nor U26722 (N_26722,N_25569,N_25091);
xor U26723 (N_26723,N_25997,N_25200);
or U26724 (N_26724,N_25128,N_25396);
xor U26725 (N_26725,N_25088,N_25279);
or U26726 (N_26726,N_25871,N_25967);
and U26727 (N_26727,N_25485,N_25229);
nand U26728 (N_26728,N_25929,N_25054);
nand U26729 (N_26729,N_25299,N_25393);
xnor U26730 (N_26730,N_25987,N_25026);
and U26731 (N_26731,N_25598,N_25457);
and U26732 (N_26732,N_25957,N_25641);
and U26733 (N_26733,N_25977,N_25314);
and U26734 (N_26734,N_25331,N_25329);
and U26735 (N_26735,N_25105,N_25564);
xor U26736 (N_26736,N_25832,N_25930);
nand U26737 (N_26737,N_25632,N_25369);
nand U26738 (N_26738,N_25724,N_25005);
and U26739 (N_26739,N_25005,N_25088);
nand U26740 (N_26740,N_25540,N_25535);
nor U26741 (N_26741,N_25356,N_25012);
or U26742 (N_26742,N_25487,N_25967);
nor U26743 (N_26743,N_25726,N_25779);
nor U26744 (N_26744,N_25233,N_25235);
xnor U26745 (N_26745,N_25032,N_25043);
or U26746 (N_26746,N_25386,N_25655);
nor U26747 (N_26747,N_25461,N_25796);
and U26748 (N_26748,N_25048,N_25572);
xnor U26749 (N_26749,N_25925,N_25369);
nor U26750 (N_26750,N_25548,N_25294);
nor U26751 (N_26751,N_25568,N_25575);
or U26752 (N_26752,N_25810,N_25441);
and U26753 (N_26753,N_25923,N_25886);
or U26754 (N_26754,N_25217,N_25563);
xnor U26755 (N_26755,N_25888,N_25205);
nand U26756 (N_26756,N_25948,N_25992);
nand U26757 (N_26757,N_25026,N_25980);
or U26758 (N_26758,N_25446,N_25527);
nor U26759 (N_26759,N_25802,N_25731);
nor U26760 (N_26760,N_25549,N_25465);
nor U26761 (N_26761,N_25644,N_25960);
or U26762 (N_26762,N_25069,N_25001);
nor U26763 (N_26763,N_25971,N_25487);
xor U26764 (N_26764,N_25280,N_25870);
and U26765 (N_26765,N_25871,N_25662);
and U26766 (N_26766,N_25709,N_25744);
and U26767 (N_26767,N_25404,N_25287);
and U26768 (N_26768,N_25964,N_25452);
nor U26769 (N_26769,N_25297,N_25045);
nor U26770 (N_26770,N_25192,N_25916);
or U26771 (N_26771,N_25025,N_25887);
nand U26772 (N_26772,N_25364,N_25267);
and U26773 (N_26773,N_25406,N_25206);
xnor U26774 (N_26774,N_25364,N_25385);
or U26775 (N_26775,N_25762,N_25520);
and U26776 (N_26776,N_25988,N_25263);
xor U26777 (N_26777,N_25207,N_25280);
xnor U26778 (N_26778,N_25324,N_25264);
xor U26779 (N_26779,N_25369,N_25668);
xor U26780 (N_26780,N_25865,N_25596);
nand U26781 (N_26781,N_25369,N_25310);
xor U26782 (N_26782,N_25827,N_25413);
xor U26783 (N_26783,N_25668,N_25621);
xnor U26784 (N_26784,N_25915,N_25227);
nand U26785 (N_26785,N_25520,N_25331);
and U26786 (N_26786,N_25676,N_25075);
nor U26787 (N_26787,N_25069,N_25697);
nand U26788 (N_26788,N_25715,N_25698);
nand U26789 (N_26789,N_25481,N_25047);
and U26790 (N_26790,N_25699,N_25971);
nand U26791 (N_26791,N_25317,N_25096);
xor U26792 (N_26792,N_25944,N_25430);
nor U26793 (N_26793,N_25525,N_25271);
nor U26794 (N_26794,N_25723,N_25201);
and U26795 (N_26795,N_25174,N_25602);
or U26796 (N_26796,N_25547,N_25127);
xor U26797 (N_26797,N_25411,N_25263);
nor U26798 (N_26798,N_25027,N_25382);
and U26799 (N_26799,N_25945,N_25791);
xnor U26800 (N_26800,N_25916,N_25233);
and U26801 (N_26801,N_25464,N_25917);
xor U26802 (N_26802,N_25283,N_25515);
nand U26803 (N_26803,N_25200,N_25145);
or U26804 (N_26804,N_25662,N_25546);
nand U26805 (N_26805,N_25022,N_25766);
or U26806 (N_26806,N_25824,N_25638);
nand U26807 (N_26807,N_25442,N_25666);
xnor U26808 (N_26808,N_25515,N_25668);
nor U26809 (N_26809,N_25150,N_25721);
nor U26810 (N_26810,N_25613,N_25573);
xnor U26811 (N_26811,N_25966,N_25557);
or U26812 (N_26812,N_25739,N_25416);
xor U26813 (N_26813,N_25592,N_25107);
and U26814 (N_26814,N_25881,N_25904);
nand U26815 (N_26815,N_25050,N_25311);
nand U26816 (N_26816,N_25039,N_25235);
nor U26817 (N_26817,N_25620,N_25133);
nand U26818 (N_26818,N_25378,N_25452);
nor U26819 (N_26819,N_25773,N_25236);
or U26820 (N_26820,N_25444,N_25017);
xor U26821 (N_26821,N_25542,N_25849);
and U26822 (N_26822,N_25381,N_25220);
xnor U26823 (N_26823,N_25409,N_25428);
nand U26824 (N_26824,N_25582,N_25354);
and U26825 (N_26825,N_25782,N_25171);
xor U26826 (N_26826,N_25028,N_25249);
or U26827 (N_26827,N_25839,N_25636);
or U26828 (N_26828,N_25315,N_25117);
and U26829 (N_26829,N_25883,N_25526);
and U26830 (N_26830,N_25327,N_25070);
nor U26831 (N_26831,N_25400,N_25987);
nand U26832 (N_26832,N_25352,N_25554);
nand U26833 (N_26833,N_25650,N_25561);
or U26834 (N_26834,N_25405,N_25625);
and U26835 (N_26835,N_25560,N_25875);
xor U26836 (N_26836,N_25882,N_25312);
and U26837 (N_26837,N_25575,N_25148);
xor U26838 (N_26838,N_25721,N_25771);
and U26839 (N_26839,N_25738,N_25713);
nand U26840 (N_26840,N_25163,N_25191);
or U26841 (N_26841,N_25092,N_25146);
xnor U26842 (N_26842,N_25392,N_25016);
or U26843 (N_26843,N_25390,N_25607);
nand U26844 (N_26844,N_25766,N_25191);
nor U26845 (N_26845,N_25200,N_25339);
and U26846 (N_26846,N_25810,N_25857);
xnor U26847 (N_26847,N_25454,N_25513);
xnor U26848 (N_26848,N_25029,N_25268);
nand U26849 (N_26849,N_25556,N_25212);
xor U26850 (N_26850,N_25362,N_25173);
nor U26851 (N_26851,N_25123,N_25344);
or U26852 (N_26852,N_25925,N_25240);
and U26853 (N_26853,N_25682,N_25433);
and U26854 (N_26854,N_25661,N_25434);
nor U26855 (N_26855,N_25998,N_25524);
or U26856 (N_26856,N_25324,N_25695);
xnor U26857 (N_26857,N_25365,N_25412);
nor U26858 (N_26858,N_25530,N_25315);
and U26859 (N_26859,N_25023,N_25116);
nand U26860 (N_26860,N_25428,N_25856);
or U26861 (N_26861,N_25513,N_25064);
nor U26862 (N_26862,N_25681,N_25416);
nor U26863 (N_26863,N_25110,N_25469);
or U26864 (N_26864,N_25082,N_25576);
nor U26865 (N_26865,N_25156,N_25897);
or U26866 (N_26866,N_25068,N_25227);
nor U26867 (N_26867,N_25716,N_25942);
or U26868 (N_26868,N_25261,N_25496);
nor U26869 (N_26869,N_25434,N_25190);
xnor U26870 (N_26870,N_25146,N_25253);
or U26871 (N_26871,N_25908,N_25122);
nand U26872 (N_26872,N_25341,N_25834);
nor U26873 (N_26873,N_25634,N_25533);
nand U26874 (N_26874,N_25137,N_25687);
nand U26875 (N_26875,N_25689,N_25648);
nand U26876 (N_26876,N_25539,N_25893);
and U26877 (N_26877,N_25586,N_25799);
nand U26878 (N_26878,N_25662,N_25622);
and U26879 (N_26879,N_25070,N_25206);
and U26880 (N_26880,N_25264,N_25680);
nand U26881 (N_26881,N_25943,N_25522);
nor U26882 (N_26882,N_25960,N_25305);
nor U26883 (N_26883,N_25587,N_25501);
xnor U26884 (N_26884,N_25418,N_25976);
nor U26885 (N_26885,N_25424,N_25906);
or U26886 (N_26886,N_25756,N_25724);
nand U26887 (N_26887,N_25192,N_25512);
and U26888 (N_26888,N_25067,N_25335);
and U26889 (N_26889,N_25900,N_25695);
or U26890 (N_26890,N_25055,N_25947);
or U26891 (N_26891,N_25162,N_25967);
nor U26892 (N_26892,N_25821,N_25980);
nand U26893 (N_26893,N_25554,N_25623);
nor U26894 (N_26894,N_25899,N_25957);
nor U26895 (N_26895,N_25287,N_25839);
or U26896 (N_26896,N_25201,N_25465);
nor U26897 (N_26897,N_25065,N_25645);
nor U26898 (N_26898,N_25862,N_25660);
nand U26899 (N_26899,N_25829,N_25442);
nand U26900 (N_26900,N_25979,N_25413);
and U26901 (N_26901,N_25533,N_25566);
nand U26902 (N_26902,N_25187,N_25180);
nand U26903 (N_26903,N_25079,N_25062);
nand U26904 (N_26904,N_25898,N_25016);
nor U26905 (N_26905,N_25292,N_25120);
nand U26906 (N_26906,N_25490,N_25510);
nand U26907 (N_26907,N_25416,N_25861);
and U26908 (N_26908,N_25373,N_25144);
and U26909 (N_26909,N_25215,N_25856);
or U26910 (N_26910,N_25916,N_25784);
and U26911 (N_26911,N_25366,N_25410);
xor U26912 (N_26912,N_25849,N_25845);
nor U26913 (N_26913,N_25430,N_25969);
nand U26914 (N_26914,N_25301,N_25860);
nor U26915 (N_26915,N_25323,N_25894);
or U26916 (N_26916,N_25118,N_25590);
xor U26917 (N_26917,N_25904,N_25380);
nor U26918 (N_26918,N_25413,N_25138);
nor U26919 (N_26919,N_25045,N_25741);
xnor U26920 (N_26920,N_25213,N_25260);
nor U26921 (N_26921,N_25228,N_25443);
and U26922 (N_26922,N_25602,N_25046);
or U26923 (N_26923,N_25327,N_25818);
or U26924 (N_26924,N_25156,N_25193);
nand U26925 (N_26925,N_25007,N_25161);
and U26926 (N_26926,N_25224,N_25831);
nand U26927 (N_26927,N_25560,N_25791);
nor U26928 (N_26928,N_25212,N_25767);
or U26929 (N_26929,N_25992,N_25381);
nor U26930 (N_26930,N_25745,N_25959);
nor U26931 (N_26931,N_25331,N_25199);
xnor U26932 (N_26932,N_25862,N_25785);
xnor U26933 (N_26933,N_25250,N_25824);
or U26934 (N_26934,N_25243,N_25879);
nand U26935 (N_26935,N_25303,N_25044);
nand U26936 (N_26936,N_25536,N_25972);
or U26937 (N_26937,N_25812,N_25719);
xnor U26938 (N_26938,N_25009,N_25848);
and U26939 (N_26939,N_25195,N_25802);
and U26940 (N_26940,N_25630,N_25510);
nand U26941 (N_26941,N_25452,N_25310);
or U26942 (N_26942,N_25256,N_25172);
or U26943 (N_26943,N_25171,N_25824);
xnor U26944 (N_26944,N_25139,N_25545);
or U26945 (N_26945,N_25311,N_25599);
or U26946 (N_26946,N_25575,N_25415);
and U26947 (N_26947,N_25739,N_25451);
nand U26948 (N_26948,N_25441,N_25525);
nand U26949 (N_26949,N_25779,N_25962);
nor U26950 (N_26950,N_25774,N_25492);
nand U26951 (N_26951,N_25343,N_25150);
and U26952 (N_26952,N_25389,N_25215);
or U26953 (N_26953,N_25808,N_25865);
nand U26954 (N_26954,N_25906,N_25684);
or U26955 (N_26955,N_25314,N_25843);
nand U26956 (N_26956,N_25133,N_25863);
xor U26957 (N_26957,N_25042,N_25584);
xnor U26958 (N_26958,N_25126,N_25063);
and U26959 (N_26959,N_25301,N_25812);
and U26960 (N_26960,N_25925,N_25342);
or U26961 (N_26961,N_25506,N_25219);
nor U26962 (N_26962,N_25957,N_25988);
and U26963 (N_26963,N_25724,N_25888);
nand U26964 (N_26964,N_25931,N_25284);
xor U26965 (N_26965,N_25849,N_25639);
nor U26966 (N_26966,N_25869,N_25028);
xor U26967 (N_26967,N_25764,N_25702);
nand U26968 (N_26968,N_25434,N_25811);
nand U26969 (N_26969,N_25179,N_25932);
nand U26970 (N_26970,N_25885,N_25610);
xnor U26971 (N_26971,N_25691,N_25911);
and U26972 (N_26972,N_25218,N_25861);
nor U26973 (N_26973,N_25178,N_25896);
nor U26974 (N_26974,N_25678,N_25148);
nand U26975 (N_26975,N_25069,N_25302);
or U26976 (N_26976,N_25488,N_25272);
nor U26977 (N_26977,N_25842,N_25802);
nand U26978 (N_26978,N_25711,N_25442);
nor U26979 (N_26979,N_25975,N_25452);
xor U26980 (N_26980,N_25298,N_25279);
or U26981 (N_26981,N_25463,N_25867);
xor U26982 (N_26982,N_25973,N_25668);
xnor U26983 (N_26983,N_25982,N_25232);
and U26984 (N_26984,N_25867,N_25406);
or U26985 (N_26985,N_25402,N_25707);
or U26986 (N_26986,N_25598,N_25539);
nand U26987 (N_26987,N_25666,N_25717);
or U26988 (N_26988,N_25074,N_25198);
nand U26989 (N_26989,N_25582,N_25956);
or U26990 (N_26990,N_25972,N_25477);
xnor U26991 (N_26991,N_25954,N_25040);
nor U26992 (N_26992,N_25865,N_25895);
nor U26993 (N_26993,N_25645,N_25907);
and U26994 (N_26994,N_25074,N_25542);
and U26995 (N_26995,N_25384,N_25241);
xnor U26996 (N_26996,N_25734,N_25096);
nand U26997 (N_26997,N_25399,N_25207);
or U26998 (N_26998,N_25423,N_25752);
and U26999 (N_26999,N_25960,N_25870);
nor U27000 (N_27000,N_26341,N_26760);
and U27001 (N_27001,N_26369,N_26506);
nand U27002 (N_27002,N_26105,N_26025);
nor U27003 (N_27003,N_26168,N_26792);
nor U27004 (N_27004,N_26597,N_26040);
or U27005 (N_27005,N_26729,N_26265);
nand U27006 (N_27006,N_26741,N_26733);
and U27007 (N_27007,N_26171,N_26237);
nand U27008 (N_27008,N_26344,N_26063);
nor U27009 (N_27009,N_26103,N_26348);
nor U27010 (N_27010,N_26579,N_26130);
and U27011 (N_27011,N_26921,N_26926);
or U27012 (N_27012,N_26319,N_26032);
xor U27013 (N_27013,N_26007,N_26363);
nand U27014 (N_27014,N_26997,N_26540);
nand U27015 (N_27015,N_26084,N_26659);
and U27016 (N_27016,N_26952,N_26875);
nor U27017 (N_27017,N_26093,N_26894);
or U27018 (N_27018,N_26799,N_26927);
nand U27019 (N_27019,N_26351,N_26727);
or U27020 (N_27020,N_26177,N_26527);
nor U27021 (N_27021,N_26394,N_26607);
xnor U27022 (N_27022,N_26408,N_26212);
and U27023 (N_27023,N_26648,N_26384);
and U27024 (N_27024,N_26305,N_26944);
xor U27025 (N_27025,N_26091,N_26210);
nor U27026 (N_27026,N_26877,N_26737);
xnor U27027 (N_27027,N_26698,N_26477);
nand U27028 (N_27028,N_26950,N_26514);
and U27029 (N_27029,N_26669,N_26656);
nand U27030 (N_27030,N_26757,N_26021);
nor U27031 (N_27031,N_26419,N_26249);
nand U27032 (N_27032,N_26423,N_26629);
xnor U27033 (N_27033,N_26273,N_26189);
xor U27034 (N_27034,N_26452,N_26417);
nor U27035 (N_27035,N_26936,N_26484);
nor U27036 (N_27036,N_26414,N_26404);
xor U27037 (N_27037,N_26738,N_26876);
or U27038 (N_27038,N_26705,N_26052);
xor U27039 (N_27039,N_26548,N_26769);
nor U27040 (N_27040,N_26914,N_26957);
and U27041 (N_27041,N_26571,N_26498);
xor U27042 (N_27042,N_26697,N_26780);
or U27043 (N_27043,N_26288,N_26614);
xnor U27044 (N_27044,N_26541,N_26897);
nand U27045 (N_27045,N_26572,N_26263);
and U27046 (N_27046,N_26128,N_26524);
nand U27047 (N_27047,N_26062,N_26368);
nor U27048 (N_27048,N_26984,N_26012);
nand U27049 (N_27049,N_26179,N_26181);
and U27050 (N_27050,N_26829,N_26674);
nand U27051 (N_27051,N_26577,N_26213);
nor U27052 (N_27052,N_26662,N_26018);
and U27053 (N_27053,N_26990,N_26569);
or U27054 (N_27054,N_26775,N_26359);
nand U27055 (N_27055,N_26497,N_26592);
xnor U27056 (N_27056,N_26334,N_26898);
or U27057 (N_27057,N_26071,N_26338);
and U27058 (N_27058,N_26753,N_26901);
or U27059 (N_27059,N_26557,N_26186);
or U27060 (N_27060,N_26896,N_26630);
and U27061 (N_27061,N_26616,N_26217);
nor U27062 (N_27062,N_26904,N_26440);
xor U27063 (N_27063,N_26617,N_26050);
nor U27064 (N_27064,N_26061,N_26429);
and U27065 (N_27065,N_26045,N_26689);
or U27066 (N_27066,N_26406,N_26499);
and U27067 (N_27067,N_26204,N_26343);
nor U27068 (N_27068,N_26717,N_26401);
and U27069 (N_27069,N_26768,N_26468);
and U27070 (N_27070,N_26488,N_26231);
or U27071 (N_27071,N_26112,N_26388);
nand U27072 (N_27072,N_26542,N_26123);
nand U27073 (N_27073,N_26358,N_26730);
nand U27074 (N_27074,N_26519,N_26657);
or U27075 (N_27075,N_26076,N_26395);
nand U27076 (N_27076,N_26166,N_26236);
and U27077 (N_27077,N_26507,N_26838);
and U27078 (N_27078,N_26908,N_26449);
xor U27079 (N_27079,N_26244,N_26126);
and U27080 (N_27080,N_26972,N_26042);
nor U27081 (N_27081,N_26392,N_26596);
xnor U27082 (N_27082,N_26871,N_26975);
and U27083 (N_27083,N_26794,N_26664);
or U27084 (N_27084,N_26378,N_26276);
nand U27085 (N_27085,N_26354,N_26841);
xnor U27086 (N_27086,N_26307,N_26810);
xnor U27087 (N_27087,N_26203,N_26136);
nand U27088 (N_27088,N_26391,N_26795);
nor U27089 (N_27089,N_26887,N_26919);
or U27090 (N_27090,N_26880,N_26459);
nand U27091 (N_27091,N_26330,N_26081);
and U27092 (N_27092,N_26293,N_26781);
or U27093 (N_27093,N_26773,N_26325);
and U27094 (N_27094,N_26470,N_26458);
xnor U27095 (N_27095,N_26732,N_26655);
nor U27096 (N_27096,N_26986,N_26530);
or U27097 (N_27097,N_26056,N_26644);
and U27098 (N_27098,N_26409,N_26886);
and U27099 (N_27099,N_26329,N_26779);
nand U27100 (N_27100,N_26920,N_26554);
xor U27101 (N_27101,N_26934,N_26869);
or U27102 (N_27102,N_26874,N_26397);
nand U27103 (N_27103,N_26024,N_26182);
nor U27104 (N_27104,N_26937,N_26114);
or U27105 (N_27105,N_26744,N_26367);
nand U27106 (N_27106,N_26620,N_26653);
and U27107 (N_27107,N_26627,N_26218);
xor U27108 (N_27108,N_26190,N_26254);
nor U27109 (N_27109,N_26808,N_26745);
nand U27110 (N_27110,N_26782,N_26193);
or U27111 (N_27111,N_26016,N_26820);
nand U27112 (N_27112,N_26313,N_26039);
xnor U27113 (N_27113,N_26512,N_26537);
xnor U27114 (N_27114,N_26603,N_26743);
nand U27115 (N_27115,N_26930,N_26543);
nand U27116 (N_27116,N_26508,N_26583);
and U27117 (N_27117,N_26684,N_26115);
nand U27118 (N_27118,N_26762,N_26977);
and U27119 (N_27119,N_26376,N_26366);
nor U27120 (N_27120,N_26108,N_26312);
nand U27121 (N_27121,N_26800,N_26591);
xnor U27122 (N_27122,N_26173,N_26723);
and U27123 (N_27123,N_26188,N_26558);
xnor U27124 (N_27124,N_26422,N_26899);
and U27125 (N_27125,N_26523,N_26194);
nand U27126 (N_27126,N_26030,N_26710);
and U27127 (N_27127,N_26615,N_26197);
or U27128 (N_27128,N_26666,N_26682);
nor U27129 (N_27129,N_26260,N_26353);
nand U27130 (N_27130,N_26259,N_26839);
and U27131 (N_27131,N_26308,N_26846);
or U27132 (N_27132,N_26234,N_26503);
or U27133 (N_27133,N_26481,N_26547);
xnor U27134 (N_27134,N_26298,N_26584);
nand U27135 (N_27135,N_26885,N_26825);
or U27136 (N_27136,N_26278,N_26362);
and U27137 (N_27137,N_26604,N_26865);
and U27138 (N_27138,N_26702,N_26501);
xnor U27139 (N_27139,N_26335,N_26479);
xnor U27140 (N_27140,N_26055,N_26457);
nor U27141 (N_27141,N_26106,N_26700);
and U27142 (N_27142,N_26001,N_26529);
xnor U27143 (N_27143,N_26824,N_26725);
and U27144 (N_27144,N_26285,N_26574);
or U27145 (N_27145,N_26955,N_26412);
nand U27146 (N_27146,N_26639,N_26478);
xnor U27147 (N_27147,N_26559,N_26491);
or U27148 (N_27148,N_26500,N_26783);
nor U27149 (N_27149,N_26834,N_26538);
nand U27150 (N_27150,N_26752,N_26451);
nor U27151 (N_27151,N_26631,N_26502);
nor U27152 (N_27152,N_26649,N_26987);
xor U27153 (N_27153,N_26555,N_26157);
or U27154 (N_27154,N_26946,N_26686);
nor U27155 (N_27155,N_26706,N_26881);
nand U27156 (N_27156,N_26956,N_26010);
and U27157 (N_27157,N_26742,N_26318);
nor U27158 (N_27158,N_26301,N_26690);
or U27159 (N_27159,N_26437,N_26192);
or U27160 (N_27160,N_26640,N_26372);
or U27161 (N_27161,N_26153,N_26772);
nand U27162 (N_27162,N_26601,N_26916);
nor U27163 (N_27163,N_26033,N_26801);
nor U27164 (N_27164,N_26836,N_26228);
or U27165 (N_27165,N_26465,N_26685);
xnor U27166 (N_27166,N_26043,N_26731);
xnor U27167 (N_27167,N_26389,N_26968);
or U27168 (N_27168,N_26870,N_26096);
xor U27169 (N_27169,N_26515,N_26804);
xor U27170 (N_27170,N_26954,N_26890);
or U27171 (N_27171,N_26859,N_26867);
and U27172 (N_27172,N_26152,N_26147);
nor U27173 (N_27173,N_26207,N_26077);
nand U27174 (N_27174,N_26943,N_26020);
nand U27175 (N_27175,N_26421,N_26945);
or U27176 (N_27176,N_26361,N_26940);
and U27177 (N_27177,N_26856,N_26080);
or U27178 (N_27178,N_26905,N_26645);
or U27179 (N_27179,N_26211,N_26480);
nor U27180 (N_27180,N_26059,N_26658);
xor U27181 (N_27181,N_26332,N_26066);
nand U27182 (N_27182,N_26694,N_26712);
nand U27183 (N_27183,N_26903,N_26140);
and U27184 (N_27184,N_26942,N_26120);
and U27185 (N_27185,N_26552,N_26400);
or U27186 (N_27186,N_26974,N_26195);
nand U27187 (N_27187,N_26239,N_26430);
or U27188 (N_27188,N_26766,N_26067);
or U27189 (N_27189,N_26017,N_26970);
or U27190 (N_27190,N_26340,N_26879);
nor U27191 (N_27191,N_26746,N_26525);
xnor U27192 (N_27192,N_26843,N_26761);
or U27193 (N_27193,N_26988,N_26602);
xnor U27194 (N_27194,N_26352,N_26082);
xnor U27195 (N_27195,N_26910,N_26089);
or U27196 (N_27196,N_26411,N_26835);
xor U27197 (N_27197,N_26551,N_26665);
nand U27198 (N_27198,N_26013,N_26981);
or U27199 (N_27199,N_26214,N_26982);
xor U27200 (N_27200,N_26466,N_26979);
nor U27201 (N_27201,N_26815,N_26420);
nand U27202 (N_27202,N_26156,N_26283);
or U27203 (N_27203,N_26822,N_26961);
nor U27204 (N_27204,N_26976,N_26224);
or U27205 (N_27205,N_26439,N_26492);
and U27206 (N_27206,N_26405,N_26814);
nand U27207 (N_27207,N_26661,N_26118);
and U27208 (N_27208,N_26246,N_26200);
and U27209 (N_27209,N_26842,N_26959);
nand U27210 (N_27210,N_26300,N_26410);
and U27211 (N_27211,N_26011,N_26504);
xor U27212 (N_27212,N_26832,N_26037);
and U27213 (N_27213,N_26159,N_26763);
and U27214 (N_27214,N_26522,N_26403);
nor U27215 (N_27215,N_26594,N_26688);
xnor U27216 (N_27216,N_26337,N_26994);
nor U27217 (N_27217,N_26670,N_26187);
nor U27218 (N_27218,N_26111,N_26549);
nor U27219 (N_27219,N_26754,N_26446);
nor U27220 (N_27220,N_26432,N_26315);
nand U27221 (N_27221,N_26888,N_26912);
nor U27222 (N_27222,N_26964,N_26223);
nor U27223 (N_27223,N_26023,N_26280);
nand U27224 (N_27224,N_26535,N_26428);
and U27225 (N_27225,N_26269,N_26328);
xor U27226 (N_27226,N_26238,N_26232);
nand U27227 (N_27227,N_26216,N_26855);
nor U27228 (N_27228,N_26463,N_26333);
or U27229 (N_27229,N_26486,N_26078);
nand U27230 (N_27230,N_26336,N_26845);
or U27231 (N_27231,N_26438,N_26626);
nor U27232 (N_27232,N_26349,N_26100);
xor U27233 (N_27233,N_26651,N_26509);
nor U27234 (N_27234,N_26643,N_26893);
nand U27235 (N_27235,N_26296,N_26844);
xor U27236 (N_27236,N_26819,N_26787);
nand U27237 (N_27237,N_26948,N_26487);
nand U27238 (N_27238,N_26104,N_26131);
or U27239 (N_27239,N_26711,N_26471);
nand U27240 (N_27240,N_26146,N_26826);
nand U27241 (N_27241,N_26483,N_26241);
nand U27242 (N_27242,N_26749,N_26517);
nor U27243 (N_27243,N_26386,N_26590);
xnor U27244 (N_27244,N_26811,N_26510);
nor U27245 (N_27245,N_26637,N_26208);
or U27246 (N_27246,N_26314,N_26545);
nor U27247 (N_27247,N_26321,N_26381);
nor U27248 (N_27248,N_26132,N_26174);
nand U27249 (N_27249,N_26015,N_26185);
and U27250 (N_27250,N_26550,N_26713);
and U27251 (N_27251,N_26793,N_26461);
xnor U27252 (N_27252,N_26747,N_26048);
nor U27253 (N_27253,N_26274,N_26947);
xnor U27254 (N_27254,N_26693,N_26802);
nand U27255 (N_27255,N_26135,N_26691);
and U27256 (N_27256,N_26133,N_26632);
and U27257 (N_27257,N_26206,N_26014);
nor U27258 (N_27258,N_26180,N_26191);
and U27259 (N_27259,N_26247,N_26764);
nand U27260 (N_27260,N_26673,N_26539);
xor U27261 (N_27261,N_26911,N_26331);
nor U27262 (N_27262,N_26567,N_26287);
or U27263 (N_27263,N_26447,N_26472);
nand U27264 (N_27264,N_26728,N_26528);
xor U27265 (N_27265,N_26143,N_26074);
or U27266 (N_27266,N_26939,N_26310);
xor U27267 (N_27267,N_26692,N_26427);
and U27268 (N_27268,N_26083,N_26242);
or U27269 (N_27269,N_26003,N_26935);
or U27270 (N_27270,N_26812,N_26272);
and U27271 (N_27271,N_26041,N_26004);
nand U27272 (N_27272,N_26586,N_26612);
nor U27273 (N_27273,N_26065,N_26064);
and U27274 (N_27274,N_26292,N_26380);
or U27275 (N_27275,N_26474,N_26364);
or U27276 (N_27276,N_26460,N_26060);
nor U27277 (N_27277,N_26714,N_26606);
nor U27278 (N_27278,N_26489,N_26960);
xnor U27279 (N_27279,N_26165,N_26668);
nor U27280 (N_27280,N_26683,N_26789);
nand U27281 (N_27281,N_26892,N_26144);
nand U27282 (N_27282,N_26496,N_26605);
xnor U27283 (N_27283,N_26306,N_26161);
nor U27284 (N_27284,N_26813,N_26075);
xor U27285 (N_27285,N_26791,N_26137);
nand U27286 (N_27286,N_26291,N_26220);
nor U27287 (N_27287,N_26513,N_26008);
nand U27288 (N_27288,N_26676,N_26347);
nor U27289 (N_27289,N_26243,N_26134);
or U27290 (N_27290,N_26719,N_26357);
and U27291 (N_27291,N_26758,N_26070);
nor U27292 (N_27292,N_26734,N_26121);
and U27293 (N_27293,N_26124,N_26383);
nand U27294 (N_27294,N_26847,N_26275);
nor U27295 (N_27295,N_26476,N_26613);
and U27296 (N_27296,N_26122,N_26784);
nand U27297 (N_27297,N_26739,N_26151);
nand U27298 (N_27298,N_26374,N_26323);
or U27299 (N_27299,N_26294,N_26989);
or U27300 (N_27300,N_26917,N_26178);
nor U27301 (N_27301,N_26467,N_26360);
or U27302 (N_27302,N_26086,N_26909);
nor U27303 (N_27303,N_26924,N_26227);
nand U27304 (N_27304,N_26895,N_26932);
xnor U27305 (N_27305,N_26371,N_26026);
xnor U27306 (N_27306,N_26495,N_26805);
nand U27307 (N_27307,N_26407,N_26915);
nand U27308 (N_27308,N_26953,N_26176);
nor U27309 (N_27309,N_26051,N_26533);
nand U27310 (N_27310,N_26303,N_26991);
or U27311 (N_27311,N_26473,N_26046);
xor U27312 (N_27312,N_26054,N_26038);
or U27313 (N_27313,N_26767,N_26951);
nor U27314 (N_27314,N_26235,N_26145);
nor U27315 (N_27315,N_26490,N_26866);
nand U27316 (N_27316,N_26980,N_26005);
and U27317 (N_27317,N_26258,N_26563);
or U27318 (N_27318,N_26324,N_26240);
or U27319 (N_27319,N_26588,N_26677);
or U27320 (N_27320,N_26493,N_26261);
nor U27321 (N_27321,N_26598,N_26327);
or U27322 (N_27322,N_26028,N_26776);
xnor U27323 (N_27323,N_26277,N_26678);
xnor U27324 (N_27324,N_26183,N_26701);
xor U27325 (N_27325,N_26009,N_26069);
and U27326 (N_27326,N_26628,N_26141);
xor U27327 (N_27327,N_26289,N_26851);
nor U27328 (N_27328,N_26850,N_26262);
nor U27329 (N_27329,N_26393,N_26993);
or U27330 (N_27330,N_26636,N_26219);
or U27331 (N_27331,N_26965,N_26848);
and U27332 (N_27332,N_26907,N_26933);
xor U27333 (N_27333,N_26209,N_26454);
or U27334 (N_27334,N_26582,N_26229);
nor U27335 (N_27335,N_26169,N_26095);
xor U27336 (N_27336,N_26175,N_26110);
nor U27337 (N_27337,N_26778,N_26671);
and U27338 (N_27338,N_26827,N_26650);
nand U27339 (N_27339,N_26770,N_26862);
and U27340 (N_27340,N_26906,N_26771);
xnor U27341 (N_27341,N_26425,N_26350);
nand U27342 (N_27342,N_26828,N_26355);
nor U27343 (N_27343,N_26608,N_26382);
nand U27344 (N_27344,N_26652,N_26356);
nand U27345 (N_27345,N_26370,N_26849);
or U27346 (N_27346,N_26647,N_26049);
and U27347 (N_27347,N_26575,N_26225);
or U27348 (N_27348,N_26599,N_26149);
or U27349 (N_27349,N_26581,N_26565);
or U27350 (N_27350,N_26585,N_26019);
xnor U27351 (N_27351,N_26090,N_26823);
nor U27352 (N_27352,N_26047,N_26999);
or U27353 (N_27353,N_26087,N_26268);
nand U27354 (N_27354,N_26044,N_26675);
nor U27355 (N_27355,N_26142,N_26162);
nand U27356 (N_27356,N_26863,N_26002);
nand U27357 (N_27357,N_26923,N_26101);
nand U27358 (N_27358,N_26623,N_26546);
or U27359 (N_27359,N_26079,N_26873);
and U27360 (N_27360,N_26797,N_26088);
nand U27361 (N_27361,N_26184,N_26922);
or U27362 (N_27362,N_26456,N_26736);
nand U27363 (N_27363,N_26129,N_26816);
nand U27364 (N_27364,N_26469,N_26304);
xnor U27365 (N_27365,N_26872,N_26316);
nand U27366 (N_27366,N_26696,N_26297);
and U27367 (N_27367,N_26938,N_26595);
nor U27368 (N_27368,N_26704,N_26611);
or U27369 (N_27369,N_26482,N_26443);
or U27370 (N_27370,N_26092,N_26672);
or U27371 (N_27371,N_26610,N_26929);
or U27372 (N_27372,N_26751,N_26619);
and U27373 (N_27373,N_26570,N_26703);
nor U27374 (N_27374,N_26663,N_26807);
nand U27375 (N_27375,N_26416,N_26634);
or U27376 (N_27376,N_26155,N_26415);
nand U27377 (N_27377,N_26852,N_26726);
or U27378 (N_27378,N_26777,N_26036);
nand U27379 (N_27379,N_26442,N_26435);
or U27380 (N_27380,N_26464,N_26450);
nor U27381 (N_27381,N_26695,N_26164);
nand U27382 (N_27382,N_26000,N_26320);
nand U27383 (N_27383,N_26996,N_26282);
and U27384 (N_27384,N_26568,N_26638);
or U27385 (N_27385,N_26853,N_26266);
nor U27386 (N_27386,N_26593,N_26109);
xor U27387 (N_27387,N_26399,N_26167);
nand U27388 (N_27388,N_26803,N_26034);
nor U27389 (N_27389,N_26475,N_26505);
or U27390 (N_27390,N_26854,N_26098);
nand U27391 (N_27391,N_26600,N_26715);
or U27392 (N_27392,N_26969,N_26646);
and U27393 (N_27393,N_26431,N_26365);
nor U27394 (N_27394,N_26253,N_26798);
and U27395 (N_27395,N_26958,N_26564);
or U27396 (N_27396,N_26099,N_26221);
nand U27397 (N_27397,N_26884,N_26967);
nand U27398 (N_27398,N_26271,N_26245);
nand U27399 (N_27399,N_26750,N_26840);
nand U27400 (N_27400,N_26441,N_26281);
nor U27401 (N_27401,N_26113,N_26641);
or U27402 (N_27402,N_26127,N_26963);
xor U27403 (N_27403,N_26154,N_26150);
nand U27404 (N_27404,N_26622,N_26251);
nand U27405 (N_27405,N_26837,N_26821);
and U27406 (N_27406,N_26027,N_26448);
nor U27407 (N_27407,N_26279,N_26818);
xor U27408 (N_27408,N_26196,N_26444);
and U27409 (N_27409,N_26326,N_26573);
and U27410 (N_27410,N_26660,N_26735);
or U27411 (N_27411,N_26436,N_26198);
or U27412 (N_27412,N_26716,N_26889);
nand U27413 (N_27413,N_26566,N_26205);
and U27414 (N_27414,N_26256,N_26925);
or U27415 (N_27415,N_26809,N_26831);
nand U27416 (N_27416,N_26992,N_26708);
or U27417 (N_27417,N_26724,N_26817);
nor U27418 (N_27418,N_26973,N_26788);
and U27419 (N_27419,N_26578,N_26345);
nor U27420 (N_27420,N_26534,N_26759);
nand U27421 (N_27421,N_26531,N_26526);
or U27422 (N_27422,N_26707,N_26721);
xnor U27423 (N_27423,N_26290,N_26830);
xnor U27424 (N_27424,N_26913,N_26158);
and U27425 (N_27425,N_26295,N_26445);
and U27426 (N_27426,N_26576,N_26765);
and U27427 (N_27427,N_26796,N_26006);
nand U27428 (N_27428,N_26299,N_26536);
or U27429 (N_27429,N_26931,N_26250);
and U27430 (N_27430,N_26097,N_26978);
nand U27431 (N_27431,N_26373,N_26868);
or U27432 (N_27432,N_26962,N_26561);
xor U27433 (N_27433,N_26681,N_26941);
or U27434 (N_27434,N_26201,N_26317);
xnor U27435 (N_27435,N_26094,N_26139);
and U27436 (N_27436,N_26125,N_26532);
nand U27437 (N_27437,N_26398,N_26022);
nand U27438 (N_27438,N_26857,N_26068);
xnor U27439 (N_27439,N_26433,N_26774);
nor U27440 (N_27440,N_26621,N_26485);
or U27441 (N_27441,N_26058,N_26160);
xnor U27442 (N_27442,N_26518,N_26864);
or U27443 (N_27443,N_26107,N_26971);
xor U27444 (N_27444,N_26722,N_26635);
or U27445 (N_27445,N_26402,N_26709);
xnor U27446 (N_27446,N_26396,N_26858);
xor U27447 (N_27447,N_26424,N_26560);
nand U27448 (N_27448,N_26138,N_26654);
or U27449 (N_27449,N_26053,N_26453);
xnor U27450 (N_27450,N_26587,N_26462);
nor U27451 (N_27451,N_26642,N_26516);
or U27452 (N_27452,N_26117,N_26878);
nor U27453 (N_27453,N_26248,N_26589);
xor U27454 (N_27454,N_26385,N_26035);
nor U27455 (N_27455,N_26346,N_26085);
nand U27456 (N_27456,N_26199,N_26494);
nor U27457 (N_27457,N_26609,N_26072);
nor U27458 (N_27458,N_26342,N_26222);
or U27459 (N_27459,N_26520,N_26387);
nor U27460 (N_27460,N_26233,N_26434);
or U27461 (N_27461,N_26902,N_26928);
and U27462 (N_27462,N_26891,N_26861);
xor U27463 (N_27463,N_26580,N_26995);
nor U27464 (N_27464,N_26170,N_26679);
or U27465 (N_27465,N_26748,N_26720);
nand U27466 (N_27466,N_26264,N_26029);
and U27467 (N_27467,N_26102,N_26882);
nor U27468 (N_27468,N_26116,N_26311);
nand U27469 (N_27469,N_26918,N_26163);
xnor U27470 (N_27470,N_26966,N_26284);
xor U27471 (N_27471,N_26562,N_26379);
xor U27472 (N_27472,N_26949,N_26756);
xor U27473 (N_27473,N_26833,N_26618);
and U27474 (N_27474,N_26148,N_26302);
nand U27475 (N_27475,N_26860,N_26544);
xnor U27476 (N_27476,N_26286,N_26985);
nand U27477 (N_27477,N_26309,N_26699);
nand U27478 (N_27478,N_26339,N_26983);
nor U27479 (N_27479,N_26267,N_26553);
nor U27480 (N_27480,N_26073,N_26031);
or U27481 (N_27481,N_26390,N_26900);
nor U27482 (N_27482,N_26680,N_26215);
nor U27483 (N_27483,N_26687,N_26270);
or U27484 (N_27484,N_26455,N_26377);
xnor U27485 (N_27485,N_26556,N_26521);
nand U27486 (N_27486,N_26375,N_26625);
nor U27487 (N_27487,N_26226,N_26119);
nand U27488 (N_27488,N_26257,N_26667);
xor U27489 (N_27489,N_26511,N_26322);
nand U27490 (N_27490,N_26806,N_26252);
or U27491 (N_27491,N_26230,N_26998);
nand U27492 (N_27492,N_26413,N_26790);
and U27493 (N_27493,N_26624,N_26883);
nand U27494 (N_27494,N_26202,N_26057);
nor U27495 (N_27495,N_26426,N_26755);
nor U27496 (N_27496,N_26172,N_26785);
nor U27497 (N_27497,N_26633,N_26740);
and U27498 (N_27498,N_26255,N_26786);
nor U27499 (N_27499,N_26718,N_26418);
nor U27500 (N_27500,N_26134,N_26672);
and U27501 (N_27501,N_26576,N_26098);
and U27502 (N_27502,N_26362,N_26636);
xnor U27503 (N_27503,N_26875,N_26722);
or U27504 (N_27504,N_26006,N_26903);
nor U27505 (N_27505,N_26143,N_26562);
and U27506 (N_27506,N_26189,N_26868);
nand U27507 (N_27507,N_26465,N_26103);
xor U27508 (N_27508,N_26921,N_26009);
nor U27509 (N_27509,N_26406,N_26323);
xnor U27510 (N_27510,N_26732,N_26556);
or U27511 (N_27511,N_26480,N_26806);
nor U27512 (N_27512,N_26193,N_26832);
or U27513 (N_27513,N_26830,N_26322);
xor U27514 (N_27514,N_26250,N_26142);
or U27515 (N_27515,N_26104,N_26751);
xnor U27516 (N_27516,N_26393,N_26540);
and U27517 (N_27517,N_26061,N_26784);
xnor U27518 (N_27518,N_26450,N_26920);
nand U27519 (N_27519,N_26811,N_26763);
and U27520 (N_27520,N_26611,N_26818);
and U27521 (N_27521,N_26291,N_26460);
and U27522 (N_27522,N_26190,N_26322);
nand U27523 (N_27523,N_26477,N_26449);
xnor U27524 (N_27524,N_26774,N_26556);
nand U27525 (N_27525,N_26041,N_26533);
and U27526 (N_27526,N_26069,N_26193);
xor U27527 (N_27527,N_26914,N_26105);
and U27528 (N_27528,N_26902,N_26692);
or U27529 (N_27529,N_26862,N_26480);
nand U27530 (N_27530,N_26671,N_26333);
or U27531 (N_27531,N_26991,N_26208);
and U27532 (N_27532,N_26195,N_26657);
xnor U27533 (N_27533,N_26519,N_26795);
nor U27534 (N_27534,N_26429,N_26463);
nor U27535 (N_27535,N_26410,N_26495);
or U27536 (N_27536,N_26728,N_26586);
xor U27537 (N_27537,N_26231,N_26938);
or U27538 (N_27538,N_26753,N_26132);
xnor U27539 (N_27539,N_26804,N_26139);
and U27540 (N_27540,N_26651,N_26237);
xor U27541 (N_27541,N_26908,N_26380);
or U27542 (N_27542,N_26862,N_26236);
xor U27543 (N_27543,N_26737,N_26008);
or U27544 (N_27544,N_26256,N_26018);
and U27545 (N_27545,N_26819,N_26612);
nor U27546 (N_27546,N_26214,N_26236);
xnor U27547 (N_27547,N_26510,N_26197);
or U27548 (N_27548,N_26398,N_26388);
xnor U27549 (N_27549,N_26474,N_26596);
nand U27550 (N_27550,N_26714,N_26125);
nand U27551 (N_27551,N_26276,N_26745);
nand U27552 (N_27552,N_26480,N_26061);
and U27553 (N_27553,N_26735,N_26410);
and U27554 (N_27554,N_26288,N_26435);
and U27555 (N_27555,N_26618,N_26955);
or U27556 (N_27556,N_26989,N_26559);
nor U27557 (N_27557,N_26507,N_26920);
nor U27558 (N_27558,N_26092,N_26749);
or U27559 (N_27559,N_26775,N_26023);
or U27560 (N_27560,N_26977,N_26556);
xnor U27561 (N_27561,N_26650,N_26720);
or U27562 (N_27562,N_26058,N_26654);
nand U27563 (N_27563,N_26287,N_26595);
and U27564 (N_27564,N_26493,N_26658);
or U27565 (N_27565,N_26307,N_26654);
or U27566 (N_27566,N_26147,N_26164);
and U27567 (N_27567,N_26118,N_26344);
xor U27568 (N_27568,N_26624,N_26898);
nor U27569 (N_27569,N_26814,N_26720);
nor U27570 (N_27570,N_26814,N_26938);
xnor U27571 (N_27571,N_26031,N_26732);
or U27572 (N_27572,N_26819,N_26727);
nand U27573 (N_27573,N_26549,N_26008);
or U27574 (N_27574,N_26702,N_26722);
or U27575 (N_27575,N_26125,N_26409);
and U27576 (N_27576,N_26493,N_26996);
nand U27577 (N_27577,N_26474,N_26587);
xnor U27578 (N_27578,N_26373,N_26967);
nor U27579 (N_27579,N_26725,N_26726);
and U27580 (N_27580,N_26233,N_26357);
xor U27581 (N_27581,N_26550,N_26298);
and U27582 (N_27582,N_26479,N_26163);
and U27583 (N_27583,N_26470,N_26639);
and U27584 (N_27584,N_26946,N_26194);
or U27585 (N_27585,N_26003,N_26006);
and U27586 (N_27586,N_26092,N_26871);
xor U27587 (N_27587,N_26962,N_26352);
or U27588 (N_27588,N_26651,N_26973);
and U27589 (N_27589,N_26697,N_26434);
nand U27590 (N_27590,N_26854,N_26413);
nand U27591 (N_27591,N_26512,N_26851);
nor U27592 (N_27592,N_26616,N_26734);
xnor U27593 (N_27593,N_26356,N_26773);
xor U27594 (N_27594,N_26072,N_26847);
and U27595 (N_27595,N_26347,N_26234);
or U27596 (N_27596,N_26214,N_26150);
or U27597 (N_27597,N_26094,N_26694);
and U27598 (N_27598,N_26263,N_26672);
or U27599 (N_27599,N_26655,N_26155);
and U27600 (N_27600,N_26272,N_26341);
nand U27601 (N_27601,N_26234,N_26080);
or U27602 (N_27602,N_26372,N_26608);
and U27603 (N_27603,N_26551,N_26310);
xor U27604 (N_27604,N_26707,N_26528);
xor U27605 (N_27605,N_26477,N_26521);
nand U27606 (N_27606,N_26247,N_26096);
xnor U27607 (N_27607,N_26595,N_26706);
or U27608 (N_27608,N_26395,N_26655);
or U27609 (N_27609,N_26274,N_26169);
or U27610 (N_27610,N_26642,N_26313);
xor U27611 (N_27611,N_26165,N_26399);
or U27612 (N_27612,N_26550,N_26456);
xor U27613 (N_27613,N_26316,N_26418);
xnor U27614 (N_27614,N_26318,N_26963);
nand U27615 (N_27615,N_26198,N_26794);
nor U27616 (N_27616,N_26978,N_26706);
and U27617 (N_27617,N_26695,N_26251);
or U27618 (N_27618,N_26360,N_26846);
nand U27619 (N_27619,N_26962,N_26621);
nand U27620 (N_27620,N_26212,N_26314);
xnor U27621 (N_27621,N_26734,N_26760);
xor U27622 (N_27622,N_26527,N_26624);
nor U27623 (N_27623,N_26362,N_26167);
or U27624 (N_27624,N_26877,N_26074);
or U27625 (N_27625,N_26910,N_26505);
or U27626 (N_27626,N_26816,N_26943);
nor U27627 (N_27627,N_26316,N_26554);
nor U27628 (N_27628,N_26861,N_26275);
or U27629 (N_27629,N_26255,N_26434);
nor U27630 (N_27630,N_26555,N_26204);
nand U27631 (N_27631,N_26031,N_26150);
nor U27632 (N_27632,N_26807,N_26296);
nor U27633 (N_27633,N_26306,N_26801);
and U27634 (N_27634,N_26382,N_26943);
and U27635 (N_27635,N_26197,N_26229);
or U27636 (N_27636,N_26538,N_26544);
xnor U27637 (N_27637,N_26123,N_26602);
or U27638 (N_27638,N_26933,N_26786);
and U27639 (N_27639,N_26890,N_26031);
nand U27640 (N_27640,N_26912,N_26345);
xnor U27641 (N_27641,N_26518,N_26092);
nand U27642 (N_27642,N_26524,N_26748);
or U27643 (N_27643,N_26130,N_26494);
nor U27644 (N_27644,N_26300,N_26244);
nand U27645 (N_27645,N_26981,N_26234);
nand U27646 (N_27646,N_26559,N_26080);
and U27647 (N_27647,N_26989,N_26467);
nand U27648 (N_27648,N_26519,N_26474);
or U27649 (N_27649,N_26066,N_26713);
or U27650 (N_27650,N_26895,N_26969);
nor U27651 (N_27651,N_26306,N_26279);
xnor U27652 (N_27652,N_26590,N_26821);
xor U27653 (N_27653,N_26709,N_26935);
xor U27654 (N_27654,N_26117,N_26457);
xor U27655 (N_27655,N_26261,N_26759);
and U27656 (N_27656,N_26062,N_26409);
or U27657 (N_27657,N_26912,N_26872);
or U27658 (N_27658,N_26680,N_26484);
nand U27659 (N_27659,N_26321,N_26330);
nand U27660 (N_27660,N_26637,N_26324);
or U27661 (N_27661,N_26305,N_26268);
xor U27662 (N_27662,N_26737,N_26161);
nor U27663 (N_27663,N_26953,N_26187);
xor U27664 (N_27664,N_26091,N_26403);
or U27665 (N_27665,N_26403,N_26772);
xnor U27666 (N_27666,N_26847,N_26544);
xor U27667 (N_27667,N_26577,N_26915);
xnor U27668 (N_27668,N_26441,N_26038);
nand U27669 (N_27669,N_26461,N_26903);
nand U27670 (N_27670,N_26579,N_26446);
and U27671 (N_27671,N_26737,N_26473);
nor U27672 (N_27672,N_26680,N_26056);
xnor U27673 (N_27673,N_26660,N_26827);
nor U27674 (N_27674,N_26951,N_26175);
nor U27675 (N_27675,N_26134,N_26469);
or U27676 (N_27676,N_26325,N_26046);
or U27677 (N_27677,N_26321,N_26699);
xor U27678 (N_27678,N_26539,N_26478);
and U27679 (N_27679,N_26918,N_26225);
or U27680 (N_27680,N_26600,N_26294);
or U27681 (N_27681,N_26328,N_26164);
or U27682 (N_27682,N_26878,N_26589);
nand U27683 (N_27683,N_26360,N_26218);
and U27684 (N_27684,N_26905,N_26991);
or U27685 (N_27685,N_26640,N_26885);
and U27686 (N_27686,N_26954,N_26668);
nand U27687 (N_27687,N_26776,N_26934);
xnor U27688 (N_27688,N_26016,N_26697);
or U27689 (N_27689,N_26754,N_26923);
nand U27690 (N_27690,N_26746,N_26811);
xnor U27691 (N_27691,N_26338,N_26518);
or U27692 (N_27692,N_26994,N_26711);
or U27693 (N_27693,N_26385,N_26203);
and U27694 (N_27694,N_26523,N_26145);
nor U27695 (N_27695,N_26907,N_26771);
nand U27696 (N_27696,N_26254,N_26120);
xnor U27697 (N_27697,N_26284,N_26579);
xnor U27698 (N_27698,N_26242,N_26982);
xnor U27699 (N_27699,N_26865,N_26297);
nand U27700 (N_27700,N_26992,N_26467);
nand U27701 (N_27701,N_26184,N_26107);
xor U27702 (N_27702,N_26666,N_26875);
and U27703 (N_27703,N_26029,N_26726);
xnor U27704 (N_27704,N_26815,N_26963);
nand U27705 (N_27705,N_26084,N_26281);
or U27706 (N_27706,N_26724,N_26492);
nand U27707 (N_27707,N_26109,N_26079);
and U27708 (N_27708,N_26359,N_26202);
xnor U27709 (N_27709,N_26424,N_26845);
or U27710 (N_27710,N_26619,N_26165);
xor U27711 (N_27711,N_26968,N_26466);
or U27712 (N_27712,N_26999,N_26548);
nor U27713 (N_27713,N_26411,N_26776);
and U27714 (N_27714,N_26667,N_26981);
nor U27715 (N_27715,N_26562,N_26152);
and U27716 (N_27716,N_26314,N_26116);
xor U27717 (N_27717,N_26792,N_26505);
nor U27718 (N_27718,N_26054,N_26934);
nand U27719 (N_27719,N_26027,N_26299);
nor U27720 (N_27720,N_26271,N_26448);
xor U27721 (N_27721,N_26308,N_26042);
and U27722 (N_27722,N_26867,N_26864);
or U27723 (N_27723,N_26771,N_26682);
nor U27724 (N_27724,N_26538,N_26738);
and U27725 (N_27725,N_26381,N_26739);
nor U27726 (N_27726,N_26831,N_26070);
and U27727 (N_27727,N_26521,N_26446);
or U27728 (N_27728,N_26869,N_26609);
xor U27729 (N_27729,N_26029,N_26160);
nor U27730 (N_27730,N_26556,N_26316);
xor U27731 (N_27731,N_26664,N_26232);
or U27732 (N_27732,N_26486,N_26972);
nor U27733 (N_27733,N_26491,N_26701);
or U27734 (N_27734,N_26458,N_26010);
nor U27735 (N_27735,N_26936,N_26496);
and U27736 (N_27736,N_26526,N_26705);
xnor U27737 (N_27737,N_26940,N_26752);
nor U27738 (N_27738,N_26880,N_26504);
nor U27739 (N_27739,N_26097,N_26628);
nand U27740 (N_27740,N_26245,N_26911);
nand U27741 (N_27741,N_26916,N_26909);
and U27742 (N_27742,N_26162,N_26896);
or U27743 (N_27743,N_26835,N_26447);
nor U27744 (N_27744,N_26143,N_26203);
xnor U27745 (N_27745,N_26407,N_26061);
or U27746 (N_27746,N_26797,N_26059);
nand U27747 (N_27747,N_26400,N_26256);
or U27748 (N_27748,N_26095,N_26044);
nor U27749 (N_27749,N_26574,N_26946);
or U27750 (N_27750,N_26245,N_26834);
and U27751 (N_27751,N_26275,N_26002);
nand U27752 (N_27752,N_26822,N_26326);
nor U27753 (N_27753,N_26789,N_26436);
nor U27754 (N_27754,N_26944,N_26169);
nand U27755 (N_27755,N_26309,N_26029);
nand U27756 (N_27756,N_26122,N_26741);
or U27757 (N_27757,N_26444,N_26230);
xor U27758 (N_27758,N_26662,N_26827);
or U27759 (N_27759,N_26090,N_26659);
xor U27760 (N_27760,N_26800,N_26094);
nor U27761 (N_27761,N_26242,N_26776);
nand U27762 (N_27762,N_26301,N_26894);
xnor U27763 (N_27763,N_26213,N_26245);
and U27764 (N_27764,N_26997,N_26014);
and U27765 (N_27765,N_26580,N_26975);
nand U27766 (N_27766,N_26001,N_26147);
nor U27767 (N_27767,N_26590,N_26197);
nand U27768 (N_27768,N_26180,N_26301);
nor U27769 (N_27769,N_26650,N_26464);
or U27770 (N_27770,N_26987,N_26819);
xnor U27771 (N_27771,N_26475,N_26222);
nand U27772 (N_27772,N_26039,N_26783);
or U27773 (N_27773,N_26104,N_26936);
or U27774 (N_27774,N_26191,N_26440);
or U27775 (N_27775,N_26339,N_26367);
nand U27776 (N_27776,N_26418,N_26938);
nand U27777 (N_27777,N_26794,N_26110);
nor U27778 (N_27778,N_26307,N_26803);
or U27779 (N_27779,N_26187,N_26752);
xnor U27780 (N_27780,N_26782,N_26530);
or U27781 (N_27781,N_26832,N_26339);
or U27782 (N_27782,N_26333,N_26103);
xor U27783 (N_27783,N_26103,N_26162);
and U27784 (N_27784,N_26293,N_26996);
nand U27785 (N_27785,N_26741,N_26145);
and U27786 (N_27786,N_26332,N_26364);
xor U27787 (N_27787,N_26987,N_26522);
xnor U27788 (N_27788,N_26329,N_26986);
nand U27789 (N_27789,N_26065,N_26916);
xnor U27790 (N_27790,N_26854,N_26173);
nand U27791 (N_27791,N_26232,N_26073);
nor U27792 (N_27792,N_26628,N_26369);
nor U27793 (N_27793,N_26051,N_26818);
nand U27794 (N_27794,N_26333,N_26945);
xor U27795 (N_27795,N_26037,N_26215);
and U27796 (N_27796,N_26543,N_26166);
or U27797 (N_27797,N_26365,N_26670);
nand U27798 (N_27798,N_26035,N_26625);
or U27799 (N_27799,N_26474,N_26466);
and U27800 (N_27800,N_26305,N_26452);
xor U27801 (N_27801,N_26715,N_26773);
nor U27802 (N_27802,N_26082,N_26272);
xnor U27803 (N_27803,N_26182,N_26641);
nand U27804 (N_27804,N_26368,N_26355);
and U27805 (N_27805,N_26033,N_26533);
nand U27806 (N_27806,N_26396,N_26052);
nor U27807 (N_27807,N_26224,N_26747);
xnor U27808 (N_27808,N_26338,N_26971);
nand U27809 (N_27809,N_26257,N_26872);
nand U27810 (N_27810,N_26121,N_26609);
or U27811 (N_27811,N_26589,N_26933);
nor U27812 (N_27812,N_26781,N_26546);
or U27813 (N_27813,N_26577,N_26885);
xnor U27814 (N_27814,N_26148,N_26314);
and U27815 (N_27815,N_26898,N_26035);
nor U27816 (N_27816,N_26995,N_26981);
and U27817 (N_27817,N_26988,N_26410);
nor U27818 (N_27818,N_26433,N_26471);
nor U27819 (N_27819,N_26589,N_26800);
nor U27820 (N_27820,N_26026,N_26070);
or U27821 (N_27821,N_26654,N_26325);
nor U27822 (N_27822,N_26202,N_26447);
nor U27823 (N_27823,N_26800,N_26929);
nor U27824 (N_27824,N_26831,N_26351);
nand U27825 (N_27825,N_26519,N_26948);
and U27826 (N_27826,N_26635,N_26272);
nor U27827 (N_27827,N_26823,N_26020);
xnor U27828 (N_27828,N_26582,N_26481);
nor U27829 (N_27829,N_26386,N_26853);
and U27830 (N_27830,N_26578,N_26996);
nor U27831 (N_27831,N_26222,N_26587);
nand U27832 (N_27832,N_26090,N_26430);
and U27833 (N_27833,N_26512,N_26359);
nand U27834 (N_27834,N_26996,N_26171);
nor U27835 (N_27835,N_26707,N_26519);
nand U27836 (N_27836,N_26597,N_26565);
and U27837 (N_27837,N_26720,N_26931);
and U27838 (N_27838,N_26097,N_26269);
or U27839 (N_27839,N_26497,N_26609);
and U27840 (N_27840,N_26941,N_26287);
or U27841 (N_27841,N_26823,N_26155);
nand U27842 (N_27842,N_26422,N_26430);
and U27843 (N_27843,N_26638,N_26582);
nor U27844 (N_27844,N_26871,N_26814);
or U27845 (N_27845,N_26107,N_26868);
and U27846 (N_27846,N_26662,N_26729);
xor U27847 (N_27847,N_26419,N_26651);
xnor U27848 (N_27848,N_26064,N_26047);
nand U27849 (N_27849,N_26669,N_26218);
nor U27850 (N_27850,N_26470,N_26028);
and U27851 (N_27851,N_26811,N_26986);
xnor U27852 (N_27852,N_26625,N_26817);
or U27853 (N_27853,N_26649,N_26998);
nand U27854 (N_27854,N_26835,N_26321);
nor U27855 (N_27855,N_26582,N_26533);
nand U27856 (N_27856,N_26434,N_26371);
nor U27857 (N_27857,N_26888,N_26613);
or U27858 (N_27858,N_26136,N_26392);
nand U27859 (N_27859,N_26523,N_26660);
or U27860 (N_27860,N_26864,N_26924);
xnor U27861 (N_27861,N_26356,N_26143);
nand U27862 (N_27862,N_26232,N_26199);
and U27863 (N_27863,N_26629,N_26500);
xnor U27864 (N_27864,N_26096,N_26582);
or U27865 (N_27865,N_26027,N_26742);
nor U27866 (N_27866,N_26124,N_26989);
xnor U27867 (N_27867,N_26898,N_26538);
xor U27868 (N_27868,N_26339,N_26907);
nand U27869 (N_27869,N_26098,N_26753);
nand U27870 (N_27870,N_26654,N_26699);
and U27871 (N_27871,N_26099,N_26391);
xnor U27872 (N_27872,N_26932,N_26705);
or U27873 (N_27873,N_26098,N_26447);
or U27874 (N_27874,N_26988,N_26969);
nor U27875 (N_27875,N_26274,N_26095);
xor U27876 (N_27876,N_26675,N_26639);
and U27877 (N_27877,N_26376,N_26683);
or U27878 (N_27878,N_26265,N_26838);
xor U27879 (N_27879,N_26409,N_26675);
or U27880 (N_27880,N_26840,N_26603);
xnor U27881 (N_27881,N_26804,N_26321);
nand U27882 (N_27882,N_26364,N_26998);
nor U27883 (N_27883,N_26391,N_26349);
nor U27884 (N_27884,N_26564,N_26824);
nor U27885 (N_27885,N_26133,N_26865);
nand U27886 (N_27886,N_26267,N_26769);
and U27887 (N_27887,N_26910,N_26620);
or U27888 (N_27888,N_26243,N_26054);
nand U27889 (N_27889,N_26537,N_26208);
nand U27890 (N_27890,N_26267,N_26696);
or U27891 (N_27891,N_26682,N_26034);
nand U27892 (N_27892,N_26697,N_26603);
xor U27893 (N_27893,N_26594,N_26214);
and U27894 (N_27894,N_26559,N_26711);
or U27895 (N_27895,N_26614,N_26912);
xnor U27896 (N_27896,N_26835,N_26359);
or U27897 (N_27897,N_26185,N_26386);
xor U27898 (N_27898,N_26204,N_26396);
and U27899 (N_27899,N_26818,N_26249);
and U27900 (N_27900,N_26046,N_26556);
nand U27901 (N_27901,N_26714,N_26816);
xnor U27902 (N_27902,N_26033,N_26380);
nand U27903 (N_27903,N_26958,N_26581);
nor U27904 (N_27904,N_26799,N_26685);
xnor U27905 (N_27905,N_26801,N_26038);
xor U27906 (N_27906,N_26433,N_26987);
and U27907 (N_27907,N_26277,N_26788);
nand U27908 (N_27908,N_26698,N_26601);
xnor U27909 (N_27909,N_26895,N_26906);
or U27910 (N_27910,N_26276,N_26562);
nand U27911 (N_27911,N_26951,N_26609);
xnor U27912 (N_27912,N_26827,N_26049);
or U27913 (N_27913,N_26664,N_26939);
and U27914 (N_27914,N_26506,N_26723);
or U27915 (N_27915,N_26082,N_26960);
nand U27916 (N_27916,N_26382,N_26165);
or U27917 (N_27917,N_26237,N_26657);
nand U27918 (N_27918,N_26623,N_26827);
and U27919 (N_27919,N_26862,N_26918);
nand U27920 (N_27920,N_26481,N_26691);
and U27921 (N_27921,N_26139,N_26696);
and U27922 (N_27922,N_26077,N_26553);
xnor U27923 (N_27923,N_26834,N_26953);
or U27924 (N_27924,N_26625,N_26094);
or U27925 (N_27925,N_26428,N_26854);
nand U27926 (N_27926,N_26418,N_26337);
or U27927 (N_27927,N_26663,N_26424);
xor U27928 (N_27928,N_26652,N_26753);
xnor U27929 (N_27929,N_26910,N_26470);
xor U27930 (N_27930,N_26969,N_26721);
or U27931 (N_27931,N_26063,N_26923);
and U27932 (N_27932,N_26738,N_26015);
or U27933 (N_27933,N_26146,N_26460);
nand U27934 (N_27934,N_26530,N_26825);
nand U27935 (N_27935,N_26388,N_26308);
or U27936 (N_27936,N_26276,N_26578);
or U27937 (N_27937,N_26157,N_26873);
nor U27938 (N_27938,N_26068,N_26244);
or U27939 (N_27939,N_26693,N_26314);
nand U27940 (N_27940,N_26269,N_26795);
and U27941 (N_27941,N_26273,N_26227);
xor U27942 (N_27942,N_26277,N_26053);
nor U27943 (N_27943,N_26671,N_26298);
and U27944 (N_27944,N_26826,N_26552);
nor U27945 (N_27945,N_26048,N_26690);
or U27946 (N_27946,N_26955,N_26734);
nand U27947 (N_27947,N_26517,N_26365);
or U27948 (N_27948,N_26487,N_26872);
and U27949 (N_27949,N_26945,N_26230);
nor U27950 (N_27950,N_26179,N_26286);
nand U27951 (N_27951,N_26152,N_26849);
xor U27952 (N_27952,N_26149,N_26718);
or U27953 (N_27953,N_26614,N_26040);
and U27954 (N_27954,N_26340,N_26911);
xor U27955 (N_27955,N_26186,N_26730);
nand U27956 (N_27956,N_26759,N_26313);
nor U27957 (N_27957,N_26733,N_26897);
nand U27958 (N_27958,N_26575,N_26270);
nor U27959 (N_27959,N_26914,N_26006);
or U27960 (N_27960,N_26499,N_26918);
or U27961 (N_27961,N_26668,N_26013);
and U27962 (N_27962,N_26896,N_26444);
or U27963 (N_27963,N_26880,N_26980);
nor U27964 (N_27964,N_26098,N_26253);
or U27965 (N_27965,N_26136,N_26934);
or U27966 (N_27966,N_26066,N_26072);
nand U27967 (N_27967,N_26732,N_26986);
nand U27968 (N_27968,N_26275,N_26820);
xnor U27969 (N_27969,N_26067,N_26969);
nor U27970 (N_27970,N_26816,N_26258);
xor U27971 (N_27971,N_26287,N_26171);
nand U27972 (N_27972,N_26184,N_26474);
xor U27973 (N_27973,N_26303,N_26204);
xnor U27974 (N_27974,N_26277,N_26188);
nor U27975 (N_27975,N_26423,N_26965);
nand U27976 (N_27976,N_26454,N_26513);
and U27977 (N_27977,N_26232,N_26583);
nor U27978 (N_27978,N_26902,N_26192);
nand U27979 (N_27979,N_26016,N_26341);
xnor U27980 (N_27980,N_26572,N_26960);
or U27981 (N_27981,N_26791,N_26039);
nor U27982 (N_27982,N_26685,N_26167);
nor U27983 (N_27983,N_26642,N_26501);
or U27984 (N_27984,N_26307,N_26814);
xor U27985 (N_27985,N_26198,N_26837);
and U27986 (N_27986,N_26228,N_26608);
and U27987 (N_27987,N_26412,N_26593);
nor U27988 (N_27988,N_26330,N_26210);
and U27989 (N_27989,N_26322,N_26281);
xnor U27990 (N_27990,N_26010,N_26835);
nor U27991 (N_27991,N_26472,N_26060);
or U27992 (N_27992,N_26901,N_26149);
nor U27993 (N_27993,N_26985,N_26569);
xnor U27994 (N_27994,N_26047,N_26667);
and U27995 (N_27995,N_26069,N_26907);
or U27996 (N_27996,N_26455,N_26164);
nor U27997 (N_27997,N_26406,N_26353);
and U27998 (N_27998,N_26909,N_26230);
nand U27999 (N_27999,N_26680,N_26912);
xnor U28000 (N_28000,N_27537,N_27070);
xor U28001 (N_28001,N_27243,N_27607);
or U28002 (N_28002,N_27965,N_27720);
xnor U28003 (N_28003,N_27928,N_27896);
nor U28004 (N_28004,N_27980,N_27557);
and U28005 (N_28005,N_27509,N_27016);
nor U28006 (N_28006,N_27769,N_27358);
and U28007 (N_28007,N_27879,N_27741);
xor U28008 (N_28008,N_27080,N_27411);
nor U28009 (N_28009,N_27838,N_27356);
or U28010 (N_28010,N_27245,N_27929);
and U28011 (N_28011,N_27757,N_27440);
nand U28012 (N_28012,N_27620,N_27298);
nor U28013 (N_28013,N_27864,N_27469);
nor U28014 (N_28014,N_27359,N_27340);
nand U28015 (N_28015,N_27944,N_27427);
nor U28016 (N_28016,N_27746,N_27289);
xnor U28017 (N_28017,N_27898,N_27744);
xor U28018 (N_28018,N_27074,N_27584);
and U28019 (N_28019,N_27131,N_27903);
nand U28020 (N_28020,N_27522,N_27867);
or U28021 (N_28021,N_27303,N_27514);
nand U28022 (N_28022,N_27486,N_27508);
xnor U28023 (N_28023,N_27588,N_27192);
nor U28024 (N_28024,N_27994,N_27028);
and U28025 (N_28025,N_27548,N_27265);
and U28026 (N_28026,N_27329,N_27585);
nor U28027 (N_28027,N_27462,N_27546);
and U28028 (N_28028,N_27609,N_27996);
or U28029 (N_28029,N_27800,N_27873);
nand U28030 (N_28030,N_27060,N_27085);
nand U28031 (N_28031,N_27404,N_27180);
nand U28032 (N_28032,N_27433,N_27513);
and U28033 (N_28033,N_27815,N_27376);
xor U28034 (N_28034,N_27268,N_27266);
nand U28035 (N_28035,N_27910,N_27498);
nor U28036 (N_28036,N_27906,N_27130);
nor U28037 (N_28037,N_27687,N_27912);
nand U28038 (N_28038,N_27354,N_27051);
or U28039 (N_28039,N_27064,N_27895);
nor U28040 (N_28040,N_27317,N_27567);
nand U28041 (N_28041,N_27461,N_27009);
and U28042 (N_28042,N_27869,N_27738);
nand U28043 (N_28043,N_27295,N_27342);
nand U28044 (N_28044,N_27553,N_27050);
nor U28045 (N_28045,N_27856,N_27690);
and U28046 (N_28046,N_27883,N_27021);
nor U28047 (N_28047,N_27715,N_27586);
nor U28048 (N_28048,N_27076,N_27111);
nor U28049 (N_28049,N_27971,N_27463);
xor U28050 (N_28050,N_27940,N_27497);
or U28051 (N_28051,N_27067,N_27972);
xnor U28052 (N_28052,N_27652,N_27413);
nand U28053 (N_28053,N_27917,N_27791);
nor U28054 (N_28054,N_27097,N_27332);
and U28055 (N_28055,N_27391,N_27885);
nor U28056 (N_28056,N_27015,N_27890);
or U28057 (N_28057,N_27273,N_27538);
xnor U28058 (N_28058,N_27642,N_27673);
nand U28059 (N_28059,N_27197,N_27569);
xor U28060 (N_28060,N_27333,N_27783);
or U28061 (N_28061,N_27252,N_27580);
and U28062 (N_28062,N_27119,N_27065);
nor U28063 (N_28063,N_27478,N_27357);
xor U28064 (N_28064,N_27520,N_27098);
nor U28065 (N_28065,N_27563,N_27312);
or U28066 (N_28066,N_27978,N_27694);
and U28067 (N_28067,N_27795,N_27045);
nand U28068 (N_28068,N_27169,N_27679);
nor U28069 (N_28069,N_27701,N_27026);
nor U28070 (N_28070,N_27682,N_27794);
and U28071 (N_28071,N_27108,N_27785);
nor U28072 (N_28072,N_27886,N_27379);
nand U28073 (N_28073,N_27825,N_27345);
and U28074 (N_28074,N_27594,N_27331);
and U28075 (N_28075,N_27846,N_27240);
or U28076 (N_28076,N_27324,N_27849);
nor U28077 (N_28077,N_27079,N_27836);
nand U28078 (N_28078,N_27595,N_27933);
xnor U28079 (N_28079,N_27658,N_27742);
or U28080 (N_28080,N_27488,N_27048);
nand U28081 (N_28081,N_27540,N_27090);
nand U28082 (N_28082,N_27824,N_27258);
nor U28083 (N_28083,N_27439,N_27942);
xor U28084 (N_28084,N_27308,N_27422);
or U28085 (N_28085,N_27179,N_27985);
and U28086 (N_28086,N_27292,N_27128);
or U28087 (N_28087,N_27750,N_27274);
and U28088 (N_28088,N_27449,N_27804);
nand U28089 (N_28089,N_27539,N_27704);
or U28090 (N_28090,N_27407,N_27531);
or U28091 (N_28091,N_27611,N_27362);
and U28092 (N_28092,N_27955,N_27001);
xnor U28093 (N_28093,N_27646,N_27394);
and U28094 (N_28094,N_27475,N_27801);
xor U28095 (N_28095,N_27773,N_27979);
or U28096 (N_28096,N_27444,N_27161);
nand U28097 (N_28097,N_27623,N_27091);
xor U28098 (N_28098,N_27392,N_27094);
nor U28099 (N_28099,N_27645,N_27571);
and U28100 (N_28100,N_27878,N_27326);
or U28101 (N_28101,N_27970,N_27071);
or U28102 (N_28102,N_27668,N_27894);
nand U28103 (N_28103,N_27854,N_27605);
and U28104 (N_28104,N_27663,N_27655);
nor U28105 (N_28105,N_27230,N_27374);
xnor U28106 (N_28106,N_27707,N_27525);
nand U28107 (N_28107,N_27100,N_27235);
nand U28108 (N_28108,N_27175,N_27466);
nand U28109 (N_28109,N_27448,N_27226);
xor U28110 (N_28110,N_27981,N_27352);
xnor U28111 (N_28111,N_27116,N_27556);
or U28112 (N_28112,N_27541,N_27176);
xor U28113 (N_28113,N_27321,N_27477);
and U28114 (N_28114,N_27195,N_27968);
nand U28115 (N_28115,N_27964,N_27617);
and U28116 (N_28116,N_27877,N_27950);
or U28117 (N_28117,N_27241,N_27960);
and U28118 (N_28118,N_27671,N_27012);
nand U28119 (N_28119,N_27523,N_27061);
nor U28120 (N_28120,N_27660,N_27386);
and U28121 (N_28121,N_27966,N_27405);
nand U28122 (N_28122,N_27634,N_27155);
nor U28123 (N_28123,N_27889,N_27731);
or U28124 (N_28124,N_27992,N_27231);
and U28125 (N_28125,N_27844,N_27493);
and U28126 (N_28126,N_27249,N_27749);
nand U28127 (N_28127,N_27246,N_27976);
nand U28128 (N_28128,N_27925,N_27082);
xor U28129 (N_28129,N_27023,N_27625);
xnor U28130 (N_28130,N_27202,N_27587);
nand U28131 (N_28131,N_27465,N_27763);
xor U28132 (N_28132,N_27272,N_27761);
and U28133 (N_28133,N_27115,N_27693);
xor U28134 (N_28134,N_27811,N_27712);
nand U28135 (N_28135,N_27217,N_27304);
nor U28136 (N_28136,N_27892,N_27207);
and U28137 (N_28137,N_27828,N_27166);
xor U28138 (N_28138,N_27796,N_27043);
and U28139 (N_28139,N_27963,N_27181);
xor U28140 (N_28140,N_27482,N_27766);
xor U28141 (N_28141,N_27410,N_27771);
or U28142 (N_28142,N_27888,N_27740);
xnor U28143 (N_28143,N_27492,N_27852);
xnor U28144 (N_28144,N_27095,N_27135);
and U28145 (N_28145,N_27904,N_27423);
or U28146 (N_28146,N_27053,N_27913);
or U28147 (N_28147,N_27284,N_27042);
and U28148 (N_28148,N_27511,N_27914);
and U28149 (N_28149,N_27535,N_27821);
nand U28150 (N_28150,N_27574,N_27237);
and U28151 (N_28151,N_27490,N_27121);
nor U28152 (N_28152,N_27114,N_27417);
nor U28153 (N_28153,N_27283,N_27174);
and U28154 (N_28154,N_27103,N_27911);
and U28155 (N_28155,N_27568,N_27677);
nand U28156 (N_28156,N_27491,N_27057);
and U28157 (N_28157,N_27562,N_27680);
xor U28158 (N_28158,N_27613,N_27743);
nor U28159 (N_28159,N_27455,N_27089);
or U28160 (N_28160,N_27020,N_27809);
or U28161 (N_28161,N_27058,N_27558);
nand U28162 (N_28162,N_27191,N_27120);
and U28163 (N_28163,N_27615,N_27722);
nor U28164 (N_28164,N_27907,N_27714);
nor U28165 (N_28165,N_27827,N_27918);
or U28166 (N_28166,N_27361,N_27393);
xor U28167 (N_28167,N_27142,N_27154);
nor U28168 (N_28168,N_27922,N_27036);
or U28169 (N_28169,N_27375,N_27242);
nor U28170 (N_28170,N_27755,N_27019);
or U28171 (N_28171,N_27691,N_27054);
xor U28172 (N_28172,N_27807,N_27112);
or U28173 (N_28173,N_27816,N_27034);
or U28174 (N_28174,N_27203,N_27117);
xor U28175 (N_28175,N_27624,N_27654);
xnor U28176 (N_28176,N_27573,N_27382);
xor U28177 (N_28177,N_27871,N_27257);
xor U28178 (N_28178,N_27941,N_27335);
xor U28179 (N_28179,N_27052,N_27832);
nand U28180 (N_28180,N_27962,N_27592);
and U28181 (N_28181,N_27544,N_27432);
nand U28182 (N_28182,N_27631,N_27075);
nor U28183 (N_28183,N_27850,N_27589);
nand U28184 (N_28184,N_27279,N_27096);
or U28185 (N_28185,N_27576,N_27723);
nand U28186 (N_28186,N_27480,N_27774);
nor U28187 (N_28187,N_27819,N_27733);
xnor U28188 (N_28188,N_27296,N_27088);
nand U28189 (N_28189,N_27572,N_27087);
nand U28190 (N_28190,N_27126,N_27024);
nand U28191 (N_28191,N_27734,N_27545);
or U28192 (N_28192,N_27281,N_27891);
and U28193 (N_28193,N_27365,N_27737);
and U28194 (N_28194,N_27177,N_27772);
or U28195 (N_28195,N_27378,N_27834);
or U28196 (N_28196,N_27014,N_27225);
or U28197 (N_28197,N_27270,N_27923);
xor U28198 (N_28198,N_27990,N_27718);
nand U28199 (N_28199,N_27046,N_27775);
nand U28200 (N_28200,N_27041,N_27288);
nor U28201 (N_28201,N_27355,N_27218);
nor U28202 (N_28202,N_27614,N_27697);
or U28203 (N_28203,N_27047,N_27063);
nor U28204 (N_28204,N_27152,N_27496);
nand U28205 (N_28205,N_27833,N_27908);
and U28206 (N_28206,N_27618,N_27030);
or U28207 (N_28207,N_27729,N_27140);
and U28208 (N_28208,N_27073,N_27487);
nor U28209 (N_28209,N_27211,N_27946);
nand U28210 (N_28210,N_27322,N_27300);
nor U28211 (N_28211,N_27032,N_27204);
xnor U28212 (N_28212,N_27670,N_27591);
xor U28213 (N_28213,N_27336,N_27829);
or U28214 (N_28214,N_27228,N_27993);
and U28215 (N_28215,N_27022,N_27629);
and U28216 (N_28216,N_27689,N_27706);
xnor U28217 (N_28217,N_27752,N_27485);
xnor U28218 (N_28218,N_27987,N_27380);
nor U28219 (N_28219,N_27789,N_27414);
nand U28220 (N_28220,N_27975,N_27010);
xnor U28221 (N_28221,N_27899,N_27708);
xor U28222 (N_28222,N_27453,N_27748);
and U28223 (N_28223,N_27632,N_27710);
nand U28224 (N_28224,N_27650,N_27859);
and U28225 (N_28225,N_27244,N_27639);
nand U28226 (N_28226,N_27503,N_27307);
or U28227 (N_28227,N_27805,N_27921);
xnor U28228 (N_28228,N_27839,N_27713);
and U28229 (N_28229,N_27530,N_27612);
or U28230 (N_28230,N_27139,N_27719);
nor U28231 (N_28231,N_27068,N_27973);
nor U28232 (N_28232,N_27893,N_27472);
xor U28233 (N_28233,N_27346,N_27776);
nor U28234 (N_28234,N_27408,N_27986);
and U28235 (N_28235,N_27025,N_27875);
and U28236 (N_28236,N_27982,N_27703);
nor U28237 (N_28237,N_27419,N_27418);
or U28238 (N_28238,N_27649,N_27328);
nor U28239 (N_28239,N_27797,N_27297);
xnor U28240 (N_28240,N_27118,N_27446);
and U28241 (N_28241,N_27364,N_27932);
and U28242 (N_28242,N_27313,N_27939);
nor U28243 (N_28243,N_27997,N_27915);
and U28244 (N_28244,N_27644,N_27726);
nor U28245 (N_28245,N_27311,N_27178);
or U28246 (N_28246,N_27262,N_27847);
nand U28247 (N_28247,N_27387,N_27919);
or U28248 (N_28248,N_27113,N_27189);
nand U28249 (N_28249,N_27788,N_27764);
xnor U28250 (N_28250,N_27759,N_27143);
nand U28251 (N_28251,N_27212,N_27006);
or U28252 (N_28252,N_27138,N_27709);
xor U28253 (N_28253,N_27206,N_27843);
or U28254 (N_28254,N_27861,N_27167);
or U28255 (N_28255,N_27483,N_27429);
xor U28256 (N_28256,N_27552,N_27106);
nand U28257 (N_28257,N_27153,N_27467);
nor U28258 (N_28258,N_27782,N_27123);
xor U28259 (N_28259,N_27416,N_27450);
xor U28260 (N_28260,N_27216,N_27842);
xor U28261 (N_28261,N_27855,N_27033);
nand U28262 (N_28262,N_27435,N_27817);
or U28263 (N_28263,N_27686,N_27724);
and U28264 (N_28264,N_27610,N_27661);
and U28265 (N_28265,N_27575,N_27157);
nor U28266 (N_28266,N_27255,N_27725);
xnor U28267 (N_28267,N_27334,N_27698);
nand U28268 (N_28268,N_27314,N_27367);
and U28269 (N_28269,N_27412,N_27991);
nor U28270 (N_28270,N_27659,N_27578);
and U28271 (N_28271,N_27129,N_27995);
or U28272 (N_28272,N_27758,N_27347);
or U28273 (N_28273,N_27388,N_27264);
and U28274 (N_28274,N_27793,N_27002);
nand U28275 (N_28275,N_27762,N_27674);
nand U28276 (N_28276,N_27183,N_27348);
nor U28277 (N_28277,N_27747,N_27302);
nand U28278 (N_28278,N_27648,N_27389);
nor U28279 (N_28279,N_27507,N_27188);
nand U28280 (N_28280,N_27837,N_27851);
or U28281 (N_28281,N_27059,N_27489);
xor U28282 (N_28282,N_27187,N_27056);
and U28283 (N_28283,N_27325,N_27251);
xor U28284 (N_28284,N_27366,N_27476);
and U28285 (N_28285,N_27236,N_27865);
and U28286 (N_28286,N_27484,N_27299);
xor U28287 (N_28287,N_27456,N_27224);
nand U28288 (N_28288,N_27445,N_27261);
nand U28289 (N_28289,N_27579,N_27900);
or U28290 (N_28290,N_27559,N_27518);
nor U28291 (N_28291,N_27826,N_27603);
xnor U28292 (N_28292,N_27527,N_27437);
nor U28293 (N_28293,N_27868,N_27803);
xnor U28294 (N_28294,N_27606,N_27699);
and U28295 (N_28295,N_27370,N_27409);
and U28296 (N_28296,N_27007,N_27381);
nor U28297 (N_28297,N_27937,N_27641);
nor U28298 (N_28298,N_27049,N_27802);
xnor U28299 (N_28299,N_27813,N_27027);
xnor U28300 (N_28300,N_27777,N_27474);
xor U28301 (N_28301,N_27506,N_27627);
nor U28302 (N_28302,N_27306,N_27685);
and U28303 (N_28303,N_27460,N_27201);
nor U28304 (N_28304,N_27239,N_27555);
nor U28305 (N_28305,N_27711,N_27735);
nor U28306 (N_28306,N_27069,N_27424);
or U28307 (N_28307,N_27814,N_27526);
nand U28308 (N_28308,N_27044,N_27510);
and U28309 (N_28309,N_27521,N_27608);
nand U28310 (N_28310,N_27442,N_27248);
nor U28311 (N_28311,N_27227,N_27092);
and U28312 (N_28312,N_27055,N_27666);
and U28313 (N_28313,N_27305,N_27186);
nand U28314 (N_28314,N_27125,N_27728);
nand U28315 (N_28315,N_27502,N_27672);
and U28316 (N_28316,N_27247,N_27193);
or U28317 (N_28317,N_27280,N_27101);
nor U28318 (N_28318,N_27170,N_27294);
nor U28319 (N_28319,N_27458,N_27099);
xor U28320 (N_28320,N_27542,N_27209);
and U28321 (N_28321,N_27233,N_27372);
or U28322 (N_28322,N_27678,N_27371);
or U28323 (N_28323,N_27667,N_27754);
nand U28324 (N_28324,N_27337,N_27945);
nand U28325 (N_28325,N_27368,N_27549);
or U28326 (N_28326,N_27881,N_27451);
nor U28327 (N_28327,N_27554,N_27882);
xor U28328 (N_28328,N_27286,N_27078);
nor U28329 (N_28329,N_27160,N_27397);
nor U28330 (N_28330,N_27823,N_27626);
nor U28331 (N_28331,N_27086,N_27127);
nand U28332 (N_28332,N_27499,N_27778);
nand U28333 (N_28333,N_27401,N_27136);
and U28334 (N_28334,N_27700,N_27122);
nor U28335 (N_28335,N_27210,N_27818);
xnor U28336 (N_28336,N_27947,N_27820);
nand U28337 (N_28337,N_27341,N_27403);
xor U28338 (N_28338,N_27684,N_27145);
nor U28339 (N_28339,N_27384,N_27385);
xnor U28340 (N_28340,N_27692,N_27969);
xor U28341 (N_28341,N_27756,N_27504);
nor U28342 (N_28342,N_27884,N_27721);
nor U28343 (N_28343,N_27132,N_27452);
and U28344 (N_28344,N_27547,N_27038);
nor U28345 (N_28345,N_27105,N_27768);
nand U28346 (N_28346,N_27619,N_27560);
or U28347 (N_28347,N_27431,N_27287);
and U28348 (N_28348,N_27653,N_27159);
nor U28349 (N_28349,N_27256,N_27102);
or U28350 (N_28350,N_27315,N_27415);
and U28351 (N_28351,N_27172,N_27870);
nand U28352 (N_28352,N_27515,N_27581);
and U28353 (N_28353,N_27989,N_27214);
or U28354 (N_28354,N_27533,N_27936);
nor U28355 (N_28355,N_27219,N_27470);
nor U28356 (N_28356,N_27909,N_27200);
and U28357 (N_28357,N_27141,N_27013);
and U28358 (N_28358,N_27285,N_27164);
or U28359 (N_28359,N_27162,N_27146);
nor U28360 (N_28360,N_27902,N_27254);
nand U28361 (N_28361,N_27561,N_27271);
nand U28362 (N_28362,N_27309,N_27784);
nor U28363 (N_28363,N_27858,N_27039);
nor U28364 (N_28364,N_27320,N_27008);
nand U28365 (N_28365,N_27876,N_27812);
or U28366 (N_28366,N_27905,N_27590);
and U28367 (N_28367,N_27602,N_27999);
or U28368 (N_28368,N_27158,N_27003);
and U28369 (N_28369,N_27622,N_27327);
nor U28370 (N_28370,N_27948,N_27862);
or U28371 (N_28371,N_27635,N_27109);
xor U28372 (N_28372,N_27353,N_27926);
xnor U28373 (N_28373,N_27872,N_27434);
or U28374 (N_28374,N_27730,N_27494);
or U28375 (N_28375,N_27727,N_27360);
or U28376 (N_28376,N_27031,N_27293);
nand U28377 (N_28377,N_27165,N_27808);
and U28378 (N_28378,N_27151,N_27275);
nor U28379 (N_28379,N_27213,N_27880);
xnor U28380 (N_28380,N_27822,N_27840);
or U28381 (N_28381,N_27640,N_27363);
xor U28382 (N_28382,N_27396,N_27349);
nand U28383 (N_28383,N_27780,N_27443);
or U28384 (N_28384,N_27806,N_27339);
and U28385 (N_28385,N_27468,N_27390);
xnor U28386 (N_28386,N_27582,N_27564);
nor U28387 (N_28387,N_27150,N_27529);
nor U28388 (N_28388,N_27977,N_27799);
or U28389 (N_28389,N_27953,N_27077);
nor U28390 (N_28390,N_27695,N_27810);
and U28391 (N_28391,N_27208,N_27084);
or U28392 (N_28392,N_27998,N_27954);
nor U28393 (N_28393,N_27232,N_27536);
or U28394 (N_28394,N_27600,N_27534);
xnor U28395 (N_28395,N_27194,N_27519);
nand U28396 (N_28396,N_27853,N_27267);
or U28397 (N_28397,N_27938,N_27931);
and U28398 (N_28398,N_27464,N_27651);
xor U28399 (N_28399,N_27436,N_27278);
and U28400 (N_28400,N_27696,N_27596);
xnor U28401 (N_28401,N_27040,N_27643);
or U28402 (N_28402,N_27767,N_27301);
nand U28403 (N_28403,N_27438,N_27665);
nor U28404 (N_28404,N_27190,N_27290);
and U28405 (N_28405,N_27630,N_27330);
nor U28406 (N_28406,N_27133,N_27156);
or U28407 (N_28407,N_27583,N_27344);
or U28408 (N_28408,N_27501,N_27831);
nand U28409 (N_28409,N_27473,N_27705);
and U28410 (N_28410,N_27662,N_27983);
or U28411 (N_28411,N_27291,N_27454);
nor U28412 (N_28412,N_27551,N_27751);
or U28413 (N_28413,N_27683,N_27110);
nand U28414 (N_28414,N_27927,N_27798);
and U28415 (N_28415,N_27934,N_27171);
or U28416 (N_28416,N_27916,N_27253);
nor U28417 (N_28417,N_27282,N_27399);
or U28418 (N_28418,N_27184,N_27459);
or U28419 (N_28419,N_27787,N_27457);
and U28420 (N_28420,N_27952,N_27338);
nor U28421 (N_28421,N_27664,N_27637);
and U28422 (N_28422,N_27897,N_27481);
or U28423 (N_28423,N_27512,N_27182);
and U28424 (N_28424,N_27597,N_27163);
nand U28425 (N_28425,N_27018,N_27638);
and U28426 (N_28426,N_27835,N_27516);
nor U28427 (N_28427,N_27524,N_27269);
xor U28428 (N_28428,N_27598,N_27736);
or U28429 (N_28429,N_27657,N_27259);
xor U28430 (N_28430,N_27420,N_27628);
and U28431 (N_28431,N_27168,N_27570);
or U28432 (N_28432,N_27395,N_27000);
nor U28433 (N_28433,N_27185,N_27656);
or U28434 (N_28434,N_27250,N_27319);
xor U28435 (N_28435,N_27732,N_27958);
nand U28436 (N_28436,N_27550,N_27528);
nand U28437 (N_28437,N_27669,N_27426);
nand U28438 (N_28438,N_27149,N_27318);
or U28439 (N_28439,N_27316,N_27425);
xor U28440 (N_28440,N_27430,N_27500);
xnor U28441 (N_28441,N_27857,N_27702);
and U28442 (N_28442,N_27072,N_27517);
nand U28443 (N_28443,N_27441,N_27029);
and U28444 (N_28444,N_27398,N_27350);
and U28445 (N_28445,N_27633,N_27949);
or U28446 (N_28446,N_27848,N_27066);
and U28447 (N_28447,N_27004,N_27011);
nand U28448 (N_28448,N_27505,N_27343);
or U28449 (N_28449,N_27636,N_27383);
nand U28450 (N_28450,N_27765,N_27196);
nand U28451 (N_28451,N_27471,N_27323);
nor U28452 (N_28452,N_27745,N_27148);
and U28453 (N_28453,N_27215,N_27593);
and U28454 (N_28454,N_27104,N_27961);
and U28455 (N_28455,N_27221,N_27781);
or U28456 (N_28456,N_27173,N_27421);
and U28457 (N_28457,N_27310,N_27543);
or U28458 (N_28458,N_27428,N_27676);
nand U28459 (N_28459,N_27035,N_27901);
and U28460 (N_28460,N_27790,N_27037);
nand U28461 (N_28461,N_27377,N_27863);
nor U28462 (N_28462,N_27647,N_27234);
nand U28463 (N_28463,N_27577,N_27276);
xor U28464 (N_28464,N_27351,N_27565);
xor U28465 (N_28465,N_27083,N_27830);
xor U28466 (N_28466,N_27532,N_27124);
and U28467 (N_28467,N_27717,N_27753);
xor U28468 (N_28468,N_27841,N_27760);
nand U28469 (N_28469,N_27144,N_27984);
or U28470 (N_28470,N_27599,N_27222);
xor U28471 (N_28471,N_27716,N_27920);
nor U28472 (N_28472,N_27495,N_27974);
nor U28473 (N_28473,N_27681,N_27107);
or U28474 (N_28474,N_27134,N_27959);
and U28475 (N_28475,N_27220,N_27447);
or U28476 (N_28476,N_27988,N_27601);
or U28477 (N_28477,N_27845,N_27260);
nand U28478 (N_28478,N_27621,N_27223);
nand U28479 (N_28479,N_27229,N_27277);
xnor U28480 (N_28480,N_27616,N_27779);
and U28481 (N_28481,N_27369,N_27198);
nand U28482 (N_28482,N_27951,N_27373);
nand U28483 (N_28483,N_27943,N_27406);
xor U28484 (N_28484,N_27479,N_27935);
or U28485 (N_28485,N_27930,N_27263);
xor U28486 (N_28486,N_27238,N_27137);
or U28487 (N_28487,N_27062,N_27147);
nand U28488 (N_28488,N_27924,N_27786);
xor U28489 (N_28489,N_27957,N_27866);
and U28490 (N_28490,N_27739,N_27402);
nor U28491 (N_28491,N_27005,N_27792);
xor U28492 (N_28492,N_27675,N_27770);
and U28493 (N_28493,N_27081,N_27093);
nand U28494 (N_28494,N_27199,N_27205);
nor U28495 (N_28495,N_27400,N_27967);
xor U28496 (N_28496,N_27604,N_27887);
and U28497 (N_28497,N_27566,N_27860);
and U28498 (N_28498,N_27956,N_27017);
and U28499 (N_28499,N_27688,N_27874);
and U28500 (N_28500,N_27859,N_27315);
or U28501 (N_28501,N_27065,N_27429);
xnor U28502 (N_28502,N_27503,N_27331);
nand U28503 (N_28503,N_27744,N_27468);
nand U28504 (N_28504,N_27696,N_27949);
and U28505 (N_28505,N_27916,N_27136);
or U28506 (N_28506,N_27567,N_27980);
nand U28507 (N_28507,N_27942,N_27100);
nor U28508 (N_28508,N_27878,N_27785);
and U28509 (N_28509,N_27597,N_27982);
and U28510 (N_28510,N_27495,N_27647);
xor U28511 (N_28511,N_27511,N_27590);
nand U28512 (N_28512,N_27391,N_27211);
nor U28513 (N_28513,N_27364,N_27814);
xnor U28514 (N_28514,N_27069,N_27819);
nor U28515 (N_28515,N_27165,N_27451);
and U28516 (N_28516,N_27336,N_27257);
nand U28517 (N_28517,N_27753,N_27601);
xor U28518 (N_28518,N_27169,N_27543);
nor U28519 (N_28519,N_27211,N_27547);
xor U28520 (N_28520,N_27650,N_27517);
and U28521 (N_28521,N_27089,N_27334);
or U28522 (N_28522,N_27292,N_27558);
xor U28523 (N_28523,N_27820,N_27694);
nor U28524 (N_28524,N_27882,N_27438);
nand U28525 (N_28525,N_27991,N_27064);
nor U28526 (N_28526,N_27502,N_27255);
nor U28527 (N_28527,N_27581,N_27084);
xnor U28528 (N_28528,N_27465,N_27895);
xor U28529 (N_28529,N_27533,N_27532);
or U28530 (N_28530,N_27452,N_27392);
and U28531 (N_28531,N_27082,N_27729);
nor U28532 (N_28532,N_27660,N_27178);
xnor U28533 (N_28533,N_27169,N_27854);
and U28534 (N_28534,N_27251,N_27854);
nand U28535 (N_28535,N_27490,N_27548);
nand U28536 (N_28536,N_27643,N_27817);
nor U28537 (N_28537,N_27380,N_27272);
or U28538 (N_28538,N_27826,N_27933);
nor U28539 (N_28539,N_27279,N_27738);
and U28540 (N_28540,N_27684,N_27835);
or U28541 (N_28541,N_27244,N_27069);
nor U28542 (N_28542,N_27698,N_27311);
and U28543 (N_28543,N_27281,N_27834);
xor U28544 (N_28544,N_27374,N_27683);
xor U28545 (N_28545,N_27469,N_27533);
and U28546 (N_28546,N_27915,N_27667);
or U28547 (N_28547,N_27261,N_27506);
nor U28548 (N_28548,N_27455,N_27583);
or U28549 (N_28549,N_27531,N_27058);
and U28550 (N_28550,N_27915,N_27446);
xnor U28551 (N_28551,N_27899,N_27796);
nor U28552 (N_28552,N_27207,N_27969);
and U28553 (N_28553,N_27697,N_27994);
and U28554 (N_28554,N_27762,N_27947);
or U28555 (N_28555,N_27430,N_27492);
nand U28556 (N_28556,N_27062,N_27024);
nand U28557 (N_28557,N_27255,N_27513);
or U28558 (N_28558,N_27588,N_27360);
and U28559 (N_28559,N_27798,N_27716);
xor U28560 (N_28560,N_27738,N_27668);
nand U28561 (N_28561,N_27725,N_27530);
xor U28562 (N_28562,N_27590,N_27058);
or U28563 (N_28563,N_27290,N_27588);
xor U28564 (N_28564,N_27694,N_27165);
and U28565 (N_28565,N_27181,N_27973);
and U28566 (N_28566,N_27701,N_27160);
nand U28567 (N_28567,N_27871,N_27920);
and U28568 (N_28568,N_27683,N_27233);
nand U28569 (N_28569,N_27173,N_27954);
and U28570 (N_28570,N_27081,N_27217);
xnor U28571 (N_28571,N_27759,N_27118);
xor U28572 (N_28572,N_27971,N_27448);
nor U28573 (N_28573,N_27655,N_27842);
nand U28574 (N_28574,N_27076,N_27151);
nand U28575 (N_28575,N_27968,N_27216);
or U28576 (N_28576,N_27528,N_27360);
or U28577 (N_28577,N_27077,N_27689);
and U28578 (N_28578,N_27729,N_27010);
xnor U28579 (N_28579,N_27398,N_27086);
xnor U28580 (N_28580,N_27326,N_27427);
nor U28581 (N_28581,N_27476,N_27834);
and U28582 (N_28582,N_27278,N_27627);
xnor U28583 (N_28583,N_27753,N_27705);
and U28584 (N_28584,N_27040,N_27215);
nand U28585 (N_28585,N_27591,N_27814);
nand U28586 (N_28586,N_27325,N_27891);
and U28587 (N_28587,N_27181,N_27982);
xor U28588 (N_28588,N_27162,N_27371);
and U28589 (N_28589,N_27187,N_27406);
xor U28590 (N_28590,N_27823,N_27095);
nand U28591 (N_28591,N_27491,N_27308);
xnor U28592 (N_28592,N_27021,N_27699);
nor U28593 (N_28593,N_27893,N_27643);
xor U28594 (N_28594,N_27370,N_27237);
or U28595 (N_28595,N_27647,N_27480);
nand U28596 (N_28596,N_27376,N_27871);
xor U28597 (N_28597,N_27883,N_27604);
nand U28598 (N_28598,N_27657,N_27222);
or U28599 (N_28599,N_27962,N_27417);
nand U28600 (N_28600,N_27326,N_27954);
xnor U28601 (N_28601,N_27373,N_27141);
or U28602 (N_28602,N_27643,N_27651);
and U28603 (N_28603,N_27293,N_27285);
and U28604 (N_28604,N_27389,N_27313);
or U28605 (N_28605,N_27163,N_27238);
or U28606 (N_28606,N_27305,N_27200);
nor U28607 (N_28607,N_27868,N_27917);
xnor U28608 (N_28608,N_27117,N_27086);
and U28609 (N_28609,N_27866,N_27721);
nor U28610 (N_28610,N_27652,N_27539);
nor U28611 (N_28611,N_27720,N_27263);
nor U28612 (N_28612,N_27644,N_27097);
xor U28613 (N_28613,N_27372,N_27595);
nor U28614 (N_28614,N_27018,N_27890);
nand U28615 (N_28615,N_27116,N_27608);
nor U28616 (N_28616,N_27222,N_27331);
or U28617 (N_28617,N_27956,N_27088);
or U28618 (N_28618,N_27541,N_27768);
nor U28619 (N_28619,N_27822,N_27541);
and U28620 (N_28620,N_27638,N_27955);
nor U28621 (N_28621,N_27735,N_27528);
xor U28622 (N_28622,N_27043,N_27341);
nand U28623 (N_28623,N_27787,N_27124);
and U28624 (N_28624,N_27319,N_27245);
and U28625 (N_28625,N_27016,N_27282);
nor U28626 (N_28626,N_27485,N_27960);
xor U28627 (N_28627,N_27356,N_27526);
xor U28628 (N_28628,N_27344,N_27677);
nor U28629 (N_28629,N_27801,N_27171);
xnor U28630 (N_28630,N_27212,N_27358);
xor U28631 (N_28631,N_27542,N_27401);
nand U28632 (N_28632,N_27399,N_27169);
and U28633 (N_28633,N_27145,N_27225);
nor U28634 (N_28634,N_27096,N_27322);
xor U28635 (N_28635,N_27376,N_27851);
xor U28636 (N_28636,N_27840,N_27343);
nor U28637 (N_28637,N_27740,N_27219);
and U28638 (N_28638,N_27405,N_27960);
and U28639 (N_28639,N_27445,N_27542);
nor U28640 (N_28640,N_27131,N_27550);
nand U28641 (N_28641,N_27031,N_27672);
nand U28642 (N_28642,N_27339,N_27561);
nand U28643 (N_28643,N_27142,N_27953);
nand U28644 (N_28644,N_27677,N_27060);
xnor U28645 (N_28645,N_27963,N_27983);
and U28646 (N_28646,N_27875,N_27307);
nor U28647 (N_28647,N_27504,N_27293);
nor U28648 (N_28648,N_27507,N_27963);
or U28649 (N_28649,N_27355,N_27552);
xor U28650 (N_28650,N_27994,N_27873);
nor U28651 (N_28651,N_27624,N_27275);
and U28652 (N_28652,N_27190,N_27956);
xnor U28653 (N_28653,N_27229,N_27934);
xnor U28654 (N_28654,N_27651,N_27576);
nor U28655 (N_28655,N_27183,N_27140);
nand U28656 (N_28656,N_27465,N_27980);
nor U28657 (N_28657,N_27086,N_27653);
xor U28658 (N_28658,N_27256,N_27144);
or U28659 (N_28659,N_27543,N_27407);
nand U28660 (N_28660,N_27103,N_27487);
nand U28661 (N_28661,N_27098,N_27102);
nor U28662 (N_28662,N_27759,N_27625);
nor U28663 (N_28663,N_27113,N_27442);
nor U28664 (N_28664,N_27977,N_27560);
nand U28665 (N_28665,N_27414,N_27281);
and U28666 (N_28666,N_27573,N_27771);
nor U28667 (N_28667,N_27452,N_27339);
nand U28668 (N_28668,N_27058,N_27178);
and U28669 (N_28669,N_27779,N_27447);
or U28670 (N_28670,N_27424,N_27833);
or U28671 (N_28671,N_27526,N_27832);
nor U28672 (N_28672,N_27672,N_27431);
or U28673 (N_28673,N_27891,N_27603);
xnor U28674 (N_28674,N_27595,N_27092);
nand U28675 (N_28675,N_27199,N_27214);
or U28676 (N_28676,N_27286,N_27479);
nand U28677 (N_28677,N_27700,N_27509);
or U28678 (N_28678,N_27764,N_27154);
xor U28679 (N_28679,N_27120,N_27984);
nand U28680 (N_28680,N_27000,N_27515);
and U28681 (N_28681,N_27380,N_27904);
xor U28682 (N_28682,N_27602,N_27673);
nor U28683 (N_28683,N_27441,N_27577);
and U28684 (N_28684,N_27038,N_27122);
nor U28685 (N_28685,N_27018,N_27654);
nor U28686 (N_28686,N_27600,N_27743);
or U28687 (N_28687,N_27722,N_27899);
and U28688 (N_28688,N_27551,N_27852);
and U28689 (N_28689,N_27760,N_27607);
nand U28690 (N_28690,N_27112,N_27867);
nor U28691 (N_28691,N_27064,N_27356);
nand U28692 (N_28692,N_27239,N_27761);
xor U28693 (N_28693,N_27496,N_27879);
nor U28694 (N_28694,N_27256,N_27529);
and U28695 (N_28695,N_27873,N_27329);
xor U28696 (N_28696,N_27461,N_27724);
nor U28697 (N_28697,N_27295,N_27152);
or U28698 (N_28698,N_27116,N_27364);
nor U28699 (N_28699,N_27264,N_27875);
nor U28700 (N_28700,N_27821,N_27975);
or U28701 (N_28701,N_27063,N_27247);
nor U28702 (N_28702,N_27894,N_27202);
nand U28703 (N_28703,N_27657,N_27543);
or U28704 (N_28704,N_27900,N_27066);
nand U28705 (N_28705,N_27161,N_27137);
or U28706 (N_28706,N_27415,N_27955);
nor U28707 (N_28707,N_27515,N_27479);
and U28708 (N_28708,N_27261,N_27113);
or U28709 (N_28709,N_27636,N_27117);
and U28710 (N_28710,N_27285,N_27454);
or U28711 (N_28711,N_27284,N_27031);
and U28712 (N_28712,N_27247,N_27642);
nand U28713 (N_28713,N_27469,N_27007);
nor U28714 (N_28714,N_27728,N_27267);
nor U28715 (N_28715,N_27957,N_27232);
and U28716 (N_28716,N_27434,N_27137);
nand U28717 (N_28717,N_27500,N_27663);
xnor U28718 (N_28718,N_27744,N_27415);
or U28719 (N_28719,N_27251,N_27933);
nand U28720 (N_28720,N_27749,N_27923);
nand U28721 (N_28721,N_27878,N_27158);
xnor U28722 (N_28722,N_27392,N_27079);
nor U28723 (N_28723,N_27784,N_27088);
and U28724 (N_28724,N_27916,N_27182);
nor U28725 (N_28725,N_27114,N_27828);
and U28726 (N_28726,N_27362,N_27878);
or U28727 (N_28727,N_27829,N_27153);
xnor U28728 (N_28728,N_27100,N_27075);
nand U28729 (N_28729,N_27363,N_27346);
and U28730 (N_28730,N_27393,N_27366);
nand U28731 (N_28731,N_27796,N_27505);
nor U28732 (N_28732,N_27515,N_27497);
or U28733 (N_28733,N_27025,N_27687);
and U28734 (N_28734,N_27298,N_27474);
nand U28735 (N_28735,N_27764,N_27256);
and U28736 (N_28736,N_27225,N_27315);
and U28737 (N_28737,N_27033,N_27381);
and U28738 (N_28738,N_27426,N_27990);
nand U28739 (N_28739,N_27928,N_27163);
xor U28740 (N_28740,N_27337,N_27299);
nand U28741 (N_28741,N_27785,N_27509);
or U28742 (N_28742,N_27300,N_27256);
and U28743 (N_28743,N_27349,N_27350);
nand U28744 (N_28744,N_27191,N_27385);
and U28745 (N_28745,N_27558,N_27801);
nand U28746 (N_28746,N_27873,N_27480);
nor U28747 (N_28747,N_27757,N_27088);
nand U28748 (N_28748,N_27358,N_27512);
nand U28749 (N_28749,N_27496,N_27750);
or U28750 (N_28750,N_27529,N_27907);
nand U28751 (N_28751,N_27349,N_27939);
and U28752 (N_28752,N_27063,N_27866);
nor U28753 (N_28753,N_27309,N_27649);
and U28754 (N_28754,N_27161,N_27609);
nand U28755 (N_28755,N_27269,N_27715);
and U28756 (N_28756,N_27198,N_27174);
nor U28757 (N_28757,N_27359,N_27396);
xor U28758 (N_28758,N_27102,N_27248);
nand U28759 (N_28759,N_27258,N_27543);
nand U28760 (N_28760,N_27793,N_27921);
xor U28761 (N_28761,N_27397,N_27092);
and U28762 (N_28762,N_27606,N_27266);
or U28763 (N_28763,N_27068,N_27273);
or U28764 (N_28764,N_27061,N_27674);
and U28765 (N_28765,N_27763,N_27080);
xnor U28766 (N_28766,N_27004,N_27860);
xor U28767 (N_28767,N_27305,N_27793);
and U28768 (N_28768,N_27471,N_27189);
and U28769 (N_28769,N_27794,N_27894);
nor U28770 (N_28770,N_27880,N_27651);
or U28771 (N_28771,N_27054,N_27480);
and U28772 (N_28772,N_27061,N_27691);
xor U28773 (N_28773,N_27125,N_27603);
and U28774 (N_28774,N_27522,N_27483);
and U28775 (N_28775,N_27586,N_27634);
nand U28776 (N_28776,N_27370,N_27700);
or U28777 (N_28777,N_27328,N_27931);
nor U28778 (N_28778,N_27559,N_27239);
nor U28779 (N_28779,N_27854,N_27009);
xnor U28780 (N_28780,N_27930,N_27375);
or U28781 (N_28781,N_27605,N_27282);
xnor U28782 (N_28782,N_27611,N_27397);
xnor U28783 (N_28783,N_27962,N_27924);
and U28784 (N_28784,N_27551,N_27304);
xnor U28785 (N_28785,N_27338,N_27770);
or U28786 (N_28786,N_27141,N_27462);
nand U28787 (N_28787,N_27322,N_27345);
nor U28788 (N_28788,N_27345,N_27348);
xnor U28789 (N_28789,N_27785,N_27581);
xnor U28790 (N_28790,N_27348,N_27603);
and U28791 (N_28791,N_27758,N_27844);
nand U28792 (N_28792,N_27043,N_27898);
nand U28793 (N_28793,N_27533,N_27415);
xnor U28794 (N_28794,N_27755,N_27637);
nand U28795 (N_28795,N_27548,N_27074);
nor U28796 (N_28796,N_27567,N_27713);
nand U28797 (N_28797,N_27539,N_27821);
nor U28798 (N_28798,N_27489,N_27815);
and U28799 (N_28799,N_27008,N_27935);
nor U28800 (N_28800,N_27764,N_27134);
nor U28801 (N_28801,N_27683,N_27204);
and U28802 (N_28802,N_27334,N_27551);
and U28803 (N_28803,N_27098,N_27970);
and U28804 (N_28804,N_27447,N_27412);
or U28805 (N_28805,N_27160,N_27209);
and U28806 (N_28806,N_27427,N_27422);
and U28807 (N_28807,N_27343,N_27451);
nand U28808 (N_28808,N_27377,N_27502);
xnor U28809 (N_28809,N_27397,N_27897);
nor U28810 (N_28810,N_27402,N_27786);
or U28811 (N_28811,N_27856,N_27061);
nor U28812 (N_28812,N_27930,N_27127);
xnor U28813 (N_28813,N_27195,N_27616);
or U28814 (N_28814,N_27574,N_27037);
xnor U28815 (N_28815,N_27751,N_27565);
and U28816 (N_28816,N_27045,N_27498);
or U28817 (N_28817,N_27618,N_27006);
nor U28818 (N_28818,N_27359,N_27111);
nand U28819 (N_28819,N_27531,N_27936);
and U28820 (N_28820,N_27644,N_27900);
and U28821 (N_28821,N_27989,N_27203);
xor U28822 (N_28822,N_27030,N_27021);
xor U28823 (N_28823,N_27564,N_27043);
and U28824 (N_28824,N_27787,N_27355);
and U28825 (N_28825,N_27483,N_27461);
and U28826 (N_28826,N_27134,N_27656);
xnor U28827 (N_28827,N_27453,N_27052);
xnor U28828 (N_28828,N_27410,N_27099);
xor U28829 (N_28829,N_27847,N_27712);
and U28830 (N_28830,N_27902,N_27976);
and U28831 (N_28831,N_27511,N_27648);
xor U28832 (N_28832,N_27008,N_27941);
or U28833 (N_28833,N_27822,N_27328);
or U28834 (N_28834,N_27552,N_27008);
and U28835 (N_28835,N_27700,N_27189);
or U28836 (N_28836,N_27830,N_27620);
and U28837 (N_28837,N_27830,N_27694);
nor U28838 (N_28838,N_27282,N_27777);
or U28839 (N_28839,N_27701,N_27950);
nand U28840 (N_28840,N_27698,N_27041);
or U28841 (N_28841,N_27199,N_27584);
nand U28842 (N_28842,N_27453,N_27676);
nor U28843 (N_28843,N_27837,N_27644);
nand U28844 (N_28844,N_27353,N_27706);
xor U28845 (N_28845,N_27615,N_27974);
nor U28846 (N_28846,N_27580,N_27240);
or U28847 (N_28847,N_27631,N_27183);
or U28848 (N_28848,N_27036,N_27555);
nor U28849 (N_28849,N_27126,N_27858);
and U28850 (N_28850,N_27254,N_27703);
nor U28851 (N_28851,N_27431,N_27683);
and U28852 (N_28852,N_27930,N_27447);
and U28853 (N_28853,N_27009,N_27665);
nand U28854 (N_28854,N_27580,N_27830);
xor U28855 (N_28855,N_27958,N_27512);
nand U28856 (N_28856,N_27964,N_27885);
nand U28857 (N_28857,N_27935,N_27826);
or U28858 (N_28858,N_27601,N_27740);
xnor U28859 (N_28859,N_27223,N_27591);
nor U28860 (N_28860,N_27459,N_27306);
nor U28861 (N_28861,N_27631,N_27751);
nand U28862 (N_28862,N_27319,N_27678);
nor U28863 (N_28863,N_27019,N_27051);
and U28864 (N_28864,N_27208,N_27380);
xor U28865 (N_28865,N_27621,N_27310);
xor U28866 (N_28866,N_27406,N_27504);
and U28867 (N_28867,N_27704,N_27125);
nor U28868 (N_28868,N_27991,N_27583);
nor U28869 (N_28869,N_27714,N_27040);
and U28870 (N_28870,N_27187,N_27396);
nand U28871 (N_28871,N_27738,N_27704);
or U28872 (N_28872,N_27825,N_27778);
nand U28873 (N_28873,N_27548,N_27058);
nor U28874 (N_28874,N_27288,N_27647);
xnor U28875 (N_28875,N_27970,N_27559);
xnor U28876 (N_28876,N_27221,N_27356);
nor U28877 (N_28877,N_27287,N_27512);
nor U28878 (N_28878,N_27765,N_27327);
nand U28879 (N_28879,N_27124,N_27856);
xnor U28880 (N_28880,N_27127,N_27828);
nor U28881 (N_28881,N_27371,N_27372);
or U28882 (N_28882,N_27491,N_27116);
and U28883 (N_28883,N_27652,N_27749);
or U28884 (N_28884,N_27815,N_27501);
or U28885 (N_28885,N_27098,N_27995);
nand U28886 (N_28886,N_27284,N_27167);
nand U28887 (N_28887,N_27239,N_27972);
or U28888 (N_28888,N_27394,N_27456);
nand U28889 (N_28889,N_27998,N_27462);
nor U28890 (N_28890,N_27814,N_27551);
nor U28891 (N_28891,N_27682,N_27022);
nor U28892 (N_28892,N_27805,N_27993);
xor U28893 (N_28893,N_27463,N_27462);
nor U28894 (N_28894,N_27094,N_27020);
or U28895 (N_28895,N_27079,N_27888);
xor U28896 (N_28896,N_27968,N_27485);
and U28897 (N_28897,N_27142,N_27026);
or U28898 (N_28898,N_27393,N_27704);
and U28899 (N_28899,N_27948,N_27916);
and U28900 (N_28900,N_27922,N_27240);
nand U28901 (N_28901,N_27485,N_27115);
xor U28902 (N_28902,N_27487,N_27924);
and U28903 (N_28903,N_27023,N_27396);
nand U28904 (N_28904,N_27991,N_27272);
xnor U28905 (N_28905,N_27249,N_27074);
nor U28906 (N_28906,N_27349,N_27723);
or U28907 (N_28907,N_27082,N_27084);
nor U28908 (N_28908,N_27310,N_27659);
and U28909 (N_28909,N_27395,N_27369);
nor U28910 (N_28910,N_27399,N_27941);
and U28911 (N_28911,N_27717,N_27810);
xnor U28912 (N_28912,N_27800,N_27607);
nand U28913 (N_28913,N_27885,N_27234);
xor U28914 (N_28914,N_27032,N_27687);
xnor U28915 (N_28915,N_27277,N_27518);
or U28916 (N_28916,N_27354,N_27670);
xor U28917 (N_28917,N_27267,N_27847);
xor U28918 (N_28918,N_27619,N_27427);
and U28919 (N_28919,N_27834,N_27818);
and U28920 (N_28920,N_27748,N_27200);
and U28921 (N_28921,N_27423,N_27045);
xor U28922 (N_28922,N_27708,N_27424);
xor U28923 (N_28923,N_27656,N_27699);
and U28924 (N_28924,N_27713,N_27198);
xnor U28925 (N_28925,N_27661,N_27031);
and U28926 (N_28926,N_27995,N_27492);
xor U28927 (N_28927,N_27086,N_27130);
xor U28928 (N_28928,N_27603,N_27772);
or U28929 (N_28929,N_27850,N_27017);
or U28930 (N_28930,N_27213,N_27398);
nor U28931 (N_28931,N_27684,N_27091);
xnor U28932 (N_28932,N_27126,N_27211);
and U28933 (N_28933,N_27965,N_27139);
nor U28934 (N_28934,N_27087,N_27666);
or U28935 (N_28935,N_27869,N_27251);
xor U28936 (N_28936,N_27877,N_27125);
nand U28937 (N_28937,N_27106,N_27656);
and U28938 (N_28938,N_27352,N_27686);
nor U28939 (N_28939,N_27458,N_27646);
xor U28940 (N_28940,N_27355,N_27198);
or U28941 (N_28941,N_27307,N_27531);
or U28942 (N_28942,N_27928,N_27670);
and U28943 (N_28943,N_27600,N_27343);
or U28944 (N_28944,N_27807,N_27488);
xnor U28945 (N_28945,N_27245,N_27183);
nor U28946 (N_28946,N_27695,N_27576);
nor U28947 (N_28947,N_27861,N_27397);
nor U28948 (N_28948,N_27048,N_27955);
xor U28949 (N_28949,N_27728,N_27112);
nand U28950 (N_28950,N_27666,N_27097);
and U28951 (N_28951,N_27039,N_27111);
and U28952 (N_28952,N_27559,N_27561);
and U28953 (N_28953,N_27946,N_27724);
nand U28954 (N_28954,N_27258,N_27644);
or U28955 (N_28955,N_27413,N_27934);
and U28956 (N_28956,N_27222,N_27714);
or U28957 (N_28957,N_27713,N_27092);
and U28958 (N_28958,N_27773,N_27968);
and U28959 (N_28959,N_27962,N_27817);
xor U28960 (N_28960,N_27949,N_27046);
nor U28961 (N_28961,N_27078,N_27712);
xnor U28962 (N_28962,N_27714,N_27943);
and U28963 (N_28963,N_27056,N_27300);
nand U28964 (N_28964,N_27732,N_27553);
nand U28965 (N_28965,N_27905,N_27174);
nor U28966 (N_28966,N_27226,N_27308);
nand U28967 (N_28967,N_27982,N_27323);
nor U28968 (N_28968,N_27628,N_27020);
nor U28969 (N_28969,N_27675,N_27185);
and U28970 (N_28970,N_27090,N_27862);
xnor U28971 (N_28971,N_27814,N_27506);
xor U28972 (N_28972,N_27643,N_27911);
xnor U28973 (N_28973,N_27602,N_27306);
nand U28974 (N_28974,N_27063,N_27205);
nor U28975 (N_28975,N_27077,N_27284);
nor U28976 (N_28976,N_27912,N_27398);
or U28977 (N_28977,N_27918,N_27965);
nand U28978 (N_28978,N_27041,N_27981);
nor U28979 (N_28979,N_27928,N_27152);
or U28980 (N_28980,N_27745,N_27468);
nand U28981 (N_28981,N_27343,N_27494);
and U28982 (N_28982,N_27325,N_27063);
xor U28983 (N_28983,N_27900,N_27578);
nor U28984 (N_28984,N_27469,N_27467);
nand U28985 (N_28985,N_27348,N_27550);
or U28986 (N_28986,N_27792,N_27896);
xnor U28987 (N_28987,N_27604,N_27849);
and U28988 (N_28988,N_27341,N_27959);
and U28989 (N_28989,N_27918,N_27915);
nor U28990 (N_28990,N_27516,N_27969);
and U28991 (N_28991,N_27397,N_27970);
xnor U28992 (N_28992,N_27748,N_27986);
or U28993 (N_28993,N_27479,N_27625);
or U28994 (N_28994,N_27000,N_27034);
nand U28995 (N_28995,N_27838,N_27006);
or U28996 (N_28996,N_27396,N_27752);
and U28997 (N_28997,N_27997,N_27560);
or U28998 (N_28998,N_27315,N_27696);
or U28999 (N_28999,N_27748,N_27822);
or U29000 (N_29000,N_28077,N_28976);
xnor U29001 (N_29001,N_28031,N_28904);
nand U29002 (N_29002,N_28241,N_28875);
nand U29003 (N_29003,N_28089,N_28217);
or U29004 (N_29004,N_28910,N_28826);
xnor U29005 (N_29005,N_28994,N_28026);
nand U29006 (N_29006,N_28638,N_28522);
nand U29007 (N_29007,N_28003,N_28810);
xnor U29008 (N_29008,N_28476,N_28289);
nand U29009 (N_29009,N_28788,N_28629);
nor U29010 (N_29010,N_28211,N_28943);
nand U29011 (N_29011,N_28283,N_28847);
nor U29012 (N_29012,N_28093,N_28667);
and U29013 (N_29013,N_28423,N_28070);
nand U29014 (N_29014,N_28563,N_28562);
xor U29015 (N_29015,N_28533,N_28059);
xnor U29016 (N_29016,N_28133,N_28959);
or U29017 (N_29017,N_28596,N_28650);
nor U29018 (N_29018,N_28416,N_28907);
or U29019 (N_29019,N_28671,N_28584);
or U29020 (N_29020,N_28891,N_28061);
xor U29021 (N_29021,N_28684,N_28484);
and U29022 (N_29022,N_28948,N_28090);
and U29023 (N_29023,N_28012,N_28102);
nor U29024 (N_29024,N_28431,N_28115);
or U29025 (N_29025,N_28420,N_28051);
xnor U29026 (N_29026,N_28570,N_28338);
and U29027 (N_29027,N_28621,N_28574);
xor U29028 (N_29028,N_28333,N_28183);
nand U29029 (N_29029,N_28571,N_28016);
nor U29030 (N_29030,N_28554,N_28421);
nor U29031 (N_29031,N_28354,N_28912);
nor U29032 (N_29032,N_28393,N_28256);
xnor U29033 (N_29033,N_28504,N_28259);
nor U29034 (N_29034,N_28634,N_28908);
and U29035 (N_29035,N_28855,N_28231);
nand U29036 (N_29036,N_28889,N_28772);
nand U29037 (N_29037,N_28770,N_28332);
nor U29038 (N_29038,N_28877,N_28940);
nand U29039 (N_29039,N_28326,N_28457);
nor U29040 (N_29040,N_28397,N_28378);
xor U29041 (N_29041,N_28730,N_28191);
or U29042 (N_29042,N_28148,N_28525);
or U29043 (N_29043,N_28180,N_28581);
and U29044 (N_29044,N_28185,N_28124);
xnor U29045 (N_29045,N_28456,N_28011);
nor U29046 (N_29046,N_28527,N_28021);
or U29047 (N_29047,N_28549,N_28695);
nand U29048 (N_29048,N_28654,N_28294);
or U29049 (N_29049,N_28560,N_28239);
nand U29050 (N_29050,N_28529,N_28376);
nor U29051 (N_29051,N_28194,N_28931);
nand U29052 (N_29052,N_28464,N_28744);
or U29053 (N_29053,N_28139,N_28727);
and U29054 (N_29054,N_28552,N_28900);
xnor U29055 (N_29055,N_28279,N_28780);
nand U29056 (N_29056,N_28215,N_28884);
and U29057 (N_29057,N_28822,N_28475);
xnor U29058 (N_29058,N_28761,N_28488);
xnor U29059 (N_29059,N_28843,N_28829);
xor U29060 (N_29060,N_28199,N_28415);
and U29061 (N_29061,N_28807,N_28756);
or U29062 (N_29062,N_28972,N_28656);
nor U29063 (N_29063,N_28374,N_28555);
or U29064 (N_29064,N_28508,N_28883);
nand U29065 (N_29065,N_28974,N_28127);
xor U29066 (N_29066,N_28930,N_28020);
nor U29067 (N_29067,N_28387,N_28144);
xor U29068 (N_29068,N_28251,N_28165);
xor U29069 (N_29069,N_28882,N_28379);
nand U29070 (N_29070,N_28334,N_28359);
nand U29071 (N_29071,N_28128,N_28921);
or U29072 (N_29072,N_28384,N_28938);
or U29073 (N_29073,N_28646,N_28499);
and U29074 (N_29074,N_28632,N_28500);
nand U29075 (N_29075,N_28116,N_28373);
and U29076 (N_29076,N_28966,N_28944);
xor U29077 (N_29077,N_28202,N_28121);
nor U29078 (N_29078,N_28773,N_28301);
and U29079 (N_29079,N_28842,N_28608);
xnor U29080 (N_29080,N_28543,N_28075);
nor U29081 (N_29081,N_28697,N_28742);
nand U29082 (N_29082,N_28542,N_28166);
or U29083 (N_29083,N_28960,N_28942);
or U29084 (N_29084,N_28518,N_28888);
or U29085 (N_29085,N_28794,N_28065);
and U29086 (N_29086,N_28107,N_28440);
nor U29087 (N_29087,N_28335,N_28098);
xor U29088 (N_29088,N_28811,N_28762);
and U29089 (N_29089,N_28273,N_28396);
or U29090 (N_29090,N_28964,N_28315);
xor U29091 (N_29091,N_28445,N_28685);
or U29092 (N_29092,N_28894,N_28443);
nand U29093 (N_29093,N_28517,N_28360);
or U29094 (N_29094,N_28028,N_28967);
and U29095 (N_29095,N_28899,N_28640);
nor U29096 (N_29096,N_28493,N_28222);
or U29097 (N_29097,N_28411,N_28749);
nor U29098 (N_29098,N_28019,N_28564);
nand U29099 (N_29099,N_28253,N_28268);
nand U29100 (N_29100,N_28796,N_28293);
and U29101 (N_29101,N_28758,N_28362);
and U29102 (N_29102,N_28696,N_28363);
xor U29103 (N_29103,N_28466,N_28419);
or U29104 (N_29104,N_28603,N_28598);
xor U29105 (N_29105,N_28680,N_28909);
nand U29106 (N_29106,N_28895,N_28663);
nand U29107 (N_29107,N_28108,N_28845);
or U29108 (N_29108,N_28274,N_28502);
nor U29109 (N_29109,N_28859,N_28665);
nand U29110 (N_29110,N_28862,N_28472);
nor U29111 (N_29111,N_28427,N_28062);
nor U29112 (N_29112,N_28911,N_28649);
xnor U29113 (N_29113,N_28590,N_28595);
xnor U29114 (N_29114,N_28186,N_28893);
and U29115 (N_29115,N_28833,N_28187);
nand U29116 (N_29116,N_28181,N_28519);
nor U29117 (N_29117,N_28804,N_28125);
nand U29118 (N_29118,N_28438,N_28080);
or U29119 (N_29119,N_28782,N_28439);
xnor U29120 (N_29120,N_28110,N_28470);
and U29121 (N_29121,N_28023,N_28970);
xor U29122 (N_29122,N_28870,N_28155);
and U29123 (N_29123,N_28715,N_28197);
nor U29124 (N_29124,N_28983,N_28903);
xor U29125 (N_29125,N_28666,N_28722);
xor U29126 (N_29126,N_28025,N_28099);
and U29127 (N_29127,N_28164,N_28325);
xnor U29128 (N_29128,N_28131,N_28004);
or U29129 (N_29129,N_28609,N_28731);
or U29130 (N_29130,N_28495,N_28006);
xnor U29131 (N_29131,N_28229,N_28798);
and U29132 (N_29132,N_28790,N_28138);
nor U29133 (N_29133,N_28896,N_28577);
nand U29134 (N_29134,N_28151,N_28204);
or U29135 (N_29135,N_28235,N_28515);
or U29136 (N_29136,N_28083,N_28069);
and U29137 (N_29137,N_28037,N_28856);
or U29138 (N_29138,N_28310,N_28612);
and U29139 (N_29139,N_28218,N_28914);
nand U29140 (N_29140,N_28364,N_28769);
nor U29141 (N_29141,N_28482,N_28838);
nor U29142 (N_29142,N_28447,N_28746);
and U29143 (N_29143,N_28986,N_28787);
nand U29144 (N_29144,N_28216,N_28147);
and U29145 (N_29145,N_28280,N_28477);
and U29146 (N_29146,N_28820,N_28965);
nor U29147 (N_29147,N_28192,N_28078);
nand U29148 (N_29148,N_28617,N_28648);
nor U29149 (N_29149,N_28361,N_28248);
nor U29150 (N_29150,N_28880,N_28161);
and U29151 (N_29151,N_28371,N_28481);
and U29152 (N_29152,N_28196,N_28342);
xnor U29153 (N_29153,N_28979,N_28568);
xnor U29154 (N_29154,N_28752,N_28206);
xor U29155 (N_29155,N_28536,N_28540);
or U29156 (N_29156,N_28669,N_28352);
xnor U29157 (N_29157,N_28072,N_28783);
xor U29158 (N_29158,N_28238,N_28436);
or U29159 (N_29159,N_28551,N_28945);
or U29160 (N_29160,N_28177,N_28048);
nand U29161 (N_29161,N_28823,N_28786);
or U29162 (N_29162,N_28002,N_28611);
and U29163 (N_29163,N_28316,N_28057);
or U29164 (N_29164,N_28084,N_28989);
and U29165 (N_29165,N_28813,N_28610);
and U29166 (N_29166,N_28998,N_28592);
nor U29167 (N_29167,N_28915,N_28614);
nand U29168 (N_29168,N_28835,N_28708);
nand U29169 (N_29169,N_28821,N_28840);
xnor U29170 (N_29170,N_28081,N_28693);
xor U29171 (N_29171,N_28027,N_28531);
and U29172 (N_29172,N_28729,N_28321);
xnor U29173 (N_29173,N_28045,N_28507);
or U29174 (N_29174,N_28626,N_28789);
nand U29175 (N_29175,N_28395,N_28692);
xor U29176 (N_29176,N_28444,N_28262);
xor U29177 (N_29177,N_28105,N_28628);
or U29178 (N_29178,N_28569,N_28633);
xor U29179 (N_29179,N_28721,N_28455);
nor U29180 (N_29180,N_28459,N_28819);
xor U29181 (N_29181,N_28463,N_28038);
nand U29182 (N_29182,N_28314,N_28996);
xnor U29183 (N_29183,N_28478,N_28732);
nor U29184 (N_29184,N_28936,N_28391);
and U29185 (N_29185,N_28890,N_28990);
nor U29186 (N_29186,N_28154,N_28160);
or U29187 (N_29187,N_28403,N_28818);
nor U29188 (N_29188,N_28828,N_28237);
nor U29189 (N_29189,N_28501,N_28451);
nand U29190 (N_29190,N_28267,N_28657);
nand U29191 (N_29191,N_28673,N_28600);
and U29192 (N_29192,N_28446,N_28625);
nand U29193 (N_29193,N_28358,N_28526);
xnor U29194 (N_29194,N_28257,N_28739);
and U29195 (N_29195,N_28349,N_28660);
and U29196 (N_29196,N_28997,N_28977);
xor U29197 (N_29197,N_28503,N_28547);
xnor U29198 (N_29198,N_28702,N_28348);
nor U29199 (N_29199,N_28042,N_28565);
or U29200 (N_29200,N_28954,N_28242);
xnor U29201 (N_29201,N_28001,N_28013);
nor U29202 (N_29202,N_28658,N_28897);
nand U29203 (N_29203,N_28506,N_28971);
nor U29204 (N_29204,N_28465,N_28771);
and U29205 (N_29205,N_28700,N_28973);
and U29206 (N_29206,N_28982,N_28035);
nand U29207 (N_29207,N_28291,N_28171);
nor U29208 (N_29208,N_28240,N_28869);
nand U29209 (N_29209,N_28462,N_28471);
and U29210 (N_29210,N_28193,N_28926);
and U29211 (N_29211,N_28987,N_28097);
and U29212 (N_29212,N_28760,N_28981);
nand U29213 (N_29213,N_28417,N_28946);
xor U29214 (N_29214,N_28801,N_28340);
and U29215 (N_29215,N_28249,N_28800);
nand U29216 (N_29216,N_28740,N_28489);
xnor U29217 (N_29217,N_28688,N_28430);
xor U29218 (N_29218,N_28227,N_28313);
xor U29219 (N_29219,N_28714,N_28641);
and U29220 (N_29220,N_28433,N_28132);
nor U29221 (N_29221,N_28765,N_28635);
or U29222 (N_29222,N_28824,N_28932);
xnor U29223 (N_29223,N_28486,N_28651);
nand U29224 (N_29224,N_28776,N_28246);
nor U29225 (N_29225,N_28033,N_28902);
nor U29226 (N_29226,N_28901,N_28143);
and U29227 (N_29227,N_28311,N_28661);
and U29228 (N_29228,N_28567,N_28831);
or U29229 (N_29229,N_28167,N_28873);
xor U29230 (N_29230,N_28343,N_28245);
xnor U29231 (N_29231,N_28631,N_28728);
and U29232 (N_29232,N_28599,N_28285);
nand U29233 (N_29233,N_28030,N_28425);
nand U29234 (N_29234,N_28520,N_28049);
nor U29235 (N_29235,N_28566,N_28054);
nand U29236 (N_29236,N_28345,N_28544);
or U29237 (N_29237,N_28919,N_28918);
xor U29238 (N_29238,N_28337,N_28136);
or U29239 (N_29239,N_28591,N_28292);
nand U29240 (N_29240,N_28350,N_28175);
nand U29241 (N_29241,N_28305,N_28985);
nand U29242 (N_29242,N_28705,N_28750);
or U29243 (N_29243,N_28975,N_28659);
nand U29244 (N_29244,N_28422,N_28734);
and U29245 (N_29245,N_28009,N_28830);
nand U29246 (N_29246,N_28468,N_28329);
nor U29247 (N_29247,N_28636,N_28513);
nand U29248 (N_29248,N_28169,N_28347);
nor U29249 (N_29249,N_28434,N_28219);
or U29250 (N_29250,N_28370,N_28432);
xnor U29251 (N_29251,N_28100,N_28587);
xnor U29252 (N_29252,N_28812,N_28939);
nand U29253 (N_29253,N_28955,N_28735);
xor U29254 (N_29254,N_28260,N_28140);
and U29255 (N_29255,N_28064,N_28137);
nor U29256 (N_29256,N_28763,N_28454);
nand U29257 (N_29257,N_28214,N_28920);
or U29258 (N_29258,N_28073,N_28718);
and U29259 (N_29259,N_28221,N_28528);
and U29260 (N_29260,N_28068,N_28353);
nor U29261 (N_29261,N_28043,N_28799);
and U29262 (N_29262,N_28809,N_28076);
nand U29263 (N_29263,N_28207,N_28679);
nand U29264 (N_29264,N_28887,N_28872);
xor U29265 (N_29265,N_28168,N_28159);
or U29266 (N_29266,N_28736,N_28441);
nand U29267 (N_29267,N_28173,N_28254);
nand U29268 (N_29268,N_28174,N_28586);
and U29269 (N_29269,N_28426,N_28923);
or U29270 (N_29270,N_28868,N_28530);
and U29271 (N_29271,N_28056,N_28546);
nor U29272 (N_29272,N_28510,N_28198);
nand U29273 (N_29273,N_28400,N_28953);
xor U29274 (N_29274,N_28392,N_28866);
xor U29275 (N_29275,N_28863,N_28929);
nor U29276 (N_29276,N_28613,N_28851);
nand U29277 (N_29277,N_28269,N_28233);
xnor U29278 (N_29278,N_28690,N_28230);
nor U29279 (N_29279,N_28178,N_28490);
nor U29280 (N_29280,N_28778,N_28505);
and U29281 (N_29281,N_28664,N_28272);
and U29282 (N_29282,N_28103,N_28548);
nor U29283 (N_29283,N_28791,N_28647);
or U29284 (N_29284,N_28244,N_28741);
nor U29285 (N_29285,N_28278,N_28858);
nand U29286 (N_29286,N_28309,N_28683);
nor U29287 (N_29287,N_28757,N_28123);
nor U29288 (N_29288,N_28119,N_28024);
xor U29289 (N_29289,N_28803,N_28336);
xor U29290 (N_29290,N_28879,N_28643);
xor U29291 (N_29291,N_28999,N_28738);
nand U29292 (N_29292,N_28748,N_28550);
nand U29293 (N_29293,N_28618,N_28355);
xor U29294 (N_29294,N_28594,N_28766);
and U29295 (N_29295,N_28220,N_28460);
and U29296 (N_29296,N_28898,N_28106);
xor U29297 (N_29297,N_28958,N_28067);
or U29298 (N_29298,N_28601,N_28947);
nor U29299 (N_29299,N_28492,N_28941);
nor U29300 (N_29300,N_28117,N_28827);
xnor U29301 (N_29301,N_28992,N_28817);
nor U29302 (N_29302,N_28346,N_28474);
nand U29303 (N_29303,N_28052,N_28935);
nor U29304 (N_29304,N_28096,N_28324);
xor U29305 (N_29305,N_28687,N_28113);
nor U29306 (N_29306,N_28952,N_28496);
nand U29307 (N_29307,N_28553,N_28327);
or U29308 (N_29308,N_28308,N_28356);
and U29309 (N_29309,N_28582,N_28545);
and U29310 (N_29310,N_28616,N_28114);
nand U29311 (N_29311,N_28226,N_28523);
xor U29312 (N_29312,N_28184,N_28825);
and U29313 (N_29313,N_28250,N_28878);
nand U29314 (N_29314,N_28968,N_28849);
xnor U29315 (N_29315,N_28322,N_28126);
or U29316 (N_29316,N_28389,N_28428);
or U29317 (N_29317,N_28271,N_28537);
nor U29318 (N_29318,N_28303,N_28699);
or U29319 (N_29319,N_28753,N_28644);
xor U29320 (N_29320,N_28754,N_28129);
nand U29321 (N_29321,N_28007,N_28717);
or U29322 (N_29322,N_28266,N_28892);
or U29323 (N_29323,N_28118,N_28320);
nand U29324 (N_29324,N_28710,N_28201);
nand U29325 (N_29325,N_28764,N_28864);
and U29326 (N_29326,N_28304,N_28706);
and U29327 (N_29327,N_28775,N_28082);
or U29328 (N_29328,N_28203,N_28086);
and U29329 (N_29329,N_28619,N_28120);
or U29330 (N_29330,N_28814,N_28145);
and U29331 (N_29331,N_28485,N_28158);
and U29332 (N_29332,N_28575,N_28176);
and U29333 (N_29333,N_28622,N_28276);
or U29334 (N_29334,N_28916,N_28055);
nor U29335 (N_29335,N_28281,N_28652);
nor U29336 (N_29336,N_28275,N_28190);
or U29337 (N_29337,N_28713,N_28319);
and U29338 (N_29338,N_28991,N_28010);
or U29339 (N_29339,N_28917,N_28725);
and U29340 (N_29340,N_28223,N_28607);
xor U29341 (N_29341,N_28341,N_28795);
or U29342 (N_29342,N_28934,N_28208);
nand U29343 (N_29343,N_28834,N_28745);
or U29344 (N_29344,N_28234,N_28576);
xor U29345 (N_29345,N_28212,N_28104);
xnor U29346 (N_29346,N_28409,N_28816);
or U29347 (N_29347,N_28405,N_28874);
xor U29348 (N_29348,N_28995,N_28228);
nand U29349 (N_29349,N_28993,N_28850);
nor U29350 (N_29350,N_28394,N_28861);
nor U29351 (N_29351,N_28297,N_28109);
and U29352 (N_29352,N_28146,N_28258);
nand U29353 (N_29353,N_28963,N_28841);
nor U29354 (N_29354,N_28593,N_28933);
and U29355 (N_29355,N_28534,N_28195);
or U29356 (N_29356,N_28719,N_28808);
nand U29357 (N_29357,N_28539,N_28302);
nand U29358 (N_29358,N_28385,N_28046);
nor U29359 (N_29359,N_28514,N_28142);
nand U29360 (N_29360,N_28284,N_28681);
nor U29361 (N_29361,N_28205,N_28905);
or U29362 (N_29362,N_28044,N_28282);
or U29363 (N_29363,N_28232,N_28662);
xor U29364 (N_29364,N_28922,N_28017);
nand U29365 (N_29365,N_28768,N_28060);
xnor U29366 (N_29366,N_28682,N_28881);
and U29367 (N_29367,N_28639,N_28642);
nor U29368 (N_29368,N_28367,N_28209);
nand U29369 (N_29369,N_28630,N_28802);
or U29370 (N_29370,N_28572,N_28704);
xor U29371 (N_29371,N_28264,N_28015);
nand U29372 (N_29372,N_28255,N_28295);
or U29373 (N_29373,N_28698,N_28511);
nor U29374 (N_29374,N_28413,N_28401);
nor U29375 (N_29375,N_28390,N_28053);
nor U29376 (N_29376,N_28694,N_28095);
xor U29377 (N_29377,N_28703,N_28779);
xnor U29378 (N_29378,N_28604,N_28627);
xor U29379 (N_29379,N_28837,N_28645);
nor U29380 (N_29380,N_28956,N_28743);
and U29381 (N_29381,N_28034,N_28668);
nand U29382 (N_29382,N_28388,N_28066);
nor U29383 (N_29383,N_28724,N_28767);
nor U29384 (N_29384,N_28461,N_28399);
nor U29385 (N_29385,N_28369,N_28263);
nand U29386 (N_29386,N_28759,N_28521);
nor U29387 (N_29387,N_28357,N_28000);
and U29388 (N_29388,N_28913,N_28094);
nand U29389 (N_29389,N_28793,N_28805);
xor U29390 (N_29390,N_28381,N_28398);
nor U29391 (N_29391,N_28236,N_28247);
nor U29392 (N_29392,N_28008,N_28134);
or U29393 (N_29393,N_28962,N_28050);
xor U29394 (N_29394,N_28298,N_28200);
and U29395 (N_29395,N_28130,N_28152);
and U29396 (N_29396,N_28224,N_28737);
nand U29397 (N_29397,N_28815,N_28330);
or U29398 (N_29398,N_28122,N_28135);
xnor U29399 (N_29399,N_28404,N_28848);
nand U29400 (N_29400,N_28323,N_28620);
nand U29401 (N_29401,N_28414,N_28453);
xnor U29402 (N_29402,N_28886,N_28516);
or U29403 (N_29403,N_28988,N_28984);
nor U29404 (N_29404,N_28844,N_28689);
and U29405 (N_29405,N_28210,N_28328);
xor U29406 (N_29406,N_28365,N_28605);
nand U29407 (N_29407,N_28382,N_28018);
nand U29408 (N_29408,N_28290,N_28491);
and U29409 (N_29409,N_28300,N_28344);
and U29410 (N_29410,N_28781,N_28961);
nor U29411 (N_29411,N_28836,N_28846);
xnor U29412 (N_29412,N_28871,N_28509);
xor U29413 (N_29413,N_28832,N_28951);
xor U29414 (N_29414,N_28747,N_28243);
nor U29415 (N_29415,N_28307,N_28318);
xor U29416 (N_29416,N_28150,N_28676);
nand U29417 (N_29417,N_28580,N_28265);
and U29418 (N_29418,N_28678,N_28296);
xor U29419 (N_29419,N_28597,N_28777);
xor U29420 (N_29420,N_28071,N_28860);
xor U29421 (N_29421,N_28408,N_28980);
and U29422 (N_29422,N_28189,N_28583);
xor U29423 (N_29423,N_28906,N_28458);
nand U29424 (N_29424,N_28418,N_28162);
nor U29425 (N_29425,N_28339,N_28467);
or U29426 (N_29426,N_28261,N_28558);
or U29427 (N_29427,N_28473,N_28172);
and U29428 (N_29428,N_28386,N_28853);
nand U29429 (N_29429,N_28733,N_28317);
or U29430 (N_29430,N_28410,N_28691);
xor U29431 (N_29431,N_28039,N_28573);
xnor U29432 (N_29432,N_28624,N_28448);
xnor U29433 (N_29433,N_28557,N_28366);
and U29434 (N_29434,N_28377,N_28774);
xnor U29435 (N_29435,N_28589,N_28375);
or U29436 (N_29436,N_28479,N_28494);
xor U29437 (N_29437,N_28559,N_28637);
nand U29438 (N_29438,N_28442,N_28925);
and U29439 (N_29439,N_28452,N_28927);
xnor U29440 (N_29440,N_28532,N_28412);
nor U29441 (N_29441,N_28351,N_28865);
or U29442 (N_29442,N_28579,N_28435);
nand U29443 (N_29443,N_28079,N_28924);
xor U29444 (N_29444,N_28036,N_28606);
nor U29445 (N_29445,N_28675,N_28074);
xor U29446 (N_29446,N_28857,N_28449);
xor U29447 (N_29447,N_28541,N_28653);
xnor U29448 (N_29448,N_28711,N_28270);
nand U29449 (N_29449,N_28372,N_28312);
nor U29450 (N_29450,N_28792,N_28538);
nand U29451 (N_29451,N_28085,N_28091);
xor U29452 (N_29452,N_28672,N_28111);
xor U29453 (N_29453,N_28029,N_28720);
and U29454 (N_29454,N_28402,N_28429);
and U29455 (N_29455,N_28885,N_28876);
xor U29456 (N_29456,N_28112,N_28022);
or U29457 (N_29457,N_28483,N_28286);
xor U29458 (N_29458,N_28040,N_28487);
nand U29459 (N_29459,N_28383,N_28707);
nor U29460 (N_29460,N_28852,N_28179);
nor U29461 (N_29461,N_28709,N_28153);
or U29462 (N_29462,N_28213,N_28969);
nand U29463 (N_29463,N_28623,N_28615);
or U29464 (N_29464,N_28677,N_28978);
nor U29465 (N_29465,N_28141,N_28784);
nor U29466 (N_29466,N_28380,N_28149);
xor U29467 (N_29467,N_28854,N_28407);
and U29468 (N_29468,N_28497,N_28670);
nor U29469 (N_29469,N_28032,N_28450);
nor U29470 (N_29470,N_28101,N_28188);
nand U29471 (N_29471,N_28712,N_28751);
and U29472 (N_29472,N_28928,N_28524);
nand U29473 (N_29473,N_28058,N_28087);
xnor U29474 (N_29474,N_28252,N_28163);
nand U29475 (N_29475,N_28437,N_28726);
nand U29476 (N_29476,N_28585,N_28041);
xor U29477 (N_29477,N_28588,N_28182);
nor U29478 (N_29478,N_28797,N_28170);
xnor U29479 (N_29479,N_28088,N_28331);
xor U29480 (N_29480,N_28287,N_28157);
xnor U29481 (N_29481,N_28716,N_28306);
xor U29482 (N_29482,N_28014,N_28674);
xnor U29483 (N_29483,N_28561,N_28655);
or U29484 (N_29484,N_28806,N_28701);
or U29485 (N_29485,N_28535,N_28047);
and U29486 (N_29486,N_28556,N_28480);
nor U29487 (N_29487,N_28424,N_28498);
or U29488 (N_29488,N_28950,N_28277);
or U29489 (N_29489,N_28602,N_28723);
or U29490 (N_29490,N_28785,N_28867);
nand U29491 (N_29491,N_28299,N_28225);
or U29492 (N_29492,N_28937,N_28839);
nor U29493 (N_29493,N_28578,N_28755);
and U29494 (N_29494,N_28949,N_28406);
nor U29495 (N_29495,N_28368,N_28469);
and U29496 (N_29496,N_28005,N_28512);
nor U29497 (N_29497,N_28063,N_28288);
xnor U29498 (N_29498,N_28686,N_28156);
nand U29499 (N_29499,N_28957,N_28092);
and U29500 (N_29500,N_28281,N_28766);
nand U29501 (N_29501,N_28007,N_28951);
nand U29502 (N_29502,N_28542,N_28523);
nor U29503 (N_29503,N_28562,N_28872);
xor U29504 (N_29504,N_28706,N_28561);
and U29505 (N_29505,N_28709,N_28027);
nor U29506 (N_29506,N_28129,N_28969);
nor U29507 (N_29507,N_28031,N_28554);
and U29508 (N_29508,N_28906,N_28374);
nand U29509 (N_29509,N_28655,N_28670);
nand U29510 (N_29510,N_28888,N_28970);
nand U29511 (N_29511,N_28330,N_28582);
nor U29512 (N_29512,N_28532,N_28492);
or U29513 (N_29513,N_28544,N_28867);
xor U29514 (N_29514,N_28031,N_28439);
and U29515 (N_29515,N_28750,N_28889);
or U29516 (N_29516,N_28866,N_28110);
or U29517 (N_29517,N_28149,N_28562);
xor U29518 (N_29518,N_28837,N_28086);
xor U29519 (N_29519,N_28156,N_28707);
xnor U29520 (N_29520,N_28130,N_28102);
xnor U29521 (N_29521,N_28990,N_28770);
nor U29522 (N_29522,N_28495,N_28749);
xnor U29523 (N_29523,N_28639,N_28500);
or U29524 (N_29524,N_28852,N_28876);
and U29525 (N_29525,N_28957,N_28963);
nor U29526 (N_29526,N_28481,N_28780);
nor U29527 (N_29527,N_28775,N_28524);
and U29528 (N_29528,N_28734,N_28022);
xnor U29529 (N_29529,N_28855,N_28851);
or U29530 (N_29530,N_28094,N_28207);
or U29531 (N_29531,N_28698,N_28244);
nor U29532 (N_29532,N_28932,N_28071);
nand U29533 (N_29533,N_28544,N_28187);
and U29534 (N_29534,N_28412,N_28293);
or U29535 (N_29535,N_28090,N_28539);
or U29536 (N_29536,N_28004,N_28047);
xor U29537 (N_29537,N_28410,N_28883);
nor U29538 (N_29538,N_28679,N_28227);
nand U29539 (N_29539,N_28137,N_28937);
nor U29540 (N_29540,N_28663,N_28014);
and U29541 (N_29541,N_28590,N_28094);
nor U29542 (N_29542,N_28102,N_28444);
xnor U29543 (N_29543,N_28331,N_28897);
or U29544 (N_29544,N_28539,N_28232);
or U29545 (N_29545,N_28862,N_28433);
nor U29546 (N_29546,N_28718,N_28672);
and U29547 (N_29547,N_28133,N_28530);
or U29548 (N_29548,N_28646,N_28638);
and U29549 (N_29549,N_28703,N_28504);
nand U29550 (N_29550,N_28687,N_28716);
nand U29551 (N_29551,N_28330,N_28041);
nand U29552 (N_29552,N_28498,N_28286);
nor U29553 (N_29553,N_28227,N_28997);
or U29554 (N_29554,N_28097,N_28029);
xnor U29555 (N_29555,N_28686,N_28689);
nor U29556 (N_29556,N_28749,N_28172);
and U29557 (N_29557,N_28606,N_28690);
or U29558 (N_29558,N_28976,N_28528);
nand U29559 (N_29559,N_28706,N_28158);
nand U29560 (N_29560,N_28727,N_28673);
xnor U29561 (N_29561,N_28817,N_28697);
and U29562 (N_29562,N_28910,N_28732);
nor U29563 (N_29563,N_28251,N_28824);
and U29564 (N_29564,N_28814,N_28012);
nand U29565 (N_29565,N_28788,N_28641);
nand U29566 (N_29566,N_28371,N_28715);
or U29567 (N_29567,N_28030,N_28062);
xor U29568 (N_29568,N_28995,N_28030);
and U29569 (N_29569,N_28037,N_28427);
and U29570 (N_29570,N_28226,N_28236);
nor U29571 (N_29571,N_28497,N_28186);
xor U29572 (N_29572,N_28087,N_28969);
nor U29573 (N_29573,N_28209,N_28388);
nand U29574 (N_29574,N_28834,N_28055);
nor U29575 (N_29575,N_28991,N_28203);
or U29576 (N_29576,N_28612,N_28053);
xnor U29577 (N_29577,N_28946,N_28415);
xor U29578 (N_29578,N_28128,N_28134);
or U29579 (N_29579,N_28860,N_28304);
or U29580 (N_29580,N_28530,N_28873);
or U29581 (N_29581,N_28073,N_28440);
and U29582 (N_29582,N_28187,N_28758);
and U29583 (N_29583,N_28428,N_28450);
or U29584 (N_29584,N_28774,N_28583);
or U29585 (N_29585,N_28281,N_28857);
and U29586 (N_29586,N_28734,N_28499);
or U29587 (N_29587,N_28023,N_28992);
xnor U29588 (N_29588,N_28659,N_28918);
or U29589 (N_29589,N_28966,N_28324);
and U29590 (N_29590,N_28528,N_28978);
nand U29591 (N_29591,N_28193,N_28713);
and U29592 (N_29592,N_28108,N_28317);
or U29593 (N_29593,N_28365,N_28440);
or U29594 (N_29594,N_28220,N_28619);
and U29595 (N_29595,N_28037,N_28943);
and U29596 (N_29596,N_28818,N_28408);
xnor U29597 (N_29597,N_28843,N_28600);
xor U29598 (N_29598,N_28221,N_28448);
or U29599 (N_29599,N_28358,N_28121);
nor U29600 (N_29600,N_28957,N_28914);
nor U29601 (N_29601,N_28365,N_28578);
and U29602 (N_29602,N_28727,N_28556);
xnor U29603 (N_29603,N_28516,N_28063);
or U29604 (N_29604,N_28333,N_28772);
and U29605 (N_29605,N_28318,N_28603);
nand U29606 (N_29606,N_28571,N_28557);
or U29607 (N_29607,N_28367,N_28773);
nand U29608 (N_29608,N_28608,N_28072);
or U29609 (N_29609,N_28034,N_28240);
xnor U29610 (N_29610,N_28666,N_28230);
xor U29611 (N_29611,N_28252,N_28733);
or U29612 (N_29612,N_28599,N_28382);
nor U29613 (N_29613,N_28057,N_28998);
nor U29614 (N_29614,N_28016,N_28481);
and U29615 (N_29615,N_28075,N_28620);
and U29616 (N_29616,N_28864,N_28562);
xnor U29617 (N_29617,N_28077,N_28665);
nor U29618 (N_29618,N_28977,N_28291);
nor U29619 (N_29619,N_28830,N_28960);
and U29620 (N_29620,N_28647,N_28380);
and U29621 (N_29621,N_28756,N_28702);
xor U29622 (N_29622,N_28918,N_28644);
nor U29623 (N_29623,N_28033,N_28885);
or U29624 (N_29624,N_28504,N_28938);
or U29625 (N_29625,N_28349,N_28871);
nand U29626 (N_29626,N_28153,N_28455);
nand U29627 (N_29627,N_28015,N_28895);
nand U29628 (N_29628,N_28121,N_28016);
xor U29629 (N_29629,N_28451,N_28566);
xnor U29630 (N_29630,N_28799,N_28828);
nand U29631 (N_29631,N_28543,N_28441);
xor U29632 (N_29632,N_28478,N_28598);
or U29633 (N_29633,N_28493,N_28994);
xor U29634 (N_29634,N_28589,N_28711);
or U29635 (N_29635,N_28671,N_28578);
nand U29636 (N_29636,N_28852,N_28698);
and U29637 (N_29637,N_28396,N_28506);
nand U29638 (N_29638,N_28868,N_28103);
nand U29639 (N_29639,N_28123,N_28662);
xnor U29640 (N_29640,N_28690,N_28857);
or U29641 (N_29641,N_28824,N_28004);
and U29642 (N_29642,N_28838,N_28303);
or U29643 (N_29643,N_28875,N_28214);
or U29644 (N_29644,N_28712,N_28671);
and U29645 (N_29645,N_28366,N_28928);
nand U29646 (N_29646,N_28090,N_28388);
nor U29647 (N_29647,N_28800,N_28928);
and U29648 (N_29648,N_28407,N_28341);
nor U29649 (N_29649,N_28028,N_28671);
nor U29650 (N_29650,N_28673,N_28367);
xor U29651 (N_29651,N_28754,N_28337);
nand U29652 (N_29652,N_28131,N_28143);
nor U29653 (N_29653,N_28519,N_28493);
xnor U29654 (N_29654,N_28817,N_28993);
nand U29655 (N_29655,N_28800,N_28427);
or U29656 (N_29656,N_28174,N_28257);
xnor U29657 (N_29657,N_28206,N_28904);
or U29658 (N_29658,N_28706,N_28732);
or U29659 (N_29659,N_28560,N_28131);
nand U29660 (N_29660,N_28396,N_28669);
or U29661 (N_29661,N_28560,N_28330);
nand U29662 (N_29662,N_28185,N_28036);
nor U29663 (N_29663,N_28827,N_28516);
nor U29664 (N_29664,N_28494,N_28781);
and U29665 (N_29665,N_28871,N_28715);
or U29666 (N_29666,N_28708,N_28072);
and U29667 (N_29667,N_28153,N_28136);
nand U29668 (N_29668,N_28841,N_28395);
or U29669 (N_29669,N_28436,N_28399);
and U29670 (N_29670,N_28704,N_28117);
and U29671 (N_29671,N_28640,N_28121);
nor U29672 (N_29672,N_28978,N_28325);
or U29673 (N_29673,N_28484,N_28491);
nand U29674 (N_29674,N_28677,N_28447);
nand U29675 (N_29675,N_28873,N_28177);
xnor U29676 (N_29676,N_28804,N_28173);
xor U29677 (N_29677,N_28588,N_28708);
and U29678 (N_29678,N_28620,N_28354);
xnor U29679 (N_29679,N_28060,N_28043);
xnor U29680 (N_29680,N_28429,N_28735);
xor U29681 (N_29681,N_28097,N_28983);
xor U29682 (N_29682,N_28008,N_28593);
nand U29683 (N_29683,N_28934,N_28043);
nand U29684 (N_29684,N_28450,N_28566);
nor U29685 (N_29685,N_28821,N_28393);
nor U29686 (N_29686,N_28349,N_28269);
nor U29687 (N_29687,N_28264,N_28435);
and U29688 (N_29688,N_28827,N_28195);
nor U29689 (N_29689,N_28343,N_28697);
nand U29690 (N_29690,N_28048,N_28971);
nand U29691 (N_29691,N_28639,N_28689);
or U29692 (N_29692,N_28846,N_28971);
xnor U29693 (N_29693,N_28800,N_28748);
nand U29694 (N_29694,N_28720,N_28902);
or U29695 (N_29695,N_28508,N_28131);
nor U29696 (N_29696,N_28759,N_28500);
nand U29697 (N_29697,N_28625,N_28199);
nor U29698 (N_29698,N_28975,N_28095);
xnor U29699 (N_29699,N_28932,N_28431);
nor U29700 (N_29700,N_28335,N_28021);
nand U29701 (N_29701,N_28029,N_28998);
nor U29702 (N_29702,N_28814,N_28953);
nand U29703 (N_29703,N_28151,N_28542);
and U29704 (N_29704,N_28136,N_28553);
and U29705 (N_29705,N_28274,N_28314);
xor U29706 (N_29706,N_28061,N_28804);
nand U29707 (N_29707,N_28564,N_28682);
nor U29708 (N_29708,N_28876,N_28088);
and U29709 (N_29709,N_28657,N_28265);
or U29710 (N_29710,N_28648,N_28786);
or U29711 (N_29711,N_28602,N_28382);
nand U29712 (N_29712,N_28087,N_28735);
or U29713 (N_29713,N_28541,N_28021);
and U29714 (N_29714,N_28639,N_28892);
nor U29715 (N_29715,N_28517,N_28042);
nor U29716 (N_29716,N_28486,N_28100);
nand U29717 (N_29717,N_28413,N_28858);
and U29718 (N_29718,N_28338,N_28351);
xor U29719 (N_29719,N_28589,N_28080);
and U29720 (N_29720,N_28908,N_28659);
nor U29721 (N_29721,N_28380,N_28582);
nand U29722 (N_29722,N_28064,N_28374);
and U29723 (N_29723,N_28831,N_28993);
xnor U29724 (N_29724,N_28050,N_28203);
or U29725 (N_29725,N_28584,N_28791);
and U29726 (N_29726,N_28584,N_28564);
xnor U29727 (N_29727,N_28218,N_28223);
and U29728 (N_29728,N_28655,N_28951);
nor U29729 (N_29729,N_28357,N_28324);
xor U29730 (N_29730,N_28592,N_28521);
nor U29731 (N_29731,N_28912,N_28169);
xnor U29732 (N_29732,N_28269,N_28035);
xnor U29733 (N_29733,N_28449,N_28393);
nand U29734 (N_29734,N_28851,N_28600);
nor U29735 (N_29735,N_28130,N_28516);
and U29736 (N_29736,N_28921,N_28328);
or U29737 (N_29737,N_28846,N_28804);
nor U29738 (N_29738,N_28433,N_28637);
nor U29739 (N_29739,N_28579,N_28764);
nand U29740 (N_29740,N_28065,N_28810);
and U29741 (N_29741,N_28491,N_28206);
or U29742 (N_29742,N_28182,N_28791);
nor U29743 (N_29743,N_28729,N_28335);
nor U29744 (N_29744,N_28620,N_28948);
or U29745 (N_29745,N_28391,N_28069);
nor U29746 (N_29746,N_28873,N_28789);
or U29747 (N_29747,N_28037,N_28922);
or U29748 (N_29748,N_28124,N_28437);
and U29749 (N_29749,N_28953,N_28330);
and U29750 (N_29750,N_28696,N_28044);
nor U29751 (N_29751,N_28241,N_28908);
or U29752 (N_29752,N_28414,N_28638);
nand U29753 (N_29753,N_28549,N_28929);
and U29754 (N_29754,N_28254,N_28163);
nor U29755 (N_29755,N_28991,N_28768);
and U29756 (N_29756,N_28905,N_28181);
and U29757 (N_29757,N_28253,N_28403);
nand U29758 (N_29758,N_28317,N_28826);
and U29759 (N_29759,N_28245,N_28623);
or U29760 (N_29760,N_28138,N_28294);
and U29761 (N_29761,N_28942,N_28248);
nor U29762 (N_29762,N_28454,N_28713);
nor U29763 (N_29763,N_28103,N_28475);
nor U29764 (N_29764,N_28446,N_28767);
or U29765 (N_29765,N_28331,N_28127);
nor U29766 (N_29766,N_28457,N_28607);
and U29767 (N_29767,N_28996,N_28232);
xor U29768 (N_29768,N_28623,N_28224);
or U29769 (N_29769,N_28541,N_28373);
or U29770 (N_29770,N_28858,N_28952);
nand U29771 (N_29771,N_28407,N_28725);
xor U29772 (N_29772,N_28706,N_28211);
nor U29773 (N_29773,N_28140,N_28826);
nor U29774 (N_29774,N_28039,N_28508);
or U29775 (N_29775,N_28505,N_28247);
and U29776 (N_29776,N_28746,N_28942);
xnor U29777 (N_29777,N_28309,N_28834);
nor U29778 (N_29778,N_28435,N_28526);
and U29779 (N_29779,N_28662,N_28590);
and U29780 (N_29780,N_28464,N_28891);
nand U29781 (N_29781,N_28577,N_28151);
xor U29782 (N_29782,N_28230,N_28775);
or U29783 (N_29783,N_28661,N_28196);
xor U29784 (N_29784,N_28809,N_28768);
nor U29785 (N_29785,N_28407,N_28837);
nor U29786 (N_29786,N_28081,N_28679);
and U29787 (N_29787,N_28945,N_28880);
nor U29788 (N_29788,N_28761,N_28269);
and U29789 (N_29789,N_28608,N_28010);
xor U29790 (N_29790,N_28632,N_28711);
nand U29791 (N_29791,N_28338,N_28814);
or U29792 (N_29792,N_28354,N_28471);
and U29793 (N_29793,N_28063,N_28313);
nor U29794 (N_29794,N_28103,N_28689);
nor U29795 (N_29795,N_28116,N_28510);
and U29796 (N_29796,N_28947,N_28711);
nor U29797 (N_29797,N_28033,N_28627);
and U29798 (N_29798,N_28946,N_28349);
and U29799 (N_29799,N_28081,N_28963);
nor U29800 (N_29800,N_28745,N_28146);
and U29801 (N_29801,N_28886,N_28342);
or U29802 (N_29802,N_28844,N_28627);
nor U29803 (N_29803,N_28125,N_28939);
or U29804 (N_29804,N_28732,N_28976);
xnor U29805 (N_29805,N_28216,N_28243);
and U29806 (N_29806,N_28605,N_28168);
nand U29807 (N_29807,N_28722,N_28006);
or U29808 (N_29808,N_28653,N_28315);
nand U29809 (N_29809,N_28327,N_28001);
xor U29810 (N_29810,N_28210,N_28515);
and U29811 (N_29811,N_28859,N_28593);
and U29812 (N_29812,N_28561,N_28012);
and U29813 (N_29813,N_28195,N_28570);
and U29814 (N_29814,N_28424,N_28369);
or U29815 (N_29815,N_28595,N_28627);
nor U29816 (N_29816,N_28870,N_28175);
or U29817 (N_29817,N_28829,N_28091);
xor U29818 (N_29818,N_28128,N_28866);
xor U29819 (N_29819,N_28649,N_28806);
nand U29820 (N_29820,N_28471,N_28792);
nand U29821 (N_29821,N_28545,N_28447);
xor U29822 (N_29822,N_28835,N_28807);
or U29823 (N_29823,N_28877,N_28891);
and U29824 (N_29824,N_28077,N_28746);
or U29825 (N_29825,N_28232,N_28951);
nand U29826 (N_29826,N_28075,N_28223);
or U29827 (N_29827,N_28932,N_28543);
xnor U29828 (N_29828,N_28606,N_28459);
and U29829 (N_29829,N_28763,N_28182);
and U29830 (N_29830,N_28846,N_28941);
or U29831 (N_29831,N_28170,N_28188);
nor U29832 (N_29832,N_28075,N_28261);
nor U29833 (N_29833,N_28743,N_28170);
nand U29834 (N_29834,N_28183,N_28878);
nor U29835 (N_29835,N_28671,N_28889);
or U29836 (N_29836,N_28546,N_28481);
and U29837 (N_29837,N_28749,N_28150);
or U29838 (N_29838,N_28777,N_28700);
xor U29839 (N_29839,N_28895,N_28353);
and U29840 (N_29840,N_28082,N_28162);
xor U29841 (N_29841,N_28868,N_28691);
nand U29842 (N_29842,N_28480,N_28205);
nand U29843 (N_29843,N_28617,N_28673);
or U29844 (N_29844,N_28249,N_28432);
xnor U29845 (N_29845,N_28013,N_28115);
xor U29846 (N_29846,N_28582,N_28086);
or U29847 (N_29847,N_28322,N_28436);
nand U29848 (N_29848,N_28120,N_28071);
nand U29849 (N_29849,N_28336,N_28988);
and U29850 (N_29850,N_28620,N_28113);
xor U29851 (N_29851,N_28312,N_28266);
and U29852 (N_29852,N_28870,N_28011);
nand U29853 (N_29853,N_28749,N_28540);
nand U29854 (N_29854,N_28226,N_28535);
nor U29855 (N_29855,N_28970,N_28034);
or U29856 (N_29856,N_28333,N_28812);
or U29857 (N_29857,N_28914,N_28972);
nand U29858 (N_29858,N_28635,N_28212);
nor U29859 (N_29859,N_28009,N_28996);
nor U29860 (N_29860,N_28234,N_28271);
nor U29861 (N_29861,N_28427,N_28064);
nor U29862 (N_29862,N_28695,N_28718);
xor U29863 (N_29863,N_28504,N_28544);
nand U29864 (N_29864,N_28149,N_28514);
nor U29865 (N_29865,N_28847,N_28792);
or U29866 (N_29866,N_28692,N_28156);
xor U29867 (N_29867,N_28091,N_28930);
and U29868 (N_29868,N_28936,N_28852);
xnor U29869 (N_29869,N_28864,N_28522);
nand U29870 (N_29870,N_28834,N_28000);
nor U29871 (N_29871,N_28633,N_28642);
nor U29872 (N_29872,N_28459,N_28443);
nand U29873 (N_29873,N_28075,N_28946);
and U29874 (N_29874,N_28530,N_28644);
and U29875 (N_29875,N_28043,N_28530);
or U29876 (N_29876,N_28710,N_28773);
and U29877 (N_29877,N_28393,N_28296);
nor U29878 (N_29878,N_28120,N_28154);
and U29879 (N_29879,N_28014,N_28508);
nand U29880 (N_29880,N_28721,N_28525);
nand U29881 (N_29881,N_28993,N_28406);
and U29882 (N_29882,N_28736,N_28240);
nand U29883 (N_29883,N_28317,N_28736);
or U29884 (N_29884,N_28924,N_28101);
or U29885 (N_29885,N_28594,N_28811);
nor U29886 (N_29886,N_28423,N_28688);
nor U29887 (N_29887,N_28864,N_28702);
nand U29888 (N_29888,N_28683,N_28965);
xnor U29889 (N_29889,N_28040,N_28126);
nand U29890 (N_29890,N_28159,N_28555);
xnor U29891 (N_29891,N_28745,N_28749);
nor U29892 (N_29892,N_28961,N_28504);
or U29893 (N_29893,N_28876,N_28954);
nand U29894 (N_29894,N_28342,N_28542);
and U29895 (N_29895,N_28672,N_28732);
or U29896 (N_29896,N_28482,N_28087);
xor U29897 (N_29897,N_28776,N_28420);
nand U29898 (N_29898,N_28405,N_28848);
nor U29899 (N_29899,N_28951,N_28554);
xnor U29900 (N_29900,N_28419,N_28434);
nor U29901 (N_29901,N_28022,N_28994);
nor U29902 (N_29902,N_28999,N_28074);
or U29903 (N_29903,N_28776,N_28568);
and U29904 (N_29904,N_28102,N_28378);
xor U29905 (N_29905,N_28434,N_28093);
and U29906 (N_29906,N_28714,N_28332);
nand U29907 (N_29907,N_28450,N_28121);
and U29908 (N_29908,N_28958,N_28910);
or U29909 (N_29909,N_28451,N_28704);
nand U29910 (N_29910,N_28071,N_28066);
nor U29911 (N_29911,N_28737,N_28938);
nand U29912 (N_29912,N_28593,N_28869);
nor U29913 (N_29913,N_28598,N_28408);
xor U29914 (N_29914,N_28453,N_28974);
nand U29915 (N_29915,N_28606,N_28852);
nor U29916 (N_29916,N_28091,N_28407);
nand U29917 (N_29917,N_28056,N_28470);
nand U29918 (N_29918,N_28083,N_28455);
nand U29919 (N_29919,N_28115,N_28593);
and U29920 (N_29920,N_28138,N_28278);
nor U29921 (N_29921,N_28944,N_28918);
nor U29922 (N_29922,N_28240,N_28518);
nor U29923 (N_29923,N_28113,N_28664);
xnor U29924 (N_29924,N_28745,N_28562);
nor U29925 (N_29925,N_28351,N_28115);
or U29926 (N_29926,N_28062,N_28059);
xor U29927 (N_29927,N_28966,N_28759);
nor U29928 (N_29928,N_28947,N_28987);
nor U29929 (N_29929,N_28277,N_28778);
xor U29930 (N_29930,N_28641,N_28766);
xor U29931 (N_29931,N_28516,N_28563);
xor U29932 (N_29932,N_28043,N_28052);
nor U29933 (N_29933,N_28391,N_28523);
nand U29934 (N_29934,N_28134,N_28605);
or U29935 (N_29935,N_28669,N_28107);
or U29936 (N_29936,N_28544,N_28602);
nand U29937 (N_29937,N_28623,N_28020);
xor U29938 (N_29938,N_28331,N_28007);
or U29939 (N_29939,N_28601,N_28336);
nor U29940 (N_29940,N_28590,N_28091);
nor U29941 (N_29941,N_28576,N_28966);
nand U29942 (N_29942,N_28748,N_28589);
xnor U29943 (N_29943,N_28942,N_28938);
xor U29944 (N_29944,N_28463,N_28465);
nor U29945 (N_29945,N_28146,N_28754);
or U29946 (N_29946,N_28568,N_28271);
nand U29947 (N_29947,N_28901,N_28680);
and U29948 (N_29948,N_28272,N_28171);
nor U29949 (N_29949,N_28983,N_28966);
and U29950 (N_29950,N_28979,N_28232);
nand U29951 (N_29951,N_28711,N_28933);
xnor U29952 (N_29952,N_28016,N_28363);
and U29953 (N_29953,N_28457,N_28927);
nor U29954 (N_29954,N_28993,N_28748);
xor U29955 (N_29955,N_28272,N_28636);
nor U29956 (N_29956,N_28831,N_28192);
and U29957 (N_29957,N_28229,N_28094);
xnor U29958 (N_29958,N_28130,N_28054);
and U29959 (N_29959,N_28403,N_28395);
xnor U29960 (N_29960,N_28922,N_28431);
nand U29961 (N_29961,N_28670,N_28783);
and U29962 (N_29962,N_28783,N_28288);
or U29963 (N_29963,N_28583,N_28687);
xnor U29964 (N_29964,N_28653,N_28613);
or U29965 (N_29965,N_28710,N_28592);
xnor U29966 (N_29966,N_28879,N_28191);
and U29967 (N_29967,N_28215,N_28668);
xnor U29968 (N_29968,N_28435,N_28897);
nand U29969 (N_29969,N_28859,N_28036);
and U29970 (N_29970,N_28538,N_28547);
nor U29971 (N_29971,N_28914,N_28839);
nor U29972 (N_29972,N_28977,N_28828);
and U29973 (N_29973,N_28174,N_28490);
or U29974 (N_29974,N_28263,N_28117);
and U29975 (N_29975,N_28174,N_28739);
nor U29976 (N_29976,N_28668,N_28949);
nand U29977 (N_29977,N_28160,N_28888);
nand U29978 (N_29978,N_28676,N_28037);
and U29979 (N_29979,N_28309,N_28884);
xor U29980 (N_29980,N_28336,N_28579);
or U29981 (N_29981,N_28529,N_28675);
and U29982 (N_29982,N_28060,N_28935);
nor U29983 (N_29983,N_28617,N_28710);
or U29984 (N_29984,N_28236,N_28857);
xnor U29985 (N_29985,N_28079,N_28020);
and U29986 (N_29986,N_28793,N_28777);
nor U29987 (N_29987,N_28601,N_28629);
and U29988 (N_29988,N_28584,N_28260);
or U29989 (N_29989,N_28313,N_28851);
nand U29990 (N_29990,N_28332,N_28181);
nand U29991 (N_29991,N_28286,N_28337);
nand U29992 (N_29992,N_28548,N_28255);
nor U29993 (N_29993,N_28557,N_28538);
nor U29994 (N_29994,N_28962,N_28393);
xor U29995 (N_29995,N_28458,N_28899);
or U29996 (N_29996,N_28939,N_28536);
or U29997 (N_29997,N_28855,N_28147);
or U29998 (N_29998,N_28574,N_28612);
xor U29999 (N_29999,N_28662,N_28441);
nor UO_0 (O_0,N_29385,N_29201);
or UO_1 (O_1,N_29244,N_29156);
nand UO_2 (O_2,N_29188,N_29184);
nand UO_3 (O_3,N_29087,N_29794);
xor UO_4 (O_4,N_29718,N_29799);
and UO_5 (O_5,N_29704,N_29935);
or UO_6 (O_6,N_29538,N_29822);
xnor UO_7 (O_7,N_29610,N_29532);
or UO_8 (O_8,N_29369,N_29120);
xor UO_9 (O_9,N_29068,N_29672);
nand UO_10 (O_10,N_29350,N_29435);
or UO_11 (O_11,N_29409,N_29906);
nand UO_12 (O_12,N_29119,N_29000);
xnor UO_13 (O_13,N_29050,N_29354);
xnor UO_14 (O_14,N_29142,N_29631);
or UO_15 (O_15,N_29203,N_29918);
nand UO_16 (O_16,N_29782,N_29242);
nor UO_17 (O_17,N_29079,N_29995);
and UO_18 (O_18,N_29828,N_29613);
or UO_19 (O_19,N_29544,N_29487);
nand UO_20 (O_20,N_29246,N_29753);
and UO_21 (O_21,N_29909,N_29829);
or UO_22 (O_22,N_29449,N_29167);
xor UO_23 (O_23,N_29980,N_29343);
nand UO_24 (O_24,N_29543,N_29023);
and UO_25 (O_25,N_29739,N_29571);
and UO_26 (O_26,N_29216,N_29611);
xor UO_27 (O_27,N_29910,N_29762);
nor UO_28 (O_28,N_29364,N_29045);
xnor UO_29 (O_29,N_29838,N_29197);
and UO_30 (O_30,N_29576,N_29312);
xnor UO_31 (O_31,N_29844,N_29735);
nand UO_32 (O_32,N_29225,N_29259);
nand UO_33 (O_33,N_29545,N_29671);
xor UO_34 (O_34,N_29027,N_29204);
nand UO_35 (O_35,N_29526,N_29057);
nor UO_36 (O_36,N_29490,N_29442);
xor UO_37 (O_37,N_29467,N_29626);
or UO_38 (O_38,N_29876,N_29491);
nor UO_39 (O_39,N_29726,N_29236);
and UO_40 (O_40,N_29265,N_29881);
nor UO_41 (O_41,N_29878,N_29560);
xor UO_42 (O_42,N_29701,N_29509);
nand UO_43 (O_43,N_29921,N_29306);
nand UO_44 (O_44,N_29984,N_29607);
nor UO_45 (O_45,N_29564,N_29378);
nand UO_46 (O_46,N_29417,N_29159);
xor UO_47 (O_47,N_29269,N_29714);
xnor UO_48 (O_48,N_29373,N_29473);
and UO_49 (O_49,N_29220,N_29933);
nor UO_50 (O_50,N_29934,N_29235);
or UO_51 (O_51,N_29664,N_29665);
nor UO_52 (O_52,N_29189,N_29334);
or UO_53 (O_53,N_29808,N_29796);
xnor UO_54 (O_54,N_29932,N_29697);
or UO_55 (O_55,N_29415,N_29929);
xnor UO_56 (O_56,N_29586,N_29508);
nor UO_57 (O_57,N_29317,N_29698);
or UO_58 (O_58,N_29699,N_29251);
or UO_59 (O_59,N_29541,N_29474);
or UO_60 (O_60,N_29195,N_29460);
nand UO_61 (O_61,N_29318,N_29107);
nor UO_62 (O_62,N_29919,N_29255);
or UO_63 (O_63,N_29049,N_29954);
nor UO_64 (O_64,N_29895,N_29622);
xor UO_65 (O_65,N_29103,N_29847);
and UO_66 (O_66,N_29992,N_29136);
or UO_67 (O_67,N_29951,N_29254);
xnor UO_68 (O_68,N_29835,N_29010);
nor UO_69 (O_69,N_29342,N_29732);
or UO_70 (O_70,N_29238,N_29507);
and UO_71 (O_71,N_29429,N_29810);
and UO_72 (O_72,N_29472,N_29897);
or UO_73 (O_73,N_29080,N_29192);
or UO_74 (O_74,N_29675,N_29521);
and UO_75 (O_75,N_29450,N_29754);
xnor UO_76 (O_76,N_29781,N_29695);
or UO_77 (O_77,N_29104,N_29553);
xor UO_78 (O_78,N_29258,N_29520);
or UO_79 (O_79,N_29076,N_29169);
nand UO_80 (O_80,N_29062,N_29958);
xor UO_81 (O_81,N_29061,N_29060);
and UO_82 (O_82,N_29670,N_29971);
nor UO_83 (O_83,N_29777,N_29466);
nand UO_84 (O_84,N_29879,N_29839);
or UO_85 (O_85,N_29964,N_29293);
and UO_86 (O_86,N_29431,N_29396);
xor UO_87 (O_87,N_29546,N_29639);
and UO_88 (O_88,N_29655,N_29166);
or UO_89 (O_89,N_29268,N_29232);
nor UO_90 (O_90,N_29091,N_29996);
or UO_91 (O_91,N_29619,N_29451);
or UO_92 (O_92,N_29746,N_29633);
nor UO_93 (O_93,N_29004,N_29733);
nor UO_94 (O_94,N_29021,N_29492);
and UO_95 (O_95,N_29848,N_29206);
nand UO_96 (O_96,N_29423,N_29355);
xnor UO_97 (O_97,N_29230,N_29444);
and UO_98 (O_98,N_29372,N_29960);
nor UO_99 (O_99,N_29406,N_29171);
xnor UO_100 (O_100,N_29748,N_29677);
nand UO_101 (O_101,N_29081,N_29755);
and UO_102 (O_102,N_29277,N_29574);
or UO_103 (O_103,N_29086,N_29055);
xor UO_104 (O_104,N_29016,N_29694);
nand UO_105 (O_105,N_29131,N_29617);
nor UO_106 (O_106,N_29005,N_29987);
xnor UO_107 (O_107,N_29551,N_29924);
or UO_108 (O_108,N_29809,N_29866);
and UO_109 (O_109,N_29529,N_29593);
or UO_110 (O_110,N_29801,N_29158);
nor UO_111 (O_111,N_29597,N_29180);
nand UO_112 (O_112,N_29757,N_29300);
and UO_113 (O_113,N_29437,N_29900);
nand UO_114 (O_114,N_29747,N_29273);
nor UO_115 (O_115,N_29124,N_29253);
xor UO_116 (O_116,N_29892,N_29123);
or UO_117 (O_117,N_29788,N_29448);
or UO_118 (O_118,N_29713,N_29302);
xnor UO_119 (O_119,N_29535,N_29191);
xor UO_120 (O_120,N_29994,N_29290);
nand UO_121 (O_121,N_29604,N_29074);
or UO_122 (O_122,N_29584,N_29630);
or UO_123 (O_123,N_29001,N_29547);
xor UO_124 (O_124,N_29920,N_29495);
and UO_125 (O_125,N_29820,N_29427);
nor UO_126 (O_126,N_29070,N_29646);
xor UO_127 (O_127,N_29562,N_29568);
nor UO_128 (O_128,N_29627,N_29245);
nand UO_129 (O_129,N_29684,N_29020);
or UO_130 (O_130,N_29834,N_29145);
and UO_131 (O_131,N_29861,N_29751);
nand UO_132 (O_132,N_29970,N_29744);
or UO_133 (O_133,N_29014,N_29149);
xor UO_134 (O_134,N_29727,N_29514);
nand UO_135 (O_135,N_29053,N_29217);
xor UO_136 (O_136,N_29653,N_29331);
or UO_137 (O_137,N_29615,N_29842);
or UO_138 (O_138,N_29375,N_29715);
and UO_139 (O_139,N_29286,N_29767);
nand UO_140 (O_140,N_29341,N_29802);
nand UO_141 (O_141,N_29982,N_29886);
and UO_142 (O_142,N_29497,N_29575);
nand UO_143 (O_143,N_29384,N_29457);
nor UO_144 (O_144,N_29849,N_29281);
and UO_145 (O_145,N_29193,N_29832);
xnor UO_146 (O_146,N_29038,N_29518);
and UO_147 (O_147,N_29634,N_29421);
or UO_148 (O_148,N_29445,N_29494);
xnor UO_149 (O_149,N_29374,N_29650);
nor UO_150 (O_150,N_29099,N_29291);
nand UO_151 (O_151,N_29882,N_29064);
and UO_152 (O_152,N_29931,N_29516);
nor UO_153 (O_153,N_29006,N_29168);
and UO_154 (O_154,N_29032,N_29309);
xnor UO_155 (O_155,N_29357,N_29654);
nand UO_156 (O_156,N_29395,N_29214);
or UO_157 (O_157,N_29303,N_29566);
and UO_158 (O_158,N_29267,N_29493);
nand UO_159 (O_159,N_29443,N_29322);
nor UO_160 (O_160,N_29824,N_29223);
xnor UO_161 (O_161,N_29552,N_29034);
nor UO_162 (O_162,N_29304,N_29307);
and UO_163 (O_163,N_29877,N_29563);
nand UO_164 (O_164,N_29326,N_29771);
nor UO_165 (O_165,N_29132,N_29738);
nor UO_166 (O_166,N_29690,N_29983);
or UO_167 (O_167,N_29094,N_29608);
nor UO_168 (O_168,N_29389,N_29390);
xnor UO_169 (O_169,N_29769,N_29948);
nand UO_170 (O_170,N_29843,N_29565);
xor UO_171 (O_171,N_29875,N_29452);
or UO_172 (O_172,N_29616,N_29815);
nor UO_173 (O_173,N_29764,N_29262);
nand UO_174 (O_174,N_29144,N_29531);
nand UO_175 (O_175,N_29807,N_29786);
and UO_176 (O_176,N_29187,N_29348);
or UO_177 (O_177,N_29862,N_29985);
nor UO_178 (O_178,N_29674,N_29219);
nor UO_179 (O_179,N_29336,N_29359);
and UO_180 (O_180,N_29414,N_29162);
or UO_181 (O_181,N_29972,N_29702);
xnor UO_182 (O_182,N_29202,N_29666);
and UO_183 (O_183,N_29779,N_29089);
or UO_184 (O_184,N_29105,N_29393);
and UO_185 (O_185,N_29656,N_29524);
or UO_186 (O_186,N_29661,N_29696);
nor UO_187 (O_187,N_29805,N_29205);
and UO_188 (O_188,N_29583,N_29248);
nor UO_189 (O_189,N_29856,N_29963);
xor UO_190 (O_190,N_29891,N_29092);
nand UO_191 (O_191,N_29555,N_29816);
or UO_192 (O_192,N_29383,N_29645);
and UO_193 (O_193,N_29352,N_29864);
xor UO_194 (O_194,N_29377,N_29917);
nor UO_195 (O_195,N_29629,N_29311);
and UO_196 (O_196,N_29595,N_29305);
nand UO_197 (O_197,N_29585,N_29030);
nand UO_198 (O_198,N_29231,N_29632);
nand UO_199 (O_199,N_29250,N_29228);
or UO_200 (O_200,N_29768,N_29871);
nand UO_201 (O_201,N_29425,N_29257);
xnor UO_202 (O_202,N_29109,N_29976);
and UO_203 (O_203,N_29082,N_29851);
or UO_204 (O_204,N_29209,N_29075);
nand UO_205 (O_205,N_29823,N_29922);
or UO_206 (O_206,N_29275,N_29537);
and UO_207 (O_207,N_29540,N_29837);
nand UO_208 (O_208,N_29519,N_29657);
nor UO_209 (O_209,N_29720,N_29182);
xnor UO_210 (O_210,N_29237,N_29048);
nor UO_211 (O_211,N_29459,N_29461);
xnor UO_212 (O_212,N_29707,N_29539);
or UO_213 (O_213,N_29424,N_29386);
nand UO_214 (O_214,N_29358,N_29040);
or UO_215 (O_215,N_29643,N_29037);
and UO_216 (O_216,N_29841,N_29763);
nand UO_217 (O_217,N_29914,N_29868);
nor UO_218 (O_218,N_29330,N_29590);
nor UO_219 (O_219,N_29637,N_29790);
nor UO_220 (O_220,N_29997,N_29436);
nand UO_221 (O_221,N_29140,N_29234);
nor UO_222 (O_222,N_29721,N_29949);
and UO_223 (O_223,N_29337,N_29432);
xnor UO_224 (O_224,N_29161,N_29722);
and UO_225 (O_225,N_29282,N_29101);
nand UO_226 (O_226,N_29153,N_29090);
nand UO_227 (O_227,N_29042,N_29335);
nor UO_228 (O_228,N_29458,N_29649);
xnor UO_229 (O_229,N_29798,N_29515);
xor UO_230 (O_230,N_29150,N_29941);
and UO_231 (O_231,N_29172,N_29088);
xor UO_232 (O_232,N_29405,N_29663);
or UO_233 (O_233,N_29527,N_29367);
or UO_234 (O_234,N_29190,N_29100);
or UO_235 (O_235,N_29957,N_29106);
nand UO_236 (O_236,N_29213,N_29511);
and UO_237 (O_237,N_29624,N_29003);
or UO_238 (O_238,N_29692,N_29712);
and UO_239 (O_239,N_29554,N_29410);
and UO_240 (O_240,N_29438,N_29199);
and UO_241 (O_241,N_29376,N_29365);
nor UO_242 (O_242,N_29469,N_29319);
nor UO_243 (O_243,N_29218,N_29827);
nor UO_244 (O_244,N_29709,N_29752);
or UO_245 (O_245,N_29969,N_29279);
nor UO_246 (O_246,N_29758,N_29464);
nor UO_247 (O_247,N_29513,N_29440);
xor UO_248 (O_248,N_29818,N_29381);
or UO_249 (O_249,N_29127,N_29271);
or UO_250 (O_250,N_29502,N_29737);
xor UO_251 (O_251,N_29859,N_29683);
nand UO_252 (O_252,N_29778,N_29623);
nand UO_253 (O_253,N_29394,N_29561);
nor UO_254 (O_254,N_29981,N_29679);
and UO_255 (O_255,N_29908,N_29940);
nor UO_256 (O_256,N_29484,N_29447);
and UO_257 (O_257,N_29635,N_29528);
xnor UO_258 (O_258,N_29078,N_29241);
nor UO_259 (O_259,N_29899,N_29453);
xnor UO_260 (O_260,N_29743,N_29356);
nand UO_261 (O_261,N_29719,N_29605);
or UO_262 (O_262,N_29146,N_29904);
and UO_263 (O_263,N_29239,N_29731);
or UO_264 (O_264,N_29852,N_29428);
nand UO_265 (O_265,N_29911,N_29887);
nor UO_266 (O_266,N_29860,N_29780);
xnor UO_267 (O_267,N_29155,N_29693);
and UO_268 (O_268,N_29783,N_29351);
and UO_269 (O_269,N_29893,N_29967);
xnor UO_270 (O_270,N_29789,N_29745);
xnor UO_271 (O_271,N_29229,N_29299);
xnor UO_272 (O_272,N_29681,N_29558);
nand UO_273 (O_273,N_29791,N_29361);
nand UO_274 (O_274,N_29470,N_29975);
or UO_275 (O_275,N_29569,N_29462);
or UO_276 (O_276,N_29134,N_29885);
xor UO_277 (O_277,N_29434,N_29112);
xnor UO_278 (O_278,N_29700,N_29803);
nor UO_279 (O_279,N_29488,N_29456);
and UO_280 (O_280,N_29125,N_29363);
nand UO_281 (O_281,N_29894,N_29121);
xnor UO_282 (O_282,N_29013,N_29750);
xor UO_283 (O_283,N_29974,N_29991);
nor UO_284 (O_284,N_29489,N_29108);
xnor UO_285 (O_285,N_29730,N_29135);
or UO_286 (O_286,N_29582,N_29111);
nand UO_287 (O_287,N_29669,N_29591);
xnor UO_288 (O_288,N_29380,N_29716);
or UO_289 (O_289,N_29194,N_29703);
xnor UO_290 (O_290,N_29196,N_29362);
and UO_291 (O_291,N_29797,N_29294);
or UO_292 (O_292,N_29198,N_29505);
xor UO_293 (O_293,N_29455,N_29705);
xnor UO_294 (O_294,N_29966,N_29599);
and UO_295 (O_295,N_29770,N_29734);
or UO_296 (O_296,N_29594,N_29051);
xor UO_297 (O_297,N_29784,N_29240);
and UO_298 (O_298,N_29179,N_29243);
xor UO_299 (O_299,N_29990,N_29479);
xnor UO_300 (O_300,N_29641,N_29402);
nor UO_301 (O_301,N_29164,N_29295);
nand UO_302 (O_302,N_29017,N_29308);
and UO_303 (O_303,N_29333,N_29298);
and UO_304 (O_304,N_29360,N_29706);
and UO_305 (O_305,N_29925,N_29927);
or UO_306 (O_306,N_29316,N_29041);
xor UO_307 (O_307,N_29533,N_29636);
nor UO_308 (O_308,N_29148,N_29058);
nand UO_309 (O_309,N_29612,N_29212);
or UO_310 (O_310,N_29072,N_29411);
nand UO_311 (O_311,N_29115,N_29329);
xor UO_312 (O_312,N_29071,N_29117);
and UO_313 (O_313,N_29077,N_29160);
xor UO_314 (O_314,N_29025,N_29039);
nor UO_315 (O_315,N_29471,N_29804);
nor UO_316 (O_316,N_29339,N_29313);
or UO_317 (O_317,N_29031,N_29478);
nor UO_318 (O_318,N_29603,N_29840);
xor UO_319 (O_319,N_29141,N_29338);
nand UO_320 (O_320,N_29542,N_29968);
and UO_321 (O_321,N_29181,N_29667);
xor UO_322 (O_322,N_29647,N_29600);
xnor UO_323 (O_323,N_29854,N_29648);
or UO_324 (O_324,N_29741,N_29913);
nor UO_325 (O_325,N_29717,N_29480);
and UO_326 (O_326,N_29019,N_29151);
xor UO_327 (O_327,N_29496,N_29178);
xnor UO_328 (O_328,N_29912,N_29157);
and UO_329 (O_329,N_29773,N_29403);
nand UO_330 (O_330,N_29143,N_29278);
or UO_331 (O_331,N_29930,N_29618);
and UO_332 (O_332,N_29662,N_29800);
xor UO_333 (O_333,N_29033,N_29602);
or UO_334 (O_334,N_29118,N_29280);
and UO_335 (O_335,N_29962,N_29978);
nand UO_336 (O_336,N_29126,N_29550);
nor UO_337 (O_337,N_29740,N_29430);
nand UO_338 (O_338,N_29468,N_29793);
nor UO_339 (O_339,N_29046,N_29486);
xnor UO_340 (O_340,N_29548,N_29128);
nor UO_341 (O_341,N_29956,N_29977);
or UO_342 (O_342,N_29907,N_29549);
nand UO_343 (O_343,N_29869,N_29400);
or UO_344 (O_344,N_29475,N_29073);
and UO_345 (O_345,N_29412,N_29578);
or UO_346 (O_346,N_29093,N_29408);
and UO_347 (O_347,N_29580,N_29742);
nand UO_348 (O_348,N_29523,N_29325);
nand UO_349 (O_349,N_29943,N_29708);
and UO_350 (O_350,N_29792,N_29512);
nor UO_351 (O_351,N_29283,N_29371);
xnor UO_352 (O_352,N_29266,N_29133);
nor UO_353 (O_353,N_29207,N_29441);
xor UO_354 (O_354,N_29353,N_29154);
nor UO_355 (O_355,N_29660,N_29501);
xor UO_356 (O_356,N_29130,N_29301);
nor UO_357 (O_357,N_29588,N_29297);
and UO_358 (O_358,N_29260,N_29573);
or UO_359 (O_359,N_29765,N_29836);
nand UO_360 (O_360,N_29853,N_29819);
nand UO_361 (O_361,N_29825,N_29296);
nor UO_362 (O_362,N_29270,N_29147);
xnor UO_363 (O_363,N_29211,N_29577);
nor UO_364 (O_364,N_29454,N_29939);
and UO_365 (O_365,N_29233,N_29688);
xor UO_366 (O_366,N_29397,N_29831);
or UO_367 (O_367,N_29926,N_29399);
nor UO_368 (O_368,N_29658,N_29676);
or UO_369 (O_369,N_29614,N_29936);
nor UO_370 (O_370,N_29022,N_29570);
xnor UO_371 (O_371,N_29938,N_29601);
xor UO_372 (O_372,N_29084,N_29098);
nand UO_373 (O_373,N_29056,N_29937);
or UO_374 (O_374,N_29596,N_29047);
xnor UO_375 (O_375,N_29002,N_29476);
and UO_376 (O_376,N_29059,N_29340);
xor UO_377 (O_377,N_29517,N_29830);
xnor UO_378 (O_378,N_29026,N_29606);
or UO_379 (O_379,N_29845,N_29500);
or UO_380 (O_380,N_29506,N_29401);
nor UO_381 (O_381,N_29973,N_29955);
nand UO_382 (O_382,N_29227,N_29723);
and UO_383 (O_383,N_29680,N_29678);
nand UO_384 (O_384,N_29986,N_29426);
xor UO_385 (O_385,N_29152,N_29775);
nor UO_386 (O_386,N_29776,N_29332);
xnor UO_387 (O_387,N_29012,N_29889);
and UO_388 (O_388,N_29256,N_29863);
xnor UO_389 (O_389,N_29884,N_29177);
xor UO_390 (O_390,N_29965,N_29640);
xnor UO_391 (O_391,N_29028,N_29224);
xor UO_392 (O_392,N_29961,N_29766);
or UO_393 (O_393,N_29264,N_29556);
or UO_394 (O_394,N_29621,N_29175);
and UO_395 (O_395,N_29817,N_29785);
nor UO_396 (O_396,N_29018,N_29756);
xor UO_397 (O_397,N_29867,N_29183);
nand UO_398 (O_398,N_29043,N_29952);
or UO_399 (O_399,N_29821,N_29221);
and UO_400 (O_400,N_29366,N_29054);
xor UO_401 (O_401,N_29903,N_29557);
nor UO_402 (O_402,N_29029,N_29905);
and UO_403 (O_403,N_29289,N_29418);
and UO_404 (O_404,N_29226,N_29287);
or UO_405 (O_405,N_29222,N_29525);
nor UO_406 (O_406,N_29063,N_29320);
nand UO_407 (O_407,N_29404,N_29208);
nor UO_408 (O_408,N_29463,N_29292);
or UO_409 (O_409,N_29083,N_29485);
xor UO_410 (O_410,N_29176,N_29498);
or UO_411 (O_411,N_29979,N_29483);
or UO_412 (O_412,N_29651,N_29883);
xnor UO_413 (O_413,N_29272,N_29944);
nor UO_414 (O_414,N_29873,N_29890);
and UO_415 (O_415,N_29953,N_29609);
and UO_416 (O_416,N_29686,N_29170);
nand UO_417 (O_417,N_29346,N_29587);
xnor UO_418 (O_418,N_29122,N_29185);
or UO_419 (O_419,N_29276,N_29249);
or UO_420 (O_420,N_29388,N_29814);
or UO_421 (O_421,N_29114,N_29247);
and UO_422 (O_422,N_29947,N_29035);
nand UO_423 (O_423,N_29252,N_29314);
and UO_424 (O_424,N_29638,N_29685);
and UO_425 (O_425,N_29044,N_29581);
nor UO_426 (O_426,N_29687,N_29999);
nand UO_427 (O_427,N_29067,N_29419);
and UO_428 (O_428,N_29285,N_29321);
nor UO_429 (O_429,N_29066,N_29481);
nor UO_430 (O_430,N_29065,N_29345);
xnor UO_431 (O_431,N_29888,N_29759);
nand UO_432 (O_432,N_29407,N_29422);
or UO_433 (O_433,N_29186,N_29116);
or UO_434 (O_434,N_29711,N_29096);
xor UO_435 (O_435,N_29477,N_29813);
and UO_436 (O_436,N_29379,N_29392);
xnor UO_437 (O_437,N_29902,N_29870);
xor UO_438 (O_438,N_29139,N_29668);
or UO_439 (O_439,N_29880,N_29261);
or UO_440 (O_440,N_29344,N_29811);
xor UO_441 (O_441,N_29642,N_29534);
xor UO_442 (O_442,N_29846,N_29567);
nor UO_443 (O_443,N_29673,N_29416);
xor UO_444 (O_444,N_29998,N_29138);
xnor UO_445 (O_445,N_29988,N_29774);
xor UO_446 (O_446,N_29598,N_29069);
nand UO_447 (O_447,N_29826,N_29787);
nand UO_448 (O_448,N_29812,N_29263);
xor UO_449 (O_449,N_29085,N_29689);
nor UO_450 (O_450,N_29446,N_29865);
nand UO_451 (O_451,N_29129,N_29760);
or UO_452 (O_452,N_29323,N_29433);
nor UO_453 (O_453,N_29368,N_29008);
or UO_454 (O_454,N_29009,N_29945);
nand UO_455 (O_455,N_29536,N_29011);
nand UO_456 (O_456,N_29928,N_29215);
nand UO_457 (O_457,N_29898,N_29439);
xor UO_458 (O_458,N_29901,N_29324);
nor UO_459 (O_459,N_29315,N_29310);
nand UO_460 (O_460,N_29620,N_29413);
nand UO_461 (O_461,N_29833,N_29095);
nand UO_462 (O_462,N_29288,N_29625);
nand UO_463 (O_463,N_29522,N_29200);
nor UO_464 (O_464,N_29959,N_29387);
xnor UO_465 (O_465,N_29857,N_29173);
and UO_466 (O_466,N_29391,N_29559);
and UO_467 (O_467,N_29328,N_29163);
xnor UO_468 (O_468,N_29465,N_29993);
or UO_469 (O_469,N_29682,N_29724);
nor UO_470 (O_470,N_29165,N_29174);
nand UO_471 (O_471,N_29659,N_29806);
xnor UO_472 (O_472,N_29015,N_29510);
nand UO_473 (O_473,N_29007,N_29284);
nand UO_474 (O_474,N_29710,N_29482);
nor UO_475 (O_475,N_29872,N_29896);
or UO_476 (O_476,N_29725,N_29736);
and UO_477 (O_477,N_29036,N_29728);
and UO_478 (O_478,N_29772,N_29097);
and UO_479 (O_479,N_29946,N_29858);
and UO_480 (O_480,N_29349,N_29024);
xor UO_481 (O_481,N_29110,N_29572);
nand UO_482 (O_482,N_29589,N_29102);
and UO_483 (O_483,N_29327,N_29989);
nand UO_484 (O_484,N_29644,N_29950);
nor UO_485 (O_485,N_29503,N_29691);
or UO_486 (O_486,N_29210,N_29592);
or UO_487 (O_487,N_29579,N_29855);
or UO_488 (O_488,N_29420,N_29628);
or UO_489 (O_489,N_29530,N_29761);
and UO_490 (O_490,N_29274,N_29504);
nor UO_491 (O_491,N_29749,N_29398);
or UO_492 (O_492,N_29137,N_29113);
or UO_493 (O_493,N_29347,N_29915);
nand UO_494 (O_494,N_29729,N_29942);
or UO_495 (O_495,N_29499,N_29382);
nand UO_496 (O_496,N_29370,N_29795);
nand UO_497 (O_497,N_29923,N_29916);
xnor UO_498 (O_498,N_29652,N_29850);
nand UO_499 (O_499,N_29052,N_29874);
and UO_500 (O_500,N_29188,N_29593);
nor UO_501 (O_501,N_29791,N_29260);
xor UO_502 (O_502,N_29120,N_29891);
nor UO_503 (O_503,N_29220,N_29848);
xnor UO_504 (O_504,N_29471,N_29058);
or UO_505 (O_505,N_29752,N_29616);
or UO_506 (O_506,N_29266,N_29565);
xnor UO_507 (O_507,N_29744,N_29131);
or UO_508 (O_508,N_29567,N_29587);
nand UO_509 (O_509,N_29245,N_29007);
and UO_510 (O_510,N_29268,N_29142);
nand UO_511 (O_511,N_29138,N_29317);
nor UO_512 (O_512,N_29035,N_29286);
or UO_513 (O_513,N_29041,N_29523);
and UO_514 (O_514,N_29519,N_29929);
and UO_515 (O_515,N_29878,N_29337);
and UO_516 (O_516,N_29699,N_29647);
and UO_517 (O_517,N_29098,N_29685);
and UO_518 (O_518,N_29878,N_29170);
and UO_519 (O_519,N_29914,N_29318);
and UO_520 (O_520,N_29533,N_29934);
xor UO_521 (O_521,N_29960,N_29078);
nor UO_522 (O_522,N_29250,N_29754);
nor UO_523 (O_523,N_29327,N_29812);
xor UO_524 (O_524,N_29310,N_29149);
or UO_525 (O_525,N_29923,N_29460);
xnor UO_526 (O_526,N_29410,N_29846);
or UO_527 (O_527,N_29714,N_29641);
or UO_528 (O_528,N_29174,N_29906);
and UO_529 (O_529,N_29204,N_29533);
nand UO_530 (O_530,N_29387,N_29216);
nor UO_531 (O_531,N_29930,N_29267);
nand UO_532 (O_532,N_29365,N_29287);
or UO_533 (O_533,N_29057,N_29574);
or UO_534 (O_534,N_29964,N_29412);
and UO_535 (O_535,N_29268,N_29431);
nand UO_536 (O_536,N_29184,N_29479);
nor UO_537 (O_537,N_29943,N_29807);
and UO_538 (O_538,N_29702,N_29394);
nor UO_539 (O_539,N_29246,N_29496);
xnor UO_540 (O_540,N_29287,N_29449);
and UO_541 (O_541,N_29265,N_29604);
xnor UO_542 (O_542,N_29141,N_29410);
nand UO_543 (O_543,N_29639,N_29672);
nor UO_544 (O_544,N_29197,N_29914);
xor UO_545 (O_545,N_29945,N_29066);
or UO_546 (O_546,N_29719,N_29033);
or UO_547 (O_547,N_29910,N_29291);
and UO_548 (O_548,N_29316,N_29490);
xnor UO_549 (O_549,N_29573,N_29047);
or UO_550 (O_550,N_29612,N_29249);
nor UO_551 (O_551,N_29009,N_29704);
or UO_552 (O_552,N_29087,N_29535);
or UO_553 (O_553,N_29612,N_29211);
nor UO_554 (O_554,N_29475,N_29925);
xor UO_555 (O_555,N_29963,N_29554);
nand UO_556 (O_556,N_29153,N_29704);
nor UO_557 (O_557,N_29126,N_29559);
nand UO_558 (O_558,N_29330,N_29989);
nand UO_559 (O_559,N_29128,N_29261);
and UO_560 (O_560,N_29295,N_29887);
or UO_561 (O_561,N_29505,N_29436);
xor UO_562 (O_562,N_29719,N_29738);
xor UO_563 (O_563,N_29197,N_29998);
or UO_564 (O_564,N_29256,N_29211);
xor UO_565 (O_565,N_29280,N_29570);
nor UO_566 (O_566,N_29850,N_29346);
nand UO_567 (O_567,N_29654,N_29460);
nand UO_568 (O_568,N_29130,N_29892);
and UO_569 (O_569,N_29871,N_29738);
xor UO_570 (O_570,N_29424,N_29915);
xnor UO_571 (O_571,N_29611,N_29324);
nand UO_572 (O_572,N_29981,N_29494);
or UO_573 (O_573,N_29815,N_29835);
and UO_574 (O_574,N_29488,N_29714);
and UO_575 (O_575,N_29004,N_29395);
xnor UO_576 (O_576,N_29696,N_29986);
xor UO_577 (O_577,N_29291,N_29629);
or UO_578 (O_578,N_29003,N_29087);
or UO_579 (O_579,N_29967,N_29882);
nor UO_580 (O_580,N_29328,N_29139);
or UO_581 (O_581,N_29985,N_29854);
or UO_582 (O_582,N_29444,N_29434);
or UO_583 (O_583,N_29056,N_29258);
and UO_584 (O_584,N_29808,N_29415);
nand UO_585 (O_585,N_29762,N_29474);
and UO_586 (O_586,N_29476,N_29640);
and UO_587 (O_587,N_29622,N_29435);
xnor UO_588 (O_588,N_29622,N_29060);
and UO_589 (O_589,N_29113,N_29950);
nor UO_590 (O_590,N_29971,N_29067);
xor UO_591 (O_591,N_29532,N_29913);
and UO_592 (O_592,N_29315,N_29887);
or UO_593 (O_593,N_29980,N_29529);
or UO_594 (O_594,N_29505,N_29517);
xnor UO_595 (O_595,N_29196,N_29063);
nor UO_596 (O_596,N_29643,N_29203);
nor UO_597 (O_597,N_29140,N_29797);
or UO_598 (O_598,N_29982,N_29498);
and UO_599 (O_599,N_29995,N_29774);
and UO_600 (O_600,N_29846,N_29916);
xnor UO_601 (O_601,N_29725,N_29505);
nand UO_602 (O_602,N_29035,N_29645);
and UO_603 (O_603,N_29990,N_29427);
nor UO_604 (O_604,N_29849,N_29436);
nand UO_605 (O_605,N_29189,N_29548);
nand UO_606 (O_606,N_29632,N_29249);
nand UO_607 (O_607,N_29400,N_29990);
or UO_608 (O_608,N_29478,N_29699);
nand UO_609 (O_609,N_29220,N_29638);
and UO_610 (O_610,N_29766,N_29612);
nor UO_611 (O_611,N_29699,N_29337);
nor UO_612 (O_612,N_29708,N_29915);
and UO_613 (O_613,N_29242,N_29008);
or UO_614 (O_614,N_29034,N_29423);
and UO_615 (O_615,N_29693,N_29395);
xnor UO_616 (O_616,N_29601,N_29814);
or UO_617 (O_617,N_29087,N_29232);
xnor UO_618 (O_618,N_29670,N_29606);
and UO_619 (O_619,N_29219,N_29334);
or UO_620 (O_620,N_29562,N_29432);
nand UO_621 (O_621,N_29409,N_29785);
or UO_622 (O_622,N_29204,N_29349);
nor UO_623 (O_623,N_29057,N_29691);
xnor UO_624 (O_624,N_29779,N_29459);
nand UO_625 (O_625,N_29420,N_29860);
and UO_626 (O_626,N_29133,N_29017);
or UO_627 (O_627,N_29479,N_29509);
and UO_628 (O_628,N_29785,N_29404);
or UO_629 (O_629,N_29406,N_29477);
and UO_630 (O_630,N_29447,N_29054);
nor UO_631 (O_631,N_29543,N_29345);
and UO_632 (O_632,N_29962,N_29049);
nand UO_633 (O_633,N_29729,N_29971);
nor UO_634 (O_634,N_29535,N_29101);
nand UO_635 (O_635,N_29583,N_29001);
nor UO_636 (O_636,N_29948,N_29190);
xor UO_637 (O_637,N_29881,N_29478);
nand UO_638 (O_638,N_29588,N_29804);
and UO_639 (O_639,N_29746,N_29972);
or UO_640 (O_640,N_29607,N_29020);
and UO_641 (O_641,N_29801,N_29932);
nor UO_642 (O_642,N_29687,N_29600);
or UO_643 (O_643,N_29098,N_29730);
or UO_644 (O_644,N_29413,N_29920);
xnor UO_645 (O_645,N_29716,N_29591);
nand UO_646 (O_646,N_29861,N_29316);
nand UO_647 (O_647,N_29455,N_29003);
or UO_648 (O_648,N_29627,N_29908);
xor UO_649 (O_649,N_29463,N_29433);
xnor UO_650 (O_650,N_29121,N_29748);
or UO_651 (O_651,N_29290,N_29631);
or UO_652 (O_652,N_29919,N_29009);
nor UO_653 (O_653,N_29412,N_29773);
nand UO_654 (O_654,N_29864,N_29446);
and UO_655 (O_655,N_29393,N_29303);
nor UO_656 (O_656,N_29704,N_29014);
and UO_657 (O_657,N_29216,N_29204);
nor UO_658 (O_658,N_29787,N_29389);
and UO_659 (O_659,N_29272,N_29132);
xnor UO_660 (O_660,N_29006,N_29542);
or UO_661 (O_661,N_29373,N_29457);
xor UO_662 (O_662,N_29946,N_29716);
and UO_663 (O_663,N_29941,N_29830);
nor UO_664 (O_664,N_29623,N_29207);
nor UO_665 (O_665,N_29228,N_29112);
nand UO_666 (O_666,N_29142,N_29330);
and UO_667 (O_667,N_29977,N_29242);
and UO_668 (O_668,N_29189,N_29208);
nand UO_669 (O_669,N_29890,N_29901);
nor UO_670 (O_670,N_29036,N_29974);
nand UO_671 (O_671,N_29374,N_29666);
xor UO_672 (O_672,N_29043,N_29935);
and UO_673 (O_673,N_29544,N_29111);
nor UO_674 (O_674,N_29841,N_29789);
nand UO_675 (O_675,N_29720,N_29360);
nor UO_676 (O_676,N_29468,N_29388);
and UO_677 (O_677,N_29030,N_29534);
xor UO_678 (O_678,N_29956,N_29715);
and UO_679 (O_679,N_29749,N_29957);
nand UO_680 (O_680,N_29362,N_29191);
xnor UO_681 (O_681,N_29712,N_29541);
and UO_682 (O_682,N_29146,N_29203);
and UO_683 (O_683,N_29621,N_29940);
and UO_684 (O_684,N_29472,N_29397);
nand UO_685 (O_685,N_29801,N_29392);
and UO_686 (O_686,N_29581,N_29968);
and UO_687 (O_687,N_29567,N_29806);
nor UO_688 (O_688,N_29306,N_29512);
nand UO_689 (O_689,N_29660,N_29991);
or UO_690 (O_690,N_29869,N_29963);
and UO_691 (O_691,N_29559,N_29330);
xnor UO_692 (O_692,N_29045,N_29285);
and UO_693 (O_693,N_29648,N_29871);
nor UO_694 (O_694,N_29515,N_29498);
or UO_695 (O_695,N_29118,N_29585);
nor UO_696 (O_696,N_29684,N_29034);
xor UO_697 (O_697,N_29566,N_29671);
nand UO_698 (O_698,N_29244,N_29762);
nor UO_699 (O_699,N_29443,N_29671);
or UO_700 (O_700,N_29777,N_29378);
nor UO_701 (O_701,N_29863,N_29027);
nand UO_702 (O_702,N_29980,N_29988);
nor UO_703 (O_703,N_29668,N_29082);
nand UO_704 (O_704,N_29220,N_29334);
or UO_705 (O_705,N_29532,N_29751);
or UO_706 (O_706,N_29443,N_29083);
nand UO_707 (O_707,N_29883,N_29499);
xor UO_708 (O_708,N_29270,N_29857);
and UO_709 (O_709,N_29662,N_29525);
xor UO_710 (O_710,N_29789,N_29254);
xor UO_711 (O_711,N_29324,N_29247);
xnor UO_712 (O_712,N_29556,N_29215);
xnor UO_713 (O_713,N_29513,N_29738);
and UO_714 (O_714,N_29321,N_29392);
and UO_715 (O_715,N_29081,N_29794);
or UO_716 (O_716,N_29739,N_29241);
and UO_717 (O_717,N_29921,N_29072);
nor UO_718 (O_718,N_29957,N_29652);
nor UO_719 (O_719,N_29133,N_29417);
nand UO_720 (O_720,N_29138,N_29723);
or UO_721 (O_721,N_29928,N_29420);
or UO_722 (O_722,N_29595,N_29546);
nand UO_723 (O_723,N_29151,N_29023);
nor UO_724 (O_724,N_29894,N_29505);
nand UO_725 (O_725,N_29023,N_29769);
nor UO_726 (O_726,N_29144,N_29173);
nor UO_727 (O_727,N_29529,N_29996);
and UO_728 (O_728,N_29392,N_29593);
nand UO_729 (O_729,N_29143,N_29305);
and UO_730 (O_730,N_29921,N_29366);
xnor UO_731 (O_731,N_29652,N_29591);
or UO_732 (O_732,N_29937,N_29347);
nor UO_733 (O_733,N_29275,N_29885);
and UO_734 (O_734,N_29922,N_29687);
nor UO_735 (O_735,N_29629,N_29020);
nand UO_736 (O_736,N_29479,N_29864);
nor UO_737 (O_737,N_29948,N_29524);
or UO_738 (O_738,N_29327,N_29960);
xnor UO_739 (O_739,N_29631,N_29820);
or UO_740 (O_740,N_29462,N_29524);
nor UO_741 (O_741,N_29739,N_29322);
and UO_742 (O_742,N_29244,N_29527);
xnor UO_743 (O_743,N_29948,N_29193);
and UO_744 (O_744,N_29962,N_29233);
nand UO_745 (O_745,N_29429,N_29944);
and UO_746 (O_746,N_29154,N_29007);
and UO_747 (O_747,N_29091,N_29599);
xnor UO_748 (O_748,N_29679,N_29200);
xor UO_749 (O_749,N_29027,N_29812);
xnor UO_750 (O_750,N_29084,N_29571);
or UO_751 (O_751,N_29720,N_29803);
xnor UO_752 (O_752,N_29144,N_29337);
nand UO_753 (O_753,N_29654,N_29743);
nor UO_754 (O_754,N_29253,N_29846);
nor UO_755 (O_755,N_29145,N_29930);
xor UO_756 (O_756,N_29537,N_29332);
nand UO_757 (O_757,N_29709,N_29178);
xnor UO_758 (O_758,N_29054,N_29657);
xnor UO_759 (O_759,N_29067,N_29590);
and UO_760 (O_760,N_29500,N_29066);
xnor UO_761 (O_761,N_29605,N_29234);
or UO_762 (O_762,N_29514,N_29313);
nand UO_763 (O_763,N_29718,N_29708);
xnor UO_764 (O_764,N_29800,N_29062);
nor UO_765 (O_765,N_29903,N_29955);
nand UO_766 (O_766,N_29790,N_29001);
and UO_767 (O_767,N_29063,N_29468);
or UO_768 (O_768,N_29407,N_29145);
or UO_769 (O_769,N_29590,N_29087);
or UO_770 (O_770,N_29679,N_29879);
and UO_771 (O_771,N_29720,N_29032);
nand UO_772 (O_772,N_29870,N_29931);
or UO_773 (O_773,N_29149,N_29327);
nor UO_774 (O_774,N_29823,N_29786);
or UO_775 (O_775,N_29844,N_29399);
and UO_776 (O_776,N_29621,N_29091);
nand UO_777 (O_777,N_29822,N_29630);
nand UO_778 (O_778,N_29408,N_29067);
nand UO_779 (O_779,N_29603,N_29711);
xnor UO_780 (O_780,N_29425,N_29903);
xor UO_781 (O_781,N_29303,N_29849);
or UO_782 (O_782,N_29518,N_29807);
or UO_783 (O_783,N_29671,N_29751);
nand UO_784 (O_784,N_29587,N_29069);
nor UO_785 (O_785,N_29256,N_29574);
and UO_786 (O_786,N_29443,N_29008);
and UO_787 (O_787,N_29557,N_29104);
or UO_788 (O_788,N_29594,N_29924);
and UO_789 (O_789,N_29755,N_29704);
or UO_790 (O_790,N_29274,N_29472);
nor UO_791 (O_791,N_29767,N_29807);
nand UO_792 (O_792,N_29710,N_29912);
nand UO_793 (O_793,N_29851,N_29146);
and UO_794 (O_794,N_29671,N_29982);
xor UO_795 (O_795,N_29252,N_29597);
nand UO_796 (O_796,N_29608,N_29199);
or UO_797 (O_797,N_29347,N_29262);
nand UO_798 (O_798,N_29812,N_29598);
or UO_799 (O_799,N_29479,N_29353);
or UO_800 (O_800,N_29494,N_29861);
xor UO_801 (O_801,N_29306,N_29421);
xor UO_802 (O_802,N_29829,N_29296);
xor UO_803 (O_803,N_29971,N_29049);
or UO_804 (O_804,N_29172,N_29545);
or UO_805 (O_805,N_29861,N_29341);
or UO_806 (O_806,N_29567,N_29324);
nand UO_807 (O_807,N_29439,N_29465);
nor UO_808 (O_808,N_29669,N_29439);
nor UO_809 (O_809,N_29581,N_29301);
or UO_810 (O_810,N_29684,N_29146);
nor UO_811 (O_811,N_29992,N_29174);
xor UO_812 (O_812,N_29818,N_29781);
nor UO_813 (O_813,N_29028,N_29189);
nor UO_814 (O_814,N_29046,N_29807);
xnor UO_815 (O_815,N_29660,N_29371);
nor UO_816 (O_816,N_29286,N_29280);
nand UO_817 (O_817,N_29885,N_29519);
nand UO_818 (O_818,N_29896,N_29959);
nand UO_819 (O_819,N_29528,N_29334);
and UO_820 (O_820,N_29438,N_29695);
nand UO_821 (O_821,N_29944,N_29189);
nor UO_822 (O_822,N_29964,N_29396);
nor UO_823 (O_823,N_29552,N_29043);
and UO_824 (O_824,N_29728,N_29998);
nor UO_825 (O_825,N_29528,N_29611);
and UO_826 (O_826,N_29614,N_29179);
or UO_827 (O_827,N_29132,N_29873);
nor UO_828 (O_828,N_29374,N_29204);
xor UO_829 (O_829,N_29385,N_29089);
nand UO_830 (O_830,N_29226,N_29761);
nand UO_831 (O_831,N_29321,N_29292);
nor UO_832 (O_832,N_29216,N_29745);
and UO_833 (O_833,N_29240,N_29535);
and UO_834 (O_834,N_29292,N_29521);
and UO_835 (O_835,N_29156,N_29487);
nand UO_836 (O_836,N_29341,N_29237);
xor UO_837 (O_837,N_29457,N_29672);
nor UO_838 (O_838,N_29832,N_29222);
nor UO_839 (O_839,N_29302,N_29095);
nor UO_840 (O_840,N_29458,N_29890);
xor UO_841 (O_841,N_29616,N_29493);
or UO_842 (O_842,N_29806,N_29542);
xnor UO_843 (O_843,N_29248,N_29856);
nand UO_844 (O_844,N_29676,N_29352);
nand UO_845 (O_845,N_29791,N_29184);
xnor UO_846 (O_846,N_29144,N_29777);
xor UO_847 (O_847,N_29080,N_29616);
xnor UO_848 (O_848,N_29958,N_29407);
and UO_849 (O_849,N_29519,N_29583);
xor UO_850 (O_850,N_29441,N_29393);
nor UO_851 (O_851,N_29988,N_29859);
or UO_852 (O_852,N_29747,N_29580);
nor UO_853 (O_853,N_29586,N_29217);
nand UO_854 (O_854,N_29030,N_29551);
nand UO_855 (O_855,N_29030,N_29176);
and UO_856 (O_856,N_29218,N_29628);
nor UO_857 (O_857,N_29547,N_29971);
or UO_858 (O_858,N_29244,N_29898);
nand UO_859 (O_859,N_29402,N_29449);
and UO_860 (O_860,N_29445,N_29415);
or UO_861 (O_861,N_29508,N_29751);
and UO_862 (O_862,N_29055,N_29669);
xor UO_863 (O_863,N_29141,N_29816);
or UO_864 (O_864,N_29721,N_29216);
nand UO_865 (O_865,N_29514,N_29119);
or UO_866 (O_866,N_29061,N_29053);
nand UO_867 (O_867,N_29508,N_29575);
or UO_868 (O_868,N_29120,N_29582);
nand UO_869 (O_869,N_29976,N_29784);
xnor UO_870 (O_870,N_29758,N_29332);
nand UO_871 (O_871,N_29604,N_29475);
or UO_872 (O_872,N_29464,N_29190);
and UO_873 (O_873,N_29970,N_29477);
nand UO_874 (O_874,N_29183,N_29550);
or UO_875 (O_875,N_29133,N_29758);
nand UO_876 (O_876,N_29054,N_29146);
nor UO_877 (O_877,N_29076,N_29564);
nor UO_878 (O_878,N_29232,N_29338);
and UO_879 (O_879,N_29360,N_29662);
nand UO_880 (O_880,N_29085,N_29936);
xor UO_881 (O_881,N_29467,N_29146);
nand UO_882 (O_882,N_29467,N_29912);
xor UO_883 (O_883,N_29123,N_29057);
xor UO_884 (O_884,N_29440,N_29988);
xnor UO_885 (O_885,N_29199,N_29246);
and UO_886 (O_886,N_29865,N_29716);
nand UO_887 (O_887,N_29742,N_29158);
and UO_888 (O_888,N_29446,N_29721);
or UO_889 (O_889,N_29724,N_29298);
nor UO_890 (O_890,N_29637,N_29795);
or UO_891 (O_891,N_29989,N_29816);
or UO_892 (O_892,N_29688,N_29162);
nand UO_893 (O_893,N_29745,N_29881);
nand UO_894 (O_894,N_29604,N_29343);
xor UO_895 (O_895,N_29734,N_29306);
nor UO_896 (O_896,N_29564,N_29520);
nand UO_897 (O_897,N_29127,N_29655);
and UO_898 (O_898,N_29234,N_29518);
nand UO_899 (O_899,N_29975,N_29110);
xnor UO_900 (O_900,N_29619,N_29174);
and UO_901 (O_901,N_29135,N_29171);
or UO_902 (O_902,N_29636,N_29337);
or UO_903 (O_903,N_29674,N_29489);
and UO_904 (O_904,N_29117,N_29804);
or UO_905 (O_905,N_29541,N_29245);
nand UO_906 (O_906,N_29390,N_29357);
nor UO_907 (O_907,N_29387,N_29504);
xnor UO_908 (O_908,N_29331,N_29638);
nor UO_909 (O_909,N_29257,N_29233);
nand UO_910 (O_910,N_29144,N_29082);
and UO_911 (O_911,N_29526,N_29985);
nor UO_912 (O_912,N_29876,N_29584);
xor UO_913 (O_913,N_29080,N_29460);
xor UO_914 (O_914,N_29630,N_29631);
nor UO_915 (O_915,N_29943,N_29727);
and UO_916 (O_916,N_29974,N_29390);
xor UO_917 (O_917,N_29994,N_29572);
xor UO_918 (O_918,N_29397,N_29979);
or UO_919 (O_919,N_29091,N_29667);
nor UO_920 (O_920,N_29027,N_29142);
and UO_921 (O_921,N_29713,N_29070);
and UO_922 (O_922,N_29238,N_29451);
and UO_923 (O_923,N_29868,N_29776);
and UO_924 (O_924,N_29144,N_29832);
or UO_925 (O_925,N_29197,N_29495);
and UO_926 (O_926,N_29531,N_29008);
nor UO_927 (O_927,N_29324,N_29531);
nor UO_928 (O_928,N_29963,N_29524);
nand UO_929 (O_929,N_29722,N_29111);
nor UO_930 (O_930,N_29675,N_29483);
nand UO_931 (O_931,N_29836,N_29056);
nand UO_932 (O_932,N_29544,N_29038);
xor UO_933 (O_933,N_29905,N_29862);
or UO_934 (O_934,N_29271,N_29166);
or UO_935 (O_935,N_29195,N_29154);
xnor UO_936 (O_936,N_29035,N_29981);
and UO_937 (O_937,N_29161,N_29811);
and UO_938 (O_938,N_29320,N_29522);
nand UO_939 (O_939,N_29699,N_29390);
nor UO_940 (O_940,N_29332,N_29216);
or UO_941 (O_941,N_29938,N_29805);
or UO_942 (O_942,N_29913,N_29886);
and UO_943 (O_943,N_29013,N_29515);
xnor UO_944 (O_944,N_29280,N_29589);
or UO_945 (O_945,N_29780,N_29346);
nor UO_946 (O_946,N_29766,N_29040);
and UO_947 (O_947,N_29887,N_29359);
xor UO_948 (O_948,N_29969,N_29230);
nand UO_949 (O_949,N_29211,N_29912);
xnor UO_950 (O_950,N_29711,N_29330);
or UO_951 (O_951,N_29036,N_29156);
or UO_952 (O_952,N_29970,N_29552);
or UO_953 (O_953,N_29785,N_29661);
nand UO_954 (O_954,N_29976,N_29403);
xor UO_955 (O_955,N_29822,N_29989);
xor UO_956 (O_956,N_29837,N_29285);
or UO_957 (O_957,N_29400,N_29820);
and UO_958 (O_958,N_29554,N_29299);
nor UO_959 (O_959,N_29544,N_29708);
xor UO_960 (O_960,N_29624,N_29009);
or UO_961 (O_961,N_29726,N_29020);
and UO_962 (O_962,N_29908,N_29696);
nand UO_963 (O_963,N_29895,N_29260);
xnor UO_964 (O_964,N_29304,N_29945);
and UO_965 (O_965,N_29790,N_29099);
nand UO_966 (O_966,N_29219,N_29374);
or UO_967 (O_967,N_29939,N_29381);
nand UO_968 (O_968,N_29486,N_29826);
and UO_969 (O_969,N_29767,N_29215);
and UO_970 (O_970,N_29328,N_29529);
and UO_971 (O_971,N_29863,N_29917);
nor UO_972 (O_972,N_29979,N_29176);
and UO_973 (O_973,N_29878,N_29211);
xor UO_974 (O_974,N_29210,N_29133);
and UO_975 (O_975,N_29895,N_29764);
nand UO_976 (O_976,N_29541,N_29743);
xnor UO_977 (O_977,N_29259,N_29591);
xnor UO_978 (O_978,N_29171,N_29381);
nand UO_979 (O_979,N_29105,N_29068);
xnor UO_980 (O_980,N_29645,N_29601);
xnor UO_981 (O_981,N_29958,N_29847);
and UO_982 (O_982,N_29224,N_29704);
and UO_983 (O_983,N_29752,N_29570);
and UO_984 (O_984,N_29318,N_29233);
nand UO_985 (O_985,N_29526,N_29909);
xnor UO_986 (O_986,N_29384,N_29923);
nand UO_987 (O_987,N_29979,N_29672);
xnor UO_988 (O_988,N_29903,N_29287);
or UO_989 (O_989,N_29662,N_29772);
or UO_990 (O_990,N_29298,N_29066);
nor UO_991 (O_991,N_29729,N_29161);
xor UO_992 (O_992,N_29118,N_29085);
or UO_993 (O_993,N_29795,N_29211);
or UO_994 (O_994,N_29761,N_29001);
or UO_995 (O_995,N_29479,N_29017);
xnor UO_996 (O_996,N_29739,N_29707);
xor UO_997 (O_997,N_29883,N_29760);
nor UO_998 (O_998,N_29743,N_29901);
and UO_999 (O_999,N_29093,N_29742);
nand UO_1000 (O_1000,N_29262,N_29731);
or UO_1001 (O_1001,N_29472,N_29235);
nor UO_1002 (O_1002,N_29935,N_29871);
or UO_1003 (O_1003,N_29785,N_29497);
nand UO_1004 (O_1004,N_29358,N_29383);
nand UO_1005 (O_1005,N_29106,N_29114);
nand UO_1006 (O_1006,N_29207,N_29757);
nor UO_1007 (O_1007,N_29538,N_29510);
xor UO_1008 (O_1008,N_29784,N_29277);
nand UO_1009 (O_1009,N_29306,N_29640);
xor UO_1010 (O_1010,N_29277,N_29825);
and UO_1011 (O_1011,N_29660,N_29382);
nand UO_1012 (O_1012,N_29468,N_29656);
or UO_1013 (O_1013,N_29589,N_29531);
xnor UO_1014 (O_1014,N_29100,N_29053);
or UO_1015 (O_1015,N_29804,N_29406);
nand UO_1016 (O_1016,N_29620,N_29707);
xor UO_1017 (O_1017,N_29088,N_29563);
and UO_1018 (O_1018,N_29894,N_29063);
or UO_1019 (O_1019,N_29715,N_29317);
xor UO_1020 (O_1020,N_29740,N_29583);
nor UO_1021 (O_1021,N_29094,N_29679);
xnor UO_1022 (O_1022,N_29350,N_29314);
xor UO_1023 (O_1023,N_29594,N_29019);
nand UO_1024 (O_1024,N_29052,N_29646);
and UO_1025 (O_1025,N_29679,N_29742);
nor UO_1026 (O_1026,N_29348,N_29071);
or UO_1027 (O_1027,N_29049,N_29798);
nand UO_1028 (O_1028,N_29903,N_29946);
and UO_1029 (O_1029,N_29687,N_29512);
xnor UO_1030 (O_1030,N_29259,N_29992);
or UO_1031 (O_1031,N_29975,N_29867);
xor UO_1032 (O_1032,N_29584,N_29608);
xor UO_1033 (O_1033,N_29214,N_29158);
xnor UO_1034 (O_1034,N_29507,N_29975);
nand UO_1035 (O_1035,N_29968,N_29090);
and UO_1036 (O_1036,N_29017,N_29987);
nor UO_1037 (O_1037,N_29454,N_29003);
and UO_1038 (O_1038,N_29280,N_29163);
nor UO_1039 (O_1039,N_29672,N_29426);
or UO_1040 (O_1040,N_29136,N_29407);
nor UO_1041 (O_1041,N_29463,N_29871);
and UO_1042 (O_1042,N_29691,N_29950);
nand UO_1043 (O_1043,N_29317,N_29844);
or UO_1044 (O_1044,N_29606,N_29610);
nor UO_1045 (O_1045,N_29795,N_29337);
nand UO_1046 (O_1046,N_29405,N_29775);
xnor UO_1047 (O_1047,N_29694,N_29763);
or UO_1048 (O_1048,N_29580,N_29498);
nand UO_1049 (O_1049,N_29579,N_29403);
or UO_1050 (O_1050,N_29261,N_29112);
xnor UO_1051 (O_1051,N_29740,N_29102);
nor UO_1052 (O_1052,N_29339,N_29509);
nand UO_1053 (O_1053,N_29299,N_29761);
or UO_1054 (O_1054,N_29563,N_29556);
xor UO_1055 (O_1055,N_29617,N_29826);
xor UO_1056 (O_1056,N_29244,N_29396);
and UO_1057 (O_1057,N_29847,N_29653);
xor UO_1058 (O_1058,N_29827,N_29904);
nand UO_1059 (O_1059,N_29223,N_29347);
and UO_1060 (O_1060,N_29457,N_29029);
and UO_1061 (O_1061,N_29432,N_29087);
nor UO_1062 (O_1062,N_29147,N_29882);
or UO_1063 (O_1063,N_29020,N_29682);
and UO_1064 (O_1064,N_29236,N_29810);
nor UO_1065 (O_1065,N_29832,N_29961);
nor UO_1066 (O_1066,N_29494,N_29827);
nand UO_1067 (O_1067,N_29677,N_29834);
and UO_1068 (O_1068,N_29816,N_29127);
or UO_1069 (O_1069,N_29798,N_29376);
nor UO_1070 (O_1070,N_29696,N_29198);
nor UO_1071 (O_1071,N_29188,N_29428);
and UO_1072 (O_1072,N_29335,N_29024);
xnor UO_1073 (O_1073,N_29339,N_29437);
or UO_1074 (O_1074,N_29260,N_29040);
nor UO_1075 (O_1075,N_29006,N_29012);
and UO_1076 (O_1076,N_29939,N_29016);
nand UO_1077 (O_1077,N_29975,N_29238);
nor UO_1078 (O_1078,N_29887,N_29489);
nand UO_1079 (O_1079,N_29180,N_29171);
xnor UO_1080 (O_1080,N_29990,N_29816);
and UO_1081 (O_1081,N_29200,N_29364);
nand UO_1082 (O_1082,N_29790,N_29548);
nor UO_1083 (O_1083,N_29092,N_29083);
xor UO_1084 (O_1084,N_29827,N_29927);
and UO_1085 (O_1085,N_29043,N_29531);
nor UO_1086 (O_1086,N_29571,N_29418);
nand UO_1087 (O_1087,N_29837,N_29814);
nor UO_1088 (O_1088,N_29484,N_29138);
or UO_1089 (O_1089,N_29487,N_29957);
nand UO_1090 (O_1090,N_29307,N_29115);
or UO_1091 (O_1091,N_29208,N_29229);
nor UO_1092 (O_1092,N_29012,N_29418);
or UO_1093 (O_1093,N_29728,N_29763);
nor UO_1094 (O_1094,N_29990,N_29720);
nor UO_1095 (O_1095,N_29408,N_29880);
xnor UO_1096 (O_1096,N_29792,N_29557);
and UO_1097 (O_1097,N_29464,N_29216);
nand UO_1098 (O_1098,N_29362,N_29410);
nor UO_1099 (O_1099,N_29630,N_29949);
xnor UO_1100 (O_1100,N_29553,N_29017);
nand UO_1101 (O_1101,N_29995,N_29949);
nor UO_1102 (O_1102,N_29755,N_29211);
xnor UO_1103 (O_1103,N_29242,N_29514);
xor UO_1104 (O_1104,N_29245,N_29410);
nand UO_1105 (O_1105,N_29117,N_29970);
nor UO_1106 (O_1106,N_29311,N_29005);
or UO_1107 (O_1107,N_29721,N_29255);
or UO_1108 (O_1108,N_29129,N_29922);
and UO_1109 (O_1109,N_29428,N_29976);
nor UO_1110 (O_1110,N_29773,N_29699);
nor UO_1111 (O_1111,N_29427,N_29503);
nand UO_1112 (O_1112,N_29746,N_29771);
or UO_1113 (O_1113,N_29263,N_29270);
xnor UO_1114 (O_1114,N_29017,N_29160);
xnor UO_1115 (O_1115,N_29846,N_29635);
or UO_1116 (O_1116,N_29939,N_29299);
or UO_1117 (O_1117,N_29371,N_29629);
or UO_1118 (O_1118,N_29637,N_29797);
nand UO_1119 (O_1119,N_29940,N_29414);
or UO_1120 (O_1120,N_29662,N_29527);
xnor UO_1121 (O_1121,N_29985,N_29887);
xor UO_1122 (O_1122,N_29173,N_29662);
or UO_1123 (O_1123,N_29965,N_29263);
and UO_1124 (O_1124,N_29418,N_29666);
xor UO_1125 (O_1125,N_29213,N_29485);
nand UO_1126 (O_1126,N_29704,N_29698);
nor UO_1127 (O_1127,N_29134,N_29041);
xnor UO_1128 (O_1128,N_29411,N_29293);
and UO_1129 (O_1129,N_29562,N_29138);
nor UO_1130 (O_1130,N_29778,N_29462);
or UO_1131 (O_1131,N_29797,N_29174);
and UO_1132 (O_1132,N_29492,N_29660);
xnor UO_1133 (O_1133,N_29940,N_29318);
or UO_1134 (O_1134,N_29021,N_29789);
nand UO_1135 (O_1135,N_29884,N_29860);
or UO_1136 (O_1136,N_29168,N_29159);
nand UO_1137 (O_1137,N_29660,N_29103);
and UO_1138 (O_1138,N_29070,N_29519);
nand UO_1139 (O_1139,N_29963,N_29619);
or UO_1140 (O_1140,N_29058,N_29184);
xor UO_1141 (O_1141,N_29769,N_29619);
nand UO_1142 (O_1142,N_29664,N_29435);
nor UO_1143 (O_1143,N_29442,N_29581);
nor UO_1144 (O_1144,N_29590,N_29711);
nor UO_1145 (O_1145,N_29892,N_29821);
and UO_1146 (O_1146,N_29839,N_29427);
or UO_1147 (O_1147,N_29002,N_29347);
and UO_1148 (O_1148,N_29057,N_29295);
nand UO_1149 (O_1149,N_29416,N_29748);
or UO_1150 (O_1150,N_29755,N_29667);
or UO_1151 (O_1151,N_29720,N_29767);
xor UO_1152 (O_1152,N_29537,N_29777);
nor UO_1153 (O_1153,N_29032,N_29713);
and UO_1154 (O_1154,N_29020,N_29633);
nor UO_1155 (O_1155,N_29437,N_29794);
nor UO_1156 (O_1156,N_29209,N_29503);
nor UO_1157 (O_1157,N_29850,N_29715);
or UO_1158 (O_1158,N_29617,N_29938);
and UO_1159 (O_1159,N_29766,N_29024);
xnor UO_1160 (O_1160,N_29325,N_29720);
nor UO_1161 (O_1161,N_29457,N_29929);
nor UO_1162 (O_1162,N_29861,N_29922);
and UO_1163 (O_1163,N_29124,N_29596);
and UO_1164 (O_1164,N_29539,N_29614);
or UO_1165 (O_1165,N_29131,N_29892);
or UO_1166 (O_1166,N_29004,N_29259);
nor UO_1167 (O_1167,N_29129,N_29245);
nor UO_1168 (O_1168,N_29528,N_29405);
xor UO_1169 (O_1169,N_29449,N_29684);
xnor UO_1170 (O_1170,N_29817,N_29653);
nor UO_1171 (O_1171,N_29555,N_29581);
nand UO_1172 (O_1172,N_29231,N_29230);
or UO_1173 (O_1173,N_29350,N_29098);
nor UO_1174 (O_1174,N_29648,N_29594);
or UO_1175 (O_1175,N_29131,N_29007);
nand UO_1176 (O_1176,N_29911,N_29262);
nor UO_1177 (O_1177,N_29632,N_29654);
xor UO_1178 (O_1178,N_29784,N_29179);
or UO_1179 (O_1179,N_29324,N_29834);
xor UO_1180 (O_1180,N_29432,N_29010);
and UO_1181 (O_1181,N_29896,N_29380);
and UO_1182 (O_1182,N_29289,N_29354);
or UO_1183 (O_1183,N_29682,N_29717);
nor UO_1184 (O_1184,N_29976,N_29451);
nor UO_1185 (O_1185,N_29251,N_29227);
or UO_1186 (O_1186,N_29212,N_29441);
or UO_1187 (O_1187,N_29432,N_29505);
or UO_1188 (O_1188,N_29849,N_29704);
nor UO_1189 (O_1189,N_29941,N_29444);
and UO_1190 (O_1190,N_29593,N_29723);
nand UO_1191 (O_1191,N_29816,N_29850);
nand UO_1192 (O_1192,N_29256,N_29043);
nand UO_1193 (O_1193,N_29624,N_29262);
nor UO_1194 (O_1194,N_29157,N_29482);
nand UO_1195 (O_1195,N_29065,N_29234);
nand UO_1196 (O_1196,N_29817,N_29028);
nor UO_1197 (O_1197,N_29383,N_29721);
xor UO_1198 (O_1198,N_29861,N_29300);
nand UO_1199 (O_1199,N_29027,N_29954);
xor UO_1200 (O_1200,N_29968,N_29172);
or UO_1201 (O_1201,N_29891,N_29475);
nor UO_1202 (O_1202,N_29882,N_29383);
nand UO_1203 (O_1203,N_29098,N_29907);
xnor UO_1204 (O_1204,N_29291,N_29038);
and UO_1205 (O_1205,N_29154,N_29978);
xor UO_1206 (O_1206,N_29571,N_29863);
xor UO_1207 (O_1207,N_29869,N_29165);
or UO_1208 (O_1208,N_29846,N_29396);
and UO_1209 (O_1209,N_29740,N_29711);
nand UO_1210 (O_1210,N_29809,N_29821);
nor UO_1211 (O_1211,N_29474,N_29484);
nor UO_1212 (O_1212,N_29715,N_29966);
nor UO_1213 (O_1213,N_29863,N_29757);
nor UO_1214 (O_1214,N_29903,N_29258);
xor UO_1215 (O_1215,N_29294,N_29520);
or UO_1216 (O_1216,N_29037,N_29904);
and UO_1217 (O_1217,N_29174,N_29899);
and UO_1218 (O_1218,N_29373,N_29308);
nand UO_1219 (O_1219,N_29957,N_29474);
nand UO_1220 (O_1220,N_29483,N_29621);
nor UO_1221 (O_1221,N_29802,N_29481);
nor UO_1222 (O_1222,N_29957,N_29657);
and UO_1223 (O_1223,N_29040,N_29848);
and UO_1224 (O_1224,N_29462,N_29723);
nor UO_1225 (O_1225,N_29952,N_29222);
or UO_1226 (O_1226,N_29973,N_29465);
xnor UO_1227 (O_1227,N_29007,N_29059);
and UO_1228 (O_1228,N_29119,N_29537);
nor UO_1229 (O_1229,N_29283,N_29545);
nor UO_1230 (O_1230,N_29758,N_29127);
or UO_1231 (O_1231,N_29272,N_29830);
nand UO_1232 (O_1232,N_29921,N_29256);
nor UO_1233 (O_1233,N_29617,N_29802);
or UO_1234 (O_1234,N_29076,N_29782);
and UO_1235 (O_1235,N_29701,N_29856);
nor UO_1236 (O_1236,N_29876,N_29525);
and UO_1237 (O_1237,N_29899,N_29852);
xor UO_1238 (O_1238,N_29595,N_29400);
nand UO_1239 (O_1239,N_29459,N_29431);
nand UO_1240 (O_1240,N_29142,N_29856);
nand UO_1241 (O_1241,N_29498,N_29502);
nor UO_1242 (O_1242,N_29101,N_29124);
nand UO_1243 (O_1243,N_29402,N_29321);
nand UO_1244 (O_1244,N_29428,N_29552);
and UO_1245 (O_1245,N_29397,N_29824);
nand UO_1246 (O_1246,N_29745,N_29072);
or UO_1247 (O_1247,N_29218,N_29894);
and UO_1248 (O_1248,N_29549,N_29325);
nand UO_1249 (O_1249,N_29762,N_29735);
xor UO_1250 (O_1250,N_29985,N_29903);
nand UO_1251 (O_1251,N_29500,N_29746);
xnor UO_1252 (O_1252,N_29215,N_29508);
nand UO_1253 (O_1253,N_29352,N_29109);
nor UO_1254 (O_1254,N_29162,N_29820);
nand UO_1255 (O_1255,N_29661,N_29319);
nor UO_1256 (O_1256,N_29854,N_29375);
and UO_1257 (O_1257,N_29323,N_29813);
xor UO_1258 (O_1258,N_29344,N_29703);
xnor UO_1259 (O_1259,N_29042,N_29865);
or UO_1260 (O_1260,N_29223,N_29020);
xnor UO_1261 (O_1261,N_29506,N_29487);
or UO_1262 (O_1262,N_29482,N_29746);
nor UO_1263 (O_1263,N_29070,N_29226);
nand UO_1264 (O_1264,N_29396,N_29996);
nand UO_1265 (O_1265,N_29980,N_29571);
xnor UO_1266 (O_1266,N_29745,N_29183);
nand UO_1267 (O_1267,N_29951,N_29284);
nor UO_1268 (O_1268,N_29708,N_29118);
nor UO_1269 (O_1269,N_29635,N_29949);
nor UO_1270 (O_1270,N_29995,N_29393);
xor UO_1271 (O_1271,N_29124,N_29532);
nand UO_1272 (O_1272,N_29690,N_29992);
and UO_1273 (O_1273,N_29374,N_29740);
and UO_1274 (O_1274,N_29484,N_29504);
xnor UO_1275 (O_1275,N_29067,N_29987);
nor UO_1276 (O_1276,N_29469,N_29902);
nand UO_1277 (O_1277,N_29039,N_29878);
nor UO_1278 (O_1278,N_29281,N_29542);
or UO_1279 (O_1279,N_29802,N_29819);
and UO_1280 (O_1280,N_29563,N_29943);
and UO_1281 (O_1281,N_29576,N_29568);
nand UO_1282 (O_1282,N_29132,N_29344);
nor UO_1283 (O_1283,N_29275,N_29530);
nor UO_1284 (O_1284,N_29719,N_29379);
xnor UO_1285 (O_1285,N_29973,N_29447);
nand UO_1286 (O_1286,N_29612,N_29899);
nand UO_1287 (O_1287,N_29773,N_29253);
or UO_1288 (O_1288,N_29977,N_29618);
nor UO_1289 (O_1289,N_29034,N_29797);
or UO_1290 (O_1290,N_29268,N_29368);
and UO_1291 (O_1291,N_29741,N_29218);
nor UO_1292 (O_1292,N_29613,N_29141);
and UO_1293 (O_1293,N_29329,N_29013);
nor UO_1294 (O_1294,N_29740,N_29142);
and UO_1295 (O_1295,N_29565,N_29616);
or UO_1296 (O_1296,N_29851,N_29704);
or UO_1297 (O_1297,N_29061,N_29873);
and UO_1298 (O_1298,N_29979,N_29529);
nand UO_1299 (O_1299,N_29000,N_29990);
and UO_1300 (O_1300,N_29611,N_29582);
nand UO_1301 (O_1301,N_29319,N_29495);
nand UO_1302 (O_1302,N_29266,N_29803);
or UO_1303 (O_1303,N_29937,N_29678);
nand UO_1304 (O_1304,N_29003,N_29527);
or UO_1305 (O_1305,N_29834,N_29184);
xor UO_1306 (O_1306,N_29600,N_29149);
nand UO_1307 (O_1307,N_29665,N_29291);
nand UO_1308 (O_1308,N_29129,N_29040);
or UO_1309 (O_1309,N_29506,N_29421);
nor UO_1310 (O_1310,N_29704,N_29373);
or UO_1311 (O_1311,N_29777,N_29762);
xnor UO_1312 (O_1312,N_29075,N_29004);
and UO_1313 (O_1313,N_29763,N_29372);
nor UO_1314 (O_1314,N_29141,N_29687);
or UO_1315 (O_1315,N_29798,N_29150);
xor UO_1316 (O_1316,N_29010,N_29375);
nor UO_1317 (O_1317,N_29576,N_29777);
nand UO_1318 (O_1318,N_29574,N_29980);
nand UO_1319 (O_1319,N_29873,N_29305);
nor UO_1320 (O_1320,N_29804,N_29279);
or UO_1321 (O_1321,N_29409,N_29093);
xnor UO_1322 (O_1322,N_29976,N_29083);
xnor UO_1323 (O_1323,N_29325,N_29267);
nor UO_1324 (O_1324,N_29032,N_29276);
and UO_1325 (O_1325,N_29275,N_29389);
or UO_1326 (O_1326,N_29180,N_29796);
nor UO_1327 (O_1327,N_29682,N_29502);
and UO_1328 (O_1328,N_29019,N_29148);
and UO_1329 (O_1329,N_29328,N_29102);
xor UO_1330 (O_1330,N_29834,N_29618);
or UO_1331 (O_1331,N_29334,N_29882);
and UO_1332 (O_1332,N_29897,N_29781);
xor UO_1333 (O_1333,N_29748,N_29739);
or UO_1334 (O_1334,N_29560,N_29515);
and UO_1335 (O_1335,N_29812,N_29471);
nand UO_1336 (O_1336,N_29382,N_29169);
nor UO_1337 (O_1337,N_29653,N_29788);
or UO_1338 (O_1338,N_29664,N_29641);
or UO_1339 (O_1339,N_29301,N_29519);
xor UO_1340 (O_1340,N_29790,N_29689);
nor UO_1341 (O_1341,N_29400,N_29626);
nand UO_1342 (O_1342,N_29675,N_29373);
nor UO_1343 (O_1343,N_29991,N_29391);
and UO_1344 (O_1344,N_29617,N_29314);
nand UO_1345 (O_1345,N_29700,N_29202);
nor UO_1346 (O_1346,N_29862,N_29556);
xor UO_1347 (O_1347,N_29720,N_29277);
or UO_1348 (O_1348,N_29285,N_29885);
and UO_1349 (O_1349,N_29983,N_29512);
xnor UO_1350 (O_1350,N_29386,N_29571);
xnor UO_1351 (O_1351,N_29174,N_29877);
and UO_1352 (O_1352,N_29916,N_29820);
and UO_1353 (O_1353,N_29488,N_29820);
and UO_1354 (O_1354,N_29945,N_29168);
or UO_1355 (O_1355,N_29039,N_29466);
or UO_1356 (O_1356,N_29425,N_29188);
nor UO_1357 (O_1357,N_29146,N_29782);
xor UO_1358 (O_1358,N_29929,N_29883);
or UO_1359 (O_1359,N_29166,N_29035);
and UO_1360 (O_1360,N_29301,N_29118);
and UO_1361 (O_1361,N_29766,N_29987);
nor UO_1362 (O_1362,N_29419,N_29203);
xor UO_1363 (O_1363,N_29417,N_29146);
or UO_1364 (O_1364,N_29405,N_29869);
nand UO_1365 (O_1365,N_29406,N_29956);
and UO_1366 (O_1366,N_29432,N_29878);
xnor UO_1367 (O_1367,N_29607,N_29063);
or UO_1368 (O_1368,N_29588,N_29881);
nand UO_1369 (O_1369,N_29969,N_29533);
or UO_1370 (O_1370,N_29468,N_29230);
nand UO_1371 (O_1371,N_29385,N_29074);
nor UO_1372 (O_1372,N_29194,N_29207);
xnor UO_1373 (O_1373,N_29686,N_29855);
and UO_1374 (O_1374,N_29434,N_29399);
xnor UO_1375 (O_1375,N_29713,N_29176);
xor UO_1376 (O_1376,N_29768,N_29437);
and UO_1377 (O_1377,N_29131,N_29763);
nand UO_1378 (O_1378,N_29564,N_29543);
or UO_1379 (O_1379,N_29612,N_29521);
and UO_1380 (O_1380,N_29913,N_29675);
xor UO_1381 (O_1381,N_29956,N_29033);
nor UO_1382 (O_1382,N_29571,N_29787);
nor UO_1383 (O_1383,N_29505,N_29256);
and UO_1384 (O_1384,N_29421,N_29064);
nand UO_1385 (O_1385,N_29877,N_29329);
and UO_1386 (O_1386,N_29795,N_29097);
xor UO_1387 (O_1387,N_29660,N_29217);
xnor UO_1388 (O_1388,N_29664,N_29155);
and UO_1389 (O_1389,N_29191,N_29510);
xor UO_1390 (O_1390,N_29329,N_29819);
xnor UO_1391 (O_1391,N_29406,N_29267);
xnor UO_1392 (O_1392,N_29824,N_29640);
nand UO_1393 (O_1393,N_29445,N_29657);
nand UO_1394 (O_1394,N_29240,N_29062);
nand UO_1395 (O_1395,N_29451,N_29788);
and UO_1396 (O_1396,N_29120,N_29191);
xor UO_1397 (O_1397,N_29840,N_29844);
nor UO_1398 (O_1398,N_29243,N_29467);
nor UO_1399 (O_1399,N_29336,N_29846);
and UO_1400 (O_1400,N_29142,N_29165);
nor UO_1401 (O_1401,N_29593,N_29201);
xor UO_1402 (O_1402,N_29437,N_29042);
and UO_1403 (O_1403,N_29604,N_29027);
and UO_1404 (O_1404,N_29394,N_29220);
and UO_1405 (O_1405,N_29951,N_29969);
or UO_1406 (O_1406,N_29399,N_29178);
or UO_1407 (O_1407,N_29789,N_29850);
or UO_1408 (O_1408,N_29069,N_29360);
or UO_1409 (O_1409,N_29183,N_29836);
nor UO_1410 (O_1410,N_29254,N_29939);
nor UO_1411 (O_1411,N_29269,N_29020);
xnor UO_1412 (O_1412,N_29208,N_29016);
nand UO_1413 (O_1413,N_29831,N_29888);
nand UO_1414 (O_1414,N_29644,N_29678);
nor UO_1415 (O_1415,N_29293,N_29804);
xor UO_1416 (O_1416,N_29748,N_29004);
and UO_1417 (O_1417,N_29693,N_29840);
nor UO_1418 (O_1418,N_29879,N_29693);
nand UO_1419 (O_1419,N_29941,N_29415);
nor UO_1420 (O_1420,N_29520,N_29674);
and UO_1421 (O_1421,N_29151,N_29537);
nand UO_1422 (O_1422,N_29901,N_29865);
nand UO_1423 (O_1423,N_29172,N_29816);
nor UO_1424 (O_1424,N_29905,N_29793);
and UO_1425 (O_1425,N_29561,N_29924);
nor UO_1426 (O_1426,N_29005,N_29026);
nor UO_1427 (O_1427,N_29195,N_29591);
nand UO_1428 (O_1428,N_29443,N_29830);
xnor UO_1429 (O_1429,N_29048,N_29515);
and UO_1430 (O_1430,N_29707,N_29670);
nor UO_1431 (O_1431,N_29672,N_29262);
and UO_1432 (O_1432,N_29725,N_29102);
xnor UO_1433 (O_1433,N_29153,N_29580);
and UO_1434 (O_1434,N_29929,N_29396);
and UO_1435 (O_1435,N_29011,N_29634);
or UO_1436 (O_1436,N_29117,N_29782);
nand UO_1437 (O_1437,N_29185,N_29585);
nand UO_1438 (O_1438,N_29060,N_29283);
nand UO_1439 (O_1439,N_29066,N_29750);
nor UO_1440 (O_1440,N_29842,N_29738);
xor UO_1441 (O_1441,N_29527,N_29972);
xnor UO_1442 (O_1442,N_29720,N_29828);
and UO_1443 (O_1443,N_29270,N_29039);
xnor UO_1444 (O_1444,N_29460,N_29661);
nor UO_1445 (O_1445,N_29360,N_29843);
nand UO_1446 (O_1446,N_29793,N_29711);
xor UO_1447 (O_1447,N_29678,N_29785);
or UO_1448 (O_1448,N_29453,N_29574);
nor UO_1449 (O_1449,N_29214,N_29233);
and UO_1450 (O_1450,N_29062,N_29276);
nand UO_1451 (O_1451,N_29859,N_29313);
or UO_1452 (O_1452,N_29206,N_29885);
nand UO_1453 (O_1453,N_29075,N_29108);
nor UO_1454 (O_1454,N_29700,N_29438);
or UO_1455 (O_1455,N_29013,N_29890);
nor UO_1456 (O_1456,N_29386,N_29887);
nand UO_1457 (O_1457,N_29539,N_29097);
nand UO_1458 (O_1458,N_29624,N_29510);
nor UO_1459 (O_1459,N_29392,N_29232);
nor UO_1460 (O_1460,N_29834,N_29826);
or UO_1461 (O_1461,N_29437,N_29636);
and UO_1462 (O_1462,N_29096,N_29267);
nand UO_1463 (O_1463,N_29610,N_29561);
nand UO_1464 (O_1464,N_29796,N_29991);
nor UO_1465 (O_1465,N_29737,N_29893);
nand UO_1466 (O_1466,N_29635,N_29502);
nand UO_1467 (O_1467,N_29929,N_29367);
and UO_1468 (O_1468,N_29198,N_29206);
or UO_1469 (O_1469,N_29184,N_29248);
and UO_1470 (O_1470,N_29253,N_29732);
or UO_1471 (O_1471,N_29398,N_29422);
or UO_1472 (O_1472,N_29916,N_29515);
nand UO_1473 (O_1473,N_29752,N_29996);
and UO_1474 (O_1474,N_29059,N_29064);
or UO_1475 (O_1475,N_29588,N_29933);
xor UO_1476 (O_1476,N_29792,N_29365);
xor UO_1477 (O_1477,N_29470,N_29743);
or UO_1478 (O_1478,N_29673,N_29865);
xor UO_1479 (O_1479,N_29205,N_29409);
nand UO_1480 (O_1480,N_29004,N_29909);
or UO_1481 (O_1481,N_29910,N_29438);
and UO_1482 (O_1482,N_29307,N_29623);
nor UO_1483 (O_1483,N_29093,N_29109);
or UO_1484 (O_1484,N_29220,N_29296);
nand UO_1485 (O_1485,N_29354,N_29006);
nand UO_1486 (O_1486,N_29278,N_29534);
and UO_1487 (O_1487,N_29743,N_29333);
or UO_1488 (O_1488,N_29359,N_29661);
xor UO_1489 (O_1489,N_29406,N_29346);
nor UO_1490 (O_1490,N_29002,N_29980);
and UO_1491 (O_1491,N_29572,N_29307);
and UO_1492 (O_1492,N_29873,N_29726);
nand UO_1493 (O_1493,N_29646,N_29942);
and UO_1494 (O_1494,N_29980,N_29591);
xor UO_1495 (O_1495,N_29897,N_29728);
nor UO_1496 (O_1496,N_29544,N_29232);
and UO_1497 (O_1497,N_29816,N_29196);
or UO_1498 (O_1498,N_29652,N_29509);
or UO_1499 (O_1499,N_29196,N_29628);
xnor UO_1500 (O_1500,N_29297,N_29061);
and UO_1501 (O_1501,N_29730,N_29165);
xor UO_1502 (O_1502,N_29857,N_29625);
nand UO_1503 (O_1503,N_29505,N_29588);
nand UO_1504 (O_1504,N_29635,N_29867);
and UO_1505 (O_1505,N_29109,N_29178);
xnor UO_1506 (O_1506,N_29287,N_29669);
and UO_1507 (O_1507,N_29500,N_29575);
or UO_1508 (O_1508,N_29116,N_29984);
and UO_1509 (O_1509,N_29211,N_29003);
or UO_1510 (O_1510,N_29801,N_29622);
xnor UO_1511 (O_1511,N_29001,N_29208);
or UO_1512 (O_1512,N_29254,N_29136);
nand UO_1513 (O_1513,N_29986,N_29635);
xnor UO_1514 (O_1514,N_29031,N_29151);
and UO_1515 (O_1515,N_29326,N_29657);
nor UO_1516 (O_1516,N_29022,N_29366);
or UO_1517 (O_1517,N_29889,N_29272);
and UO_1518 (O_1518,N_29560,N_29476);
xnor UO_1519 (O_1519,N_29099,N_29393);
nor UO_1520 (O_1520,N_29007,N_29667);
and UO_1521 (O_1521,N_29376,N_29384);
xnor UO_1522 (O_1522,N_29036,N_29902);
xnor UO_1523 (O_1523,N_29785,N_29964);
xor UO_1524 (O_1524,N_29324,N_29304);
nand UO_1525 (O_1525,N_29155,N_29455);
nor UO_1526 (O_1526,N_29665,N_29075);
and UO_1527 (O_1527,N_29082,N_29970);
nor UO_1528 (O_1528,N_29996,N_29414);
nand UO_1529 (O_1529,N_29210,N_29557);
xor UO_1530 (O_1530,N_29647,N_29127);
xor UO_1531 (O_1531,N_29212,N_29369);
or UO_1532 (O_1532,N_29301,N_29472);
nand UO_1533 (O_1533,N_29188,N_29793);
and UO_1534 (O_1534,N_29229,N_29715);
nor UO_1535 (O_1535,N_29503,N_29211);
or UO_1536 (O_1536,N_29771,N_29861);
nor UO_1537 (O_1537,N_29989,N_29918);
nand UO_1538 (O_1538,N_29532,N_29310);
xor UO_1539 (O_1539,N_29237,N_29837);
and UO_1540 (O_1540,N_29109,N_29996);
or UO_1541 (O_1541,N_29575,N_29849);
and UO_1542 (O_1542,N_29524,N_29227);
and UO_1543 (O_1543,N_29286,N_29670);
nand UO_1544 (O_1544,N_29614,N_29822);
and UO_1545 (O_1545,N_29960,N_29060);
nor UO_1546 (O_1546,N_29551,N_29752);
and UO_1547 (O_1547,N_29583,N_29925);
nand UO_1548 (O_1548,N_29858,N_29074);
nand UO_1549 (O_1549,N_29109,N_29583);
nor UO_1550 (O_1550,N_29111,N_29474);
nand UO_1551 (O_1551,N_29656,N_29490);
nor UO_1552 (O_1552,N_29732,N_29303);
nor UO_1553 (O_1553,N_29760,N_29049);
or UO_1554 (O_1554,N_29423,N_29544);
nor UO_1555 (O_1555,N_29046,N_29998);
nand UO_1556 (O_1556,N_29706,N_29251);
and UO_1557 (O_1557,N_29972,N_29593);
xor UO_1558 (O_1558,N_29009,N_29994);
or UO_1559 (O_1559,N_29621,N_29770);
and UO_1560 (O_1560,N_29370,N_29098);
and UO_1561 (O_1561,N_29344,N_29288);
nand UO_1562 (O_1562,N_29216,N_29767);
xor UO_1563 (O_1563,N_29227,N_29591);
xnor UO_1564 (O_1564,N_29261,N_29167);
or UO_1565 (O_1565,N_29447,N_29738);
nor UO_1566 (O_1566,N_29654,N_29280);
nand UO_1567 (O_1567,N_29897,N_29284);
xor UO_1568 (O_1568,N_29030,N_29102);
or UO_1569 (O_1569,N_29012,N_29635);
and UO_1570 (O_1570,N_29275,N_29616);
and UO_1571 (O_1571,N_29861,N_29310);
and UO_1572 (O_1572,N_29263,N_29850);
nor UO_1573 (O_1573,N_29542,N_29893);
xor UO_1574 (O_1574,N_29887,N_29144);
or UO_1575 (O_1575,N_29908,N_29338);
xor UO_1576 (O_1576,N_29661,N_29126);
nand UO_1577 (O_1577,N_29389,N_29852);
xnor UO_1578 (O_1578,N_29305,N_29390);
xor UO_1579 (O_1579,N_29088,N_29339);
nand UO_1580 (O_1580,N_29770,N_29274);
nor UO_1581 (O_1581,N_29093,N_29813);
xnor UO_1582 (O_1582,N_29365,N_29498);
nor UO_1583 (O_1583,N_29620,N_29775);
and UO_1584 (O_1584,N_29399,N_29721);
nand UO_1585 (O_1585,N_29865,N_29749);
nand UO_1586 (O_1586,N_29159,N_29388);
xnor UO_1587 (O_1587,N_29819,N_29889);
nand UO_1588 (O_1588,N_29175,N_29447);
xnor UO_1589 (O_1589,N_29137,N_29062);
nor UO_1590 (O_1590,N_29042,N_29957);
and UO_1591 (O_1591,N_29570,N_29342);
and UO_1592 (O_1592,N_29788,N_29808);
nand UO_1593 (O_1593,N_29428,N_29426);
or UO_1594 (O_1594,N_29266,N_29502);
nor UO_1595 (O_1595,N_29946,N_29070);
nor UO_1596 (O_1596,N_29332,N_29878);
xnor UO_1597 (O_1597,N_29422,N_29544);
nand UO_1598 (O_1598,N_29119,N_29163);
or UO_1599 (O_1599,N_29215,N_29756);
nand UO_1600 (O_1600,N_29342,N_29895);
xor UO_1601 (O_1601,N_29117,N_29346);
and UO_1602 (O_1602,N_29317,N_29705);
or UO_1603 (O_1603,N_29480,N_29381);
nor UO_1604 (O_1604,N_29751,N_29734);
or UO_1605 (O_1605,N_29348,N_29991);
nor UO_1606 (O_1606,N_29775,N_29281);
and UO_1607 (O_1607,N_29370,N_29852);
nand UO_1608 (O_1608,N_29059,N_29113);
or UO_1609 (O_1609,N_29449,N_29966);
nand UO_1610 (O_1610,N_29251,N_29368);
and UO_1611 (O_1611,N_29565,N_29125);
or UO_1612 (O_1612,N_29301,N_29570);
and UO_1613 (O_1613,N_29037,N_29150);
nor UO_1614 (O_1614,N_29077,N_29792);
xor UO_1615 (O_1615,N_29932,N_29371);
and UO_1616 (O_1616,N_29374,N_29634);
and UO_1617 (O_1617,N_29517,N_29148);
nor UO_1618 (O_1618,N_29954,N_29524);
nand UO_1619 (O_1619,N_29982,N_29053);
nor UO_1620 (O_1620,N_29688,N_29963);
nand UO_1621 (O_1621,N_29558,N_29786);
and UO_1622 (O_1622,N_29696,N_29588);
or UO_1623 (O_1623,N_29899,N_29513);
or UO_1624 (O_1624,N_29406,N_29232);
xnor UO_1625 (O_1625,N_29488,N_29232);
and UO_1626 (O_1626,N_29149,N_29203);
nand UO_1627 (O_1627,N_29446,N_29955);
or UO_1628 (O_1628,N_29607,N_29899);
or UO_1629 (O_1629,N_29805,N_29047);
nor UO_1630 (O_1630,N_29748,N_29908);
nand UO_1631 (O_1631,N_29510,N_29539);
nor UO_1632 (O_1632,N_29470,N_29995);
or UO_1633 (O_1633,N_29911,N_29375);
or UO_1634 (O_1634,N_29586,N_29193);
nor UO_1635 (O_1635,N_29343,N_29645);
nor UO_1636 (O_1636,N_29530,N_29818);
nand UO_1637 (O_1637,N_29228,N_29723);
nand UO_1638 (O_1638,N_29957,N_29737);
or UO_1639 (O_1639,N_29762,N_29922);
and UO_1640 (O_1640,N_29086,N_29668);
nor UO_1641 (O_1641,N_29695,N_29544);
or UO_1642 (O_1642,N_29076,N_29976);
nor UO_1643 (O_1643,N_29889,N_29003);
nand UO_1644 (O_1644,N_29354,N_29070);
nor UO_1645 (O_1645,N_29692,N_29540);
nor UO_1646 (O_1646,N_29548,N_29420);
xor UO_1647 (O_1647,N_29806,N_29231);
xor UO_1648 (O_1648,N_29582,N_29804);
and UO_1649 (O_1649,N_29504,N_29407);
and UO_1650 (O_1650,N_29679,N_29018);
xnor UO_1651 (O_1651,N_29310,N_29672);
and UO_1652 (O_1652,N_29390,N_29135);
nor UO_1653 (O_1653,N_29392,N_29065);
xnor UO_1654 (O_1654,N_29591,N_29024);
nand UO_1655 (O_1655,N_29281,N_29777);
or UO_1656 (O_1656,N_29267,N_29251);
nor UO_1657 (O_1657,N_29821,N_29371);
nand UO_1658 (O_1658,N_29590,N_29449);
nor UO_1659 (O_1659,N_29358,N_29577);
nor UO_1660 (O_1660,N_29608,N_29727);
nor UO_1661 (O_1661,N_29736,N_29439);
nor UO_1662 (O_1662,N_29074,N_29042);
or UO_1663 (O_1663,N_29337,N_29459);
xnor UO_1664 (O_1664,N_29148,N_29880);
nor UO_1665 (O_1665,N_29963,N_29849);
nor UO_1666 (O_1666,N_29321,N_29639);
nor UO_1667 (O_1667,N_29354,N_29473);
and UO_1668 (O_1668,N_29823,N_29674);
xor UO_1669 (O_1669,N_29324,N_29535);
or UO_1670 (O_1670,N_29081,N_29028);
or UO_1671 (O_1671,N_29407,N_29299);
nor UO_1672 (O_1672,N_29109,N_29808);
nor UO_1673 (O_1673,N_29599,N_29653);
and UO_1674 (O_1674,N_29909,N_29348);
nand UO_1675 (O_1675,N_29055,N_29748);
nor UO_1676 (O_1676,N_29456,N_29956);
and UO_1677 (O_1677,N_29951,N_29164);
xnor UO_1678 (O_1678,N_29662,N_29793);
nand UO_1679 (O_1679,N_29309,N_29092);
nor UO_1680 (O_1680,N_29150,N_29623);
and UO_1681 (O_1681,N_29800,N_29567);
and UO_1682 (O_1682,N_29800,N_29935);
nand UO_1683 (O_1683,N_29592,N_29705);
and UO_1684 (O_1684,N_29355,N_29956);
xnor UO_1685 (O_1685,N_29608,N_29269);
and UO_1686 (O_1686,N_29340,N_29080);
xor UO_1687 (O_1687,N_29760,N_29774);
nand UO_1688 (O_1688,N_29422,N_29621);
xor UO_1689 (O_1689,N_29760,N_29256);
nand UO_1690 (O_1690,N_29524,N_29535);
xnor UO_1691 (O_1691,N_29239,N_29223);
nand UO_1692 (O_1692,N_29483,N_29744);
or UO_1693 (O_1693,N_29656,N_29357);
and UO_1694 (O_1694,N_29448,N_29912);
nor UO_1695 (O_1695,N_29810,N_29524);
xnor UO_1696 (O_1696,N_29553,N_29377);
or UO_1697 (O_1697,N_29988,N_29924);
or UO_1698 (O_1698,N_29745,N_29939);
nor UO_1699 (O_1699,N_29917,N_29102);
nand UO_1700 (O_1700,N_29756,N_29837);
or UO_1701 (O_1701,N_29015,N_29697);
or UO_1702 (O_1702,N_29044,N_29984);
and UO_1703 (O_1703,N_29540,N_29440);
xor UO_1704 (O_1704,N_29589,N_29466);
xor UO_1705 (O_1705,N_29742,N_29136);
nand UO_1706 (O_1706,N_29131,N_29989);
and UO_1707 (O_1707,N_29484,N_29126);
xor UO_1708 (O_1708,N_29892,N_29090);
xnor UO_1709 (O_1709,N_29301,N_29034);
or UO_1710 (O_1710,N_29210,N_29781);
or UO_1711 (O_1711,N_29553,N_29879);
xor UO_1712 (O_1712,N_29727,N_29484);
nor UO_1713 (O_1713,N_29524,N_29785);
nand UO_1714 (O_1714,N_29046,N_29532);
and UO_1715 (O_1715,N_29598,N_29709);
nand UO_1716 (O_1716,N_29102,N_29020);
or UO_1717 (O_1717,N_29002,N_29295);
or UO_1718 (O_1718,N_29650,N_29326);
xnor UO_1719 (O_1719,N_29983,N_29374);
xnor UO_1720 (O_1720,N_29408,N_29899);
nor UO_1721 (O_1721,N_29907,N_29522);
and UO_1722 (O_1722,N_29643,N_29593);
nor UO_1723 (O_1723,N_29011,N_29132);
xnor UO_1724 (O_1724,N_29331,N_29501);
xnor UO_1725 (O_1725,N_29971,N_29337);
nor UO_1726 (O_1726,N_29456,N_29486);
and UO_1727 (O_1727,N_29798,N_29955);
nand UO_1728 (O_1728,N_29856,N_29263);
nand UO_1729 (O_1729,N_29188,N_29359);
and UO_1730 (O_1730,N_29770,N_29260);
and UO_1731 (O_1731,N_29870,N_29331);
xor UO_1732 (O_1732,N_29901,N_29629);
xor UO_1733 (O_1733,N_29054,N_29979);
nand UO_1734 (O_1734,N_29069,N_29554);
or UO_1735 (O_1735,N_29748,N_29803);
xnor UO_1736 (O_1736,N_29880,N_29719);
nand UO_1737 (O_1737,N_29762,N_29559);
nand UO_1738 (O_1738,N_29995,N_29653);
and UO_1739 (O_1739,N_29437,N_29150);
nand UO_1740 (O_1740,N_29099,N_29764);
xnor UO_1741 (O_1741,N_29081,N_29516);
nor UO_1742 (O_1742,N_29153,N_29536);
nand UO_1743 (O_1743,N_29071,N_29326);
nand UO_1744 (O_1744,N_29764,N_29686);
and UO_1745 (O_1745,N_29145,N_29613);
and UO_1746 (O_1746,N_29755,N_29085);
nor UO_1747 (O_1747,N_29611,N_29936);
and UO_1748 (O_1748,N_29258,N_29821);
and UO_1749 (O_1749,N_29740,N_29906);
nor UO_1750 (O_1750,N_29217,N_29323);
nand UO_1751 (O_1751,N_29532,N_29063);
or UO_1752 (O_1752,N_29371,N_29461);
nor UO_1753 (O_1753,N_29649,N_29927);
nand UO_1754 (O_1754,N_29314,N_29658);
xor UO_1755 (O_1755,N_29146,N_29100);
nand UO_1756 (O_1756,N_29500,N_29835);
nand UO_1757 (O_1757,N_29496,N_29776);
or UO_1758 (O_1758,N_29411,N_29013);
xnor UO_1759 (O_1759,N_29666,N_29108);
nand UO_1760 (O_1760,N_29969,N_29629);
nand UO_1761 (O_1761,N_29104,N_29679);
and UO_1762 (O_1762,N_29630,N_29035);
xor UO_1763 (O_1763,N_29674,N_29808);
xnor UO_1764 (O_1764,N_29395,N_29466);
nand UO_1765 (O_1765,N_29376,N_29833);
nor UO_1766 (O_1766,N_29376,N_29840);
or UO_1767 (O_1767,N_29223,N_29898);
or UO_1768 (O_1768,N_29375,N_29420);
nor UO_1769 (O_1769,N_29628,N_29720);
nor UO_1770 (O_1770,N_29492,N_29174);
and UO_1771 (O_1771,N_29966,N_29381);
nor UO_1772 (O_1772,N_29784,N_29187);
and UO_1773 (O_1773,N_29082,N_29031);
nor UO_1774 (O_1774,N_29000,N_29635);
nand UO_1775 (O_1775,N_29466,N_29102);
nor UO_1776 (O_1776,N_29378,N_29752);
and UO_1777 (O_1777,N_29816,N_29478);
xor UO_1778 (O_1778,N_29660,N_29483);
and UO_1779 (O_1779,N_29331,N_29759);
and UO_1780 (O_1780,N_29046,N_29659);
xnor UO_1781 (O_1781,N_29026,N_29890);
and UO_1782 (O_1782,N_29391,N_29342);
nand UO_1783 (O_1783,N_29904,N_29424);
or UO_1784 (O_1784,N_29726,N_29636);
or UO_1785 (O_1785,N_29753,N_29407);
nor UO_1786 (O_1786,N_29534,N_29733);
and UO_1787 (O_1787,N_29387,N_29017);
nand UO_1788 (O_1788,N_29374,N_29409);
or UO_1789 (O_1789,N_29485,N_29501);
and UO_1790 (O_1790,N_29986,N_29022);
xnor UO_1791 (O_1791,N_29717,N_29323);
nor UO_1792 (O_1792,N_29077,N_29378);
or UO_1793 (O_1793,N_29977,N_29820);
or UO_1794 (O_1794,N_29631,N_29827);
and UO_1795 (O_1795,N_29825,N_29324);
and UO_1796 (O_1796,N_29887,N_29571);
nor UO_1797 (O_1797,N_29803,N_29609);
and UO_1798 (O_1798,N_29554,N_29790);
xor UO_1799 (O_1799,N_29778,N_29167);
nor UO_1800 (O_1800,N_29752,N_29626);
and UO_1801 (O_1801,N_29779,N_29534);
nand UO_1802 (O_1802,N_29112,N_29206);
and UO_1803 (O_1803,N_29536,N_29168);
and UO_1804 (O_1804,N_29788,N_29824);
or UO_1805 (O_1805,N_29881,N_29898);
xor UO_1806 (O_1806,N_29415,N_29522);
and UO_1807 (O_1807,N_29994,N_29767);
nor UO_1808 (O_1808,N_29243,N_29028);
xor UO_1809 (O_1809,N_29526,N_29026);
and UO_1810 (O_1810,N_29293,N_29081);
nand UO_1811 (O_1811,N_29040,N_29724);
nand UO_1812 (O_1812,N_29114,N_29402);
and UO_1813 (O_1813,N_29261,N_29021);
xor UO_1814 (O_1814,N_29256,N_29840);
and UO_1815 (O_1815,N_29767,N_29713);
nand UO_1816 (O_1816,N_29413,N_29250);
nor UO_1817 (O_1817,N_29709,N_29837);
xnor UO_1818 (O_1818,N_29555,N_29905);
nor UO_1819 (O_1819,N_29533,N_29806);
nor UO_1820 (O_1820,N_29442,N_29508);
nand UO_1821 (O_1821,N_29932,N_29621);
or UO_1822 (O_1822,N_29474,N_29227);
and UO_1823 (O_1823,N_29362,N_29555);
or UO_1824 (O_1824,N_29111,N_29752);
nand UO_1825 (O_1825,N_29420,N_29377);
or UO_1826 (O_1826,N_29607,N_29844);
and UO_1827 (O_1827,N_29031,N_29616);
nor UO_1828 (O_1828,N_29935,N_29373);
or UO_1829 (O_1829,N_29267,N_29015);
or UO_1830 (O_1830,N_29967,N_29812);
nor UO_1831 (O_1831,N_29229,N_29317);
or UO_1832 (O_1832,N_29975,N_29416);
and UO_1833 (O_1833,N_29025,N_29005);
nor UO_1834 (O_1834,N_29922,N_29956);
nor UO_1835 (O_1835,N_29671,N_29154);
nor UO_1836 (O_1836,N_29964,N_29384);
nor UO_1837 (O_1837,N_29856,N_29029);
xor UO_1838 (O_1838,N_29504,N_29456);
nand UO_1839 (O_1839,N_29990,N_29983);
nand UO_1840 (O_1840,N_29391,N_29436);
xor UO_1841 (O_1841,N_29304,N_29587);
nand UO_1842 (O_1842,N_29685,N_29534);
nand UO_1843 (O_1843,N_29417,N_29989);
and UO_1844 (O_1844,N_29013,N_29553);
xnor UO_1845 (O_1845,N_29622,N_29216);
nor UO_1846 (O_1846,N_29689,N_29126);
xor UO_1847 (O_1847,N_29842,N_29289);
or UO_1848 (O_1848,N_29646,N_29912);
nor UO_1849 (O_1849,N_29515,N_29583);
nor UO_1850 (O_1850,N_29333,N_29391);
nor UO_1851 (O_1851,N_29561,N_29312);
and UO_1852 (O_1852,N_29810,N_29729);
and UO_1853 (O_1853,N_29089,N_29315);
and UO_1854 (O_1854,N_29155,N_29900);
and UO_1855 (O_1855,N_29751,N_29968);
and UO_1856 (O_1856,N_29284,N_29287);
nand UO_1857 (O_1857,N_29878,N_29398);
nand UO_1858 (O_1858,N_29407,N_29743);
nor UO_1859 (O_1859,N_29703,N_29793);
nand UO_1860 (O_1860,N_29801,N_29235);
nor UO_1861 (O_1861,N_29070,N_29985);
and UO_1862 (O_1862,N_29257,N_29028);
nor UO_1863 (O_1863,N_29683,N_29732);
or UO_1864 (O_1864,N_29411,N_29580);
xnor UO_1865 (O_1865,N_29190,N_29733);
nand UO_1866 (O_1866,N_29939,N_29708);
or UO_1867 (O_1867,N_29591,N_29107);
and UO_1868 (O_1868,N_29145,N_29783);
nor UO_1869 (O_1869,N_29052,N_29025);
nand UO_1870 (O_1870,N_29787,N_29716);
or UO_1871 (O_1871,N_29295,N_29463);
nand UO_1872 (O_1872,N_29232,N_29387);
or UO_1873 (O_1873,N_29974,N_29661);
nand UO_1874 (O_1874,N_29879,N_29412);
and UO_1875 (O_1875,N_29249,N_29850);
or UO_1876 (O_1876,N_29819,N_29418);
xnor UO_1877 (O_1877,N_29040,N_29069);
nand UO_1878 (O_1878,N_29620,N_29215);
nand UO_1879 (O_1879,N_29408,N_29251);
nor UO_1880 (O_1880,N_29573,N_29811);
nand UO_1881 (O_1881,N_29085,N_29453);
or UO_1882 (O_1882,N_29875,N_29489);
nor UO_1883 (O_1883,N_29318,N_29968);
or UO_1884 (O_1884,N_29148,N_29900);
and UO_1885 (O_1885,N_29971,N_29984);
xor UO_1886 (O_1886,N_29912,N_29431);
and UO_1887 (O_1887,N_29617,N_29338);
or UO_1888 (O_1888,N_29937,N_29286);
xnor UO_1889 (O_1889,N_29644,N_29701);
and UO_1890 (O_1890,N_29880,N_29711);
or UO_1891 (O_1891,N_29806,N_29883);
or UO_1892 (O_1892,N_29612,N_29030);
xnor UO_1893 (O_1893,N_29545,N_29869);
nor UO_1894 (O_1894,N_29827,N_29222);
and UO_1895 (O_1895,N_29201,N_29078);
and UO_1896 (O_1896,N_29421,N_29741);
nand UO_1897 (O_1897,N_29177,N_29278);
nor UO_1898 (O_1898,N_29772,N_29848);
nor UO_1899 (O_1899,N_29695,N_29982);
nand UO_1900 (O_1900,N_29633,N_29630);
and UO_1901 (O_1901,N_29390,N_29203);
nand UO_1902 (O_1902,N_29492,N_29240);
nand UO_1903 (O_1903,N_29600,N_29797);
nor UO_1904 (O_1904,N_29150,N_29448);
or UO_1905 (O_1905,N_29350,N_29204);
xnor UO_1906 (O_1906,N_29468,N_29642);
xnor UO_1907 (O_1907,N_29046,N_29096);
and UO_1908 (O_1908,N_29084,N_29749);
xor UO_1909 (O_1909,N_29667,N_29410);
xnor UO_1910 (O_1910,N_29385,N_29273);
xnor UO_1911 (O_1911,N_29977,N_29708);
or UO_1912 (O_1912,N_29249,N_29527);
or UO_1913 (O_1913,N_29826,N_29876);
nor UO_1914 (O_1914,N_29426,N_29704);
xnor UO_1915 (O_1915,N_29308,N_29201);
xor UO_1916 (O_1916,N_29520,N_29088);
nor UO_1917 (O_1917,N_29299,N_29277);
or UO_1918 (O_1918,N_29307,N_29278);
nand UO_1919 (O_1919,N_29762,N_29044);
or UO_1920 (O_1920,N_29525,N_29942);
and UO_1921 (O_1921,N_29509,N_29190);
nor UO_1922 (O_1922,N_29768,N_29027);
nand UO_1923 (O_1923,N_29304,N_29578);
nand UO_1924 (O_1924,N_29080,N_29574);
or UO_1925 (O_1925,N_29707,N_29854);
and UO_1926 (O_1926,N_29581,N_29256);
nand UO_1927 (O_1927,N_29208,N_29023);
and UO_1928 (O_1928,N_29710,N_29066);
nand UO_1929 (O_1929,N_29749,N_29612);
xnor UO_1930 (O_1930,N_29566,N_29774);
and UO_1931 (O_1931,N_29890,N_29324);
or UO_1932 (O_1932,N_29186,N_29536);
xnor UO_1933 (O_1933,N_29394,N_29086);
nand UO_1934 (O_1934,N_29955,N_29574);
and UO_1935 (O_1935,N_29321,N_29211);
nand UO_1936 (O_1936,N_29056,N_29658);
or UO_1937 (O_1937,N_29159,N_29389);
or UO_1938 (O_1938,N_29027,N_29320);
xnor UO_1939 (O_1939,N_29770,N_29243);
xor UO_1940 (O_1940,N_29068,N_29102);
and UO_1941 (O_1941,N_29095,N_29211);
and UO_1942 (O_1942,N_29855,N_29944);
and UO_1943 (O_1943,N_29395,N_29076);
nand UO_1944 (O_1944,N_29432,N_29883);
and UO_1945 (O_1945,N_29434,N_29095);
nor UO_1946 (O_1946,N_29168,N_29858);
nor UO_1947 (O_1947,N_29863,N_29333);
and UO_1948 (O_1948,N_29589,N_29070);
and UO_1949 (O_1949,N_29623,N_29467);
xor UO_1950 (O_1950,N_29044,N_29278);
nor UO_1951 (O_1951,N_29360,N_29262);
or UO_1952 (O_1952,N_29049,N_29684);
and UO_1953 (O_1953,N_29003,N_29293);
or UO_1954 (O_1954,N_29780,N_29512);
nand UO_1955 (O_1955,N_29376,N_29516);
nand UO_1956 (O_1956,N_29667,N_29303);
or UO_1957 (O_1957,N_29835,N_29572);
or UO_1958 (O_1958,N_29008,N_29189);
and UO_1959 (O_1959,N_29252,N_29028);
or UO_1960 (O_1960,N_29672,N_29149);
or UO_1961 (O_1961,N_29042,N_29866);
or UO_1962 (O_1962,N_29072,N_29618);
and UO_1963 (O_1963,N_29404,N_29944);
xor UO_1964 (O_1964,N_29032,N_29789);
xor UO_1965 (O_1965,N_29134,N_29496);
or UO_1966 (O_1966,N_29574,N_29148);
and UO_1967 (O_1967,N_29462,N_29545);
nor UO_1968 (O_1968,N_29897,N_29326);
nor UO_1969 (O_1969,N_29648,N_29690);
or UO_1970 (O_1970,N_29949,N_29932);
xnor UO_1971 (O_1971,N_29802,N_29164);
and UO_1972 (O_1972,N_29320,N_29716);
or UO_1973 (O_1973,N_29132,N_29979);
nor UO_1974 (O_1974,N_29413,N_29455);
nor UO_1975 (O_1975,N_29054,N_29779);
nor UO_1976 (O_1976,N_29221,N_29337);
nor UO_1977 (O_1977,N_29622,N_29175);
or UO_1978 (O_1978,N_29254,N_29878);
and UO_1979 (O_1979,N_29185,N_29075);
and UO_1980 (O_1980,N_29676,N_29568);
nor UO_1981 (O_1981,N_29912,N_29911);
or UO_1982 (O_1982,N_29459,N_29898);
xor UO_1983 (O_1983,N_29642,N_29905);
nand UO_1984 (O_1984,N_29309,N_29049);
xor UO_1985 (O_1985,N_29817,N_29748);
nor UO_1986 (O_1986,N_29804,N_29165);
nor UO_1987 (O_1987,N_29097,N_29188);
or UO_1988 (O_1988,N_29520,N_29531);
or UO_1989 (O_1989,N_29981,N_29864);
xor UO_1990 (O_1990,N_29516,N_29386);
and UO_1991 (O_1991,N_29175,N_29876);
nand UO_1992 (O_1992,N_29312,N_29684);
nor UO_1993 (O_1993,N_29516,N_29427);
and UO_1994 (O_1994,N_29620,N_29425);
nor UO_1995 (O_1995,N_29164,N_29836);
nand UO_1996 (O_1996,N_29581,N_29552);
xor UO_1997 (O_1997,N_29754,N_29535);
nor UO_1998 (O_1998,N_29934,N_29519);
and UO_1999 (O_1999,N_29469,N_29174);
or UO_2000 (O_2000,N_29414,N_29205);
xor UO_2001 (O_2001,N_29398,N_29548);
and UO_2002 (O_2002,N_29217,N_29205);
nor UO_2003 (O_2003,N_29877,N_29890);
and UO_2004 (O_2004,N_29107,N_29453);
and UO_2005 (O_2005,N_29100,N_29744);
nand UO_2006 (O_2006,N_29274,N_29838);
or UO_2007 (O_2007,N_29351,N_29944);
nor UO_2008 (O_2008,N_29268,N_29541);
or UO_2009 (O_2009,N_29994,N_29375);
xnor UO_2010 (O_2010,N_29630,N_29863);
or UO_2011 (O_2011,N_29313,N_29360);
or UO_2012 (O_2012,N_29820,N_29580);
or UO_2013 (O_2013,N_29844,N_29176);
and UO_2014 (O_2014,N_29766,N_29523);
nor UO_2015 (O_2015,N_29878,N_29742);
or UO_2016 (O_2016,N_29834,N_29726);
xor UO_2017 (O_2017,N_29341,N_29100);
xnor UO_2018 (O_2018,N_29750,N_29088);
or UO_2019 (O_2019,N_29727,N_29253);
nand UO_2020 (O_2020,N_29944,N_29632);
xnor UO_2021 (O_2021,N_29541,N_29761);
and UO_2022 (O_2022,N_29339,N_29518);
xnor UO_2023 (O_2023,N_29672,N_29406);
and UO_2024 (O_2024,N_29672,N_29497);
nor UO_2025 (O_2025,N_29615,N_29006);
nor UO_2026 (O_2026,N_29547,N_29508);
xor UO_2027 (O_2027,N_29942,N_29201);
or UO_2028 (O_2028,N_29489,N_29923);
xor UO_2029 (O_2029,N_29045,N_29630);
or UO_2030 (O_2030,N_29540,N_29368);
nor UO_2031 (O_2031,N_29946,N_29673);
or UO_2032 (O_2032,N_29348,N_29454);
or UO_2033 (O_2033,N_29548,N_29868);
nand UO_2034 (O_2034,N_29054,N_29569);
or UO_2035 (O_2035,N_29055,N_29076);
or UO_2036 (O_2036,N_29590,N_29377);
nand UO_2037 (O_2037,N_29663,N_29424);
xnor UO_2038 (O_2038,N_29864,N_29155);
xor UO_2039 (O_2039,N_29022,N_29193);
nor UO_2040 (O_2040,N_29298,N_29643);
nor UO_2041 (O_2041,N_29082,N_29368);
xnor UO_2042 (O_2042,N_29885,N_29524);
and UO_2043 (O_2043,N_29354,N_29976);
and UO_2044 (O_2044,N_29681,N_29620);
or UO_2045 (O_2045,N_29775,N_29456);
or UO_2046 (O_2046,N_29088,N_29211);
nor UO_2047 (O_2047,N_29715,N_29518);
or UO_2048 (O_2048,N_29810,N_29956);
xor UO_2049 (O_2049,N_29803,N_29829);
nor UO_2050 (O_2050,N_29890,N_29948);
nor UO_2051 (O_2051,N_29116,N_29765);
or UO_2052 (O_2052,N_29910,N_29580);
xnor UO_2053 (O_2053,N_29083,N_29121);
nor UO_2054 (O_2054,N_29296,N_29069);
and UO_2055 (O_2055,N_29167,N_29420);
xor UO_2056 (O_2056,N_29617,N_29591);
and UO_2057 (O_2057,N_29286,N_29679);
nand UO_2058 (O_2058,N_29615,N_29634);
and UO_2059 (O_2059,N_29771,N_29811);
xnor UO_2060 (O_2060,N_29519,N_29770);
xor UO_2061 (O_2061,N_29580,N_29249);
nand UO_2062 (O_2062,N_29464,N_29310);
nor UO_2063 (O_2063,N_29592,N_29348);
and UO_2064 (O_2064,N_29132,N_29462);
xor UO_2065 (O_2065,N_29420,N_29537);
nand UO_2066 (O_2066,N_29533,N_29212);
xor UO_2067 (O_2067,N_29824,N_29814);
xnor UO_2068 (O_2068,N_29507,N_29417);
xnor UO_2069 (O_2069,N_29185,N_29894);
nor UO_2070 (O_2070,N_29794,N_29814);
and UO_2071 (O_2071,N_29157,N_29144);
or UO_2072 (O_2072,N_29129,N_29369);
and UO_2073 (O_2073,N_29551,N_29273);
nand UO_2074 (O_2074,N_29146,N_29729);
xnor UO_2075 (O_2075,N_29936,N_29892);
or UO_2076 (O_2076,N_29441,N_29757);
or UO_2077 (O_2077,N_29686,N_29065);
or UO_2078 (O_2078,N_29910,N_29381);
and UO_2079 (O_2079,N_29226,N_29469);
nand UO_2080 (O_2080,N_29985,N_29656);
nor UO_2081 (O_2081,N_29163,N_29804);
or UO_2082 (O_2082,N_29589,N_29419);
nor UO_2083 (O_2083,N_29239,N_29036);
and UO_2084 (O_2084,N_29478,N_29592);
xnor UO_2085 (O_2085,N_29405,N_29455);
xnor UO_2086 (O_2086,N_29330,N_29148);
xor UO_2087 (O_2087,N_29972,N_29325);
xnor UO_2088 (O_2088,N_29035,N_29020);
or UO_2089 (O_2089,N_29510,N_29560);
nor UO_2090 (O_2090,N_29854,N_29447);
nand UO_2091 (O_2091,N_29772,N_29635);
nand UO_2092 (O_2092,N_29648,N_29769);
nor UO_2093 (O_2093,N_29789,N_29414);
nand UO_2094 (O_2094,N_29938,N_29837);
and UO_2095 (O_2095,N_29426,N_29522);
or UO_2096 (O_2096,N_29960,N_29989);
nor UO_2097 (O_2097,N_29729,N_29567);
nand UO_2098 (O_2098,N_29790,N_29378);
nor UO_2099 (O_2099,N_29609,N_29818);
nor UO_2100 (O_2100,N_29324,N_29508);
nor UO_2101 (O_2101,N_29393,N_29588);
nand UO_2102 (O_2102,N_29535,N_29370);
or UO_2103 (O_2103,N_29452,N_29256);
and UO_2104 (O_2104,N_29645,N_29833);
xor UO_2105 (O_2105,N_29145,N_29411);
and UO_2106 (O_2106,N_29694,N_29740);
or UO_2107 (O_2107,N_29494,N_29075);
and UO_2108 (O_2108,N_29872,N_29108);
nor UO_2109 (O_2109,N_29964,N_29984);
or UO_2110 (O_2110,N_29372,N_29077);
or UO_2111 (O_2111,N_29201,N_29945);
nor UO_2112 (O_2112,N_29243,N_29905);
xor UO_2113 (O_2113,N_29483,N_29528);
or UO_2114 (O_2114,N_29122,N_29997);
xor UO_2115 (O_2115,N_29261,N_29411);
nand UO_2116 (O_2116,N_29030,N_29602);
nor UO_2117 (O_2117,N_29015,N_29045);
xor UO_2118 (O_2118,N_29553,N_29628);
nor UO_2119 (O_2119,N_29298,N_29428);
and UO_2120 (O_2120,N_29579,N_29560);
nor UO_2121 (O_2121,N_29127,N_29020);
xnor UO_2122 (O_2122,N_29806,N_29382);
and UO_2123 (O_2123,N_29516,N_29605);
nand UO_2124 (O_2124,N_29101,N_29118);
xor UO_2125 (O_2125,N_29065,N_29525);
xnor UO_2126 (O_2126,N_29872,N_29254);
nor UO_2127 (O_2127,N_29149,N_29990);
or UO_2128 (O_2128,N_29543,N_29709);
nor UO_2129 (O_2129,N_29995,N_29718);
nand UO_2130 (O_2130,N_29483,N_29608);
nor UO_2131 (O_2131,N_29198,N_29862);
nand UO_2132 (O_2132,N_29238,N_29621);
nor UO_2133 (O_2133,N_29438,N_29470);
or UO_2134 (O_2134,N_29776,N_29495);
xnor UO_2135 (O_2135,N_29477,N_29542);
xor UO_2136 (O_2136,N_29262,N_29033);
nand UO_2137 (O_2137,N_29831,N_29005);
nor UO_2138 (O_2138,N_29123,N_29575);
or UO_2139 (O_2139,N_29267,N_29029);
nor UO_2140 (O_2140,N_29386,N_29748);
xnor UO_2141 (O_2141,N_29566,N_29768);
nand UO_2142 (O_2142,N_29271,N_29575);
and UO_2143 (O_2143,N_29807,N_29763);
nand UO_2144 (O_2144,N_29548,N_29838);
nor UO_2145 (O_2145,N_29118,N_29797);
nor UO_2146 (O_2146,N_29342,N_29291);
xnor UO_2147 (O_2147,N_29655,N_29030);
and UO_2148 (O_2148,N_29213,N_29336);
and UO_2149 (O_2149,N_29753,N_29659);
or UO_2150 (O_2150,N_29766,N_29349);
nand UO_2151 (O_2151,N_29995,N_29864);
xor UO_2152 (O_2152,N_29641,N_29970);
or UO_2153 (O_2153,N_29550,N_29676);
and UO_2154 (O_2154,N_29495,N_29949);
and UO_2155 (O_2155,N_29310,N_29277);
xor UO_2156 (O_2156,N_29554,N_29226);
and UO_2157 (O_2157,N_29169,N_29481);
nor UO_2158 (O_2158,N_29268,N_29915);
xor UO_2159 (O_2159,N_29394,N_29061);
nor UO_2160 (O_2160,N_29851,N_29549);
nor UO_2161 (O_2161,N_29389,N_29837);
and UO_2162 (O_2162,N_29810,N_29324);
and UO_2163 (O_2163,N_29356,N_29545);
and UO_2164 (O_2164,N_29710,N_29874);
and UO_2165 (O_2165,N_29036,N_29582);
and UO_2166 (O_2166,N_29517,N_29130);
or UO_2167 (O_2167,N_29694,N_29949);
nand UO_2168 (O_2168,N_29437,N_29301);
nand UO_2169 (O_2169,N_29591,N_29856);
nand UO_2170 (O_2170,N_29898,N_29025);
and UO_2171 (O_2171,N_29644,N_29905);
or UO_2172 (O_2172,N_29567,N_29257);
nor UO_2173 (O_2173,N_29284,N_29436);
xnor UO_2174 (O_2174,N_29696,N_29084);
nor UO_2175 (O_2175,N_29424,N_29543);
nand UO_2176 (O_2176,N_29478,N_29866);
xnor UO_2177 (O_2177,N_29975,N_29831);
nor UO_2178 (O_2178,N_29606,N_29507);
nand UO_2179 (O_2179,N_29965,N_29005);
or UO_2180 (O_2180,N_29628,N_29430);
nand UO_2181 (O_2181,N_29820,N_29610);
xnor UO_2182 (O_2182,N_29277,N_29119);
nand UO_2183 (O_2183,N_29039,N_29811);
nor UO_2184 (O_2184,N_29814,N_29646);
xnor UO_2185 (O_2185,N_29283,N_29219);
or UO_2186 (O_2186,N_29718,N_29106);
xnor UO_2187 (O_2187,N_29808,N_29017);
nand UO_2188 (O_2188,N_29382,N_29141);
nand UO_2189 (O_2189,N_29279,N_29401);
xnor UO_2190 (O_2190,N_29417,N_29083);
and UO_2191 (O_2191,N_29338,N_29044);
nand UO_2192 (O_2192,N_29544,N_29597);
or UO_2193 (O_2193,N_29120,N_29273);
and UO_2194 (O_2194,N_29353,N_29169);
xnor UO_2195 (O_2195,N_29605,N_29146);
nor UO_2196 (O_2196,N_29985,N_29592);
or UO_2197 (O_2197,N_29841,N_29922);
xor UO_2198 (O_2198,N_29527,N_29279);
and UO_2199 (O_2199,N_29842,N_29347);
and UO_2200 (O_2200,N_29513,N_29339);
nand UO_2201 (O_2201,N_29813,N_29538);
nor UO_2202 (O_2202,N_29403,N_29264);
nand UO_2203 (O_2203,N_29283,N_29455);
nand UO_2204 (O_2204,N_29476,N_29217);
nor UO_2205 (O_2205,N_29913,N_29193);
nor UO_2206 (O_2206,N_29775,N_29729);
xor UO_2207 (O_2207,N_29401,N_29744);
nand UO_2208 (O_2208,N_29666,N_29620);
nor UO_2209 (O_2209,N_29371,N_29536);
xnor UO_2210 (O_2210,N_29406,N_29515);
nand UO_2211 (O_2211,N_29539,N_29508);
nand UO_2212 (O_2212,N_29403,N_29497);
and UO_2213 (O_2213,N_29149,N_29675);
nand UO_2214 (O_2214,N_29607,N_29641);
and UO_2215 (O_2215,N_29067,N_29764);
and UO_2216 (O_2216,N_29879,N_29822);
or UO_2217 (O_2217,N_29423,N_29104);
or UO_2218 (O_2218,N_29167,N_29890);
nor UO_2219 (O_2219,N_29207,N_29588);
nor UO_2220 (O_2220,N_29900,N_29958);
xnor UO_2221 (O_2221,N_29790,N_29701);
and UO_2222 (O_2222,N_29249,N_29004);
or UO_2223 (O_2223,N_29386,N_29663);
nor UO_2224 (O_2224,N_29650,N_29524);
or UO_2225 (O_2225,N_29092,N_29135);
or UO_2226 (O_2226,N_29137,N_29395);
nor UO_2227 (O_2227,N_29277,N_29450);
xnor UO_2228 (O_2228,N_29359,N_29082);
or UO_2229 (O_2229,N_29182,N_29633);
nor UO_2230 (O_2230,N_29459,N_29213);
nor UO_2231 (O_2231,N_29132,N_29570);
or UO_2232 (O_2232,N_29859,N_29451);
nor UO_2233 (O_2233,N_29828,N_29491);
and UO_2234 (O_2234,N_29945,N_29772);
and UO_2235 (O_2235,N_29099,N_29655);
xor UO_2236 (O_2236,N_29858,N_29935);
or UO_2237 (O_2237,N_29216,N_29357);
or UO_2238 (O_2238,N_29930,N_29829);
nor UO_2239 (O_2239,N_29605,N_29167);
or UO_2240 (O_2240,N_29837,N_29148);
nand UO_2241 (O_2241,N_29624,N_29395);
xor UO_2242 (O_2242,N_29373,N_29929);
xnor UO_2243 (O_2243,N_29185,N_29800);
nor UO_2244 (O_2244,N_29294,N_29007);
or UO_2245 (O_2245,N_29870,N_29742);
nor UO_2246 (O_2246,N_29556,N_29860);
and UO_2247 (O_2247,N_29114,N_29532);
and UO_2248 (O_2248,N_29437,N_29760);
or UO_2249 (O_2249,N_29140,N_29335);
and UO_2250 (O_2250,N_29129,N_29412);
nor UO_2251 (O_2251,N_29887,N_29443);
or UO_2252 (O_2252,N_29541,N_29107);
nor UO_2253 (O_2253,N_29698,N_29795);
xnor UO_2254 (O_2254,N_29017,N_29050);
or UO_2255 (O_2255,N_29675,N_29150);
xnor UO_2256 (O_2256,N_29869,N_29832);
nor UO_2257 (O_2257,N_29490,N_29686);
and UO_2258 (O_2258,N_29310,N_29536);
or UO_2259 (O_2259,N_29383,N_29164);
nand UO_2260 (O_2260,N_29373,N_29090);
or UO_2261 (O_2261,N_29979,N_29739);
nand UO_2262 (O_2262,N_29521,N_29691);
nor UO_2263 (O_2263,N_29234,N_29957);
or UO_2264 (O_2264,N_29333,N_29550);
xnor UO_2265 (O_2265,N_29798,N_29349);
xor UO_2266 (O_2266,N_29735,N_29629);
or UO_2267 (O_2267,N_29680,N_29806);
nor UO_2268 (O_2268,N_29533,N_29328);
or UO_2269 (O_2269,N_29659,N_29271);
nand UO_2270 (O_2270,N_29023,N_29933);
or UO_2271 (O_2271,N_29408,N_29603);
nor UO_2272 (O_2272,N_29186,N_29469);
nor UO_2273 (O_2273,N_29409,N_29962);
nor UO_2274 (O_2274,N_29356,N_29559);
nand UO_2275 (O_2275,N_29144,N_29608);
xnor UO_2276 (O_2276,N_29987,N_29965);
nand UO_2277 (O_2277,N_29842,N_29532);
or UO_2278 (O_2278,N_29272,N_29529);
nor UO_2279 (O_2279,N_29571,N_29147);
nor UO_2280 (O_2280,N_29871,N_29867);
or UO_2281 (O_2281,N_29307,N_29659);
nor UO_2282 (O_2282,N_29064,N_29700);
or UO_2283 (O_2283,N_29068,N_29973);
and UO_2284 (O_2284,N_29381,N_29843);
xnor UO_2285 (O_2285,N_29020,N_29353);
nor UO_2286 (O_2286,N_29487,N_29266);
nor UO_2287 (O_2287,N_29998,N_29548);
nor UO_2288 (O_2288,N_29700,N_29340);
nor UO_2289 (O_2289,N_29296,N_29649);
and UO_2290 (O_2290,N_29702,N_29434);
nor UO_2291 (O_2291,N_29338,N_29815);
nand UO_2292 (O_2292,N_29491,N_29471);
xor UO_2293 (O_2293,N_29311,N_29866);
and UO_2294 (O_2294,N_29395,N_29923);
nor UO_2295 (O_2295,N_29249,N_29603);
and UO_2296 (O_2296,N_29797,N_29206);
xnor UO_2297 (O_2297,N_29009,N_29023);
nand UO_2298 (O_2298,N_29687,N_29061);
and UO_2299 (O_2299,N_29997,N_29870);
or UO_2300 (O_2300,N_29855,N_29319);
nand UO_2301 (O_2301,N_29115,N_29591);
nand UO_2302 (O_2302,N_29220,N_29942);
or UO_2303 (O_2303,N_29946,N_29670);
and UO_2304 (O_2304,N_29141,N_29446);
nand UO_2305 (O_2305,N_29416,N_29223);
and UO_2306 (O_2306,N_29954,N_29561);
xnor UO_2307 (O_2307,N_29951,N_29354);
nand UO_2308 (O_2308,N_29840,N_29404);
and UO_2309 (O_2309,N_29850,N_29335);
nor UO_2310 (O_2310,N_29206,N_29280);
xor UO_2311 (O_2311,N_29988,N_29047);
nand UO_2312 (O_2312,N_29911,N_29575);
xor UO_2313 (O_2313,N_29633,N_29915);
and UO_2314 (O_2314,N_29553,N_29044);
nor UO_2315 (O_2315,N_29579,N_29232);
xor UO_2316 (O_2316,N_29931,N_29824);
or UO_2317 (O_2317,N_29382,N_29841);
xnor UO_2318 (O_2318,N_29486,N_29567);
or UO_2319 (O_2319,N_29129,N_29398);
nand UO_2320 (O_2320,N_29285,N_29879);
or UO_2321 (O_2321,N_29098,N_29315);
xor UO_2322 (O_2322,N_29948,N_29235);
nand UO_2323 (O_2323,N_29373,N_29154);
and UO_2324 (O_2324,N_29413,N_29389);
xor UO_2325 (O_2325,N_29892,N_29051);
nor UO_2326 (O_2326,N_29352,N_29563);
nor UO_2327 (O_2327,N_29527,N_29173);
nand UO_2328 (O_2328,N_29604,N_29858);
or UO_2329 (O_2329,N_29100,N_29925);
or UO_2330 (O_2330,N_29054,N_29903);
nand UO_2331 (O_2331,N_29612,N_29002);
nand UO_2332 (O_2332,N_29082,N_29893);
xnor UO_2333 (O_2333,N_29998,N_29553);
nor UO_2334 (O_2334,N_29301,N_29509);
nand UO_2335 (O_2335,N_29647,N_29081);
or UO_2336 (O_2336,N_29899,N_29390);
nand UO_2337 (O_2337,N_29680,N_29044);
nor UO_2338 (O_2338,N_29505,N_29336);
nand UO_2339 (O_2339,N_29419,N_29021);
nand UO_2340 (O_2340,N_29660,N_29452);
nor UO_2341 (O_2341,N_29385,N_29450);
xor UO_2342 (O_2342,N_29932,N_29022);
nand UO_2343 (O_2343,N_29799,N_29355);
nand UO_2344 (O_2344,N_29619,N_29516);
nand UO_2345 (O_2345,N_29578,N_29815);
or UO_2346 (O_2346,N_29710,N_29036);
nor UO_2347 (O_2347,N_29590,N_29791);
or UO_2348 (O_2348,N_29828,N_29248);
or UO_2349 (O_2349,N_29521,N_29909);
nor UO_2350 (O_2350,N_29895,N_29312);
nand UO_2351 (O_2351,N_29532,N_29698);
and UO_2352 (O_2352,N_29171,N_29671);
and UO_2353 (O_2353,N_29360,N_29480);
nand UO_2354 (O_2354,N_29993,N_29463);
or UO_2355 (O_2355,N_29292,N_29926);
xnor UO_2356 (O_2356,N_29742,N_29939);
nor UO_2357 (O_2357,N_29723,N_29984);
nand UO_2358 (O_2358,N_29033,N_29144);
nor UO_2359 (O_2359,N_29744,N_29510);
xor UO_2360 (O_2360,N_29507,N_29481);
xnor UO_2361 (O_2361,N_29972,N_29274);
or UO_2362 (O_2362,N_29443,N_29155);
xor UO_2363 (O_2363,N_29749,N_29305);
and UO_2364 (O_2364,N_29157,N_29845);
nand UO_2365 (O_2365,N_29935,N_29786);
nor UO_2366 (O_2366,N_29981,N_29186);
nand UO_2367 (O_2367,N_29871,N_29156);
and UO_2368 (O_2368,N_29924,N_29322);
nor UO_2369 (O_2369,N_29253,N_29946);
nor UO_2370 (O_2370,N_29429,N_29180);
nor UO_2371 (O_2371,N_29620,N_29180);
xnor UO_2372 (O_2372,N_29494,N_29583);
or UO_2373 (O_2373,N_29307,N_29176);
and UO_2374 (O_2374,N_29454,N_29184);
and UO_2375 (O_2375,N_29573,N_29692);
xor UO_2376 (O_2376,N_29571,N_29962);
nor UO_2377 (O_2377,N_29953,N_29156);
or UO_2378 (O_2378,N_29623,N_29673);
nand UO_2379 (O_2379,N_29346,N_29408);
or UO_2380 (O_2380,N_29867,N_29284);
nand UO_2381 (O_2381,N_29614,N_29043);
or UO_2382 (O_2382,N_29728,N_29166);
xnor UO_2383 (O_2383,N_29587,N_29906);
or UO_2384 (O_2384,N_29046,N_29580);
and UO_2385 (O_2385,N_29976,N_29574);
nor UO_2386 (O_2386,N_29528,N_29367);
or UO_2387 (O_2387,N_29322,N_29735);
or UO_2388 (O_2388,N_29432,N_29047);
nand UO_2389 (O_2389,N_29115,N_29654);
xor UO_2390 (O_2390,N_29625,N_29411);
xor UO_2391 (O_2391,N_29019,N_29404);
and UO_2392 (O_2392,N_29365,N_29651);
nand UO_2393 (O_2393,N_29917,N_29694);
or UO_2394 (O_2394,N_29419,N_29866);
and UO_2395 (O_2395,N_29349,N_29502);
or UO_2396 (O_2396,N_29020,N_29852);
nand UO_2397 (O_2397,N_29087,N_29231);
nor UO_2398 (O_2398,N_29500,N_29144);
or UO_2399 (O_2399,N_29441,N_29984);
nand UO_2400 (O_2400,N_29850,N_29225);
and UO_2401 (O_2401,N_29378,N_29412);
and UO_2402 (O_2402,N_29318,N_29944);
nor UO_2403 (O_2403,N_29906,N_29015);
or UO_2404 (O_2404,N_29052,N_29418);
nand UO_2405 (O_2405,N_29047,N_29224);
xnor UO_2406 (O_2406,N_29840,N_29688);
or UO_2407 (O_2407,N_29674,N_29885);
or UO_2408 (O_2408,N_29064,N_29353);
nand UO_2409 (O_2409,N_29428,N_29670);
xor UO_2410 (O_2410,N_29802,N_29339);
nor UO_2411 (O_2411,N_29905,N_29908);
nor UO_2412 (O_2412,N_29356,N_29680);
xor UO_2413 (O_2413,N_29950,N_29810);
xor UO_2414 (O_2414,N_29151,N_29915);
nand UO_2415 (O_2415,N_29378,N_29349);
nand UO_2416 (O_2416,N_29103,N_29857);
or UO_2417 (O_2417,N_29333,N_29989);
nand UO_2418 (O_2418,N_29312,N_29861);
nand UO_2419 (O_2419,N_29011,N_29440);
or UO_2420 (O_2420,N_29635,N_29546);
xor UO_2421 (O_2421,N_29168,N_29123);
nand UO_2422 (O_2422,N_29307,N_29206);
nand UO_2423 (O_2423,N_29956,N_29362);
nor UO_2424 (O_2424,N_29329,N_29817);
nor UO_2425 (O_2425,N_29910,N_29634);
xor UO_2426 (O_2426,N_29442,N_29833);
and UO_2427 (O_2427,N_29072,N_29578);
nor UO_2428 (O_2428,N_29267,N_29959);
nand UO_2429 (O_2429,N_29121,N_29667);
nand UO_2430 (O_2430,N_29713,N_29509);
nor UO_2431 (O_2431,N_29740,N_29799);
or UO_2432 (O_2432,N_29477,N_29785);
nand UO_2433 (O_2433,N_29999,N_29026);
nor UO_2434 (O_2434,N_29049,N_29508);
nor UO_2435 (O_2435,N_29652,N_29864);
nand UO_2436 (O_2436,N_29511,N_29960);
or UO_2437 (O_2437,N_29838,N_29101);
and UO_2438 (O_2438,N_29343,N_29867);
xnor UO_2439 (O_2439,N_29854,N_29570);
nand UO_2440 (O_2440,N_29661,N_29479);
or UO_2441 (O_2441,N_29029,N_29911);
xor UO_2442 (O_2442,N_29047,N_29608);
or UO_2443 (O_2443,N_29806,N_29061);
and UO_2444 (O_2444,N_29746,N_29486);
and UO_2445 (O_2445,N_29432,N_29795);
or UO_2446 (O_2446,N_29500,N_29065);
xor UO_2447 (O_2447,N_29173,N_29218);
nand UO_2448 (O_2448,N_29500,N_29914);
xor UO_2449 (O_2449,N_29481,N_29023);
nand UO_2450 (O_2450,N_29054,N_29017);
or UO_2451 (O_2451,N_29158,N_29238);
and UO_2452 (O_2452,N_29807,N_29846);
nor UO_2453 (O_2453,N_29172,N_29457);
nor UO_2454 (O_2454,N_29802,N_29374);
or UO_2455 (O_2455,N_29671,N_29585);
and UO_2456 (O_2456,N_29150,N_29200);
nor UO_2457 (O_2457,N_29288,N_29425);
or UO_2458 (O_2458,N_29330,N_29163);
xor UO_2459 (O_2459,N_29439,N_29077);
and UO_2460 (O_2460,N_29828,N_29659);
nor UO_2461 (O_2461,N_29478,N_29027);
or UO_2462 (O_2462,N_29801,N_29187);
and UO_2463 (O_2463,N_29945,N_29382);
nand UO_2464 (O_2464,N_29921,N_29879);
nor UO_2465 (O_2465,N_29437,N_29563);
or UO_2466 (O_2466,N_29838,N_29915);
nor UO_2467 (O_2467,N_29054,N_29088);
xnor UO_2468 (O_2468,N_29255,N_29858);
nor UO_2469 (O_2469,N_29989,N_29058);
xor UO_2470 (O_2470,N_29567,N_29755);
and UO_2471 (O_2471,N_29552,N_29056);
nor UO_2472 (O_2472,N_29698,N_29797);
and UO_2473 (O_2473,N_29874,N_29311);
nor UO_2474 (O_2474,N_29732,N_29203);
xnor UO_2475 (O_2475,N_29477,N_29974);
and UO_2476 (O_2476,N_29952,N_29635);
nand UO_2477 (O_2477,N_29447,N_29472);
and UO_2478 (O_2478,N_29776,N_29854);
or UO_2479 (O_2479,N_29545,N_29023);
nand UO_2480 (O_2480,N_29934,N_29109);
or UO_2481 (O_2481,N_29527,N_29958);
or UO_2482 (O_2482,N_29958,N_29122);
xnor UO_2483 (O_2483,N_29921,N_29316);
nand UO_2484 (O_2484,N_29386,N_29276);
nor UO_2485 (O_2485,N_29938,N_29734);
xor UO_2486 (O_2486,N_29819,N_29897);
or UO_2487 (O_2487,N_29126,N_29967);
xnor UO_2488 (O_2488,N_29490,N_29717);
and UO_2489 (O_2489,N_29065,N_29970);
nand UO_2490 (O_2490,N_29290,N_29171);
xnor UO_2491 (O_2491,N_29086,N_29028);
nor UO_2492 (O_2492,N_29087,N_29417);
nand UO_2493 (O_2493,N_29666,N_29157);
xnor UO_2494 (O_2494,N_29907,N_29169);
xnor UO_2495 (O_2495,N_29865,N_29235);
nand UO_2496 (O_2496,N_29765,N_29473);
or UO_2497 (O_2497,N_29655,N_29907);
xnor UO_2498 (O_2498,N_29229,N_29249);
xnor UO_2499 (O_2499,N_29730,N_29420);
nand UO_2500 (O_2500,N_29588,N_29127);
nand UO_2501 (O_2501,N_29403,N_29617);
and UO_2502 (O_2502,N_29916,N_29922);
and UO_2503 (O_2503,N_29361,N_29630);
xnor UO_2504 (O_2504,N_29217,N_29807);
nor UO_2505 (O_2505,N_29982,N_29915);
nand UO_2506 (O_2506,N_29510,N_29644);
nor UO_2507 (O_2507,N_29911,N_29883);
and UO_2508 (O_2508,N_29782,N_29970);
nand UO_2509 (O_2509,N_29858,N_29501);
and UO_2510 (O_2510,N_29275,N_29980);
nand UO_2511 (O_2511,N_29424,N_29362);
or UO_2512 (O_2512,N_29813,N_29049);
or UO_2513 (O_2513,N_29425,N_29233);
and UO_2514 (O_2514,N_29502,N_29354);
nand UO_2515 (O_2515,N_29550,N_29485);
nor UO_2516 (O_2516,N_29835,N_29501);
or UO_2517 (O_2517,N_29000,N_29778);
nor UO_2518 (O_2518,N_29733,N_29161);
nand UO_2519 (O_2519,N_29380,N_29866);
or UO_2520 (O_2520,N_29853,N_29683);
nor UO_2521 (O_2521,N_29567,N_29434);
and UO_2522 (O_2522,N_29780,N_29181);
nand UO_2523 (O_2523,N_29946,N_29487);
and UO_2524 (O_2524,N_29130,N_29073);
nor UO_2525 (O_2525,N_29462,N_29112);
or UO_2526 (O_2526,N_29378,N_29357);
or UO_2527 (O_2527,N_29531,N_29656);
or UO_2528 (O_2528,N_29815,N_29140);
and UO_2529 (O_2529,N_29947,N_29294);
nor UO_2530 (O_2530,N_29723,N_29040);
and UO_2531 (O_2531,N_29884,N_29121);
nor UO_2532 (O_2532,N_29444,N_29873);
nand UO_2533 (O_2533,N_29288,N_29775);
or UO_2534 (O_2534,N_29613,N_29500);
xnor UO_2535 (O_2535,N_29999,N_29659);
or UO_2536 (O_2536,N_29041,N_29390);
or UO_2537 (O_2537,N_29863,N_29862);
and UO_2538 (O_2538,N_29717,N_29057);
nand UO_2539 (O_2539,N_29474,N_29609);
xnor UO_2540 (O_2540,N_29022,N_29904);
or UO_2541 (O_2541,N_29728,N_29223);
nor UO_2542 (O_2542,N_29089,N_29210);
or UO_2543 (O_2543,N_29307,N_29766);
and UO_2544 (O_2544,N_29461,N_29735);
xor UO_2545 (O_2545,N_29908,N_29806);
nand UO_2546 (O_2546,N_29550,N_29590);
nand UO_2547 (O_2547,N_29217,N_29814);
nor UO_2548 (O_2548,N_29361,N_29192);
xor UO_2549 (O_2549,N_29446,N_29010);
and UO_2550 (O_2550,N_29685,N_29600);
nand UO_2551 (O_2551,N_29162,N_29758);
xor UO_2552 (O_2552,N_29116,N_29008);
xnor UO_2553 (O_2553,N_29892,N_29562);
nor UO_2554 (O_2554,N_29970,N_29730);
xnor UO_2555 (O_2555,N_29030,N_29418);
or UO_2556 (O_2556,N_29346,N_29994);
and UO_2557 (O_2557,N_29654,N_29326);
or UO_2558 (O_2558,N_29969,N_29896);
nand UO_2559 (O_2559,N_29441,N_29653);
xor UO_2560 (O_2560,N_29643,N_29623);
xnor UO_2561 (O_2561,N_29463,N_29501);
nor UO_2562 (O_2562,N_29590,N_29451);
xor UO_2563 (O_2563,N_29726,N_29531);
xnor UO_2564 (O_2564,N_29117,N_29813);
nand UO_2565 (O_2565,N_29794,N_29784);
or UO_2566 (O_2566,N_29257,N_29595);
nor UO_2567 (O_2567,N_29836,N_29250);
xnor UO_2568 (O_2568,N_29443,N_29539);
nor UO_2569 (O_2569,N_29139,N_29259);
and UO_2570 (O_2570,N_29314,N_29308);
xor UO_2571 (O_2571,N_29129,N_29089);
nor UO_2572 (O_2572,N_29287,N_29112);
or UO_2573 (O_2573,N_29435,N_29136);
or UO_2574 (O_2574,N_29625,N_29359);
nor UO_2575 (O_2575,N_29264,N_29641);
and UO_2576 (O_2576,N_29225,N_29710);
nand UO_2577 (O_2577,N_29888,N_29368);
or UO_2578 (O_2578,N_29333,N_29173);
nor UO_2579 (O_2579,N_29814,N_29323);
or UO_2580 (O_2580,N_29834,N_29284);
xor UO_2581 (O_2581,N_29340,N_29044);
or UO_2582 (O_2582,N_29673,N_29430);
or UO_2583 (O_2583,N_29981,N_29076);
xor UO_2584 (O_2584,N_29602,N_29253);
and UO_2585 (O_2585,N_29211,N_29105);
nand UO_2586 (O_2586,N_29935,N_29609);
or UO_2587 (O_2587,N_29078,N_29085);
nand UO_2588 (O_2588,N_29052,N_29363);
nand UO_2589 (O_2589,N_29812,N_29821);
xor UO_2590 (O_2590,N_29338,N_29211);
or UO_2591 (O_2591,N_29767,N_29655);
or UO_2592 (O_2592,N_29690,N_29113);
or UO_2593 (O_2593,N_29501,N_29542);
nand UO_2594 (O_2594,N_29264,N_29927);
nor UO_2595 (O_2595,N_29930,N_29110);
nand UO_2596 (O_2596,N_29042,N_29614);
and UO_2597 (O_2597,N_29518,N_29025);
xnor UO_2598 (O_2598,N_29477,N_29727);
xnor UO_2599 (O_2599,N_29327,N_29706);
nand UO_2600 (O_2600,N_29620,N_29386);
and UO_2601 (O_2601,N_29836,N_29579);
nor UO_2602 (O_2602,N_29679,N_29999);
xnor UO_2603 (O_2603,N_29485,N_29033);
xnor UO_2604 (O_2604,N_29364,N_29335);
and UO_2605 (O_2605,N_29191,N_29397);
nor UO_2606 (O_2606,N_29450,N_29184);
or UO_2607 (O_2607,N_29824,N_29096);
xnor UO_2608 (O_2608,N_29174,N_29965);
nor UO_2609 (O_2609,N_29889,N_29041);
xnor UO_2610 (O_2610,N_29451,N_29230);
xor UO_2611 (O_2611,N_29436,N_29345);
xor UO_2612 (O_2612,N_29479,N_29291);
and UO_2613 (O_2613,N_29845,N_29807);
and UO_2614 (O_2614,N_29867,N_29676);
nand UO_2615 (O_2615,N_29639,N_29472);
and UO_2616 (O_2616,N_29740,N_29672);
or UO_2617 (O_2617,N_29377,N_29535);
nand UO_2618 (O_2618,N_29567,N_29152);
and UO_2619 (O_2619,N_29086,N_29071);
nand UO_2620 (O_2620,N_29493,N_29745);
nand UO_2621 (O_2621,N_29522,N_29358);
nand UO_2622 (O_2622,N_29354,N_29642);
nor UO_2623 (O_2623,N_29763,N_29865);
nor UO_2624 (O_2624,N_29681,N_29001);
nor UO_2625 (O_2625,N_29071,N_29915);
nand UO_2626 (O_2626,N_29029,N_29252);
or UO_2627 (O_2627,N_29988,N_29233);
nor UO_2628 (O_2628,N_29892,N_29460);
xor UO_2629 (O_2629,N_29901,N_29121);
xnor UO_2630 (O_2630,N_29657,N_29653);
xnor UO_2631 (O_2631,N_29234,N_29100);
nand UO_2632 (O_2632,N_29211,N_29665);
nor UO_2633 (O_2633,N_29876,N_29156);
nor UO_2634 (O_2634,N_29912,N_29073);
nand UO_2635 (O_2635,N_29797,N_29362);
xor UO_2636 (O_2636,N_29816,N_29443);
xor UO_2637 (O_2637,N_29709,N_29184);
nor UO_2638 (O_2638,N_29286,N_29708);
nand UO_2639 (O_2639,N_29307,N_29080);
or UO_2640 (O_2640,N_29302,N_29471);
nand UO_2641 (O_2641,N_29903,N_29409);
or UO_2642 (O_2642,N_29223,N_29952);
or UO_2643 (O_2643,N_29806,N_29890);
nand UO_2644 (O_2644,N_29111,N_29020);
nor UO_2645 (O_2645,N_29940,N_29196);
or UO_2646 (O_2646,N_29142,N_29766);
xnor UO_2647 (O_2647,N_29892,N_29026);
and UO_2648 (O_2648,N_29628,N_29137);
and UO_2649 (O_2649,N_29590,N_29178);
xor UO_2650 (O_2650,N_29367,N_29963);
or UO_2651 (O_2651,N_29829,N_29054);
nand UO_2652 (O_2652,N_29939,N_29094);
xnor UO_2653 (O_2653,N_29074,N_29177);
or UO_2654 (O_2654,N_29725,N_29266);
xnor UO_2655 (O_2655,N_29774,N_29120);
and UO_2656 (O_2656,N_29451,N_29390);
nor UO_2657 (O_2657,N_29362,N_29509);
or UO_2658 (O_2658,N_29089,N_29898);
xnor UO_2659 (O_2659,N_29811,N_29636);
and UO_2660 (O_2660,N_29577,N_29882);
or UO_2661 (O_2661,N_29653,N_29964);
nand UO_2662 (O_2662,N_29956,N_29266);
and UO_2663 (O_2663,N_29316,N_29516);
or UO_2664 (O_2664,N_29919,N_29954);
nand UO_2665 (O_2665,N_29374,N_29312);
and UO_2666 (O_2666,N_29221,N_29477);
xnor UO_2667 (O_2667,N_29571,N_29394);
xnor UO_2668 (O_2668,N_29144,N_29253);
nand UO_2669 (O_2669,N_29462,N_29494);
nor UO_2670 (O_2670,N_29442,N_29682);
and UO_2671 (O_2671,N_29945,N_29475);
nor UO_2672 (O_2672,N_29517,N_29507);
and UO_2673 (O_2673,N_29178,N_29028);
and UO_2674 (O_2674,N_29692,N_29814);
xnor UO_2675 (O_2675,N_29301,N_29395);
and UO_2676 (O_2676,N_29574,N_29430);
nand UO_2677 (O_2677,N_29593,N_29817);
or UO_2678 (O_2678,N_29280,N_29904);
nand UO_2679 (O_2679,N_29025,N_29412);
and UO_2680 (O_2680,N_29617,N_29934);
nor UO_2681 (O_2681,N_29851,N_29417);
nor UO_2682 (O_2682,N_29295,N_29311);
or UO_2683 (O_2683,N_29028,N_29605);
nor UO_2684 (O_2684,N_29502,N_29484);
and UO_2685 (O_2685,N_29206,N_29029);
xor UO_2686 (O_2686,N_29041,N_29542);
and UO_2687 (O_2687,N_29037,N_29626);
and UO_2688 (O_2688,N_29788,N_29456);
nor UO_2689 (O_2689,N_29748,N_29398);
nor UO_2690 (O_2690,N_29991,N_29987);
xor UO_2691 (O_2691,N_29325,N_29596);
or UO_2692 (O_2692,N_29022,N_29696);
and UO_2693 (O_2693,N_29025,N_29463);
nand UO_2694 (O_2694,N_29980,N_29458);
nand UO_2695 (O_2695,N_29584,N_29466);
nand UO_2696 (O_2696,N_29793,N_29724);
or UO_2697 (O_2697,N_29448,N_29298);
xnor UO_2698 (O_2698,N_29340,N_29839);
or UO_2699 (O_2699,N_29634,N_29004);
xor UO_2700 (O_2700,N_29061,N_29762);
or UO_2701 (O_2701,N_29640,N_29845);
nand UO_2702 (O_2702,N_29125,N_29800);
and UO_2703 (O_2703,N_29649,N_29121);
nand UO_2704 (O_2704,N_29787,N_29525);
or UO_2705 (O_2705,N_29183,N_29899);
and UO_2706 (O_2706,N_29538,N_29869);
or UO_2707 (O_2707,N_29082,N_29270);
xor UO_2708 (O_2708,N_29925,N_29718);
nor UO_2709 (O_2709,N_29405,N_29615);
or UO_2710 (O_2710,N_29142,N_29497);
and UO_2711 (O_2711,N_29537,N_29451);
xor UO_2712 (O_2712,N_29072,N_29084);
xnor UO_2713 (O_2713,N_29032,N_29037);
xnor UO_2714 (O_2714,N_29719,N_29405);
nand UO_2715 (O_2715,N_29533,N_29427);
and UO_2716 (O_2716,N_29519,N_29760);
or UO_2717 (O_2717,N_29794,N_29196);
and UO_2718 (O_2718,N_29042,N_29794);
xor UO_2719 (O_2719,N_29241,N_29815);
and UO_2720 (O_2720,N_29683,N_29081);
and UO_2721 (O_2721,N_29402,N_29288);
nand UO_2722 (O_2722,N_29276,N_29359);
nand UO_2723 (O_2723,N_29332,N_29951);
or UO_2724 (O_2724,N_29060,N_29879);
nor UO_2725 (O_2725,N_29346,N_29710);
or UO_2726 (O_2726,N_29811,N_29477);
nor UO_2727 (O_2727,N_29881,N_29613);
nor UO_2728 (O_2728,N_29295,N_29662);
nor UO_2729 (O_2729,N_29883,N_29697);
nor UO_2730 (O_2730,N_29348,N_29390);
nor UO_2731 (O_2731,N_29031,N_29099);
and UO_2732 (O_2732,N_29204,N_29757);
nor UO_2733 (O_2733,N_29728,N_29290);
and UO_2734 (O_2734,N_29118,N_29956);
nand UO_2735 (O_2735,N_29718,N_29329);
or UO_2736 (O_2736,N_29758,N_29453);
nor UO_2737 (O_2737,N_29921,N_29583);
xnor UO_2738 (O_2738,N_29288,N_29589);
nor UO_2739 (O_2739,N_29238,N_29540);
nor UO_2740 (O_2740,N_29474,N_29217);
or UO_2741 (O_2741,N_29068,N_29618);
or UO_2742 (O_2742,N_29866,N_29708);
and UO_2743 (O_2743,N_29833,N_29001);
xor UO_2744 (O_2744,N_29879,N_29193);
and UO_2745 (O_2745,N_29881,N_29389);
nand UO_2746 (O_2746,N_29043,N_29410);
or UO_2747 (O_2747,N_29057,N_29629);
nand UO_2748 (O_2748,N_29993,N_29572);
and UO_2749 (O_2749,N_29966,N_29231);
nand UO_2750 (O_2750,N_29403,N_29647);
nor UO_2751 (O_2751,N_29728,N_29312);
and UO_2752 (O_2752,N_29225,N_29525);
or UO_2753 (O_2753,N_29926,N_29992);
nor UO_2754 (O_2754,N_29512,N_29233);
nand UO_2755 (O_2755,N_29785,N_29496);
or UO_2756 (O_2756,N_29762,N_29595);
and UO_2757 (O_2757,N_29019,N_29469);
nor UO_2758 (O_2758,N_29671,N_29194);
nor UO_2759 (O_2759,N_29840,N_29285);
or UO_2760 (O_2760,N_29386,N_29363);
nand UO_2761 (O_2761,N_29535,N_29644);
nor UO_2762 (O_2762,N_29306,N_29036);
xnor UO_2763 (O_2763,N_29418,N_29878);
and UO_2764 (O_2764,N_29696,N_29981);
and UO_2765 (O_2765,N_29149,N_29591);
nand UO_2766 (O_2766,N_29291,N_29752);
nor UO_2767 (O_2767,N_29498,N_29208);
xor UO_2768 (O_2768,N_29999,N_29214);
and UO_2769 (O_2769,N_29453,N_29890);
xnor UO_2770 (O_2770,N_29566,N_29769);
nand UO_2771 (O_2771,N_29563,N_29016);
and UO_2772 (O_2772,N_29045,N_29745);
nand UO_2773 (O_2773,N_29227,N_29909);
and UO_2774 (O_2774,N_29470,N_29725);
nor UO_2775 (O_2775,N_29895,N_29893);
xor UO_2776 (O_2776,N_29883,N_29419);
nand UO_2777 (O_2777,N_29209,N_29676);
nand UO_2778 (O_2778,N_29642,N_29275);
or UO_2779 (O_2779,N_29153,N_29456);
nor UO_2780 (O_2780,N_29493,N_29261);
nor UO_2781 (O_2781,N_29553,N_29513);
nand UO_2782 (O_2782,N_29185,N_29664);
and UO_2783 (O_2783,N_29332,N_29698);
nor UO_2784 (O_2784,N_29262,N_29857);
nand UO_2785 (O_2785,N_29419,N_29059);
and UO_2786 (O_2786,N_29510,N_29220);
or UO_2787 (O_2787,N_29065,N_29628);
and UO_2788 (O_2788,N_29006,N_29695);
or UO_2789 (O_2789,N_29045,N_29309);
and UO_2790 (O_2790,N_29086,N_29376);
nand UO_2791 (O_2791,N_29218,N_29767);
xnor UO_2792 (O_2792,N_29663,N_29474);
and UO_2793 (O_2793,N_29698,N_29388);
xnor UO_2794 (O_2794,N_29906,N_29822);
or UO_2795 (O_2795,N_29538,N_29597);
xor UO_2796 (O_2796,N_29242,N_29452);
and UO_2797 (O_2797,N_29841,N_29722);
and UO_2798 (O_2798,N_29352,N_29529);
xor UO_2799 (O_2799,N_29082,N_29740);
nand UO_2800 (O_2800,N_29929,N_29846);
or UO_2801 (O_2801,N_29514,N_29515);
nor UO_2802 (O_2802,N_29697,N_29367);
nand UO_2803 (O_2803,N_29081,N_29282);
nand UO_2804 (O_2804,N_29604,N_29881);
and UO_2805 (O_2805,N_29923,N_29771);
or UO_2806 (O_2806,N_29573,N_29677);
nor UO_2807 (O_2807,N_29731,N_29809);
xnor UO_2808 (O_2808,N_29814,N_29717);
or UO_2809 (O_2809,N_29398,N_29551);
nand UO_2810 (O_2810,N_29755,N_29965);
and UO_2811 (O_2811,N_29906,N_29813);
and UO_2812 (O_2812,N_29569,N_29430);
nor UO_2813 (O_2813,N_29592,N_29848);
or UO_2814 (O_2814,N_29419,N_29931);
nor UO_2815 (O_2815,N_29446,N_29593);
nand UO_2816 (O_2816,N_29241,N_29745);
and UO_2817 (O_2817,N_29882,N_29935);
or UO_2818 (O_2818,N_29470,N_29530);
and UO_2819 (O_2819,N_29923,N_29603);
xnor UO_2820 (O_2820,N_29057,N_29766);
nor UO_2821 (O_2821,N_29437,N_29777);
xor UO_2822 (O_2822,N_29934,N_29740);
and UO_2823 (O_2823,N_29240,N_29150);
or UO_2824 (O_2824,N_29320,N_29338);
nor UO_2825 (O_2825,N_29628,N_29068);
nor UO_2826 (O_2826,N_29696,N_29288);
nor UO_2827 (O_2827,N_29981,N_29391);
or UO_2828 (O_2828,N_29984,N_29950);
or UO_2829 (O_2829,N_29014,N_29583);
nand UO_2830 (O_2830,N_29661,N_29205);
nor UO_2831 (O_2831,N_29431,N_29631);
xnor UO_2832 (O_2832,N_29826,N_29732);
and UO_2833 (O_2833,N_29442,N_29130);
nand UO_2834 (O_2834,N_29691,N_29068);
nor UO_2835 (O_2835,N_29672,N_29296);
or UO_2836 (O_2836,N_29563,N_29151);
nand UO_2837 (O_2837,N_29632,N_29085);
nand UO_2838 (O_2838,N_29361,N_29394);
nand UO_2839 (O_2839,N_29818,N_29416);
nand UO_2840 (O_2840,N_29277,N_29295);
nor UO_2841 (O_2841,N_29852,N_29877);
or UO_2842 (O_2842,N_29960,N_29868);
nand UO_2843 (O_2843,N_29891,N_29308);
xor UO_2844 (O_2844,N_29462,N_29823);
and UO_2845 (O_2845,N_29699,N_29211);
and UO_2846 (O_2846,N_29950,N_29330);
nor UO_2847 (O_2847,N_29897,N_29824);
or UO_2848 (O_2848,N_29317,N_29632);
xor UO_2849 (O_2849,N_29322,N_29436);
xor UO_2850 (O_2850,N_29858,N_29430);
or UO_2851 (O_2851,N_29774,N_29674);
or UO_2852 (O_2852,N_29584,N_29727);
xor UO_2853 (O_2853,N_29458,N_29927);
nand UO_2854 (O_2854,N_29105,N_29688);
xor UO_2855 (O_2855,N_29661,N_29467);
and UO_2856 (O_2856,N_29280,N_29011);
nor UO_2857 (O_2857,N_29244,N_29367);
nor UO_2858 (O_2858,N_29066,N_29949);
nand UO_2859 (O_2859,N_29483,N_29433);
nand UO_2860 (O_2860,N_29250,N_29078);
xor UO_2861 (O_2861,N_29364,N_29862);
nor UO_2862 (O_2862,N_29928,N_29610);
and UO_2863 (O_2863,N_29074,N_29100);
nand UO_2864 (O_2864,N_29158,N_29292);
and UO_2865 (O_2865,N_29770,N_29649);
nand UO_2866 (O_2866,N_29156,N_29708);
or UO_2867 (O_2867,N_29946,N_29052);
nand UO_2868 (O_2868,N_29766,N_29246);
and UO_2869 (O_2869,N_29075,N_29902);
xnor UO_2870 (O_2870,N_29113,N_29743);
nor UO_2871 (O_2871,N_29310,N_29214);
and UO_2872 (O_2872,N_29823,N_29726);
xor UO_2873 (O_2873,N_29570,N_29942);
nor UO_2874 (O_2874,N_29686,N_29669);
xnor UO_2875 (O_2875,N_29415,N_29619);
or UO_2876 (O_2876,N_29990,N_29409);
xnor UO_2877 (O_2877,N_29893,N_29800);
nor UO_2878 (O_2878,N_29649,N_29609);
nand UO_2879 (O_2879,N_29261,N_29704);
or UO_2880 (O_2880,N_29854,N_29586);
or UO_2881 (O_2881,N_29005,N_29826);
nand UO_2882 (O_2882,N_29350,N_29449);
or UO_2883 (O_2883,N_29262,N_29882);
nand UO_2884 (O_2884,N_29291,N_29920);
and UO_2885 (O_2885,N_29322,N_29698);
nand UO_2886 (O_2886,N_29344,N_29154);
nor UO_2887 (O_2887,N_29513,N_29241);
nor UO_2888 (O_2888,N_29099,N_29119);
nand UO_2889 (O_2889,N_29511,N_29781);
xor UO_2890 (O_2890,N_29442,N_29222);
or UO_2891 (O_2891,N_29669,N_29665);
nand UO_2892 (O_2892,N_29230,N_29258);
or UO_2893 (O_2893,N_29818,N_29467);
and UO_2894 (O_2894,N_29357,N_29787);
xor UO_2895 (O_2895,N_29551,N_29211);
and UO_2896 (O_2896,N_29733,N_29674);
and UO_2897 (O_2897,N_29828,N_29604);
xnor UO_2898 (O_2898,N_29785,N_29916);
nor UO_2899 (O_2899,N_29637,N_29355);
xnor UO_2900 (O_2900,N_29415,N_29272);
nor UO_2901 (O_2901,N_29635,N_29905);
xor UO_2902 (O_2902,N_29202,N_29524);
xor UO_2903 (O_2903,N_29923,N_29609);
xor UO_2904 (O_2904,N_29470,N_29440);
or UO_2905 (O_2905,N_29066,N_29927);
or UO_2906 (O_2906,N_29905,N_29563);
xnor UO_2907 (O_2907,N_29584,N_29050);
or UO_2908 (O_2908,N_29783,N_29003);
xor UO_2909 (O_2909,N_29031,N_29535);
nor UO_2910 (O_2910,N_29815,N_29068);
or UO_2911 (O_2911,N_29623,N_29298);
xnor UO_2912 (O_2912,N_29804,N_29960);
xor UO_2913 (O_2913,N_29339,N_29195);
and UO_2914 (O_2914,N_29903,N_29913);
and UO_2915 (O_2915,N_29039,N_29691);
nand UO_2916 (O_2916,N_29312,N_29041);
and UO_2917 (O_2917,N_29878,N_29996);
and UO_2918 (O_2918,N_29717,N_29382);
nor UO_2919 (O_2919,N_29961,N_29435);
or UO_2920 (O_2920,N_29823,N_29382);
xor UO_2921 (O_2921,N_29455,N_29647);
or UO_2922 (O_2922,N_29844,N_29661);
or UO_2923 (O_2923,N_29737,N_29222);
or UO_2924 (O_2924,N_29459,N_29223);
xnor UO_2925 (O_2925,N_29080,N_29818);
nor UO_2926 (O_2926,N_29264,N_29132);
nand UO_2927 (O_2927,N_29121,N_29698);
nand UO_2928 (O_2928,N_29083,N_29236);
or UO_2929 (O_2929,N_29143,N_29266);
nand UO_2930 (O_2930,N_29949,N_29458);
nor UO_2931 (O_2931,N_29070,N_29367);
nand UO_2932 (O_2932,N_29485,N_29767);
nor UO_2933 (O_2933,N_29807,N_29326);
nand UO_2934 (O_2934,N_29038,N_29868);
xor UO_2935 (O_2935,N_29682,N_29881);
and UO_2936 (O_2936,N_29688,N_29013);
nand UO_2937 (O_2937,N_29320,N_29682);
nand UO_2938 (O_2938,N_29807,N_29374);
and UO_2939 (O_2939,N_29896,N_29337);
and UO_2940 (O_2940,N_29914,N_29756);
and UO_2941 (O_2941,N_29877,N_29821);
and UO_2942 (O_2942,N_29861,N_29211);
nor UO_2943 (O_2943,N_29067,N_29098);
and UO_2944 (O_2944,N_29241,N_29009);
xnor UO_2945 (O_2945,N_29586,N_29649);
or UO_2946 (O_2946,N_29701,N_29742);
or UO_2947 (O_2947,N_29197,N_29809);
nand UO_2948 (O_2948,N_29327,N_29061);
nor UO_2949 (O_2949,N_29706,N_29040);
or UO_2950 (O_2950,N_29349,N_29906);
nor UO_2951 (O_2951,N_29019,N_29312);
nand UO_2952 (O_2952,N_29528,N_29863);
nor UO_2953 (O_2953,N_29650,N_29217);
xor UO_2954 (O_2954,N_29773,N_29553);
and UO_2955 (O_2955,N_29591,N_29143);
nor UO_2956 (O_2956,N_29017,N_29366);
or UO_2957 (O_2957,N_29912,N_29585);
and UO_2958 (O_2958,N_29175,N_29088);
nor UO_2959 (O_2959,N_29729,N_29800);
nand UO_2960 (O_2960,N_29855,N_29128);
and UO_2961 (O_2961,N_29144,N_29288);
xor UO_2962 (O_2962,N_29345,N_29524);
and UO_2963 (O_2963,N_29645,N_29425);
and UO_2964 (O_2964,N_29703,N_29795);
xnor UO_2965 (O_2965,N_29054,N_29714);
and UO_2966 (O_2966,N_29000,N_29927);
nand UO_2967 (O_2967,N_29327,N_29714);
or UO_2968 (O_2968,N_29510,N_29961);
nand UO_2969 (O_2969,N_29566,N_29952);
nand UO_2970 (O_2970,N_29670,N_29414);
or UO_2971 (O_2971,N_29528,N_29494);
or UO_2972 (O_2972,N_29677,N_29750);
or UO_2973 (O_2973,N_29440,N_29077);
xor UO_2974 (O_2974,N_29680,N_29318);
nor UO_2975 (O_2975,N_29383,N_29893);
or UO_2976 (O_2976,N_29341,N_29716);
and UO_2977 (O_2977,N_29212,N_29672);
nand UO_2978 (O_2978,N_29144,N_29271);
xnor UO_2979 (O_2979,N_29327,N_29772);
nor UO_2980 (O_2980,N_29205,N_29626);
and UO_2981 (O_2981,N_29517,N_29622);
nand UO_2982 (O_2982,N_29667,N_29819);
nand UO_2983 (O_2983,N_29368,N_29312);
xor UO_2984 (O_2984,N_29868,N_29965);
nand UO_2985 (O_2985,N_29135,N_29771);
or UO_2986 (O_2986,N_29144,N_29963);
nor UO_2987 (O_2987,N_29101,N_29428);
or UO_2988 (O_2988,N_29979,N_29445);
nor UO_2989 (O_2989,N_29438,N_29018);
nand UO_2990 (O_2990,N_29380,N_29536);
and UO_2991 (O_2991,N_29105,N_29322);
and UO_2992 (O_2992,N_29476,N_29053);
and UO_2993 (O_2993,N_29559,N_29696);
and UO_2994 (O_2994,N_29261,N_29792);
nand UO_2995 (O_2995,N_29155,N_29701);
nor UO_2996 (O_2996,N_29907,N_29117);
or UO_2997 (O_2997,N_29933,N_29274);
or UO_2998 (O_2998,N_29955,N_29987);
or UO_2999 (O_2999,N_29757,N_29743);
xor UO_3000 (O_3000,N_29453,N_29609);
nor UO_3001 (O_3001,N_29417,N_29198);
and UO_3002 (O_3002,N_29106,N_29282);
xor UO_3003 (O_3003,N_29507,N_29634);
xnor UO_3004 (O_3004,N_29839,N_29214);
nor UO_3005 (O_3005,N_29647,N_29661);
xnor UO_3006 (O_3006,N_29499,N_29881);
nor UO_3007 (O_3007,N_29788,N_29793);
nor UO_3008 (O_3008,N_29390,N_29957);
nor UO_3009 (O_3009,N_29731,N_29768);
nand UO_3010 (O_3010,N_29664,N_29563);
xor UO_3011 (O_3011,N_29536,N_29929);
xor UO_3012 (O_3012,N_29161,N_29858);
and UO_3013 (O_3013,N_29194,N_29058);
nor UO_3014 (O_3014,N_29023,N_29222);
nand UO_3015 (O_3015,N_29342,N_29187);
nand UO_3016 (O_3016,N_29660,N_29993);
xnor UO_3017 (O_3017,N_29161,N_29452);
xnor UO_3018 (O_3018,N_29820,N_29691);
or UO_3019 (O_3019,N_29127,N_29495);
or UO_3020 (O_3020,N_29249,N_29747);
nand UO_3021 (O_3021,N_29737,N_29930);
or UO_3022 (O_3022,N_29603,N_29549);
and UO_3023 (O_3023,N_29645,N_29073);
and UO_3024 (O_3024,N_29825,N_29183);
nand UO_3025 (O_3025,N_29438,N_29382);
nand UO_3026 (O_3026,N_29392,N_29501);
nand UO_3027 (O_3027,N_29366,N_29709);
and UO_3028 (O_3028,N_29224,N_29505);
nor UO_3029 (O_3029,N_29365,N_29165);
nand UO_3030 (O_3030,N_29334,N_29030);
nand UO_3031 (O_3031,N_29072,N_29390);
or UO_3032 (O_3032,N_29403,N_29629);
nor UO_3033 (O_3033,N_29898,N_29415);
xor UO_3034 (O_3034,N_29473,N_29930);
xnor UO_3035 (O_3035,N_29719,N_29867);
nand UO_3036 (O_3036,N_29115,N_29948);
and UO_3037 (O_3037,N_29889,N_29141);
nor UO_3038 (O_3038,N_29122,N_29891);
xnor UO_3039 (O_3039,N_29996,N_29012);
nand UO_3040 (O_3040,N_29718,N_29557);
nor UO_3041 (O_3041,N_29057,N_29029);
nand UO_3042 (O_3042,N_29259,N_29767);
and UO_3043 (O_3043,N_29540,N_29986);
or UO_3044 (O_3044,N_29429,N_29066);
xnor UO_3045 (O_3045,N_29367,N_29967);
nand UO_3046 (O_3046,N_29059,N_29622);
or UO_3047 (O_3047,N_29859,N_29032);
and UO_3048 (O_3048,N_29324,N_29548);
xnor UO_3049 (O_3049,N_29766,N_29832);
nand UO_3050 (O_3050,N_29900,N_29321);
and UO_3051 (O_3051,N_29478,N_29714);
or UO_3052 (O_3052,N_29847,N_29287);
nand UO_3053 (O_3053,N_29670,N_29844);
and UO_3054 (O_3054,N_29592,N_29540);
nand UO_3055 (O_3055,N_29815,N_29376);
and UO_3056 (O_3056,N_29771,N_29375);
nand UO_3057 (O_3057,N_29065,N_29812);
nor UO_3058 (O_3058,N_29025,N_29781);
nand UO_3059 (O_3059,N_29554,N_29200);
nand UO_3060 (O_3060,N_29550,N_29461);
nand UO_3061 (O_3061,N_29210,N_29924);
xnor UO_3062 (O_3062,N_29012,N_29503);
nand UO_3063 (O_3063,N_29891,N_29759);
and UO_3064 (O_3064,N_29448,N_29457);
nor UO_3065 (O_3065,N_29531,N_29326);
xor UO_3066 (O_3066,N_29588,N_29797);
nor UO_3067 (O_3067,N_29472,N_29024);
and UO_3068 (O_3068,N_29011,N_29924);
and UO_3069 (O_3069,N_29083,N_29316);
or UO_3070 (O_3070,N_29045,N_29339);
nand UO_3071 (O_3071,N_29404,N_29645);
or UO_3072 (O_3072,N_29494,N_29760);
and UO_3073 (O_3073,N_29542,N_29289);
nand UO_3074 (O_3074,N_29881,N_29941);
nand UO_3075 (O_3075,N_29861,N_29620);
nor UO_3076 (O_3076,N_29656,N_29595);
and UO_3077 (O_3077,N_29565,N_29953);
or UO_3078 (O_3078,N_29538,N_29235);
and UO_3079 (O_3079,N_29387,N_29641);
xnor UO_3080 (O_3080,N_29898,N_29666);
or UO_3081 (O_3081,N_29363,N_29501);
nand UO_3082 (O_3082,N_29591,N_29795);
and UO_3083 (O_3083,N_29908,N_29606);
xor UO_3084 (O_3084,N_29121,N_29586);
and UO_3085 (O_3085,N_29723,N_29785);
nand UO_3086 (O_3086,N_29099,N_29141);
or UO_3087 (O_3087,N_29543,N_29903);
or UO_3088 (O_3088,N_29736,N_29337);
and UO_3089 (O_3089,N_29737,N_29878);
and UO_3090 (O_3090,N_29456,N_29395);
or UO_3091 (O_3091,N_29284,N_29439);
or UO_3092 (O_3092,N_29557,N_29878);
or UO_3093 (O_3093,N_29985,N_29118);
nor UO_3094 (O_3094,N_29777,N_29145);
or UO_3095 (O_3095,N_29761,N_29310);
or UO_3096 (O_3096,N_29296,N_29892);
and UO_3097 (O_3097,N_29201,N_29295);
or UO_3098 (O_3098,N_29573,N_29823);
nand UO_3099 (O_3099,N_29775,N_29204);
or UO_3100 (O_3100,N_29576,N_29203);
or UO_3101 (O_3101,N_29019,N_29310);
nor UO_3102 (O_3102,N_29842,N_29210);
and UO_3103 (O_3103,N_29333,N_29148);
xor UO_3104 (O_3104,N_29002,N_29180);
xor UO_3105 (O_3105,N_29423,N_29840);
or UO_3106 (O_3106,N_29297,N_29688);
and UO_3107 (O_3107,N_29758,N_29655);
nand UO_3108 (O_3108,N_29753,N_29586);
and UO_3109 (O_3109,N_29659,N_29591);
and UO_3110 (O_3110,N_29492,N_29145);
nor UO_3111 (O_3111,N_29525,N_29646);
nand UO_3112 (O_3112,N_29624,N_29891);
nor UO_3113 (O_3113,N_29052,N_29656);
and UO_3114 (O_3114,N_29815,N_29595);
or UO_3115 (O_3115,N_29004,N_29607);
and UO_3116 (O_3116,N_29075,N_29748);
nand UO_3117 (O_3117,N_29845,N_29536);
or UO_3118 (O_3118,N_29083,N_29344);
or UO_3119 (O_3119,N_29151,N_29350);
or UO_3120 (O_3120,N_29027,N_29350);
nand UO_3121 (O_3121,N_29031,N_29810);
or UO_3122 (O_3122,N_29692,N_29048);
and UO_3123 (O_3123,N_29192,N_29914);
nand UO_3124 (O_3124,N_29911,N_29769);
nand UO_3125 (O_3125,N_29278,N_29211);
nand UO_3126 (O_3126,N_29227,N_29871);
and UO_3127 (O_3127,N_29250,N_29861);
nor UO_3128 (O_3128,N_29435,N_29347);
or UO_3129 (O_3129,N_29259,N_29399);
or UO_3130 (O_3130,N_29037,N_29770);
or UO_3131 (O_3131,N_29718,N_29423);
nand UO_3132 (O_3132,N_29169,N_29593);
nor UO_3133 (O_3133,N_29567,N_29284);
and UO_3134 (O_3134,N_29918,N_29975);
xnor UO_3135 (O_3135,N_29762,N_29082);
xor UO_3136 (O_3136,N_29643,N_29731);
xnor UO_3137 (O_3137,N_29562,N_29763);
nand UO_3138 (O_3138,N_29913,N_29174);
nor UO_3139 (O_3139,N_29051,N_29657);
and UO_3140 (O_3140,N_29115,N_29790);
xnor UO_3141 (O_3141,N_29229,N_29005);
xnor UO_3142 (O_3142,N_29032,N_29331);
nand UO_3143 (O_3143,N_29979,N_29346);
nand UO_3144 (O_3144,N_29338,N_29085);
and UO_3145 (O_3145,N_29001,N_29967);
or UO_3146 (O_3146,N_29491,N_29687);
and UO_3147 (O_3147,N_29074,N_29699);
nand UO_3148 (O_3148,N_29606,N_29520);
nand UO_3149 (O_3149,N_29627,N_29578);
xor UO_3150 (O_3150,N_29402,N_29457);
or UO_3151 (O_3151,N_29831,N_29351);
and UO_3152 (O_3152,N_29943,N_29438);
and UO_3153 (O_3153,N_29063,N_29310);
or UO_3154 (O_3154,N_29897,N_29992);
xor UO_3155 (O_3155,N_29543,N_29472);
nand UO_3156 (O_3156,N_29629,N_29806);
xnor UO_3157 (O_3157,N_29188,N_29376);
nand UO_3158 (O_3158,N_29935,N_29849);
nand UO_3159 (O_3159,N_29834,N_29665);
nand UO_3160 (O_3160,N_29215,N_29964);
nand UO_3161 (O_3161,N_29292,N_29934);
nor UO_3162 (O_3162,N_29538,N_29337);
nand UO_3163 (O_3163,N_29589,N_29719);
nor UO_3164 (O_3164,N_29938,N_29566);
nor UO_3165 (O_3165,N_29072,N_29356);
nand UO_3166 (O_3166,N_29496,N_29843);
or UO_3167 (O_3167,N_29703,N_29866);
xor UO_3168 (O_3168,N_29221,N_29536);
nor UO_3169 (O_3169,N_29849,N_29350);
nor UO_3170 (O_3170,N_29015,N_29331);
or UO_3171 (O_3171,N_29611,N_29584);
nor UO_3172 (O_3172,N_29184,N_29311);
nor UO_3173 (O_3173,N_29823,N_29077);
nand UO_3174 (O_3174,N_29692,N_29083);
xor UO_3175 (O_3175,N_29727,N_29281);
nor UO_3176 (O_3176,N_29026,N_29113);
or UO_3177 (O_3177,N_29120,N_29818);
nor UO_3178 (O_3178,N_29220,N_29692);
xor UO_3179 (O_3179,N_29282,N_29309);
xnor UO_3180 (O_3180,N_29286,N_29221);
nor UO_3181 (O_3181,N_29772,N_29260);
or UO_3182 (O_3182,N_29111,N_29140);
nor UO_3183 (O_3183,N_29281,N_29564);
or UO_3184 (O_3184,N_29857,N_29206);
nand UO_3185 (O_3185,N_29881,N_29532);
and UO_3186 (O_3186,N_29298,N_29688);
xnor UO_3187 (O_3187,N_29468,N_29414);
nand UO_3188 (O_3188,N_29222,N_29343);
or UO_3189 (O_3189,N_29363,N_29768);
nor UO_3190 (O_3190,N_29922,N_29879);
nor UO_3191 (O_3191,N_29361,N_29379);
and UO_3192 (O_3192,N_29567,N_29258);
nand UO_3193 (O_3193,N_29341,N_29551);
and UO_3194 (O_3194,N_29391,N_29874);
xnor UO_3195 (O_3195,N_29706,N_29717);
xnor UO_3196 (O_3196,N_29043,N_29293);
or UO_3197 (O_3197,N_29853,N_29602);
or UO_3198 (O_3198,N_29900,N_29072);
xnor UO_3199 (O_3199,N_29308,N_29538);
nand UO_3200 (O_3200,N_29777,N_29311);
nand UO_3201 (O_3201,N_29646,N_29315);
nand UO_3202 (O_3202,N_29658,N_29393);
nor UO_3203 (O_3203,N_29269,N_29494);
xnor UO_3204 (O_3204,N_29517,N_29720);
and UO_3205 (O_3205,N_29046,N_29098);
xor UO_3206 (O_3206,N_29168,N_29367);
or UO_3207 (O_3207,N_29728,N_29443);
xnor UO_3208 (O_3208,N_29403,N_29869);
nand UO_3209 (O_3209,N_29168,N_29369);
nand UO_3210 (O_3210,N_29268,N_29921);
xor UO_3211 (O_3211,N_29940,N_29802);
xnor UO_3212 (O_3212,N_29554,N_29693);
xor UO_3213 (O_3213,N_29583,N_29153);
and UO_3214 (O_3214,N_29750,N_29735);
nand UO_3215 (O_3215,N_29189,N_29280);
and UO_3216 (O_3216,N_29639,N_29060);
nand UO_3217 (O_3217,N_29622,N_29901);
and UO_3218 (O_3218,N_29412,N_29488);
and UO_3219 (O_3219,N_29421,N_29281);
nand UO_3220 (O_3220,N_29433,N_29218);
or UO_3221 (O_3221,N_29526,N_29924);
and UO_3222 (O_3222,N_29816,N_29588);
nand UO_3223 (O_3223,N_29255,N_29600);
nand UO_3224 (O_3224,N_29101,N_29587);
nor UO_3225 (O_3225,N_29502,N_29282);
nand UO_3226 (O_3226,N_29797,N_29392);
nor UO_3227 (O_3227,N_29382,N_29835);
nor UO_3228 (O_3228,N_29903,N_29366);
or UO_3229 (O_3229,N_29220,N_29711);
or UO_3230 (O_3230,N_29101,N_29416);
xor UO_3231 (O_3231,N_29799,N_29200);
nand UO_3232 (O_3232,N_29839,N_29527);
and UO_3233 (O_3233,N_29172,N_29742);
or UO_3234 (O_3234,N_29183,N_29733);
nand UO_3235 (O_3235,N_29660,N_29394);
xor UO_3236 (O_3236,N_29054,N_29573);
nand UO_3237 (O_3237,N_29058,N_29434);
nor UO_3238 (O_3238,N_29443,N_29920);
or UO_3239 (O_3239,N_29325,N_29292);
nand UO_3240 (O_3240,N_29056,N_29319);
xor UO_3241 (O_3241,N_29305,N_29990);
nand UO_3242 (O_3242,N_29013,N_29972);
nand UO_3243 (O_3243,N_29889,N_29641);
xor UO_3244 (O_3244,N_29868,N_29676);
or UO_3245 (O_3245,N_29595,N_29345);
and UO_3246 (O_3246,N_29414,N_29681);
nand UO_3247 (O_3247,N_29317,N_29449);
xor UO_3248 (O_3248,N_29361,N_29562);
xor UO_3249 (O_3249,N_29665,N_29492);
xnor UO_3250 (O_3250,N_29731,N_29598);
or UO_3251 (O_3251,N_29313,N_29771);
nor UO_3252 (O_3252,N_29482,N_29896);
or UO_3253 (O_3253,N_29019,N_29423);
nor UO_3254 (O_3254,N_29155,N_29821);
and UO_3255 (O_3255,N_29924,N_29600);
nand UO_3256 (O_3256,N_29193,N_29330);
or UO_3257 (O_3257,N_29024,N_29777);
nor UO_3258 (O_3258,N_29309,N_29520);
and UO_3259 (O_3259,N_29023,N_29017);
nand UO_3260 (O_3260,N_29016,N_29581);
or UO_3261 (O_3261,N_29849,N_29429);
and UO_3262 (O_3262,N_29713,N_29798);
or UO_3263 (O_3263,N_29713,N_29547);
or UO_3264 (O_3264,N_29388,N_29069);
xor UO_3265 (O_3265,N_29770,N_29755);
nor UO_3266 (O_3266,N_29259,N_29677);
nand UO_3267 (O_3267,N_29816,N_29554);
nor UO_3268 (O_3268,N_29915,N_29752);
or UO_3269 (O_3269,N_29351,N_29821);
xnor UO_3270 (O_3270,N_29534,N_29750);
and UO_3271 (O_3271,N_29358,N_29248);
xor UO_3272 (O_3272,N_29237,N_29313);
or UO_3273 (O_3273,N_29456,N_29939);
xor UO_3274 (O_3274,N_29586,N_29077);
nor UO_3275 (O_3275,N_29074,N_29240);
xor UO_3276 (O_3276,N_29577,N_29636);
and UO_3277 (O_3277,N_29317,N_29447);
xor UO_3278 (O_3278,N_29353,N_29200);
and UO_3279 (O_3279,N_29124,N_29326);
or UO_3280 (O_3280,N_29287,N_29784);
and UO_3281 (O_3281,N_29317,N_29056);
xor UO_3282 (O_3282,N_29727,N_29797);
nor UO_3283 (O_3283,N_29040,N_29782);
and UO_3284 (O_3284,N_29170,N_29603);
xnor UO_3285 (O_3285,N_29019,N_29035);
and UO_3286 (O_3286,N_29383,N_29618);
and UO_3287 (O_3287,N_29133,N_29960);
nand UO_3288 (O_3288,N_29908,N_29467);
and UO_3289 (O_3289,N_29489,N_29768);
and UO_3290 (O_3290,N_29841,N_29046);
and UO_3291 (O_3291,N_29813,N_29397);
nand UO_3292 (O_3292,N_29747,N_29499);
nand UO_3293 (O_3293,N_29428,N_29720);
and UO_3294 (O_3294,N_29847,N_29357);
and UO_3295 (O_3295,N_29623,N_29058);
or UO_3296 (O_3296,N_29667,N_29264);
nand UO_3297 (O_3297,N_29977,N_29125);
xnor UO_3298 (O_3298,N_29909,N_29828);
xor UO_3299 (O_3299,N_29428,N_29403);
or UO_3300 (O_3300,N_29239,N_29140);
nand UO_3301 (O_3301,N_29675,N_29060);
nand UO_3302 (O_3302,N_29633,N_29255);
xor UO_3303 (O_3303,N_29382,N_29151);
nor UO_3304 (O_3304,N_29325,N_29617);
or UO_3305 (O_3305,N_29426,N_29165);
nor UO_3306 (O_3306,N_29100,N_29018);
and UO_3307 (O_3307,N_29073,N_29065);
and UO_3308 (O_3308,N_29093,N_29800);
and UO_3309 (O_3309,N_29339,N_29366);
xnor UO_3310 (O_3310,N_29266,N_29640);
xor UO_3311 (O_3311,N_29747,N_29991);
nor UO_3312 (O_3312,N_29492,N_29825);
xnor UO_3313 (O_3313,N_29862,N_29883);
nand UO_3314 (O_3314,N_29887,N_29853);
and UO_3315 (O_3315,N_29115,N_29112);
nor UO_3316 (O_3316,N_29646,N_29340);
and UO_3317 (O_3317,N_29362,N_29650);
nor UO_3318 (O_3318,N_29938,N_29134);
nand UO_3319 (O_3319,N_29515,N_29230);
xor UO_3320 (O_3320,N_29769,N_29248);
and UO_3321 (O_3321,N_29724,N_29886);
xor UO_3322 (O_3322,N_29137,N_29740);
or UO_3323 (O_3323,N_29732,N_29163);
nand UO_3324 (O_3324,N_29414,N_29997);
or UO_3325 (O_3325,N_29969,N_29028);
nand UO_3326 (O_3326,N_29528,N_29812);
xor UO_3327 (O_3327,N_29862,N_29438);
nor UO_3328 (O_3328,N_29889,N_29895);
or UO_3329 (O_3329,N_29505,N_29029);
or UO_3330 (O_3330,N_29535,N_29366);
xor UO_3331 (O_3331,N_29499,N_29681);
xnor UO_3332 (O_3332,N_29648,N_29743);
or UO_3333 (O_3333,N_29002,N_29197);
or UO_3334 (O_3334,N_29125,N_29017);
and UO_3335 (O_3335,N_29373,N_29215);
or UO_3336 (O_3336,N_29434,N_29119);
or UO_3337 (O_3337,N_29036,N_29419);
xnor UO_3338 (O_3338,N_29293,N_29657);
or UO_3339 (O_3339,N_29657,N_29974);
and UO_3340 (O_3340,N_29990,N_29725);
xor UO_3341 (O_3341,N_29355,N_29272);
xor UO_3342 (O_3342,N_29198,N_29259);
xor UO_3343 (O_3343,N_29517,N_29561);
and UO_3344 (O_3344,N_29337,N_29579);
and UO_3345 (O_3345,N_29845,N_29396);
nor UO_3346 (O_3346,N_29690,N_29789);
xor UO_3347 (O_3347,N_29167,N_29303);
nand UO_3348 (O_3348,N_29110,N_29009);
and UO_3349 (O_3349,N_29646,N_29405);
xor UO_3350 (O_3350,N_29816,N_29722);
xor UO_3351 (O_3351,N_29900,N_29533);
nand UO_3352 (O_3352,N_29302,N_29301);
or UO_3353 (O_3353,N_29421,N_29545);
and UO_3354 (O_3354,N_29583,N_29844);
or UO_3355 (O_3355,N_29914,N_29873);
or UO_3356 (O_3356,N_29312,N_29006);
xor UO_3357 (O_3357,N_29408,N_29008);
and UO_3358 (O_3358,N_29862,N_29067);
or UO_3359 (O_3359,N_29188,N_29870);
and UO_3360 (O_3360,N_29897,N_29288);
nor UO_3361 (O_3361,N_29863,N_29544);
xor UO_3362 (O_3362,N_29322,N_29053);
and UO_3363 (O_3363,N_29651,N_29272);
and UO_3364 (O_3364,N_29270,N_29763);
and UO_3365 (O_3365,N_29864,N_29028);
and UO_3366 (O_3366,N_29264,N_29811);
and UO_3367 (O_3367,N_29092,N_29452);
nor UO_3368 (O_3368,N_29111,N_29948);
or UO_3369 (O_3369,N_29830,N_29845);
or UO_3370 (O_3370,N_29864,N_29616);
and UO_3371 (O_3371,N_29494,N_29666);
nand UO_3372 (O_3372,N_29445,N_29029);
nor UO_3373 (O_3373,N_29700,N_29649);
xor UO_3374 (O_3374,N_29950,N_29392);
nor UO_3375 (O_3375,N_29195,N_29321);
nand UO_3376 (O_3376,N_29996,N_29168);
xnor UO_3377 (O_3377,N_29901,N_29926);
or UO_3378 (O_3378,N_29441,N_29411);
nand UO_3379 (O_3379,N_29858,N_29019);
or UO_3380 (O_3380,N_29450,N_29683);
xor UO_3381 (O_3381,N_29756,N_29343);
and UO_3382 (O_3382,N_29792,N_29423);
or UO_3383 (O_3383,N_29480,N_29487);
nand UO_3384 (O_3384,N_29223,N_29290);
nor UO_3385 (O_3385,N_29684,N_29005);
nor UO_3386 (O_3386,N_29679,N_29552);
nand UO_3387 (O_3387,N_29593,N_29212);
or UO_3388 (O_3388,N_29246,N_29307);
or UO_3389 (O_3389,N_29173,N_29539);
xor UO_3390 (O_3390,N_29403,N_29255);
nor UO_3391 (O_3391,N_29406,N_29009);
and UO_3392 (O_3392,N_29731,N_29372);
xnor UO_3393 (O_3393,N_29314,N_29608);
or UO_3394 (O_3394,N_29779,N_29240);
or UO_3395 (O_3395,N_29168,N_29907);
and UO_3396 (O_3396,N_29194,N_29768);
xnor UO_3397 (O_3397,N_29433,N_29398);
xor UO_3398 (O_3398,N_29914,N_29826);
and UO_3399 (O_3399,N_29534,N_29681);
xnor UO_3400 (O_3400,N_29417,N_29707);
nand UO_3401 (O_3401,N_29280,N_29255);
or UO_3402 (O_3402,N_29198,N_29669);
nor UO_3403 (O_3403,N_29026,N_29066);
nor UO_3404 (O_3404,N_29928,N_29854);
xor UO_3405 (O_3405,N_29962,N_29715);
nand UO_3406 (O_3406,N_29649,N_29845);
xor UO_3407 (O_3407,N_29271,N_29670);
and UO_3408 (O_3408,N_29614,N_29519);
nand UO_3409 (O_3409,N_29209,N_29183);
and UO_3410 (O_3410,N_29908,N_29351);
or UO_3411 (O_3411,N_29383,N_29983);
nand UO_3412 (O_3412,N_29281,N_29259);
nor UO_3413 (O_3413,N_29583,N_29193);
nor UO_3414 (O_3414,N_29082,N_29959);
or UO_3415 (O_3415,N_29919,N_29441);
nand UO_3416 (O_3416,N_29535,N_29401);
and UO_3417 (O_3417,N_29310,N_29568);
nor UO_3418 (O_3418,N_29183,N_29783);
or UO_3419 (O_3419,N_29512,N_29941);
and UO_3420 (O_3420,N_29973,N_29830);
nand UO_3421 (O_3421,N_29836,N_29654);
and UO_3422 (O_3422,N_29533,N_29117);
and UO_3423 (O_3423,N_29469,N_29771);
or UO_3424 (O_3424,N_29920,N_29273);
nand UO_3425 (O_3425,N_29310,N_29238);
nor UO_3426 (O_3426,N_29579,N_29119);
nor UO_3427 (O_3427,N_29749,N_29807);
and UO_3428 (O_3428,N_29491,N_29781);
nand UO_3429 (O_3429,N_29571,N_29020);
and UO_3430 (O_3430,N_29986,N_29334);
nand UO_3431 (O_3431,N_29650,N_29884);
nand UO_3432 (O_3432,N_29311,N_29293);
or UO_3433 (O_3433,N_29195,N_29227);
nand UO_3434 (O_3434,N_29374,N_29116);
nor UO_3435 (O_3435,N_29172,N_29379);
nor UO_3436 (O_3436,N_29636,N_29402);
xnor UO_3437 (O_3437,N_29093,N_29177);
or UO_3438 (O_3438,N_29512,N_29372);
nand UO_3439 (O_3439,N_29790,N_29478);
nand UO_3440 (O_3440,N_29452,N_29083);
nor UO_3441 (O_3441,N_29630,N_29988);
xnor UO_3442 (O_3442,N_29626,N_29914);
or UO_3443 (O_3443,N_29435,N_29358);
or UO_3444 (O_3444,N_29660,N_29160);
and UO_3445 (O_3445,N_29545,N_29118);
xor UO_3446 (O_3446,N_29392,N_29152);
or UO_3447 (O_3447,N_29271,N_29911);
nand UO_3448 (O_3448,N_29373,N_29641);
or UO_3449 (O_3449,N_29926,N_29921);
and UO_3450 (O_3450,N_29484,N_29808);
nand UO_3451 (O_3451,N_29679,N_29696);
nand UO_3452 (O_3452,N_29636,N_29876);
nor UO_3453 (O_3453,N_29310,N_29764);
and UO_3454 (O_3454,N_29905,N_29547);
nand UO_3455 (O_3455,N_29835,N_29052);
and UO_3456 (O_3456,N_29569,N_29929);
or UO_3457 (O_3457,N_29285,N_29221);
xnor UO_3458 (O_3458,N_29712,N_29793);
xnor UO_3459 (O_3459,N_29620,N_29514);
nor UO_3460 (O_3460,N_29044,N_29449);
or UO_3461 (O_3461,N_29485,N_29999);
nand UO_3462 (O_3462,N_29383,N_29583);
and UO_3463 (O_3463,N_29351,N_29263);
xor UO_3464 (O_3464,N_29143,N_29465);
xor UO_3465 (O_3465,N_29124,N_29633);
xor UO_3466 (O_3466,N_29327,N_29898);
nand UO_3467 (O_3467,N_29949,N_29449);
nor UO_3468 (O_3468,N_29473,N_29139);
or UO_3469 (O_3469,N_29363,N_29649);
or UO_3470 (O_3470,N_29389,N_29238);
nor UO_3471 (O_3471,N_29016,N_29019);
nor UO_3472 (O_3472,N_29088,N_29341);
nor UO_3473 (O_3473,N_29998,N_29464);
and UO_3474 (O_3474,N_29410,N_29298);
xnor UO_3475 (O_3475,N_29804,N_29651);
or UO_3476 (O_3476,N_29948,N_29046);
nor UO_3477 (O_3477,N_29108,N_29890);
nand UO_3478 (O_3478,N_29158,N_29928);
and UO_3479 (O_3479,N_29642,N_29294);
and UO_3480 (O_3480,N_29842,N_29416);
and UO_3481 (O_3481,N_29234,N_29508);
nor UO_3482 (O_3482,N_29167,N_29827);
and UO_3483 (O_3483,N_29940,N_29236);
nor UO_3484 (O_3484,N_29533,N_29473);
xor UO_3485 (O_3485,N_29602,N_29790);
nand UO_3486 (O_3486,N_29038,N_29454);
nand UO_3487 (O_3487,N_29620,N_29073);
nor UO_3488 (O_3488,N_29859,N_29024);
and UO_3489 (O_3489,N_29491,N_29188);
and UO_3490 (O_3490,N_29567,N_29626);
or UO_3491 (O_3491,N_29157,N_29982);
xor UO_3492 (O_3492,N_29558,N_29566);
nor UO_3493 (O_3493,N_29582,N_29972);
nor UO_3494 (O_3494,N_29970,N_29880);
nand UO_3495 (O_3495,N_29705,N_29159);
nor UO_3496 (O_3496,N_29445,N_29162);
nor UO_3497 (O_3497,N_29932,N_29540);
xnor UO_3498 (O_3498,N_29902,N_29028);
nor UO_3499 (O_3499,N_29536,N_29477);
endmodule