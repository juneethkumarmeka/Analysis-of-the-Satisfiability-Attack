module basic_1000_10000_1500_50_levels_2xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_907,In_802);
nor U1 (N_1,In_758,In_805);
or U2 (N_2,In_478,In_86);
nor U3 (N_3,In_161,In_354);
nand U4 (N_4,In_69,In_494);
or U5 (N_5,In_465,In_303);
nand U6 (N_6,In_729,In_233);
nor U7 (N_7,In_825,In_838);
nand U8 (N_8,In_366,In_435);
nand U9 (N_9,In_851,In_502);
or U10 (N_10,In_650,In_603);
nand U11 (N_11,In_318,In_510);
or U12 (N_12,In_865,In_448);
xnor U13 (N_13,In_596,In_163);
and U14 (N_14,In_364,In_826);
nor U15 (N_15,In_594,In_289);
or U16 (N_16,In_271,In_269);
nand U17 (N_17,In_212,In_706);
and U18 (N_18,In_716,In_126);
nand U19 (N_19,In_299,In_198);
nor U20 (N_20,In_844,In_800);
and U21 (N_21,In_97,In_636);
nor U22 (N_22,In_22,In_947);
and U23 (N_23,In_760,In_374);
nand U24 (N_24,In_846,In_95);
nand U25 (N_25,In_182,In_81);
and U26 (N_26,In_931,In_797);
or U27 (N_27,In_262,In_455);
nand U28 (N_28,In_246,In_668);
or U29 (N_29,In_382,In_499);
or U30 (N_30,In_576,In_14);
nand U31 (N_31,In_121,In_138);
or U32 (N_32,In_350,In_273);
and U33 (N_33,In_935,In_599);
nor U34 (N_34,In_98,In_39);
nor U35 (N_35,In_590,In_993);
or U36 (N_36,In_215,In_996);
nand U37 (N_37,In_443,In_445);
xnor U38 (N_38,In_660,In_131);
nor U39 (N_39,In_609,In_737);
nor U40 (N_40,In_971,In_595);
and U41 (N_41,In_724,In_120);
nor U42 (N_42,In_910,In_591);
and U43 (N_43,In_437,In_646);
nand U44 (N_44,In_224,In_125);
nor U45 (N_45,In_777,In_308);
nor U46 (N_46,In_249,In_190);
nor U47 (N_47,In_235,In_567);
and U48 (N_48,In_475,In_765);
or U49 (N_49,In_624,In_171);
or U50 (N_50,In_44,In_261);
nand U51 (N_51,In_294,In_889);
nor U52 (N_52,In_201,In_543);
and U53 (N_53,In_183,In_420);
nand U54 (N_54,In_887,In_283);
or U55 (N_55,In_962,In_714);
nor U56 (N_56,In_167,In_547);
nor U57 (N_57,In_157,In_997);
and U58 (N_58,In_701,In_979);
nor U59 (N_59,In_741,In_438);
and U60 (N_60,In_504,In_360);
nor U61 (N_61,In_762,In_440);
or U62 (N_62,In_598,In_527);
or U63 (N_63,In_221,In_373);
and U64 (N_64,In_690,In_693);
nor U65 (N_65,In_639,In_775);
or U66 (N_66,In_89,In_684);
and U67 (N_67,In_732,In_425);
nor U68 (N_68,In_414,In_343);
or U69 (N_69,In_835,In_384);
and U70 (N_70,In_827,In_123);
nor U71 (N_71,In_640,In_881);
nor U72 (N_72,In_327,In_164);
nand U73 (N_73,In_862,In_179);
or U74 (N_74,In_549,In_62);
nor U75 (N_75,In_76,In_472);
or U76 (N_76,In_24,In_357);
nand U77 (N_77,In_930,In_616);
nor U78 (N_78,In_509,In_730);
or U79 (N_79,In_305,In_788);
and U80 (N_80,In_534,In_927);
nand U81 (N_81,In_561,In_105);
nand U82 (N_82,In_874,In_434);
nand U83 (N_83,In_255,In_752);
or U84 (N_84,In_584,In_491);
and U85 (N_85,In_109,In_924);
nor U86 (N_86,In_687,In_340);
nand U87 (N_87,In_515,In_857);
nand U88 (N_88,In_217,In_13);
or U89 (N_89,In_77,In_520);
nor U90 (N_90,In_557,In_866);
nor U91 (N_91,In_29,In_270);
nor U92 (N_92,In_454,In_681);
nand U93 (N_93,In_321,In_498);
or U94 (N_94,In_275,In_310);
or U95 (N_95,In_667,In_771);
nor U96 (N_96,In_942,In_877);
nand U97 (N_97,In_136,In_0);
or U98 (N_98,In_586,In_755);
or U99 (N_99,In_150,In_407);
nand U100 (N_100,In_140,In_416);
nand U101 (N_101,In_585,In_670);
nand U102 (N_102,In_348,In_296);
nand U103 (N_103,In_113,In_694);
nor U104 (N_104,In_917,In_961);
and U105 (N_105,In_159,In_511);
nor U106 (N_106,In_422,In_958);
or U107 (N_107,In_885,In_411);
and U108 (N_108,In_849,In_756);
and U109 (N_109,In_144,In_837);
nand U110 (N_110,In_367,In_52);
or U111 (N_111,In_776,In_256);
nor U112 (N_112,In_923,In_814);
and U113 (N_113,In_808,In_82);
and U114 (N_114,In_908,In_879);
nor U115 (N_115,In_747,In_241);
xor U116 (N_116,In_540,In_54);
nand U117 (N_117,In_238,In_749);
or U118 (N_118,In_858,In_535);
xnor U119 (N_119,In_631,In_780);
nand U120 (N_120,In_368,In_3);
and U121 (N_121,In_751,In_733);
nand U122 (N_122,In_116,In_976);
nor U123 (N_123,In_477,In_371);
nand U124 (N_124,In_978,In_46);
and U125 (N_125,In_850,In_983);
nand U126 (N_126,In_365,In_564);
nand U127 (N_127,In_876,In_583);
nor U128 (N_128,In_331,In_968);
nor U129 (N_129,In_61,In_723);
and U130 (N_130,In_873,In_127);
nor U131 (N_131,In_7,In_896);
nor U132 (N_132,In_871,In_298);
nand U133 (N_133,In_252,In_801);
nor U134 (N_134,In_550,In_840);
nor U135 (N_135,In_482,In_655);
nor U136 (N_136,In_102,In_951);
nor U137 (N_137,In_339,In_115);
or U138 (N_138,In_767,In_146);
or U139 (N_139,In_73,In_117);
nor U140 (N_140,In_152,In_390);
or U141 (N_141,In_325,In_165);
and U142 (N_142,In_114,In_592);
and U143 (N_143,In_848,In_854);
and U144 (N_144,In_59,In_88);
nand U145 (N_145,In_490,In_828);
and U146 (N_146,In_948,In_139);
nand U147 (N_147,In_539,In_789);
nor U148 (N_148,In_259,In_194);
nor U149 (N_149,In_284,In_719);
nand U150 (N_150,In_991,In_56);
or U151 (N_151,In_292,In_408);
and U152 (N_152,In_530,In_174);
nand U153 (N_153,In_912,In_613);
nor U154 (N_154,In_891,In_973);
and U155 (N_155,In_143,In_597);
and U156 (N_156,In_155,In_832);
or U157 (N_157,In_572,In_565);
nand U158 (N_158,In_717,In_313);
and U159 (N_159,In_806,In_64);
nand U160 (N_160,In_169,In_607);
nand U161 (N_161,In_944,In_404);
or U162 (N_162,In_427,In_734);
and U163 (N_163,In_992,In_742);
or U164 (N_164,In_381,In_459);
xor U165 (N_165,In_421,In_600);
nor U166 (N_166,In_754,In_798);
nor U167 (N_167,In_41,In_769);
and U168 (N_168,In_329,In_265);
and U169 (N_169,In_492,In_35);
and U170 (N_170,In_675,In_847);
or U171 (N_171,In_919,In_671);
nand U172 (N_172,In_254,In_322);
or U173 (N_173,In_248,In_987);
nand U174 (N_174,In_503,In_111);
and U175 (N_175,In_937,In_526);
and U176 (N_176,In_225,In_615);
and U177 (N_177,In_78,In_47);
xnor U178 (N_178,In_23,In_359);
nand U179 (N_179,In_712,In_264);
nand U180 (N_180,In_18,In_2);
or U181 (N_181,In_185,In_48);
nand U182 (N_182,In_93,In_929);
nand U183 (N_183,In_816,In_34);
and U184 (N_184,In_410,In_575);
xnor U185 (N_185,In_822,In_451);
or U186 (N_186,In_207,In_861);
nand U187 (N_187,In_998,In_38);
nand U188 (N_188,In_622,In_932);
nor U189 (N_189,In_785,In_954);
or U190 (N_190,In_933,In_376);
and U191 (N_191,In_999,In_618);
and U192 (N_192,In_629,In_500);
or U193 (N_193,In_938,In_778);
nor U194 (N_194,In_845,In_279);
and U195 (N_195,In_20,In_909);
and U196 (N_196,In_952,In_178);
or U197 (N_197,In_955,In_884);
or U198 (N_198,In_630,In_635);
nand U199 (N_199,In_211,In_718);
nand U200 (N_200,In_532,N_157);
nor U201 (N_201,In_319,N_124);
and U202 (N_202,In_517,In_324);
and U203 (N_203,N_170,In_841);
nor U204 (N_204,In_405,In_725);
nor U205 (N_205,N_31,N_179);
nor U206 (N_206,N_111,In_393);
xnor U207 (N_207,N_25,In_197);
nor U208 (N_208,N_19,In_379);
nand U209 (N_209,In_202,In_260);
nor U210 (N_210,In_957,N_17);
or U211 (N_211,In_456,N_32);
and U212 (N_212,N_39,In_748);
nor U213 (N_213,In_479,In_824);
nor U214 (N_214,In_1,In_84);
nand U215 (N_215,N_104,In_960);
nor U216 (N_216,In_941,N_167);
and U217 (N_217,In_469,In_295);
or U218 (N_218,In_579,In_297);
or U219 (N_219,In_45,N_10);
nor U220 (N_220,In_715,In_461);
nand U221 (N_221,In_55,In_134);
and U222 (N_222,In_672,In_489);
nand U223 (N_223,In_634,In_272);
nand U224 (N_224,In_108,In_316);
nor U225 (N_225,In_188,In_524);
and U226 (N_226,In_419,In_247);
nand U227 (N_227,In_394,In_356);
nand U228 (N_228,N_97,N_171);
nand U229 (N_229,In_314,In_49);
xor U230 (N_230,In_175,N_60);
and U231 (N_231,In_153,In_276);
nand U232 (N_232,N_106,N_5);
and U233 (N_233,In_263,In_145);
nand U234 (N_234,In_107,In_554);
or U235 (N_235,In_523,In_112);
and U236 (N_236,In_464,In_430);
nor U237 (N_237,In_287,In_137);
nor U238 (N_238,In_74,In_428);
nor U239 (N_239,In_245,In_395);
and U240 (N_240,In_770,In_85);
or U241 (N_241,In_677,In_66);
nand U242 (N_242,N_168,In_58);
nor U243 (N_243,In_546,N_108);
nor U244 (N_244,In_555,N_128);
nand U245 (N_245,In_617,In_433);
nor U246 (N_246,In_282,In_656);
nand U247 (N_247,In_423,In_400);
or U248 (N_248,In_432,N_59);
and U249 (N_249,N_110,In_429);
nor U250 (N_250,In_463,In_323);
or U251 (N_251,In_811,In_817);
nand U252 (N_252,In_810,In_286);
and U253 (N_253,In_135,N_137);
and U254 (N_254,N_177,N_155);
or U255 (N_255,In_19,N_56);
or U256 (N_256,In_214,In_306);
nand U257 (N_257,N_152,In_649);
or U258 (N_258,In_32,N_35);
or U259 (N_259,In_658,In_644);
and U260 (N_260,N_29,N_142);
nand U261 (N_261,In_229,In_57);
nor U262 (N_262,In_385,In_704);
nor U263 (N_263,In_637,In_506);
or U264 (N_264,In_562,In_815);
nor U265 (N_265,In_665,In_903);
and U266 (N_266,N_112,In_856);
nand U267 (N_267,In_389,In_956);
nor U268 (N_268,In_409,In_790);
or U269 (N_269,In_199,N_85);
and U270 (N_270,N_145,N_12);
nor U271 (N_271,N_162,N_20);
and U272 (N_272,In_870,In_80);
nand U273 (N_273,N_61,In_606);
nand U274 (N_274,In_4,N_166);
or U275 (N_275,In_28,In_669);
nor U276 (N_276,In_466,In_882);
nor U277 (N_277,In_36,In_556);
nand U278 (N_278,In_787,In_449);
or U279 (N_279,In_542,N_30);
nor U280 (N_280,N_113,In_290);
and U281 (N_281,In_333,In_441);
or U282 (N_282,In_552,N_86);
nor U283 (N_283,N_185,In_731);
and U284 (N_284,N_175,N_140);
nand U285 (N_285,In_415,In_580);
and U286 (N_286,N_36,N_184);
or U287 (N_287,In_766,In_982);
and U288 (N_288,In_657,In_156);
xor U289 (N_289,In_945,N_91);
and U290 (N_290,In_15,In_70);
nand U291 (N_291,In_601,In_743);
or U292 (N_292,N_53,In_989);
nand U293 (N_293,In_231,In_959);
and U294 (N_294,In_819,In_237);
nor U295 (N_295,In_699,In_574);
nand U296 (N_296,N_52,In_501);
nor U297 (N_297,In_42,N_0);
and U298 (N_298,In_711,N_150);
or U299 (N_299,In_654,In_738);
nand U300 (N_300,In_351,N_173);
nand U301 (N_301,In_151,N_82);
and U302 (N_302,N_195,N_28);
nand U303 (N_303,In_759,N_44);
and U304 (N_304,In_83,In_162);
nor U305 (N_305,N_54,N_37);
or U306 (N_306,In_674,In_892);
or U307 (N_307,N_138,In_147);
or U308 (N_308,In_234,In_678);
and U309 (N_309,N_27,In_274);
nor U310 (N_310,In_403,In_521);
nor U311 (N_311,In_218,In_496);
or U312 (N_312,N_109,N_165);
and U313 (N_313,N_58,In_709);
and U314 (N_314,In_981,In_529);
nand U315 (N_315,In_133,In_370);
or U316 (N_316,N_43,In_739);
and U317 (N_317,In_589,N_172);
and U318 (N_318,In_872,In_372);
or U319 (N_319,N_55,N_123);
or U320 (N_320,In_488,N_26);
and U321 (N_321,In_533,N_63);
nand U322 (N_322,N_45,In_67);
and U323 (N_323,N_182,In_12);
or U324 (N_324,In_573,N_164);
nor U325 (N_325,In_605,In_280);
or U326 (N_326,In_210,In_544);
nor U327 (N_327,N_180,In_807);
and U328 (N_328,In_926,In_782);
and U329 (N_329,In_966,In_713);
nand U330 (N_330,In_803,N_158);
nand U331 (N_331,In_326,In_158);
nand U332 (N_332,In_344,N_181);
and U333 (N_333,In_764,In_925);
or U334 (N_334,In_336,In_842);
nand U335 (N_335,In_285,N_190);
nor U336 (N_336,N_2,In_642);
nor U337 (N_337,N_186,In_679);
or U338 (N_338,In_936,In_783);
nor U339 (N_339,In_17,In_883);
xnor U340 (N_340,N_197,In_588);
nand U341 (N_341,N_4,In_700);
and U342 (N_342,In_514,In_666);
nor U343 (N_343,In_10,In_195);
nor U344 (N_344,N_114,N_153);
nor U345 (N_345,In_895,N_89);
and U346 (N_346,In_898,N_105);
or U347 (N_347,In_820,N_116);
and U348 (N_348,In_795,In_369);
nand U349 (N_349,In_177,In_792);
xor U350 (N_350,N_194,N_193);
or U351 (N_351,N_198,In_239);
nor U352 (N_352,N_154,In_453);
and U353 (N_353,In_347,In_467);
nand U354 (N_354,In_31,In_988);
or U355 (N_355,N_8,In_781);
nand U356 (N_356,In_11,In_16);
or U357 (N_357,In_843,In_916);
xor U358 (N_358,In_99,In_906);
xor U359 (N_359,In_242,In_399);
nand U360 (N_360,N_131,In_307);
xor U361 (N_361,In_266,N_126);
or U362 (N_362,N_41,N_73);
nand U363 (N_363,In_722,In_869);
nor U364 (N_364,N_64,In_537);
xnor U365 (N_365,In_582,In_302);
nand U366 (N_366,In_812,In_516);
or U367 (N_367,In_831,N_47);
nand U368 (N_368,In_149,In_934);
or U369 (N_369,In_864,N_46);
nand U370 (N_370,In_375,In_627);
and U371 (N_371,In_648,In_558);
or U372 (N_372,N_199,In_581);
nor U373 (N_373,In_943,In_142);
and U374 (N_374,In_184,In_967);
and U375 (N_375,N_51,In_386);
and U376 (N_376,N_75,In_257);
or U377 (N_377,In_474,In_972);
xnor U378 (N_378,In_563,In_628);
nor U379 (N_379,In_708,In_226);
nand U380 (N_380,In_969,In_860);
or U381 (N_381,In_974,In_72);
nor U382 (N_382,In_745,In_774);
and U383 (N_383,In_335,N_62);
nand U384 (N_384,N_7,In_380);
nand U385 (N_385,In_383,N_48);
or U386 (N_386,N_121,In_702);
nand U387 (N_387,In_328,In_559);
and U388 (N_388,In_222,In_5);
and U389 (N_389,In_462,In_43);
nor U390 (N_390,In_446,In_949);
nor U391 (N_391,N_80,In_101);
and U392 (N_392,In_33,In_553);
and U393 (N_393,In_196,In_40);
or U394 (N_394,N_188,In_338);
and U395 (N_395,In_103,In_560);
and U396 (N_396,N_143,In_878);
and U397 (N_397,In_705,In_258);
nor U398 (N_398,In_320,In_975);
or U399 (N_399,In_661,In_625);
or U400 (N_400,N_33,In_431);
nor U401 (N_401,N_280,In_990);
nand U402 (N_402,N_397,In_977);
and U403 (N_403,In_25,N_327);
nand U404 (N_404,N_289,N_222);
xnor U405 (N_405,In_703,In_676);
or U406 (N_406,N_3,In_697);
or U407 (N_407,N_341,In_426);
or U408 (N_408,In_880,N_318);
xnor U409 (N_409,In_794,N_296);
nor U410 (N_410,In_578,In_913);
xor U411 (N_411,In_181,N_232);
and U412 (N_412,In_897,In_119);
or U413 (N_413,N_216,In_964);
or U414 (N_414,N_283,In_643);
nor U415 (N_415,In_939,N_276);
and U416 (N_416,In_888,N_14);
and U417 (N_417,In_688,In_900);
xnor U418 (N_418,In_91,N_24);
nor U419 (N_419,N_81,In_508);
and U420 (N_420,N_156,In_412);
or U421 (N_421,N_208,N_203);
or U422 (N_422,In_487,N_117);
or U423 (N_423,N_141,In_193);
or U424 (N_424,In_250,In_545);
nand U425 (N_425,In_902,In_346);
or U426 (N_426,In_154,N_343);
and U427 (N_427,In_953,In_483);
and U428 (N_428,N_187,N_220);
and U429 (N_429,In_965,In_548);
nor U430 (N_430,In_619,In_950);
or U431 (N_431,N_250,N_320);
and U432 (N_432,N_129,In_911);
nor U433 (N_433,N_253,N_68);
and U434 (N_434,N_16,In_986);
or U435 (N_435,In_519,N_391);
nor U436 (N_436,N_396,N_322);
or U437 (N_437,N_311,In_349);
nor U438 (N_438,N_50,N_78);
or U439 (N_439,In_779,N_281);
nand U440 (N_440,In_387,N_371);
nand U441 (N_441,In_92,In_632);
or U442 (N_442,N_313,N_238);
or U443 (N_443,In_401,In_614);
or U444 (N_444,N_102,In_392);
and U445 (N_445,N_144,N_65);
xor U446 (N_446,In_172,N_252);
and U447 (N_447,N_77,In_970);
and U448 (N_448,In_570,N_139);
nand U449 (N_449,In_623,In_875);
and U450 (N_450,N_288,N_210);
nor U451 (N_451,In_784,N_248);
nand U452 (N_452,In_406,N_72);
nand U453 (N_453,In_87,In_768);
nor U454 (N_454,N_254,N_386);
nor U455 (N_455,In_823,In_645);
nor U456 (N_456,N_42,N_96);
nor U457 (N_457,In_963,In_569);
nand U458 (N_458,In_304,N_382);
nand U459 (N_459,In_200,In_398);
or U460 (N_460,N_270,In_21);
or U461 (N_461,N_119,In_641);
nand U462 (N_462,N_130,In_791);
and U463 (N_463,N_265,N_242);
nand U464 (N_464,In_353,In_189);
or U465 (N_465,In_662,In_311);
or U466 (N_466,N_321,N_277);
or U467 (N_467,In_485,In_130);
nor U468 (N_468,N_209,N_135);
or U469 (N_469,N_107,In_587);
nor U470 (N_470,In_922,In_209);
or U471 (N_471,N_178,In_278);
nor U472 (N_472,In_638,In_852);
nor U473 (N_473,In_692,N_340);
nor U474 (N_474,N_390,N_367);
or U475 (N_475,N_151,N_346);
nand U476 (N_476,N_368,N_363);
and U477 (N_477,In_26,N_260);
or U478 (N_478,N_330,N_373);
and U479 (N_479,In_894,In_460);
and U480 (N_480,In_493,N_337);
or U481 (N_481,N_101,N_103);
nand U482 (N_482,N_268,In_621);
nand U483 (N_483,N_206,In_863);
nor U484 (N_484,In_205,N_11);
nor U485 (N_485,N_134,In_799);
nor U486 (N_486,In_740,In_480);
or U487 (N_487,N_348,In_689);
and U488 (N_488,N_161,N_307);
nand U489 (N_489,In_148,In_9);
nor U490 (N_490,In_682,In_836);
nand U491 (N_491,In_859,N_83);
or U492 (N_492,In_481,N_237);
and U493 (N_493,N_71,N_84);
or U494 (N_494,In_735,In_680);
nand U495 (N_495,In_786,In_352);
or U496 (N_496,N_353,N_217);
nor U497 (N_497,N_319,In_129);
and U498 (N_498,N_40,N_393);
or U499 (N_499,In_170,N_282);
and U500 (N_500,N_122,In_180);
or U501 (N_501,In_744,N_258);
and U502 (N_502,N_95,In_696);
nor U503 (N_503,N_302,N_100);
nor U504 (N_504,In_763,N_364);
and U505 (N_505,In_612,In_341);
and U506 (N_506,N_192,In_721);
and U507 (N_507,In_355,N_240);
nor U508 (N_508,In_663,N_356);
nor U509 (N_509,N_324,N_269);
xor U510 (N_510,N_74,In_63);
and U511 (N_511,In_447,N_176);
nor U512 (N_512,N_274,In_551);
nand U513 (N_513,In_30,In_94);
and U514 (N_514,In_757,In_602);
nor U515 (N_515,N_377,N_329);
and U516 (N_516,N_230,N_136);
nand U517 (N_517,In_928,N_132);
nand U518 (N_518,N_18,N_272);
xnor U519 (N_519,In_813,N_169);
nand U520 (N_520,In_834,In_685);
and U521 (N_521,In_51,N_127);
nor U522 (N_522,In_505,N_354);
nor U523 (N_523,In_27,In_173);
nand U524 (N_524,In_223,In_664);
or U525 (N_525,N_314,N_385);
nand U526 (N_526,In_362,In_8);
and U527 (N_527,In_686,In_868);
nor U528 (N_528,In_568,In_452);
and U529 (N_529,In_243,N_148);
or U530 (N_530,In_337,In_293);
nor U531 (N_531,N_372,N_304);
and U532 (N_532,N_94,N_9);
or U533 (N_533,In_402,In_904);
nand U534 (N_534,N_160,In_914);
or U535 (N_535,N_146,In_358);
nor U536 (N_536,N_338,N_159);
nand U537 (N_537,N_333,N_221);
nor U538 (N_538,N_388,N_369);
nand U539 (N_539,In_809,In_980);
nor U540 (N_540,N_214,N_202);
and U541 (N_541,N_264,N_133);
nor U542 (N_542,N_392,N_278);
nor U543 (N_543,In_439,In_315);
and U544 (N_544,In_436,N_125);
and U545 (N_545,In_710,In_268);
and U546 (N_546,In_291,In_905);
and U547 (N_547,In_213,N_300);
or U548 (N_548,In_334,In_330);
nand U549 (N_549,In_604,N_271);
or U550 (N_550,N_201,In_166);
or U551 (N_551,N_251,In_830);
and U552 (N_552,N_355,In_985);
and U553 (N_553,In_458,N_34);
nor U554 (N_554,In_720,In_470);
nor U555 (N_555,N_239,N_273);
nor U556 (N_556,In_450,In_71);
or U557 (N_557,In_727,In_128);
or U558 (N_558,N_213,In_946);
nor U559 (N_559,In_610,In_396);
nand U560 (N_560,In_995,In_361);
and U561 (N_561,N_266,N_183);
and U562 (N_562,In_829,In_444);
and U563 (N_563,In_388,In_818);
or U564 (N_564,N_394,N_21);
or U565 (N_565,In_471,N_339);
or U566 (N_566,In_994,In_940);
nor U567 (N_567,N_310,In_691);
or U568 (N_568,N_376,N_228);
nand U569 (N_569,N_92,In_317);
nand U570 (N_570,In_240,N_98);
nand U571 (N_571,N_211,In_75);
nand U572 (N_572,N_352,N_285);
nor U573 (N_573,N_244,N_303);
or U574 (N_574,In_921,N_205);
nand U575 (N_575,In_186,N_378);
nor U576 (N_576,In_6,N_374);
nor U577 (N_577,N_115,N_233);
or U578 (N_578,In_473,N_196);
nor U579 (N_579,In_611,N_66);
and U580 (N_580,In_659,In_442);
or U581 (N_581,In_484,N_347);
nand U582 (N_582,N_49,N_189);
or U583 (N_583,In_853,In_309);
or U584 (N_584,N_342,In_79);
nor U585 (N_585,In_68,In_65);
nand U586 (N_586,In_633,In_528);
xor U587 (N_587,In_251,N_370);
nand U588 (N_588,In_378,In_203);
nor U589 (N_589,N_236,N_224);
and U590 (N_590,N_357,N_286);
nand U591 (N_591,N_6,N_200);
or U592 (N_592,In_683,N_249);
and U593 (N_593,N_381,N_79);
nand U594 (N_594,In_391,In_124);
nand U595 (N_595,In_698,N_334);
or U596 (N_596,N_88,N_389);
nand U597 (N_597,In_867,N_290);
nor U598 (N_598,N_247,In_855);
and U599 (N_599,In_522,In_397);
and U600 (N_600,In_60,In_100);
and U601 (N_601,N_455,N_474);
and U602 (N_602,N_583,N_421);
nand U603 (N_603,N_463,N_577);
or U604 (N_604,In_53,N_588);
and U605 (N_605,N_241,N_325);
nor U606 (N_606,N_326,N_564);
or U607 (N_607,N_562,In_773);
and U608 (N_608,N_443,N_500);
nor U609 (N_609,N_596,In_486);
nand U610 (N_610,N_23,N_528);
and U611 (N_611,N_479,N_470);
nor U612 (N_612,In_750,N_543);
nor U613 (N_613,N_519,N_399);
or U614 (N_614,N_556,N_408);
and U615 (N_615,N_529,N_308);
xnor U616 (N_616,N_478,N_545);
nand U617 (N_617,N_416,N_438);
nand U618 (N_618,N_323,N_571);
xor U619 (N_619,N_526,N_306);
nand U620 (N_620,In_707,In_232);
or U621 (N_621,N_542,N_229);
nor U622 (N_622,N_493,N_505);
and U623 (N_623,N_552,N_418);
nand U624 (N_624,N_405,N_293);
nor U625 (N_625,In_106,In_566);
xor U626 (N_626,In_288,N_548);
nand U627 (N_627,N_350,In_695);
and U628 (N_628,In_50,In_236);
or U629 (N_629,N_301,N_263);
and U630 (N_630,N_406,N_459);
nor U631 (N_631,N_453,N_549);
or U632 (N_632,N_585,N_379);
nand U633 (N_633,N_279,N_380);
and U634 (N_634,In_512,N_533);
nor U635 (N_635,N_568,In_424);
or U636 (N_636,N_511,N_473);
nor U637 (N_637,N_447,In_413);
nor U638 (N_638,N_362,N_335);
or U639 (N_639,N_538,In_653);
nor U640 (N_640,N_422,N_420);
xor U641 (N_641,N_557,N_521);
nor U642 (N_642,N_365,N_572);
xnor U643 (N_643,N_57,N_581);
or U644 (N_644,N_331,In_332);
or U645 (N_645,N_457,N_336);
nand U646 (N_646,N_471,N_223);
or U647 (N_647,N_361,In_230);
nand U648 (N_648,In_168,N_553);
nand U649 (N_649,In_228,N_480);
nor U650 (N_650,N_524,N_219);
and U651 (N_651,N_87,N_584);
nor U652 (N_652,N_433,N_448);
or U653 (N_653,N_70,In_804);
nand U654 (N_654,N_498,N_435);
nor U655 (N_655,N_445,In_216);
nand U656 (N_656,N_535,N_358);
and U657 (N_657,N_560,N_427);
nand U658 (N_658,N_496,N_586);
nand U659 (N_659,In_513,N_467);
nor U660 (N_660,In_531,In_187);
or U661 (N_661,N_512,In_495);
nor U662 (N_662,N_149,N_458);
or U663 (N_663,N_404,N_551);
nor U664 (N_664,N_316,N_559);
nand U665 (N_665,N_409,N_256);
nand U666 (N_666,N_507,N_477);
nand U667 (N_667,N_578,N_487);
or U668 (N_668,N_503,N_423);
nand U669 (N_669,N_461,In_518);
nor U670 (N_670,N_434,N_554);
and U671 (N_671,N_573,In_984);
or U672 (N_672,N_536,N_429);
and U673 (N_673,N_525,N_317);
nand U674 (N_674,N_502,N_432);
xnor U675 (N_675,In_160,N_328);
nand U676 (N_676,N_527,N_570);
and U677 (N_677,N_1,N_481);
and U678 (N_678,N_591,N_451);
and U679 (N_679,N_212,N_403);
nor U680 (N_680,N_287,In_219);
or U681 (N_681,N_514,N_257);
and U682 (N_682,N_579,N_417);
nand U683 (N_683,N_69,N_563);
and U684 (N_684,N_345,In_342);
or U685 (N_685,In_220,N_309);
and U686 (N_686,In_300,N_469);
and U687 (N_687,In_736,N_598);
nand U688 (N_688,N_517,N_509);
nor U689 (N_689,N_450,In_37);
or U690 (N_690,N_499,N_539);
nor U691 (N_691,N_495,In_345);
or U692 (N_692,In_626,In_673);
and U693 (N_693,In_227,N_426);
or U694 (N_694,N_235,N_547);
nand U695 (N_695,In_110,In_577);
nor U696 (N_696,In_893,In_890);
nand U697 (N_697,N_490,N_226);
xor U698 (N_698,In_525,N_440);
and U699 (N_699,In_593,N_315);
and U700 (N_700,N_465,N_513);
or U701 (N_701,N_444,In_652);
nor U702 (N_702,N_531,In_301);
or U703 (N_703,In_915,In_538);
nand U704 (N_704,N_246,N_291);
nor U705 (N_705,In_839,N_218);
and U706 (N_706,N_413,N_439);
or U707 (N_707,N_147,N_489);
or U708 (N_708,N_387,N_411);
xnor U709 (N_709,N_15,N_437);
nand U710 (N_710,In_821,N_259);
nor U711 (N_711,N_580,N_599);
or U712 (N_712,N_592,In_476);
or U713 (N_713,N_234,N_541);
nor U714 (N_714,In_920,N_225);
nor U715 (N_715,In_104,In_281);
or U716 (N_716,N_501,In_541);
or U717 (N_717,N_456,N_401);
and U718 (N_718,In_753,N_402);
nor U719 (N_719,N_540,N_13);
or U720 (N_720,N_460,N_398);
or U721 (N_721,In_418,N_76);
nor U722 (N_722,N_595,N_464);
and U723 (N_723,In_96,N_174);
nand U724 (N_724,N_476,In_468);
nand U725 (N_725,In_726,N_530);
and U726 (N_726,In_728,N_332);
and U727 (N_727,N_561,N_412);
nand U728 (N_728,N_261,N_67);
nor U729 (N_729,N_589,In_267);
or U730 (N_730,N_497,N_99);
and U731 (N_731,In_746,N_407);
or U732 (N_732,N_410,In_497);
or U733 (N_733,N_452,N_400);
or U734 (N_734,N_305,N_243);
or U735 (N_735,N_506,N_298);
or U736 (N_736,In_206,In_651);
and U737 (N_737,In_647,N_510);
nand U738 (N_738,N_294,In_277);
nor U739 (N_739,N_295,N_582);
or U740 (N_740,N_482,In_192);
or U741 (N_741,N_284,In_886);
and U742 (N_742,N_516,N_449);
nand U743 (N_743,In_833,N_520);
nor U744 (N_744,N_515,In_761);
nand U745 (N_745,N_430,N_475);
or U746 (N_746,N_227,N_344);
nor U747 (N_747,N_587,N_163);
nor U748 (N_748,N_90,N_366);
nand U749 (N_749,In_90,N_436);
xor U750 (N_750,N_360,In_899);
nand U751 (N_751,N_255,N_566);
nor U752 (N_752,In_571,In_118);
nor U753 (N_753,N_215,N_590);
and U754 (N_754,N_550,N_574);
and U755 (N_755,N_245,N_446);
nand U756 (N_756,N_532,N_22);
xnor U757 (N_757,N_120,N_375);
nand U758 (N_758,N_292,N_569);
and U759 (N_759,N_204,N_38);
or U760 (N_760,In_253,N_593);
nand U761 (N_761,In_793,N_576);
or U762 (N_762,In_122,N_312);
or U763 (N_763,N_558,In_176);
nor U764 (N_764,In_312,N_424);
and U765 (N_765,N_468,N_508);
or U766 (N_766,N_472,In_208);
or U767 (N_767,N_518,N_567);
nand U768 (N_768,N_534,In_132);
and U769 (N_769,N_491,N_575);
nor U770 (N_770,In_918,In_901);
nand U771 (N_771,N_207,N_93);
nor U772 (N_772,N_262,In_620);
nor U773 (N_773,N_442,In_377);
nor U774 (N_774,In_608,N_395);
or U775 (N_775,N_414,N_419);
and U776 (N_776,N_466,N_546);
nor U777 (N_777,N_118,N_351);
nor U778 (N_778,N_415,In_191);
nand U779 (N_779,N_483,N_594);
nand U780 (N_780,N_462,N_523);
and U781 (N_781,N_555,N_349);
or U782 (N_782,In_507,In_363);
or U783 (N_783,N_383,N_565);
or U784 (N_784,N_485,N_299);
or U785 (N_785,N_297,In_417);
and U786 (N_786,In_204,N_431);
nand U787 (N_787,N_231,In_244);
and U788 (N_788,N_544,N_486);
and U789 (N_789,In_796,N_441);
nand U790 (N_790,N_191,N_504);
and U791 (N_791,N_597,N_537);
or U792 (N_792,N_494,In_772);
nor U793 (N_793,N_384,N_492);
or U794 (N_794,N_428,In_457);
nand U795 (N_795,In_141,N_275);
or U796 (N_796,In_536,N_522);
nand U797 (N_797,N_454,N_488);
nand U798 (N_798,N_484,N_425);
nand U799 (N_799,N_359,N_267);
nand U800 (N_800,N_731,N_630);
nand U801 (N_801,N_645,N_760);
nand U802 (N_802,N_653,N_764);
nand U803 (N_803,N_759,N_701);
or U804 (N_804,N_770,N_756);
or U805 (N_805,N_690,N_682);
and U806 (N_806,N_743,N_611);
or U807 (N_807,N_672,N_621);
and U808 (N_808,N_684,N_692);
nand U809 (N_809,N_703,N_732);
and U810 (N_810,N_625,N_602);
xor U811 (N_811,N_699,N_716);
or U812 (N_812,N_723,N_689);
and U813 (N_813,N_778,N_719);
nand U814 (N_814,N_691,N_776);
or U815 (N_815,N_705,N_658);
and U816 (N_816,N_730,N_761);
or U817 (N_817,N_706,N_679);
nor U818 (N_818,N_744,N_720);
nor U819 (N_819,N_644,N_704);
and U820 (N_820,N_628,N_792);
nand U821 (N_821,N_726,N_781);
nor U822 (N_822,N_702,N_608);
nand U823 (N_823,N_668,N_772);
nor U824 (N_824,N_638,N_717);
or U825 (N_825,N_721,N_662);
and U826 (N_826,N_788,N_623);
or U827 (N_827,N_746,N_605);
nand U828 (N_828,N_799,N_748);
nand U829 (N_829,N_675,N_707);
or U830 (N_830,N_750,N_652);
and U831 (N_831,N_661,N_613);
or U832 (N_832,N_734,N_656);
nor U833 (N_833,N_765,N_774);
nor U834 (N_834,N_678,N_620);
nor U835 (N_835,N_695,N_729);
nor U836 (N_836,N_694,N_629);
nand U837 (N_837,N_722,N_796);
nor U838 (N_838,N_791,N_631);
nand U839 (N_839,N_612,N_790);
and U840 (N_840,N_784,N_768);
and U841 (N_841,N_789,N_738);
nand U842 (N_842,N_670,N_604);
nand U843 (N_843,N_657,N_713);
and U844 (N_844,N_758,N_642);
nand U845 (N_845,N_632,N_600);
or U846 (N_846,N_766,N_673);
and U847 (N_847,N_777,N_637);
nand U848 (N_848,N_659,N_727);
and U849 (N_849,N_785,N_681);
or U850 (N_850,N_626,N_634);
nor U851 (N_851,N_618,N_718);
and U852 (N_852,N_633,N_769);
nand U853 (N_853,N_725,N_715);
xnor U854 (N_854,N_683,N_609);
or U855 (N_855,N_780,N_724);
nand U856 (N_856,N_763,N_709);
or U857 (N_857,N_677,N_794);
or U858 (N_858,N_798,N_601);
or U859 (N_859,N_669,N_749);
nor U860 (N_860,N_664,N_775);
nor U861 (N_861,N_753,N_708);
xnor U862 (N_862,N_617,N_619);
and U863 (N_863,N_773,N_736);
nand U864 (N_864,N_616,N_747);
or U865 (N_865,N_696,N_636);
nor U866 (N_866,N_742,N_735);
or U867 (N_867,N_714,N_643);
nand U868 (N_868,N_741,N_755);
nand U869 (N_869,N_737,N_676);
or U870 (N_870,N_651,N_680);
and U871 (N_871,N_710,N_740);
and U872 (N_872,N_693,N_687);
or U873 (N_873,N_635,N_795);
or U874 (N_874,N_771,N_603);
and U875 (N_875,N_666,N_697);
nor U876 (N_876,N_786,N_779);
nor U877 (N_877,N_674,N_671);
or U878 (N_878,N_751,N_712);
xor U879 (N_879,N_739,N_615);
or U880 (N_880,N_700,N_688);
or U881 (N_881,N_639,N_614);
nand U882 (N_882,N_647,N_787);
or U883 (N_883,N_650,N_667);
or U884 (N_884,N_757,N_646);
nand U885 (N_885,N_754,N_745);
nand U886 (N_886,N_665,N_698);
nor U887 (N_887,N_641,N_797);
and U888 (N_888,N_640,N_686);
or U889 (N_889,N_622,N_782);
or U890 (N_890,N_793,N_606);
or U891 (N_891,N_711,N_660);
nor U892 (N_892,N_627,N_655);
nor U893 (N_893,N_610,N_752);
or U894 (N_894,N_783,N_648);
or U895 (N_895,N_733,N_654);
and U896 (N_896,N_649,N_663);
nor U897 (N_897,N_767,N_607);
or U898 (N_898,N_624,N_762);
xor U899 (N_899,N_728,N_685);
nor U900 (N_900,N_692,N_719);
and U901 (N_901,N_710,N_687);
and U902 (N_902,N_723,N_709);
nand U903 (N_903,N_799,N_729);
or U904 (N_904,N_792,N_692);
nor U905 (N_905,N_646,N_703);
nand U906 (N_906,N_725,N_673);
or U907 (N_907,N_653,N_740);
or U908 (N_908,N_705,N_677);
or U909 (N_909,N_616,N_782);
or U910 (N_910,N_727,N_678);
or U911 (N_911,N_777,N_728);
nand U912 (N_912,N_686,N_601);
and U913 (N_913,N_661,N_673);
nand U914 (N_914,N_732,N_711);
or U915 (N_915,N_697,N_649);
or U916 (N_916,N_668,N_774);
nand U917 (N_917,N_688,N_790);
and U918 (N_918,N_795,N_629);
nand U919 (N_919,N_614,N_771);
nand U920 (N_920,N_767,N_641);
or U921 (N_921,N_737,N_772);
or U922 (N_922,N_634,N_769);
or U923 (N_923,N_612,N_632);
or U924 (N_924,N_708,N_707);
nor U925 (N_925,N_684,N_662);
and U926 (N_926,N_672,N_636);
and U927 (N_927,N_762,N_660);
nor U928 (N_928,N_644,N_616);
or U929 (N_929,N_602,N_706);
nand U930 (N_930,N_629,N_637);
nor U931 (N_931,N_770,N_701);
nor U932 (N_932,N_704,N_799);
nor U933 (N_933,N_719,N_600);
nor U934 (N_934,N_755,N_628);
nand U935 (N_935,N_658,N_788);
and U936 (N_936,N_780,N_715);
nor U937 (N_937,N_635,N_705);
xnor U938 (N_938,N_620,N_705);
nor U939 (N_939,N_658,N_671);
or U940 (N_940,N_772,N_686);
nor U941 (N_941,N_675,N_693);
or U942 (N_942,N_607,N_623);
or U943 (N_943,N_786,N_782);
or U944 (N_944,N_685,N_716);
nand U945 (N_945,N_716,N_791);
or U946 (N_946,N_767,N_652);
or U947 (N_947,N_646,N_714);
nor U948 (N_948,N_612,N_785);
or U949 (N_949,N_645,N_751);
xnor U950 (N_950,N_650,N_625);
or U951 (N_951,N_607,N_612);
nor U952 (N_952,N_621,N_684);
nand U953 (N_953,N_615,N_631);
and U954 (N_954,N_667,N_784);
nor U955 (N_955,N_792,N_752);
or U956 (N_956,N_679,N_747);
and U957 (N_957,N_721,N_799);
and U958 (N_958,N_796,N_757);
xor U959 (N_959,N_726,N_632);
nor U960 (N_960,N_606,N_652);
nor U961 (N_961,N_657,N_740);
or U962 (N_962,N_677,N_610);
xor U963 (N_963,N_628,N_659);
nand U964 (N_964,N_694,N_653);
and U965 (N_965,N_621,N_780);
or U966 (N_966,N_694,N_640);
and U967 (N_967,N_697,N_653);
or U968 (N_968,N_624,N_652);
or U969 (N_969,N_707,N_740);
nor U970 (N_970,N_707,N_774);
or U971 (N_971,N_638,N_739);
or U972 (N_972,N_610,N_663);
or U973 (N_973,N_795,N_690);
nand U974 (N_974,N_721,N_616);
and U975 (N_975,N_689,N_690);
or U976 (N_976,N_648,N_707);
or U977 (N_977,N_752,N_750);
or U978 (N_978,N_706,N_753);
nor U979 (N_979,N_613,N_666);
nor U980 (N_980,N_616,N_612);
nand U981 (N_981,N_776,N_766);
nor U982 (N_982,N_725,N_744);
xnor U983 (N_983,N_725,N_739);
and U984 (N_984,N_612,N_779);
nand U985 (N_985,N_603,N_785);
and U986 (N_986,N_767,N_645);
and U987 (N_987,N_720,N_763);
or U988 (N_988,N_689,N_699);
or U989 (N_989,N_654,N_683);
nand U990 (N_990,N_698,N_720);
and U991 (N_991,N_776,N_731);
nor U992 (N_992,N_783,N_748);
or U993 (N_993,N_606,N_798);
or U994 (N_994,N_641,N_677);
or U995 (N_995,N_756,N_685);
or U996 (N_996,N_670,N_774);
and U997 (N_997,N_722,N_734);
nand U998 (N_998,N_739,N_720);
and U999 (N_999,N_681,N_795);
nand U1000 (N_1000,N_931,N_939);
nand U1001 (N_1001,N_801,N_909);
and U1002 (N_1002,N_960,N_817);
and U1003 (N_1003,N_908,N_934);
xnor U1004 (N_1004,N_879,N_861);
and U1005 (N_1005,N_911,N_962);
xor U1006 (N_1006,N_930,N_901);
nor U1007 (N_1007,N_948,N_886);
and U1008 (N_1008,N_816,N_863);
nor U1009 (N_1009,N_874,N_980);
nand U1010 (N_1010,N_958,N_912);
nand U1011 (N_1011,N_964,N_828);
nand U1012 (N_1012,N_803,N_894);
nor U1013 (N_1013,N_916,N_904);
and U1014 (N_1014,N_830,N_970);
nor U1015 (N_1015,N_866,N_975);
nand U1016 (N_1016,N_932,N_870);
and U1017 (N_1017,N_915,N_895);
and U1018 (N_1018,N_835,N_988);
or U1019 (N_1019,N_867,N_890);
xor U1020 (N_1020,N_846,N_954);
or U1021 (N_1021,N_938,N_822);
and U1022 (N_1022,N_971,N_900);
or U1023 (N_1023,N_985,N_815);
nand U1024 (N_1024,N_812,N_955);
or U1025 (N_1025,N_831,N_840);
nor U1026 (N_1026,N_913,N_808);
nor U1027 (N_1027,N_972,N_860);
nand U1028 (N_1028,N_882,N_829);
nand U1029 (N_1029,N_850,N_877);
nor U1030 (N_1030,N_824,N_876);
nor U1031 (N_1031,N_887,N_992);
nand U1032 (N_1032,N_818,N_959);
or U1033 (N_1033,N_907,N_814);
nand U1034 (N_1034,N_947,N_827);
and U1035 (N_1035,N_924,N_961);
nor U1036 (N_1036,N_996,N_883);
nand U1037 (N_1037,N_837,N_906);
nand U1038 (N_1038,N_905,N_889);
or U1039 (N_1039,N_898,N_806);
and U1040 (N_1040,N_997,N_914);
and U1041 (N_1041,N_859,N_892);
or U1042 (N_1042,N_966,N_884);
nand U1043 (N_1043,N_945,N_953);
xor U1044 (N_1044,N_833,N_853);
nand U1045 (N_1045,N_977,N_813);
nand U1046 (N_1046,N_893,N_897);
nor U1047 (N_1047,N_919,N_839);
nor U1048 (N_1048,N_848,N_881);
or U1049 (N_1049,N_922,N_844);
or U1050 (N_1050,N_841,N_946);
xor U1051 (N_1051,N_805,N_986);
xor U1052 (N_1052,N_868,N_902);
or U1053 (N_1053,N_956,N_856);
nor U1054 (N_1054,N_855,N_927);
or U1055 (N_1055,N_836,N_918);
or U1056 (N_1056,N_878,N_888);
and U1057 (N_1057,N_845,N_978);
nor U1058 (N_1058,N_957,N_858);
or U1059 (N_1059,N_826,N_823);
xor U1060 (N_1060,N_821,N_951);
and U1061 (N_1061,N_969,N_802);
nand U1062 (N_1062,N_872,N_920);
nand U1063 (N_1063,N_973,N_923);
nor U1064 (N_1064,N_869,N_994);
nand U1065 (N_1065,N_963,N_937);
and U1066 (N_1066,N_989,N_933);
nor U1067 (N_1067,N_979,N_832);
or U1068 (N_1068,N_849,N_885);
and U1069 (N_1069,N_917,N_896);
nand U1070 (N_1070,N_981,N_999);
and U1071 (N_1071,N_854,N_929);
and U1072 (N_1072,N_800,N_950);
nor U1073 (N_1073,N_838,N_809);
nor U1074 (N_1074,N_880,N_976);
or U1075 (N_1075,N_847,N_873);
or U1076 (N_1076,N_910,N_965);
or U1077 (N_1077,N_834,N_998);
xnor U1078 (N_1078,N_899,N_967);
nand U1079 (N_1079,N_949,N_983);
nor U1080 (N_1080,N_843,N_943);
nand U1081 (N_1081,N_857,N_807);
and U1082 (N_1082,N_811,N_921);
and U1083 (N_1083,N_942,N_941);
nor U1084 (N_1084,N_820,N_974);
and U1085 (N_1085,N_862,N_852);
or U1086 (N_1086,N_891,N_925);
or U1087 (N_1087,N_935,N_984);
nor U1088 (N_1088,N_991,N_944);
and U1089 (N_1089,N_940,N_952);
xnor U1090 (N_1090,N_865,N_851);
nor U1091 (N_1091,N_987,N_995);
or U1092 (N_1092,N_871,N_864);
and U1093 (N_1093,N_993,N_968);
or U1094 (N_1094,N_903,N_875);
or U1095 (N_1095,N_819,N_842);
nand U1096 (N_1096,N_825,N_928);
and U1097 (N_1097,N_810,N_982);
and U1098 (N_1098,N_926,N_936);
nand U1099 (N_1099,N_804,N_990);
and U1100 (N_1100,N_921,N_806);
nor U1101 (N_1101,N_879,N_880);
nand U1102 (N_1102,N_877,N_842);
nor U1103 (N_1103,N_872,N_902);
and U1104 (N_1104,N_898,N_993);
nand U1105 (N_1105,N_853,N_898);
nand U1106 (N_1106,N_904,N_985);
nor U1107 (N_1107,N_943,N_862);
nor U1108 (N_1108,N_932,N_886);
and U1109 (N_1109,N_811,N_994);
or U1110 (N_1110,N_976,N_809);
nor U1111 (N_1111,N_947,N_882);
nand U1112 (N_1112,N_991,N_863);
or U1113 (N_1113,N_913,N_987);
or U1114 (N_1114,N_973,N_959);
or U1115 (N_1115,N_805,N_879);
nand U1116 (N_1116,N_842,N_861);
nand U1117 (N_1117,N_878,N_913);
or U1118 (N_1118,N_917,N_909);
nor U1119 (N_1119,N_937,N_841);
nor U1120 (N_1120,N_908,N_887);
or U1121 (N_1121,N_897,N_815);
nor U1122 (N_1122,N_944,N_885);
or U1123 (N_1123,N_889,N_808);
nand U1124 (N_1124,N_884,N_816);
nand U1125 (N_1125,N_898,N_929);
nor U1126 (N_1126,N_923,N_885);
or U1127 (N_1127,N_980,N_811);
nand U1128 (N_1128,N_875,N_842);
nand U1129 (N_1129,N_936,N_935);
or U1130 (N_1130,N_959,N_827);
or U1131 (N_1131,N_935,N_843);
and U1132 (N_1132,N_920,N_878);
or U1133 (N_1133,N_894,N_843);
and U1134 (N_1134,N_924,N_838);
and U1135 (N_1135,N_974,N_940);
and U1136 (N_1136,N_816,N_910);
and U1137 (N_1137,N_908,N_811);
nor U1138 (N_1138,N_822,N_878);
or U1139 (N_1139,N_815,N_942);
nand U1140 (N_1140,N_854,N_997);
and U1141 (N_1141,N_924,N_856);
and U1142 (N_1142,N_848,N_851);
xor U1143 (N_1143,N_861,N_807);
nand U1144 (N_1144,N_840,N_811);
and U1145 (N_1145,N_806,N_875);
nand U1146 (N_1146,N_812,N_928);
and U1147 (N_1147,N_901,N_820);
and U1148 (N_1148,N_930,N_828);
nand U1149 (N_1149,N_930,N_830);
nor U1150 (N_1150,N_809,N_981);
or U1151 (N_1151,N_825,N_915);
or U1152 (N_1152,N_826,N_945);
nand U1153 (N_1153,N_887,N_897);
and U1154 (N_1154,N_970,N_974);
and U1155 (N_1155,N_840,N_817);
nor U1156 (N_1156,N_963,N_919);
or U1157 (N_1157,N_835,N_865);
nor U1158 (N_1158,N_995,N_950);
and U1159 (N_1159,N_868,N_925);
and U1160 (N_1160,N_964,N_850);
and U1161 (N_1161,N_990,N_808);
xor U1162 (N_1162,N_944,N_851);
nor U1163 (N_1163,N_871,N_886);
nand U1164 (N_1164,N_981,N_879);
and U1165 (N_1165,N_981,N_867);
nor U1166 (N_1166,N_874,N_867);
and U1167 (N_1167,N_977,N_860);
nor U1168 (N_1168,N_800,N_986);
nand U1169 (N_1169,N_834,N_802);
nor U1170 (N_1170,N_862,N_827);
nor U1171 (N_1171,N_934,N_823);
nand U1172 (N_1172,N_830,N_824);
nand U1173 (N_1173,N_900,N_965);
or U1174 (N_1174,N_914,N_900);
nand U1175 (N_1175,N_809,N_916);
xor U1176 (N_1176,N_800,N_867);
and U1177 (N_1177,N_942,N_805);
or U1178 (N_1178,N_907,N_887);
nand U1179 (N_1179,N_866,N_956);
nand U1180 (N_1180,N_806,N_873);
or U1181 (N_1181,N_973,N_819);
nor U1182 (N_1182,N_952,N_873);
or U1183 (N_1183,N_808,N_985);
nor U1184 (N_1184,N_969,N_961);
nand U1185 (N_1185,N_933,N_896);
or U1186 (N_1186,N_939,N_942);
nor U1187 (N_1187,N_887,N_929);
xnor U1188 (N_1188,N_901,N_828);
or U1189 (N_1189,N_904,N_890);
nand U1190 (N_1190,N_812,N_885);
nor U1191 (N_1191,N_902,N_815);
or U1192 (N_1192,N_929,N_885);
and U1193 (N_1193,N_927,N_897);
nand U1194 (N_1194,N_871,N_988);
nand U1195 (N_1195,N_867,N_960);
nor U1196 (N_1196,N_914,N_824);
or U1197 (N_1197,N_839,N_972);
or U1198 (N_1198,N_962,N_855);
nor U1199 (N_1199,N_978,N_914);
or U1200 (N_1200,N_1132,N_1199);
and U1201 (N_1201,N_1119,N_1181);
and U1202 (N_1202,N_1035,N_1068);
nor U1203 (N_1203,N_1173,N_1071);
nand U1204 (N_1204,N_1041,N_1110);
and U1205 (N_1205,N_1124,N_1040);
or U1206 (N_1206,N_1046,N_1197);
and U1207 (N_1207,N_1175,N_1114);
and U1208 (N_1208,N_1145,N_1017);
nand U1209 (N_1209,N_1096,N_1147);
nand U1210 (N_1210,N_1195,N_1077);
nand U1211 (N_1211,N_1164,N_1006);
and U1212 (N_1212,N_1090,N_1062);
and U1213 (N_1213,N_1083,N_1030);
and U1214 (N_1214,N_1036,N_1196);
nand U1215 (N_1215,N_1022,N_1031);
nand U1216 (N_1216,N_1058,N_1134);
or U1217 (N_1217,N_1162,N_1142);
nand U1218 (N_1218,N_1156,N_1008);
and U1219 (N_1219,N_1144,N_1101);
and U1220 (N_1220,N_1176,N_1100);
nor U1221 (N_1221,N_1168,N_1191);
or U1222 (N_1222,N_1067,N_1021);
or U1223 (N_1223,N_1174,N_1037);
nor U1224 (N_1224,N_1117,N_1053);
nand U1225 (N_1225,N_1169,N_1120);
nor U1226 (N_1226,N_1158,N_1188);
xnor U1227 (N_1227,N_1042,N_1066);
nor U1228 (N_1228,N_1087,N_1039);
nor U1229 (N_1229,N_1085,N_1179);
nor U1230 (N_1230,N_1009,N_1118);
and U1231 (N_1231,N_1126,N_1018);
nand U1232 (N_1232,N_1076,N_1154);
nand U1233 (N_1233,N_1127,N_1026);
and U1234 (N_1234,N_1038,N_1102);
or U1235 (N_1235,N_1024,N_1082);
or U1236 (N_1236,N_1084,N_1138);
and U1237 (N_1237,N_1032,N_1052);
or U1238 (N_1238,N_1109,N_1178);
nor U1239 (N_1239,N_1048,N_1170);
and U1240 (N_1240,N_1113,N_1152);
and U1241 (N_1241,N_1094,N_1148);
nor U1242 (N_1242,N_1140,N_1146);
nor U1243 (N_1243,N_1060,N_1001);
or U1244 (N_1244,N_1157,N_1141);
or U1245 (N_1245,N_1064,N_1044);
or U1246 (N_1246,N_1054,N_1091);
nor U1247 (N_1247,N_1194,N_1081);
nand U1248 (N_1248,N_1128,N_1005);
and U1249 (N_1249,N_1165,N_1003);
and U1250 (N_1250,N_1004,N_1092);
and U1251 (N_1251,N_1099,N_1079);
or U1252 (N_1252,N_1065,N_1088);
or U1253 (N_1253,N_1028,N_1027);
and U1254 (N_1254,N_1080,N_1093);
or U1255 (N_1255,N_1043,N_1183);
nor U1256 (N_1256,N_1089,N_1015);
or U1257 (N_1257,N_1122,N_1045);
nor U1258 (N_1258,N_1104,N_1150);
nand U1259 (N_1259,N_1025,N_1057);
and U1260 (N_1260,N_1070,N_1002);
nand U1261 (N_1261,N_1185,N_1155);
xor U1262 (N_1262,N_1073,N_1131);
or U1263 (N_1263,N_1153,N_1184);
and U1264 (N_1264,N_1166,N_1029);
nor U1265 (N_1265,N_1047,N_1159);
or U1266 (N_1266,N_1034,N_1049);
and U1267 (N_1267,N_1167,N_1171);
nor U1268 (N_1268,N_1149,N_1056);
xor U1269 (N_1269,N_1106,N_1095);
nand U1270 (N_1270,N_1069,N_1180);
nor U1271 (N_1271,N_1123,N_1163);
and U1272 (N_1272,N_1086,N_1010);
xor U1273 (N_1273,N_1193,N_1097);
nor U1274 (N_1274,N_1019,N_1139);
nand U1275 (N_1275,N_1137,N_1023);
nor U1276 (N_1276,N_1161,N_1011);
nor U1277 (N_1277,N_1186,N_1177);
nand U1278 (N_1278,N_1121,N_1190);
nand U1279 (N_1279,N_1074,N_1007);
or U1280 (N_1280,N_1103,N_1059);
nand U1281 (N_1281,N_1133,N_1198);
nand U1282 (N_1282,N_1151,N_1108);
nand U1283 (N_1283,N_1160,N_1116);
nand U1284 (N_1284,N_1135,N_1072);
or U1285 (N_1285,N_1172,N_1136);
or U1286 (N_1286,N_1061,N_1078);
and U1287 (N_1287,N_1192,N_1143);
nand U1288 (N_1288,N_1055,N_1098);
nor U1289 (N_1289,N_1051,N_1129);
or U1290 (N_1290,N_1063,N_1130);
nor U1291 (N_1291,N_1020,N_1107);
and U1292 (N_1292,N_1187,N_1033);
xor U1293 (N_1293,N_1182,N_1115);
and U1294 (N_1294,N_1050,N_1075);
and U1295 (N_1295,N_1189,N_1000);
or U1296 (N_1296,N_1112,N_1014);
or U1297 (N_1297,N_1013,N_1016);
nor U1298 (N_1298,N_1111,N_1105);
nand U1299 (N_1299,N_1012,N_1125);
and U1300 (N_1300,N_1000,N_1130);
nand U1301 (N_1301,N_1139,N_1065);
and U1302 (N_1302,N_1128,N_1074);
or U1303 (N_1303,N_1029,N_1162);
or U1304 (N_1304,N_1155,N_1000);
nand U1305 (N_1305,N_1049,N_1127);
or U1306 (N_1306,N_1031,N_1057);
and U1307 (N_1307,N_1005,N_1013);
nand U1308 (N_1308,N_1006,N_1071);
or U1309 (N_1309,N_1137,N_1165);
nand U1310 (N_1310,N_1126,N_1150);
nor U1311 (N_1311,N_1159,N_1008);
nand U1312 (N_1312,N_1058,N_1155);
nor U1313 (N_1313,N_1050,N_1060);
and U1314 (N_1314,N_1162,N_1161);
or U1315 (N_1315,N_1127,N_1033);
or U1316 (N_1316,N_1049,N_1010);
or U1317 (N_1317,N_1044,N_1114);
and U1318 (N_1318,N_1009,N_1142);
and U1319 (N_1319,N_1107,N_1141);
nand U1320 (N_1320,N_1140,N_1147);
and U1321 (N_1321,N_1096,N_1098);
nand U1322 (N_1322,N_1196,N_1035);
or U1323 (N_1323,N_1158,N_1041);
nand U1324 (N_1324,N_1119,N_1183);
nor U1325 (N_1325,N_1102,N_1031);
and U1326 (N_1326,N_1171,N_1189);
or U1327 (N_1327,N_1181,N_1017);
nand U1328 (N_1328,N_1137,N_1155);
nor U1329 (N_1329,N_1121,N_1169);
nor U1330 (N_1330,N_1089,N_1009);
nand U1331 (N_1331,N_1088,N_1054);
nand U1332 (N_1332,N_1119,N_1156);
nand U1333 (N_1333,N_1120,N_1192);
nor U1334 (N_1334,N_1178,N_1017);
and U1335 (N_1335,N_1101,N_1127);
nor U1336 (N_1336,N_1146,N_1197);
or U1337 (N_1337,N_1077,N_1030);
and U1338 (N_1338,N_1068,N_1144);
or U1339 (N_1339,N_1064,N_1069);
and U1340 (N_1340,N_1134,N_1047);
nand U1341 (N_1341,N_1102,N_1071);
nand U1342 (N_1342,N_1084,N_1071);
and U1343 (N_1343,N_1136,N_1119);
or U1344 (N_1344,N_1049,N_1135);
nor U1345 (N_1345,N_1194,N_1108);
nor U1346 (N_1346,N_1169,N_1006);
or U1347 (N_1347,N_1156,N_1116);
nor U1348 (N_1348,N_1162,N_1056);
and U1349 (N_1349,N_1141,N_1023);
nor U1350 (N_1350,N_1177,N_1075);
nor U1351 (N_1351,N_1110,N_1034);
nor U1352 (N_1352,N_1194,N_1096);
nor U1353 (N_1353,N_1175,N_1014);
or U1354 (N_1354,N_1167,N_1155);
or U1355 (N_1355,N_1193,N_1181);
nand U1356 (N_1356,N_1112,N_1085);
or U1357 (N_1357,N_1021,N_1139);
or U1358 (N_1358,N_1020,N_1134);
nand U1359 (N_1359,N_1104,N_1078);
and U1360 (N_1360,N_1035,N_1161);
nand U1361 (N_1361,N_1146,N_1158);
or U1362 (N_1362,N_1079,N_1131);
nor U1363 (N_1363,N_1091,N_1075);
or U1364 (N_1364,N_1016,N_1039);
nand U1365 (N_1365,N_1177,N_1184);
and U1366 (N_1366,N_1128,N_1052);
and U1367 (N_1367,N_1083,N_1179);
and U1368 (N_1368,N_1040,N_1008);
nand U1369 (N_1369,N_1040,N_1002);
nand U1370 (N_1370,N_1189,N_1145);
nor U1371 (N_1371,N_1090,N_1051);
nor U1372 (N_1372,N_1120,N_1196);
or U1373 (N_1373,N_1067,N_1095);
and U1374 (N_1374,N_1199,N_1091);
or U1375 (N_1375,N_1192,N_1151);
nand U1376 (N_1376,N_1174,N_1048);
nor U1377 (N_1377,N_1018,N_1069);
nand U1378 (N_1378,N_1047,N_1014);
or U1379 (N_1379,N_1097,N_1185);
nor U1380 (N_1380,N_1091,N_1111);
and U1381 (N_1381,N_1156,N_1004);
nand U1382 (N_1382,N_1122,N_1172);
nor U1383 (N_1383,N_1067,N_1153);
and U1384 (N_1384,N_1176,N_1104);
or U1385 (N_1385,N_1068,N_1055);
nor U1386 (N_1386,N_1016,N_1083);
and U1387 (N_1387,N_1080,N_1187);
or U1388 (N_1388,N_1149,N_1032);
nor U1389 (N_1389,N_1054,N_1192);
or U1390 (N_1390,N_1061,N_1188);
nor U1391 (N_1391,N_1060,N_1071);
nand U1392 (N_1392,N_1126,N_1017);
or U1393 (N_1393,N_1134,N_1103);
nand U1394 (N_1394,N_1150,N_1106);
or U1395 (N_1395,N_1081,N_1098);
or U1396 (N_1396,N_1048,N_1146);
nor U1397 (N_1397,N_1165,N_1107);
nand U1398 (N_1398,N_1002,N_1063);
and U1399 (N_1399,N_1106,N_1062);
and U1400 (N_1400,N_1206,N_1243);
and U1401 (N_1401,N_1351,N_1246);
nor U1402 (N_1402,N_1380,N_1263);
nor U1403 (N_1403,N_1288,N_1283);
or U1404 (N_1404,N_1238,N_1370);
nand U1405 (N_1405,N_1212,N_1249);
nor U1406 (N_1406,N_1265,N_1259);
or U1407 (N_1407,N_1269,N_1231);
nand U1408 (N_1408,N_1376,N_1359);
nand U1409 (N_1409,N_1285,N_1322);
nor U1410 (N_1410,N_1366,N_1346);
or U1411 (N_1411,N_1270,N_1253);
nand U1412 (N_1412,N_1377,N_1382);
and U1413 (N_1413,N_1205,N_1345);
xor U1414 (N_1414,N_1298,N_1349);
and U1415 (N_1415,N_1267,N_1297);
nand U1416 (N_1416,N_1391,N_1342);
or U1417 (N_1417,N_1241,N_1354);
and U1418 (N_1418,N_1328,N_1291);
nor U1419 (N_1419,N_1200,N_1373);
nand U1420 (N_1420,N_1242,N_1282);
and U1421 (N_1421,N_1316,N_1209);
and U1422 (N_1422,N_1289,N_1287);
or U1423 (N_1423,N_1293,N_1394);
nor U1424 (N_1424,N_1224,N_1386);
nor U1425 (N_1425,N_1341,N_1215);
and U1426 (N_1426,N_1303,N_1308);
nor U1427 (N_1427,N_1397,N_1385);
nand U1428 (N_1428,N_1256,N_1367);
nand U1429 (N_1429,N_1294,N_1389);
nor U1430 (N_1430,N_1378,N_1362);
nor U1431 (N_1431,N_1277,N_1324);
nor U1432 (N_1432,N_1239,N_1290);
or U1433 (N_1433,N_1326,N_1276);
nand U1434 (N_1434,N_1353,N_1286);
nand U1435 (N_1435,N_1396,N_1315);
or U1436 (N_1436,N_1240,N_1201);
and U1437 (N_1437,N_1363,N_1333);
and U1438 (N_1438,N_1344,N_1255);
nand U1439 (N_1439,N_1340,N_1251);
nand U1440 (N_1440,N_1300,N_1372);
and U1441 (N_1441,N_1321,N_1379);
nor U1442 (N_1442,N_1233,N_1331);
nor U1443 (N_1443,N_1273,N_1247);
nand U1444 (N_1444,N_1325,N_1252);
nand U1445 (N_1445,N_1334,N_1335);
nor U1446 (N_1446,N_1218,N_1284);
and U1447 (N_1447,N_1371,N_1260);
nand U1448 (N_1448,N_1207,N_1272);
nor U1449 (N_1449,N_1220,N_1262);
or U1450 (N_1450,N_1358,N_1398);
and U1451 (N_1451,N_1343,N_1234);
and U1452 (N_1452,N_1395,N_1271);
or U1453 (N_1453,N_1365,N_1202);
and U1454 (N_1454,N_1214,N_1318);
and U1455 (N_1455,N_1313,N_1274);
and U1456 (N_1456,N_1387,N_1330);
nor U1457 (N_1457,N_1227,N_1307);
nand U1458 (N_1458,N_1299,N_1381);
nand U1459 (N_1459,N_1230,N_1314);
nor U1460 (N_1460,N_1383,N_1257);
nand U1461 (N_1461,N_1232,N_1369);
xor U1462 (N_1462,N_1319,N_1302);
nor U1463 (N_1463,N_1245,N_1350);
and U1464 (N_1464,N_1355,N_1361);
nand U1465 (N_1465,N_1248,N_1235);
nand U1466 (N_1466,N_1301,N_1266);
and U1467 (N_1467,N_1312,N_1305);
nand U1468 (N_1468,N_1304,N_1210);
nand U1469 (N_1469,N_1275,N_1368);
nor U1470 (N_1470,N_1356,N_1250);
nand U1471 (N_1471,N_1216,N_1211);
nand U1472 (N_1472,N_1237,N_1204);
nand U1473 (N_1473,N_1279,N_1261);
and U1474 (N_1474,N_1311,N_1352);
or U1475 (N_1475,N_1332,N_1208);
nand U1476 (N_1476,N_1236,N_1222);
and U1477 (N_1477,N_1296,N_1228);
or U1478 (N_1478,N_1219,N_1392);
and U1479 (N_1479,N_1384,N_1339);
nor U1480 (N_1480,N_1244,N_1306);
and U1481 (N_1481,N_1278,N_1292);
and U1482 (N_1482,N_1374,N_1217);
nor U1483 (N_1483,N_1360,N_1348);
and U1484 (N_1484,N_1254,N_1309);
or U1485 (N_1485,N_1390,N_1375);
or U1486 (N_1486,N_1388,N_1310);
nand U1487 (N_1487,N_1364,N_1338);
or U1488 (N_1488,N_1295,N_1327);
nand U1489 (N_1489,N_1223,N_1347);
and U1490 (N_1490,N_1320,N_1213);
nand U1491 (N_1491,N_1203,N_1317);
or U1492 (N_1492,N_1393,N_1268);
nor U1493 (N_1493,N_1280,N_1399);
or U1494 (N_1494,N_1258,N_1229);
nor U1495 (N_1495,N_1225,N_1336);
and U1496 (N_1496,N_1329,N_1221);
nand U1497 (N_1497,N_1281,N_1337);
nand U1498 (N_1498,N_1323,N_1226);
and U1499 (N_1499,N_1264,N_1357);
and U1500 (N_1500,N_1202,N_1390);
nand U1501 (N_1501,N_1226,N_1256);
and U1502 (N_1502,N_1357,N_1284);
nand U1503 (N_1503,N_1263,N_1244);
or U1504 (N_1504,N_1321,N_1242);
nor U1505 (N_1505,N_1368,N_1292);
or U1506 (N_1506,N_1314,N_1377);
nor U1507 (N_1507,N_1246,N_1251);
and U1508 (N_1508,N_1296,N_1274);
nand U1509 (N_1509,N_1339,N_1286);
and U1510 (N_1510,N_1399,N_1384);
nor U1511 (N_1511,N_1265,N_1329);
nor U1512 (N_1512,N_1283,N_1329);
nand U1513 (N_1513,N_1339,N_1360);
nor U1514 (N_1514,N_1231,N_1298);
and U1515 (N_1515,N_1226,N_1287);
xnor U1516 (N_1516,N_1279,N_1372);
and U1517 (N_1517,N_1387,N_1213);
and U1518 (N_1518,N_1294,N_1368);
or U1519 (N_1519,N_1310,N_1206);
and U1520 (N_1520,N_1289,N_1371);
nor U1521 (N_1521,N_1370,N_1240);
nand U1522 (N_1522,N_1283,N_1313);
or U1523 (N_1523,N_1364,N_1217);
or U1524 (N_1524,N_1394,N_1253);
and U1525 (N_1525,N_1222,N_1364);
nand U1526 (N_1526,N_1281,N_1377);
or U1527 (N_1527,N_1295,N_1340);
nor U1528 (N_1528,N_1288,N_1356);
nand U1529 (N_1529,N_1327,N_1233);
and U1530 (N_1530,N_1276,N_1368);
or U1531 (N_1531,N_1380,N_1336);
nand U1532 (N_1532,N_1202,N_1376);
and U1533 (N_1533,N_1370,N_1226);
nand U1534 (N_1534,N_1286,N_1372);
or U1535 (N_1535,N_1307,N_1303);
or U1536 (N_1536,N_1326,N_1333);
and U1537 (N_1537,N_1318,N_1387);
or U1538 (N_1538,N_1244,N_1272);
and U1539 (N_1539,N_1396,N_1250);
xnor U1540 (N_1540,N_1205,N_1258);
or U1541 (N_1541,N_1332,N_1399);
nand U1542 (N_1542,N_1298,N_1218);
nor U1543 (N_1543,N_1327,N_1363);
nand U1544 (N_1544,N_1304,N_1372);
and U1545 (N_1545,N_1262,N_1205);
nor U1546 (N_1546,N_1387,N_1223);
nand U1547 (N_1547,N_1369,N_1376);
and U1548 (N_1548,N_1266,N_1279);
nor U1549 (N_1549,N_1250,N_1317);
or U1550 (N_1550,N_1300,N_1226);
xor U1551 (N_1551,N_1293,N_1278);
and U1552 (N_1552,N_1345,N_1287);
and U1553 (N_1553,N_1304,N_1281);
and U1554 (N_1554,N_1335,N_1372);
and U1555 (N_1555,N_1268,N_1352);
or U1556 (N_1556,N_1365,N_1262);
nor U1557 (N_1557,N_1373,N_1202);
xnor U1558 (N_1558,N_1335,N_1293);
nand U1559 (N_1559,N_1218,N_1335);
or U1560 (N_1560,N_1304,N_1287);
nor U1561 (N_1561,N_1253,N_1299);
and U1562 (N_1562,N_1361,N_1335);
or U1563 (N_1563,N_1363,N_1240);
nand U1564 (N_1564,N_1236,N_1381);
and U1565 (N_1565,N_1372,N_1203);
and U1566 (N_1566,N_1346,N_1363);
nor U1567 (N_1567,N_1327,N_1365);
nand U1568 (N_1568,N_1283,N_1334);
nand U1569 (N_1569,N_1344,N_1372);
nand U1570 (N_1570,N_1362,N_1296);
nand U1571 (N_1571,N_1397,N_1256);
nand U1572 (N_1572,N_1225,N_1244);
or U1573 (N_1573,N_1304,N_1264);
and U1574 (N_1574,N_1270,N_1339);
nor U1575 (N_1575,N_1282,N_1211);
nand U1576 (N_1576,N_1220,N_1203);
nor U1577 (N_1577,N_1392,N_1339);
nand U1578 (N_1578,N_1368,N_1204);
nor U1579 (N_1579,N_1222,N_1243);
nor U1580 (N_1580,N_1222,N_1256);
and U1581 (N_1581,N_1390,N_1328);
or U1582 (N_1582,N_1315,N_1371);
xor U1583 (N_1583,N_1302,N_1225);
nor U1584 (N_1584,N_1287,N_1268);
or U1585 (N_1585,N_1349,N_1267);
and U1586 (N_1586,N_1287,N_1312);
nand U1587 (N_1587,N_1315,N_1232);
and U1588 (N_1588,N_1284,N_1372);
nand U1589 (N_1589,N_1367,N_1376);
or U1590 (N_1590,N_1373,N_1353);
nor U1591 (N_1591,N_1283,N_1272);
or U1592 (N_1592,N_1334,N_1256);
xor U1593 (N_1593,N_1282,N_1334);
nand U1594 (N_1594,N_1229,N_1334);
nor U1595 (N_1595,N_1293,N_1262);
and U1596 (N_1596,N_1362,N_1359);
nor U1597 (N_1597,N_1274,N_1247);
or U1598 (N_1598,N_1394,N_1306);
nor U1599 (N_1599,N_1270,N_1279);
or U1600 (N_1600,N_1484,N_1461);
or U1601 (N_1601,N_1569,N_1564);
nor U1602 (N_1602,N_1485,N_1503);
and U1603 (N_1603,N_1550,N_1472);
xnor U1604 (N_1604,N_1568,N_1437);
and U1605 (N_1605,N_1508,N_1496);
or U1606 (N_1606,N_1506,N_1478);
nor U1607 (N_1607,N_1452,N_1521);
nand U1608 (N_1608,N_1583,N_1440);
and U1609 (N_1609,N_1571,N_1557);
and U1610 (N_1610,N_1431,N_1597);
or U1611 (N_1611,N_1523,N_1507);
nand U1612 (N_1612,N_1559,N_1519);
nor U1613 (N_1613,N_1544,N_1509);
or U1614 (N_1614,N_1490,N_1426);
or U1615 (N_1615,N_1466,N_1546);
or U1616 (N_1616,N_1560,N_1486);
and U1617 (N_1617,N_1448,N_1551);
and U1618 (N_1618,N_1579,N_1463);
and U1619 (N_1619,N_1558,N_1539);
and U1620 (N_1620,N_1574,N_1567);
nand U1621 (N_1621,N_1411,N_1445);
or U1622 (N_1622,N_1512,N_1465);
xor U1623 (N_1623,N_1402,N_1554);
and U1624 (N_1624,N_1493,N_1407);
and U1625 (N_1625,N_1421,N_1598);
or U1626 (N_1626,N_1410,N_1581);
and U1627 (N_1627,N_1499,N_1572);
nand U1628 (N_1628,N_1500,N_1533);
and U1629 (N_1629,N_1427,N_1538);
or U1630 (N_1630,N_1430,N_1475);
nand U1631 (N_1631,N_1451,N_1436);
nand U1632 (N_1632,N_1545,N_1473);
nand U1633 (N_1633,N_1514,N_1488);
nor U1634 (N_1634,N_1495,N_1428);
nand U1635 (N_1635,N_1497,N_1522);
and U1636 (N_1636,N_1491,N_1513);
nand U1637 (N_1637,N_1565,N_1458);
nor U1638 (N_1638,N_1480,N_1439);
or U1639 (N_1639,N_1462,N_1595);
and U1640 (N_1640,N_1470,N_1457);
or U1641 (N_1641,N_1556,N_1453);
and U1642 (N_1642,N_1404,N_1599);
or U1643 (N_1643,N_1578,N_1501);
nor U1644 (N_1644,N_1580,N_1494);
nor U1645 (N_1645,N_1449,N_1415);
nand U1646 (N_1646,N_1518,N_1406);
and U1647 (N_1647,N_1530,N_1528);
nor U1648 (N_1648,N_1416,N_1590);
and U1649 (N_1649,N_1563,N_1433);
and U1650 (N_1650,N_1438,N_1540);
and U1651 (N_1651,N_1477,N_1573);
nor U1652 (N_1652,N_1403,N_1467);
and U1653 (N_1653,N_1587,N_1584);
nand U1654 (N_1654,N_1535,N_1515);
or U1655 (N_1655,N_1537,N_1593);
or U1656 (N_1656,N_1586,N_1562);
nor U1657 (N_1657,N_1460,N_1450);
and U1658 (N_1658,N_1520,N_1549);
and U1659 (N_1659,N_1511,N_1504);
or U1660 (N_1660,N_1469,N_1553);
or U1661 (N_1661,N_1543,N_1570);
nor U1662 (N_1662,N_1585,N_1502);
nand U1663 (N_1663,N_1487,N_1425);
nor U1664 (N_1664,N_1405,N_1541);
nor U1665 (N_1665,N_1412,N_1561);
nand U1666 (N_1666,N_1435,N_1596);
nor U1667 (N_1667,N_1527,N_1498);
nor U1668 (N_1668,N_1447,N_1505);
and U1669 (N_1669,N_1417,N_1479);
and U1670 (N_1670,N_1422,N_1526);
nand U1671 (N_1671,N_1443,N_1552);
xor U1672 (N_1672,N_1456,N_1401);
nor U1673 (N_1673,N_1582,N_1492);
and U1674 (N_1674,N_1413,N_1408);
nor U1675 (N_1675,N_1483,N_1534);
nand U1676 (N_1676,N_1420,N_1481);
or U1677 (N_1677,N_1548,N_1517);
nor U1678 (N_1678,N_1442,N_1446);
nor U1679 (N_1679,N_1566,N_1444);
or U1680 (N_1680,N_1532,N_1575);
and U1681 (N_1681,N_1529,N_1542);
or U1682 (N_1682,N_1576,N_1577);
and U1683 (N_1683,N_1424,N_1400);
and U1684 (N_1684,N_1464,N_1423);
nand U1685 (N_1685,N_1516,N_1531);
nand U1686 (N_1686,N_1591,N_1454);
nor U1687 (N_1687,N_1489,N_1588);
or U1688 (N_1688,N_1592,N_1547);
and U1689 (N_1689,N_1555,N_1429);
nand U1690 (N_1690,N_1474,N_1471);
and U1691 (N_1691,N_1409,N_1468);
nand U1692 (N_1692,N_1476,N_1418);
nand U1693 (N_1693,N_1589,N_1510);
and U1694 (N_1694,N_1536,N_1419);
and U1695 (N_1695,N_1459,N_1455);
or U1696 (N_1696,N_1524,N_1525);
or U1697 (N_1697,N_1594,N_1441);
or U1698 (N_1698,N_1414,N_1434);
xnor U1699 (N_1699,N_1482,N_1432);
nor U1700 (N_1700,N_1451,N_1570);
nor U1701 (N_1701,N_1594,N_1513);
or U1702 (N_1702,N_1416,N_1514);
and U1703 (N_1703,N_1450,N_1523);
nor U1704 (N_1704,N_1407,N_1520);
nor U1705 (N_1705,N_1499,N_1413);
nand U1706 (N_1706,N_1446,N_1576);
nand U1707 (N_1707,N_1571,N_1475);
or U1708 (N_1708,N_1561,N_1588);
nor U1709 (N_1709,N_1485,N_1457);
or U1710 (N_1710,N_1513,N_1591);
and U1711 (N_1711,N_1518,N_1524);
nand U1712 (N_1712,N_1574,N_1469);
and U1713 (N_1713,N_1449,N_1430);
nor U1714 (N_1714,N_1517,N_1525);
or U1715 (N_1715,N_1540,N_1459);
nand U1716 (N_1716,N_1538,N_1542);
nor U1717 (N_1717,N_1483,N_1463);
and U1718 (N_1718,N_1569,N_1406);
and U1719 (N_1719,N_1568,N_1510);
nor U1720 (N_1720,N_1446,N_1415);
nor U1721 (N_1721,N_1511,N_1576);
and U1722 (N_1722,N_1453,N_1542);
and U1723 (N_1723,N_1509,N_1421);
or U1724 (N_1724,N_1504,N_1552);
nor U1725 (N_1725,N_1540,N_1532);
nor U1726 (N_1726,N_1457,N_1420);
nand U1727 (N_1727,N_1545,N_1457);
xnor U1728 (N_1728,N_1495,N_1543);
and U1729 (N_1729,N_1577,N_1471);
and U1730 (N_1730,N_1400,N_1442);
nand U1731 (N_1731,N_1439,N_1536);
or U1732 (N_1732,N_1467,N_1504);
and U1733 (N_1733,N_1440,N_1574);
or U1734 (N_1734,N_1420,N_1514);
nand U1735 (N_1735,N_1434,N_1442);
nand U1736 (N_1736,N_1421,N_1420);
nor U1737 (N_1737,N_1424,N_1533);
and U1738 (N_1738,N_1573,N_1419);
xor U1739 (N_1739,N_1508,N_1521);
or U1740 (N_1740,N_1416,N_1404);
or U1741 (N_1741,N_1553,N_1466);
or U1742 (N_1742,N_1563,N_1579);
and U1743 (N_1743,N_1403,N_1469);
and U1744 (N_1744,N_1578,N_1403);
nand U1745 (N_1745,N_1417,N_1553);
and U1746 (N_1746,N_1485,N_1410);
nor U1747 (N_1747,N_1542,N_1420);
nand U1748 (N_1748,N_1527,N_1467);
nor U1749 (N_1749,N_1591,N_1424);
or U1750 (N_1750,N_1453,N_1522);
or U1751 (N_1751,N_1424,N_1407);
or U1752 (N_1752,N_1410,N_1453);
nand U1753 (N_1753,N_1538,N_1458);
nand U1754 (N_1754,N_1533,N_1468);
nor U1755 (N_1755,N_1544,N_1527);
or U1756 (N_1756,N_1527,N_1564);
or U1757 (N_1757,N_1541,N_1473);
nor U1758 (N_1758,N_1564,N_1500);
or U1759 (N_1759,N_1515,N_1504);
and U1760 (N_1760,N_1466,N_1452);
and U1761 (N_1761,N_1433,N_1518);
xor U1762 (N_1762,N_1434,N_1483);
or U1763 (N_1763,N_1402,N_1501);
and U1764 (N_1764,N_1521,N_1496);
or U1765 (N_1765,N_1407,N_1567);
or U1766 (N_1766,N_1423,N_1597);
nand U1767 (N_1767,N_1474,N_1580);
or U1768 (N_1768,N_1518,N_1467);
or U1769 (N_1769,N_1510,N_1449);
and U1770 (N_1770,N_1406,N_1471);
or U1771 (N_1771,N_1518,N_1498);
nor U1772 (N_1772,N_1584,N_1573);
and U1773 (N_1773,N_1474,N_1490);
and U1774 (N_1774,N_1452,N_1577);
nand U1775 (N_1775,N_1471,N_1429);
or U1776 (N_1776,N_1430,N_1431);
and U1777 (N_1777,N_1431,N_1407);
and U1778 (N_1778,N_1417,N_1438);
nand U1779 (N_1779,N_1430,N_1486);
and U1780 (N_1780,N_1453,N_1408);
or U1781 (N_1781,N_1553,N_1460);
nand U1782 (N_1782,N_1559,N_1534);
nand U1783 (N_1783,N_1509,N_1405);
and U1784 (N_1784,N_1401,N_1443);
and U1785 (N_1785,N_1491,N_1559);
nand U1786 (N_1786,N_1421,N_1476);
or U1787 (N_1787,N_1469,N_1472);
and U1788 (N_1788,N_1462,N_1478);
nor U1789 (N_1789,N_1477,N_1519);
nand U1790 (N_1790,N_1440,N_1491);
xor U1791 (N_1791,N_1492,N_1507);
or U1792 (N_1792,N_1578,N_1416);
and U1793 (N_1793,N_1580,N_1505);
nand U1794 (N_1794,N_1519,N_1571);
or U1795 (N_1795,N_1489,N_1595);
or U1796 (N_1796,N_1427,N_1480);
or U1797 (N_1797,N_1446,N_1406);
or U1798 (N_1798,N_1540,N_1468);
and U1799 (N_1799,N_1450,N_1543);
and U1800 (N_1800,N_1641,N_1745);
nor U1801 (N_1801,N_1717,N_1651);
nor U1802 (N_1802,N_1665,N_1724);
nand U1803 (N_1803,N_1607,N_1635);
or U1804 (N_1804,N_1663,N_1684);
or U1805 (N_1805,N_1688,N_1661);
nor U1806 (N_1806,N_1751,N_1644);
or U1807 (N_1807,N_1730,N_1741);
nor U1808 (N_1808,N_1615,N_1772);
and U1809 (N_1809,N_1675,N_1773);
and U1810 (N_1810,N_1746,N_1791);
nor U1811 (N_1811,N_1617,N_1756);
or U1812 (N_1812,N_1642,N_1696);
xor U1813 (N_1813,N_1723,N_1796);
nand U1814 (N_1814,N_1689,N_1779);
nand U1815 (N_1815,N_1762,N_1695);
and U1816 (N_1816,N_1792,N_1613);
nand U1817 (N_1817,N_1782,N_1609);
nand U1818 (N_1818,N_1759,N_1740);
or U1819 (N_1819,N_1768,N_1707);
nand U1820 (N_1820,N_1781,N_1783);
nand U1821 (N_1821,N_1650,N_1660);
and U1822 (N_1822,N_1602,N_1739);
xnor U1823 (N_1823,N_1713,N_1700);
or U1824 (N_1824,N_1763,N_1706);
and U1825 (N_1825,N_1799,N_1657);
nor U1826 (N_1826,N_1787,N_1712);
or U1827 (N_1827,N_1727,N_1780);
and U1828 (N_1828,N_1682,N_1735);
nand U1829 (N_1829,N_1620,N_1680);
and U1830 (N_1830,N_1624,N_1679);
nor U1831 (N_1831,N_1685,N_1738);
nand U1832 (N_1832,N_1691,N_1729);
and U1833 (N_1833,N_1765,N_1640);
nand U1834 (N_1834,N_1770,N_1670);
and U1835 (N_1835,N_1631,N_1619);
and U1836 (N_1836,N_1639,N_1633);
and U1837 (N_1837,N_1702,N_1721);
or U1838 (N_1838,N_1618,N_1622);
or U1839 (N_1839,N_1666,N_1761);
and U1840 (N_1840,N_1715,N_1720);
and U1841 (N_1841,N_1752,N_1734);
nor U1842 (N_1842,N_1697,N_1671);
nor U1843 (N_1843,N_1760,N_1748);
or U1844 (N_1844,N_1608,N_1626);
nor U1845 (N_1845,N_1636,N_1648);
nor U1846 (N_1846,N_1652,N_1672);
or U1847 (N_1847,N_1647,N_1699);
nor U1848 (N_1848,N_1774,N_1743);
or U1849 (N_1849,N_1793,N_1726);
nor U1850 (N_1850,N_1764,N_1654);
nor U1851 (N_1851,N_1630,N_1794);
nor U1852 (N_1852,N_1758,N_1676);
or U1853 (N_1853,N_1718,N_1690);
or U1854 (N_1854,N_1668,N_1643);
nor U1855 (N_1855,N_1605,N_1634);
or U1856 (N_1856,N_1673,N_1653);
nand U1857 (N_1857,N_1662,N_1692);
nor U1858 (N_1858,N_1693,N_1686);
nor U1859 (N_1859,N_1674,N_1766);
nand U1860 (N_1860,N_1646,N_1737);
and U1861 (N_1861,N_1681,N_1784);
xnor U1862 (N_1862,N_1710,N_1701);
and U1863 (N_1863,N_1600,N_1664);
nor U1864 (N_1864,N_1606,N_1777);
nand U1865 (N_1865,N_1629,N_1722);
or U1866 (N_1866,N_1612,N_1638);
nor U1867 (N_1867,N_1709,N_1789);
and U1868 (N_1868,N_1601,N_1797);
or U1869 (N_1869,N_1669,N_1790);
and U1870 (N_1870,N_1610,N_1747);
nand U1871 (N_1871,N_1623,N_1733);
nor U1872 (N_1872,N_1616,N_1604);
and U1873 (N_1873,N_1656,N_1716);
and U1874 (N_1874,N_1798,N_1754);
and U1875 (N_1875,N_1621,N_1785);
nand U1876 (N_1876,N_1769,N_1775);
nand U1877 (N_1877,N_1753,N_1719);
or U1878 (N_1878,N_1725,N_1704);
and U1879 (N_1879,N_1732,N_1757);
nand U1880 (N_1880,N_1683,N_1698);
or U1881 (N_1881,N_1708,N_1655);
nand U1882 (N_1882,N_1728,N_1755);
nand U1883 (N_1883,N_1736,N_1677);
nor U1884 (N_1884,N_1678,N_1637);
nor U1885 (N_1885,N_1611,N_1667);
or U1886 (N_1886,N_1778,N_1711);
nand U1887 (N_1887,N_1750,N_1749);
nand U1888 (N_1888,N_1628,N_1786);
nand U1889 (N_1889,N_1742,N_1632);
nand U1890 (N_1890,N_1659,N_1703);
nand U1891 (N_1891,N_1687,N_1771);
or U1892 (N_1892,N_1714,N_1658);
or U1893 (N_1893,N_1645,N_1795);
nor U1894 (N_1894,N_1603,N_1788);
and U1895 (N_1895,N_1649,N_1694);
or U1896 (N_1896,N_1731,N_1744);
nand U1897 (N_1897,N_1614,N_1776);
nand U1898 (N_1898,N_1767,N_1705);
nand U1899 (N_1899,N_1625,N_1627);
nand U1900 (N_1900,N_1720,N_1671);
nor U1901 (N_1901,N_1602,N_1638);
nor U1902 (N_1902,N_1767,N_1661);
nand U1903 (N_1903,N_1624,N_1771);
or U1904 (N_1904,N_1641,N_1695);
and U1905 (N_1905,N_1720,N_1708);
and U1906 (N_1906,N_1625,N_1650);
and U1907 (N_1907,N_1709,N_1612);
or U1908 (N_1908,N_1713,N_1613);
nand U1909 (N_1909,N_1681,N_1686);
nor U1910 (N_1910,N_1691,N_1721);
and U1911 (N_1911,N_1744,N_1793);
and U1912 (N_1912,N_1664,N_1709);
nor U1913 (N_1913,N_1734,N_1647);
nor U1914 (N_1914,N_1670,N_1724);
and U1915 (N_1915,N_1776,N_1644);
nand U1916 (N_1916,N_1746,N_1687);
or U1917 (N_1917,N_1604,N_1637);
and U1918 (N_1918,N_1672,N_1774);
and U1919 (N_1919,N_1600,N_1642);
nor U1920 (N_1920,N_1642,N_1605);
or U1921 (N_1921,N_1686,N_1776);
xor U1922 (N_1922,N_1746,N_1758);
and U1923 (N_1923,N_1755,N_1799);
nor U1924 (N_1924,N_1708,N_1715);
and U1925 (N_1925,N_1623,N_1795);
or U1926 (N_1926,N_1629,N_1655);
and U1927 (N_1927,N_1766,N_1743);
nand U1928 (N_1928,N_1779,N_1694);
nor U1929 (N_1929,N_1758,N_1781);
or U1930 (N_1930,N_1616,N_1621);
nand U1931 (N_1931,N_1777,N_1717);
and U1932 (N_1932,N_1688,N_1674);
nor U1933 (N_1933,N_1676,N_1738);
or U1934 (N_1934,N_1743,N_1642);
nor U1935 (N_1935,N_1744,N_1754);
nor U1936 (N_1936,N_1663,N_1614);
or U1937 (N_1937,N_1606,N_1735);
or U1938 (N_1938,N_1641,N_1699);
nand U1939 (N_1939,N_1738,N_1722);
or U1940 (N_1940,N_1700,N_1777);
or U1941 (N_1941,N_1651,N_1634);
or U1942 (N_1942,N_1710,N_1646);
or U1943 (N_1943,N_1766,N_1718);
or U1944 (N_1944,N_1653,N_1717);
or U1945 (N_1945,N_1789,N_1624);
nor U1946 (N_1946,N_1699,N_1632);
or U1947 (N_1947,N_1763,N_1643);
and U1948 (N_1948,N_1762,N_1753);
nor U1949 (N_1949,N_1721,N_1728);
and U1950 (N_1950,N_1702,N_1776);
nor U1951 (N_1951,N_1645,N_1730);
nor U1952 (N_1952,N_1629,N_1745);
nand U1953 (N_1953,N_1724,N_1662);
and U1954 (N_1954,N_1666,N_1613);
nand U1955 (N_1955,N_1680,N_1797);
nor U1956 (N_1956,N_1765,N_1768);
nand U1957 (N_1957,N_1793,N_1607);
and U1958 (N_1958,N_1752,N_1758);
and U1959 (N_1959,N_1773,N_1688);
and U1960 (N_1960,N_1763,N_1665);
nand U1961 (N_1961,N_1780,N_1697);
and U1962 (N_1962,N_1740,N_1672);
nand U1963 (N_1963,N_1730,N_1770);
nand U1964 (N_1964,N_1699,N_1673);
and U1965 (N_1965,N_1678,N_1797);
and U1966 (N_1966,N_1681,N_1776);
and U1967 (N_1967,N_1755,N_1678);
nand U1968 (N_1968,N_1712,N_1614);
or U1969 (N_1969,N_1650,N_1747);
and U1970 (N_1970,N_1789,N_1700);
nor U1971 (N_1971,N_1652,N_1671);
and U1972 (N_1972,N_1664,N_1776);
nor U1973 (N_1973,N_1617,N_1740);
or U1974 (N_1974,N_1667,N_1602);
nor U1975 (N_1975,N_1794,N_1626);
and U1976 (N_1976,N_1600,N_1728);
nand U1977 (N_1977,N_1613,N_1646);
or U1978 (N_1978,N_1648,N_1717);
and U1979 (N_1979,N_1797,N_1761);
or U1980 (N_1980,N_1664,N_1798);
nor U1981 (N_1981,N_1605,N_1738);
nand U1982 (N_1982,N_1729,N_1605);
and U1983 (N_1983,N_1712,N_1600);
or U1984 (N_1984,N_1741,N_1665);
and U1985 (N_1985,N_1624,N_1669);
nor U1986 (N_1986,N_1774,N_1648);
nand U1987 (N_1987,N_1623,N_1791);
and U1988 (N_1988,N_1702,N_1701);
and U1989 (N_1989,N_1627,N_1764);
or U1990 (N_1990,N_1692,N_1706);
nor U1991 (N_1991,N_1607,N_1689);
and U1992 (N_1992,N_1717,N_1794);
nand U1993 (N_1993,N_1745,N_1790);
nor U1994 (N_1994,N_1727,N_1688);
and U1995 (N_1995,N_1770,N_1764);
nor U1996 (N_1996,N_1785,N_1764);
nor U1997 (N_1997,N_1708,N_1669);
nor U1998 (N_1998,N_1711,N_1760);
and U1999 (N_1999,N_1648,N_1637);
or U2000 (N_2000,N_1852,N_1876);
nor U2001 (N_2001,N_1805,N_1879);
nor U2002 (N_2002,N_1954,N_1821);
nor U2003 (N_2003,N_1922,N_1806);
nor U2004 (N_2004,N_1895,N_1964);
and U2005 (N_2005,N_1938,N_1944);
or U2006 (N_2006,N_1856,N_1886);
nand U2007 (N_2007,N_1961,N_1847);
nand U2008 (N_2008,N_1953,N_1842);
and U2009 (N_2009,N_1940,N_1889);
and U2010 (N_2010,N_1880,N_1872);
or U2011 (N_2011,N_1991,N_1990);
nor U2012 (N_2012,N_1823,N_1900);
nand U2013 (N_2013,N_1892,N_1859);
or U2014 (N_2014,N_1808,N_1910);
nor U2015 (N_2015,N_1937,N_1832);
nor U2016 (N_2016,N_1897,N_1841);
or U2017 (N_2017,N_1827,N_1836);
xnor U2018 (N_2018,N_1845,N_1973);
nor U2019 (N_2019,N_1851,N_1955);
nand U2020 (N_2020,N_1812,N_1869);
nand U2021 (N_2021,N_1833,N_1920);
nand U2022 (N_2022,N_1941,N_1914);
nand U2023 (N_2023,N_1863,N_1804);
or U2024 (N_2024,N_1873,N_1919);
nor U2025 (N_2025,N_1989,N_1891);
nand U2026 (N_2026,N_1997,N_1800);
or U2027 (N_2027,N_1890,N_1868);
nor U2028 (N_2028,N_1967,N_1849);
nor U2029 (N_2029,N_1934,N_1916);
or U2030 (N_2030,N_1932,N_1903);
nand U2031 (N_2031,N_1896,N_1957);
nand U2032 (N_2032,N_1994,N_1913);
and U2033 (N_2033,N_1883,N_1998);
and U2034 (N_2034,N_1950,N_1894);
or U2035 (N_2035,N_1958,N_1871);
and U2036 (N_2036,N_1905,N_1815);
or U2037 (N_2037,N_1816,N_1855);
nor U2038 (N_2038,N_1906,N_1986);
nor U2039 (N_2039,N_1843,N_1899);
nor U2040 (N_2040,N_1942,N_1981);
nor U2041 (N_2041,N_1947,N_1881);
or U2042 (N_2042,N_1877,N_1930);
nand U2043 (N_2043,N_1860,N_1927);
and U2044 (N_2044,N_1918,N_1854);
and U2045 (N_2045,N_1817,N_1825);
nand U2046 (N_2046,N_1962,N_1908);
nand U2047 (N_2047,N_1875,N_1814);
and U2048 (N_2048,N_1819,N_1893);
xor U2049 (N_2049,N_1831,N_1933);
xnor U2050 (N_2050,N_1975,N_1963);
nand U2051 (N_2051,N_1884,N_1923);
nand U2052 (N_2052,N_1874,N_1966);
nand U2053 (N_2053,N_1987,N_1902);
xnor U2054 (N_2054,N_1822,N_1838);
nor U2055 (N_2055,N_1870,N_1952);
and U2056 (N_2056,N_1946,N_1960);
and U2057 (N_2057,N_1901,N_1943);
nand U2058 (N_2058,N_1861,N_1848);
nand U2059 (N_2059,N_1826,N_1904);
or U2060 (N_2060,N_1813,N_1965);
nand U2061 (N_2061,N_1988,N_1976);
or U2062 (N_2062,N_1850,N_1912);
or U2063 (N_2063,N_1969,N_1865);
or U2064 (N_2064,N_1939,N_1978);
or U2065 (N_2065,N_1835,N_1907);
or U2066 (N_2066,N_1971,N_1885);
nand U2067 (N_2067,N_1931,N_1810);
or U2068 (N_2068,N_1996,N_1985);
and U2069 (N_2069,N_1974,N_1830);
nand U2070 (N_2070,N_1917,N_1915);
nor U2071 (N_2071,N_1995,N_1984);
and U2072 (N_2072,N_1970,N_1811);
and U2073 (N_2073,N_1925,N_1935);
or U2074 (N_2074,N_1924,N_1807);
nor U2075 (N_2075,N_1982,N_1837);
or U2076 (N_2076,N_1911,N_1979);
or U2077 (N_2077,N_1834,N_1844);
and U2078 (N_2078,N_1867,N_1803);
nor U2079 (N_2079,N_1993,N_1949);
or U2080 (N_2080,N_1992,N_1983);
and U2081 (N_2081,N_1828,N_1929);
nand U2082 (N_2082,N_1959,N_1846);
or U2083 (N_2083,N_1928,N_1809);
nor U2084 (N_2084,N_1909,N_1945);
nand U2085 (N_2085,N_1824,N_1921);
nor U2086 (N_2086,N_1864,N_1980);
and U2087 (N_2087,N_1818,N_1898);
or U2088 (N_2088,N_1972,N_1820);
nor U2089 (N_2089,N_1968,N_1951);
or U2090 (N_2090,N_1948,N_1853);
and U2091 (N_2091,N_1801,N_1888);
and U2092 (N_2092,N_1862,N_1956);
nor U2093 (N_2093,N_1829,N_1857);
xor U2094 (N_2094,N_1840,N_1926);
nand U2095 (N_2095,N_1936,N_1839);
and U2096 (N_2096,N_1858,N_1878);
nand U2097 (N_2097,N_1802,N_1882);
nor U2098 (N_2098,N_1866,N_1977);
nor U2099 (N_2099,N_1999,N_1887);
or U2100 (N_2100,N_1899,N_1930);
nor U2101 (N_2101,N_1861,N_1966);
xnor U2102 (N_2102,N_1942,N_1923);
nor U2103 (N_2103,N_1809,N_1842);
and U2104 (N_2104,N_1892,N_1921);
and U2105 (N_2105,N_1845,N_1871);
or U2106 (N_2106,N_1920,N_1999);
or U2107 (N_2107,N_1836,N_1991);
xnor U2108 (N_2108,N_1952,N_1902);
nand U2109 (N_2109,N_1860,N_1926);
nor U2110 (N_2110,N_1929,N_1875);
nand U2111 (N_2111,N_1970,N_1924);
nand U2112 (N_2112,N_1866,N_1860);
nor U2113 (N_2113,N_1979,N_1978);
nor U2114 (N_2114,N_1882,N_1874);
or U2115 (N_2115,N_1936,N_1880);
nor U2116 (N_2116,N_1851,N_1896);
or U2117 (N_2117,N_1858,N_1814);
nand U2118 (N_2118,N_1808,N_1822);
nand U2119 (N_2119,N_1891,N_1910);
and U2120 (N_2120,N_1830,N_1986);
nor U2121 (N_2121,N_1807,N_1834);
nand U2122 (N_2122,N_1830,N_1904);
nand U2123 (N_2123,N_1913,N_1876);
nor U2124 (N_2124,N_1967,N_1841);
or U2125 (N_2125,N_1847,N_1878);
and U2126 (N_2126,N_1857,N_1840);
or U2127 (N_2127,N_1881,N_1855);
and U2128 (N_2128,N_1811,N_1953);
or U2129 (N_2129,N_1915,N_1986);
or U2130 (N_2130,N_1813,N_1870);
nor U2131 (N_2131,N_1822,N_1889);
nand U2132 (N_2132,N_1854,N_1983);
or U2133 (N_2133,N_1988,N_1874);
and U2134 (N_2134,N_1861,N_1818);
nand U2135 (N_2135,N_1925,N_1810);
nand U2136 (N_2136,N_1989,N_1851);
nor U2137 (N_2137,N_1977,N_1809);
nor U2138 (N_2138,N_1821,N_1826);
or U2139 (N_2139,N_1991,N_1935);
nand U2140 (N_2140,N_1802,N_1925);
nor U2141 (N_2141,N_1803,N_1812);
xnor U2142 (N_2142,N_1801,N_1929);
or U2143 (N_2143,N_1969,N_1844);
xor U2144 (N_2144,N_1902,N_1847);
nand U2145 (N_2145,N_1941,N_1983);
or U2146 (N_2146,N_1984,N_1951);
nor U2147 (N_2147,N_1831,N_1909);
nor U2148 (N_2148,N_1815,N_1928);
or U2149 (N_2149,N_1924,N_1890);
nand U2150 (N_2150,N_1915,N_1836);
or U2151 (N_2151,N_1810,N_1952);
or U2152 (N_2152,N_1905,N_1869);
and U2153 (N_2153,N_1864,N_1963);
or U2154 (N_2154,N_1912,N_1922);
and U2155 (N_2155,N_1808,N_1953);
nor U2156 (N_2156,N_1976,N_1958);
and U2157 (N_2157,N_1918,N_1831);
or U2158 (N_2158,N_1877,N_1882);
nor U2159 (N_2159,N_1930,N_1822);
and U2160 (N_2160,N_1886,N_1997);
and U2161 (N_2161,N_1804,N_1938);
and U2162 (N_2162,N_1823,N_1939);
or U2163 (N_2163,N_1942,N_1866);
nand U2164 (N_2164,N_1959,N_1875);
or U2165 (N_2165,N_1872,N_1819);
nor U2166 (N_2166,N_1961,N_1914);
and U2167 (N_2167,N_1848,N_1894);
nor U2168 (N_2168,N_1806,N_1800);
or U2169 (N_2169,N_1959,N_1969);
nand U2170 (N_2170,N_1821,N_1891);
nand U2171 (N_2171,N_1802,N_1820);
nor U2172 (N_2172,N_1803,N_1945);
or U2173 (N_2173,N_1991,N_1973);
nand U2174 (N_2174,N_1825,N_1869);
nor U2175 (N_2175,N_1835,N_1898);
or U2176 (N_2176,N_1851,N_1835);
nor U2177 (N_2177,N_1866,N_1820);
nor U2178 (N_2178,N_1957,N_1810);
or U2179 (N_2179,N_1894,N_1818);
nor U2180 (N_2180,N_1865,N_1895);
and U2181 (N_2181,N_1964,N_1982);
nor U2182 (N_2182,N_1890,N_1870);
nand U2183 (N_2183,N_1997,N_1827);
nor U2184 (N_2184,N_1991,N_1984);
and U2185 (N_2185,N_1898,N_1985);
and U2186 (N_2186,N_1943,N_1958);
nand U2187 (N_2187,N_1971,N_1940);
nor U2188 (N_2188,N_1876,N_1880);
or U2189 (N_2189,N_1873,N_1971);
nand U2190 (N_2190,N_1857,N_1838);
nand U2191 (N_2191,N_1964,N_1867);
or U2192 (N_2192,N_1975,N_1871);
or U2193 (N_2193,N_1983,N_1979);
xor U2194 (N_2194,N_1825,N_1823);
nor U2195 (N_2195,N_1829,N_1827);
and U2196 (N_2196,N_1966,N_1987);
or U2197 (N_2197,N_1883,N_1812);
or U2198 (N_2198,N_1926,N_1838);
nand U2199 (N_2199,N_1881,N_1880);
xor U2200 (N_2200,N_2103,N_2113);
and U2201 (N_2201,N_2162,N_2029);
and U2202 (N_2202,N_2196,N_2036);
or U2203 (N_2203,N_2011,N_2146);
xor U2204 (N_2204,N_2074,N_2182);
nor U2205 (N_2205,N_2129,N_2063);
nand U2206 (N_2206,N_2123,N_2032);
and U2207 (N_2207,N_2104,N_2060);
or U2208 (N_2208,N_2030,N_2086);
and U2209 (N_2209,N_2000,N_2093);
nand U2210 (N_2210,N_2066,N_2041);
or U2211 (N_2211,N_2018,N_2010);
nand U2212 (N_2212,N_2112,N_2140);
or U2213 (N_2213,N_2145,N_2124);
nand U2214 (N_2214,N_2147,N_2185);
nand U2215 (N_2215,N_2168,N_2007);
nor U2216 (N_2216,N_2133,N_2023);
nor U2217 (N_2217,N_2149,N_2002);
and U2218 (N_2218,N_2122,N_2025);
nand U2219 (N_2219,N_2096,N_2120);
nor U2220 (N_2220,N_2035,N_2083);
or U2221 (N_2221,N_2198,N_2087);
nor U2222 (N_2222,N_2097,N_2142);
nor U2223 (N_2223,N_2152,N_2056);
nor U2224 (N_2224,N_2057,N_2085);
or U2225 (N_2225,N_2115,N_2155);
nand U2226 (N_2226,N_2068,N_2090);
or U2227 (N_2227,N_2121,N_2038);
nor U2228 (N_2228,N_2079,N_2050);
nand U2229 (N_2229,N_2062,N_2101);
nor U2230 (N_2230,N_2191,N_2070);
nor U2231 (N_2231,N_2055,N_2033);
nor U2232 (N_2232,N_2179,N_2046);
and U2233 (N_2233,N_2110,N_2004);
nand U2234 (N_2234,N_2013,N_2001);
nand U2235 (N_2235,N_2137,N_2118);
nor U2236 (N_2236,N_2167,N_2020);
or U2237 (N_2237,N_2028,N_2067);
nand U2238 (N_2238,N_2014,N_2069);
nor U2239 (N_2239,N_2156,N_2178);
nor U2240 (N_2240,N_2027,N_2024);
and U2241 (N_2241,N_2106,N_2026);
or U2242 (N_2242,N_2076,N_2051);
or U2243 (N_2243,N_2190,N_2016);
nor U2244 (N_2244,N_2130,N_2095);
and U2245 (N_2245,N_2177,N_2009);
or U2246 (N_2246,N_2174,N_2037);
nand U2247 (N_2247,N_2102,N_2075);
nand U2248 (N_2248,N_2169,N_2164);
nand U2249 (N_2249,N_2126,N_2071);
nand U2250 (N_2250,N_2065,N_2089);
or U2251 (N_2251,N_2107,N_2144);
or U2252 (N_2252,N_2072,N_2015);
nor U2253 (N_2253,N_2143,N_2077);
or U2254 (N_2254,N_2170,N_2058);
and U2255 (N_2255,N_2100,N_2176);
nand U2256 (N_2256,N_2194,N_2134);
or U2257 (N_2257,N_2187,N_2017);
nand U2258 (N_2258,N_2084,N_2184);
or U2259 (N_2259,N_2091,N_2148);
nand U2260 (N_2260,N_2003,N_2008);
and U2261 (N_2261,N_2161,N_2098);
nor U2262 (N_2262,N_2138,N_2159);
and U2263 (N_2263,N_2158,N_2053);
nor U2264 (N_2264,N_2081,N_2078);
nor U2265 (N_2265,N_2111,N_2039);
and U2266 (N_2266,N_2092,N_2141);
nor U2267 (N_2267,N_2094,N_2189);
and U2268 (N_2268,N_2105,N_2108);
xor U2269 (N_2269,N_2054,N_2116);
or U2270 (N_2270,N_2193,N_2064);
nor U2271 (N_2271,N_2043,N_2151);
or U2272 (N_2272,N_2175,N_2042);
and U2273 (N_2273,N_2195,N_2173);
nand U2274 (N_2274,N_2199,N_2192);
or U2275 (N_2275,N_2136,N_2040);
nor U2276 (N_2276,N_2172,N_2031);
xnor U2277 (N_2277,N_2157,N_2127);
and U2278 (N_2278,N_2154,N_2135);
nor U2279 (N_2279,N_2153,N_2166);
and U2280 (N_2280,N_2171,N_2005);
or U2281 (N_2281,N_2006,N_2019);
nand U2282 (N_2282,N_2048,N_2049);
nor U2283 (N_2283,N_2099,N_2052);
xor U2284 (N_2284,N_2139,N_2119);
nand U2285 (N_2285,N_2163,N_2183);
and U2286 (N_2286,N_2047,N_2186);
or U2287 (N_2287,N_2117,N_2188);
nand U2288 (N_2288,N_2114,N_2131);
xor U2289 (N_2289,N_2180,N_2045);
and U2290 (N_2290,N_2128,N_2197);
or U2291 (N_2291,N_2165,N_2022);
or U2292 (N_2292,N_2109,N_2080);
or U2293 (N_2293,N_2132,N_2125);
nand U2294 (N_2294,N_2059,N_2021);
nand U2295 (N_2295,N_2044,N_2073);
nand U2296 (N_2296,N_2181,N_2088);
nand U2297 (N_2297,N_2150,N_2012);
nor U2298 (N_2298,N_2082,N_2061);
and U2299 (N_2299,N_2034,N_2160);
nor U2300 (N_2300,N_2186,N_2129);
or U2301 (N_2301,N_2025,N_2174);
nand U2302 (N_2302,N_2140,N_2192);
nand U2303 (N_2303,N_2015,N_2154);
or U2304 (N_2304,N_2137,N_2188);
nand U2305 (N_2305,N_2157,N_2120);
nand U2306 (N_2306,N_2154,N_2149);
or U2307 (N_2307,N_2171,N_2069);
or U2308 (N_2308,N_2156,N_2005);
xor U2309 (N_2309,N_2112,N_2072);
and U2310 (N_2310,N_2170,N_2038);
or U2311 (N_2311,N_2152,N_2150);
or U2312 (N_2312,N_2023,N_2055);
or U2313 (N_2313,N_2028,N_2094);
or U2314 (N_2314,N_2051,N_2010);
and U2315 (N_2315,N_2147,N_2001);
nand U2316 (N_2316,N_2138,N_2031);
and U2317 (N_2317,N_2038,N_2150);
and U2318 (N_2318,N_2060,N_2007);
or U2319 (N_2319,N_2156,N_2172);
or U2320 (N_2320,N_2043,N_2062);
and U2321 (N_2321,N_2037,N_2060);
or U2322 (N_2322,N_2180,N_2069);
or U2323 (N_2323,N_2157,N_2175);
and U2324 (N_2324,N_2081,N_2054);
nand U2325 (N_2325,N_2184,N_2081);
nand U2326 (N_2326,N_2016,N_2163);
nor U2327 (N_2327,N_2155,N_2101);
nor U2328 (N_2328,N_2120,N_2044);
and U2329 (N_2329,N_2048,N_2026);
nand U2330 (N_2330,N_2010,N_2082);
nor U2331 (N_2331,N_2172,N_2005);
or U2332 (N_2332,N_2143,N_2121);
nor U2333 (N_2333,N_2031,N_2098);
nand U2334 (N_2334,N_2086,N_2193);
or U2335 (N_2335,N_2183,N_2125);
nand U2336 (N_2336,N_2179,N_2018);
nand U2337 (N_2337,N_2011,N_2025);
nor U2338 (N_2338,N_2069,N_2135);
nor U2339 (N_2339,N_2021,N_2194);
nand U2340 (N_2340,N_2038,N_2084);
or U2341 (N_2341,N_2071,N_2129);
xnor U2342 (N_2342,N_2181,N_2121);
nor U2343 (N_2343,N_2190,N_2129);
or U2344 (N_2344,N_2096,N_2182);
nor U2345 (N_2345,N_2018,N_2136);
or U2346 (N_2346,N_2075,N_2087);
nor U2347 (N_2347,N_2156,N_2174);
nor U2348 (N_2348,N_2117,N_2034);
nor U2349 (N_2349,N_2049,N_2163);
and U2350 (N_2350,N_2092,N_2090);
nand U2351 (N_2351,N_2156,N_2085);
and U2352 (N_2352,N_2112,N_2002);
or U2353 (N_2353,N_2037,N_2073);
and U2354 (N_2354,N_2064,N_2035);
nand U2355 (N_2355,N_2190,N_2041);
or U2356 (N_2356,N_2106,N_2170);
or U2357 (N_2357,N_2075,N_2152);
nor U2358 (N_2358,N_2081,N_2101);
nor U2359 (N_2359,N_2119,N_2064);
nor U2360 (N_2360,N_2099,N_2144);
or U2361 (N_2361,N_2105,N_2114);
or U2362 (N_2362,N_2076,N_2110);
xor U2363 (N_2363,N_2058,N_2009);
nor U2364 (N_2364,N_2187,N_2042);
or U2365 (N_2365,N_2039,N_2103);
nor U2366 (N_2366,N_2091,N_2153);
xor U2367 (N_2367,N_2127,N_2021);
nor U2368 (N_2368,N_2082,N_2020);
and U2369 (N_2369,N_2130,N_2154);
nor U2370 (N_2370,N_2161,N_2017);
nand U2371 (N_2371,N_2066,N_2129);
nor U2372 (N_2372,N_2136,N_2001);
nand U2373 (N_2373,N_2107,N_2017);
nand U2374 (N_2374,N_2062,N_2171);
nand U2375 (N_2375,N_2016,N_2054);
and U2376 (N_2376,N_2051,N_2086);
or U2377 (N_2377,N_2120,N_2059);
and U2378 (N_2378,N_2122,N_2010);
or U2379 (N_2379,N_2117,N_2052);
and U2380 (N_2380,N_2163,N_2136);
nor U2381 (N_2381,N_2003,N_2028);
or U2382 (N_2382,N_2027,N_2011);
and U2383 (N_2383,N_2167,N_2032);
nand U2384 (N_2384,N_2193,N_2083);
nor U2385 (N_2385,N_2019,N_2151);
and U2386 (N_2386,N_2002,N_2057);
and U2387 (N_2387,N_2117,N_2028);
nand U2388 (N_2388,N_2094,N_2147);
nand U2389 (N_2389,N_2199,N_2051);
nand U2390 (N_2390,N_2086,N_2110);
and U2391 (N_2391,N_2060,N_2112);
nor U2392 (N_2392,N_2042,N_2129);
nand U2393 (N_2393,N_2086,N_2153);
nand U2394 (N_2394,N_2199,N_2170);
nand U2395 (N_2395,N_2104,N_2066);
nand U2396 (N_2396,N_2164,N_2023);
or U2397 (N_2397,N_2198,N_2068);
and U2398 (N_2398,N_2007,N_2142);
nand U2399 (N_2399,N_2192,N_2151);
or U2400 (N_2400,N_2205,N_2386);
and U2401 (N_2401,N_2223,N_2384);
and U2402 (N_2402,N_2275,N_2373);
nor U2403 (N_2403,N_2243,N_2244);
nor U2404 (N_2404,N_2310,N_2246);
nor U2405 (N_2405,N_2251,N_2370);
xnor U2406 (N_2406,N_2253,N_2250);
and U2407 (N_2407,N_2342,N_2258);
nor U2408 (N_2408,N_2354,N_2255);
nor U2409 (N_2409,N_2312,N_2378);
nand U2410 (N_2410,N_2278,N_2339);
nand U2411 (N_2411,N_2229,N_2272);
and U2412 (N_2412,N_2208,N_2252);
and U2413 (N_2413,N_2388,N_2376);
nor U2414 (N_2414,N_2207,N_2287);
and U2415 (N_2415,N_2303,N_2201);
or U2416 (N_2416,N_2397,N_2353);
nor U2417 (N_2417,N_2290,N_2351);
or U2418 (N_2418,N_2337,N_2359);
nand U2419 (N_2419,N_2219,N_2263);
and U2420 (N_2420,N_2295,N_2203);
nand U2421 (N_2421,N_2230,N_2349);
or U2422 (N_2422,N_2224,N_2227);
or U2423 (N_2423,N_2330,N_2281);
nand U2424 (N_2424,N_2276,N_2274);
and U2425 (N_2425,N_2222,N_2344);
or U2426 (N_2426,N_2226,N_2288);
and U2427 (N_2427,N_2273,N_2238);
or U2428 (N_2428,N_2316,N_2328);
nand U2429 (N_2429,N_2200,N_2338);
nand U2430 (N_2430,N_2358,N_2268);
nand U2431 (N_2431,N_2247,N_2314);
nor U2432 (N_2432,N_2379,N_2204);
or U2433 (N_2433,N_2395,N_2361);
nand U2434 (N_2434,N_2383,N_2266);
and U2435 (N_2435,N_2368,N_2225);
xnor U2436 (N_2436,N_2381,N_2367);
or U2437 (N_2437,N_2382,N_2257);
xor U2438 (N_2438,N_2236,N_2347);
nand U2439 (N_2439,N_2283,N_2341);
nand U2440 (N_2440,N_2309,N_2277);
nor U2441 (N_2441,N_2299,N_2391);
nand U2442 (N_2442,N_2389,N_2377);
and U2443 (N_2443,N_2321,N_2327);
or U2444 (N_2444,N_2352,N_2390);
or U2445 (N_2445,N_2302,N_2211);
or U2446 (N_2446,N_2322,N_2260);
and U2447 (N_2447,N_2256,N_2374);
nor U2448 (N_2448,N_2387,N_2325);
or U2449 (N_2449,N_2291,N_2311);
or U2450 (N_2450,N_2293,N_2210);
or U2451 (N_2451,N_2315,N_2217);
and U2452 (N_2452,N_2396,N_2215);
nor U2453 (N_2453,N_2228,N_2317);
nand U2454 (N_2454,N_2232,N_2369);
and U2455 (N_2455,N_2221,N_2362);
or U2456 (N_2456,N_2304,N_2394);
nand U2457 (N_2457,N_2267,N_2206);
nand U2458 (N_2458,N_2264,N_2297);
nand U2459 (N_2459,N_2305,N_2242);
nand U2460 (N_2460,N_2319,N_2346);
or U2461 (N_2461,N_2340,N_2216);
nand U2462 (N_2462,N_2218,N_2307);
or U2463 (N_2463,N_2331,N_2363);
or U2464 (N_2464,N_2350,N_2333);
nand U2465 (N_2465,N_2392,N_2393);
and U2466 (N_2466,N_2356,N_2240);
nand U2467 (N_2467,N_2294,N_2329);
nand U2468 (N_2468,N_2345,N_2237);
nand U2469 (N_2469,N_2231,N_2343);
nor U2470 (N_2470,N_2332,N_2323);
or U2471 (N_2471,N_2261,N_2360);
nand U2472 (N_2472,N_2245,N_2326);
or U2473 (N_2473,N_2259,N_2306);
nor U2474 (N_2474,N_2313,N_2300);
nand U2475 (N_2475,N_2213,N_2355);
nor U2476 (N_2476,N_2289,N_2399);
or U2477 (N_2477,N_2280,N_2398);
and U2478 (N_2478,N_2212,N_2241);
nor U2479 (N_2479,N_2336,N_2233);
or U2480 (N_2480,N_2282,N_2286);
nor U2481 (N_2481,N_2318,N_2234);
nor U2482 (N_2482,N_2269,N_2334);
or U2483 (N_2483,N_2371,N_2271);
or U2484 (N_2484,N_2301,N_2364);
xor U2485 (N_2485,N_2249,N_2335);
nor U2486 (N_2486,N_2284,N_2366);
or U2487 (N_2487,N_2385,N_2375);
or U2488 (N_2488,N_2254,N_2357);
nand U2489 (N_2489,N_2380,N_2308);
and U2490 (N_2490,N_2220,N_2270);
nor U2491 (N_2491,N_2285,N_2265);
or U2492 (N_2492,N_2214,N_2202);
and U2493 (N_2493,N_2324,N_2298);
or U2494 (N_2494,N_2296,N_2262);
and U2495 (N_2495,N_2320,N_2348);
nand U2496 (N_2496,N_2279,N_2235);
or U2497 (N_2497,N_2292,N_2365);
and U2498 (N_2498,N_2209,N_2372);
and U2499 (N_2499,N_2248,N_2239);
nor U2500 (N_2500,N_2348,N_2288);
nor U2501 (N_2501,N_2338,N_2264);
nand U2502 (N_2502,N_2239,N_2218);
nand U2503 (N_2503,N_2296,N_2376);
nor U2504 (N_2504,N_2290,N_2261);
or U2505 (N_2505,N_2384,N_2289);
nor U2506 (N_2506,N_2210,N_2358);
nor U2507 (N_2507,N_2335,N_2236);
nand U2508 (N_2508,N_2310,N_2248);
nand U2509 (N_2509,N_2247,N_2232);
nor U2510 (N_2510,N_2312,N_2229);
nand U2511 (N_2511,N_2241,N_2382);
nor U2512 (N_2512,N_2389,N_2358);
or U2513 (N_2513,N_2315,N_2267);
nand U2514 (N_2514,N_2332,N_2374);
nor U2515 (N_2515,N_2262,N_2359);
or U2516 (N_2516,N_2204,N_2215);
nand U2517 (N_2517,N_2314,N_2304);
nor U2518 (N_2518,N_2303,N_2293);
and U2519 (N_2519,N_2334,N_2328);
and U2520 (N_2520,N_2390,N_2294);
nand U2521 (N_2521,N_2271,N_2211);
nand U2522 (N_2522,N_2265,N_2271);
and U2523 (N_2523,N_2225,N_2348);
nand U2524 (N_2524,N_2200,N_2377);
nand U2525 (N_2525,N_2353,N_2369);
or U2526 (N_2526,N_2255,N_2344);
nor U2527 (N_2527,N_2299,N_2205);
or U2528 (N_2528,N_2297,N_2353);
nand U2529 (N_2529,N_2343,N_2249);
and U2530 (N_2530,N_2396,N_2310);
and U2531 (N_2531,N_2309,N_2247);
nor U2532 (N_2532,N_2318,N_2352);
nand U2533 (N_2533,N_2331,N_2377);
nor U2534 (N_2534,N_2364,N_2352);
or U2535 (N_2535,N_2290,N_2339);
nand U2536 (N_2536,N_2226,N_2269);
or U2537 (N_2537,N_2393,N_2201);
xnor U2538 (N_2538,N_2368,N_2267);
or U2539 (N_2539,N_2214,N_2300);
and U2540 (N_2540,N_2305,N_2338);
and U2541 (N_2541,N_2202,N_2336);
nand U2542 (N_2542,N_2273,N_2268);
nand U2543 (N_2543,N_2330,N_2271);
nand U2544 (N_2544,N_2393,N_2352);
or U2545 (N_2545,N_2335,N_2269);
and U2546 (N_2546,N_2340,N_2259);
nand U2547 (N_2547,N_2387,N_2353);
nor U2548 (N_2548,N_2202,N_2215);
or U2549 (N_2549,N_2257,N_2285);
and U2550 (N_2550,N_2359,N_2239);
nor U2551 (N_2551,N_2202,N_2349);
or U2552 (N_2552,N_2214,N_2367);
and U2553 (N_2553,N_2356,N_2340);
nand U2554 (N_2554,N_2209,N_2336);
nor U2555 (N_2555,N_2290,N_2285);
nand U2556 (N_2556,N_2388,N_2313);
nand U2557 (N_2557,N_2351,N_2267);
nor U2558 (N_2558,N_2268,N_2264);
nand U2559 (N_2559,N_2276,N_2278);
xnor U2560 (N_2560,N_2259,N_2318);
and U2561 (N_2561,N_2277,N_2326);
nor U2562 (N_2562,N_2248,N_2254);
nand U2563 (N_2563,N_2396,N_2326);
nand U2564 (N_2564,N_2258,N_2275);
xor U2565 (N_2565,N_2242,N_2288);
and U2566 (N_2566,N_2291,N_2362);
or U2567 (N_2567,N_2393,N_2229);
and U2568 (N_2568,N_2294,N_2354);
or U2569 (N_2569,N_2278,N_2309);
and U2570 (N_2570,N_2329,N_2206);
nor U2571 (N_2571,N_2235,N_2393);
or U2572 (N_2572,N_2376,N_2339);
xnor U2573 (N_2573,N_2280,N_2336);
nand U2574 (N_2574,N_2385,N_2393);
nand U2575 (N_2575,N_2318,N_2203);
or U2576 (N_2576,N_2232,N_2208);
nor U2577 (N_2577,N_2208,N_2235);
or U2578 (N_2578,N_2280,N_2239);
nand U2579 (N_2579,N_2329,N_2216);
or U2580 (N_2580,N_2239,N_2249);
nor U2581 (N_2581,N_2240,N_2310);
nor U2582 (N_2582,N_2361,N_2375);
or U2583 (N_2583,N_2209,N_2393);
nor U2584 (N_2584,N_2385,N_2212);
or U2585 (N_2585,N_2367,N_2281);
nand U2586 (N_2586,N_2332,N_2283);
nor U2587 (N_2587,N_2302,N_2221);
nor U2588 (N_2588,N_2269,N_2353);
nand U2589 (N_2589,N_2262,N_2252);
xor U2590 (N_2590,N_2381,N_2373);
xnor U2591 (N_2591,N_2208,N_2202);
nand U2592 (N_2592,N_2368,N_2377);
and U2593 (N_2593,N_2297,N_2391);
nor U2594 (N_2594,N_2371,N_2275);
and U2595 (N_2595,N_2281,N_2212);
or U2596 (N_2596,N_2358,N_2264);
nand U2597 (N_2597,N_2389,N_2310);
or U2598 (N_2598,N_2269,N_2288);
nor U2599 (N_2599,N_2281,N_2393);
nand U2600 (N_2600,N_2489,N_2423);
and U2601 (N_2601,N_2509,N_2422);
nor U2602 (N_2602,N_2451,N_2404);
nand U2603 (N_2603,N_2526,N_2513);
and U2604 (N_2604,N_2493,N_2510);
nand U2605 (N_2605,N_2420,N_2574);
nand U2606 (N_2606,N_2432,N_2563);
or U2607 (N_2607,N_2545,N_2441);
nor U2608 (N_2608,N_2477,N_2452);
nand U2609 (N_2609,N_2401,N_2400);
nor U2610 (N_2610,N_2425,N_2564);
or U2611 (N_2611,N_2478,N_2487);
nand U2612 (N_2612,N_2462,N_2507);
or U2613 (N_2613,N_2483,N_2557);
and U2614 (N_2614,N_2529,N_2535);
nand U2615 (N_2615,N_2435,N_2490);
and U2616 (N_2616,N_2572,N_2496);
nor U2617 (N_2617,N_2543,N_2522);
nand U2618 (N_2618,N_2499,N_2485);
nand U2619 (N_2619,N_2559,N_2537);
or U2620 (N_2620,N_2551,N_2542);
and U2621 (N_2621,N_2455,N_2494);
nand U2622 (N_2622,N_2411,N_2479);
nor U2623 (N_2623,N_2544,N_2514);
nand U2624 (N_2624,N_2589,N_2586);
nor U2625 (N_2625,N_2488,N_2474);
nor U2626 (N_2626,N_2556,N_2534);
and U2627 (N_2627,N_2596,N_2502);
and U2628 (N_2628,N_2426,N_2541);
nand U2629 (N_2629,N_2481,N_2443);
nand U2630 (N_2630,N_2552,N_2464);
nor U2631 (N_2631,N_2469,N_2466);
nand U2632 (N_2632,N_2566,N_2593);
nor U2633 (N_2633,N_2573,N_2444);
nand U2634 (N_2634,N_2575,N_2491);
nand U2635 (N_2635,N_2471,N_2583);
or U2636 (N_2636,N_2506,N_2528);
nor U2637 (N_2637,N_2533,N_2503);
or U2638 (N_2638,N_2431,N_2584);
and U2639 (N_2639,N_2531,N_2456);
nor U2640 (N_2640,N_2550,N_2585);
and U2641 (N_2641,N_2473,N_2580);
and U2642 (N_2642,N_2438,N_2412);
or U2643 (N_2643,N_2591,N_2418);
or U2644 (N_2644,N_2517,N_2549);
or U2645 (N_2645,N_2414,N_2495);
or U2646 (N_2646,N_2527,N_2558);
and U2647 (N_2647,N_2470,N_2520);
nor U2648 (N_2648,N_2599,N_2565);
and U2649 (N_2649,N_2597,N_2561);
nor U2650 (N_2650,N_2467,N_2486);
or U2651 (N_2651,N_2468,N_2571);
or U2652 (N_2652,N_2595,N_2447);
or U2653 (N_2653,N_2405,N_2454);
and U2654 (N_2654,N_2523,N_2582);
nand U2655 (N_2655,N_2560,N_2568);
and U2656 (N_2656,N_2419,N_2449);
nand U2657 (N_2657,N_2436,N_2590);
nor U2658 (N_2658,N_2463,N_2465);
or U2659 (N_2659,N_2592,N_2539);
nor U2660 (N_2660,N_2407,N_2415);
nand U2661 (N_2661,N_2598,N_2480);
or U2662 (N_2662,N_2555,N_2588);
nand U2663 (N_2663,N_2554,N_2525);
xor U2664 (N_2664,N_2562,N_2428);
nand U2665 (N_2665,N_2538,N_2413);
xnor U2666 (N_2666,N_2442,N_2578);
or U2667 (N_2667,N_2475,N_2433);
or U2668 (N_2668,N_2516,N_2421);
nor U2669 (N_2669,N_2448,N_2445);
nand U2670 (N_2670,N_2492,N_2505);
nand U2671 (N_2671,N_2403,N_2417);
and U2672 (N_2672,N_2524,N_2532);
or U2673 (N_2673,N_2504,N_2406);
or U2674 (N_2674,N_2547,N_2446);
nand U2675 (N_2675,N_2437,N_2472);
and U2676 (N_2676,N_2546,N_2515);
nor U2677 (N_2677,N_2461,N_2427);
nand U2678 (N_2678,N_2594,N_2484);
xor U2679 (N_2679,N_2518,N_2453);
nor U2680 (N_2680,N_2577,N_2587);
and U2681 (N_2681,N_2458,N_2530);
nand U2682 (N_2682,N_2576,N_2402);
nand U2683 (N_2683,N_2459,N_2540);
or U2684 (N_2684,N_2553,N_2511);
nand U2685 (N_2685,N_2439,N_2536);
nand U2686 (N_2686,N_2429,N_2424);
and U2687 (N_2687,N_2460,N_2498);
nor U2688 (N_2688,N_2476,N_2567);
and U2689 (N_2689,N_2521,N_2434);
and U2690 (N_2690,N_2416,N_2497);
and U2691 (N_2691,N_2457,N_2450);
nand U2692 (N_2692,N_2501,N_2500);
and U2693 (N_2693,N_2519,N_2430);
or U2694 (N_2694,N_2569,N_2508);
and U2695 (N_2695,N_2548,N_2409);
and U2696 (N_2696,N_2581,N_2482);
and U2697 (N_2697,N_2408,N_2570);
nor U2698 (N_2698,N_2410,N_2440);
nand U2699 (N_2699,N_2579,N_2512);
nor U2700 (N_2700,N_2430,N_2523);
nor U2701 (N_2701,N_2536,N_2515);
or U2702 (N_2702,N_2480,N_2492);
nor U2703 (N_2703,N_2571,N_2537);
or U2704 (N_2704,N_2526,N_2435);
xor U2705 (N_2705,N_2536,N_2589);
nand U2706 (N_2706,N_2585,N_2514);
nor U2707 (N_2707,N_2594,N_2420);
nor U2708 (N_2708,N_2524,N_2487);
and U2709 (N_2709,N_2567,N_2406);
or U2710 (N_2710,N_2413,N_2561);
and U2711 (N_2711,N_2532,N_2467);
and U2712 (N_2712,N_2474,N_2507);
or U2713 (N_2713,N_2461,N_2482);
nor U2714 (N_2714,N_2542,N_2493);
and U2715 (N_2715,N_2483,N_2480);
nor U2716 (N_2716,N_2521,N_2557);
or U2717 (N_2717,N_2509,N_2429);
and U2718 (N_2718,N_2402,N_2505);
nor U2719 (N_2719,N_2587,N_2445);
or U2720 (N_2720,N_2480,N_2512);
or U2721 (N_2721,N_2515,N_2538);
and U2722 (N_2722,N_2594,N_2523);
nor U2723 (N_2723,N_2483,N_2425);
nand U2724 (N_2724,N_2415,N_2574);
and U2725 (N_2725,N_2444,N_2458);
nor U2726 (N_2726,N_2536,N_2413);
or U2727 (N_2727,N_2485,N_2521);
and U2728 (N_2728,N_2416,N_2477);
and U2729 (N_2729,N_2591,N_2430);
nand U2730 (N_2730,N_2517,N_2538);
nand U2731 (N_2731,N_2415,N_2432);
nor U2732 (N_2732,N_2502,N_2459);
or U2733 (N_2733,N_2475,N_2566);
and U2734 (N_2734,N_2452,N_2432);
nand U2735 (N_2735,N_2425,N_2438);
nand U2736 (N_2736,N_2594,N_2570);
nor U2737 (N_2737,N_2487,N_2461);
and U2738 (N_2738,N_2584,N_2567);
and U2739 (N_2739,N_2437,N_2507);
nor U2740 (N_2740,N_2547,N_2464);
nand U2741 (N_2741,N_2562,N_2596);
and U2742 (N_2742,N_2436,N_2516);
or U2743 (N_2743,N_2416,N_2526);
nand U2744 (N_2744,N_2436,N_2419);
and U2745 (N_2745,N_2429,N_2572);
nor U2746 (N_2746,N_2487,N_2413);
nand U2747 (N_2747,N_2423,N_2450);
or U2748 (N_2748,N_2500,N_2482);
nand U2749 (N_2749,N_2589,N_2466);
nand U2750 (N_2750,N_2478,N_2444);
or U2751 (N_2751,N_2456,N_2559);
or U2752 (N_2752,N_2567,N_2529);
nand U2753 (N_2753,N_2574,N_2449);
or U2754 (N_2754,N_2562,N_2563);
nand U2755 (N_2755,N_2553,N_2582);
nor U2756 (N_2756,N_2464,N_2585);
nand U2757 (N_2757,N_2475,N_2491);
nand U2758 (N_2758,N_2474,N_2546);
nor U2759 (N_2759,N_2507,N_2580);
nand U2760 (N_2760,N_2416,N_2506);
nand U2761 (N_2761,N_2503,N_2569);
or U2762 (N_2762,N_2574,N_2485);
nand U2763 (N_2763,N_2426,N_2439);
or U2764 (N_2764,N_2475,N_2575);
or U2765 (N_2765,N_2489,N_2491);
nor U2766 (N_2766,N_2403,N_2443);
and U2767 (N_2767,N_2538,N_2421);
nand U2768 (N_2768,N_2563,N_2575);
and U2769 (N_2769,N_2425,N_2577);
nor U2770 (N_2770,N_2417,N_2584);
nor U2771 (N_2771,N_2471,N_2527);
nor U2772 (N_2772,N_2524,N_2481);
and U2773 (N_2773,N_2482,N_2418);
nor U2774 (N_2774,N_2592,N_2408);
and U2775 (N_2775,N_2528,N_2478);
and U2776 (N_2776,N_2520,N_2501);
nand U2777 (N_2777,N_2502,N_2588);
nand U2778 (N_2778,N_2594,N_2427);
nor U2779 (N_2779,N_2506,N_2524);
nand U2780 (N_2780,N_2565,N_2436);
nor U2781 (N_2781,N_2446,N_2475);
nand U2782 (N_2782,N_2481,N_2599);
and U2783 (N_2783,N_2570,N_2540);
or U2784 (N_2784,N_2503,N_2571);
nor U2785 (N_2785,N_2499,N_2525);
nand U2786 (N_2786,N_2525,N_2458);
nor U2787 (N_2787,N_2495,N_2520);
or U2788 (N_2788,N_2545,N_2531);
or U2789 (N_2789,N_2458,N_2449);
or U2790 (N_2790,N_2568,N_2567);
or U2791 (N_2791,N_2429,N_2512);
nor U2792 (N_2792,N_2459,N_2435);
and U2793 (N_2793,N_2438,N_2543);
nor U2794 (N_2794,N_2449,N_2537);
or U2795 (N_2795,N_2577,N_2503);
nor U2796 (N_2796,N_2473,N_2555);
nor U2797 (N_2797,N_2443,N_2445);
nand U2798 (N_2798,N_2438,N_2558);
nand U2799 (N_2799,N_2402,N_2446);
or U2800 (N_2800,N_2724,N_2686);
and U2801 (N_2801,N_2655,N_2691);
nand U2802 (N_2802,N_2778,N_2782);
xnor U2803 (N_2803,N_2642,N_2768);
and U2804 (N_2804,N_2639,N_2759);
and U2805 (N_2805,N_2632,N_2758);
or U2806 (N_2806,N_2706,N_2719);
nand U2807 (N_2807,N_2659,N_2777);
and U2808 (N_2808,N_2715,N_2710);
nor U2809 (N_2809,N_2722,N_2741);
nor U2810 (N_2810,N_2701,N_2736);
nand U2811 (N_2811,N_2776,N_2646);
or U2812 (N_2812,N_2631,N_2624);
nor U2813 (N_2813,N_2652,N_2713);
nand U2814 (N_2814,N_2723,N_2638);
nor U2815 (N_2815,N_2791,N_2618);
and U2816 (N_2816,N_2787,N_2679);
nor U2817 (N_2817,N_2697,N_2752);
and U2818 (N_2818,N_2689,N_2767);
nand U2819 (N_2819,N_2772,N_2685);
nand U2820 (N_2820,N_2643,N_2771);
nor U2821 (N_2821,N_2673,N_2727);
and U2822 (N_2822,N_2645,N_2731);
and U2823 (N_2823,N_2790,N_2665);
and U2824 (N_2824,N_2675,N_2725);
and U2825 (N_2825,N_2792,N_2661);
or U2826 (N_2826,N_2630,N_2784);
nor U2827 (N_2827,N_2766,N_2795);
xor U2828 (N_2828,N_2677,N_2636);
and U2829 (N_2829,N_2781,N_2640);
and U2830 (N_2830,N_2696,N_2730);
nor U2831 (N_2831,N_2743,N_2605);
or U2832 (N_2832,N_2705,N_2666);
nor U2833 (N_2833,N_2756,N_2693);
nand U2834 (N_2834,N_2692,N_2629);
and U2835 (N_2835,N_2680,N_2797);
nand U2836 (N_2836,N_2603,N_2614);
and U2837 (N_2837,N_2793,N_2600);
nor U2838 (N_2838,N_2746,N_2647);
nor U2839 (N_2839,N_2670,N_2611);
nor U2840 (N_2840,N_2668,N_2607);
nand U2841 (N_2841,N_2601,N_2667);
or U2842 (N_2842,N_2606,N_2775);
or U2843 (N_2843,N_2729,N_2650);
nand U2844 (N_2844,N_2742,N_2712);
and U2845 (N_2845,N_2763,N_2751);
nor U2846 (N_2846,N_2699,N_2684);
and U2847 (N_2847,N_2663,N_2740);
nor U2848 (N_2848,N_2760,N_2744);
xor U2849 (N_2849,N_2608,N_2604);
nor U2850 (N_2850,N_2620,N_2602);
or U2851 (N_2851,N_2621,N_2613);
or U2852 (N_2852,N_2669,N_2714);
nand U2853 (N_2853,N_2798,N_2779);
nand U2854 (N_2854,N_2735,N_2757);
nand U2855 (N_2855,N_2783,N_2657);
and U2856 (N_2856,N_2644,N_2754);
nand U2857 (N_2857,N_2761,N_2788);
or U2858 (N_2858,N_2609,N_2702);
nor U2859 (N_2859,N_2635,N_2708);
or U2860 (N_2860,N_2648,N_2749);
nor U2861 (N_2861,N_2615,N_2733);
or U2862 (N_2862,N_2739,N_2785);
and U2863 (N_2863,N_2682,N_2617);
nand U2864 (N_2864,N_2726,N_2737);
and U2865 (N_2865,N_2773,N_2745);
and U2866 (N_2866,N_2678,N_2695);
or U2867 (N_2867,N_2641,N_2672);
nor U2868 (N_2868,N_2738,N_2664);
or U2869 (N_2869,N_2780,N_2703);
or U2870 (N_2870,N_2654,N_2720);
and U2871 (N_2871,N_2612,N_2649);
nor U2872 (N_2872,N_2626,N_2616);
nor U2873 (N_2873,N_2764,N_2694);
or U2874 (N_2874,N_2681,N_2799);
and U2875 (N_2875,N_2707,N_2728);
nand U2876 (N_2876,N_2747,N_2765);
nand U2877 (N_2877,N_2688,N_2789);
nor U2878 (N_2878,N_2674,N_2623);
nand U2879 (N_2879,N_2671,N_2721);
and U2880 (N_2880,N_2748,N_2633);
or U2881 (N_2881,N_2716,N_2734);
nand U2882 (N_2882,N_2711,N_2676);
nand U2883 (N_2883,N_2619,N_2651);
nand U2884 (N_2884,N_2774,N_2660);
or U2885 (N_2885,N_2750,N_2622);
nand U2886 (N_2886,N_2794,N_2770);
or U2887 (N_2887,N_2717,N_2718);
nand U2888 (N_2888,N_2796,N_2656);
nor U2889 (N_2889,N_2653,N_2786);
and U2890 (N_2890,N_2662,N_2610);
and U2891 (N_2891,N_2753,N_2634);
nand U2892 (N_2892,N_2683,N_2658);
or U2893 (N_2893,N_2769,N_2627);
or U2894 (N_2894,N_2732,N_2625);
or U2895 (N_2895,N_2762,N_2698);
nand U2896 (N_2896,N_2628,N_2755);
nor U2897 (N_2897,N_2704,N_2709);
or U2898 (N_2898,N_2637,N_2690);
nor U2899 (N_2899,N_2700,N_2687);
nor U2900 (N_2900,N_2764,N_2769);
nor U2901 (N_2901,N_2797,N_2676);
nor U2902 (N_2902,N_2667,N_2727);
or U2903 (N_2903,N_2628,N_2766);
nor U2904 (N_2904,N_2656,N_2600);
nand U2905 (N_2905,N_2620,N_2755);
nand U2906 (N_2906,N_2680,N_2666);
or U2907 (N_2907,N_2789,N_2761);
nor U2908 (N_2908,N_2638,N_2710);
and U2909 (N_2909,N_2642,N_2705);
nand U2910 (N_2910,N_2665,N_2619);
nand U2911 (N_2911,N_2772,N_2730);
and U2912 (N_2912,N_2701,N_2772);
or U2913 (N_2913,N_2647,N_2629);
nand U2914 (N_2914,N_2781,N_2635);
xnor U2915 (N_2915,N_2665,N_2689);
nand U2916 (N_2916,N_2634,N_2736);
and U2917 (N_2917,N_2620,N_2735);
and U2918 (N_2918,N_2776,N_2774);
nand U2919 (N_2919,N_2644,N_2797);
or U2920 (N_2920,N_2798,N_2785);
nand U2921 (N_2921,N_2750,N_2674);
nor U2922 (N_2922,N_2777,N_2713);
and U2923 (N_2923,N_2746,N_2643);
nand U2924 (N_2924,N_2605,N_2711);
or U2925 (N_2925,N_2766,N_2602);
nand U2926 (N_2926,N_2786,N_2761);
nand U2927 (N_2927,N_2747,N_2626);
or U2928 (N_2928,N_2657,N_2662);
or U2929 (N_2929,N_2702,N_2698);
and U2930 (N_2930,N_2697,N_2786);
or U2931 (N_2931,N_2666,N_2653);
nor U2932 (N_2932,N_2785,N_2689);
nor U2933 (N_2933,N_2740,N_2708);
and U2934 (N_2934,N_2622,N_2798);
nand U2935 (N_2935,N_2637,N_2720);
nand U2936 (N_2936,N_2703,N_2608);
or U2937 (N_2937,N_2734,N_2702);
and U2938 (N_2938,N_2671,N_2708);
or U2939 (N_2939,N_2657,N_2616);
or U2940 (N_2940,N_2714,N_2654);
or U2941 (N_2941,N_2703,N_2664);
xor U2942 (N_2942,N_2798,N_2792);
nor U2943 (N_2943,N_2724,N_2768);
nand U2944 (N_2944,N_2639,N_2641);
nand U2945 (N_2945,N_2660,N_2698);
and U2946 (N_2946,N_2724,N_2783);
nand U2947 (N_2947,N_2731,N_2791);
and U2948 (N_2948,N_2709,N_2697);
and U2949 (N_2949,N_2784,N_2796);
nor U2950 (N_2950,N_2787,N_2714);
and U2951 (N_2951,N_2765,N_2775);
or U2952 (N_2952,N_2608,N_2689);
and U2953 (N_2953,N_2720,N_2757);
or U2954 (N_2954,N_2735,N_2649);
nor U2955 (N_2955,N_2635,N_2764);
or U2956 (N_2956,N_2736,N_2779);
and U2957 (N_2957,N_2744,N_2627);
nand U2958 (N_2958,N_2697,N_2674);
nand U2959 (N_2959,N_2642,N_2666);
nor U2960 (N_2960,N_2600,N_2746);
nand U2961 (N_2961,N_2677,N_2731);
or U2962 (N_2962,N_2753,N_2796);
and U2963 (N_2963,N_2763,N_2646);
and U2964 (N_2964,N_2792,N_2789);
nand U2965 (N_2965,N_2695,N_2719);
and U2966 (N_2966,N_2716,N_2698);
nor U2967 (N_2967,N_2719,N_2609);
or U2968 (N_2968,N_2667,N_2750);
nor U2969 (N_2969,N_2790,N_2641);
nand U2970 (N_2970,N_2628,N_2774);
and U2971 (N_2971,N_2693,N_2620);
nor U2972 (N_2972,N_2721,N_2775);
nor U2973 (N_2973,N_2690,N_2602);
and U2974 (N_2974,N_2690,N_2723);
nand U2975 (N_2975,N_2761,N_2703);
nor U2976 (N_2976,N_2653,N_2778);
nand U2977 (N_2977,N_2637,N_2613);
or U2978 (N_2978,N_2713,N_2778);
and U2979 (N_2979,N_2795,N_2724);
or U2980 (N_2980,N_2694,N_2621);
or U2981 (N_2981,N_2690,N_2726);
nand U2982 (N_2982,N_2673,N_2772);
xnor U2983 (N_2983,N_2606,N_2619);
nand U2984 (N_2984,N_2798,N_2791);
nand U2985 (N_2985,N_2673,N_2661);
nor U2986 (N_2986,N_2646,N_2645);
nor U2987 (N_2987,N_2748,N_2681);
and U2988 (N_2988,N_2628,N_2717);
or U2989 (N_2989,N_2792,N_2719);
or U2990 (N_2990,N_2691,N_2716);
nand U2991 (N_2991,N_2638,N_2670);
and U2992 (N_2992,N_2799,N_2685);
or U2993 (N_2993,N_2607,N_2795);
and U2994 (N_2994,N_2612,N_2781);
or U2995 (N_2995,N_2666,N_2678);
nand U2996 (N_2996,N_2716,N_2632);
or U2997 (N_2997,N_2708,N_2640);
nor U2998 (N_2998,N_2637,N_2644);
and U2999 (N_2999,N_2767,N_2742);
nand U3000 (N_3000,N_2989,N_2923);
and U3001 (N_3001,N_2850,N_2926);
and U3002 (N_3002,N_2965,N_2939);
xor U3003 (N_3003,N_2916,N_2909);
xnor U3004 (N_3004,N_2897,N_2979);
nand U3005 (N_3005,N_2818,N_2996);
nand U3006 (N_3006,N_2900,N_2912);
and U3007 (N_3007,N_2822,N_2882);
and U3008 (N_3008,N_2869,N_2920);
and U3009 (N_3009,N_2870,N_2927);
and U3010 (N_3010,N_2984,N_2852);
nand U3011 (N_3011,N_2956,N_2821);
or U3012 (N_3012,N_2834,N_2857);
nand U3013 (N_3013,N_2884,N_2831);
nor U3014 (N_3014,N_2978,N_2964);
nor U3015 (N_3015,N_2854,N_2801);
nand U3016 (N_3016,N_2843,N_2995);
or U3017 (N_3017,N_2981,N_2893);
nor U3018 (N_3018,N_2890,N_2911);
xor U3019 (N_3019,N_2986,N_2875);
and U3020 (N_3020,N_2864,N_2949);
and U3021 (N_3021,N_2967,N_2840);
or U3022 (N_3022,N_2874,N_2826);
and U3023 (N_3023,N_2809,N_2837);
nor U3024 (N_3024,N_2928,N_2881);
nand U3025 (N_3025,N_2896,N_2901);
or U3026 (N_3026,N_2955,N_2952);
and U3027 (N_3027,N_2867,N_2971);
nor U3028 (N_3028,N_2905,N_2962);
nand U3029 (N_3029,N_2929,N_2877);
and U3030 (N_3030,N_2853,N_2904);
nand U3031 (N_3031,N_2985,N_2816);
nor U3032 (N_3032,N_2812,N_2950);
nor U3033 (N_3033,N_2942,N_2963);
and U3034 (N_3034,N_2915,N_2876);
or U3035 (N_3035,N_2806,N_2935);
nand U3036 (N_3036,N_2800,N_2974);
or U3037 (N_3037,N_2810,N_2941);
and U3038 (N_3038,N_2878,N_2879);
nand U3039 (N_3039,N_2990,N_2888);
and U3040 (N_3040,N_2991,N_2841);
and U3041 (N_3041,N_2815,N_2824);
nand U3042 (N_3042,N_2980,N_2885);
nor U3043 (N_3043,N_2998,N_2883);
or U3044 (N_3044,N_2859,N_2871);
and U3045 (N_3045,N_2865,N_2866);
or U3046 (N_3046,N_2898,N_2993);
nor U3047 (N_3047,N_2994,N_2861);
or U3048 (N_3048,N_2903,N_2936);
nand U3049 (N_3049,N_2940,N_2913);
or U3050 (N_3050,N_2892,N_2947);
or U3051 (N_3051,N_2959,N_2906);
or U3052 (N_3052,N_2975,N_2988);
nor U3053 (N_3053,N_2839,N_2842);
and U3054 (N_3054,N_2804,N_2899);
nand U3055 (N_3055,N_2891,N_2972);
or U3056 (N_3056,N_2830,N_2860);
or U3057 (N_3057,N_2945,N_2807);
nor U3058 (N_3058,N_2820,N_2895);
and U3059 (N_3059,N_2808,N_2880);
nand U3060 (N_3060,N_2937,N_2973);
and U3061 (N_3061,N_2919,N_2961);
or U3062 (N_3062,N_2846,N_2908);
nand U3063 (N_3063,N_2873,N_2838);
or U3064 (N_3064,N_2953,N_2970);
nand U3065 (N_3065,N_2907,N_2946);
and U3066 (N_3066,N_2856,N_2933);
nand U3067 (N_3067,N_2827,N_2954);
or U3068 (N_3068,N_2983,N_2997);
and U3069 (N_3069,N_2805,N_2958);
or U3070 (N_3070,N_2847,N_2960);
or U3071 (N_3071,N_2894,N_2811);
or U3072 (N_3072,N_2833,N_2951);
or U3073 (N_3073,N_2817,N_2930);
nor U3074 (N_3074,N_2931,N_2976);
nor U3075 (N_3075,N_2813,N_2855);
nor U3076 (N_3076,N_2814,N_2948);
or U3077 (N_3077,N_2872,N_2966);
nand U3078 (N_3078,N_2823,N_2914);
or U3079 (N_3079,N_2977,N_2858);
nand U3080 (N_3080,N_2922,N_2849);
or U3081 (N_3081,N_2802,N_2863);
or U3082 (N_3082,N_2944,N_2918);
and U3083 (N_3083,N_2845,N_2987);
or U3084 (N_3084,N_2921,N_2982);
xnor U3085 (N_3085,N_2925,N_2957);
nand U3086 (N_3086,N_2992,N_2969);
nand U3087 (N_3087,N_2848,N_2999);
and U3088 (N_3088,N_2910,N_2887);
or U3089 (N_3089,N_2938,N_2932);
nor U3090 (N_3090,N_2902,N_2868);
nand U3091 (N_3091,N_2828,N_2819);
nand U3092 (N_3092,N_2862,N_2934);
and U3093 (N_3093,N_2832,N_2829);
and U3094 (N_3094,N_2835,N_2844);
or U3095 (N_3095,N_2917,N_2943);
or U3096 (N_3096,N_2886,N_2851);
and U3097 (N_3097,N_2889,N_2825);
and U3098 (N_3098,N_2968,N_2803);
and U3099 (N_3099,N_2924,N_2836);
or U3100 (N_3100,N_2941,N_2914);
or U3101 (N_3101,N_2812,N_2959);
or U3102 (N_3102,N_2858,N_2902);
nor U3103 (N_3103,N_2853,N_2833);
nand U3104 (N_3104,N_2874,N_2994);
and U3105 (N_3105,N_2936,N_2821);
nor U3106 (N_3106,N_2939,N_2856);
nand U3107 (N_3107,N_2852,N_2908);
and U3108 (N_3108,N_2854,N_2816);
nor U3109 (N_3109,N_2840,N_2941);
and U3110 (N_3110,N_2967,N_2958);
nand U3111 (N_3111,N_2912,N_2835);
nand U3112 (N_3112,N_2930,N_2996);
nand U3113 (N_3113,N_2885,N_2970);
and U3114 (N_3114,N_2824,N_2933);
nand U3115 (N_3115,N_2812,N_2981);
nand U3116 (N_3116,N_2980,N_2928);
nand U3117 (N_3117,N_2846,N_2928);
nand U3118 (N_3118,N_2913,N_2996);
and U3119 (N_3119,N_2856,N_2929);
or U3120 (N_3120,N_2904,N_2831);
and U3121 (N_3121,N_2847,N_2979);
or U3122 (N_3122,N_2842,N_2853);
or U3123 (N_3123,N_2837,N_2804);
nand U3124 (N_3124,N_2899,N_2949);
and U3125 (N_3125,N_2860,N_2937);
or U3126 (N_3126,N_2936,N_2984);
nand U3127 (N_3127,N_2852,N_2964);
and U3128 (N_3128,N_2884,N_2999);
and U3129 (N_3129,N_2988,N_2818);
nor U3130 (N_3130,N_2991,N_2809);
and U3131 (N_3131,N_2895,N_2961);
nor U3132 (N_3132,N_2901,N_2835);
nor U3133 (N_3133,N_2859,N_2995);
and U3134 (N_3134,N_2880,N_2911);
or U3135 (N_3135,N_2926,N_2813);
nor U3136 (N_3136,N_2969,N_2967);
and U3137 (N_3137,N_2883,N_2940);
and U3138 (N_3138,N_2948,N_2888);
nor U3139 (N_3139,N_2854,N_2977);
and U3140 (N_3140,N_2926,N_2862);
and U3141 (N_3141,N_2882,N_2886);
and U3142 (N_3142,N_2934,N_2960);
or U3143 (N_3143,N_2823,N_2822);
nand U3144 (N_3144,N_2968,N_2917);
or U3145 (N_3145,N_2927,N_2858);
nand U3146 (N_3146,N_2902,N_2907);
or U3147 (N_3147,N_2863,N_2852);
and U3148 (N_3148,N_2946,N_2877);
and U3149 (N_3149,N_2805,N_2912);
and U3150 (N_3150,N_2843,N_2808);
or U3151 (N_3151,N_2916,N_2903);
nand U3152 (N_3152,N_2982,N_2873);
or U3153 (N_3153,N_2889,N_2814);
nand U3154 (N_3154,N_2911,N_2919);
and U3155 (N_3155,N_2953,N_2825);
and U3156 (N_3156,N_2924,N_2928);
nand U3157 (N_3157,N_2848,N_2880);
and U3158 (N_3158,N_2953,N_2888);
and U3159 (N_3159,N_2821,N_2945);
nor U3160 (N_3160,N_2871,N_2826);
nor U3161 (N_3161,N_2950,N_2923);
and U3162 (N_3162,N_2872,N_2979);
nor U3163 (N_3163,N_2997,N_2995);
and U3164 (N_3164,N_2938,N_2879);
nor U3165 (N_3165,N_2850,N_2976);
xor U3166 (N_3166,N_2906,N_2981);
or U3167 (N_3167,N_2848,N_2850);
nand U3168 (N_3168,N_2833,N_2924);
and U3169 (N_3169,N_2968,N_2800);
nand U3170 (N_3170,N_2943,N_2816);
nand U3171 (N_3171,N_2883,N_2824);
xor U3172 (N_3172,N_2890,N_2946);
or U3173 (N_3173,N_2933,N_2910);
nand U3174 (N_3174,N_2819,N_2948);
nand U3175 (N_3175,N_2913,N_2952);
nor U3176 (N_3176,N_2991,N_2808);
and U3177 (N_3177,N_2830,N_2977);
and U3178 (N_3178,N_2995,N_2802);
nand U3179 (N_3179,N_2996,N_2951);
or U3180 (N_3180,N_2898,N_2864);
or U3181 (N_3181,N_2952,N_2972);
or U3182 (N_3182,N_2879,N_2902);
or U3183 (N_3183,N_2917,N_2920);
and U3184 (N_3184,N_2929,N_2903);
nand U3185 (N_3185,N_2883,N_2984);
nor U3186 (N_3186,N_2945,N_2837);
and U3187 (N_3187,N_2866,N_2804);
and U3188 (N_3188,N_2921,N_2810);
or U3189 (N_3189,N_2894,N_2945);
nand U3190 (N_3190,N_2931,N_2968);
nor U3191 (N_3191,N_2934,N_2825);
nand U3192 (N_3192,N_2850,N_2888);
nand U3193 (N_3193,N_2918,N_2815);
nor U3194 (N_3194,N_2985,N_2862);
nor U3195 (N_3195,N_2806,N_2999);
nor U3196 (N_3196,N_2829,N_2875);
and U3197 (N_3197,N_2908,N_2988);
xor U3198 (N_3198,N_2859,N_2963);
or U3199 (N_3199,N_2998,N_2922);
or U3200 (N_3200,N_3026,N_3175);
or U3201 (N_3201,N_3024,N_3031);
or U3202 (N_3202,N_3115,N_3157);
nor U3203 (N_3203,N_3192,N_3150);
nor U3204 (N_3204,N_3112,N_3134);
or U3205 (N_3205,N_3130,N_3057);
and U3206 (N_3206,N_3091,N_3077);
nor U3207 (N_3207,N_3189,N_3123);
nor U3208 (N_3208,N_3119,N_3173);
or U3209 (N_3209,N_3045,N_3059);
nand U3210 (N_3210,N_3147,N_3195);
xor U3211 (N_3211,N_3097,N_3078);
and U3212 (N_3212,N_3073,N_3060);
nor U3213 (N_3213,N_3050,N_3144);
or U3214 (N_3214,N_3108,N_3135);
nor U3215 (N_3215,N_3141,N_3171);
nand U3216 (N_3216,N_3027,N_3064);
nand U3217 (N_3217,N_3166,N_3092);
or U3218 (N_3218,N_3133,N_3098);
nor U3219 (N_3219,N_3096,N_3025);
nor U3220 (N_3220,N_3075,N_3034);
nor U3221 (N_3221,N_3004,N_3158);
and U3222 (N_3222,N_3087,N_3020);
nor U3223 (N_3223,N_3088,N_3156);
nor U3224 (N_3224,N_3053,N_3137);
nand U3225 (N_3225,N_3120,N_3164);
or U3226 (N_3226,N_3048,N_3022);
and U3227 (N_3227,N_3183,N_3043);
and U3228 (N_3228,N_3013,N_3070);
nand U3229 (N_3229,N_3111,N_3149);
and U3230 (N_3230,N_3003,N_3121);
or U3231 (N_3231,N_3186,N_3107);
or U3232 (N_3232,N_3029,N_3145);
nor U3233 (N_3233,N_3032,N_3066);
or U3234 (N_3234,N_3076,N_3058);
nand U3235 (N_3235,N_3069,N_3193);
nor U3236 (N_3236,N_3198,N_3063);
nor U3237 (N_3237,N_3178,N_3170);
nand U3238 (N_3238,N_3041,N_3104);
nor U3239 (N_3239,N_3113,N_3179);
nor U3240 (N_3240,N_3190,N_3046);
and U3241 (N_3241,N_3172,N_3000);
and U3242 (N_3242,N_3129,N_3062);
or U3243 (N_3243,N_3008,N_3160);
and U3244 (N_3244,N_3090,N_3083);
nor U3245 (N_3245,N_3094,N_3188);
nand U3246 (N_3246,N_3176,N_3159);
nand U3247 (N_3247,N_3184,N_3122);
nand U3248 (N_3248,N_3197,N_3127);
nor U3249 (N_3249,N_3015,N_3044);
nand U3250 (N_3250,N_3177,N_3124);
or U3251 (N_3251,N_3061,N_3072);
and U3252 (N_3252,N_3047,N_3152);
nand U3253 (N_3253,N_3131,N_3039);
nand U3254 (N_3254,N_3011,N_3030);
or U3255 (N_3255,N_3082,N_3017);
or U3256 (N_3256,N_3146,N_3038);
nor U3257 (N_3257,N_3002,N_3110);
and U3258 (N_3258,N_3084,N_3071);
nand U3259 (N_3259,N_3035,N_3036);
nand U3260 (N_3260,N_3165,N_3067);
and U3261 (N_3261,N_3128,N_3142);
or U3262 (N_3262,N_3140,N_3099);
nand U3263 (N_3263,N_3089,N_3016);
or U3264 (N_3264,N_3182,N_3052);
nor U3265 (N_3265,N_3180,N_3021);
or U3266 (N_3266,N_3185,N_3101);
or U3267 (N_3267,N_3106,N_3116);
and U3268 (N_3268,N_3074,N_3153);
or U3269 (N_3269,N_3079,N_3138);
or U3270 (N_3270,N_3005,N_3065);
or U3271 (N_3271,N_3161,N_3191);
and U3272 (N_3272,N_3136,N_3095);
and U3273 (N_3273,N_3109,N_3196);
or U3274 (N_3274,N_3174,N_3114);
nand U3275 (N_3275,N_3023,N_3118);
and U3276 (N_3276,N_3055,N_3194);
and U3277 (N_3277,N_3100,N_3162);
or U3278 (N_3278,N_3010,N_3006);
or U3279 (N_3279,N_3154,N_3051);
or U3280 (N_3280,N_3014,N_3169);
or U3281 (N_3281,N_3163,N_3148);
nand U3282 (N_3282,N_3103,N_3187);
nor U3283 (N_3283,N_3001,N_3081);
nor U3284 (N_3284,N_3012,N_3085);
or U3285 (N_3285,N_3037,N_3125);
and U3286 (N_3286,N_3139,N_3080);
nand U3287 (N_3287,N_3068,N_3018);
nand U3288 (N_3288,N_3105,N_3019);
nand U3289 (N_3289,N_3132,N_3126);
nand U3290 (N_3290,N_3007,N_3151);
nand U3291 (N_3291,N_3033,N_3056);
or U3292 (N_3292,N_3028,N_3199);
nor U3293 (N_3293,N_3086,N_3042);
nor U3294 (N_3294,N_3143,N_3117);
nor U3295 (N_3295,N_3009,N_3155);
and U3296 (N_3296,N_3040,N_3181);
or U3297 (N_3297,N_3093,N_3168);
nand U3298 (N_3298,N_3167,N_3049);
nor U3299 (N_3299,N_3102,N_3054);
and U3300 (N_3300,N_3103,N_3194);
or U3301 (N_3301,N_3084,N_3125);
and U3302 (N_3302,N_3059,N_3172);
and U3303 (N_3303,N_3107,N_3124);
nand U3304 (N_3304,N_3002,N_3019);
and U3305 (N_3305,N_3165,N_3104);
and U3306 (N_3306,N_3107,N_3007);
and U3307 (N_3307,N_3163,N_3075);
nand U3308 (N_3308,N_3027,N_3120);
or U3309 (N_3309,N_3108,N_3025);
nor U3310 (N_3310,N_3169,N_3064);
and U3311 (N_3311,N_3163,N_3055);
nor U3312 (N_3312,N_3029,N_3189);
and U3313 (N_3313,N_3045,N_3049);
nor U3314 (N_3314,N_3099,N_3193);
or U3315 (N_3315,N_3129,N_3189);
or U3316 (N_3316,N_3181,N_3131);
nor U3317 (N_3317,N_3153,N_3000);
nand U3318 (N_3318,N_3122,N_3192);
and U3319 (N_3319,N_3071,N_3048);
or U3320 (N_3320,N_3199,N_3165);
nor U3321 (N_3321,N_3151,N_3053);
nand U3322 (N_3322,N_3188,N_3169);
and U3323 (N_3323,N_3106,N_3104);
or U3324 (N_3324,N_3181,N_3103);
and U3325 (N_3325,N_3049,N_3171);
nor U3326 (N_3326,N_3121,N_3059);
nor U3327 (N_3327,N_3111,N_3196);
xor U3328 (N_3328,N_3096,N_3135);
nand U3329 (N_3329,N_3143,N_3193);
or U3330 (N_3330,N_3194,N_3182);
nand U3331 (N_3331,N_3011,N_3055);
or U3332 (N_3332,N_3038,N_3075);
and U3333 (N_3333,N_3004,N_3143);
or U3334 (N_3334,N_3154,N_3069);
nor U3335 (N_3335,N_3015,N_3066);
and U3336 (N_3336,N_3116,N_3166);
or U3337 (N_3337,N_3014,N_3050);
nor U3338 (N_3338,N_3160,N_3053);
nor U3339 (N_3339,N_3187,N_3076);
nor U3340 (N_3340,N_3193,N_3168);
nor U3341 (N_3341,N_3113,N_3029);
nor U3342 (N_3342,N_3124,N_3171);
nand U3343 (N_3343,N_3046,N_3199);
nand U3344 (N_3344,N_3027,N_3046);
nor U3345 (N_3345,N_3188,N_3168);
or U3346 (N_3346,N_3140,N_3044);
and U3347 (N_3347,N_3158,N_3000);
or U3348 (N_3348,N_3036,N_3098);
nand U3349 (N_3349,N_3021,N_3141);
nand U3350 (N_3350,N_3157,N_3144);
and U3351 (N_3351,N_3045,N_3082);
nor U3352 (N_3352,N_3013,N_3127);
or U3353 (N_3353,N_3015,N_3148);
and U3354 (N_3354,N_3110,N_3103);
and U3355 (N_3355,N_3081,N_3010);
or U3356 (N_3356,N_3089,N_3125);
and U3357 (N_3357,N_3179,N_3166);
and U3358 (N_3358,N_3180,N_3122);
nor U3359 (N_3359,N_3093,N_3115);
nand U3360 (N_3360,N_3181,N_3167);
nand U3361 (N_3361,N_3028,N_3070);
nand U3362 (N_3362,N_3170,N_3108);
nor U3363 (N_3363,N_3055,N_3076);
nor U3364 (N_3364,N_3114,N_3000);
or U3365 (N_3365,N_3176,N_3131);
nor U3366 (N_3366,N_3019,N_3123);
nand U3367 (N_3367,N_3072,N_3069);
nor U3368 (N_3368,N_3172,N_3125);
or U3369 (N_3369,N_3130,N_3175);
and U3370 (N_3370,N_3070,N_3153);
nand U3371 (N_3371,N_3065,N_3028);
xor U3372 (N_3372,N_3057,N_3038);
or U3373 (N_3373,N_3113,N_3128);
nand U3374 (N_3374,N_3199,N_3191);
or U3375 (N_3375,N_3130,N_3172);
nor U3376 (N_3376,N_3055,N_3110);
or U3377 (N_3377,N_3010,N_3140);
nand U3378 (N_3378,N_3181,N_3025);
nor U3379 (N_3379,N_3015,N_3029);
and U3380 (N_3380,N_3092,N_3002);
and U3381 (N_3381,N_3121,N_3019);
and U3382 (N_3382,N_3153,N_3043);
or U3383 (N_3383,N_3177,N_3123);
and U3384 (N_3384,N_3147,N_3159);
nor U3385 (N_3385,N_3047,N_3082);
nand U3386 (N_3386,N_3102,N_3111);
nor U3387 (N_3387,N_3087,N_3113);
or U3388 (N_3388,N_3047,N_3101);
nand U3389 (N_3389,N_3091,N_3111);
or U3390 (N_3390,N_3087,N_3013);
nor U3391 (N_3391,N_3115,N_3152);
or U3392 (N_3392,N_3084,N_3099);
or U3393 (N_3393,N_3038,N_3130);
nor U3394 (N_3394,N_3196,N_3017);
or U3395 (N_3395,N_3129,N_3039);
or U3396 (N_3396,N_3113,N_3047);
and U3397 (N_3397,N_3172,N_3154);
xor U3398 (N_3398,N_3079,N_3011);
nand U3399 (N_3399,N_3191,N_3175);
nand U3400 (N_3400,N_3397,N_3312);
and U3401 (N_3401,N_3306,N_3236);
nand U3402 (N_3402,N_3321,N_3304);
or U3403 (N_3403,N_3200,N_3245);
nand U3404 (N_3404,N_3316,N_3359);
nand U3405 (N_3405,N_3299,N_3264);
nor U3406 (N_3406,N_3287,N_3297);
nand U3407 (N_3407,N_3239,N_3229);
or U3408 (N_3408,N_3203,N_3225);
nand U3409 (N_3409,N_3231,N_3249);
nand U3410 (N_3410,N_3283,N_3221);
and U3411 (N_3411,N_3372,N_3387);
nor U3412 (N_3412,N_3346,N_3320);
and U3413 (N_3413,N_3218,N_3232);
nor U3414 (N_3414,N_3250,N_3235);
and U3415 (N_3415,N_3282,N_3237);
nor U3416 (N_3416,N_3205,N_3340);
nand U3417 (N_3417,N_3277,N_3391);
nor U3418 (N_3418,N_3275,N_3220);
and U3419 (N_3419,N_3389,N_3271);
and U3420 (N_3420,N_3222,N_3351);
or U3421 (N_3421,N_3366,N_3255);
and U3422 (N_3422,N_3303,N_3284);
nor U3423 (N_3423,N_3367,N_3352);
or U3424 (N_3424,N_3311,N_3327);
xnor U3425 (N_3425,N_3214,N_3382);
and U3426 (N_3426,N_3319,N_3357);
nand U3427 (N_3427,N_3383,N_3212);
nand U3428 (N_3428,N_3385,N_3226);
or U3429 (N_3429,N_3305,N_3337);
and U3430 (N_3430,N_3213,N_3301);
nand U3431 (N_3431,N_3268,N_3396);
nor U3432 (N_3432,N_3234,N_3330);
or U3433 (N_3433,N_3228,N_3251);
and U3434 (N_3434,N_3238,N_3261);
or U3435 (N_3435,N_3329,N_3292);
and U3436 (N_3436,N_3210,N_3368);
and U3437 (N_3437,N_3376,N_3267);
or U3438 (N_3438,N_3332,N_3286);
and U3439 (N_3439,N_3298,N_3375);
or U3440 (N_3440,N_3243,N_3215);
nor U3441 (N_3441,N_3230,N_3296);
nor U3442 (N_3442,N_3333,N_3354);
nand U3443 (N_3443,N_3342,N_3328);
or U3444 (N_3444,N_3241,N_3269);
or U3445 (N_3445,N_3364,N_3219);
nand U3446 (N_3446,N_3361,N_3302);
xnor U3447 (N_3447,N_3349,N_3390);
nand U3448 (N_3448,N_3207,N_3223);
and U3449 (N_3449,N_3276,N_3347);
or U3450 (N_3450,N_3317,N_3209);
or U3451 (N_3451,N_3370,N_3386);
xor U3452 (N_3452,N_3323,N_3378);
or U3453 (N_3453,N_3285,N_3363);
nand U3454 (N_3454,N_3392,N_3227);
nor U3455 (N_3455,N_3308,N_3211);
nand U3456 (N_3456,N_3374,N_3379);
nor U3457 (N_3457,N_3345,N_3233);
nand U3458 (N_3458,N_3315,N_3256);
nor U3459 (N_3459,N_3270,N_3338);
nand U3460 (N_3460,N_3300,N_3377);
nand U3461 (N_3461,N_3313,N_3381);
xnor U3462 (N_3462,N_3278,N_3395);
nor U3463 (N_3463,N_3365,N_3388);
nand U3464 (N_3464,N_3310,N_3260);
nor U3465 (N_3465,N_3380,N_3336);
and U3466 (N_3466,N_3280,N_3294);
nand U3467 (N_3467,N_3398,N_3208);
nor U3468 (N_3468,N_3259,N_3295);
and U3469 (N_3469,N_3242,N_3355);
and U3470 (N_3470,N_3348,N_3263);
nor U3471 (N_3471,N_3202,N_3353);
and U3472 (N_3472,N_3322,N_3265);
and U3473 (N_3473,N_3343,N_3371);
and U3474 (N_3474,N_3216,N_3324);
or U3475 (N_3475,N_3360,N_3358);
nor U3476 (N_3476,N_3335,N_3266);
nand U3477 (N_3477,N_3253,N_3362);
or U3478 (N_3478,N_3217,N_3394);
or U3479 (N_3479,N_3279,N_3262);
nor U3480 (N_3480,N_3399,N_3204);
nand U3481 (N_3481,N_3272,N_3244);
nor U3482 (N_3482,N_3293,N_3318);
or U3483 (N_3483,N_3254,N_3350);
nand U3484 (N_3484,N_3289,N_3288);
or U3485 (N_3485,N_3326,N_3334);
nand U3486 (N_3486,N_3281,N_3240);
nand U3487 (N_3487,N_3274,N_3344);
or U3488 (N_3488,N_3248,N_3201);
nand U3489 (N_3489,N_3369,N_3307);
nand U3490 (N_3490,N_3291,N_3252);
or U3491 (N_3491,N_3339,N_3247);
nor U3492 (N_3492,N_3325,N_3257);
and U3493 (N_3493,N_3373,N_3258);
nand U3494 (N_3494,N_3384,N_3246);
or U3495 (N_3495,N_3341,N_3331);
nor U3496 (N_3496,N_3206,N_3393);
and U3497 (N_3497,N_3314,N_3309);
nand U3498 (N_3498,N_3356,N_3290);
xnor U3499 (N_3499,N_3224,N_3273);
and U3500 (N_3500,N_3299,N_3342);
and U3501 (N_3501,N_3315,N_3342);
nor U3502 (N_3502,N_3352,N_3265);
or U3503 (N_3503,N_3319,N_3385);
nand U3504 (N_3504,N_3319,N_3382);
or U3505 (N_3505,N_3338,N_3229);
and U3506 (N_3506,N_3352,N_3259);
and U3507 (N_3507,N_3394,N_3291);
nand U3508 (N_3508,N_3251,N_3365);
or U3509 (N_3509,N_3350,N_3204);
nand U3510 (N_3510,N_3209,N_3354);
nor U3511 (N_3511,N_3240,N_3278);
nand U3512 (N_3512,N_3289,N_3303);
nand U3513 (N_3513,N_3246,N_3249);
nand U3514 (N_3514,N_3275,N_3228);
xnor U3515 (N_3515,N_3246,N_3369);
nand U3516 (N_3516,N_3294,N_3389);
and U3517 (N_3517,N_3350,N_3209);
and U3518 (N_3518,N_3344,N_3247);
and U3519 (N_3519,N_3380,N_3238);
nor U3520 (N_3520,N_3312,N_3395);
and U3521 (N_3521,N_3369,N_3383);
nand U3522 (N_3522,N_3310,N_3315);
and U3523 (N_3523,N_3396,N_3235);
nor U3524 (N_3524,N_3377,N_3380);
or U3525 (N_3525,N_3310,N_3283);
nor U3526 (N_3526,N_3318,N_3264);
or U3527 (N_3527,N_3276,N_3289);
nor U3528 (N_3528,N_3265,N_3235);
and U3529 (N_3529,N_3288,N_3370);
nor U3530 (N_3530,N_3372,N_3308);
or U3531 (N_3531,N_3304,N_3399);
nand U3532 (N_3532,N_3352,N_3356);
or U3533 (N_3533,N_3209,N_3386);
nand U3534 (N_3534,N_3352,N_3241);
or U3535 (N_3535,N_3277,N_3386);
nor U3536 (N_3536,N_3286,N_3347);
nor U3537 (N_3537,N_3365,N_3286);
or U3538 (N_3538,N_3395,N_3353);
and U3539 (N_3539,N_3277,N_3271);
and U3540 (N_3540,N_3325,N_3236);
and U3541 (N_3541,N_3208,N_3325);
and U3542 (N_3542,N_3381,N_3205);
or U3543 (N_3543,N_3387,N_3375);
and U3544 (N_3544,N_3200,N_3379);
and U3545 (N_3545,N_3377,N_3249);
nand U3546 (N_3546,N_3302,N_3255);
and U3547 (N_3547,N_3352,N_3383);
nand U3548 (N_3548,N_3368,N_3200);
nor U3549 (N_3549,N_3285,N_3361);
nor U3550 (N_3550,N_3328,N_3327);
nand U3551 (N_3551,N_3398,N_3290);
or U3552 (N_3552,N_3231,N_3247);
nand U3553 (N_3553,N_3290,N_3220);
nand U3554 (N_3554,N_3223,N_3253);
or U3555 (N_3555,N_3283,N_3364);
or U3556 (N_3556,N_3384,N_3395);
nor U3557 (N_3557,N_3225,N_3229);
and U3558 (N_3558,N_3325,N_3227);
and U3559 (N_3559,N_3315,N_3372);
xor U3560 (N_3560,N_3373,N_3286);
and U3561 (N_3561,N_3206,N_3339);
or U3562 (N_3562,N_3257,N_3389);
and U3563 (N_3563,N_3260,N_3313);
nor U3564 (N_3564,N_3264,N_3284);
nand U3565 (N_3565,N_3280,N_3223);
nor U3566 (N_3566,N_3299,N_3209);
nand U3567 (N_3567,N_3272,N_3351);
and U3568 (N_3568,N_3210,N_3340);
nand U3569 (N_3569,N_3225,N_3287);
nor U3570 (N_3570,N_3360,N_3349);
nand U3571 (N_3571,N_3212,N_3369);
nor U3572 (N_3572,N_3267,N_3243);
and U3573 (N_3573,N_3363,N_3342);
nand U3574 (N_3574,N_3267,N_3252);
nand U3575 (N_3575,N_3352,N_3201);
and U3576 (N_3576,N_3366,N_3324);
and U3577 (N_3577,N_3255,N_3259);
xnor U3578 (N_3578,N_3351,N_3340);
nand U3579 (N_3579,N_3263,N_3352);
and U3580 (N_3580,N_3204,N_3265);
or U3581 (N_3581,N_3291,N_3302);
nor U3582 (N_3582,N_3344,N_3392);
nor U3583 (N_3583,N_3280,N_3352);
or U3584 (N_3584,N_3276,N_3293);
nor U3585 (N_3585,N_3384,N_3350);
nor U3586 (N_3586,N_3358,N_3355);
nor U3587 (N_3587,N_3281,N_3349);
nand U3588 (N_3588,N_3221,N_3386);
xnor U3589 (N_3589,N_3331,N_3374);
or U3590 (N_3590,N_3293,N_3397);
nand U3591 (N_3591,N_3200,N_3338);
nor U3592 (N_3592,N_3300,N_3362);
nor U3593 (N_3593,N_3341,N_3210);
and U3594 (N_3594,N_3364,N_3314);
nor U3595 (N_3595,N_3205,N_3233);
and U3596 (N_3596,N_3352,N_3299);
nand U3597 (N_3597,N_3370,N_3313);
nor U3598 (N_3598,N_3322,N_3344);
or U3599 (N_3599,N_3249,N_3214);
or U3600 (N_3600,N_3543,N_3567);
nand U3601 (N_3601,N_3570,N_3566);
nor U3602 (N_3602,N_3569,N_3408);
nand U3603 (N_3603,N_3534,N_3451);
nor U3604 (N_3604,N_3520,N_3470);
nor U3605 (N_3605,N_3416,N_3439);
and U3606 (N_3606,N_3498,N_3450);
and U3607 (N_3607,N_3515,N_3487);
nand U3608 (N_3608,N_3500,N_3577);
xnor U3609 (N_3609,N_3598,N_3533);
and U3610 (N_3610,N_3538,N_3406);
or U3611 (N_3611,N_3468,N_3556);
and U3612 (N_3612,N_3428,N_3529);
and U3613 (N_3613,N_3434,N_3481);
nor U3614 (N_3614,N_3443,N_3550);
nor U3615 (N_3615,N_3547,N_3463);
nand U3616 (N_3616,N_3411,N_3413);
nor U3617 (N_3617,N_3422,N_3492);
xor U3618 (N_3618,N_3525,N_3446);
nor U3619 (N_3619,N_3578,N_3561);
or U3620 (N_3620,N_3444,N_3400);
and U3621 (N_3621,N_3507,N_3549);
or U3622 (N_3622,N_3506,N_3562);
nor U3623 (N_3623,N_3404,N_3474);
and U3624 (N_3624,N_3438,N_3539);
and U3625 (N_3625,N_3403,N_3593);
and U3626 (N_3626,N_3502,N_3469);
nor U3627 (N_3627,N_3447,N_3594);
nand U3628 (N_3628,N_3558,N_3559);
and U3629 (N_3629,N_3579,N_3417);
nand U3630 (N_3630,N_3518,N_3595);
nand U3631 (N_3631,N_3541,N_3530);
or U3632 (N_3632,N_3575,N_3585);
nand U3633 (N_3633,N_3528,N_3453);
or U3634 (N_3634,N_3546,N_3401);
nand U3635 (N_3635,N_3471,N_3563);
or U3636 (N_3636,N_3418,N_3419);
and U3637 (N_3637,N_3531,N_3526);
nand U3638 (N_3638,N_3524,N_3484);
or U3639 (N_3639,N_3405,N_3425);
or U3640 (N_3640,N_3499,N_3519);
nor U3641 (N_3641,N_3496,N_3465);
and U3642 (N_3642,N_3426,N_3591);
or U3643 (N_3643,N_3449,N_3480);
nand U3644 (N_3644,N_3414,N_3574);
nor U3645 (N_3645,N_3521,N_3552);
and U3646 (N_3646,N_3435,N_3494);
nor U3647 (N_3647,N_3483,N_3564);
and U3648 (N_3648,N_3491,N_3560);
and U3649 (N_3649,N_3421,N_3420);
or U3650 (N_3650,N_3479,N_3457);
or U3651 (N_3651,N_3587,N_3581);
or U3652 (N_3652,N_3555,N_3431);
nand U3653 (N_3653,N_3544,N_3512);
nor U3654 (N_3654,N_3427,N_3407);
nand U3655 (N_3655,N_3497,N_3493);
nor U3656 (N_3656,N_3584,N_3596);
and U3657 (N_3657,N_3554,N_3462);
nor U3658 (N_3658,N_3464,N_3448);
nor U3659 (N_3659,N_3537,N_3489);
and U3660 (N_3660,N_3580,N_3430);
nor U3661 (N_3661,N_3505,N_3523);
nor U3662 (N_3662,N_3527,N_3459);
nor U3663 (N_3663,N_3410,N_3424);
nor U3664 (N_3664,N_3553,N_3514);
xnor U3665 (N_3665,N_3503,N_3516);
nand U3666 (N_3666,N_3589,N_3572);
nor U3667 (N_3667,N_3473,N_3440);
nand U3668 (N_3668,N_3540,N_3478);
and U3669 (N_3669,N_3402,N_3476);
or U3670 (N_3670,N_3573,N_3511);
nand U3671 (N_3671,N_3467,N_3441);
and U3672 (N_3672,N_3592,N_3513);
or U3673 (N_3673,N_3458,N_3454);
and U3674 (N_3674,N_3442,N_3535);
or U3675 (N_3675,N_3485,N_3588);
and U3676 (N_3676,N_3460,N_3490);
nand U3677 (N_3677,N_3504,N_3522);
nor U3678 (N_3678,N_3495,N_3583);
nor U3679 (N_3679,N_3445,N_3461);
or U3680 (N_3680,N_3517,N_3590);
or U3681 (N_3681,N_3423,N_3437);
or U3682 (N_3682,N_3409,N_3557);
nor U3683 (N_3683,N_3433,N_3571);
or U3684 (N_3684,N_3486,N_3475);
and U3685 (N_3685,N_3582,N_3510);
or U3686 (N_3686,N_3532,N_3536);
nor U3687 (N_3687,N_3432,N_3508);
and U3688 (N_3688,N_3452,N_3456);
and U3689 (N_3689,N_3576,N_3548);
xnor U3690 (N_3690,N_3415,N_3545);
and U3691 (N_3691,N_3482,N_3586);
xnor U3692 (N_3692,N_3412,N_3565);
nand U3693 (N_3693,N_3568,N_3472);
nand U3694 (N_3694,N_3429,N_3599);
nor U3695 (N_3695,N_3466,N_3436);
or U3696 (N_3696,N_3455,N_3551);
or U3697 (N_3697,N_3477,N_3509);
xnor U3698 (N_3698,N_3488,N_3597);
nor U3699 (N_3699,N_3542,N_3501);
nand U3700 (N_3700,N_3439,N_3515);
and U3701 (N_3701,N_3464,N_3488);
nand U3702 (N_3702,N_3441,N_3409);
nand U3703 (N_3703,N_3568,N_3571);
and U3704 (N_3704,N_3584,N_3500);
or U3705 (N_3705,N_3536,N_3599);
nor U3706 (N_3706,N_3496,N_3490);
or U3707 (N_3707,N_3532,N_3554);
nand U3708 (N_3708,N_3577,N_3542);
nand U3709 (N_3709,N_3596,N_3503);
nand U3710 (N_3710,N_3511,N_3571);
nor U3711 (N_3711,N_3551,N_3518);
and U3712 (N_3712,N_3502,N_3518);
nand U3713 (N_3713,N_3507,N_3455);
or U3714 (N_3714,N_3414,N_3424);
xor U3715 (N_3715,N_3534,N_3462);
or U3716 (N_3716,N_3431,N_3556);
or U3717 (N_3717,N_3526,N_3485);
nand U3718 (N_3718,N_3502,N_3444);
xor U3719 (N_3719,N_3588,N_3484);
and U3720 (N_3720,N_3585,N_3503);
and U3721 (N_3721,N_3567,N_3434);
and U3722 (N_3722,N_3562,N_3453);
or U3723 (N_3723,N_3412,N_3406);
nand U3724 (N_3724,N_3598,N_3410);
or U3725 (N_3725,N_3401,N_3407);
or U3726 (N_3726,N_3519,N_3456);
or U3727 (N_3727,N_3499,N_3532);
nand U3728 (N_3728,N_3522,N_3578);
nand U3729 (N_3729,N_3498,N_3405);
or U3730 (N_3730,N_3509,N_3565);
or U3731 (N_3731,N_3443,N_3457);
nor U3732 (N_3732,N_3589,N_3517);
and U3733 (N_3733,N_3569,N_3557);
or U3734 (N_3734,N_3542,N_3586);
nand U3735 (N_3735,N_3584,N_3557);
and U3736 (N_3736,N_3573,N_3482);
and U3737 (N_3737,N_3514,N_3570);
nor U3738 (N_3738,N_3404,N_3464);
and U3739 (N_3739,N_3460,N_3405);
nor U3740 (N_3740,N_3447,N_3437);
nor U3741 (N_3741,N_3575,N_3439);
or U3742 (N_3742,N_3499,N_3527);
and U3743 (N_3743,N_3492,N_3534);
xor U3744 (N_3744,N_3562,N_3459);
nand U3745 (N_3745,N_3470,N_3404);
nor U3746 (N_3746,N_3576,N_3478);
nand U3747 (N_3747,N_3497,N_3577);
nand U3748 (N_3748,N_3534,N_3527);
or U3749 (N_3749,N_3553,N_3426);
or U3750 (N_3750,N_3561,N_3410);
nand U3751 (N_3751,N_3409,N_3566);
or U3752 (N_3752,N_3508,N_3574);
nand U3753 (N_3753,N_3479,N_3552);
nand U3754 (N_3754,N_3511,N_3520);
or U3755 (N_3755,N_3544,N_3571);
and U3756 (N_3756,N_3412,N_3495);
or U3757 (N_3757,N_3597,N_3428);
xnor U3758 (N_3758,N_3516,N_3426);
or U3759 (N_3759,N_3594,N_3498);
or U3760 (N_3760,N_3517,N_3485);
nand U3761 (N_3761,N_3484,N_3478);
and U3762 (N_3762,N_3520,N_3522);
or U3763 (N_3763,N_3492,N_3488);
nand U3764 (N_3764,N_3536,N_3443);
nand U3765 (N_3765,N_3541,N_3574);
nor U3766 (N_3766,N_3508,N_3596);
nor U3767 (N_3767,N_3438,N_3515);
and U3768 (N_3768,N_3501,N_3526);
and U3769 (N_3769,N_3591,N_3453);
nand U3770 (N_3770,N_3581,N_3474);
nor U3771 (N_3771,N_3485,N_3496);
and U3772 (N_3772,N_3547,N_3428);
and U3773 (N_3773,N_3574,N_3576);
or U3774 (N_3774,N_3452,N_3441);
nor U3775 (N_3775,N_3538,N_3488);
or U3776 (N_3776,N_3530,N_3465);
nand U3777 (N_3777,N_3411,N_3526);
nor U3778 (N_3778,N_3459,N_3412);
nand U3779 (N_3779,N_3408,N_3417);
nand U3780 (N_3780,N_3528,N_3510);
and U3781 (N_3781,N_3550,N_3410);
and U3782 (N_3782,N_3400,N_3556);
and U3783 (N_3783,N_3594,N_3507);
nand U3784 (N_3784,N_3546,N_3437);
nor U3785 (N_3785,N_3439,N_3440);
and U3786 (N_3786,N_3520,N_3563);
or U3787 (N_3787,N_3578,N_3533);
nand U3788 (N_3788,N_3557,N_3488);
and U3789 (N_3789,N_3506,N_3520);
or U3790 (N_3790,N_3501,N_3476);
nand U3791 (N_3791,N_3478,N_3422);
nand U3792 (N_3792,N_3561,N_3486);
and U3793 (N_3793,N_3525,N_3542);
nor U3794 (N_3794,N_3496,N_3403);
and U3795 (N_3795,N_3513,N_3594);
and U3796 (N_3796,N_3458,N_3533);
or U3797 (N_3797,N_3442,N_3589);
and U3798 (N_3798,N_3571,N_3586);
nand U3799 (N_3799,N_3519,N_3594);
nand U3800 (N_3800,N_3758,N_3761);
or U3801 (N_3801,N_3642,N_3680);
or U3802 (N_3802,N_3753,N_3685);
nand U3803 (N_3803,N_3683,N_3713);
or U3804 (N_3804,N_3626,N_3718);
nor U3805 (N_3805,N_3651,N_3676);
nor U3806 (N_3806,N_3677,N_3799);
xor U3807 (N_3807,N_3791,N_3716);
xnor U3808 (N_3808,N_3625,N_3729);
or U3809 (N_3809,N_3702,N_3619);
and U3810 (N_3810,N_3738,N_3707);
or U3811 (N_3811,N_3719,N_3645);
and U3812 (N_3812,N_3755,N_3790);
nand U3813 (N_3813,N_3709,N_3605);
nor U3814 (N_3814,N_3728,N_3665);
or U3815 (N_3815,N_3650,N_3623);
nor U3816 (N_3816,N_3724,N_3774);
nand U3817 (N_3817,N_3644,N_3693);
or U3818 (N_3818,N_3796,N_3710);
or U3819 (N_3819,N_3786,N_3788);
or U3820 (N_3820,N_3773,N_3727);
nor U3821 (N_3821,N_3778,N_3754);
or U3822 (N_3822,N_3798,N_3620);
nand U3823 (N_3823,N_3614,N_3771);
nand U3824 (N_3824,N_3632,N_3692);
or U3825 (N_3825,N_3723,N_3787);
and U3826 (N_3826,N_3684,N_3782);
or U3827 (N_3827,N_3612,N_3637);
nand U3828 (N_3828,N_3671,N_3734);
and U3829 (N_3829,N_3793,N_3781);
and U3830 (N_3830,N_3797,N_3775);
or U3831 (N_3831,N_3664,N_3674);
nor U3832 (N_3832,N_3682,N_3646);
and U3833 (N_3833,N_3748,N_3624);
or U3834 (N_3834,N_3675,N_3667);
or U3835 (N_3835,N_3760,N_3627);
nor U3836 (N_3836,N_3759,N_3631);
and U3837 (N_3837,N_3725,N_3634);
or U3838 (N_3838,N_3757,N_3750);
nor U3839 (N_3839,N_3648,N_3743);
and U3840 (N_3840,N_3714,N_3705);
nand U3841 (N_3841,N_3764,N_3601);
nand U3842 (N_3842,N_3639,N_3732);
nand U3843 (N_3843,N_3766,N_3741);
nand U3844 (N_3844,N_3770,N_3657);
and U3845 (N_3845,N_3795,N_3706);
nor U3846 (N_3846,N_3621,N_3762);
and U3847 (N_3847,N_3733,N_3660);
xnor U3848 (N_3848,N_3687,N_3703);
and U3849 (N_3849,N_3647,N_3744);
nand U3850 (N_3850,N_3780,N_3628);
nor U3851 (N_3851,N_3611,N_3737);
and U3852 (N_3852,N_3661,N_3658);
xnor U3853 (N_3853,N_3765,N_3721);
or U3854 (N_3854,N_3603,N_3740);
nand U3855 (N_3855,N_3698,N_3777);
nor U3856 (N_3856,N_3615,N_3767);
or U3857 (N_3857,N_3756,N_3636);
and U3858 (N_3858,N_3630,N_3794);
or U3859 (N_3859,N_3688,N_3700);
xor U3860 (N_3860,N_3742,N_3768);
or U3861 (N_3861,N_3679,N_3662);
and U3862 (N_3862,N_3697,N_3708);
and U3863 (N_3863,N_3752,N_3776);
or U3864 (N_3864,N_3669,N_3600);
or U3865 (N_3865,N_3613,N_3722);
or U3866 (N_3866,N_3701,N_3638);
and U3867 (N_3867,N_3704,N_3720);
and U3868 (N_3868,N_3731,N_3606);
nand U3869 (N_3869,N_3681,N_3616);
and U3870 (N_3870,N_3618,N_3686);
or U3871 (N_3871,N_3668,N_3696);
nor U3872 (N_3872,N_3643,N_3736);
or U3873 (N_3873,N_3730,N_3663);
and U3874 (N_3874,N_3717,N_3746);
nor U3875 (N_3875,N_3635,N_3653);
or U3876 (N_3876,N_3763,N_3649);
and U3877 (N_3877,N_3608,N_3694);
and U3878 (N_3878,N_3607,N_3641);
and U3879 (N_3879,N_3784,N_3712);
or U3880 (N_3880,N_3690,N_3691);
or U3881 (N_3881,N_3783,N_3609);
nor U3882 (N_3882,N_3666,N_3610);
nor U3883 (N_3883,N_3640,N_3715);
nand U3884 (N_3884,N_3602,N_3789);
nor U3885 (N_3885,N_3711,N_3622);
and U3886 (N_3886,N_3695,N_3656);
nand U3887 (N_3887,N_3633,N_3739);
or U3888 (N_3888,N_3785,N_3629);
nand U3889 (N_3889,N_3689,N_3678);
nor U3890 (N_3890,N_3747,N_3672);
nor U3891 (N_3891,N_3604,N_3749);
nand U3892 (N_3892,N_3655,N_3792);
nand U3893 (N_3893,N_3670,N_3699);
or U3894 (N_3894,N_3652,N_3772);
and U3895 (N_3895,N_3751,N_3673);
nand U3896 (N_3896,N_3779,N_3769);
or U3897 (N_3897,N_3726,N_3735);
and U3898 (N_3898,N_3745,N_3659);
nand U3899 (N_3899,N_3617,N_3654);
or U3900 (N_3900,N_3781,N_3756);
and U3901 (N_3901,N_3781,N_3727);
nor U3902 (N_3902,N_3688,N_3708);
nand U3903 (N_3903,N_3739,N_3647);
nor U3904 (N_3904,N_3611,N_3670);
nand U3905 (N_3905,N_3649,N_3620);
or U3906 (N_3906,N_3638,N_3753);
and U3907 (N_3907,N_3684,N_3757);
xor U3908 (N_3908,N_3741,N_3770);
and U3909 (N_3909,N_3725,N_3685);
and U3910 (N_3910,N_3696,N_3644);
nor U3911 (N_3911,N_3600,N_3617);
nand U3912 (N_3912,N_3737,N_3751);
or U3913 (N_3913,N_3789,N_3734);
nand U3914 (N_3914,N_3732,N_3718);
or U3915 (N_3915,N_3738,N_3728);
nor U3916 (N_3916,N_3612,N_3776);
and U3917 (N_3917,N_3653,N_3759);
nor U3918 (N_3918,N_3724,N_3753);
or U3919 (N_3919,N_3627,N_3616);
nand U3920 (N_3920,N_3685,N_3794);
nand U3921 (N_3921,N_3621,N_3697);
nand U3922 (N_3922,N_3747,N_3677);
or U3923 (N_3923,N_3704,N_3623);
or U3924 (N_3924,N_3629,N_3727);
nor U3925 (N_3925,N_3609,N_3650);
and U3926 (N_3926,N_3734,N_3609);
and U3927 (N_3927,N_3641,N_3648);
and U3928 (N_3928,N_3717,N_3644);
nor U3929 (N_3929,N_3615,N_3637);
nand U3930 (N_3930,N_3659,N_3622);
xnor U3931 (N_3931,N_3761,N_3790);
and U3932 (N_3932,N_3608,N_3697);
and U3933 (N_3933,N_3772,N_3707);
and U3934 (N_3934,N_3618,N_3720);
and U3935 (N_3935,N_3708,N_3733);
and U3936 (N_3936,N_3637,N_3711);
and U3937 (N_3937,N_3699,N_3654);
or U3938 (N_3938,N_3705,N_3793);
nor U3939 (N_3939,N_3628,N_3677);
nor U3940 (N_3940,N_3798,N_3646);
nor U3941 (N_3941,N_3673,N_3697);
nor U3942 (N_3942,N_3733,N_3786);
nor U3943 (N_3943,N_3641,N_3634);
and U3944 (N_3944,N_3695,N_3794);
or U3945 (N_3945,N_3752,N_3749);
or U3946 (N_3946,N_3621,N_3727);
and U3947 (N_3947,N_3759,N_3610);
nor U3948 (N_3948,N_3759,N_3767);
nor U3949 (N_3949,N_3731,N_3730);
nor U3950 (N_3950,N_3628,N_3724);
and U3951 (N_3951,N_3613,N_3734);
xnor U3952 (N_3952,N_3752,N_3789);
nor U3953 (N_3953,N_3639,N_3683);
nand U3954 (N_3954,N_3685,N_3796);
and U3955 (N_3955,N_3767,N_3755);
and U3956 (N_3956,N_3600,N_3750);
nor U3957 (N_3957,N_3770,N_3633);
nand U3958 (N_3958,N_3611,N_3624);
and U3959 (N_3959,N_3671,N_3741);
and U3960 (N_3960,N_3706,N_3607);
nor U3961 (N_3961,N_3709,N_3630);
and U3962 (N_3962,N_3732,N_3782);
or U3963 (N_3963,N_3794,N_3657);
and U3964 (N_3964,N_3682,N_3727);
and U3965 (N_3965,N_3758,N_3635);
nor U3966 (N_3966,N_3648,N_3682);
or U3967 (N_3967,N_3754,N_3642);
nor U3968 (N_3968,N_3714,N_3713);
nor U3969 (N_3969,N_3723,N_3741);
or U3970 (N_3970,N_3698,N_3733);
and U3971 (N_3971,N_3682,N_3603);
or U3972 (N_3972,N_3652,N_3716);
and U3973 (N_3973,N_3733,N_3696);
nor U3974 (N_3974,N_3751,N_3717);
nand U3975 (N_3975,N_3689,N_3733);
or U3976 (N_3976,N_3676,N_3659);
nand U3977 (N_3977,N_3737,N_3679);
and U3978 (N_3978,N_3621,N_3787);
or U3979 (N_3979,N_3628,N_3603);
nor U3980 (N_3980,N_3620,N_3744);
nand U3981 (N_3981,N_3623,N_3652);
nor U3982 (N_3982,N_3663,N_3629);
xnor U3983 (N_3983,N_3788,N_3610);
or U3984 (N_3984,N_3734,N_3675);
nor U3985 (N_3985,N_3676,N_3762);
and U3986 (N_3986,N_3752,N_3768);
and U3987 (N_3987,N_3795,N_3735);
xor U3988 (N_3988,N_3738,N_3763);
and U3989 (N_3989,N_3754,N_3795);
or U3990 (N_3990,N_3612,N_3696);
nor U3991 (N_3991,N_3698,N_3742);
nor U3992 (N_3992,N_3636,N_3789);
nor U3993 (N_3993,N_3670,N_3712);
and U3994 (N_3994,N_3754,N_3735);
nand U3995 (N_3995,N_3727,N_3758);
or U3996 (N_3996,N_3717,N_3787);
xnor U3997 (N_3997,N_3734,N_3757);
and U3998 (N_3998,N_3629,N_3658);
nor U3999 (N_3999,N_3716,N_3704);
nor U4000 (N_4000,N_3895,N_3903);
or U4001 (N_4001,N_3804,N_3847);
and U4002 (N_4002,N_3999,N_3884);
nand U4003 (N_4003,N_3880,N_3953);
nand U4004 (N_4004,N_3936,N_3961);
nor U4005 (N_4005,N_3835,N_3938);
and U4006 (N_4006,N_3944,N_3990);
nor U4007 (N_4007,N_3877,N_3874);
or U4008 (N_4008,N_3818,N_3948);
and U4009 (N_4009,N_3968,N_3997);
nor U4010 (N_4010,N_3969,N_3916);
nor U4011 (N_4011,N_3917,N_3933);
or U4012 (N_4012,N_3855,N_3918);
nand U4013 (N_4013,N_3977,N_3955);
or U4014 (N_4014,N_3888,N_3891);
or U4015 (N_4015,N_3849,N_3803);
nand U4016 (N_4016,N_3889,N_3947);
and U4017 (N_4017,N_3843,N_3846);
nand U4018 (N_4018,N_3975,N_3960);
nor U4019 (N_4019,N_3992,N_3870);
nor U4020 (N_4020,N_3905,N_3829);
nor U4021 (N_4021,N_3890,N_3908);
nand U4022 (N_4022,N_3812,N_3909);
and U4023 (N_4023,N_3831,N_3963);
nand U4024 (N_4024,N_3808,N_3988);
nor U4025 (N_4025,N_3876,N_3943);
nand U4026 (N_4026,N_3979,N_3817);
nor U4027 (N_4027,N_3896,N_3993);
and U4028 (N_4028,N_3851,N_3872);
nand U4029 (N_4029,N_3914,N_3920);
and U4030 (N_4030,N_3940,N_3996);
nor U4031 (N_4031,N_3815,N_3939);
nand U4032 (N_4032,N_3838,N_3930);
or U4033 (N_4033,N_3973,N_3971);
nand U4034 (N_4034,N_3964,N_3864);
nand U4035 (N_4035,N_3879,N_3816);
nor U4036 (N_4036,N_3887,N_3982);
xor U4037 (N_4037,N_3922,N_3994);
nand U4038 (N_4038,N_3910,N_3952);
nand U4039 (N_4039,N_3806,N_3929);
nor U4040 (N_4040,N_3809,N_3937);
nor U4041 (N_4041,N_3972,N_3956);
nand U4042 (N_4042,N_3998,N_3913);
nand U4043 (N_4043,N_3919,N_3859);
nor U4044 (N_4044,N_3853,N_3981);
and U4045 (N_4045,N_3901,N_3986);
or U4046 (N_4046,N_3819,N_3927);
and U4047 (N_4047,N_3946,N_3915);
or U4048 (N_4048,N_3827,N_3912);
and U4049 (N_4049,N_3902,N_3850);
or U4050 (N_4050,N_3984,N_3906);
and U4051 (N_4051,N_3823,N_3878);
and U4052 (N_4052,N_3957,N_3983);
nor U4053 (N_4053,N_3942,N_3980);
and U4054 (N_4054,N_3836,N_3951);
nand U4055 (N_4055,N_3894,N_3867);
nand U4056 (N_4056,N_3842,N_3868);
or U4057 (N_4057,N_3958,N_3935);
or U4058 (N_4058,N_3845,N_3862);
or U4059 (N_4059,N_3925,N_3826);
and U4060 (N_4060,N_3871,N_3805);
nand U4061 (N_4061,N_3813,N_3932);
nor U4062 (N_4062,N_3873,N_3856);
nand U4063 (N_4063,N_3924,N_3921);
or U4064 (N_4064,N_3950,N_3800);
nand U4065 (N_4065,N_3865,N_3885);
nor U4066 (N_4066,N_3852,N_3987);
nand U4067 (N_4067,N_3841,N_3883);
or U4068 (N_4068,N_3866,N_3834);
or U4069 (N_4069,N_3822,N_3959);
nand U4070 (N_4070,N_3810,N_3840);
and U4071 (N_4071,N_3985,N_3978);
and U4072 (N_4072,N_3898,N_3860);
or U4073 (N_4073,N_3811,N_3821);
nand U4074 (N_4074,N_3814,N_3967);
or U4075 (N_4075,N_3928,N_3854);
and U4076 (N_4076,N_3875,N_3892);
nor U4077 (N_4077,N_3825,N_3820);
or U4078 (N_4078,N_3833,N_3900);
nor U4079 (N_4079,N_3839,N_3857);
nand U4080 (N_4080,N_3844,N_3966);
nand U4081 (N_4081,N_3897,N_3881);
or U4082 (N_4082,N_3907,N_3954);
nand U4083 (N_4083,N_3869,N_3941);
and U4084 (N_4084,N_3899,N_3949);
and U4085 (N_4085,N_3807,N_3991);
or U4086 (N_4086,N_3904,N_3848);
and U4087 (N_4087,N_3863,N_3837);
or U4088 (N_4088,N_3886,N_3926);
nand U4089 (N_4089,N_3934,N_3974);
and U4090 (N_4090,N_3861,N_3911);
and U4091 (N_4091,N_3962,N_3995);
or U4092 (N_4092,N_3931,N_3976);
and U4093 (N_4093,N_3989,N_3858);
nor U4094 (N_4094,N_3923,N_3832);
or U4095 (N_4095,N_3824,N_3945);
and U4096 (N_4096,N_3882,N_3801);
or U4097 (N_4097,N_3965,N_3802);
nor U4098 (N_4098,N_3970,N_3830);
nand U4099 (N_4099,N_3828,N_3893);
nand U4100 (N_4100,N_3990,N_3997);
nor U4101 (N_4101,N_3932,N_3991);
nand U4102 (N_4102,N_3932,N_3881);
nand U4103 (N_4103,N_3850,N_3950);
or U4104 (N_4104,N_3917,N_3955);
or U4105 (N_4105,N_3897,N_3850);
nand U4106 (N_4106,N_3874,N_3884);
nand U4107 (N_4107,N_3890,N_3878);
or U4108 (N_4108,N_3800,N_3874);
or U4109 (N_4109,N_3993,N_3822);
xor U4110 (N_4110,N_3886,N_3895);
xnor U4111 (N_4111,N_3918,N_3978);
and U4112 (N_4112,N_3941,N_3864);
xor U4113 (N_4113,N_3838,N_3958);
or U4114 (N_4114,N_3879,N_3960);
or U4115 (N_4115,N_3887,N_3915);
nand U4116 (N_4116,N_3842,N_3884);
nor U4117 (N_4117,N_3880,N_3818);
or U4118 (N_4118,N_3814,N_3962);
nor U4119 (N_4119,N_3982,N_3977);
nor U4120 (N_4120,N_3837,N_3893);
nand U4121 (N_4121,N_3883,N_3818);
and U4122 (N_4122,N_3938,N_3958);
nand U4123 (N_4123,N_3981,N_3801);
nand U4124 (N_4124,N_3813,N_3968);
or U4125 (N_4125,N_3951,N_3972);
nor U4126 (N_4126,N_3991,N_3860);
or U4127 (N_4127,N_3899,N_3884);
or U4128 (N_4128,N_3849,N_3998);
and U4129 (N_4129,N_3858,N_3950);
or U4130 (N_4130,N_3890,N_3863);
nand U4131 (N_4131,N_3929,N_3983);
and U4132 (N_4132,N_3803,N_3919);
or U4133 (N_4133,N_3863,N_3937);
nand U4134 (N_4134,N_3944,N_3896);
nor U4135 (N_4135,N_3862,N_3858);
and U4136 (N_4136,N_3906,N_3968);
nand U4137 (N_4137,N_3890,N_3814);
and U4138 (N_4138,N_3916,N_3842);
xor U4139 (N_4139,N_3931,N_3820);
or U4140 (N_4140,N_3846,N_3805);
or U4141 (N_4141,N_3863,N_3952);
nor U4142 (N_4142,N_3931,N_3858);
nor U4143 (N_4143,N_3843,N_3898);
or U4144 (N_4144,N_3849,N_3935);
or U4145 (N_4145,N_3943,N_3808);
and U4146 (N_4146,N_3988,N_3947);
and U4147 (N_4147,N_3923,N_3962);
and U4148 (N_4148,N_3840,N_3955);
xnor U4149 (N_4149,N_3949,N_3982);
nor U4150 (N_4150,N_3847,N_3873);
nor U4151 (N_4151,N_3948,N_3846);
nand U4152 (N_4152,N_3999,N_3860);
or U4153 (N_4153,N_3851,N_3808);
xnor U4154 (N_4154,N_3893,N_3818);
nor U4155 (N_4155,N_3846,N_3853);
nand U4156 (N_4156,N_3940,N_3829);
and U4157 (N_4157,N_3916,N_3860);
or U4158 (N_4158,N_3928,N_3962);
and U4159 (N_4159,N_3824,N_3896);
nand U4160 (N_4160,N_3895,N_3872);
nand U4161 (N_4161,N_3801,N_3961);
or U4162 (N_4162,N_3867,N_3960);
nor U4163 (N_4163,N_3855,N_3981);
or U4164 (N_4164,N_3856,N_3854);
nand U4165 (N_4165,N_3976,N_3889);
or U4166 (N_4166,N_3982,N_3950);
or U4167 (N_4167,N_3838,N_3899);
or U4168 (N_4168,N_3901,N_3945);
or U4169 (N_4169,N_3884,N_3994);
nor U4170 (N_4170,N_3841,N_3890);
or U4171 (N_4171,N_3875,N_3882);
xor U4172 (N_4172,N_3860,N_3937);
nor U4173 (N_4173,N_3885,N_3819);
nor U4174 (N_4174,N_3876,N_3800);
or U4175 (N_4175,N_3845,N_3975);
nand U4176 (N_4176,N_3885,N_3863);
or U4177 (N_4177,N_3936,N_3830);
and U4178 (N_4178,N_3883,N_3817);
nand U4179 (N_4179,N_3955,N_3802);
nor U4180 (N_4180,N_3882,N_3866);
nor U4181 (N_4181,N_3871,N_3951);
and U4182 (N_4182,N_3822,N_3800);
nand U4183 (N_4183,N_3944,N_3809);
nand U4184 (N_4184,N_3986,N_3939);
nand U4185 (N_4185,N_3973,N_3931);
nand U4186 (N_4186,N_3937,N_3997);
nor U4187 (N_4187,N_3812,N_3829);
and U4188 (N_4188,N_3883,N_3822);
or U4189 (N_4189,N_3802,N_3900);
and U4190 (N_4190,N_3836,N_3969);
and U4191 (N_4191,N_3897,N_3964);
and U4192 (N_4192,N_3810,N_3904);
and U4193 (N_4193,N_3905,N_3892);
nand U4194 (N_4194,N_3809,N_3982);
nand U4195 (N_4195,N_3870,N_3982);
or U4196 (N_4196,N_3959,N_3802);
nor U4197 (N_4197,N_3907,N_3910);
or U4198 (N_4198,N_3861,N_3994);
and U4199 (N_4199,N_3820,N_3859);
or U4200 (N_4200,N_4041,N_4112);
nor U4201 (N_4201,N_4139,N_4126);
or U4202 (N_4202,N_4008,N_4158);
or U4203 (N_4203,N_4042,N_4070);
nor U4204 (N_4204,N_4075,N_4085);
nor U4205 (N_4205,N_4183,N_4186);
or U4206 (N_4206,N_4147,N_4095);
or U4207 (N_4207,N_4163,N_4198);
nand U4208 (N_4208,N_4048,N_4065);
and U4209 (N_4209,N_4150,N_4006);
nor U4210 (N_4210,N_4140,N_4098);
nor U4211 (N_4211,N_4014,N_4117);
and U4212 (N_4212,N_4109,N_4050);
nor U4213 (N_4213,N_4052,N_4015);
and U4214 (N_4214,N_4038,N_4174);
and U4215 (N_4215,N_4175,N_4187);
nor U4216 (N_4216,N_4011,N_4033);
nor U4217 (N_4217,N_4181,N_4137);
nor U4218 (N_4218,N_4021,N_4184);
xnor U4219 (N_4219,N_4125,N_4083);
nand U4220 (N_4220,N_4020,N_4162);
or U4221 (N_4221,N_4113,N_4111);
nor U4222 (N_4222,N_4101,N_4130);
nor U4223 (N_4223,N_4051,N_4080);
nor U4224 (N_4224,N_4012,N_4056);
nand U4225 (N_4225,N_4082,N_4149);
nand U4226 (N_4226,N_4010,N_4049);
and U4227 (N_4227,N_4122,N_4156);
and U4228 (N_4228,N_4036,N_4157);
or U4229 (N_4229,N_4058,N_4100);
nand U4230 (N_4230,N_4035,N_4005);
nand U4231 (N_4231,N_4000,N_4135);
nor U4232 (N_4232,N_4096,N_4024);
and U4233 (N_4233,N_4195,N_4031);
nand U4234 (N_4234,N_4002,N_4123);
and U4235 (N_4235,N_4099,N_4097);
or U4236 (N_4236,N_4191,N_4120);
or U4237 (N_4237,N_4182,N_4196);
or U4238 (N_4238,N_4034,N_4009);
and U4239 (N_4239,N_4061,N_4073);
nor U4240 (N_4240,N_4164,N_4040);
nor U4241 (N_4241,N_4161,N_4177);
nand U4242 (N_4242,N_4043,N_4013);
xnor U4243 (N_4243,N_4023,N_4017);
or U4244 (N_4244,N_4068,N_4172);
xor U4245 (N_4245,N_4067,N_4119);
nand U4246 (N_4246,N_4141,N_4190);
nand U4247 (N_4247,N_4054,N_4071);
nor U4248 (N_4248,N_4136,N_4094);
xor U4249 (N_4249,N_4188,N_4121);
or U4250 (N_4250,N_4108,N_4007);
nor U4251 (N_4251,N_4145,N_4084);
or U4252 (N_4252,N_4062,N_4037);
nor U4253 (N_4253,N_4151,N_4199);
and U4254 (N_4254,N_4091,N_4107);
nand U4255 (N_4255,N_4066,N_4127);
nor U4256 (N_4256,N_4060,N_4086);
nor U4257 (N_4257,N_4046,N_4001);
nand U4258 (N_4258,N_4003,N_4105);
nor U4259 (N_4259,N_4092,N_4167);
and U4260 (N_4260,N_4131,N_4078);
or U4261 (N_4261,N_4064,N_4176);
nand U4262 (N_4262,N_4045,N_4088);
nor U4263 (N_4263,N_4044,N_4178);
nor U4264 (N_4264,N_4025,N_4171);
and U4265 (N_4265,N_4133,N_4146);
or U4266 (N_4266,N_4154,N_4159);
and U4267 (N_4267,N_4197,N_4170);
nand U4268 (N_4268,N_4193,N_4155);
nand U4269 (N_4269,N_4055,N_4192);
nor U4270 (N_4270,N_4160,N_4019);
and U4271 (N_4271,N_4028,N_4004);
nand U4272 (N_4272,N_4029,N_4148);
nor U4273 (N_4273,N_4132,N_4194);
nor U4274 (N_4274,N_4018,N_4063);
or U4275 (N_4275,N_4026,N_4103);
or U4276 (N_4276,N_4134,N_4189);
and U4277 (N_4277,N_4027,N_4076);
nand U4278 (N_4278,N_4152,N_4114);
or U4279 (N_4279,N_4087,N_4169);
nor U4280 (N_4280,N_4079,N_4118);
nand U4281 (N_4281,N_4110,N_4074);
nand U4282 (N_4282,N_4168,N_4081);
and U4283 (N_4283,N_4102,N_4116);
and U4284 (N_4284,N_4153,N_4059);
and U4285 (N_4285,N_4142,N_4138);
and U4286 (N_4286,N_4129,N_4093);
and U4287 (N_4287,N_4185,N_4022);
and U4288 (N_4288,N_4104,N_4072);
or U4289 (N_4289,N_4166,N_4047);
nand U4290 (N_4290,N_4173,N_4089);
nand U4291 (N_4291,N_4180,N_4115);
or U4292 (N_4292,N_4179,N_4069);
or U4293 (N_4293,N_4144,N_4165);
or U4294 (N_4294,N_4106,N_4039);
nand U4295 (N_4295,N_4128,N_4077);
nor U4296 (N_4296,N_4030,N_4053);
and U4297 (N_4297,N_4090,N_4143);
nor U4298 (N_4298,N_4124,N_4057);
or U4299 (N_4299,N_4032,N_4016);
nor U4300 (N_4300,N_4024,N_4061);
nor U4301 (N_4301,N_4138,N_4144);
and U4302 (N_4302,N_4025,N_4038);
nand U4303 (N_4303,N_4089,N_4006);
or U4304 (N_4304,N_4018,N_4026);
nand U4305 (N_4305,N_4085,N_4003);
and U4306 (N_4306,N_4126,N_4114);
or U4307 (N_4307,N_4015,N_4002);
and U4308 (N_4308,N_4028,N_4140);
or U4309 (N_4309,N_4159,N_4100);
or U4310 (N_4310,N_4049,N_4057);
or U4311 (N_4311,N_4198,N_4010);
or U4312 (N_4312,N_4025,N_4035);
or U4313 (N_4313,N_4174,N_4070);
or U4314 (N_4314,N_4177,N_4171);
nor U4315 (N_4315,N_4160,N_4028);
and U4316 (N_4316,N_4066,N_4098);
nor U4317 (N_4317,N_4185,N_4032);
and U4318 (N_4318,N_4001,N_4094);
nand U4319 (N_4319,N_4080,N_4040);
nor U4320 (N_4320,N_4043,N_4120);
and U4321 (N_4321,N_4118,N_4175);
and U4322 (N_4322,N_4085,N_4157);
nor U4323 (N_4323,N_4061,N_4106);
and U4324 (N_4324,N_4167,N_4121);
nand U4325 (N_4325,N_4018,N_4079);
nor U4326 (N_4326,N_4093,N_4167);
nand U4327 (N_4327,N_4048,N_4154);
or U4328 (N_4328,N_4001,N_4088);
nand U4329 (N_4329,N_4086,N_4089);
and U4330 (N_4330,N_4157,N_4169);
or U4331 (N_4331,N_4088,N_4107);
and U4332 (N_4332,N_4013,N_4045);
nand U4333 (N_4333,N_4014,N_4132);
nor U4334 (N_4334,N_4104,N_4113);
nand U4335 (N_4335,N_4060,N_4116);
nor U4336 (N_4336,N_4182,N_4118);
nor U4337 (N_4337,N_4032,N_4004);
nor U4338 (N_4338,N_4155,N_4064);
nor U4339 (N_4339,N_4023,N_4065);
nor U4340 (N_4340,N_4086,N_4114);
nand U4341 (N_4341,N_4018,N_4186);
nor U4342 (N_4342,N_4123,N_4069);
nor U4343 (N_4343,N_4006,N_4025);
or U4344 (N_4344,N_4188,N_4162);
and U4345 (N_4345,N_4005,N_4108);
and U4346 (N_4346,N_4083,N_4163);
or U4347 (N_4347,N_4195,N_4114);
nand U4348 (N_4348,N_4103,N_4091);
nor U4349 (N_4349,N_4199,N_4017);
nor U4350 (N_4350,N_4104,N_4005);
nor U4351 (N_4351,N_4142,N_4157);
nor U4352 (N_4352,N_4067,N_4099);
nor U4353 (N_4353,N_4154,N_4134);
nor U4354 (N_4354,N_4113,N_4057);
and U4355 (N_4355,N_4152,N_4031);
or U4356 (N_4356,N_4072,N_4016);
nor U4357 (N_4357,N_4065,N_4032);
and U4358 (N_4358,N_4056,N_4133);
xor U4359 (N_4359,N_4087,N_4162);
nand U4360 (N_4360,N_4001,N_4081);
or U4361 (N_4361,N_4076,N_4083);
nand U4362 (N_4362,N_4178,N_4075);
nand U4363 (N_4363,N_4154,N_4120);
xnor U4364 (N_4364,N_4077,N_4161);
nor U4365 (N_4365,N_4153,N_4190);
and U4366 (N_4366,N_4060,N_4001);
or U4367 (N_4367,N_4128,N_4160);
nor U4368 (N_4368,N_4087,N_4058);
nand U4369 (N_4369,N_4137,N_4100);
and U4370 (N_4370,N_4014,N_4172);
or U4371 (N_4371,N_4133,N_4100);
nand U4372 (N_4372,N_4131,N_4006);
or U4373 (N_4373,N_4195,N_4071);
nand U4374 (N_4374,N_4146,N_4193);
nand U4375 (N_4375,N_4070,N_4177);
nor U4376 (N_4376,N_4069,N_4121);
or U4377 (N_4377,N_4061,N_4105);
and U4378 (N_4378,N_4034,N_4061);
and U4379 (N_4379,N_4185,N_4178);
and U4380 (N_4380,N_4198,N_4104);
or U4381 (N_4381,N_4078,N_4167);
or U4382 (N_4382,N_4017,N_4120);
and U4383 (N_4383,N_4083,N_4157);
or U4384 (N_4384,N_4118,N_4027);
nor U4385 (N_4385,N_4038,N_4173);
or U4386 (N_4386,N_4047,N_4113);
or U4387 (N_4387,N_4194,N_4178);
or U4388 (N_4388,N_4073,N_4072);
nor U4389 (N_4389,N_4079,N_4175);
and U4390 (N_4390,N_4034,N_4197);
xor U4391 (N_4391,N_4109,N_4117);
nor U4392 (N_4392,N_4091,N_4106);
nor U4393 (N_4393,N_4080,N_4089);
nand U4394 (N_4394,N_4083,N_4040);
nor U4395 (N_4395,N_4076,N_4067);
nand U4396 (N_4396,N_4027,N_4019);
nand U4397 (N_4397,N_4045,N_4196);
nor U4398 (N_4398,N_4105,N_4107);
nor U4399 (N_4399,N_4191,N_4002);
nand U4400 (N_4400,N_4278,N_4219);
nor U4401 (N_4401,N_4246,N_4314);
and U4402 (N_4402,N_4396,N_4300);
nand U4403 (N_4403,N_4366,N_4276);
xor U4404 (N_4404,N_4390,N_4211);
and U4405 (N_4405,N_4348,N_4372);
nand U4406 (N_4406,N_4331,N_4303);
or U4407 (N_4407,N_4251,N_4273);
nor U4408 (N_4408,N_4376,N_4228);
nor U4409 (N_4409,N_4325,N_4321);
nand U4410 (N_4410,N_4234,N_4281);
and U4411 (N_4411,N_4245,N_4326);
or U4412 (N_4412,N_4237,N_4262);
nor U4413 (N_4413,N_4227,N_4289);
and U4414 (N_4414,N_4265,N_4214);
nor U4415 (N_4415,N_4272,N_4339);
and U4416 (N_4416,N_4240,N_4296);
nor U4417 (N_4417,N_4329,N_4369);
nand U4418 (N_4418,N_4375,N_4255);
nand U4419 (N_4419,N_4288,N_4370);
and U4420 (N_4420,N_4371,N_4290);
and U4421 (N_4421,N_4304,N_4285);
nor U4422 (N_4422,N_4355,N_4308);
nor U4423 (N_4423,N_4307,N_4367);
or U4424 (N_4424,N_4384,N_4202);
and U4425 (N_4425,N_4336,N_4378);
and U4426 (N_4426,N_4381,N_4385);
nor U4427 (N_4427,N_4218,N_4226);
nor U4428 (N_4428,N_4342,N_4270);
nor U4429 (N_4429,N_4395,N_4284);
nor U4430 (N_4430,N_4264,N_4200);
nand U4431 (N_4431,N_4216,N_4244);
and U4432 (N_4432,N_4340,N_4206);
nand U4433 (N_4433,N_4324,N_4388);
nand U4434 (N_4434,N_4305,N_4221);
and U4435 (N_4435,N_4347,N_4253);
nand U4436 (N_4436,N_4256,N_4349);
nor U4437 (N_4437,N_4343,N_4287);
nor U4438 (N_4438,N_4322,N_4241);
or U4439 (N_4439,N_4391,N_4338);
and U4440 (N_4440,N_4360,N_4382);
and U4441 (N_4441,N_4350,N_4368);
or U4442 (N_4442,N_4269,N_4373);
nor U4443 (N_4443,N_4298,N_4243);
xnor U4444 (N_4444,N_4248,N_4328);
nor U4445 (N_4445,N_4271,N_4260);
or U4446 (N_4446,N_4351,N_4306);
and U4447 (N_4447,N_4389,N_4266);
and U4448 (N_4448,N_4239,N_4286);
or U4449 (N_4449,N_4359,N_4249);
nor U4450 (N_4450,N_4282,N_4380);
nor U4451 (N_4451,N_4250,N_4210);
nand U4452 (N_4452,N_4275,N_4313);
or U4453 (N_4453,N_4230,N_4365);
or U4454 (N_4454,N_4293,N_4204);
nand U4455 (N_4455,N_4398,N_4242);
or U4456 (N_4456,N_4309,N_4361);
xor U4457 (N_4457,N_4292,N_4223);
nand U4458 (N_4458,N_4315,N_4310);
or U4459 (N_4459,N_4279,N_4301);
or U4460 (N_4460,N_4252,N_4354);
xor U4461 (N_4461,N_4297,N_4217);
nand U4462 (N_4462,N_4235,N_4358);
nand U4463 (N_4463,N_4268,N_4299);
and U4464 (N_4464,N_4224,N_4316);
and U4465 (N_4465,N_4352,N_4311);
and U4466 (N_4466,N_4332,N_4220);
nand U4467 (N_4467,N_4263,N_4330);
and U4468 (N_4468,N_4319,N_4203);
nand U4469 (N_4469,N_4229,N_4222);
xor U4470 (N_4470,N_4335,N_4212);
nand U4471 (N_4471,N_4302,N_4259);
and U4472 (N_4472,N_4379,N_4267);
nor U4473 (N_4473,N_4277,N_4232);
and U4474 (N_4474,N_4387,N_4261);
nand U4475 (N_4475,N_4333,N_4394);
or U4476 (N_4476,N_4291,N_4236);
nand U4477 (N_4477,N_4392,N_4374);
nor U4478 (N_4478,N_4257,N_4208);
nand U4479 (N_4479,N_4357,N_4327);
and U4480 (N_4480,N_4207,N_4386);
nand U4481 (N_4481,N_4231,N_4399);
nor U4482 (N_4482,N_4362,N_4283);
nand U4483 (N_4483,N_4295,N_4337);
nor U4484 (N_4484,N_4274,N_4205);
or U4485 (N_4485,N_4233,N_4213);
or U4486 (N_4486,N_4377,N_4383);
or U4487 (N_4487,N_4344,N_4318);
nand U4488 (N_4488,N_4317,N_4294);
and U4489 (N_4489,N_4341,N_4346);
nand U4490 (N_4490,N_4247,N_4254);
nor U4491 (N_4491,N_4320,N_4225);
and U4492 (N_4492,N_4258,N_4215);
or U4493 (N_4493,N_4201,N_4364);
nand U4494 (N_4494,N_4238,N_4353);
and U4495 (N_4495,N_4334,N_4397);
nor U4496 (N_4496,N_4323,N_4363);
and U4497 (N_4497,N_4345,N_4312);
nand U4498 (N_4498,N_4209,N_4280);
nand U4499 (N_4499,N_4393,N_4356);
nor U4500 (N_4500,N_4372,N_4285);
nor U4501 (N_4501,N_4320,N_4239);
nand U4502 (N_4502,N_4251,N_4328);
or U4503 (N_4503,N_4394,N_4281);
nor U4504 (N_4504,N_4265,N_4399);
or U4505 (N_4505,N_4270,N_4207);
and U4506 (N_4506,N_4234,N_4296);
or U4507 (N_4507,N_4397,N_4267);
xnor U4508 (N_4508,N_4363,N_4312);
and U4509 (N_4509,N_4221,N_4377);
nor U4510 (N_4510,N_4261,N_4266);
nand U4511 (N_4511,N_4325,N_4271);
nor U4512 (N_4512,N_4386,N_4270);
nand U4513 (N_4513,N_4294,N_4203);
nor U4514 (N_4514,N_4230,N_4289);
nor U4515 (N_4515,N_4282,N_4353);
or U4516 (N_4516,N_4275,N_4350);
nand U4517 (N_4517,N_4223,N_4304);
nand U4518 (N_4518,N_4330,N_4245);
or U4519 (N_4519,N_4294,N_4376);
nor U4520 (N_4520,N_4383,N_4223);
and U4521 (N_4521,N_4366,N_4292);
nor U4522 (N_4522,N_4254,N_4364);
nor U4523 (N_4523,N_4295,N_4379);
nand U4524 (N_4524,N_4365,N_4279);
or U4525 (N_4525,N_4257,N_4342);
nand U4526 (N_4526,N_4387,N_4394);
nor U4527 (N_4527,N_4302,N_4376);
nor U4528 (N_4528,N_4212,N_4293);
nand U4529 (N_4529,N_4207,N_4373);
nand U4530 (N_4530,N_4391,N_4348);
and U4531 (N_4531,N_4366,N_4333);
and U4532 (N_4532,N_4356,N_4331);
nor U4533 (N_4533,N_4214,N_4278);
and U4534 (N_4534,N_4209,N_4272);
nand U4535 (N_4535,N_4225,N_4221);
or U4536 (N_4536,N_4372,N_4265);
nor U4537 (N_4537,N_4249,N_4340);
nand U4538 (N_4538,N_4367,N_4365);
or U4539 (N_4539,N_4213,N_4331);
nor U4540 (N_4540,N_4264,N_4309);
or U4541 (N_4541,N_4298,N_4286);
nor U4542 (N_4542,N_4335,N_4255);
nand U4543 (N_4543,N_4213,N_4235);
and U4544 (N_4544,N_4364,N_4331);
and U4545 (N_4545,N_4245,N_4258);
nand U4546 (N_4546,N_4367,N_4274);
and U4547 (N_4547,N_4222,N_4236);
nor U4548 (N_4548,N_4346,N_4231);
or U4549 (N_4549,N_4308,N_4331);
nor U4550 (N_4550,N_4264,N_4206);
or U4551 (N_4551,N_4299,N_4356);
nand U4552 (N_4552,N_4326,N_4377);
and U4553 (N_4553,N_4326,N_4313);
nor U4554 (N_4554,N_4225,N_4227);
nand U4555 (N_4555,N_4313,N_4376);
xnor U4556 (N_4556,N_4352,N_4375);
nor U4557 (N_4557,N_4211,N_4330);
and U4558 (N_4558,N_4281,N_4320);
or U4559 (N_4559,N_4346,N_4290);
or U4560 (N_4560,N_4362,N_4263);
nor U4561 (N_4561,N_4294,N_4204);
or U4562 (N_4562,N_4277,N_4268);
nor U4563 (N_4563,N_4295,N_4288);
and U4564 (N_4564,N_4326,N_4389);
nand U4565 (N_4565,N_4312,N_4394);
nor U4566 (N_4566,N_4320,N_4299);
nor U4567 (N_4567,N_4349,N_4274);
nor U4568 (N_4568,N_4202,N_4241);
nor U4569 (N_4569,N_4258,N_4318);
or U4570 (N_4570,N_4269,N_4340);
nor U4571 (N_4571,N_4260,N_4303);
nor U4572 (N_4572,N_4265,N_4285);
nand U4573 (N_4573,N_4200,N_4201);
or U4574 (N_4574,N_4211,N_4393);
and U4575 (N_4575,N_4374,N_4372);
nor U4576 (N_4576,N_4251,N_4232);
nand U4577 (N_4577,N_4210,N_4232);
or U4578 (N_4578,N_4288,N_4200);
nor U4579 (N_4579,N_4342,N_4398);
nor U4580 (N_4580,N_4211,N_4321);
nor U4581 (N_4581,N_4221,N_4313);
nand U4582 (N_4582,N_4264,N_4344);
nor U4583 (N_4583,N_4328,N_4284);
and U4584 (N_4584,N_4280,N_4325);
nand U4585 (N_4585,N_4248,N_4338);
nor U4586 (N_4586,N_4301,N_4399);
nor U4587 (N_4587,N_4310,N_4396);
nand U4588 (N_4588,N_4379,N_4266);
or U4589 (N_4589,N_4230,N_4253);
nand U4590 (N_4590,N_4322,N_4255);
nor U4591 (N_4591,N_4272,N_4344);
nand U4592 (N_4592,N_4220,N_4252);
and U4593 (N_4593,N_4257,N_4290);
and U4594 (N_4594,N_4373,N_4359);
and U4595 (N_4595,N_4233,N_4294);
or U4596 (N_4596,N_4230,N_4242);
nand U4597 (N_4597,N_4268,N_4281);
or U4598 (N_4598,N_4260,N_4317);
and U4599 (N_4599,N_4357,N_4323);
or U4600 (N_4600,N_4580,N_4505);
nand U4601 (N_4601,N_4585,N_4526);
nand U4602 (N_4602,N_4579,N_4570);
nor U4603 (N_4603,N_4592,N_4406);
nor U4604 (N_4604,N_4460,N_4556);
nor U4605 (N_4605,N_4475,N_4576);
nand U4606 (N_4606,N_4539,N_4586);
nand U4607 (N_4607,N_4495,N_4424);
and U4608 (N_4608,N_4550,N_4467);
and U4609 (N_4609,N_4498,N_4554);
or U4610 (N_4610,N_4553,N_4582);
and U4611 (N_4611,N_4490,N_4531);
nor U4612 (N_4612,N_4534,N_4519);
nor U4613 (N_4613,N_4563,N_4469);
nand U4614 (N_4614,N_4546,N_4599);
nand U4615 (N_4615,N_4464,N_4566);
nor U4616 (N_4616,N_4513,N_4412);
and U4617 (N_4617,N_4423,N_4438);
xor U4618 (N_4618,N_4597,N_4559);
nor U4619 (N_4619,N_4584,N_4588);
nor U4620 (N_4620,N_4535,N_4405);
nand U4621 (N_4621,N_4598,N_4436);
nand U4622 (N_4622,N_4596,N_4497);
or U4623 (N_4623,N_4448,N_4434);
or U4624 (N_4624,N_4451,N_4400);
or U4625 (N_4625,N_4578,N_4525);
nor U4626 (N_4626,N_4502,N_4510);
xnor U4627 (N_4627,N_4545,N_4575);
and U4628 (N_4628,N_4516,N_4453);
nor U4629 (N_4629,N_4470,N_4476);
and U4630 (N_4630,N_4521,N_4493);
nor U4631 (N_4631,N_4454,N_4547);
nor U4632 (N_4632,N_4541,N_4418);
or U4633 (N_4633,N_4552,N_4573);
nor U4634 (N_4634,N_4408,N_4428);
and U4635 (N_4635,N_4480,N_4419);
nand U4636 (N_4636,N_4549,N_4462);
nor U4637 (N_4637,N_4574,N_4414);
or U4638 (N_4638,N_4415,N_4445);
nand U4639 (N_4639,N_4427,N_4489);
nor U4640 (N_4640,N_4520,N_4407);
nand U4641 (N_4641,N_4401,N_4593);
nand U4642 (N_4642,N_4595,N_4509);
and U4643 (N_4643,N_4583,N_4536);
or U4644 (N_4644,N_4538,N_4555);
and U4645 (N_4645,N_4561,N_4416);
nor U4646 (N_4646,N_4506,N_4457);
nand U4647 (N_4647,N_4442,N_4494);
and U4648 (N_4648,N_4444,N_4523);
and U4649 (N_4649,N_4540,N_4590);
xnor U4650 (N_4650,N_4569,N_4517);
nand U4651 (N_4651,N_4459,N_4433);
nor U4652 (N_4652,N_4468,N_4560);
nor U4653 (N_4653,N_4565,N_4492);
or U4654 (N_4654,N_4487,N_4544);
nand U4655 (N_4655,N_4562,N_4591);
nand U4656 (N_4656,N_4500,N_4518);
nor U4657 (N_4657,N_4581,N_4530);
and U4658 (N_4658,N_4431,N_4482);
nand U4659 (N_4659,N_4425,N_4527);
nor U4660 (N_4660,N_4528,N_4548);
xor U4661 (N_4661,N_4413,N_4529);
and U4662 (N_4662,N_4474,N_4466);
and U4663 (N_4663,N_4488,N_4402);
nor U4664 (N_4664,N_4465,N_4594);
nand U4665 (N_4665,N_4450,N_4491);
and U4666 (N_4666,N_4440,N_4568);
xor U4667 (N_4667,N_4477,N_4567);
nor U4668 (N_4668,N_4537,N_4572);
and U4669 (N_4669,N_4504,N_4446);
and U4670 (N_4670,N_4439,N_4515);
and U4671 (N_4671,N_4478,N_4471);
and U4672 (N_4672,N_4524,N_4485);
and U4673 (N_4673,N_4542,N_4422);
nor U4674 (N_4674,N_4551,N_4486);
nand U4675 (N_4675,N_4499,N_4481);
nand U4676 (N_4676,N_4514,N_4587);
nand U4677 (N_4677,N_4456,N_4410);
or U4678 (N_4678,N_4429,N_4532);
or U4679 (N_4679,N_4479,N_4409);
and U4680 (N_4680,N_4522,N_4404);
nand U4681 (N_4681,N_4420,N_4558);
and U4682 (N_4682,N_4443,N_4411);
and U4683 (N_4683,N_4533,N_4430);
and U4684 (N_4684,N_4571,N_4501);
nand U4685 (N_4685,N_4447,N_4449);
nor U4686 (N_4686,N_4432,N_4437);
and U4687 (N_4687,N_4512,N_4403);
or U4688 (N_4688,N_4508,N_4496);
or U4689 (N_4689,N_4483,N_4511);
nor U4690 (N_4690,N_4577,N_4421);
nor U4691 (N_4691,N_4543,N_4564);
and U4692 (N_4692,N_4441,N_4503);
or U4693 (N_4693,N_4589,N_4463);
or U4694 (N_4694,N_4435,N_4426);
and U4695 (N_4695,N_4473,N_4455);
and U4696 (N_4696,N_4458,N_4417);
nand U4697 (N_4697,N_4557,N_4484);
nor U4698 (N_4698,N_4472,N_4507);
and U4699 (N_4699,N_4452,N_4461);
nand U4700 (N_4700,N_4435,N_4526);
or U4701 (N_4701,N_4481,N_4461);
and U4702 (N_4702,N_4422,N_4425);
nor U4703 (N_4703,N_4546,N_4566);
or U4704 (N_4704,N_4413,N_4522);
nand U4705 (N_4705,N_4571,N_4556);
xnor U4706 (N_4706,N_4440,N_4500);
and U4707 (N_4707,N_4565,N_4464);
and U4708 (N_4708,N_4547,N_4506);
nand U4709 (N_4709,N_4418,N_4550);
nand U4710 (N_4710,N_4486,N_4476);
and U4711 (N_4711,N_4438,N_4474);
or U4712 (N_4712,N_4470,N_4444);
nand U4713 (N_4713,N_4461,N_4450);
nand U4714 (N_4714,N_4572,N_4599);
nor U4715 (N_4715,N_4502,N_4506);
nand U4716 (N_4716,N_4420,N_4584);
nor U4717 (N_4717,N_4587,N_4449);
and U4718 (N_4718,N_4429,N_4541);
nand U4719 (N_4719,N_4532,N_4433);
and U4720 (N_4720,N_4479,N_4593);
or U4721 (N_4721,N_4590,N_4545);
xor U4722 (N_4722,N_4411,N_4511);
nor U4723 (N_4723,N_4598,N_4402);
nand U4724 (N_4724,N_4445,N_4434);
nand U4725 (N_4725,N_4537,N_4599);
and U4726 (N_4726,N_4471,N_4445);
xor U4727 (N_4727,N_4570,N_4459);
or U4728 (N_4728,N_4515,N_4442);
or U4729 (N_4729,N_4483,N_4430);
and U4730 (N_4730,N_4449,N_4450);
xnor U4731 (N_4731,N_4435,N_4548);
or U4732 (N_4732,N_4478,N_4431);
nor U4733 (N_4733,N_4404,N_4537);
nor U4734 (N_4734,N_4441,N_4457);
or U4735 (N_4735,N_4593,N_4509);
and U4736 (N_4736,N_4470,N_4560);
and U4737 (N_4737,N_4417,N_4442);
and U4738 (N_4738,N_4465,N_4501);
nand U4739 (N_4739,N_4586,N_4451);
nand U4740 (N_4740,N_4515,N_4496);
nor U4741 (N_4741,N_4502,N_4427);
and U4742 (N_4742,N_4532,N_4527);
nand U4743 (N_4743,N_4563,N_4481);
nor U4744 (N_4744,N_4565,N_4548);
or U4745 (N_4745,N_4442,N_4490);
or U4746 (N_4746,N_4473,N_4429);
and U4747 (N_4747,N_4573,N_4489);
and U4748 (N_4748,N_4438,N_4492);
and U4749 (N_4749,N_4448,N_4459);
and U4750 (N_4750,N_4520,N_4429);
nor U4751 (N_4751,N_4423,N_4487);
nand U4752 (N_4752,N_4541,N_4519);
and U4753 (N_4753,N_4538,N_4510);
nand U4754 (N_4754,N_4597,N_4438);
or U4755 (N_4755,N_4578,N_4415);
or U4756 (N_4756,N_4508,N_4468);
nand U4757 (N_4757,N_4474,N_4412);
nor U4758 (N_4758,N_4418,N_4405);
and U4759 (N_4759,N_4513,N_4539);
and U4760 (N_4760,N_4566,N_4521);
xor U4761 (N_4761,N_4564,N_4469);
or U4762 (N_4762,N_4547,N_4465);
and U4763 (N_4763,N_4498,N_4596);
nor U4764 (N_4764,N_4503,N_4464);
or U4765 (N_4765,N_4587,N_4447);
nor U4766 (N_4766,N_4437,N_4500);
nand U4767 (N_4767,N_4466,N_4449);
and U4768 (N_4768,N_4583,N_4482);
and U4769 (N_4769,N_4470,N_4488);
nor U4770 (N_4770,N_4510,N_4568);
or U4771 (N_4771,N_4517,N_4450);
nor U4772 (N_4772,N_4538,N_4578);
and U4773 (N_4773,N_4501,N_4574);
or U4774 (N_4774,N_4401,N_4581);
nor U4775 (N_4775,N_4550,N_4421);
nor U4776 (N_4776,N_4540,N_4533);
nand U4777 (N_4777,N_4470,N_4435);
nor U4778 (N_4778,N_4557,N_4552);
and U4779 (N_4779,N_4569,N_4533);
or U4780 (N_4780,N_4588,N_4492);
and U4781 (N_4781,N_4532,N_4581);
or U4782 (N_4782,N_4524,N_4406);
and U4783 (N_4783,N_4457,N_4551);
nand U4784 (N_4784,N_4573,N_4484);
nand U4785 (N_4785,N_4546,N_4452);
nand U4786 (N_4786,N_4551,N_4597);
xor U4787 (N_4787,N_4425,N_4476);
nor U4788 (N_4788,N_4461,N_4503);
nand U4789 (N_4789,N_4435,N_4510);
or U4790 (N_4790,N_4427,N_4433);
and U4791 (N_4791,N_4491,N_4543);
nand U4792 (N_4792,N_4464,N_4447);
nor U4793 (N_4793,N_4414,N_4541);
or U4794 (N_4794,N_4568,N_4402);
and U4795 (N_4795,N_4510,N_4526);
and U4796 (N_4796,N_4475,N_4533);
and U4797 (N_4797,N_4462,N_4473);
and U4798 (N_4798,N_4438,N_4525);
nor U4799 (N_4799,N_4427,N_4417);
and U4800 (N_4800,N_4655,N_4683);
nand U4801 (N_4801,N_4690,N_4774);
and U4802 (N_4802,N_4737,N_4753);
nand U4803 (N_4803,N_4799,N_4705);
and U4804 (N_4804,N_4756,N_4782);
nor U4805 (N_4805,N_4758,N_4648);
nand U4806 (N_4806,N_4712,N_4744);
or U4807 (N_4807,N_4671,N_4669);
nand U4808 (N_4808,N_4791,N_4786);
or U4809 (N_4809,N_4779,N_4717);
nand U4810 (N_4810,N_4747,N_4685);
or U4811 (N_4811,N_4738,N_4619);
nor U4812 (N_4812,N_4749,N_4759);
and U4813 (N_4813,N_4755,N_4620);
nand U4814 (N_4814,N_4780,N_4639);
and U4815 (N_4815,N_4664,N_4636);
or U4816 (N_4816,N_4617,N_4667);
nand U4817 (N_4817,N_4634,N_4661);
nor U4818 (N_4818,N_4703,N_4697);
or U4819 (N_4819,N_4775,N_4650);
or U4820 (N_4820,N_4610,N_4686);
nor U4821 (N_4821,N_4768,N_4647);
or U4822 (N_4822,N_4784,N_4675);
nand U4823 (N_4823,N_4743,N_4644);
or U4824 (N_4824,N_4613,N_4777);
nand U4825 (N_4825,N_4761,N_4704);
and U4826 (N_4826,N_4623,N_4602);
and U4827 (N_4827,N_4735,N_4673);
nor U4828 (N_4828,N_4702,N_4766);
nand U4829 (N_4829,N_4689,N_4770);
nor U4830 (N_4830,N_4733,N_4792);
nand U4831 (N_4831,N_4662,N_4652);
and U4832 (N_4832,N_4646,N_4767);
and U4833 (N_4833,N_4722,N_4754);
nor U4834 (N_4834,N_4600,N_4611);
and U4835 (N_4835,N_4640,N_4760);
and U4836 (N_4836,N_4773,N_4656);
or U4837 (N_4837,N_4778,N_4696);
and U4838 (N_4838,N_4668,N_4765);
and U4839 (N_4839,N_4763,N_4790);
nand U4840 (N_4840,N_4762,N_4627);
nand U4841 (N_4841,N_4726,N_4658);
nand U4842 (N_4842,N_4734,N_4681);
nor U4843 (N_4843,N_4659,N_4614);
nor U4844 (N_4844,N_4706,N_4701);
nand U4845 (N_4845,N_4793,N_4785);
nor U4846 (N_4846,N_4653,N_4699);
and U4847 (N_4847,N_4630,N_4641);
or U4848 (N_4848,N_4693,N_4707);
or U4849 (N_4849,N_4657,N_4632);
nand U4850 (N_4850,N_4727,N_4772);
nand U4851 (N_4851,N_4710,N_4688);
nand U4852 (N_4852,N_4750,N_4781);
nand U4853 (N_4853,N_4783,N_4679);
and U4854 (N_4854,N_4748,N_4720);
nor U4855 (N_4855,N_4628,N_4731);
nor U4856 (N_4856,N_4642,N_4609);
or U4857 (N_4857,N_4626,N_4622);
nand U4858 (N_4858,N_4666,N_4752);
nand U4859 (N_4859,N_4631,N_4618);
and U4860 (N_4860,N_4607,N_4612);
nand U4861 (N_4861,N_4719,N_4643);
nand U4862 (N_4862,N_4601,N_4740);
and U4863 (N_4863,N_4678,N_4721);
nor U4864 (N_4864,N_4660,N_4687);
nor U4865 (N_4865,N_4637,N_4670);
nand U4866 (N_4866,N_4716,N_4608);
or U4867 (N_4867,N_4715,N_4709);
nor U4868 (N_4868,N_4729,N_4708);
nand U4869 (N_4869,N_4723,N_4672);
nor U4870 (N_4870,N_4771,N_4789);
or U4871 (N_4871,N_4732,N_4684);
and U4872 (N_4872,N_4746,N_4621);
and U4873 (N_4873,N_4682,N_4680);
nand U4874 (N_4874,N_4604,N_4757);
or U4875 (N_4875,N_4700,N_4788);
or U4876 (N_4876,N_4776,N_4714);
nor U4877 (N_4877,N_4713,N_4724);
nand U4878 (N_4878,N_4798,N_4730);
nor U4879 (N_4879,N_4645,N_4694);
nor U4880 (N_4880,N_4692,N_4654);
or U4881 (N_4881,N_4624,N_4797);
nand U4882 (N_4882,N_4665,N_4676);
and U4883 (N_4883,N_4649,N_4769);
nor U4884 (N_4884,N_4638,N_4677);
or U4885 (N_4885,N_4651,N_4796);
and U4886 (N_4886,N_4728,N_4711);
nand U4887 (N_4887,N_4674,N_4718);
nand U4888 (N_4888,N_4625,N_4725);
nand U4889 (N_4889,N_4698,N_4794);
nand U4890 (N_4890,N_4616,N_4741);
and U4891 (N_4891,N_4691,N_4603);
and U4892 (N_4892,N_4605,N_4739);
and U4893 (N_4893,N_4751,N_4663);
or U4894 (N_4894,N_4742,N_4764);
and U4895 (N_4895,N_4606,N_4795);
xor U4896 (N_4896,N_4695,N_4635);
nand U4897 (N_4897,N_4787,N_4736);
and U4898 (N_4898,N_4633,N_4615);
nand U4899 (N_4899,N_4745,N_4629);
nor U4900 (N_4900,N_4677,N_4657);
nand U4901 (N_4901,N_4634,N_4672);
and U4902 (N_4902,N_4614,N_4690);
and U4903 (N_4903,N_4693,N_4695);
nand U4904 (N_4904,N_4778,N_4785);
or U4905 (N_4905,N_4758,N_4686);
or U4906 (N_4906,N_4710,N_4702);
or U4907 (N_4907,N_4679,N_4779);
or U4908 (N_4908,N_4653,N_4613);
and U4909 (N_4909,N_4669,N_4607);
nand U4910 (N_4910,N_4634,N_4612);
nand U4911 (N_4911,N_4638,N_4655);
or U4912 (N_4912,N_4762,N_4647);
nor U4913 (N_4913,N_4605,N_4675);
nor U4914 (N_4914,N_4674,N_4737);
or U4915 (N_4915,N_4695,N_4687);
and U4916 (N_4916,N_4714,N_4716);
or U4917 (N_4917,N_4652,N_4694);
and U4918 (N_4918,N_4713,N_4664);
or U4919 (N_4919,N_4706,N_4767);
nand U4920 (N_4920,N_4646,N_4609);
and U4921 (N_4921,N_4689,N_4723);
and U4922 (N_4922,N_4707,N_4747);
nor U4923 (N_4923,N_4703,N_4708);
or U4924 (N_4924,N_4781,N_4701);
or U4925 (N_4925,N_4705,N_4655);
or U4926 (N_4926,N_4624,N_4670);
nor U4927 (N_4927,N_4673,N_4749);
nor U4928 (N_4928,N_4680,N_4711);
nand U4929 (N_4929,N_4712,N_4753);
and U4930 (N_4930,N_4639,N_4609);
and U4931 (N_4931,N_4677,N_4651);
nand U4932 (N_4932,N_4750,N_4647);
or U4933 (N_4933,N_4718,N_4749);
or U4934 (N_4934,N_4655,N_4652);
nor U4935 (N_4935,N_4768,N_4727);
or U4936 (N_4936,N_4688,N_4709);
nand U4937 (N_4937,N_4666,N_4727);
nor U4938 (N_4938,N_4649,N_4663);
nor U4939 (N_4939,N_4627,N_4692);
nand U4940 (N_4940,N_4602,N_4700);
and U4941 (N_4941,N_4623,N_4619);
and U4942 (N_4942,N_4634,N_4674);
and U4943 (N_4943,N_4620,N_4625);
and U4944 (N_4944,N_4671,N_4658);
nand U4945 (N_4945,N_4641,N_4640);
or U4946 (N_4946,N_4744,N_4703);
nand U4947 (N_4947,N_4738,N_4791);
or U4948 (N_4948,N_4726,N_4679);
nand U4949 (N_4949,N_4736,N_4738);
or U4950 (N_4950,N_4695,N_4634);
xnor U4951 (N_4951,N_4631,N_4728);
and U4952 (N_4952,N_4771,N_4761);
and U4953 (N_4953,N_4625,N_4793);
nor U4954 (N_4954,N_4738,N_4795);
and U4955 (N_4955,N_4644,N_4712);
nor U4956 (N_4956,N_4672,N_4679);
or U4957 (N_4957,N_4623,N_4620);
and U4958 (N_4958,N_4680,N_4622);
and U4959 (N_4959,N_4692,N_4647);
xnor U4960 (N_4960,N_4754,N_4705);
nor U4961 (N_4961,N_4771,N_4694);
nor U4962 (N_4962,N_4638,N_4651);
nand U4963 (N_4963,N_4653,N_4616);
and U4964 (N_4964,N_4656,N_4637);
and U4965 (N_4965,N_4675,N_4748);
and U4966 (N_4966,N_4776,N_4766);
or U4967 (N_4967,N_4737,N_4638);
and U4968 (N_4968,N_4632,N_4736);
or U4969 (N_4969,N_4751,N_4607);
xnor U4970 (N_4970,N_4663,N_4757);
nor U4971 (N_4971,N_4633,N_4756);
or U4972 (N_4972,N_4632,N_4771);
or U4973 (N_4973,N_4615,N_4686);
nand U4974 (N_4974,N_4767,N_4734);
nand U4975 (N_4975,N_4753,N_4719);
and U4976 (N_4976,N_4614,N_4752);
nor U4977 (N_4977,N_4747,N_4777);
or U4978 (N_4978,N_4683,N_4757);
and U4979 (N_4979,N_4630,N_4683);
nand U4980 (N_4980,N_4678,N_4626);
and U4981 (N_4981,N_4671,N_4688);
nand U4982 (N_4982,N_4741,N_4602);
nand U4983 (N_4983,N_4634,N_4705);
nor U4984 (N_4984,N_4708,N_4725);
or U4985 (N_4985,N_4651,N_4794);
nand U4986 (N_4986,N_4626,N_4614);
or U4987 (N_4987,N_4798,N_4759);
nor U4988 (N_4988,N_4753,N_4656);
nor U4989 (N_4989,N_4613,N_4798);
or U4990 (N_4990,N_4670,N_4674);
nand U4991 (N_4991,N_4687,N_4666);
and U4992 (N_4992,N_4652,N_4780);
and U4993 (N_4993,N_4688,N_4796);
or U4994 (N_4994,N_4667,N_4770);
nand U4995 (N_4995,N_4683,N_4604);
or U4996 (N_4996,N_4637,N_4660);
nand U4997 (N_4997,N_4618,N_4628);
nor U4998 (N_4998,N_4614,N_4798);
and U4999 (N_4999,N_4789,N_4696);
or U5000 (N_5000,N_4863,N_4806);
and U5001 (N_5001,N_4994,N_4985);
nand U5002 (N_5002,N_4932,N_4803);
nor U5003 (N_5003,N_4812,N_4824);
nor U5004 (N_5004,N_4908,N_4989);
nand U5005 (N_5005,N_4838,N_4851);
nor U5006 (N_5006,N_4813,N_4894);
nor U5007 (N_5007,N_4849,N_4886);
or U5008 (N_5008,N_4842,N_4900);
or U5009 (N_5009,N_4925,N_4912);
or U5010 (N_5010,N_4976,N_4967);
nand U5011 (N_5011,N_4998,N_4896);
nor U5012 (N_5012,N_4960,N_4893);
xnor U5013 (N_5013,N_4841,N_4870);
xor U5014 (N_5014,N_4918,N_4930);
or U5015 (N_5015,N_4866,N_4897);
and U5016 (N_5016,N_4802,N_4901);
or U5017 (N_5017,N_4904,N_4865);
or U5018 (N_5018,N_4862,N_4935);
nand U5019 (N_5019,N_4883,N_4956);
xnor U5020 (N_5020,N_4833,N_4971);
nor U5021 (N_5021,N_4881,N_4853);
or U5022 (N_5022,N_4882,N_4855);
or U5023 (N_5023,N_4926,N_4848);
and U5024 (N_5024,N_4915,N_4969);
nor U5025 (N_5025,N_4857,N_4987);
and U5026 (N_5026,N_4801,N_4839);
nand U5027 (N_5027,N_4950,N_4871);
nand U5028 (N_5028,N_4949,N_4906);
xor U5029 (N_5029,N_4905,N_4809);
and U5030 (N_5030,N_4816,N_4939);
nor U5031 (N_5031,N_4843,N_4903);
nor U5032 (N_5032,N_4829,N_4872);
nor U5033 (N_5033,N_4811,N_4920);
and U5034 (N_5034,N_4953,N_4810);
and U5035 (N_5035,N_4819,N_4840);
nor U5036 (N_5036,N_4965,N_4919);
or U5037 (N_5037,N_4937,N_4888);
nand U5038 (N_5038,N_4814,N_4910);
nor U5039 (N_5039,N_4879,N_4979);
nand U5040 (N_5040,N_4907,N_4974);
or U5041 (N_5041,N_4968,N_4899);
nor U5042 (N_5042,N_4972,N_4982);
and U5043 (N_5043,N_4827,N_4807);
nor U5044 (N_5044,N_4875,N_4929);
nand U5045 (N_5045,N_4938,N_4885);
or U5046 (N_5046,N_4981,N_4852);
and U5047 (N_5047,N_4957,N_4942);
and U5048 (N_5048,N_4847,N_4946);
and U5049 (N_5049,N_4876,N_4992);
and U5050 (N_5050,N_4820,N_4948);
or U5051 (N_5051,N_4996,N_4913);
and U5052 (N_5052,N_4983,N_4878);
nand U5053 (N_5053,N_4858,N_4993);
or U5054 (N_5054,N_4954,N_4951);
nor U5055 (N_5055,N_4832,N_4856);
and U5056 (N_5056,N_4868,N_4952);
nor U5057 (N_5057,N_4818,N_4975);
or U5058 (N_5058,N_4836,N_4933);
or U5059 (N_5059,N_4823,N_4995);
xor U5060 (N_5060,N_4944,N_4831);
and U5061 (N_5061,N_4889,N_4964);
and U5062 (N_5062,N_4854,N_4923);
nand U5063 (N_5063,N_4860,N_4887);
nand U5064 (N_5064,N_4861,N_4928);
nor U5065 (N_5065,N_4850,N_4980);
nand U5066 (N_5066,N_4911,N_4970);
nor U5067 (N_5067,N_4845,N_4837);
and U5068 (N_5068,N_4834,N_4963);
and U5069 (N_5069,N_4941,N_4997);
nand U5070 (N_5070,N_4943,N_4988);
xor U5071 (N_5071,N_4961,N_4815);
nand U5072 (N_5072,N_4895,N_4927);
nor U5073 (N_5073,N_4826,N_4955);
nand U5074 (N_5074,N_4914,N_4877);
nand U5075 (N_5075,N_4817,N_4821);
and U5076 (N_5076,N_4804,N_4880);
or U5077 (N_5077,N_4867,N_4859);
and U5078 (N_5078,N_4909,N_4945);
nor U5079 (N_5079,N_4800,N_4966);
or U5080 (N_5080,N_4835,N_4978);
nand U5081 (N_5081,N_4891,N_4916);
and U5082 (N_5082,N_4890,N_4844);
xnor U5083 (N_5083,N_4984,N_4917);
or U5084 (N_5084,N_4864,N_4999);
and U5085 (N_5085,N_4958,N_4991);
and U5086 (N_5086,N_4805,N_4898);
or U5087 (N_5087,N_4892,N_4884);
and U5088 (N_5088,N_4990,N_4936);
and U5089 (N_5089,N_4846,N_4874);
nor U5090 (N_5090,N_4977,N_4830);
and U5091 (N_5091,N_4947,N_4828);
or U5092 (N_5092,N_4931,N_4825);
and U5093 (N_5093,N_4902,N_4873);
nand U5094 (N_5094,N_4934,N_4808);
nor U5095 (N_5095,N_4959,N_4924);
nor U5096 (N_5096,N_4986,N_4922);
and U5097 (N_5097,N_4869,N_4921);
and U5098 (N_5098,N_4822,N_4962);
and U5099 (N_5099,N_4973,N_4940);
xnor U5100 (N_5100,N_4871,N_4903);
nand U5101 (N_5101,N_4980,N_4862);
nor U5102 (N_5102,N_4825,N_4908);
and U5103 (N_5103,N_4817,N_4880);
nand U5104 (N_5104,N_4819,N_4823);
and U5105 (N_5105,N_4894,N_4952);
nand U5106 (N_5106,N_4993,N_4801);
and U5107 (N_5107,N_4875,N_4963);
or U5108 (N_5108,N_4974,N_4843);
nor U5109 (N_5109,N_4971,N_4835);
nand U5110 (N_5110,N_4818,N_4849);
nand U5111 (N_5111,N_4913,N_4819);
or U5112 (N_5112,N_4928,N_4866);
and U5113 (N_5113,N_4962,N_4850);
or U5114 (N_5114,N_4994,N_4911);
xnor U5115 (N_5115,N_4989,N_4999);
nand U5116 (N_5116,N_4813,N_4940);
or U5117 (N_5117,N_4900,N_4994);
or U5118 (N_5118,N_4872,N_4886);
or U5119 (N_5119,N_4882,N_4821);
nand U5120 (N_5120,N_4895,N_4801);
nand U5121 (N_5121,N_4952,N_4816);
and U5122 (N_5122,N_4836,N_4828);
and U5123 (N_5123,N_4893,N_4849);
or U5124 (N_5124,N_4987,N_4900);
nand U5125 (N_5125,N_4868,N_4807);
or U5126 (N_5126,N_4968,N_4983);
xor U5127 (N_5127,N_4982,N_4870);
nor U5128 (N_5128,N_4952,N_4878);
and U5129 (N_5129,N_4862,N_4857);
and U5130 (N_5130,N_4919,N_4809);
or U5131 (N_5131,N_4850,N_4921);
or U5132 (N_5132,N_4844,N_4835);
and U5133 (N_5133,N_4966,N_4828);
and U5134 (N_5134,N_4939,N_4854);
and U5135 (N_5135,N_4966,N_4922);
or U5136 (N_5136,N_4824,N_4914);
nand U5137 (N_5137,N_4818,N_4860);
nand U5138 (N_5138,N_4943,N_4864);
or U5139 (N_5139,N_4908,N_4821);
nor U5140 (N_5140,N_4839,N_4963);
nand U5141 (N_5141,N_4802,N_4896);
nand U5142 (N_5142,N_4893,N_4814);
or U5143 (N_5143,N_4901,N_4918);
nor U5144 (N_5144,N_4967,N_4982);
nand U5145 (N_5145,N_4903,N_4816);
and U5146 (N_5146,N_4939,N_4974);
and U5147 (N_5147,N_4849,N_4973);
or U5148 (N_5148,N_4845,N_4959);
nor U5149 (N_5149,N_4974,N_4893);
and U5150 (N_5150,N_4912,N_4899);
and U5151 (N_5151,N_4930,N_4910);
and U5152 (N_5152,N_4951,N_4823);
nand U5153 (N_5153,N_4929,N_4808);
and U5154 (N_5154,N_4820,N_4842);
and U5155 (N_5155,N_4831,N_4958);
or U5156 (N_5156,N_4976,N_4853);
xor U5157 (N_5157,N_4807,N_4968);
or U5158 (N_5158,N_4963,N_4934);
and U5159 (N_5159,N_4987,N_4956);
or U5160 (N_5160,N_4907,N_4971);
or U5161 (N_5161,N_4936,N_4953);
xnor U5162 (N_5162,N_4962,N_4868);
or U5163 (N_5163,N_4996,N_4829);
nor U5164 (N_5164,N_4902,N_4863);
nor U5165 (N_5165,N_4838,N_4968);
nand U5166 (N_5166,N_4899,N_4827);
nand U5167 (N_5167,N_4959,N_4979);
and U5168 (N_5168,N_4895,N_4994);
and U5169 (N_5169,N_4845,N_4974);
nand U5170 (N_5170,N_4948,N_4989);
xnor U5171 (N_5171,N_4943,N_4802);
nor U5172 (N_5172,N_4932,N_4807);
nand U5173 (N_5173,N_4851,N_4974);
nor U5174 (N_5174,N_4894,N_4847);
nand U5175 (N_5175,N_4843,N_4924);
nor U5176 (N_5176,N_4905,N_4912);
nor U5177 (N_5177,N_4845,N_4856);
nand U5178 (N_5178,N_4973,N_4845);
nor U5179 (N_5179,N_4816,N_4973);
nor U5180 (N_5180,N_4907,N_4988);
nor U5181 (N_5181,N_4891,N_4979);
nor U5182 (N_5182,N_4822,N_4804);
nand U5183 (N_5183,N_4882,N_4998);
or U5184 (N_5184,N_4967,N_4856);
xnor U5185 (N_5185,N_4959,N_4922);
or U5186 (N_5186,N_4959,N_4943);
nand U5187 (N_5187,N_4828,N_4951);
nor U5188 (N_5188,N_4895,N_4896);
and U5189 (N_5189,N_4905,N_4877);
nand U5190 (N_5190,N_4956,N_4865);
or U5191 (N_5191,N_4989,N_4974);
nand U5192 (N_5192,N_4853,N_4994);
nand U5193 (N_5193,N_4986,N_4907);
nor U5194 (N_5194,N_4882,N_4909);
nor U5195 (N_5195,N_4977,N_4835);
nor U5196 (N_5196,N_4820,N_4953);
and U5197 (N_5197,N_4930,N_4964);
or U5198 (N_5198,N_4890,N_4873);
nand U5199 (N_5199,N_4848,N_4832);
or U5200 (N_5200,N_5171,N_5194);
nand U5201 (N_5201,N_5067,N_5007);
and U5202 (N_5202,N_5142,N_5018);
xor U5203 (N_5203,N_5056,N_5003);
nor U5204 (N_5204,N_5150,N_5042);
and U5205 (N_5205,N_5006,N_5137);
or U5206 (N_5206,N_5039,N_5141);
or U5207 (N_5207,N_5157,N_5099);
nand U5208 (N_5208,N_5159,N_5162);
or U5209 (N_5209,N_5183,N_5103);
and U5210 (N_5210,N_5176,N_5084);
nand U5211 (N_5211,N_5189,N_5034);
and U5212 (N_5212,N_5048,N_5188);
nor U5213 (N_5213,N_5119,N_5163);
and U5214 (N_5214,N_5116,N_5181);
nor U5215 (N_5215,N_5186,N_5173);
nor U5216 (N_5216,N_5120,N_5112);
xor U5217 (N_5217,N_5136,N_5088);
nor U5218 (N_5218,N_5132,N_5149);
nor U5219 (N_5219,N_5031,N_5182);
nand U5220 (N_5220,N_5148,N_5062);
nand U5221 (N_5221,N_5168,N_5140);
nand U5222 (N_5222,N_5082,N_5087);
or U5223 (N_5223,N_5178,N_5107);
nor U5224 (N_5224,N_5123,N_5059);
or U5225 (N_5225,N_5009,N_5066);
and U5226 (N_5226,N_5055,N_5109);
xnor U5227 (N_5227,N_5094,N_5156);
nand U5228 (N_5228,N_5046,N_5061);
or U5229 (N_5229,N_5012,N_5036);
or U5230 (N_5230,N_5069,N_5097);
or U5231 (N_5231,N_5135,N_5170);
or U5232 (N_5232,N_5072,N_5106);
and U5233 (N_5233,N_5199,N_5032);
nor U5234 (N_5234,N_5030,N_5124);
and U5235 (N_5235,N_5093,N_5079);
and U5236 (N_5236,N_5058,N_5133);
nor U5237 (N_5237,N_5045,N_5198);
nand U5238 (N_5238,N_5013,N_5005);
or U5239 (N_5239,N_5144,N_5022);
and U5240 (N_5240,N_5001,N_5101);
nand U5241 (N_5241,N_5083,N_5029);
or U5242 (N_5242,N_5158,N_5020);
nor U5243 (N_5243,N_5028,N_5065);
nand U5244 (N_5244,N_5037,N_5008);
nor U5245 (N_5245,N_5060,N_5152);
or U5246 (N_5246,N_5169,N_5117);
nor U5247 (N_5247,N_5160,N_5113);
nand U5248 (N_5248,N_5075,N_5151);
or U5249 (N_5249,N_5090,N_5121);
or U5250 (N_5250,N_5078,N_5044);
and U5251 (N_5251,N_5098,N_5187);
and U5252 (N_5252,N_5196,N_5184);
nor U5253 (N_5253,N_5038,N_5010);
nand U5254 (N_5254,N_5128,N_5179);
and U5255 (N_5255,N_5175,N_5115);
or U5256 (N_5256,N_5091,N_5105);
nand U5257 (N_5257,N_5050,N_5143);
nor U5258 (N_5258,N_5153,N_5051);
nand U5259 (N_5259,N_5043,N_5025);
nor U5260 (N_5260,N_5076,N_5023);
and U5261 (N_5261,N_5054,N_5096);
nor U5262 (N_5262,N_5127,N_5195);
or U5263 (N_5263,N_5011,N_5193);
or U5264 (N_5264,N_5111,N_5154);
and U5265 (N_5265,N_5114,N_5161);
and U5266 (N_5266,N_5027,N_5130);
nand U5267 (N_5267,N_5166,N_5064);
and U5268 (N_5268,N_5014,N_5167);
or U5269 (N_5269,N_5073,N_5068);
nor U5270 (N_5270,N_5100,N_5164);
nand U5271 (N_5271,N_5102,N_5145);
nor U5272 (N_5272,N_5089,N_5104);
or U5273 (N_5273,N_5172,N_5165);
and U5274 (N_5274,N_5074,N_5155);
nand U5275 (N_5275,N_5125,N_5019);
or U5276 (N_5276,N_5035,N_5017);
or U5277 (N_5277,N_5126,N_5118);
or U5278 (N_5278,N_5057,N_5002);
or U5279 (N_5279,N_5081,N_5021);
or U5280 (N_5280,N_5015,N_5053);
nand U5281 (N_5281,N_5146,N_5000);
or U5282 (N_5282,N_5049,N_5177);
nand U5283 (N_5283,N_5185,N_5129);
nand U5284 (N_5284,N_5070,N_5180);
nand U5285 (N_5285,N_5122,N_5063);
nor U5286 (N_5286,N_5052,N_5086);
or U5287 (N_5287,N_5033,N_5174);
or U5288 (N_5288,N_5139,N_5110);
or U5289 (N_5289,N_5026,N_5131);
xor U5290 (N_5290,N_5040,N_5138);
and U5291 (N_5291,N_5095,N_5071);
nand U5292 (N_5292,N_5004,N_5077);
or U5293 (N_5293,N_5134,N_5085);
or U5294 (N_5294,N_5147,N_5191);
nor U5295 (N_5295,N_5190,N_5047);
and U5296 (N_5296,N_5080,N_5192);
or U5297 (N_5297,N_5108,N_5092);
or U5298 (N_5298,N_5016,N_5024);
or U5299 (N_5299,N_5197,N_5041);
nand U5300 (N_5300,N_5054,N_5139);
or U5301 (N_5301,N_5107,N_5011);
and U5302 (N_5302,N_5069,N_5046);
nor U5303 (N_5303,N_5017,N_5167);
and U5304 (N_5304,N_5083,N_5078);
or U5305 (N_5305,N_5124,N_5074);
nand U5306 (N_5306,N_5132,N_5145);
xor U5307 (N_5307,N_5193,N_5038);
nand U5308 (N_5308,N_5044,N_5188);
nand U5309 (N_5309,N_5095,N_5162);
and U5310 (N_5310,N_5188,N_5183);
nand U5311 (N_5311,N_5106,N_5147);
nand U5312 (N_5312,N_5135,N_5187);
and U5313 (N_5313,N_5008,N_5087);
and U5314 (N_5314,N_5170,N_5125);
nor U5315 (N_5315,N_5085,N_5179);
nor U5316 (N_5316,N_5109,N_5043);
nor U5317 (N_5317,N_5159,N_5183);
nor U5318 (N_5318,N_5071,N_5073);
or U5319 (N_5319,N_5193,N_5196);
nand U5320 (N_5320,N_5130,N_5066);
nor U5321 (N_5321,N_5105,N_5082);
nor U5322 (N_5322,N_5007,N_5073);
and U5323 (N_5323,N_5019,N_5156);
and U5324 (N_5324,N_5178,N_5104);
and U5325 (N_5325,N_5033,N_5163);
and U5326 (N_5326,N_5006,N_5001);
and U5327 (N_5327,N_5108,N_5194);
nor U5328 (N_5328,N_5175,N_5186);
or U5329 (N_5329,N_5108,N_5056);
xor U5330 (N_5330,N_5087,N_5127);
nor U5331 (N_5331,N_5106,N_5121);
nand U5332 (N_5332,N_5185,N_5155);
nor U5333 (N_5333,N_5012,N_5119);
and U5334 (N_5334,N_5175,N_5018);
nor U5335 (N_5335,N_5084,N_5057);
nand U5336 (N_5336,N_5104,N_5057);
nand U5337 (N_5337,N_5184,N_5016);
nand U5338 (N_5338,N_5037,N_5080);
or U5339 (N_5339,N_5113,N_5097);
nand U5340 (N_5340,N_5192,N_5018);
nand U5341 (N_5341,N_5160,N_5173);
or U5342 (N_5342,N_5054,N_5005);
or U5343 (N_5343,N_5163,N_5133);
nand U5344 (N_5344,N_5016,N_5080);
nand U5345 (N_5345,N_5096,N_5065);
xnor U5346 (N_5346,N_5197,N_5018);
nand U5347 (N_5347,N_5020,N_5037);
nand U5348 (N_5348,N_5195,N_5099);
or U5349 (N_5349,N_5167,N_5010);
nand U5350 (N_5350,N_5031,N_5160);
nand U5351 (N_5351,N_5100,N_5114);
or U5352 (N_5352,N_5197,N_5111);
nor U5353 (N_5353,N_5066,N_5113);
or U5354 (N_5354,N_5182,N_5134);
nand U5355 (N_5355,N_5079,N_5135);
nand U5356 (N_5356,N_5174,N_5113);
nand U5357 (N_5357,N_5079,N_5053);
nand U5358 (N_5358,N_5024,N_5026);
nand U5359 (N_5359,N_5193,N_5097);
or U5360 (N_5360,N_5191,N_5029);
nand U5361 (N_5361,N_5132,N_5128);
nand U5362 (N_5362,N_5178,N_5169);
or U5363 (N_5363,N_5194,N_5067);
nor U5364 (N_5364,N_5013,N_5037);
and U5365 (N_5365,N_5046,N_5005);
and U5366 (N_5366,N_5056,N_5146);
nand U5367 (N_5367,N_5103,N_5166);
nand U5368 (N_5368,N_5169,N_5019);
nor U5369 (N_5369,N_5020,N_5075);
or U5370 (N_5370,N_5054,N_5021);
nand U5371 (N_5371,N_5188,N_5110);
and U5372 (N_5372,N_5083,N_5066);
nor U5373 (N_5373,N_5198,N_5079);
and U5374 (N_5374,N_5032,N_5147);
or U5375 (N_5375,N_5117,N_5034);
and U5376 (N_5376,N_5038,N_5191);
or U5377 (N_5377,N_5114,N_5071);
and U5378 (N_5378,N_5018,N_5015);
xor U5379 (N_5379,N_5081,N_5047);
and U5380 (N_5380,N_5182,N_5140);
or U5381 (N_5381,N_5036,N_5125);
and U5382 (N_5382,N_5186,N_5038);
or U5383 (N_5383,N_5056,N_5166);
nand U5384 (N_5384,N_5192,N_5196);
and U5385 (N_5385,N_5014,N_5154);
or U5386 (N_5386,N_5041,N_5007);
nor U5387 (N_5387,N_5167,N_5041);
and U5388 (N_5388,N_5121,N_5041);
nand U5389 (N_5389,N_5035,N_5146);
nor U5390 (N_5390,N_5064,N_5044);
nor U5391 (N_5391,N_5185,N_5054);
nand U5392 (N_5392,N_5027,N_5072);
nand U5393 (N_5393,N_5170,N_5104);
and U5394 (N_5394,N_5112,N_5176);
or U5395 (N_5395,N_5046,N_5067);
nor U5396 (N_5396,N_5162,N_5098);
or U5397 (N_5397,N_5170,N_5176);
or U5398 (N_5398,N_5186,N_5134);
and U5399 (N_5399,N_5020,N_5153);
or U5400 (N_5400,N_5302,N_5269);
nand U5401 (N_5401,N_5206,N_5310);
and U5402 (N_5402,N_5303,N_5203);
nand U5403 (N_5403,N_5388,N_5225);
nand U5404 (N_5404,N_5399,N_5283);
or U5405 (N_5405,N_5292,N_5294);
nand U5406 (N_5406,N_5389,N_5274);
nand U5407 (N_5407,N_5240,N_5391);
and U5408 (N_5408,N_5208,N_5328);
and U5409 (N_5409,N_5335,N_5205);
and U5410 (N_5410,N_5390,N_5257);
nand U5411 (N_5411,N_5220,N_5248);
or U5412 (N_5412,N_5368,N_5266);
xor U5413 (N_5413,N_5288,N_5360);
nand U5414 (N_5414,N_5376,N_5231);
nand U5415 (N_5415,N_5207,N_5216);
nor U5416 (N_5416,N_5352,N_5314);
or U5417 (N_5417,N_5364,N_5222);
nand U5418 (N_5418,N_5270,N_5214);
or U5419 (N_5419,N_5276,N_5333);
or U5420 (N_5420,N_5347,N_5297);
or U5421 (N_5421,N_5379,N_5201);
or U5422 (N_5422,N_5359,N_5378);
nor U5423 (N_5423,N_5223,N_5278);
nor U5424 (N_5424,N_5271,N_5246);
and U5425 (N_5425,N_5371,N_5382);
nor U5426 (N_5426,N_5386,N_5285);
or U5427 (N_5427,N_5375,N_5210);
nor U5428 (N_5428,N_5398,N_5258);
xnor U5429 (N_5429,N_5202,N_5341);
and U5430 (N_5430,N_5373,N_5320);
nand U5431 (N_5431,N_5286,N_5357);
nor U5432 (N_5432,N_5291,N_5293);
nor U5433 (N_5433,N_5342,N_5256);
nand U5434 (N_5434,N_5301,N_5387);
or U5435 (N_5435,N_5281,N_5268);
or U5436 (N_5436,N_5372,N_5284);
or U5437 (N_5437,N_5337,N_5313);
or U5438 (N_5438,N_5321,N_5374);
or U5439 (N_5439,N_5330,N_5298);
nor U5440 (N_5440,N_5228,N_5385);
xnor U5441 (N_5441,N_5351,N_5215);
or U5442 (N_5442,N_5300,N_5353);
nor U5443 (N_5443,N_5273,N_5244);
nor U5444 (N_5444,N_5265,N_5332);
or U5445 (N_5445,N_5253,N_5394);
and U5446 (N_5446,N_5324,N_5242);
nor U5447 (N_5447,N_5249,N_5255);
nor U5448 (N_5448,N_5237,N_5326);
or U5449 (N_5449,N_5355,N_5261);
and U5450 (N_5450,N_5393,N_5272);
nor U5451 (N_5451,N_5299,N_5259);
nand U5452 (N_5452,N_5396,N_5331);
or U5453 (N_5453,N_5340,N_5280);
nand U5454 (N_5454,N_5356,N_5296);
or U5455 (N_5455,N_5343,N_5350);
xor U5456 (N_5456,N_5251,N_5224);
or U5457 (N_5457,N_5322,N_5377);
nor U5458 (N_5458,N_5317,N_5311);
or U5459 (N_5459,N_5334,N_5370);
or U5460 (N_5460,N_5312,N_5319);
and U5461 (N_5461,N_5236,N_5380);
and U5462 (N_5462,N_5212,N_5238);
nand U5463 (N_5463,N_5304,N_5229);
nor U5464 (N_5464,N_5260,N_5323);
or U5465 (N_5465,N_5366,N_5200);
or U5466 (N_5466,N_5383,N_5369);
and U5467 (N_5467,N_5218,N_5318);
xor U5468 (N_5468,N_5367,N_5289);
xor U5469 (N_5469,N_5233,N_5232);
and U5470 (N_5470,N_5363,N_5263);
or U5471 (N_5471,N_5295,N_5235);
or U5472 (N_5472,N_5250,N_5252);
or U5473 (N_5473,N_5339,N_5227);
nor U5474 (N_5474,N_5221,N_5325);
nand U5475 (N_5475,N_5279,N_5392);
or U5476 (N_5476,N_5254,N_5282);
nand U5477 (N_5477,N_5308,N_5245);
nand U5478 (N_5478,N_5316,N_5362);
or U5479 (N_5479,N_5348,N_5358);
nor U5480 (N_5480,N_5305,N_5226);
or U5481 (N_5481,N_5213,N_5397);
or U5482 (N_5482,N_5315,N_5204);
nand U5483 (N_5483,N_5384,N_5361);
and U5484 (N_5484,N_5349,N_5327);
nor U5485 (N_5485,N_5381,N_5336);
or U5486 (N_5486,N_5346,N_5365);
nand U5487 (N_5487,N_5247,N_5219);
and U5488 (N_5488,N_5338,N_5287);
nand U5489 (N_5489,N_5234,N_5306);
nand U5490 (N_5490,N_5241,N_5267);
nand U5491 (N_5491,N_5239,N_5345);
and U5492 (N_5492,N_5307,N_5262);
or U5493 (N_5493,N_5211,N_5264);
nand U5494 (N_5494,N_5329,N_5309);
or U5495 (N_5495,N_5230,N_5243);
or U5496 (N_5496,N_5275,N_5277);
or U5497 (N_5497,N_5395,N_5354);
and U5498 (N_5498,N_5209,N_5217);
nand U5499 (N_5499,N_5290,N_5344);
or U5500 (N_5500,N_5348,N_5279);
or U5501 (N_5501,N_5248,N_5387);
or U5502 (N_5502,N_5268,N_5230);
or U5503 (N_5503,N_5273,N_5251);
nor U5504 (N_5504,N_5398,N_5233);
nor U5505 (N_5505,N_5302,N_5211);
and U5506 (N_5506,N_5238,N_5216);
nand U5507 (N_5507,N_5258,N_5287);
nand U5508 (N_5508,N_5366,N_5290);
and U5509 (N_5509,N_5372,N_5311);
and U5510 (N_5510,N_5308,N_5386);
or U5511 (N_5511,N_5215,N_5346);
and U5512 (N_5512,N_5378,N_5305);
nand U5513 (N_5513,N_5206,N_5323);
and U5514 (N_5514,N_5327,N_5350);
and U5515 (N_5515,N_5227,N_5275);
and U5516 (N_5516,N_5205,N_5208);
nor U5517 (N_5517,N_5350,N_5213);
nand U5518 (N_5518,N_5329,N_5343);
or U5519 (N_5519,N_5258,N_5293);
and U5520 (N_5520,N_5284,N_5377);
nor U5521 (N_5521,N_5324,N_5288);
or U5522 (N_5522,N_5230,N_5272);
nand U5523 (N_5523,N_5363,N_5237);
and U5524 (N_5524,N_5318,N_5261);
nor U5525 (N_5525,N_5303,N_5305);
and U5526 (N_5526,N_5275,N_5314);
nor U5527 (N_5527,N_5296,N_5360);
nand U5528 (N_5528,N_5284,N_5225);
nor U5529 (N_5529,N_5241,N_5210);
or U5530 (N_5530,N_5222,N_5214);
and U5531 (N_5531,N_5380,N_5368);
or U5532 (N_5532,N_5224,N_5367);
or U5533 (N_5533,N_5338,N_5372);
nor U5534 (N_5534,N_5235,N_5339);
or U5535 (N_5535,N_5378,N_5255);
and U5536 (N_5536,N_5281,N_5274);
or U5537 (N_5537,N_5373,N_5250);
nand U5538 (N_5538,N_5313,N_5311);
and U5539 (N_5539,N_5341,N_5205);
nor U5540 (N_5540,N_5306,N_5348);
or U5541 (N_5541,N_5266,N_5339);
nand U5542 (N_5542,N_5227,N_5368);
and U5543 (N_5543,N_5227,N_5332);
nor U5544 (N_5544,N_5281,N_5370);
nor U5545 (N_5545,N_5212,N_5273);
or U5546 (N_5546,N_5331,N_5375);
nand U5547 (N_5547,N_5236,N_5223);
nand U5548 (N_5548,N_5214,N_5339);
nand U5549 (N_5549,N_5244,N_5272);
and U5550 (N_5550,N_5361,N_5258);
nand U5551 (N_5551,N_5353,N_5218);
and U5552 (N_5552,N_5353,N_5343);
nand U5553 (N_5553,N_5282,N_5338);
nand U5554 (N_5554,N_5387,N_5376);
or U5555 (N_5555,N_5267,N_5388);
or U5556 (N_5556,N_5287,N_5296);
or U5557 (N_5557,N_5250,N_5356);
nand U5558 (N_5558,N_5303,N_5257);
nor U5559 (N_5559,N_5352,N_5201);
and U5560 (N_5560,N_5200,N_5234);
or U5561 (N_5561,N_5326,N_5388);
and U5562 (N_5562,N_5290,N_5265);
or U5563 (N_5563,N_5348,N_5319);
nand U5564 (N_5564,N_5390,N_5329);
nand U5565 (N_5565,N_5395,N_5253);
and U5566 (N_5566,N_5261,N_5349);
nand U5567 (N_5567,N_5315,N_5351);
nand U5568 (N_5568,N_5252,N_5276);
and U5569 (N_5569,N_5283,N_5395);
nand U5570 (N_5570,N_5348,N_5374);
or U5571 (N_5571,N_5378,N_5271);
nand U5572 (N_5572,N_5205,N_5277);
nor U5573 (N_5573,N_5399,N_5300);
or U5574 (N_5574,N_5232,N_5255);
and U5575 (N_5575,N_5200,N_5390);
nand U5576 (N_5576,N_5275,N_5337);
and U5577 (N_5577,N_5300,N_5322);
nor U5578 (N_5578,N_5317,N_5219);
nor U5579 (N_5579,N_5273,N_5378);
and U5580 (N_5580,N_5344,N_5220);
and U5581 (N_5581,N_5331,N_5394);
nor U5582 (N_5582,N_5270,N_5331);
nand U5583 (N_5583,N_5372,N_5394);
or U5584 (N_5584,N_5336,N_5224);
nand U5585 (N_5585,N_5368,N_5269);
nor U5586 (N_5586,N_5310,N_5345);
nor U5587 (N_5587,N_5310,N_5248);
and U5588 (N_5588,N_5224,N_5394);
or U5589 (N_5589,N_5357,N_5323);
nand U5590 (N_5590,N_5266,N_5377);
nand U5591 (N_5591,N_5244,N_5329);
nor U5592 (N_5592,N_5220,N_5232);
nand U5593 (N_5593,N_5353,N_5329);
nand U5594 (N_5594,N_5351,N_5390);
nor U5595 (N_5595,N_5362,N_5351);
nor U5596 (N_5596,N_5261,N_5302);
or U5597 (N_5597,N_5298,N_5283);
nor U5598 (N_5598,N_5353,N_5211);
nor U5599 (N_5599,N_5305,N_5250);
nor U5600 (N_5600,N_5434,N_5562);
xor U5601 (N_5601,N_5402,N_5450);
nor U5602 (N_5602,N_5457,N_5441);
and U5603 (N_5603,N_5533,N_5459);
nor U5604 (N_5604,N_5478,N_5496);
or U5605 (N_5605,N_5498,N_5406);
and U5606 (N_5606,N_5537,N_5461);
nor U5607 (N_5607,N_5506,N_5508);
nand U5608 (N_5608,N_5427,N_5460);
and U5609 (N_5609,N_5404,N_5572);
or U5610 (N_5610,N_5577,N_5580);
or U5611 (N_5611,N_5411,N_5492);
or U5612 (N_5612,N_5437,N_5554);
and U5613 (N_5613,N_5509,N_5505);
nor U5614 (N_5614,N_5445,N_5494);
or U5615 (N_5615,N_5497,N_5431);
nand U5616 (N_5616,N_5594,N_5471);
or U5617 (N_5617,N_5477,N_5422);
and U5618 (N_5618,N_5544,N_5570);
and U5619 (N_5619,N_5532,N_5401);
nand U5620 (N_5620,N_5557,N_5535);
nor U5621 (N_5621,N_5517,N_5529);
nand U5622 (N_5622,N_5487,N_5439);
and U5623 (N_5623,N_5556,N_5489);
nor U5624 (N_5624,N_5482,N_5470);
nor U5625 (N_5625,N_5569,N_5412);
nand U5626 (N_5626,N_5481,N_5530);
nand U5627 (N_5627,N_5418,N_5410);
or U5628 (N_5628,N_5565,N_5486);
or U5629 (N_5629,N_5465,N_5444);
nand U5630 (N_5630,N_5493,N_5455);
nor U5631 (N_5631,N_5547,N_5586);
and U5632 (N_5632,N_5527,N_5588);
nor U5633 (N_5633,N_5559,N_5502);
nor U5634 (N_5634,N_5590,N_5414);
and U5635 (N_5635,N_5551,N_5526);
nor U5636 (N_5636,N_5511,N_5430);
or U5637 (N_5637,N_5574,N_5453);
and U5638 (N_5638,N_5488,N_5483);
nor U5639 (N_5639,N_5548,N_5472);
or U5640 (N_5640,N_5417,N_5582);
xor U5641 (N_5641,N_5428,N_5432);
nand U5642 (N_5642,N_5433,N_5534);
nor U5643 (N_5643,N_5584,N_5480);
and U5644 (N_5644,N_5501,N_5474);
nand U5645 (N_5645,N_5456,N_5499);
xnor U5646 (N_5646,N_5409,N_5598);
and U5647 (N_5647,N_5442,N_5416);
or U5648 (N_5648,N_5519,N_5578);
nand U5649 (N_5649,N_5553,N_5426);
and U5650 (N_5650,N_5421,N_5543);
nand U5651 (N_5651,N_5462,N_5424);
or U5652 (N_5652,N_5449,N_5500);
nor U5653 (N_5653,N_5525,N_5440);
and U5654 (N_5654,N_5429,N_5593);
or U5655 (N_5655,N_5513,N_5420);
or U5656 (N_5656,N_5520,N_5516);
nor U5657 (N_5657,N_5568,N_5435);
and U5658 (N_5658,N_5597,N_5518);
nor U5659 (N_5659,N_5581,N_5552);
and U5660 (N_5660,N_5405,N_5485);
nor U5661 (N_5661,N_5484,N_5592);
nand U5662 (N_5662,N_5558,N_5512);
nand U5663 (N_5663,N_5541,N_5436);
and U5664 (N_5664,N_5515,N_5536);
or U5665 (N_5665,N_5587,N_5571);
and U5666 (N_5666,N_5545,N_5528);
nor U5667 (N_5667,N_5540,N_5555);
and U5668 (N_5668,N_5415,N_5591);
and U5669 (N_5669,N_5561,N_5451);
nor U5670 (N_5670,N_5448,N_5503);
nor U5671 (N_5671,N_5589,N_5550);
and U5672 (N_5672,N_5400,N_5524);
and U5673 (N_5673,N_5566,N_5403);
and U5674 (N_5674,N_5495,N_5531);
nor U5675 (N_5675,N_5564,N_5423);
xor U5676 (N_5676,N_5523,N_5596);
nand U5677 (N_5677,N_5542,N_5538);
nand U5678 (N_5678,N_5463,N_5599);
or U5679 (N_5679,N_5419,N_5579);
nor U5680 (N_5680,N_5514,N_5576);
or U5681 (N_5681,N_5490,N_5546);
and U5682 (N_5682,N_5447,N_5522);
nor U5683 (N_5683,N_5491,N_5521);
nand U5684 (N_5684,N_5408,N_5507);
nand U5685 (N_5685,N_5567,N_5458);
nor U5686 (N_5686,N_5583,N_5464);
nand U5687 (N_5687,N_5595,N_5549);
nand U5688 (N_5688,N_5573,N_5443);
or U5689 (N_5689,N_5475,N_5466);
nor U5690 (N_5690,N_5469,N_5563);
or U5691 (N_5691,N_5575,N_5539);
and U5692 (N_5692,N_5476,N_5413);
nand U5693 (N_5693,N_5504,N_5407);
or U5694 (N_5694,N_5446,N_5438);
nand U5695 (N_5695,N_5452,N_5425);
xnor U5696 (N_5696,N_5468,N_5454);
and U5697 (N_5697,N_5585,N_5560);
and U5698 (N_5698,N_5510,N_5473);
nor U5699 (N_5699,N_5479,N_5467);
and U5700 (N_5700,N_5493,N_5432);
nand U5701 (N_5701,N_5445,N_5432);
nand U5702 (N_5702,N_5515,N_5442);
xor U5703 (N_5703,N_5593,N_5506);
nand U5704 (N_5704,N_5537,N_5422);
and U5705 (N_5705,N_5454,N_5429);
and U5706 (N_5706,N_5567,N_5549);
nand U5707 (N_5707,N_5495,N_5432);
nand U5708 (N_5708,N_5586,N_5418);
nand U5709 (N_5709,N_5420,N_5510);
nand U5710 (N_5710,N_5438,N_5412);
xor U5711 (N_5711,N_5487,N_5508);
nand U5712 (N_5712,N_5499,N_5586);
or U5713 (N_5713,N_5577,N_5555);
nand U5714 (N_5714,N_5468,N_5464);
nand U5715 (N_5715,N_5410,N_5488);
or U5716 (N_5716,N_5586,N_5576);
or U5717 (N_5717,N_5498,N_5462);
nor U5718 (N_5718,N_5502,N_5598);
nand U5719 (N_5719,N_5495,N_5520);
nor U5720 (N_5720,N_5531,N_5474);
or U5721 (N_5721,N_5576,N_5429);
and U5722 (N_5722,N_5568,N_5518);
nor U5723 (N_5723,N_5498,N_5411);
or U5724 (N_5724,N_5426,N_5576);
or U5725 (N_5725,N_5592,N_5506);
nor U5726 (N_5726,N_5535,N_5595);
nand U5727 (N_5727,N_5416,N_5411);
nor U5728 (N_5728,N_5508,N_5558);
and U5729 (N_5729,N_5454,N_5476);
xnor U5730 (N_5730,N_5513,N_5532);
or U5731 (N_5731,N_5545,N_5477);
nand U5732 (N_5732,N_5423,N_5533);
nor U5733 (N_5733,N_5400,N_5568);
and U5734 (N_5734,N_5404,N_5558);
and U5735 (N_5735,N_5597,N_5577);
or U5736 (N_5736,N_5591,N_5426);
and U5737 (N_5737,N_5537,N_5460);
nor U5738 (N_5738,N_5477,N_5473);
nand U5739 (N_5739,N_5456,N_5480);
and U5740 (N_5740,N_5418,N_5584);
nand U5741 (N_5741,N_5455,N_5496);
or U5742 (N_5742,N_5566,N_5518);
nand U5743 (N_5743,N_5488,N_5522);
or U5744 (N_5744,N_5528,N_5521);
or U5745 (N_5745,N_5567,N_5555);
nand U5746 (N_5746,N_5502,N_5549);
and U5747 (N_5747,N_5595,N_5558);
nand U5748 (N_5748,N_5588,N_5590);
nor U5749 (N_5749,N_5480,N_5446);
nand U5750 (N_5750,N_5492,N_5590);
nor U5751 (N_5751,N_5438,N_5561);
xnor U5752 (N_5752,N_5473,N_5558);
and U5753 (N_5753,N_5504,N_5557);
nand U5754 (N_5754,N_5542,N_5427);
nor U5755 (N_5755,N_5552,N_5443);
and U5756 (N_5756,N_5515,N_5590);
nand U5757 (N_5757,N_5425,N_5547);
nand U5758 (N_5758,N_5526,N_5423);
or U5759 (N_5759,N_5576,N_5461);
and U5760 (N_5760,N_5534,N_5561);
nand U5761 (N_5761,N_5584,N_5527);
or U5762 (N_5762,N_5508,N_5476);
or U5763 (N_5763,N_5481,N_5487);
nand U5764 (N_5764,N_5474,N_5449);
nand U5765 (N_5765,N_5451,N_5442);
nor U5766 (N_5766,N_5508,N_5421);
nor U5767 (N_5767,N_5510,N_5476);
or U5768 (N_5768,N_5436,N_5549);
and U5769 (N_5769,N_5437,N_5498);
nor U5770 (N_5770,N_5431,N_5591);
nor U5771 (N_5771,N_5560,N_5497);
or U5772 (N_5772,N_5503,N_5443);
nor U5773 (N_5773,N_5453,N_5498);
or U5774 (N_5774,N_5426,N_5419);
or U5775 (N_5775,N_5501,N_5421);
nand U5776 (N_5776,N_5555,N_5581);
nand U5777 (N_5777,N_5507,N_5442);
or U5778 (N_5778,N_5442,N_5509);
and U5779 (N_5779,N_5492,N_5510);
nand U5780 (N_5780,N_5537,N_5556);
and U5781 (N_5781,N_5598,N_5417);
and U5782 (N_5782,N_5442,N_5510);
nor U5783 (N_5783,N_5579,N_5507);
nand U5784 (N_5784,N_5553,N_5492);
nor U5785 (N_5785,N_5527,N_5518);
or U5786 (N_5786,N_5536,N_5541);
or U5787 (N_5787,N_5570,N_5500);
nor U5788 (N_5788,N_5431,N_5517);
nand U5789 (N_5789,N_5523,N_5487);
or U5790 (N_5790,N_5459,N_5488);
nor U5791 (N_5791,N_5544,N_5474);
and U5792 (N_5792,N_5454,N_5530);
and U5793 (N_5793,N_5499,N_5552);
or U5794 (N_5794,N_5531,N_5509);
xor U5795 (N_5795,N_5432,N_5588);
and U5796 (N_5796,N_5465,N_5558);
xor U5797 (N_5797,N_5401,N_5544);
and U5798 (N_5798,N_5447,N_5556);
xor U5799 (N_5799,N_5577,N_5422);
and U5800 (N_5800,N_5651,N_5797);
nand U5801 (N_5801,N_5771,N_5727);
or U5802 (N_5802,N_5704,N_5745);
or U5803 (N_5803,N_5729,N_5608);
or U5804 (N_5804,N_5732,N_5623);
and U5805 (N_5805,N_5718,N_5739);
nand U5806 (N_5806,N_5757,N_5627);
nand U5807 (N_5807,N_5721,N_5619);
nand U5808 (N_5808,N_5687,N_5786);
and U5809 (N_5809,N_5688,N_5773);
nand U5810 (N_5810,N_5620,N_5672);
nand U5811 (N_5811,N_5724,N_5740);
and U5812 (N_5812,N_5643,N_5795);
nor U5813 (N_5813,N_5639,N_5614);
or U5814 (N_5814,N_5618,N_5629);
nand U5815 (N_5815,N_5642,N_5701);
nand U5816 (N_5816,N_5603,N_5666);
nor U5817 (N_5817,N_5778,N_5783);
and U5818 (N_5818,N_5705,N_5692);
nor U5819 (N_5819,N_5612,N_5690);
nor U5820 (N_5820,N_5607,N_5706);
and U5821 (N_5821,N_5696,N_5787);
or U5822 (N_5822,N_5695,N_5645);
nand U5823 (N_5823,N_5653,N_5624);
nand U5824 (N_5824,N_5714,N_5726);
xnor U5825 (N_5825,N_5677,N_5793);
nor U5826 (N_5826,N_5678,N_5691);
or U5827 (N_5827,N_5638,N_5667);
or U5828 (N_5828,N_5790,N_5765);
nand U5829 (N_5829,N_5713,N_5799);
nand U5830 (N_5830,N_5613,N_5788);
or U5831 (N_5831,N_5676,N_5637);
nor U5832 (N_5832,N_5606,N_5716);
nand U5833 (N_5833,N_5710,N_5725);
nand U5834 (N_5834,N_5641,N_5751);
or U5835 (N_5835,N_5632,N_5763);
and U5836 (N_5836,N_5720,N_5657);
and U5837 (N_5837,N_5625,N_5700);
or U5838 (N_5838,N_5604,N_5774);
or U5839 (N_5839,N_5630,N_5600);
nor U5840 (N_5840,N_5683,N_5709);
or U5841 (N_5841,N_5753,N_5654);
nor U5842 (N_5842,N_5626,N_5752);
and U5843 (N_5843,N_5611,N_5768);
or U5844 (N_5844,N_5609,N_5723);
and U5845 (N_5845,N_5764,N_5648);
and U5846 (N_5846,N_5650,N_5798);
and U5847 (N_5847,N_5715,N_5659);
nand U5848 (N_5848,N_5747,N_5675);
or U5849 (N_5849,N_5628,N_5662);
nand U5850 (N_5850,N_5766,N_5722);
nor U5851 (N_5851,N_5686,N_5674);
or U5852 (N_5852,N_5734,N_5728);
nand U5853 (N_5853,N_5646,N_5762);
nor U5854 (N_5854,N_5731,N_5635);
nand U5855 (N_5855,N_5661,N_5616);
nor U5856 (N_5856,N_5761,N_5789);
nand U5857 (N_5857,N_5689,N_5668);
nor U5858 (N_5858,N_5703,N_5796);
and U5859 (N_5859,N_5784,N_5711);
or U5860 (N_5860,N_5776,N_5622);
and U5861 (N_5861,N_5679,N_5792);
nand U5862 (N_5862,N_5794,N_5756);
nor U5863 (N_5863,N_5707,N_5760);
and U5864 (N_5864,N_5719,N_5656);
or U5865 (N_5865,N_5750,N_5702);
xor U5866 (N_5866,N_5782,N_5655);
nor U5867 (N_5867,N_5775,N_5758);
nand U5868 (N_5868,N_5779,N_5693);
and U5869 (N_5869,N_5615,N_5736);
or U5870 (N_5870,N_5746,N_5785);
nor U5871 (N_5871,N_5755,N_5769);
and U5872 (N_5872,N_5669,N_5617);
and U5873 (N_5873,N_5749,N_5717);
or U5874 (N_5874,N_5733,N_5735);
and U5875 (N_5875,N_5647,N_5777);
nand U5876 (N_5876,N_5781,N_5759);
nand U5877 (N_5877,N_5649,N_5770);
nor U5878 (N_5878,N_5633,N_5682);
or U5879 (N_5879,N_5671,N_5791);
or U5880 (N_5880,N_5634,N_5708);
nand U5881 (N_5881,N_5712,N_5670);
nand U5882 (N_5882,N_5602,N_5605);
nand U5883 (N_5883,N_5737,N_5673);
nor U5884 (N_5884,N_5664,N_5772);
and U5885 (N_5885,N_5684,N_5681);
nor U5886 (N_5886,N_5699,N_5694);
nand U5887 (N_5887,N_5658,N_5663);
nor U5888 (N_5888,N_5636,N_5743);
or U5889 (N_5889,N_5660,N_5621);
or U5890 (N_5890,N_5644,N_5744);
xor U5891 (N_5891,N_5748,N_5631);
or U5892 (N_5892,N_5780,N_5767);
nand U5893 (N_5893,N_5754,N_5738);
or U5894 (N_5894,N_5652,N_5741);
and U5895 (N_5895,N_5730,N_5680);
and U5896 (N_5896,N_5697,N_5640);
nand U5897 (N_5897,N_5665,N_5685);
nor U5898 (N_5898,N_5698,N_5601);
and U5899 (N_5899,N_5610,N_5742);
xnor U5900 (N_5900,N_5774,N_5702);
nor U5901 (N_5901,N_5628,N_5767);
nand U5902 (N_5902,N_5775,N_5751);
nand U5903 (N_5903,N_5732,N_5736);
or U5904 (N_5904,N_5702,N_5622);
or U5905 (N_5905,N_5697,N_5686);
nor U5906 (N_5906,N_5760,N_5789);
nor U5907 (N_5907,N_5786,N_5739);
or U5908 (N_5908,N_5686,N_5662);
or U5909 (N_5909,N_5794,N_5641);
nand U5910 (N_5910,N_5623,N_5729);
nor U5911 (N_5911,N_5702,N_5749);
and U5912 (N_5912,N_5690,N_5678);
nand U5913 (N_5913,N_5702,N_5740);
and U5914 (N_5914,N_5795,N_5799);
and U5915 (N_5915,N_5780,N_5698);
nor U5916 (N_5916,N_5709,N_5670);
nor U5917 (N_5917,N_5714,N_5799);
or U5918 (N_5918,N_5679,N_5644);
or U5919 (N_5919,N_5627,N_5702);
or U5920 (N_5920,N_5644,N_5720);
or U5921 (N_5921,N_5722,N_5623);
nor U5922 (N_5922,N_5653,N_5753);
or U5923 (N_5923,N_5646,N_5785);
xnor U5924 (N_5924,N_5691,N_5706);
and U5925 (N_5925,N_5607,N_5670);
nor U5926 (N_5926,N_5640,N_5613);
nand U5927 (N_5927,N_5780,N_5710);
nor U5928 (N_5928,N_5615,N_5794);
nor U5929 (N_5929,N_5617,N_5736);
nand U5930 (N_5930,N_5688,N_5603);
and U5931 (N_5931,N_5774,N_5645);
nand U5932 (N_5932,N_5682,N_5623);
or U5933 (N_5933,N_5668,N_5776);
nand U5934 (N_5934,N_5624,N_5782);
and U5935 (N_5935,N_5606,N_5604);
nand U5936 (N_5936,N_5717,N_5657);
or U5937 (N_5937,N_5793,N_5623);
or U5938 (N_5938,N_5640,N_5653);
nand U5939 (N_5939,N_5684,N_5763);
or U5940 (N_5940,N_5621,N_5762);
nor U5941 (N_5941,N_5607,N_5712);
and U5942 (N_5942,N_5702,N_5635);
and U5943 (N_5943,N_5641,N_5625);
and U5944 (N_5944,N_5646,N_5775);
nand U5945 (N_5945,N_5758,N_5661);
nor U5946 (N_5946,N_5632,N_5787);
nand U5947 (N_5947,N_5710,N_5663);
and U5948 (N_5948,N_5671,N_5630);
or U5949 (N_5949,N_5756,N_5646);
and U5950 (N_5950,N_5737,N_5785);
or U5951 (N_5951,N_5750,N_5690);
xor U5952 (N_5952,N_5623,N_5765);
or U5953 (N_5953,N_5754,N_5798);
and U5954 (N_5954,N_5740,N_5686);
nand U5955 (N_5955,N_5648,N_5744);
nand U5956 (N_5956,N_5627,N_5720);
nand U5957 (N_5957,N_5677,N_5675);
nand U5958 (N_5958,N_5730,N_5679);
nor U5959 (N_5959,N_5648,N_5788);
nand U5960 (N_5960,N_5631,N_5600);
or U5961 (N_5961,N_5633,N_5746);
or U5962 (N_5962,N_5611,N_5782);
or U5963 (N_5963,N_5660,N_5696);
nand U5964 (N_5964,N_5636,N_5632);
nor U5965 (N_5965,N_5755,N_5638);
and U5966 (N_5966,N_5771,N_5673);
nor U5967 (N_5967,N_5631,N_5678);
or U5968 (N_5968,N_5672,N_5628);
or U5969 (N_5969,N_5746,N_5695);
xnor U5970 (N_5970,N_5679,N_5776);
nor U5971 (N_5971,N_5632,N_5794);
or U5972 (N_5972,N_5711,N_5704);
nand U5973 (N_5973,N_5602,N_5706);
nor U5974 (N_5974,N_5730,N_5601);
or U5975 (N_5975,N_5669,N_5641);
or U5976 (N_5976,N_5609,N_5700);
or U5977 (N_5977,N_5610,N_5680);
and U5978 (N_5978,N_5600,N_5763);
nor U5979 (N_5979,N_5624,N_5791);
and U5980 (N_5980,N_5786,N_5757);
and U5981 (N_5981,N_5649,N_5714);
and U5982 (N_5982,N_5764,N_5611);
and U5983 (N_5983,N_5754,N_5618);
nand U5984 (N_5984,N_5734,N_5746);
nand U5985 (N_5985,N_5713,N_5781);
nor U5986 (N_5986,N_5656,N_5610);
or U5987 (N_5987,N_5761,N_5631);
and U5988 (N_5988,N_5764,N_5760);
and U5989 (N_5989,N_5685,N_5601);
or U5990 (N_5990,N_5725,N_5705);
or U5991 (N_5991,N_5606,N_5659);
nand U5992 (N_5992,N_5770,N_5604);
and U5993 (N_5993,N_5696,N_5690);
and U5994 (N_5994,N_5669,N_5760);
or U5995 (N_5995,N_5675,N_5654);
or U5996 (N_5996,N_5624,N_5661);
nor U5997 (N_5997,N_5760,N_5606);
nand U5998 (N_5998,N_5627,N_5617);
nand U5999 (N_5999,N_5792,N_5731);
and U6000 (N_6000,N_5824,N_5926);
xor U6001 (N_6001,N_5852,N_5984);
and U6002 (N_6002,N_5973,N_5801);
and U6003 (N_6003,N_5880,N_5952);
or U6004 (N_6004,N_5871,N_5983);
xnor U6005 (N_6005,N_5883,N_5985);
nor U6006 (N_6006,N_5941,N_5830);
and U6007 (N_6007,N_5825,N_5853);
nand U6008 (N_6008,N_5818,N_5951);
nand U6009 (N_6009,N_5861,N_5970);
and U6010 (N_6010,N_5874,N_5826);
and U6011 (N_6011,N_5897,N_5997);
or U6012 (N_6012,N_5901,N_5966);
and U6013 (N_6013,N_5860,N_5930);
nand U6014 (N_6014,N_5991,N_5844);
and U6015 (N_6015,N_5831,N_5885);
nand U6016 (N_6016,N_5828,N_5854);
nand U6017 (N_6017,N_5900,N_5992);
or U6018 (N_6018,N_5922,N_5894);
xor U6019 (N_6019,N_5902,N_5817);
or U6020 (N_6020,N_5963,N_5808);
and U6021 (N_6021,N_5990,N_5890);
and U6022 (N_6022,N_5912,N_5892);
or U6023 (N_6023,N_5804,N_5971);
and U6024 (N_6024,N_5908,N_5998);
or U6025 (N_6025,N_5988,N_5867);
and U6026 (N_6026,N_5955,N_5904);
and U6027 (N_6027,N_5907,N_5843);
xnor U6028 (N_6028,N_5995,N_5823);
nor U6029 (N_6029,N_5954,N_5836);
or U6030 (N_6030,N_5862,N_5924);
nand U6031 (N_6031,N_5928,N_5875);
nand U6032 (N_6032,N_5811,N_5979);
or U6033 (N_6033,N_5977,N_5911);
nor U6034 (N_6034,N_5842,N_5986);
and U6035 (N_6035,N_5835,N_5933);
and U6036 (N_6036,N_5877,N_5993);
and U6037 (N_6037,N_5943,N_5850);
nor U6038 (N_6038,N_5962,N_5972);
and U6039 (N_6039,N_5821,N_5974);
nor U6040 (N_6040,N_5975,N_5814);
nor U6041 (N_6041,N_5919,N_5816);
nor U6042 (N_6042,N_5887,N_5849);
nand U6043 (N_6043,N_5947,N_5969);
and U6044 (N_6044,N_5964,N_5809);
xnor U6045 (N_6045,N_5967,N_5932);
and U6046 (N_6046,N_5976,N_5873);
nor U6047 (N_6047,N_5810,N_5927);
or U6048 (N_6048,N_5863,N_5936);
nor U6049 (N_6049,N_5884,N_5965);
and U6050 (N_6050,N_5978,N_5961);
or U6051 (N_6051,N_5929,N_5870);
or U6052 (N_6052,N_5888,N_5827);
xor U6053 (N_6053,N_5953,N_5858);
and U6054 (N_6054,N_5838,N_5812);
and U6055 (N_6055,N_5906,N_5848);
or U6056 (N_6056,N_5847,N_5800);
or U6057 (N_6057,N_5819,N_5968);
nor U6058 (N_6058,N_5921,N_5889);
nand U6059 (N_6059,N_5851,N_5945);
and U6060 (N_6060,N_5996,N_5931);
and U6061 (N_6061,N_5949,N_5935);
nor U6062 (N_6062,N_5958,N_5815);
and U6063 (N_6063,N_5917,N_5939);
nor U6064 (N_6064,N_5868,N_5959);
or U6065 (N_6065,N_5925,N_5946);
xnor U6066 (N_6066,N_5845,N_5857);
nor U6067 (N_6067,N_5864,N_5896);
nand U6068 (N_6068,N_5994,N_5938);
xnor U6069 (N_6069,N_5855,N_5980);
nand U6070 (N_6070,N_5840,N_5829);
and U6071 (N_6071,N_5920,N_5822);
nand U6072 (N_6072,N_5899,N_5803);
nand U6073 (N_6073,N_5999,N_5895);
and U6074 (N_6074,N_5957,N_5893);
and U6075 (N_6075,N_5918,N_5807);
or U6076 (N_6076,N_5859,N_5805);
nand U6077 (N_6077,N_5839,N_5872);
or U6078 (N_6078,N_5806,N_5802);
and U6079 (N_6079,N_5865,N_5937);
and U6080 (N_6080,N_5915,N_5948);
nand U6081 (N_6081,N_5833,N_5903);
and U6082 (N_6082,N_5891,N_5956);
nand U6083 (N_6083,N_5886,N_5942);
nand U6084 (N_6084,N_5909,N_5882);
or U6085 (N_6085,N_5813,N_5987);
nor U6086 (N_6086,N_5846,N_5989);
nand U6087 (N_6087,N_5856,N_5910);
or U6088 (N_6088,N_5878,N_5898);
nor U6089 (N_6089,N_5866,N_5940);
and U6090 (N_6090,N_5834,N_5981);
nor U6091 (N_6091,N_5820,N_5869);
nand U6092 (N_6092,N_5876,N_5841);
nand U6093 (N_6093,N_5950,N_5923);
nor U6094 (N_6094,N_5914,N_5982);
nor U6095 (N_6095,N_5879,N_5944);
or U6096 (N_6096,N_5934,N_5960);
nor U6097 (N_6097,N_5913,N_5837);
nand U6098 (N_6098,N_5832,N_5881);
nand U6099 (N_6099,N_5916,N_5905);
nor U6100 (N_6100,N_5930,N_5879);
and U6101 (N_6101,N_5962,N_5944);
and U6102 (N_6102,N_5827,N_5837);
or U6103 (N_6103,N_5992,N_5881);
xnor U6104 (N_6104,N_5912,N_5915);
nor U6105 (N_6105,N_5826,N_5877);
nand U6106 (N_6106,N_5910,N_5978);
nand U6107 (N_6107,N_5963,N_5802);
xnor U6108 (N_6108,N_5893,N_5865);
nand U6109 (N_6109,N_5823,N_5935);
xor U6110 (N_6110,N_5881,N_5844);
nand U6111 (N_6111,N_5892,N_5939);
nor U6112 (N_6112,N_5838,N_5952);
and U6113 (N_6113,N_5939,N_5849);
nor U6114 (N_6114,N_5945,N_5887);
nor U6115 (N_6115,N_5840,N_5965);
nor U6116 (N_6116,N_5948,N_5880);
nand U6117 (N_6117,N_5949,N_5839);
nand U6118 (N_6118,N_5929,N_5931);
or U6119 (N_6119,N_5898,N_5900);
and U6120 (N_6120,N_5902,N_5945);
and U6121 (N_6121,N_5910,N_5886);
nand U6122 (N_6122,N_5814,N_5858);
nand U6123 (N_6123,N_5997,N_5999);
xnor U6124 (N_6124,N_5815,N_5865);
nor U6125 (N_6125,N_5923,N_5822);
and U6126 (N_6126,N_5952,N_5892);
nor U6127 (N_6127,N_5802,N_5951);
nor U6128 (N_6128,N_5946,N_5847);
and U6129 (N_6129,N_5894,N_5992);
nand U6130 (N_6130,N_5876,N_5931);
nor U6131 (N_6131,N_5811,N_5948);
nand U6132 (N_6132,N_5960,N_5880);
nor U6133 (N_6133,N_5976,N_5912);
nand U6134 (N_6134,N_5998,N_5870);
nor U6135 (N_6135,N_5904,N_5802);
or U6136 (N_6136,N_5889,N_5969);
nand U6137 (N_6137,N_5817,N_5901);
or U6138 (N_6138,N_5826,N_5821);
or U6139 (N_6139,N_5965,N_5928);
nor U6140 (N_6140,N_5875,N_5900);
xnor U6141 (N_6141,N_5824,N_5806);
or U6142 (N_6142,N_5815,N_5936);
nand U6143 (N_6143,N_5890,N_5975);
and U6144 (N_6144,N_5990,N_5876);
or U6145 (N_6145,N_5961,N_5985);
or U6146 (N_6146,N_5972,N_5901);
nand U6147 (N_6147,N_5883,N_5911);
or U6148 (N_6148,N_5835,N_5858);
and U6149 (N_6149,N_5989,N_5901);
or U6150 (N_6150,N_5966,N_5938);
nor U6151 (N_6151,N_5945,N_5933);
nor U6152 (N_6152,N_5812,N_5860);
nand U6153 (N_6153,N_5853,N_5893);
nor U6154 (N_6154,N_5938,N_5993);
nor U6155 (N_6155,N_5971,N_5907);
nand U6156 (N_6156,N_5883,N_5877);
or U6157 (N_6157,N_5872,N_5807);
xor U6158 (N_6158,N_5848,N_5926);
and U6159 (N_6159,N_5872,N_5968);
and U6160 (N_6160,N_5924,N_5900);
or U6161 (N_6161,N_5927,N_5862);
nand U6162 (N_6162,N_5943,N_5919);
nor U6163 (N_6163,N_5840,N_5933);
nor U6164 (N_6164,N_5889,N_5905);
or U6165 (N_6165,N_5899,N_5807);
nor U6166 (N_6166,N_5932,N_5886);
nand U6167 (N_6167,N_5839,N_5901);
nand U6168 (N_6168,N_5899,N_5877);
or U6169 (N_6169,N_5910,N_5950);
xor U6170 (N_6170,N_5985,N_5861);
or U6171 (N_6171,N_5958,N_5972);
nor U6172 (N_6172,N_5880,N_5935);
and U6173 (N_6173,N_5845,N_5928);
nand U6174 (N_6174,N_5866,N_5978);
and U6175 (N_6175,N_5856,N_5878);
nand U6176 (N_6176,N_5986,N_5824);
or U6177 (N_6177,N_5849,N_5922);
nand U6178 (N_6178,N_5863,N_5827);
or U6179 (N_6179,N_5881,N_5939);
nand U6180 (N_6180,N_5811,N_5927);
nor U6181 (N_6181,N_5871,N_5874);
and U6182 (N_6182,N_5929,N_5952);
nor U6183 (N_6183,N_5898,N_5824);
and U6184 (N_6184,N_5833,N_5953);
nand U6185 (N_6185,N_5990,N_5837);
and U6186 (N_6186,N_5920,N_5827);
and U6187 (N_6187,N_5855,N_5875);
nand U6188 (N_6188,N_5967,N_5810);
or U6189 (N_6189,N_5968,N_5849);
nand U6190 (N_6190,N_5908,N_5854);
or U6191 (N_6191,N_5872,N_5857);
and U6192 (N_6192,N_5870,N_5880);
and U6193 (N_6193,N_5875,N_5957);
or U6194 (N_6194,N_5989,N_5999);
and U6195 (N_6195,N_5920,N_5842);
nand U6196 (N_6196,N_5885,N_5980);
nand U6197 (N_6197,N_5877,N_5876);
and U6198 (N_6198,N_5881,N_5807);
and U6199 (N_6199,N_5969,N_5856);
or U6200 (N_6200,N_6155,N_6082);
and U6201 (N_6201,N_6129,N_6025);
or U6202 (N_6202,N_6144,N_6104);
nand U6203 (N_6203,N_6036,N_6127);
and U6204 (N_6204,N_6106,N_6077);
nor U6205 (N_6205,N_6103,N_6074);
nand U6206 (N_6206,N_6071,N_6114);
nor U6207 (N_6207,N_6001,N_6136);
nand U6208 (N_6208,N_6131,N_6035);
xor U6209 (N_6209,N_6117,N_6064);
and U6210 (N_6210,N_6184,N_6094);
or U6211 (N_6211,N_6086,N_6034);
nor U6212 (N_6212,N_6125,N_6084);
and U6213 (N_6213,N_6047,N_6151);
nor U6214 (N_6214,N_6021,N_6121);
nor U6215 (N_6215,N_6067,N_6028);
nor U6216 (N_6216,N_6142,N_6169);
nand U6217 (N_6217,N_6081,N_6051);
nand U6218 (N_6218,N_6132,N_6032);
or U6219 (N_6219,N_6110,N_6033);
or U6220 (N_6220,N_6165,N_6143);
and U6221 (N_6221,N_6062,N_6005);
nand U6222 (N_6222,N_6056,N_6115);
nor U6223 (N_6223,N_6006,N_6146);
nand U6224 (N_6224,N_6113,N_6135);
nor U6225 (N_6225,N_6167,N_6041);
nand U6226 (N_6226,N_6099,N_6186);
and U6227 (N_6227,N_6193,N_6163);
and U6228 (N_6228,N_6160,N_6179);
nor U6229 (N_6229,N_6116,N_6171);
or U6230 (N_6230,N_6089,N_6178);
xor U6231 (N_6231,N_6076,N_6019);
nand U6232 (N_6232,N_6180,N_6137);
nand U6233 (N_6233,N_6069,N_6105);
or U6234 (N_6234,N_6055,N_6042);
or U6235 (N_6235,N_6139,N_6145);
nor U6236 (N_6236,N_6085,N_6096);
and U6237 (N_6237,N_6174,N_6101);
or U6238 (N_6238,N_6014,N_6173);
and U6239 (N_6239,N_6149,N_6053);
and U6240 (N_6240,N_6192,N_6083);
and U6241 (N_6241,N_6195,N_6112);
nor U6242 (N_6242,N_6016,N_6119);
and U6243 (N_6243,N_6128,N_6168);
and U6244 (N_6244,N_6141,N_6108);
nand U6245 (N_6245,N_6150,N_6038);
nand U6246 (N_6246,N_6176,N_6107);
or U6247 (N_6247,N_6090,N_6052);
and U6248 (N_6248,N_6102,N_6199);
and U6249 (N_6249,N_6166,N_6185);
and U6250 (N_6250,N_6189,N_6073);
or U6251 (N_6251,N_6175,N_6066);
or U6252 (N_6252,N_6087,N_6134);
nand U6253 (N_6253,N_6037,N_6177);
nor U6254 (N_6254,N_6068,N_6063);
nand U6255 (N_6255,N_6161,N_6126);
nor U6256 (N_6256,N_6003,N_6010);
or U6257 (N_6257,N_6024,N_6098);
or U6258 (N_6258,N_6188,N_6162);
or U6259 (N_6259,N_6029,N_6097);
nor U6260 (N_6260,N_6198,N_6122);
nand U6261 (N_6261,N_6123,N_6039);
nand U6262 (N_6262,N_6133,N_6046);
xor U6263 (N_6263,N_6059,N_6040);
nand U6264 (N_6264,N_6170,N_6026);
and U6265 (N_6265,N_6013,N_6031);
nand U6266 (N_6266,N_6138,N_6111);
nor U6267 (N_6267,N_6091,N_6015);
and U6268 (N_6268,N_6043,N_6183);
or U6269 (N_6269,N_6030,N_6045);
or U6270 (N_6270,N_6152,N_6118);
nand U6271 (N_6271,N_6095,N_6158);
or U6272 (N_6272,N_6148,N_6092);
and U6273 (N_6273,N_6080,N_6008);
or U6274 (N_6274,N_6002,N_6022);
nor U6275 (N_6275,N_6050,N_6156);
nand U6276 (N_6276,N_6075,N_6157);
or U6277 (N_6277,N_6182,N_6048);
or U6278 (N_6278,N_6078,N_6061);
nor U6279 (N_6279,N_6196,N_6018);
or U6280 (N_6280,N_6191,N_6023);
or U6281 (N_6281,N_6058,N_6190);
xor U6282 (N_6282,N_6004,N_6079);
or U6283 (N_6283,N_6027,N_6124);
or U6284 (N_6284,N_6044,N_6088);
or U6285 (N_6285,N_6130,N_6187);
nand U6286 (N_6286,N_6065,N_6140);
nor U6287 (N_6287,N_6197,N_6060);
and U6288 (N_6288,N_6017,N_6057);
and U6289 (N_6289,N_6009,N_6072);
nor U6290 (N_6290,N_6172,N_6054);
nor U6291 (N_6291,N_6120,N_6070);
and U6292 (N_6292,N_6164,N_6093);
nand U6293 (N_6293,N_6194,N_6159);
and U6294 (N_6294,N_6020,N_6154);
nand U6295 (N_6295,N_6049,N_6011);
or U6296 (N_6296,N_6109,N_6007);
or U6297 (N_6297,N_6153,N_6012);
nor U6298 (N_6298,N_6100,N_6147);
or U6299 (N_6299,N_6000,N_6181);
nand U6300 (N_6300,N_6006,N_6048);
nor U6301 (N_6301,N_6082,N_6061);
or U6302 (N_6302,N_6068,N_6177);
and U6303 (N_6303,N_6108,N_6048);
or U6304 (N_6304,N_6140,N_6190);
nor U6305 (N_6305,N_6008,N_6196);
and U6306 (N_6306,N_6002,N_6115);
nor U6307 (N_6307,N_6010,N_6034);
nand U6308 (N_6308,N_6153,N_6104);
or U6309 (N_6309,N_6138,N_6105);
nand U6310 (N_6310,N_6136,N_6119);
nand U6311 (N_6311,N_6058,N_6180);
or U6312 (N_6312,N_6065,N_6011);
nand U6313 (N_6313,N_6198,N_6047);
or U6314 (N_6314,N_6188,N_6199);
nand U6315 (N_6315,N_6055,N_6177);
and U6316 (N_6316,N_6124,N_6038);
nor U6317 (N_6317,N_6101,N_6080);
or U6318 (N_6318,N_6168,N_6061);
or U6319 (N_6319,N_6116,N_6160);
or U6320 (N_6320,N_6132,N_6104);
and U6321 (N_6321,N_6178,N_6193);
nor U6322 (N_6322,N_6141,N_6087);
nor U6323 (N_6323,N_6050,N_6037);
nor U6324 (N_6324,N_6099,N_6022);
xnor U6325 (N_6325,N_6185,N_6036);
nor U6326 (N_6326,N_6118,N_6113);
nor U6327 (N_6327,N_6007,N_6162);
nand U6328 (N_6328,N_6106,N_6014);
and U6329 (N_6329,N_6123,N_6025);
and U6330 (N_6330,N_6105,N_6111);
xnor U6331 (N_6331,N_6141,N_6145);
nand U6332 (N_6332,N_6082,N_6004);
nor U6333 (N_6333,N_6124,N_6025);
and U6334 (N_6334,N_6138,N_6156);
and U6335 (N_6335,N_6171,N_6062);
or U6336 (N_6336,N_6164,N_6074);
or U6337 (N_6337,N_6105,N_6042);
xor U6338 (N_6338,N_6159,N_6103);
and U6339 (N_6339,N_6026,N_6073);
or U6340 (N_6340,N_6116,N_6128);
nand U6341 (N_6341,N_6014,N_6128);
and U6342 (N_6342,N_6005,N_6163);
and U6343 (N_6343,N_6059,N_6171);
nand U6344 (N_6344,N_6125,N_6171);
nand U6345 (N_6345,N_6059,N_6005);
nand U6346 (N_6346,N_6011,N_6043);
or U6347 (N_6347,N_6119,N_6128);
nor U6348 (N_6348,N_6080,N_6123);
or U6349 (N_6349,N_6013,N_6063);
and U6350 (N_6350,N_6112,N_6168);
nand U6351 (N_6351,N_6005,N_6101);
nor U6352 (N_6352,N_6165,N_6044);
nand U6353 (N_6353,N_6013,N_6011);
or U6354 (N_6354,N_6074,N_6145);
or U6355 (N_6355,N_6071,N_6035);
nand U6356 (N_6356,N_6179,N_6014);
or U6357 (N_6357,N_6063,N_6076);
xnor U6358 (N_6358,N_6137,N_6093);
and U6359 (N_6359,N_6085,N_6190);
nor U6360 (N_6360,N_6133,N_6142);
nor U6361 (N_6361,N_6142,N_6168);
or U6362 (N_6362,N_6078,N_6023);
nor U6363 (N_6363,N_6100,N_6123);
nor U6364 (N_6364,N_6192,N_6134);
and U6365 (N_6365,N_6029,N_6099);
or U6366 (N_6366,N_6089,N_6191);
nand U6367 (N_6367,N_6199,N_6135);
and U6368 (N_6368,N_6187,N_6188);
nor U6369 (N_6369,N_6103,N_6127);
nor U6370 (N_6370,N_6175,N_6159);
and U6371 (N_6371,N_6154,N_6011);
or U6372 (N_6372,N_6173,N_6087);
and U6373 (N_6373,N_6166,N_6061);
and U6374 (N_6374,N_6035,N_6106);
nand U6375 (N_6375,N_6163,N_6125);
and U6376 (N_6376,N_6180,N_6116);
and U6377 (N_6377,N_6010,N_6048);
or U6378 (N_6378,N_6051,N_6078);
or U6379 (N_6379,N_6178,N_6099);
and U6380 (N_6380,N_6091,N_6023);
nor U6381 (N_6381,N_6037,N_6020);
nor U6382 (N_6382,N_6151,N_6022);
nor U6383 (N_6383,N_6163,N_6176);
and U6384 (N_6384,N_6079,N_6083);
or U6385 (N_6385,N_6120,N_6006);
and U6386 (N_6386,N_6043,N_6056);
or U6387 (N_6387,N_6024,N_6092);
nand U6388 (N_6388,N_6192,N_6168);
or U6389 (N_6389,N_6119,N_6184);
and U6390 (N_6390,N_6048,N_6169);
nor U6391 (N_6391,N_6176,N_6191);
nor U6392 (N_6392,N_6156,N_6108);
nand U6393 (N_6393,N_6130,N_6027);
nor U6394 (N_6394,N_6165,N_6198);
nor U6395 (N_6395,N_6017,N_6011);
or U6396 (N_6396,N_6038,N_6170);
or U6397 (N_6397,N_6072,N_6074);
xnor U6398 (N_6398,N_6067,N_6008);
nand U6399 (N_6399,N_6187,N_6145);
nand U6400 (N_6400,N_6246,N_6389);
and U6401 (N_6401,N_6250,N_6374);
and U6402 (N_6402,N_6339,N_6312);
nand U6403 (N_6403,N_6278,N_6275);
or U6404 (N_6404,N_6328,N_6218);
and U6405 (N_6405,N_6318,N_6253);
or U6406 (N_6406,N_6321,N_6364);
nand U6407 (N_6407,N_6210,N_6229);
nor U6408 (N_6408,N_6303,N_6256);
nand U6409 (N_6409,N_6348,N_6216);
and U6410 (N_6410,N_6317,N_6342);
nor U6411 (N_6411,N_6384,N_6376);
and U6412 (N_6412,N_6265,N_6322);
or U6413 (N_6413,N_6395,N_6379);
nor U6414 (N_6414,N_6300,N_6259);
and U6415 (N_6415,N_6217,N_6262);
or U6416 (N_6416,N_6288,N_6373);
nand U6417 (N_6417,N_6356,N_6249);
and U6418 (N_6418,N_6357,N_6286);
nor U6419 (N_6419,N_6241,N_6363);
or U6420 (N_6420,N_6289,N_6203);
nand U6421 (N_6421,N_6238,N_6396);
nand U6422 (N_6422,N_6244,N_6240);
xor U6423 (N_6423,N_6274,N_6263);
and U6424 (N_6424,N_6325,N_6232);
nor U6425 (N_6425,N_6360,N_6242);
nand U6426 (N_6426,N_6378,N_6316);
nand U6427 (N_6427,N_6280,N_6207);
nand U6428 (N_6428,N_6239,N_6248);
and U6429 (N_6429,N_6366,N_6313);
xor U6430 (N_6430,N_6370,N_6347);
nor U6431 (N_6431,N_6371,N_6385);
or U6432 (N_6432,N_6237,N_6230);
nor U6433 (N_6433,N_6369,N_6223);
nand U6434 (N_6434,N_6330,N_6358);
xor U6435 (N_6435,N_6226,N_6293);
nor U6436 (N_6436,N_6394,N_6386);
nor U6437 (N_6437,N_6340,N_6380);
and U6438 (N_6438,N_6255,N_6251);
or U6439 (N_6439,N_6397,N_6335);
and U6440 (N_6440,N_6326,N_6332);
or U6441 (N_6441,N_6224,N_6287);
nand U6442 (N_6442,N_6338,N_6277);
and U6443 (N_6443,N_6261,N_6390);
and U6444 (N_6444,N_6297,N_6291);
nor U6445 (N_6445,N_6204,N_6212);
or U6446 (N_6446,N_6213,N_6269);
nand U6447 (N_6447,N_6301,N_6276);
nor U6448 (N_6448,N_6341,N_6387);
and U6449 (N_6449,N_6235,N_6344);
nand U6450 (N_6450,N_6228,N_6329);
and U6451 (N_6451,N_6309,N_6343);
or U6452 (N_6452,N_6383,N_6225);
or U6453 (N_6453,N_6222,N_6302);
and U6454 (N_6454,N_6333,N_6202);
nor U6455 (N_6455,N_6252,N_6391);
nand U6456 (N_6456,N_6268,N_6382);
nor U6457 (N_6457,N_6258,N_6361);
or U6458 (N_6458,N_6272,N_6367);
or U6459 (N_6459,N_6319,N_6398);
nor U6460 (N_6460,N_6392,N_6290);
and U6461 (N_6461,N_6306,N_6345);
and U6462 (N_6462,N_6219,N_6220);
nand U6463 (N_6463,N_6282,N_6372);
nor U6464 (N_6464,N_6295,N_6311);
nor U6465 (N_6465,N_6368,N_6284);
and U6466 (N_6466,N_6211,N_6381);
and U6467 (N_6467,N_6334,N_6336);
and U6468 (N_6468,N_6200,N_6346);
and U6469 (N_6469,N_6308,N_6375);
nand U6470 (N_6470,N_6267,N_6349);
nor U6471 (N_6471,N_6377,N_6215);
xor U6472 (N_6472,N_6351,N_6320);
and U6473 (N_6473,N_6365,N_6236);
nand U6474 (N_6474,N_6307,N_6314);
or U6475 (N_6475,N_6299,N_6247);
nand U6476 (N_6476,N_6266,N_6355);
nor U6477 (N_6477,N_6201,N_6254);
and U6478 (N_6478,N_6270,N_6362);
nand U6479 (N_6479,N_6227,N_6305);
nor U6480 (N_6480,N_6206,N_6209);
xnor U6481 (N_6481,N_6359,N_6214);
or U6482 (N_6482,N_6353,N_6331);
nor U6483 (N_6483,N_6205,N_6279);
or U6484 (N_6484,N_6264,N_6281);
nor U6485 (N_6485,N_6285,N_6243);
nand U6486 (N_6486,N_6257,N_6260);
or U6487 (N_6487,N_6292,N_6273);
or U6488 (N_6488,N_6354,N_6337);
and U6489 (N_6489,N_6208,N_6234);
or U6490 (N_6490,N_6327,N_6221);
nand U6491 (N_6491,N_6352,N_6304);
and U6492 (N_6492,N_6271,N_6245);
nand U6493 (N_6493,N_6388,N_6310);
or U6494 (N_6494,N_6294,N_6296);
or U6495 (N_6495,N_6323,N_6283);
and U6496 (N_6496,N_6393,N_6298);
nor U6497 (N_6497,N_6315,N_6324);
and U6498 (N_6498,N_6350,N_6231);
or U6499 (N_6499,N_6233,N_6399);
or U6500 (N_6500,N_6374,N_6359);
or U6501 (N_6501,N_6310,N_6289);
nand U6502 (N_6502,N_6214,N_6291);
nand U6503 (N_6503,N_6323,N_6296);
and U6504 (N_6504,N_6360,N_6257);
or U6505 (N_6505,N_6294,N_6267);
nand U6506 (N_6506,N_6379,N_6216);
or U6507 (N_6507,N_6258,N_6253);
nor U6508 (N_6508,N_6258,N_6348);
nor U6509 (N_6509,N_6244,N_6258);
nand U6510 (N_6510,N_6224,N_6234);
and U6511 (N_6511,N_6234,N_6325);
and U6512 (N_6512,N_6287,N_6203);
nor U6513 (N_6513,N_6397,N_6358);
or U6514 (N_6514,N_6374,N_6263);
nor U6515 (N_6515,N_6288,N_6360);
nand U6516 (N_6516,N_6331,N_6371);
xor U6517 (N_6517,N_6281,N_6241);
or U6518 (N_6518,N_6380,N_6389);
nor U6519 (N_6519,N_6395,N_6278);
and U6520 (N_6520,N_6219,N_6367);
and U6521 (N_6521,N_6340,N_6212);
nand U6522 (N_6522,N_6261,N_6302);
nand U6523 (N_6523,N_6279,N_6368);
nor U6524 (N_6524,N_6242,N_6363);
or U6525 (N_6525,N_6338,N_6268);
nor U6526 (N_6526,N_6291,N_6395);
xnor U6527 (N_6527,N_6251,N_6332);
or U6528 (N_6528,N_6353,N_6364);
nand U6529 (N_6529,N_6297,N_6258);
and U6530 (N_6530,N_6391,N_6351);
or U6531 (N_6531,N_6218,N_6347);
and U6532 (N_6532,N_6373,N_6277);
nor U6533 (N_6533,N_6211,N_6303);
and U6534 (N_6534,N_6352,N_6367);
or U6535 (N_6535,N_6260,N_6292);
nor U6536 (N_6536,N_6312,N_6380);
and U6537 (N_6537,N_6356,N_6370);
and U6538 (N_6538,N_6319,N_6326);
nand U6539 (N_6539,N_6361,N_6262);
nand U6540 (N_6540,N_6244,N_6314);
nor U6541 (N_6541,N_6266,N_6385);
and U6542 (N_6542,N_6242,N_6333);
nor U6543 (N_6543,N_6201,N_6298);
nor U6544 (N_6544,N_6211,N_6282);
xnor U6545 (N_6545,N_6307,N_6237);
nand U6546 (N_6546,N_6393,N_6377);
or U6547 (N_6547,N_6268,N_6285);
nand U6548 (N_6548,N_6272,N_6218);
and U6549 (N_6549,N_6265,N_6320);
or U6550 (N_6550,N_6227,N_6267);
and U6551 (N_6551,N_6275,N_6316);
or U6552 (N_6552,N_6270,N_6247);
and U6553 (N_6553,N_6296,N_6328);
nand U6554 (N_6554,N_6260,N_6334);
and U6555 (N_6555,N_6272,N_6332);
nand U6556 (N_6556,N_6326,N_6262);
nand U6557 (N_6557,N_6223,N_6350);
or U6558 (N_6558,N_6371,N_6265);
nand U6559 (N_6559,N_6205,N_6328);
nand U6560 (N_6560,N_6336,N_6290);
nand U6561 (N_6561,N_6313,N_6329);
nor U6562 (N_6562,N_6357,N_6389);
or U6563 (N_6563,N_6283,N_6383);
and U6564 (N_6564,N_6328,N_6390);
xor U6565 (N_6565,N_6391,N_6320);
nor U6566 (N_6566,N_6265,N_6237);
nand U6567 (N_6567,N_6331,N_6378);
nand U6568 (N_6568,N_6334,N_6365);
nand U6569 (N_6569,N_6204,N_6221);
and U6570 (N_6570,N_6310,N_6315);
or U6571 (N_6571,N_6366,N_6367);
nor U6572 (N_6572,N_6392,N_6298);
nand U6573 (N_6573,N_6395,N_6296);
nand U6574 (N_6574,N_6243,N_6316);
and U6575 (N_6575,N_6300,N_6357);
or U6576 (N_6576,N_6345,N_6386);
nand U6577 (N_6577,N_6361,N_6249);
and U6578 (N_6578,N_6259,N_6257);
nand U6579 (N_6579,N_6285,N_6250);
nand U6580 (N_6580,N_6262,N_6257);
and U6581 (N_6581,N_6241,N_6254);
and U6582 (N_6582,N_6345,N_6361);
nor U6583 (N_6583,N_6348,N_6202);
and U6584 (N_6584,N_6294,N_6306);
or U6585 (N_6585,N_6370,N_6391);
and U6586 (N_6586,N_6291,N_6224);
nand U6587 (N_6587,N_6286,N_6245);
nand U6588 (N_6588,N_6335,N_6367);
nor U6589 (N_6589,N_6277,N_6287);
nand U6590 (N_6590,N_6205,N_6384);
nor U6591 (N_6591,N_6297,N_6206);
xnor U6592 (N_6592,N_6279,N_6208);
and U6593 (N_6593,N_6320,N_6222);
and U6594 (N_6594,N_6312,N_6201);
or U6595 (N_6595,N_6336,N_6204);
nand U6596 (N_6596,N_6288,N_6341);
nor U6597 (N_6597,N_6392,N_6356);
nand U6598 (N_6598,N_6276,N_6333);
and U6599 (N_6599,N_6323,N_6235);
nor U6600 (N_6600,N_6518,N_6595);
nand U6601 (N_6601,N_6521,N_6548);
nor U6602 (N_6602,N_6416,N_6583);
nor U6603 (N_6603,N_6542,N_6468);
or U6604 (N_6604,N_6460,N_6477);
nor U6605 (N_6605,N_6492,N_6496);
nor U6606 (N_6606,N_6424,N_6533);
and U6607 (N_6607,N_6463,N_6408);
and U6608 (N_6608,N_6598,N_6505);
and U6609 (N_6609,N_6440,N_6423);
nor U6610 (N_6610,N_6565,N_6459);
and U6611 (N_6611,N_6596,N_6462);
nor U6612 (N_6612,N_6495,N_6502);
or U6613 (N_6613,N_6453,N_6588);
nor U6614 (N_6614,N_6592,N_6488);
nand U6615 (N_6615,N_6456,N_6470);
and U6616 (N_6616,N_6524,N_6482);
or U6617 (N_6617,N_6513,N_6597);
or U6618 (N_6618,N_6486,N_6577);
nand U6619 (N_6619,N_6404,N_6479);
or U6620 (N_6620,N_6568,N_6443);
nand U6621 (N_6621,N_6579,N_6528);
nand U6622 (N_6622,N_6422,N_6428);
and U6623 (N_6623,N_6410,N_6584);
and U6624 (N_6624,N_6514,N_6447);
nor U6625 (N_6625,N_6566,N_6570);
and U6626 (N_6626,N_6498,N_6549);
nor U6627 (N_6627,N_6580,N_6523);
or U6628 (N_6628,N_6541,N_6593);
and U6629 (N_6629,N_6535,N_6575);
nor U6630 (N_6630,N_6510,N_6538);
nor U6631 (N_6631,N_6519,N_6474);
nor U6632 (N_6632,N_6411,N_6490);
and U6633 (N_6633,N_6589,N_6429);
or U6634 (N_6634,N_6517,N_6537);
nor U6635 (N_6635,N_6400,N_6473);
nor U6636 (N_6636,N_6586,N_6417);
nor U6637 (N_6637,N_6539,N_6527);
and U6638 (N_6638,N_6415,N_6525);
and U6639 (N_6639,N_6483,N_6599);
and U6640 (N_6640,N_6493,N_6434);
xor U6641 (N_6641,N_6564,N_6455);
or U6642 (N_6642,N_6469,N_6466);
and U6643 (N_6643,N_6420,N_6436);
and U6644 (N_6644,N_6438,N_6439);
or U6645 (N_6645,N_6421,N_6574);
xor U6646 (N_6646,N_6414,N_6501);
and U6647 (N_6647,N_6405,N_6557);
nand U6648 (N_6648,N_6441,N_6550);
nor U6649 (N_6649,N_6465,N_6581);
and U6650 (N_6650,N_6452,N_6431);
nand U6651 (N_6651,N_6526,N_6484);
or U6652 (N_6652,N_6426,N_6409);
nor U6653 (N_6653,N_6476,N_6532);
or U6654 (N_6654,N_6487,N_6412);
and U6655 (N_6655,N_6512,N_6552);
nor U6656 (N_6656,N_6454,N_6448);
and U6657 (N_6657,N_6427,N_6497);
or U6658 (N_6658,N_6554,N_6572);
or U6659 (N_6659,N_6500,N_6590);
nor U6660 (N_6660,N_6582,N_6445);
or U6661 (N_6661,N_6534,N_6419);
and U6662 (N_6662,N_6467,N_6413);
or U6663 (N_6663,N_6499,N_6560);
nor U6664 (N_6664,N_6418,N_6402);
nor U6665 (N_6665,N_6457,N_6444);
nor U6666 (N_6666,N_6449,N_6451);
and U6667 (N_6667,N_6585,N_6491);
and U6668 (N_6668,N_6571,N_6540);
and U6669 (N_6669,N_6458,N_6503);
or U6670 (N_6670,N_6489,N_6531);
nand U6671 (N_6671,N_6536,N_6561);
nor U6672 (N_6672,N_6558,N_6546);
and U6673 (N_6673,N_6569,N_6432);
nor U6674 (N_6674,N_6515,N_6407);
and U6675 (N_6675,N_6430,N_6506);
xor U6676 (N_6676,N_6509,N_6578);
or U6677 (N_6677,N_6401,N_6433);
or U6678 (N_6678,N_6591,N_6544);
or U6679 (N_6679,N_6480,N_6522);
nor U6680 (N_6680,N_6573,N_6547);
and U6681 (N_6681,N_6516,N_6437);
nor U6682 (N_6682,N_6511,N_6494);
and U6683 (N_6683,N_6471,N_6461);
and U6684 (N_6684,N_6485,N_6504);
and U6685 (N_6685,N_6406,N_6478);
nor U6686 (N_6686,N_6553,N_6545);
and U6687 (N_6687,N_6543,N_6464);
nor U6688 (N_6688,N_6529,N_6563);
nand U6689 (N_6689,N_6450,N_6556);
nand U6690 (N_6690,N_6435,N_6594);
or U6691 (N_6691,N_6559,N_6425);
nor U6692 (N_6692,N_6530,N_6562);
nand U6693 (N_6693,N_6507,N_6567);
nor U6694 (N_6694,N_6551,N_6555);
or U6695 (N_6695,N_6520,N_6472);
or U6696 (N_6696,N_6481,N_6475);
and U6697 (N_6697,N_6587,N_6576);
nand U6698 (N_6698,N_6442,N_6508);
or U6699 (N_6699,N_6403,N_6446);
or U6700 (N_6700,N_6599,N_6458);
nor U6701 (N_6701,N_6573,N_6583);
or U6702 (N_6702,N_6571,N_6569);
nand U6703 (N_6703,N_6570,N_6476);
nand U6704 (N_6704,N_6589,N_6585);
and U6705 (N_6705,N_6428,N_6459);
nor U6706 (N_6706,N_6501,N_6527);
or U6707 (N_6707,N_6444,N_6530);
nand U6708 (N_6708,N_6498,N_6468);
and U6709 (N_6709,N_6431,N_6426);
nor U6710 (N_6710,N_6405,N_6567);
nor U6711 (N_6711,N_6453,N_6574);
or U6712 (N_6712,N_6411,N_6529);
nand U6713 (N_6713,N_6487,N_6484);
and U6714 (N_6714,N_6469,N_6461);
nor U6715 (N_6715,N_6535,N_6572);
nor U6716 (N_6716,N_6483,N_6434);
nand U6717 (N_6717,N_6531,N_6422);
nand U6718 (N_6718,N_6516,N_6596);
nor U6719 (N_6719,N_6547,N_6570);
nand U6720 (N_6720,N_6558,N_6531);
and U6721 (N_6721,N_6505,N_6439);
nor U6722 (N_6722,N_6506,N_6528);
nand U6723 (N_6723,N_6579,N_6466);
and U6724 (N_6724,N_6587,N_6463);
nor U6725 (N_6725,N_6539,N_6520);
nor U6726 (N_6726,N_6554,N_6517);
nor U6727 (N_6727,N_6523,N_6426);
xor U6728 (N_6728,N_6525,N_6595);
nand U6729 (N_6729,N_6546,N_6463);
and U6730 (N_6730,N_6530,N_6527);
and U6731 (N_6731,N_6539,N_6406);
nand U6732 (N_6732,N_6594,N_6597);
nand U6733 (N_6733,N_6500,N_6435);
xor U6734 (N_6734,N_6515,N_6402);
or U6735 (N_6735,N_6491,N_6543);
and U6736 (N_6736,N_6405,N_6545);
nand U6737 (N_6737,N_6575,N_6587);
or U6738 (N_6738,N_6441,N_6448);
and U6739 (N_6739,N_6588,N_6568);
nand U6740 (N_6740,N_6569,N_6413);
and U6741 (N_6741,N_6463,N_6499);
nand U6742 (N_6742,N_6500,N_6429);
nor U6743 (N_6743,N_6576,N_6543);
and U6744 (N_6744,N_6466,N_6515);
and U6745 (N_6745,N_6403,N_6432);
nor U6746 (N_6746,N_6575,N_6462);
nor U6747 (N_6747,N_6538,N_6571);
or U6748 (N_6748,N_6439,N_6502);
xnor U6749 (N_6749,N_6403,N_6501);
nor U6750 (N_6750,N_6576,N_6502);
nand U6751 (N_6751,N_6424,N_6513);
nor U6752 (N_6752,N_6519,N_6556);
or U6753 (N_6753,N_6498,N_6493);
nor U6754 (N_6754,N_6529,N_6489);
and U6755 (N_6755,N_6445,N_6579);
or U6756 (N_6756,N_6475,N_6589);
nand U6757 (N_6757,N_6588,N_6526);
nand U6758 (N_6758,N_6577,N_6564);
nor U6759 (N_6759,N_6514,N_6436);
or U6760 (N_6760,N_6483,N_6475);
and U6761 (N_6761,N_6479,N_6558);
nor U6762 (N_6762,N_6496,N_6451);
nor U6763 (N_6763,N_6591,N_6520);
and U6764 (N_6764,N_6592,N_6413);
or U6765 (N_6765,N_6420,N_6447);
nand U6766 (N_6766,N_6487,N_6449);
and U6767 (N_6767,N_6572,N_6478);
and U6768 (N_6768,N_6502,N_6432);
nor U6769 (N_6769,N_6451,N_6420);
and U6770 (N_6770,N_6535,N_6422);
nor U6771 (N_6771,N_6479,N_6482);
and U6772 (N_6772,N_6557,N_6419);
and U6773 (N_6773,N_6429,N_6543);
or U6774 (N_6774,N_6575,N_6544);
nand U6775 (N_6775,N_6404,N_6490);
nand U6776 (N_6776,N_6447,N_6515);
and U6777 (N_6777,N_6532,N_6560);
nand U6778 (N_6778,N_6590,N_6406);
and U6779 (N_6779,N_6449,N_6472);
nand U6780 (N_6780,N_6577,N_6553);
nor U6781 (N_6781,N_6538,N_6464);
nand U6782 (N_6782,N_6470,N_6425);
and U6783 (N_6783,N_6431,N_6537);
nand U6784 (N_6784,N_6403,N_6460);
nand U6785 (N_6785,N_6598,N_6418);
and U6786 (N_6786,N_6447,N_6526);
nand U6787 (N_6787,N_6570,N_6560);
and U6788 (N_6788,N_6424,N_6518);
and U6789 (N_6789,N_6490,N_6458);
nor U6790 (N_6790,N_6562,N_6489);
nor U6791 (N_6791,N_6576,N_6568);
nor U6792 (N_6792,N_6543,N_6532);
xor U6793 (N_6793,N_6435,N_6491);
nand U6794 (N_6794,N_6550,N_6471);
xnor U6795 (N_6795,N_6454,N_6499);
nand U6796 (N_6796,N_6429,N_6527);
or U6797 (N_6797,N_6593,N_6517);
nor U6798 (N_6798,N_6536,N_6420);
nand U6799 (N_6799,N_6511,N_6520);
nand U6800 (N_6800,N_6654,N_6736);
nor U6801 (N_6801,N_6638,N_6608);
or U6802 (N_6802,N_6613,N_6718);
or U6803 (N_6803,N_6730,N_6672);
nor U6804 (N_6804,N_6762,N_6693);
nor U6805 (N_6805,N_6729,N_6700);
and U6806 (N_6806,N_6734,N_6680);
or U6807 (N_6807,N_6669,N_6760);
and U6808 (N_6808,N_6755,N_6685);
or U6809 (N_6809,N_6739,N_6714);
nor U6810 (N_6810,N_6664,N_6780);
nand U6811 (N_6811,N_6742,N_6645);
nand U6812 (N_6812,N_6732,N_6644);
nor U6813 (N_6813,N_6646,N_6719);
nand U6814 (N_6814,N_6773,N_6601);
and U6815 (N_6815,N_6620,N_6692);
nor U6816 (N_6816,N_6699,N_6643);
nor U6817 (N_6817,N_6765,N_6694);
and U6818 (N_6818,N_6759,N_6763);
nand U6819 (N_6819,N_6631,N_6761);
and U6820 (N_6820,N_6662,N_6658);
and U6821 (N_6821,N_6798,N_6639);
nand U6822 (N_6822,N_6673,N_6728);
or U6823 (N_6823,N_6630,N_6784);
and U6824 (N_6824,N_6782,N_6723);
and U6825 (N_6825,N_6611,N_6791);
and U6826 (N_6826,N_6726,N_6741);
nor U6827 (N_6827,N_6768,N_6797);
nor U6828 (N_6828,N_6632,N_6668);
or U6829 (N_6829,N_6657,N_6640);
nand U6830 (N_6830,N_6665,N_6628);
nor U6831 (N_6831,N_6642,N_6724);
xor U6832 (N_6832,N_6676,N_6619);
and U6833 (N_6833,N_6648,N_6747);
or U6834 (N_6834,N_6604,N_6740);
and U6835 (N_6835,N_6627,N_6677);
and U6836 (N_6836,N_6702,N_6641);
and U6837 (N_6837,N_6622,N_6637);
or U6838 (N_6838,N_6603,N_6623);
nand U6839 (N_6839,N_6647,N_6697);
and U6840 (N_6840,N_6629,N_6616);
and U6841 (N_6841,N_6793,N_6653);
or U6842 (N_6842,N_6771,N_6756);
and U6843 (N_6843,N_6781,N_6750);
or U6844 (N_6844,N_6774,N_6683);
or U6845 (N_6845,N_6789,N_6712);
nor U6846 (N_6846,N_6650,N_6704);
and U6847 (N_6847,N_6696,N_6671);
or U6848 (N_6848,N_6711,N_6749);
nand U6849 (N_6849,N_6722,N_6799);
nand U6850 (N_6850,N_6667,N_6621);
and U6851 (N_6851,N_6635,N_6686);
or U6852 (N_6852,N_6720,N_6687);
or U6853 (N_6853,N_6618,N_6752);
or U6854 (N_6854,N_6701,N_6733);
nand U6855 (N_6855,N_6666,N_6717);
nor U6856 (N_6856,N_6675,N_6767);
and U6857 (N_6857,N_6745,N_6721);
or U6858 (N_6858,N_6754,N_6737);
and U6859 (N_6859,N_6612,N_6731);
nor U6860 (N_6860,N_6695,N_6624);
nor U6861 (N_6861,N_6769,N_6690);
and U6862 (N_6862,N_6698,N_6663);
and U6863 (N_6863,N_6649,N_6785);
and U6864 (N_6864,N_6625,N_6788);
and U6865 (N_6865,N_6707,N_6777);
and U6866 (N_6866,N_6681,N_6716);
nor U6867 (N_6867,N_6626,N_6783);
nor U6868 (N_6868,N_6751,N_6614);
or U6869 (N_6869,N_6706,N_6795);
or U6870 (N_6870,N_6682,N_6602);
nor U6871 (N_6871,N_6715,N_6670);
nand U6872 (N_6872,N_6794,N_6659);
nand U6873 (N_6873,N_6651,N_6636);
nor U6874 (N_6874,N_6776,N_6753);
and U6875 (N_6875,N_6766,N_6610);
nand U6876 (N_6876,N_6778,N_6674);
nand U6877 (N_6877,N_6617,N_6688);
nand U6878 (N_6878,N_6709,N_6727);
nor U6879 (N_6879,N_6713,N_6770);
nand U6880 (N_6880,N_6710,N_6746);
or U6881 (N_6881,N_6634,N_6691);
or U6882 (N_6882,N_6703,N_6633);
or U6883 (N_6883,N_6772,N_6689);
nor U6884 (N_6884,N_6792,N_6652);
nand U6885 (N_6885,N_6679,N_6725);
nor U6886 (N_6886,N_6758,N_6678);
nand U6887 (N_6887,N_6757,N_6779);
xor U6888 (N_6888,N_6743,N_6615);
and U6889 (N_6889,N_6660,N_6606);
or U6890 (N_6890,N_6605,N_6744);
and U6891 (N_6891,N_6684,N_6748);
and U6892 (N_6892,N_6656,N_6600);
nand U6893 (N_6893,N_6735,N_6607);
and U6894 (N_6894,N_6790,N_6796);
and U6895 (N_6895,N_6764,N_6661);
and U6896 (N_6896,N_6775,N_6655);
and U6897 (N_6897,N_6786,N_6609);
or U6898 (N_6898,N_6738,N_6708);
or U6899 (N_6899,N_6787,N_6705);
and U6900 (N_6900,N_6669,N_6633);
nor U6901 (N_6901,N_6696,N_6699);
and U6902 (N_6902,N_6685,N_6784);
or U6903 (N_6903,N_6763,N_6620);
and U6904 (N_6904,N_6618,N_6710);
or U6905 (N_6905,N_6607,N_6772);
nand U6906 (N_6906,N_6654,N_6624);
nand U6907 (N_6907,N_6687,N_6608);
or U6908 (N_6908,N_6732,N_6761);
nand U6909 (N_6909,N_6625,N_6617);
or U6910 (N_6910,N_6769,N_6684);
or U6911 (N_6911,N_6752,N_6757);
and U6912 (N_6912,N_6778,N_6726);
nor U6913 (N_6913,N_6798,N_6626);
or U6914 (N_6914,N_6699,N_6691);
or U6915 (N_6915,N_6773,N_6779);
or U6916 (N_6916,N_6688,N_6707);
nand U6917 (N_6917,N_6652,N_6769);
nand U6918 (N_6918,N_6759,N_6710);
and U6919 (N_6919,N_6658,N_6604);
nand U6920 (N_6920,N_6766,N_6618);
nand U6921 (N_6921,N_6798,N_6729);
nor U6922 (N_6922,N_6611,N_6732);
nand U6923 (N_6923,N_6614,N_6794);
and U6924 (N_6924,N_6720,N_6732);
or U6925 (N_6925,N_6632,N_6604);
and U6926 (N_6926,N_6655,N_6611);
nor U6927 (N_6927,N_6776,N_6650);
or U6928 (N_6928,N_6670,N_6730);
nor U6929 (N_6929,N_6682,N_6709);
nor U6930 (N_6930,N_6600,N_6758);
nor U6931 (N_6931,N_6747,N_6791);
or U6932 (N_6932,N_6771,N_6608);
nor U6933 (N_6933,N_6750,N_6757);
nor U6934 (N_6934,N_6663,N_6731);
or U6935 (N_6935,N_6712,N_6614);
nor U6936 (N_6936,N_6635,N_6777);
nor U6937 (N_6937,N_6660,N_6600);
and U6938 (N_6938,N_6749,N_6640);
nand U6939 (N_6939,N_6688,N_6693);
nand U6940 (N_6940,N_6762,N_6689);
nand U6941 (N_6941,N_6695,N_6745);
or U6942 (N_6942,N_6731,N_6651);
xnor U6943 (N_6943,N_6724,N_6603);
or U6944 (N_6944,N_6742,N_6611);
nand U6945 (N_6945,N_6747,N_6746);
and U6946 (N_6946,N_6626,N_6746);
xnor U6947 (N_6947,N_6673,N_6782);
and U6948 (N_6948,N_6687,N_6781);
and U6949 (N_6949,N_6672,N_6768);
xor U6950 (N_6950,N_6754,N_6648);
and U6951 (N_6951,N_6701,N_6660);
and U6952 (N_6952,N_6741,N_6678);
nor U6953 (N_6953,N_6731,N_6727);
nor U6954 (N_6954,N_6648,N_6720);
nor U6955 (N_6955,N_6702,N_6654);
or U6956 (N_6956,N_6781,N_6600);
nor U6957 (N_6957,N_6738,N_6710);
or U6958 (N_6958,N_6732,N_6673);
and U6959 (N_6959,N_6657,N_6757);
or U6960 (N_6960,N_6795,N_6654);
and U6961 (N_6961,N_6694,N_6690);
nand U6962 (N_6962,N_6717,N_6698);
and U6963 (N_6963,N_6783,N_6722);
nand U6964 (N_6964,N_6734,N_6672);
or U6965 (N_6965,N_6651,N_6756);
nand U6966 (N_6966,N_6697,N_6691);
or U6967 (N_6967,N_6616,N_6656);
nand U6968 (N_6968,N_6646,N_6784);
nor U6969 (N_6969,N_6696,N_6628);
nor U6970 (N_6970,N_6639,N_6680);
nor U6971 (N_6971,N_6611,N_6692);
nor U6972 (N_6972,N_6624,N_6717);
or U6973 (N_6973,N_6791,N_6661);
nor U6974 (N_6974,N_6697,N_6769);
or U6975 (N_6975,N_6712,N_6651);
or U6976 (N_6976,N_6733,N_6667);
xnor U6977 (N_6977,N_6689,N_6678);
or U6978 (N_6978,N_6661,N_6693);
or U6979 (N_6979,N_6672,N_6735);
nor U6980 (N_6980,N_6742,N_6702);
nand U6981 (N_6981,N_6744,N_6610);
and U6982 (N_6982,N_6618,N_6761);
nand U6983 (N_6983,N_6726,N_6786);
and U6984 (N_6984,N_6730,N_6684);
nor U6985 (N_6985,N_6630,N_6793);
nor U6986 (N_6986,N_6743,N_6610);
and U6987 (N_6987,N_6769,N_6622);
or U6988 (N_6988,N_6698,N_6645);
nand U6989 (N_6989,N_6641,N_6789);
or U6990 (N_6990,N_6745,N_6707);
nand U6991 (N_6991,N_6752,N_6759);
or U6992 (N_6992,N_6708,N_6750);
xnor U6993 (N_6993,N_6777,N_6747);
and U6994 (N_6994,N_6713,N_6604);
nand U6995 (N_6995,N_6636,N_6698);
nand U6996 (N_6996,N_6738,N_6620);
xnor U6997 (N_6997,N_6689,N_6705);
nor U6998 (N_6998,N_6695,N_6719);
and U6999 (N_6999,N_6758,N_6753);
and U7000 (N_7000,N_6850,N_6889);
xor U7001 (N_7001,N_6874,N_6817);
nor U7002 (N_7002,N_6882,N_6894);
nor U7003 (N_7003,N_6860,N_6859);
nor U7004 (N_7004,N_6823,N_6966);
or U7005 (N_7005,N_6938,N_6910);
nand U7006 (N_7006,N_6901,N_6813);
xnor U7007 (N_7007,N_6847,N_6810);
nor U7008 (N_7008,N_6892,N_6825);
and U7009 (N_7009,N_6855,N_6861);
or U7010 (N_7010,N_6956,N_6964);
nor U7011 (N_7011,N_6819,N_6939);
and U7012 (N_7012,N_6816,N_6934);
or U7013 (N_7013,N_6880,N_6987);
nor U7014 (N_7014,N_6830,N_6923);
nand U7015 (N_7015,N_6862,N_6871);
nand U7016 (N_7016,N_6919,N_6804);
nand U7017 (N_7017,N_6865,N_6856);
or U7018 (N_7018,N_6972,N_6922);
nor U7019 (N_7019,N_6989,N_6867);
nand U7020 (N_7020,N_6936,N_6970);
nor U7021 (N_7021,N_6916,N_6809);
or U7022 (N_7022,N_6808,N_6866);
or U7023 (N_7023,N_6841,N_6986);
nand U7024 (N_7024,N_6974,N_6891);
nor U7025 (N_7025,N_6828,N_6975);
or U7026 (N_7026,N_6831,N_6952);
nor U7027 (N_7027,N_6877,N_6949);
nand U7028 (N_7028,N_6931,N_6800);
or U7029 (N_7029,N_6821,N_6929);
nor U7030 (N_7030,N_6979,N_6839);
and U7031 (N_7031,N_6999,N_6812);
nor U7032 (N_7032,N_6824,N_6961);
or U7033 (N_7033,N_6927,N_6953);
nand U7034 (N_7034,N_6945,N_6838);
nand U7035 (N_7035,N_6988,N_6958);
xnor U7036 (N_7036,N_6886,N_6947);
xor U7037 (N_7037,N_6982,N_6976);
or U7038 (N_7038,N_6965,N_6849);
and U7039 (N_7039,N_6924,N_6876);
or U7040 (N_7040,N_6930,N_6951);
or U7041 (N_7041,N_6888,N_6920);
nor U7042 (N_7042,N_6864,N_6932);
and U7043 (N_7043,N_6883,N_6815);
or U7044 (N_7044,N_6852,N_6943);
nand U7045 (N_7045,N_6848,N_6902);
nor U7046 (N_7046,N_6907,N_6983);
and U7047 (N_7047,N_6844,N_6857);
and U7048 (N_7048,N_6806,N_6996);
and U7049 (N_7049,N_6829,N_6834);
nor U7050 (N_7050,N_6840,N_6833);
nor U7051 (N_7051,N_6909,N_6915);
nor U7052 (N_7052,N_6969,N_6926);
xnor U7053 (N_7053,N_6863,N_6851);
nor U7054 (N_7054,N_6942,N_6873);
nor U7055 (N_7055,N_6832,N_6913);
and U7056 (N_7056,N_6978,N_6904);
nand U7057 (N_7057,N_6898,N_6995);
or U7058 (N_7058,N_6890,N_6971);
nand U7059 (N_7059,N_6807,N_6903);
nand U7060 (N_7060,N_6955,N_6994);
and U7061 (N_7061,N_6993,N_6811);
nand U7062 (N_7062,N_6899,N_6820);
or U7063 (N_7063,N_6940,N_6973);
nor U7064 (N_7064,N_6879,N_6984);
or U7065 (N_7065,N_6925,N_6917);
and U7066 (N_7066,N_6805,N_6845);
or U7067 (N_7067,N_6826,N_6950);
or U7068 (N_7068,N_6928,N_6944);
or U7069 (N_7069,N_6963,N_6985);
nand U7070 (N_7070,N_6908,N_6954);
nand U7071 (N_7071,N_6843,N_6992);
or U7072 (N_7072,N_6977,N_6827);
and U7073 (N_7073,N_6937,N_6959);
or U7074 (N_7074,N_6980,N_6941);
and U7075 (N_7075,N_6875,N_6935);
or U7076 (N_7076,N_6962,N_6835);
nor U7077 (N_7077,N_6887,N_6968);
xnor U7078 (N_7078,N_6911,N_6893);
or U7079 (N_7079,N_6991,N_6858);
or U7080 (N_7080,N_6998,N_6960);
nor U7081 (N_7081,N_6905,N_6884);
and U7082 (N_7082,N_6868,N_6933);
or U7083 (N_7083,N_6818,N_6853);
and U7084 (N_7084,N_6842,N_6869);
and U7085 (N_7085,N_6802,N_6881);
nand U7086 (N_7086,N_6990,N_6897);
and U7087 (N_7087,N_6885,N_6814);
nor U7088 (N_7088,N_6967,N_6895);
nor U7089 (N_7089,N_6912,N_6836);
nor U7090 (N_7090,N_6946,N_6981);
or U7091 (N_7091,N_6872,N_6837);
or U7092 (N_7092,N_6846,N_6878);
nand U7093 (N_7093,N_6900,N_6906);
and U7094 (N_7094,N_6822,N_6803);
and U7095 (N_7095,N_6997,N_6948);
nor U7096 (N_7096,N_6854,N_6914);
and U7097 (N_7097,N_6921,N_6957);
or U7098 (N_7098,N_6918,N_6870);
nor U7099 (N_7099,N_6896,N_6801);
and U7100 (N_7100,N_6881,N_6871);
nand U7101 (N_7101,N_6856,N_6845);
nor U7102 (N_7102,N_6804,N_6889);
or U7103 (N_7103,N_6928,N_6964);
and U7104 (N_7104,N_6903,N_6932);
nor U7105 (N_7105,N_6970,N_6812);
and U7106 (N_7106,N_6914,N_6838);
nor U7107 (N_7107,N_6922,N_6839);
nand U7108 (N_7108,N_6889,N_6970);
and U7109 (N_7109,N_6810,N_6892);
nor U7110 (N_7110,N_6983,N_6932);
nand U7111 (N_7111,N_6801,N_6961);
nand U7112 (N_7112,N_6998,N_6813);
and U7113 (N_7113,N_6977,N_6843);
nand U7114 (N_7114,N_6924,N_6850);
nand U7115 (N_7115,N_6923,N_6808);
nand U7116 (N_7116,N_6982,N_6915);
nor U7117 (N_7117,N_6881,N_6909);
xor U7118 (N_7118,N_6951,N_6848);
or U7119 (N_7119,N_6819,N_6914);
xor U7120 (N_7120,N_6811,N_6863);
nor U7121 (N_7121,N_6892,N_6952);
or U7122 (N_7122,N_6962,N_6856);
nand U7123 (N_7123,N_6874,N_6869);
nor U7124 (N_7124,N_6866,N_6969);
nor U7125 (N_7125,N_6905,N_6828);
or U7126 (N_7126,N_6825,N_6831);
nor U7127 (N_7127,N_6811,N_6810);
or U7128 (N_7128,N_6970,N_6816);
nand U7129 (N_7129,N_6840,N_6817);
nor U7130 (N_7130,N_6868,N_6952);
and U7131 (N_7131,N_6972,N_6921);
nand U7132 (N_7132,N_6805,N_6891);
nand U7133 (N_7133,N_6820,N_6861);
xnor U7134 (N_7134,N_6829,N_6912);
nand U7135 (N_7135,N_6982,N_6922);
and U7136 (N_7136,N_6880,N_6863);
or U7137 (N_7137,N_6826,N_6954);
nor U7138 (N_7138,N_6853,N_6810);
and U7139 (N_7139,N_6960,N_6961);
or U7140 (N_7140,N_6928,N_6828);
and U7141 (N_7141,N_6816,N_6847);
or U7142 (N_7142,N_6876,N_6918);
nor U7143 (N_7143,N_6902,N_6840);
or U7144 (N_7144,N_6825,N_6879);
and U7145 (N_7145,N_6884,N_6984);
or U7146 (N_7146,N_6952,N_6819);
and U7147 (N_7147,N_6828,N_6833);
nor U7148 (N_7148,N_6922,N_6874);
and U7149 (N_7149,N_6979,N_6936);
and U7150 (N_7150,N_6893,N_6945);
nor U7151 (N_7151,N_6955,N_6907);
or U7152 (N_7152,N_6848,N_6800);
nor U7153 (N_7153,N_6878,N_6887);
or U7154 (N_7154,N_6903,N_6859);
or U7155 (N_7155,N_6887,N_6888);
nor U7156 (N_7156,N_6990,N_6823);
and U7157 (N_7157,N_6930,N_6869);
nand U7158 (N_7158,N_6916,N_6993);
and U7159 (N_7159,N_6962,N_6939);
or U7160 (N_7160,N_6827,N_6904);
and U7161 (N_7161,N_6969,N_6949);
nand U7162 (N_7162,N_6902,N_6903);
and U7163 (N_7163,N_6981,N_6809);
and U7164 (N_7164,N_6834,N_6832);
xnor U7165 (N_7165,N_6910,N_6966);
or U7166 (N_7166,N_6829,N_6827);
and U7167 (N_7167,N_6849,N_6963);
nor U7168 (N_7168,N_6872,N_6949);
or U7169 (N_7169,N_6960,N_6910);
nor U7170 (N_7170,N_6929,N_6908);
and U7171 (N_7171,N_6903,N_6941);
and U7172 (N_7172,N_6877,N_6805);
nor U7173 (N_7173,N_6852,N_6978);
nor U7174 (N_7174,N_6896,N_6840);
or U7175 (N_7175,N_6977,N_6803);
xnor U7176 (N_7176,N_6940,N_6949);
and U7177 (N_7177,N_6951,N_6884);
nand U7178 (N_7178,N_6955,N_6927);
or U7179 (N_7179,N_6952,N_6821);
and U7180 (N_7180,N_6803,N_6902);
and U7181 (N_7181,N_6980,N_6819);
nand U7182 (N_7182,N_6861,N_6860);
nor U7183 (N_7183,N_6969,N_6997);
and U7184 (N_7184,N_6912,N_6828);
nand U7185 (N_7185,N_6945,N_6987);
nand U7186 (N_7186,N_6929,N_6823);
nand U7187 (N_7187,N_6957,N_6913);
or U7188 (N_7188,N_6843,N_6831);
nand U7189 (N_7189,N_6913,N_6830);
nand U7190 (N_7190,N_6987,N_6845);
nand U7191 (N_7191,N_6963,N_6881);
nand U7192 (N_7192,N_6930,N_6942);
and U7193 (N_7193,N_6929,N_6853);
or U7194 (N_7194,N_6849,N_6867);
nand U7195 (N_7195,N_6832,N_6859);
nand U7196 (N_7196,N_6937,N_6905);
and U7197 (N_7197,N_6999,N_6854);
nor U7198 (N_7198,N_6954,N_6834);
and U7199 (N_7199,N_6807,N_6951);
nand U7200 (N_7200,N_7039,N_7175);
nand U7201 (N_7201,N_7045,N_7172);
and U7202 (N_7202,N_7120,N_7068);
nand U7203 (N_7203,N_7001,N_7078);
and U7204 (N_7204,N_7171,N_7033);
or U7205 (N_7205,N_7061,N_7198);
nor U7206 (N_7206,N_7123,N_7142);
or U7207 (N_7207,N_7183,N_7153);
or U7208 (N_7208,N_7155,N_7151);
and U7209 (N_7209,N_7100,N_7020);
and U7210 (N_7210,N_7014,N_7138);
and U7211 (N_7211,N_7169,N_7057);
or U7212 (N_7212,N_7017,N_7085);
or U7213 (N_7213,N_7009,N_7192);
or U7214 (N_7214,N_7161,N_7047);
nand U7215 (N_7215,N_7102,N_7093);
and U7216 (N_7216,N_7190,N_7181);
and U7217 (N_7217,N_7187,N_7165);
nand U7218 (N_7218,N_7133,N_7177);
and U7219 (N_7219,N_7074,N_7111);
nor U7220 (N_7220,N_7130,N_7089);
or U7221 (N_7221,N_7106,N_7052);
and U7222 (N_7222,N_7013,N_7070);
nor U7223 (N_7223,N_7140,N_7135);
nor U7224 (N_7224,N_7146,N_7095);
and U7225 (N_7225,N_7159,N_7029);
nor U7226 (N_7226,N_7067,N_7096);
or U7227 (N_7227,N_7050,N_7041);
or U7228 (N_7228,N_7066,N_7031);
or U7229 (N_7229,N_7145,N_7026);
nand U7230 (N_7230,N_7122,N_7019);
nand U7231 (N_7231,N_7083,N_7079);
and U7232 (N_7232,N_7090,N_7134);
nor U7233 (N_7233,N_7035,N_7113);
nor U7234 (N_7234,N_7154,N_7160);
and U7235 (N_7235,N_7104,N_7166);
nor U7236 (N_7236,N_7034,N_7197);
nor U7237 (N_7237,N_7191,N_7005);
nand U7238 (N_7238,N_7038,N_7081);
and U7239 (N_7239,N_7099,N_7127);
and U7240 (N_7240,N_7139,N_7164);
and U7241 (N_7241,N_7162,N_7170);
nor U7242 (N_7242,N_7054,N_7037);
or U7243 (N_7243,N_7118,N_7132);
and U7244 (N_7244,N_7152,N_7024);
nand U7245 (N_7245,N_7015,N_7101);
nor U7246 (N_7246,N_7195,N_7189);
nand U7247 (N_7247,N_7023,N_7163);
and U7248 (N_7248,N_7012,N_7143);
nand U7249 (N_7249,N_7114,N_7056);
nand U7250 (N_7250,N_7109,N_7178);
or U7251 (N_7251,N_7076,N_7018);
nor U7252 (N_7252,N_7137,N_7084);
nand U7253 (N_7253,N_7124,N_7174);
or U7254 (N_7254,N_7046,N_7088);
nor U7255 (N_7255,N_7129,N_7125);
or U7256 (N_7256,N_7179,N_7149);
and U7257 (N_7257,N_7199,N_7107);
or U7258 (N_7258,N_7051,N_7021);
nor U7259 (N_7259,N_7119,N_7182);
nand U7260 (N_7260,N_7042,N_7004);
nand U7261 (N_7261,N_7011,N_7144);
nand U7262 (N_7262,N_7028,N_7006);
nand U7263 (N_7263,N_7072,N_7156);
nand U7264 (N_7264,N_7044,N_7168);
nor U7265 (N_7265,N_7116,N_7173);
or U7266 (N_7266,N_7059,N_7000);
or U7267 (N_7267,N_7105,N_7071);
nand U7268 (N_7268,N_7002,N_7049);
nor U7269 (N_7269,N_7080,N_7043);
and U7270 (N_7270,N_7087,N_7131);
nand U7271 (N_7271,N_7091,N_7053);
nor U7272 (N_7272,N_7110,N_7060);
and U7273 (N_7273,N_7128,N_7036);
and U7274 (N_7274,N_7186,N_7062);
and U7275 (N_7275,N_7196,N_7008);
and U7276 (N_7276,N_7030,N_7027);
nor U7277 (N_7277,N_7176,N_7082);
nor U7278 (N_7278,N_7077,N_7048);
nand U7279 (N_7279,N_7184,N_7188);
or U7280 (N_7280,N_7136,N_7086);
nor U7281 (N_7281,N_7016,N_7115);
nor U7282 (N_7282,N_7065,N_7003);
nand U7283 (N_7283,N_7147,N_7112);
xor U7284 (N_7284,N_7022,N_7073);
nor U7285 (N_7285,N_7007,N_7055);
nand U7286 (N_7286,N_7094,N_7069);
or U7287 (N_7287,N_7058,N_7010);
and U7288 (N_7288,N_7185,N_7040);
or U7289 (N_7289,N_7193,N_7167);
or U7290 (N_7290,N_7064,N_7063);
nor U7291 (N_7291,N_7180,N_7092);
nor U7292 (N_7292,N_7025,N_7103);
nor U7293 (N_7293,N_7121,N_7157);
nor U7294 (N_7294,N_7148,N_7194);
nand U7295 (N_7295,N_7075,N_7141);
and U7296 (N_7296,N_7126,N_7117);
nor U7297 (N_7297,N_7098,N_7150);
and U7298 (N_7298,N_7032,N_7097);
nor U7299 (N_7299,N_7158,N_7108);
nand U7300 (N_7300,N_7199,N_7118);
nor U7301 (N_7301,N_7183,N_7102);
nor U7302 (N_7302,N_7085,N_7117);
nor U7303 (N_7303,N_7186,N_7067);
xnor U7304 (N_7304,N_7112,N_7113);
or U7305 (N_7305,N_7059,N_7163);
nor U7306 (N_7306,N_7090,N_7183);
or U7307 (N_7307,N_7098,N_7045);
nand U7308 (N_7308,N_7027,N_7195);
nor U7309 (N_7309,N_7103,N_7067);
and U7310 (N_7310,N_7035,N_7174);
nand U7311 (N_7311,N_7033,N_7054);
and U7312 (N_7312,N_7133,N_7079);
and U7313 (N_7313,N_7178,N_7137);
or U7314 (N_7314,N_7120,N_7179);
and U7315 (N_7315,N_7195,N_7194);
and U7316 (N_7316,N_7196,N_7146);
nand U7317 (N_7317,N_7080,N_7134);
or U7318 (N_7318,N_7025,N_7091);
nor U7319 (N_7319,N_7032,N_7134);
nand U7320 (N_7320,N_7192,N_7077);
nand U7321 (N_7321,N_7196,N_7126);
and U7322 (N_7322,N_7039,N_7064);
and U7323 (N_7323,N_7066,N_7004);
and U7324 (N_7324,N_7159,N_7062);
nor U7325 (N_7325,N_7052,N_7143);
nand U7326 (N_7326,N_7016,N_7003);
or U7327 (N_7327,N_7002,N_7155);
and U7328 (N_7328,N_7143,N_7138);
nor U7329 (N_7329,N_7179,N_7087);
and U7330 (N_7330,N_7079,N_7005);
nor U7331 (N_7331,N_7045,N_7169);
nand U7332 (N_7332,N_7060,N_7140);
or U7333 (N_7333,N_7110,N_7113);
xor U7334 (N_7334,N_7162,N_7112);
nand U7335 (N_7335,N_7167,N_7133);
and U7336 (N_7336,N_7060,N_7067);
nand U7337 (N_7337,N_7190,N_7029);
nor U7338 (N_7338,N_7071,N_7193);
xor U7339 (N_7339,N_7117,N_7133);
nand U7340 (N_7340,N_7121,N_7099);
or U7341 (N_7341,N_7069,N_7118);
or U7342 (N_7342,N_7005,N_7106);
nand U7343 (N_7343,N_7085,N_7155);
and U7344 (N_7344,N_7114,N_7138);
or U7345 (N_7345,N_7098,N_7103);
nor U7346 (N_7346,N_7035,N_7082);
xnor U7347 (N_7347,N_7094,N_7142);
nor U7348 (N_7348,N_7167,N_7034);
and U7349 (N_7349,N_7103,N_7011);
or U7350 (N_7350,N_7056,N_7097);
nor U7351 (N_7351,N_7193,N_7137);
nand U7352 (N_7352,N_7070,N_7110);
nand U7353 (N_7353,N_7140,N_7069);
and U7354 (N_7354,N_7106,N_7003);
nand U7355 (N_7355,N_7145,N_7086);
or U7356 (N_7356,N_7072,N_7077);
or U7357 (N_7357,N_7105,N_7140);
and U7358 (N_7358,N_7034,N_7187);
or U7359 (N_7359,N_7094,N_7165);
or U7360 (N_7360,N_7162,N_7033);
or U7361 (N_7361,N_7087,N_7025);
nand U7362 (N_7362,N_7175,N_7129);
nor U7363 (N_7363,N_7052,N_7150);
and U7364 (N_7364,N_7036,N_7078);
or U7365 (N_7365,N_7100,N_7105);
nor U7366 (N_7366,N_7166,N_7172);
nor U7367 (N_7367,N_7076,N_7008);
xnor U7368 (N_7368,N_7094,N_7123);
nor U7369 (N_7369,N_7158,N_7082);
nor U7370 (N_7370,N_7118,N_7127);
nand U7371 (N_7371,N_7093,N_7068);
or U7372 (N_7372,N_7091,N_7102);
nor U7373 (N_7373,N_7020,N_7094);
or U7374 (N_7374,N_7007,N_7098);
or U7375 (N_7375,N_7110,N_7040);
and U7376 (N_7376,N_7102,N_7166);
nor U7377 (N_7377,N_7121,N_7112);
nand U7378 (N_7378,N_7055,N_7027);
nand U7379 (N_7379,N_7097,N_7121);
or U7380 (N_7380,N_7197,N_7042);
and U7381 (N_7381,N_7131,N_7133);
and U7382 (N_7382,N_7011,N_7115);
nor U7383 (N_7383,N_7143,N_7059);
nor U7384 (N_7384,N_7079,N_7120);
nand U7385 (N_7385,N_7126,N_7044);
and U7386 (N_7386,N_7003,N_7084);
nand U7387 (N_7387,N_7095,N_7100);
nand U7388 (N_7388,N_7175,N_7149);
nand U7389 (N_7389,N_7120,N_7133);
and U7390 (N_7390,N_7150,N_7007);
or U7391 (N_7391,N_7083,N_7119);
nor U7392 (N_7392,N_7016,N_7112);
nor U7393 (N_7393,N_7178,N_7048);
nand U7394 (N_7394,N_7055,N_7176);
nor U7395 (N_7395,N_7199,N_7005);
nor U7396 (N_7396,N_7096,N_7108);
and U7397 (N_7397,N_7035,N_7000);
and U7398 (N_7398,N_7129,N_7072);
nand U7399 (N_7399,N_7031,N_7003);
nand U7400 (N_7400,N_7250,N_7352);
nor U7401 (N_7401,N_7226,N_7340);
or U7402 (N_7402,N_7318,N_7269);
or U7403 (N_7403,N_7322,N_7304);
nor U7404 (N_7404,N_7234,N_7208);
nand U7405 (N_7405,N_7276,N_7378);
and U7406 (N_7406,N_7383,N_7293);
nor U7407 (N_7407,N_7274,N_7351);
nor U7408 (N_7408,N_7221,N_7331);
and U7409 (N_7409,N_7211,N_7207);
and U7410 (N_7410,N_7333,N_7225);
nor U7411 (N_7411,N_7348,N_7292);
nand U7412 (N_7412,N_7374,N_7245);
nand U7413 (N_7413,N_7372,N_7321);
or U7414 (N_7414,N_7213,N_7366);
nand U7415 (N_7415,N_7346,N_7230);
or U7416 (N_7416,N_7387,N_7364);
and U7417 (N_7417,N_7339,N_7291);
nor U7418 (N_7418,N_7359,N_7317);
and U7419 (N_7419,N_7324,N_7282);
nor U7420 (N_7420,N_7238,N_7257);
nor U7421 (N_7421,N_7268,N_7379);
nand U7422 (N_7422,N_7252,N_7216);
nand U7423 (N_7423,N_7261,N_7313);
xnor U7424 (N_7424,N_7254,N_7242);
nor U7425 (N_7425,N_7399,N_7338);
nand U7426 (N_7426,N_7278,N_7329);
and U7427 (N_7427,N_7305,N_7290);
nor U7428 (N_7428,N_7328,N_7354);
nand U7429 (N_7429,N_7214,N_7353);
and U7430 (N_7430,N_7259,N_7355);
or U7431 (N_7431,N_7382,N_7398);
or U7432 (N_7432,N_7319,N_7263);
and U7433 (N_7433,N_7251,N_7272);
nor U7434 (N_7434,N_7239,N_7336);
nor U7435 (N_7435,N_7286,N_7356);
nor U7436 (N_7436,N_7341,N_7285);
nor U7437 (N_7437,N_7397,N_7302);
nand U7438 (N_7438,N_7349,N_7206);
nor U7439 (N_7439,N_7395,N_7396);
nor U7440 (N_7440,N_7241,N_7246);
nor U7441 (N_7441,N_7265,N_7385);
nor U7442 (N_7442,N_7215,N_7391);
nand U7443 (N_7443,N_7345,N_7300);
nor U7444 (N_7444,N_7210,N_7334);
xnor U7445 (N_7445,N_7316,N_7231);
and U7446 (N_7446,N_7368,N_7381);
nand U7447 (N_7447,N_7307,N_7330);
nand U7448 (N_7448,N_7204,N_7343);
and U7449 (N_7449,N_7247,N_7280);
or U7450 (N_7450,N_7375,N_7394);
or U7451 (N_7451,N_7205,N_7299);
nand U7452 (N_7452,N_7362,N_7326);
xor U7453 (N_7453,N_7200,N_7350);
nor U7454 (N_7454,N_7219,N_7201);
nor U7455 (N_7455,N_7296,N_7303);
nor U7456 (N_7456,N_7209,N_7240);
nor U7457 (N_7457,N_7301,N_7284);
nor U7458 (N_7458,N_7377,N_7287);
nand U7459 (N_7459,N_7308,N_7357);
nor U7460 (N_7460,N_7369,N_7224);
nand U7461 (N_7461,N_7223,N_7376);
nand U7462 (N_7462,N_7327,N_7236);
nor U7463 (N_7463,N_7390,N_7271);
nand U7464 (N_7464,N_7371,N_7243);
and U7465 (N_7465,N_7235,N_7388);
or U7466 (N_7466,N_7222,N_7260);
nor U7467 (N_7467,N_7370,N_7203);
or U7468 (N_7468,N_7312,N_7320);
and U7469 (N_7469,N_7314,N_7323);
nor U7470 (N_7470,N_7279,N_7288);
xnor U7471 (N_7471,N_7229,N_7295);
or U7472 (N_7472,N_7347,N_7332);
or U7473 (N_7473,N_7281,N_7360);
nor U7474 (N_7474,N_7310,N_7335);
nand U7475 (N_7475,N_7337,N_7266);
nand U7476 (N_7476,N_7358,N_7311);
nand U7477 (N_7477,N_7393,N_7367);
nand U7478 (N_7478,N_7365,N_7277);
nand U7479 (N_7479,N_7306,N_7273);
and U7480 (N_7480,N_7228,N_7267);
or U7481 (N_7481,N_7217,N_7275);
or U7482 (N_7482,N_7249,N_7363);
nand U7483 (N_7483,N_7325,N_7386);
and U7484 (N_7484,N_7380,N_7218);
or U7485 (N_7485,N_7256,N_7248);
nor U7486 (N_7486,N_7297,N_7220);
and U7487 (N_7487,N_7298,N_7342);
nand U7488 (N_7488,N_7212,N_7244);
or U7489 (N_7489,N_7255,N_7233);
xnor U7490 (N_7490,N_7384,N_7202);
nand U7491 (N_7491,N_7373,N_7361);
and U7492 (N_7492,N_7270,N_7309);
nand U7493 (N_7493,N_7294,N_7227);
or U7494 (N_7494,N_7253,N_7232);
and U7495 (N_7495,N_7283,N_7237);
nand U7496 (N_7496,N_7289,N_7389);
nor U7497 (N_7497,N_7262,N_7344);
nand U7498 (N_7498,N_7258,N_7392);
nor U7499 (N_7499,N_7264,N_7315);
and U7500 (N_7500,N_7275,N_7374);
nand U7501 (N_7501,N_7340,N_7350);
and U7502 (N_7502,N_7313,N_7217);
nand U7503 (N_7503,N_7221,N_7363);
or U7504 (N_7504,N_7253,N_7269);
or U7505 (N_7505,N_7321,N_7273);
nand U7506 (N_7506,N_7230,N_7384);
or U7507 (N_7507,N_7291,N_7328);
or U7508 (N_7508,N_7328,N_7319);
nor U7509 (N_7509,N_7302,N_7323);
nand U7510 (N_7510,N_7389,N_7327);
and U7511 (N_7511,N_7392,N_7232);
nand U7512 (N_7512,N_7301,N_7270);
and U7513 (N_7513,N_7327,N_7226);
and U7514 (N_7514,N_7275,N_7303);
or U7515 (N_7515,N_7384,N_7386);
nand U7516 (N_7516,N_7300,N_7310);
or U7517 (N_7517,N_7229,N_7308);
nand U7518 (N_7518,N_7333,N_7302);
nor U7519 (N_7519,N_7371,N_7328);
or U7520 (N_7520,N_7326,N_7322);
and U7521 (N_7521,N_7382,N_7355);
nor U7522 (N_7522,N_7202,N_7380);
or U7523 (N_7523,N_7207,N_7307);
and U7524 (N_7524,N_7226,N_7224);
nor U7525 (N_7525,N_7203,N_7294);
or U7526 (N_7526,N_7221,N_7348);
nor U7527 (N_7527,N_7269,N_7282);
or U7528 (N_7528,N_7371,N_7290);
nand U7529 (N_7529,N_7357,N_7225);
nor U7530 (N_7530,N_7381,N_7283);
nand U7531 (N_7531,N_7230,N_7307);
and U7532 (N_7532,N_7276,N_7292);
and U7533 (N_7533,N_7306,N_7201);
nand U7534 (N_7534,N_7387,N_7235);
nand U7535 (N_7535,N_7248,N_7307);
nor U7536 (N_7536,N_7235,N_7210);
nand U7537 (N_7537,N_7291,N_7318);
xnor U7538 (N_7538,N_7223,N_7252);
nor U7539 (N_7539,N_7353,N_7303);
nor U7540 (N_7540,N_7356,N_7335);
and U7541 (N_7541,N_7369,N_7326);
nand U7542 (N_7542,N_7221,N_7283);
nand U7543 (N_7543,N_7293,N_7246);
and U7544 (N_7544,N_7367,N_7294);
nand U7545 (N_7545,N_7210,N_7304);
and U7546 (N_7546,N_7229,N_7235);
nor U7547 (N_7547,N_7376,N_7298);
nand U7548 (N_7548,N_7393,N_7255);
nor U7549 (N_7549,N_7300,N_7289);
and U7550 (N_7550,N_7342,N_7386);
or U7551 (N_7551,N_7268,N_7280);
or U7552 (N_7552,N_7263,N_7244);
or U7553 (N_7553,N_7394,N_7374);
or U7554 (N_7554,N_7397,N_7392);
nor U7555 (N_7555,N_7333,N_7369);
nor U7556 (N_7556,N_7389,N_7377);
nand U7557 (N_7557,N_7394,N_7398);
nand U7558 (N_7558,N_7313,N_7206);
or U7559 (N_7559,N_7374,N_7210);
nor U7560 (N_7560,N_7286,N_7321);
or U7561 (N_7561,N_7216,N_7239);
or U7562 (N_7562,N_7218,N_7262);
nor U7563 (N_7563,N_7201,N_7276);
nand U7564 (N_7564,N_7260,N_7281);
or U7565 (N_7565,N_7336,N_7389);
nand U7566 (N_7566,N_7334,N_7206);
nand U7567 (N_7567,N_7354,N_7351);
nor U7568 (N_7568,N_7295,N_7342);
xnor U7569 (N_7569,N_7266,N_7395);
and U7570 (N_7570,N_7398,N_7331);
nand U7571 (N_7571,N_7215,N_7265);
or U7572 (N_7572,N_7235,N_7251);
and U7573 (N_7573,N_7323,N_7344);
nor U7574 (N_7574,N_7376,N_7293);
nand U7575 (N_7575,N_7326,N_7302);
or U7576 (N_7576,N_7358,N_7234);
or U7577 (N_7577,N_7225,N_7286);
and U7578 (N_7578,N_7241,N_7359);
nand U7579 (N_7579,N_7247,N_7365);
nor U7580 (N_7580,N_7233,N_7376);
and U7581 (N_7581,N_7382,N_7208);
nand U7582 (N_7582,N_7223,N_7390);
nand U7583 (N_7583,N_7346,N_7374);
and U7584 (N_7584,N_7277,N_7366);
nor U7585 (N_7585,N_7238,N_7355);
and U7586 (N_7586,N_7208,N_7200);
nand U7587 (N_7587,N_7338,N_7273);
nand U7588 (N_7588,N_7346,N_7375);
and U7589 (N_7589,N_7350,N_7306);
nand U7590 (N_7590,N_7361,N_7360);
nor U7591 (N_7591,N_7398,N_7320);
nand U7592 (N_7592,N_7270,N_7273);
and U7593 (N_7593,N_7203,N_7212);
nor U7594 (N_7594,N_7335,N_7355);
nand U7595 (N_7595,N_7366,N_7228);
nor U7596 (N_7596,N_7338,N_7381);
nor U7597 (N_7597,N_7357,N_7252);
nor U7598 (N_7598,N_7212,N_7356);
and U7599 (N_7599,N_7381,N_7359);
nand U7600 (N_7600,N_7455,N_7552);
nor U7601 (N_7601,N_7589,N_7467);
nor U7602 (N_7602,N_7429,N_7558);
and U7603 (N_7603,N_7418,N_7427);
nor U7604 (N_7604,N_7464,N_7542);
and U7605 (N_7605,N_7413,N_7447);
nor U7606 (N_7606,N_7557,N_7595);
nor U7607 (N_7607,N_7507,N_7593);
xnor U7608 (N_7608,N_7579,N_7435);
nor U7609 (N_7609,N_7517,N_7416);
or U7610 (N_7610,N_7582,N_7443);
nor U7611 (N_7611,N_7434,N_7521);
and U7612 (N_7612,N_7597,N_7537);
and U7613 (N_7613,N_7560,N_7489);
or U7614 (N_7614,N_7472,N_7534);
nand U7615 (N_7615,N_7463,N_7504);
or U7616 (N_7616,N_7513,N_7495);
or U7617 (N_7617,N_7478,N_7514);
nand U7618 (N_7618,N_7439,N_7473);
or U7619 (N_7619,N_7576,N_7549);
or U7620 (N_7620,N_7519,N_7506);
and U7621 (N_7621,N_7437,N_7591);
or U7622 (N_7622,N_7441,N_7406);
nor U7623 (N_7623,N_7585,N_7566);
and U7624 (N_7624,N_7469,N_7491);
and U7625 (N_7625,N_7553,N_7551);
nor U7626 (N_7626,N_7512,N_7461);
nand U7627 (N_7627,N_7402,N_7404);
nand U7628 (N_7628,N_7428,N_7545);
or U7629 (N_7629,N_7479,N_7480);
nand U7630 (N_7630,N_7531,N_7527);
or U7631 (N_7631,N_7408,N_7544);
and U7632 (N_7632,N_7475,N_7538);
nand U7633 (N_7633,N_7430,N_7539);
and U7634 (N_7634,N_7452,N_7509);
or U7635 (N_7635,N_7448,N_7486);
or U7636 (N_7636,N_7508,N_7497);
or U7637 (N_7637,N_7500,N_7492);
nor U7638 (N_7638,N_7401,N_7586);
nand U7639 (N_7639,N_7420,N_7599);
and U7640 (N_7640,N_7575,N_7554);
nor U7641 (N_7641,N_7498,N_7528);
nand U7642 (N_7642,N_7564,N_7476);
nor U7643 (N_7643,N_7481,N_7563);
nand U7644 (N_7644,N_7490,N_7598);
or U7645 (N_7645,N_7451,N_7574);
and U7646 (N_7646,N_7547,N_7438);
nor U7647 (N_7647,N_7596,N_7407);
and U7648 (N_7648,N_7535,N_7590);
nor U7649 (N_7649,N_7410,N_7445);
xnor U7650 (N_7650,N_7525,N_7477);
or U7651 (N_7651,N_7580,N_7433);
nand U7652 (N_7652,N_7412,N_7515);
nor U7653 (N_7653,N_7436,N_7567);
nand U7654 (N_7654,N_7584,N_7470);
nor U7655 (N_7655,N_7449,N_7588);
and U7656 (N_7656,N_7543,N_7529);
and U7657 (N_7657,N_7530,N_7440);
or U7658 (N_7658,N_7561,N_7468);
and U7659 (N_7659,N_7570,N_7487);
nor U7660 (N_7660,N_7442,N_7405);
and U7661 (N_7661,N_7496,N_7562);
nand U7662 (N_7662,N_7499,N_7431);
and U7663 (N_7663,N_7555,N_7450);
nand U7664 (N_7664,N_7524,N_7493);
nor U7665 (N_7665,N_7532,N_7518);
nand U7666 (N_7666,N_7565,N_7400);
nor U7667 (N_7667,N_7494,N_7510);
nor U7668 (N_7668,N_7548,N_7594);
and U7669 (N_7669,N_7505,N_7424);
and U7670 (N_7670,N_7403,N_7484);
or U7671 (N_7671,N_7466,N_7503);
and U7672 (N_7672,N_7546,N_7411);
nor U7673 (N_7673,N_7453,N_7458);
or U7674 (N_7674,N_7474,N_7459);
or U7675 (N_7675,N_7550,N_7516);
xnor U7676 (N_7676,N_7419,N_7556);
or U7677 (N_7677,N_7421,N_7415);
and U7678 (N_7678,N_7581,N_7572);
nand U7679 (N_7679,N_7457,N_7577);
and U7680 (N_7680,N_7541,N_7409);
and U7681 (N_7681,N_7569,N_7444);
nor U7682 (N_7682,N_7511,N_7501);
and U7683 (N_7683,N_7533,N_7426);
nor U7684 (N_7684,N_7462,N_7522);
nor U7685 (N_7685,N_7460,N_7425);
or U7686 (N_7686,N_7414,N_7483);
nor U7687 (N_7687,N_7578,N_7446);
nand U7688 (N_7688,N_7540,N_7571);
nor U7689 (N_7689,N_7417,N_7526);
or U7690 (N_7690,N_7485,N_7423);
nor U7691 (N_7691,N_7502,N_7456);
xor U7692 (N_7692,N_7583,N_7471);
nand U7693 (N_7693,N_7432,N_7454);
or U7694 (N_7694,N_7536,N_7465);
and U7695 (N_7695,N_7482,N_7587);
nor U7696 (N_7696,N_7592,N_7559);
nand U7697 (N_7697,N_7422,N_7568);
nor U7698 (N_7698,N_7573,N_7520);
nand U7699 (N_7699,N_7523,N_7488);
nor U7700 (N_7700,N_7503,N_7439);
and U7701 (N_7701,N_7500,N_7490);
and U7702 (N_7702,N_7459,N_7457);
nand U7703 (N_7703,N_7400,N_7566);
or U7704 (N_7704,N_7519,N_7583);
and U7705 (N_7705,N_7493,N_7507);
and U7706 (N_7706,N_7514,N_7590);
and U7707 (N_7707,N_7523,N_7576);
nor U7708 (N_7708,N_7410,N_7408);
nand U7709 (N_7709,N_7514,N_7444);
nor U7710 (N_7710,N_7515,N_7484);
and U7711 (N_7711,N_7464,N_7492);
nor U7712 (N_7712,N_7552,N_7471);
or U7713 (N_7713,N_7559,N_7583);
nand U7714 (N_7714,N_7476,N_7429);
and U7715 (N_7715,N_7458,N_7508);
or U7716 (N_7716,N_7583,N_7533);
xnor U7717 (N_7717,N_7535,N_7547);
nor U7718 (N_7718,N_7471,N_7527);
and U7719 (N_7719,N_7469,N_7506);
or U7720 (N_7720,N_7580,N_7500);
or U7721 (N_7721,N_7502,N_7590);
and U7722 (N_7722,N_7520,N_7514);
and U7723 (N_7723,N_7479,N_7483);
or U7724 (N_7724,N_7422,N_7513);
nand U7725 (N_7725,N_7541,N_7462);
nand U7726 (N_7726,N_7497,N_7421);
or U7727 (N_7727,N_7506,N_7537);
or U7728 (N_7728,N_7548,N_7501);
nor U7729 (N_7729,N_7455,N_7526);
nand U7730 (N_7730,N_7513,N_7553);
nand U7731 (N_7731,N_7412,N_7598);
or U7732 (N_7732,N_7468,N_7570);
nand U7733 (N_7733,N_7420,N_7524);
or U7734 (N_7734,N_7409,N_7457);
nor U7735 (N_7735,N_7578,N_7420);
nand U7736 (N_7736,N_7516,N_7588);
nor U7737 (N_7737,N_7478,N_7470);
nor U7738 (N_7738,N_7436,N_7480);
xor U7739 (N_7739,N_7404,N_7533);
nor U7740 (N_7740,N_7434,N_7532);
nand U7741 (N_7741,N_7588,N_7478);
and U7742 (N_7742,N_7572,N_7528);
nand U7743 (N_7743,N_7488,N_7540);
nand U7744 (N_7744,N_7502,N_7405);
xor U7745 (N_7745,N_7579,N_7574);
or U7746 (N_7746,N_7430,N_7530);
and U7747 (N_7747,N_7541,N_7533);
nor U7748 (N_7748,N_7476,N_7508);
and U7749 (N_7749,N_7431,N_7506);
nor U7750 (N_7750,N_7404,N_7414);
nand U7751 (N_7751,N_7493,N_7573);
and U7752 (N_7752,N_7503,N_7501);
and U7753 (N_7753,N_7594,N_7589);
and U7754 (N_7754,N_7530,N_7480);
nor U7755 (N_7755,N_7524,N_7433);
and U7756 (N_7756,N_7598,N_7447);
or U7757 (N_7757,N_7489,N_7472);
and U7758 (N_7758,N_7555,N_7522);
nand U7759 (N_7759,N_7449,N_7538);
nor U7760 (N_7760,N_7497,N_7479);
and U7761 (N_7761,N_7548,N_7569);
nor U7762 (N_7762,N_7486,N_7540);
and U7763 (N_7763,N_7494,N_7523);
and U7764 (N_7764,N_7471,N_7572);
nor U7765 (N_7765,N_7518,N_7430);
nand U7766 (N_7766,N_7503,N_7437);
nor U7767 (N_7767,N_7450,N_7526);
or U7768 (N_7768,N_7502,N_7414);
nor U7769 (N_7769,N_7452,N_7547);
nand U7770 (N_7770,N_7517,N_7417);
and U7771 (N_7771,N_7579,N_7403);
nand U7772 (N_7772,N_7584,N_7440);
and U7773 (N_7773,N_7444,N_7582);
or U7774 (N_7774,N_7532,N_7438);
nor U7775 (N_7775,N_7548,N_7421);
and U7776 (N_7776,N_7458,N_7511);
or U7777 (N_7777,N_7557,N_7428);
nand U7778 (N_7778,N_7480,N_7591);
nand U7779 (N_7779,N_7572,N_7416);
nand U7780 (N_7780,N_7569,N_7506);
and U7781 (N_7781,N_7481,N_7527);
or U7782 (N_7782,N_7421,N_7410);
nand U7783 (N_7783,N_7493,N_7548);
and U7784 (N_7784,N_7482,N_7473);
nor U7785 (N_7785,N_7487,N_7513);
and U7786 (N_7786,N_7514,N_7555);
xor U7787 (N_7787,N_7522,N_7482);
and U7788 (N_7788,N_7446,N_7424);
nor U7789 (N_7789,N_7559,N_7477);
nand U7790 (N_7790,N_7515,N_7493);
and U7791 (N_7791,N_7452,N_7555);
nand U7792 (N_7792,N_7535,N_7520);
nor U7793 (N_7793,N_7465,N_7453);
nand U7794 (N_7794,N_7473,N_7450);
nand U7795 (N_7795,N_7540,N_7576);
or U7796 (N_7796,N_7460,N_7578);
nor U7797 (N_7797,N_7546,N_7481);
nand U7798 (N_7798,N_7525,N_7513);
and U7799 (N_7799,N_7523,N_7585);
xnor U7800 (N_7800,N_7630,N_7747);
nand U7801 (N_7801,N_7681,N_7692);
and U7802 (N_7802,N_7695,N_7743);
or U7803 (N_7803,N_7729,N_7646);
nand U7804 (N_7804,N_7788,N_7619);
nor U7805 (N_7805,N_7770,N_7777);
nand U7806 (N_7806,N_7702,N_7795);
xnor U7807 (N_7807,N_7727,N_7786);
nand U7808 (N_7808,N_7633,N_7600);
nor U7809 (N_7809,N_7704,N_7769);
and U7810 (N_7810,N_7768,N_7782);
nor U7811 (N_7811,N_7698,N_7725);
nand U7812 (N_7812,N_7601,N_7640);
nand U7813 (N_7813,N_7605,N_7669);
and U7814 (N_7814,N_7772,N_7613);
nor U7815 (N_7815,N_7703,N_7617);
nand U7816 (N_7816,N_7721,N_7738);
nor U7817 (N_7817,N_7637,N_7737);
nand U7818 (N_7818,N_7716,N_7649);
or U7819 (N_7819,N_7664,N_7739);
nor U7820 (N_7820,N_7734,N_7783);
nor U7821 (N_7821,N_7672,N_7732);
nor U7822 (N_7822,N_7756,N_7791);
or U7823 (N_7823,N_7674,N_7781);
or U7824 (N_7824,N_7684,N_7628);
or U7825 (N_7825,N_7709,N_7645);
or U7826 (N_7826,N_7762,N_7616);
nand U7827 (N_7827,N_7723,N_7618);
and U7828 (N_7828,N_7657,N_7751);
or U7829 (N_7829,N_7602,N_7708);
nor U7830 (N_7830,N_7771,N_7647);
or U7831 (N_7831,N_7745,N_7722);
and U7832 (N_7832,N_7644,N_7690);
xnor U7833 (N_7833,N_7730,N_7615);
nand U7834 (N_7834,N_7790,N_7687);
and U7835 (N_7835,N_7779,N_7686);
nand U7836 (N_7836,N_7660,N_7655);
or U7837 (N_7837,N_7662,N_7607);
or U7838 (N_7838,N_7606,N_7648);
and U7839 (N_7839,N_7668,N_7694);
nor U7840 (N_7840,N_7789,N_7629);
and U7841 (N_7841,N_7611,N_7714);
nand U7842 (N_7842,N_7742,N_7774);
nor U7843 (N_7843,N_7604,N_7706);
nor U7844 (N_7844,N_7766,N_7667);
nor U7845 (N_7845,N_7627,N_7603);
nor U7846 (N_7846,N_7659,N_7636);
nand U7847 (N_7847,N_7691,N_7713);
nand U7848 (N_7848,N_7642,N_7775);
and U7849 (N_7849,N_7639,N_7767);
and U7850 (N_7850,N_7675,N_7683);
and U7851 (N_7851,N_7631,N_7700);
nand U7852 (N_7852,N_7621,N_7753);
nor U7853 (N_7853,N_7757,N_7712);
nor U7854 (N_7854,N_7758,N_7707);
and U7855 (N_7855,N_7792,N_7744);
nand U7856 (N_7856,N_7614,N_7728);
nand U7857 (N_7857,N_7678,N_7796);
nand U7858 (N_7858,N_7719,N_7711);
and U7859 (N_7859,N_7658,N_7733);
and U7860 (N_7860,N_7760,N_7787);
and U7861 (N_7861,N_7653,N_7680);
nand U7862 (N_7862,N_7759,N_7701);
and U7863 (N_7863,N_7717,N_7705);
and U7864 (N_7864,N_7625,N_7697);
nand U7865 (N_7865,N_7785,N_7622);
and U7866 (N_7866,N_7688,N_7670);
nor U7867 (N_7867,N_7780,N_7656);
or U7868 (N_7868,N_7752,N_7740);
nor U7869 (N_7869,N_7623,N_7754);
nand U7870 (N_7870,N_7735,N_7731);
or U7871 (N_7871,N_7654,N_7726);
or U7872 (N_7872,N_7673,N_7610);
nor U7873 (N_7873,N_7661,N_7746);
or U7874 (N_7874,N_7778,N_7685);
and U7875 (N_7875,N_7763,N_7671);
or U7876 (N_7876,N_7741,N_7635);
nand U7877 (N_7877,N_7666,N_7609);
or U7878 (N_7878,N_7651,N_7650);
or U7879 (N_7879,N_7715,N_7624);
or U7880 (N_7880,N_7677,N_7710);
nor U7881 (N_7881,N_7798,N_7652);
or U7882 (N_7882,N_7718,N_7699);
and U7883 (N_7883,N_7679,N_7696);
or U7884 (N_7884,N_7773,N_7793);
nand U7885 (N_7885,N_7799,N_7749);
or U7886 (N_7886,N_7638,N_7620);
nand U7887 (N_7887,N_7776,N_7750);
nor U7888 (N_7888,N_7663,N_7797);
or U7889 (N_7889,N_7626,N_7748);
nor U7890 (N_7890,N_7765,N_7612);
nor U7891 (N_7891,N_7755,N_7724);
nor U7892 (N_7892,N_7761,N_7764);
nand U7893 (N_7893,N_7665,N_7676);
or U7894 (N_7894,N_7736,N_7794);
or U7895 (N_7895,N_7720,N_7682);
xor U7896 (N_7896,N_7643,N_7634);
and U7897 (N_7897,N_7608,N_7693);
or U7898 (N_7898,N_7689,N_7632);
nor U7899 (N_7899,N_7641,N_7784);
or U7900 (N_7900,N_7636,N_7724);
nor U7901 (N_7901,N_7671,N_7681);
or U7902 (N_7902,N_7679,N_7722);
or U7903 (N_7903,N_7782,N_7652);
or U7904 (N_7904,N_7716,N_7690);
nor U7905 (N_7905,N_7690,N_7759);
nand U7906 (N_7906,N_7705,N_7633);
and U7907 (N_7907,N_7603,N_7680);
nand U7908 (N_7908,N_7676,N_7624);
and U7909 (N_7909,N_7701,N_7648);
or U7910 (N_7910,N_7756,N_7646);
or U7911 (N_7911,N_7668,N_7617);
nor U7912 (N_7912,N_7696,N_7636);
or U7913 (N_7913,N_7732,N_7791);
or U7914 (N_7914,N_7667,N_7683);
nand U7915 (N_7915,N_7728,N_7703);
nand U7916 (N_7916,N_7795,N_7723);
or U7917 (N_7917,N_7669,N_7675);
and U7918 (N_7918,N_7604,N_7697);
and U7919 (N_7919,N_7783,N_7777);
and U7920 (N_7920,N_7700,N_7694);
or U7921 (N_7921,N_7657,N_7639);
and U7922 (N_7922,N_7710,N_7766);
nor U7923 (N_7923,N_7799,N_7600);
and U7924 (N_7924,N_7606,N_7795);
or U7925 (N_7925,N_7755,N_7763);
or U7926 (N_7926,N_7724,N_7792);
and U7927 (N_7927,N_7670,N_7600);
or U7928 (N_7928,N_7666,N_7689);
or U7929 (N_7929,N_7623,N_7782);
nand U7930 (N_7930,N_7664,N_7676);
xor U7931 (N_7931,N_7731,N_7775);
or U7932 (N_7932,N_7705,N_7712);
and U7933 (N_7933,N_7699,N_7710);
nand U7934 (N_7934,N_7652,N_7611);
nand U7935 (N_7935,N_7745,N_7796);
nor U7936 (N_7936,N_7777,N_7743);
or U7937 (N_7937,N_7796,N_7765);
nand U7938 (N_7938,N_7741,N_7647);
and U7939 (N_7939,N_7754,N_7713);
nand U7940 (N_7940,N_7742,N_7707);
nor U7941 (N_7941,N_7733,N_7719);
and U7942 (N_7942,N_7752,N_7638);
and U7943 (N_7943,N_7675,N_7755);
and U7944 (N_7944,N_7763,N_7613);
nand U7945 (N_7945,N_7631,N_7741);
or U7946 (N_7946,N_7742,N_7645);
nand U7947 (N_7947,N_7799,N_7724);
or U7948 (N_7948,N_7746,N_7786);
and U7949 (N_7949,N_7656,N_7662);
nand U7950 (N_7950,N_7741,N_7698);
nor U7951 (N_7951,N_7657,N_7779);
or U7952 (N_7952,N_7736,N_7727);
or U7953 (N_7953,N_7753,N_7604);
nand U7954 (N_7954,N_7700,N_7729);
or U7955 (N_7955,N_7632,N_7684);
nor U7956 (N_7956,N_7694,N_7636);
nand U7957 (N_7957,N_7699,N_7738);
nand U7958 (N_7958,N_7631,N_7683);
and U7959 (N_7959,N_7613,N_7659);
nand U7960 (N_7960,N_7687,N_7714);
nor U7961 (N_7961,N_7621,N_7716);
nand U7962 (N_7962,N_7695,N_7712);
nor U7963 (N_7963,N_7647,N_7621);
nand U7964 (N_7964,N_7688,N_7623);
xnor U7965 (N_7965,N_7793,N_7664);
nand U7966 (N_7966,N_7654,N_7671);
nor U7967 (N_7967,N_7632,N_7748);
nor U7968 (N_7968,N_7699,N_7752);
or U7969 (N_7969,N_7793,N_7625);
xnor U7970 (N_7970,N_7758,N_7651);
and U7971 (N_7971,N_7747,N_7757);
nand U7972 (N_7972,N_7776,N_7689);
nand U7973 (N_7973,N_7694,N_7670);
nor U7974 (N_7974,N_7614,N_7699);
and U7975 (N_7975,N_7714,N_7686);
and U7976 (N_7976,N_7679,N_7779);
or U7977 (N_7977,N_7612,N_7666);
nand U7978 (N_7978,N_7663,N_7634);
nor U7979 (N_7979,N_7630,N_7681);
nand U7980 (N_7980,N_7672,N_7799);
xnor U7981 (N_7981,N_7776,N_7664);
and U7982 (N_7982,N_7616,N_7618);
or U7983 (N_7983,N_7761,N_7688);
nand U7984 (N_7984,N_7776,N_7640);
xor U7985 (N_7985,N_7699,N_7788);
and U7986 (N_7986,N_7606,N_7761);
or U7987 (N_7987,N_7604,N_7689);
nor U7988 (N_7988,N_7601,N_7766);
nand U7989 (N_7989,N_7608,N_7758);
nor U7990 (N_7990,N_7686,N_7718);
and U7991 (N_7991,N_7777,N_7784);
and U7992 (N_7992,N_7796,N_7642);
xnor U7993 (N_7993,N_7732,N_7739);
or U7994 (N_7994,N_7701,N_7712);
xnor U7995 (N_7995,N_7630,N_7776);
nor U7996 (N_7996,N_7625,N_7672);
nand U7997 (N_7997,N_7747,N_7792);
or U7998 (N_7998,N_7708,N_7749);
xor U7999 (N_7999,N_7756,N_7792);
or U8000 (N_8000,N_7836,N_7846);
nor U8001 (N_8001,N_7940,N_7867);
nor U8002 (N_8002,N_7890,N_7932);
nand U8003 (N_8003,N_7903,N_7803);
nor U8004 (N_8004,N_7997,N_7871);
nor U8005 (N_8005,N_7918,N_7881);
nand U8006 (N_8006,N_7964,N_7902);
and U8007 (N_8007,N_7832,N_7883);
and U8008 (N_8008,N_7808,N_7886);
or U8009 (N_8009,N_7819,N_7991);
nor U8010 (N_8010,N_7875,N_7974);
nand U8011 (N_8011,N_7901,N_7952);
nand U8012 (N_8012,N_7801,N_7946);
or U8013 (N_8013,N_7870,N_7844);
or U8014 (N_8014,N_7920,N_7865);
nor U8015 (N_8015,N_7949,N_7843);
or U8016 (N_8016,N_7899,N_7965);
or U8017 (N_8017,N_7927,N_7840);
nor U8018 (N_8018,N_7897,N_7975);
xnor U8019 (N_8019,N_7914,N_7830);
and U8020 (N_8020,N_7906,N_7988);
nand U8021 (N_8021,N_7944,N_7880);
and U8022 (N_8022,N_7817,N_7851);
or U8023 (N_8023,N_7845,N_7999);
and U8024 (N_8024,N_7834,N_7885);
nor U8025 (N_8025,N_7933,N_7820);
nand U8026 (N_8026,N_7976,N_7812);
or U8027 (N_8027,N_7935,N_7937);
nor U8028 (N_8028,N_7805,N_7866);
and U8029 (N_8029,N_7986,N_7982);
nor U8030 (N_8030,N_7900,N_7876);
and U8031 (N_8031,N_7895,N_7929);
and U8032 (N_8032,N_7831,N_7981);
nor U8033 (N_8033,N_7888,N_7841);
nor U8034 (N_8034,N_7939,N_7936);
xnor U8035 (N_8035,N_7892,N_7908);
nor U8036 (N_8036,N_7913,N_7894);
or U8037 (N_8037,N_7823,N_7879);
nor U8038 (N_8038,N_7800,N_7924);
and U8039 (N_8039,N_7859,N_7923);
nand U8040 (N_8040,N_7847,N_7860);
nand U8041 (N_8041,N_7868,N_7984);
nor U8042 (N_8042,N_7978,N_7833);
and U8043 (N_8043,N_7921,N_7874);
nand U8044 (N_8044,N_7912,N_7824);
nor U8045 (N_8045,N_7905,N_7850);
and U8046 (N_8046,N_7989,N_7941);
nand U8047 (N_8047,N_7804,N_7864);
nor U8048 (N_8048,N_7926,N_7909);
nor U8049 (N_8049,N_7950,N_7838);
nor U8050 (N_8050,N_7996,N_7891);
and U8051 (N_8051,N_7943,N_7893);
nor U8052 (N_8052,N_7821,N_7960);
or U8053 (N_8053,N_7861,N_7959);
nor U8054 (N_8054,N_7977,N_7917);
nand U8055 (N_8055,N_7907,N_7818);
nor U8056 (N_8056,N_7953,N_7807);
and U8057 (N_8057,N_7969,N_7995);
nor U8058 (N_8058,N_7904,N_7948);
xnor U8059 (N_8059,N_7919,N_7966);
nor U8060 (N_8060,N_7922,N_7916);
or U8061 (N_8061,N_7884,N_7992);
and U8062 (N_8062,N_7947,N_7987);
nor U8063 (N_8063,N_7958,N_7813);
or U8064 (N_8064,N_7872,N_7815);
or U8065 (N_8065,N_7961,N_7882);
and U8066 (N_8066,N_7855,N_7915);
and U8067 (N_8067,N_7837,N_7814);
and U8068 (N_8068,N_7896,N_7955);
and U8069 (N_8069,N_7887,N_7990);
and U8070 (N_8070,N_7835,N_7972);
nor U8071 (N_8071,N_7852,N_7839);
and U8072 (N_8072,N_7848,N_7842);
or U8073 (N_8073,N_7934,N_7970);
or U8074 (N_8074,N_7827,N_7862);
and U8075 (N_8075,N_7951,N_7994);
and U8076 (N_8076,N_7931,N_7971);
or U8077 (N_8077,N_7828,N_7911);
nand U8078 (N_8078,N_7829,N_7826);
nand U8079 (N_8079,N_7993,N_7889);
nand U8080 (N_8080,N_7973,N_7816);
nand U8081 (N_8081,N_7910,N_7873);
nand U8082 (N_8082,N_7998,N_7811);
nor U8083 (N_8083,N_7858,N_7957);
nand U8084 (N_8084,N_7877,N_7928);
nor U8085 (N_8085,N_7853,N_7930);
nand U8086 (N_8086,N_7898,N_7956);
and U8087 (N_8087,N_7863,N_7942);
nor U8088 (N_8088,N_7856,N_7962);
and U8089 (N_8089,N_7806,N_7822);
nand U8090 (N_8090,N_7802,N_7825);
or U8091 (N_8091,N_7979,N_7849);
or U8092 (N_8092,N_7945,N_7854);
nor U8093 (N_8093,N_7857,N_7954);
or U8094 (N_8094,N_7938,N_7963);
nor U8095 (N_8095,N_7810,N_7878);
nand U8096 (N_8096,N_7809,N_7869);
and U8097 (N_8097,N_7967,N_7983);
or U8098 (N_8098,N_7968,N_7925);
and U8099 (N_8099,N_7980,N_7985);
nor U8100 (N_8100,N_7821,N_7976);
nor U8101 (N_8101,N_7876,N_7970);
and U8102 (N_8102,N_7873,N_7916);
nand U8103 (N_8103,N_7996,N_7858);
or U8104 (N_8104,N_7878,N_7961);
nor U8105 (N_8105,N_7832,N_7968);
nor U8106 (N_8106,N_7821,N_7887);
nand U8107 (N_8107,N_7830,N_7877);
or U8108 (N_8108,N_7956,N_7873);
nor U8109 (N_8109,N_7891,N_7892);
nand U8110 (N_8110,N_7945,N_7822);
nand U8111 (N_8111,N_7933,N_7908);
and U8112 (N_8112,N_7908,N_7810);
nand U8113 (N_8113,N_7892,N_7930);
and U8114 (N_8114,N_7986,N_7818);
or U8115 (N_8115,N_7823,N_7996);
or U8116 (N_8116,N_7977,N_7814);
or U8117 (N_8117,N_7978,N_7958);
nor U8118 (N_8118,N_7937,N_7908);
xnor U8119 (N_8119,N_7865,N_7911);
and U8120 (N_8120,N_7924,N_7997);
nor U8121 (N_8121,N_7836,N_7894);
or U8122 (N_8122,N_7974,N_7941);
nor U8123 (N_8123,N_7989,N_7806);
nor U8124 (N_8124,N_7842,N_7864);
and U8125 (N_8125,N_7806,N_7849);
nand U8126 (N_8126,N_7932,N_7892);
or U8127 (N_8127,N_7984,N_7907);
and U8128 (N_8128,N_7997,N_7881);
nor U8129 (N_8129,N_7982,N_7969);
nor U8130 (N_8130,N_7877,N_7903);
nor U8131 (N_8131,N_7964,N_7945);
nor U8132 (N_8132,N_7965,N_7902);
nand U8133 (N_8133,N_7896,N_7993);
nand U8134 (N_8134,N_7803,N_7900);
nand U8135 (N_8135,N_7879,N_7878);
nor U8136 (N_8136,N_7807,N_7964);
nor U8137 (N_8137,N_7942,N_7844);
nor U8138 (N_8138,N_7806,N_7886);
or U8139 (N_8139,N_7849,N_7818);
nor U8140 (N_8140,N_7853,N_7946);
or U8141 (N_8141,N_7935,N_7952);
nor U8142 (N_8142,N_7877,N_7810);
nand U8143 (N_8143,N_7814,N_7840);
nand U8144 (N_8144,N_7832,N_7834);
or U8145 (N_8145,N_7843,N_7982);
nor U8146 (N_8146,N_7949,N_7861);
and U8147 (N_8147,N_7956,N_7886);
nand U8148 (N_8148,N_7894,N_7953);
and U8149 (N_8149,N_7814,N_7974);
and U8150 (N_8150,N_7999,N_7883);
nor U8151 (N_8151,N_7937,N_7978);
nor U8152 (N_8152,N_7815,N_7877);
nand U8153 (N_8153,N_7815,N_7974);
and U8154 (N_8154,N_7892,N_7952);
and U8155 (N_8155,N_7914,N_7861);
or U8156 (N_8156,N_7957,N_7834);
and U8157 (N_8157,N_7944,N_7803);
and U8158 (N_8158,N_7946,N_7978);
and U8159 (N_8159,N_7834,N_7846);
nor U8160 (N_8160,N_7912,N_7862);
and U8161 (N_8161,N_7835,N_7820);
and U8162 (N_8162,N_7935,N_7894);
nor U8163 (N_8163,N_7888,N_7933);
nor U8164 (N_8164,N_7925,N_7964);
or U8165 (N_8165,N_7863,N_7867);
nor U8166 (N_8166,N_7994,N_7959);
nand U8167 (N_8167,N_7972,N_7814);
and U8168 (N_8168,N_7855,N_7889);
nor U8169 (N_8169,N_7908,N_7903);
nor U8170 (N_8170,N_7895,N_7867);
and U8171 (N_8171,N_7802,N_7936);
or U8172 (N_8172,N_7869,N_7862);
or U8173 (N_8173,N_7850,N_7846);
nand U8174 (N_8174,N_7991,N_7813);
and U8175 (N_8175,N_7858,N_7900);
and U8176 (N_8176,N_7820,N_7918);
nand U8177 (N_8177,N_7988,N_7925);
or U8178 (N_8178,N_7955,N_7906);
and U8179 (N_8179,N_7803,N_7836);
or U8180 (N_8180,N_7982,N_7803);
or U8181 (N_8181,N_7952,N_7854);
nor U8182 (N_8182,N_7812,N_7809);
or U8183 (N_8183,N_7804,N_7886);
nand U8184 (N_8184,N_7906,N_7804);
and U8185 (N_8185,N_7875,N_7837);
nor U8186 (N_8186,N_7804,N_7968);
and U8187 (N_8187,N_7925,N_7947);
or U8188 (N_8188,N_7840,N_7836);
nor U8189 (N_8189,N_7838,N_7850);
nor U8190 (N_8190,N_7966,N_7872);
nor U8191 (N_8191,N_7883,N_7877);
or U8192 (N_8192,N_7987,N_7991);
nor U8193 (N_8193,N_7818,N_7952);
or U8194 (N_8194,N_7868,N_7841);
nand U8195 (N_8195,N_7908,N_7825);
and U8196 (N_8196,N_7910,N_7823);
and U8197 (N_8197,N_7943,N_7956);
nand U8198 (N_8198,N_7880,N_7887);
or U8199 (N_8199,N_7832,N_7850);
and U8200 (N_8200,N_8097,N_8195);
and U8201 (N_8201,N_8148,N_8176);
and U8202 (N_8202,N_8099,N_8062);
or U8203 (N_8203,N_8004,N_8017);
nor U8204 (N_8204,N_8057,N_8187);
nor U8205 (N_8205,N_8128,N_8151);
nor U8206 (N_8206,N_8166,N_8173);
xor U8207 (N_8207,N_8041,N_8095);
and U8208 (N_8208,N_8016,N_8160);
nor U8209 (N_8209,N_8014,N_8009);
or U8210 (N_8210,N_8040,N_8067);
nand U8211 (N_8211,N_8010,N_8070);
or U8212 (N_8212,N_8131,N_8044);
and U8213 (N_8213,N_8172,N_8027);
or U8214 (N_8214,N_8159,N_8129);
nor U8215 (N_8215,N_8190,N_8028);
and U8216 (N_8216,N_8049,N_8154);
and U8217 (N_8217,N_8082,N_8071);
and U8218 (N_8218,N_8081,N_8119);
and U8219 (N_8219,N_8092,N_8168);
nand U8220 (N_8220,N_8075,N_8036);
nand U8221 (N_8221,N_8038,N_8026);
nand U8222 (N_8222,N_8105,N_8110);
nor U8223 (N_8223,N_8145,N_8140);
nor U8224 (N_8224,N_8127,N_8073);
and U8225 (N_8225,N_8037,N_8183);
and U8226 (N_8226,N_8132,N_8029);
or U8227 (N_8227,N_8064,N_8039);
nand U8228 (N_8228,N_8072,N_8002);
nor U8229 (N_8229,N_8135,N_8153);
nor U8230 (N_8230,N_8114,N_8011);
or U8231 (N_8231,N_8125,N_8006);
or U8232 (N_8232,N_8188,N_8141);
and U8233 (N_8233,N_8089,N_8033);
and U8234 (N_8234,N_8056,N_8170);
or U8235 (N_8235,N_8178,N_8186);
and U8236 (N_8236,N_8093,N_8196);
and U8237 (N_8237,N_8008,N_8086);
nand U8238 (N_8238,N_8118,N_8076);
nor U8239 (N_8239,N_8126,N_8152);
and U8240 (N_8240,N_8059,N_8096);
and U8241 (N_8241,N_8143,N_8007);
or U8242 (N_8242,N_8138,N_8091);
nand U8243 (N_8243,N_8083,N_8088);
nand U8244 (N_8244,N_8130,N_8050);
nor U8245 (N_8245,N_8065,N_8191);
nor U8246 (N_8246,N_8161,N_8019);
and U8247 (N_8247,N_8031,N_8074);
and U8248 (N_8248,N_8023,N_8117);
and U8249 (N_8249,N_8162,N_8030);
nor U8250 (N_8250,N_8107,N_8109);
and U8251 (N_8251,N_8024,N_8020);
and U8252 (N_8252,N_8013,N_8192);
xor U8253 (N_8253,N_8193,N_8136);
xnor U8254 (N_8254,N_8194,N_8180);
nand U8255 (N_8255,N_8102,N_8139);
nand U8256 (N_8256,N_8133,N_8025);
nand U8257 (N_8257,N_8112,N_8080);
or U8258 (N_8258,N_8184,N_8134);
nand U8259 (N_8259,N_8189,N_8069);
or U8260 (N_8260,N_8045,N_8003);
nand U8261 (N_8261,N_8174,N_8144);
nand U8262 (N_8262,N_8046,N_8063);
nor U8263 (N_8263,N_8034,N_8198);
or U8264 (N_8264,N_8156,N_8122);
or U8265 (N_8265,N_8022,N_8175);
nand U8266 (N_8266,N_8087,N_8158);
or U8267 (N_8267,N_8001,N_8101);
nor U8268 (N_8268,N_8053,N_8171);
and U8269 (N_8269,N_8155,N_8058);
nor U8270 (N_8270,N_8120,N_8197);
and U8271 (N_8271,N_8084,N_8068);
or U8272 (N_8272,N_8121,N_8179);
nand U8273 (N_8273,N_8048,N_8199);
or U8274 (N_8274,N_8079,N_8177);
nor U8275 (N_8275,N_8163,N_8054);
and U8276 (N_8276,N_8043,N_8115);
or U8277 (N_8277,N_8116,N_8047);
nor U8278 (N_8278,N_8185,N_8106);
nand U8279 (N_8279,N_8051,N_8182);
nand U8280 (N_8280,N_8142,N_8085);
or U8281 (N_8281,N_8146,N_8111);
nand U8282 (N_8282,N_8052,N_8060);
and U8283 (N_8283,N_8098,N_8021);
nand U8284 (N_8284,N_8005,N_8150);
and U8285 (N_8285,N_8165,N_8035);
nand U8286 (N_8286,N_8000,N_8104);
or U8287 (N_8287,N_8078,N_8066);
nor U8288 (N_8288,N_8100,N_8094);
nor U8289 (N_8289,N_8167,N_8149);
nand U8290 (N_8290,N_8090,N_8123);
nand U8291 (N_8291,N_8061,N_8124);
and U8292 (N_8292,N_8012,N_8055);
or U8293 (N_8293,N_8164,N_8108);
and U8294 (N_8294,N_8077,N_8137);
nor U8295 (N_8295,N_8147,N_8157);
xor U8296 (N_8296,N_8018,N_8042);
nor U8297 (N_8297,N_8181,N_8103);
and U8298 (N_8298,N_8015,N_8169);
and U8299 (N_8299,N_8113,N_8032);
and U8300 (N_8300,N_8006,N_8053);
or U8301 (N_8301,N_8018,N_8115);
nand U8302 (N_8302,N_8180,N_8182);
or U8303 (N_8303,N_8094,N_8111);
nand U8304 (N_8304,N_8136,N_8194);
nand U8305 (N_8305,N_8062,N_8096);
xnor U8306 (N_8306,N_8134,N_8002);
or U8307 (N_8307,N_8153,N_8169);
and U8308 (N_8308,N_8008,N_8088);
or U8309 (N_8309,N_8019,N_8139);
xor U8310 (N_8310,N_8063,N_8126);
nand U8311 (N_8311,N_8144,N_8115);
nand U8312 (N_8312,N_8179,N_8034);
nand U8313 (N_8313,N_8014,N_8152);
or U8314 (N_8314,N_8038,N_8133);
xor U8315 (N_8315,N_8091,N_8160);
and U8316 (N_8316,N_8101,N_8017);
nand U8317 (N_8317,N_8069,N_8041);
nand U8318 (N_8318,N_8122,N_8051);
and U8319 (N_8319,N_8084,N_8023);
or U8320 (N_8320,N_8195,N_8036);
or U8321 (N_8321,N_8068,N_8025);
and U8322 (N_8322,N_8062,N_8021);
nor U8323 (N_8323,N_8089,N_8143);
xor U8324 (N_8324,N_8033,N_8147);
and U8325 (N_8325,N_8015,N_8077);
and U8326 (N_8326,N_8157,N_8113);
nor U8327 (N_8327,N_8141,N_8014);
nor U8328 (N_8328,N_8013,N_8086);
nor U8329 (N_8329,N_8106,N_8014);
nand U8330 (N_8330,N_8141,N_8083);
or U8331 (N_8331,N_8161,N_8075);
or U8332 (N_8332,N_8145,N_8001);
or U8333 (N_8333,N_8023,N_8057);
or U8334 (N_8334,N_8091,N_8082);
or U8335 (N_8335,N_8049,N_8048);
nand U8336 (N_8336,N_8175,N_8089);
nor U8337 (N_8337,N_8134,N_8008);
and U8338 (N_8338,N_8065,N_8097);
nor U8339 (N_8339,N_8071,N_8156);
and U8340 (N_8340,N_8068,N_8197);
or U8341 (N_8341,N_8069,N_8028);
nor U8342 (N_8342,N_8001,N_8176);
nand U8343 (N_8343,N_8109,N_8121);
nand U8344 (N_8344,N_8019,N_8180);
nor U8345 (N_8345,N_8029,N_8004);
and U8346 (N_8346,N_8113,N_8034);
and U8347 (N_8347,N_8065,N_8117);
and U8348 (N_8348,N_8022,N_8189);
and U8349 (N_8349,N_8056,N_8119);
or U8350 (N_8350,N_8020,N_8049);
and U8351 (N_8351,N_8110,N_8155);
nor U8352 (N_8352,N_8010,N_8146);
or U8353 (N_8353,N_8076,N_8014);
nor U8354 (N_8354,N_8143,N_8091);
nand U8355 (N_8355,N_8127,N_8170);
nor U8356 (N_8356,N_8140,N_8124);
nor U8357 (N_8357,N_8193,N_8100);
nor U8358 (N_8358,N_8167,N_8044);
or U8359 (N_8359,N_8009,N_8138);
nor U8360 (N_8360,N_8027,N_8108);
xor U8361 (N_8361,N_8160,N_8052);
nand U8362 (N_8362,N_8035,N_8182);
and U8363 (N_8363,N_8184,N_8060);
nand U8364 (N_8364,N_8107,N_8097);
and U8365 (N_8365,N_8138,N_8104);
nand U8366 (N_8366,N_8122,N_8182);
and U8367 (N_8367,N_8105,N_8037);
and U8368 (N_8368,N_8002,N_8074);
nor U8369 (N_8369,N_8119,N_8059);
nor U8370 (N_8370,N_8143,N_8082);
nand U8371 (N_8371,N_8092,N_8000);
nor U8372 (N_8372,N_8127,N_8081);
and U8373 (N_8373,N_8030,N_8106);
nor U8374 (N_8374,N_8121,N_8113);
nor U8375 (N_8375,N_8008,N_8121);
and U8376 (N_8376,N_8077,N_8036);
nand U8377 (N_8377,N_8136,N_8158);
nand U8378 (N_8378,N_8158,N_8011);
nor U8379 (N_8379,N_8092,N_8162);
nor U8380 (N_8380,N_8160,N_8143);
nand U8381 (N_8381,N_8005,N_8082);
nor U8382 (N_8382,N_8164,N_8197);
nand U8383 (N_8383,N_8143,N_8156);
nor U8384 (N_8384,N_8185,N_8160);
xor U8385 (N_8385,N_8050,N_8062);
and U8386 (N_8386,N_8054,N_8023);
nand U8387 (N_8387,N_8113,N_8106);
or U8388 (N_8388,N_8081,N_8048);
nand U8389 (N_8389,N_8124,N_8077);
nand U8390 (N_8390,N_8031,N_8166);
or U8391 (N_8391,N_8128,N_8118);
or U8392 (N_8392,N_8109,N_8165);
nand U8393 (N_8393,N_8167,N_8143);
nor U8394 (N_8394,N_8000,N_8009);
nor U8395 (N_8395,N_8070,N_8106);
and U8396 (N_8396,N_8007,N_8058);
nand U8397 (N_8397,N_8012,N_8148);
nor U8398 (N_8398,N_8161,N_8009);
or U8399 (N_8399,N_8017,N_8134);
nand U8400 (N_8400,N_8315,N_8210);
or U8401 (N_8401,N_8243,N_8206);
xor U8402 (N_8402,N_8270,N_8331);
and U8403 (N_8403,N_8235,N_8241);
nand U8404 (N_8404,N_8324,N_8397);
nand U8405 (N_8405,N_8248,N_8321);
and U8406 (N_8406,N_8220,N_8310);
and U8407 (N_8407,N_8381,N_8377);
and U8408 (N_8408,N_8382,N_8295);
and U8409 (N_8409,N_8223,N_8246);
nand U8410 (N_8410,N_8262,N_8301);
nor U8411 (N_8411,N_8390,N_8290);
nand U8412 (N_8412,N_8352,N_8387);
nand U8413 (N_8413,N_8398,N_8392);
nor U8414 (N_8414,N_8298,N_8354);
and U8415 (N_8415,N_8329,N_8353);
nor U8416 (N_8416,N_8304,N_8244);
nand U8417 (N_8417,N_8362,N_8231);
and U8418 (N_8418,N_8372,N_8228);
nand U8419 (N_8419,N_8212,N_8396);
and U8420 (N_8420,N_8322,N_8388);
nand U8421 (N_8421,N_8303,N_8389);
or U8422 (N_8422,N_8317,N_8217);
or U8423 (N_8423,N_8211,N_8232);
and U8424 (N_8424,N_8383,N_8376);
nor U8425 (N_8425,N_8334,N_8345);
or U8426 (N_8426,N_8238,N_8374);
nand U8427 (N_8427,N_8339,N_8245);
nand U8428 (N_8428,N_8393,N_8325);
or U8429 (N_8429,N_8259,N_8332);
and U8430 (N_8430,N_8282,N_8385);
nand U8431 (N_8431,N_8313,N_8305);
nor U8432 (N_8432,N_8285,N_8263);
or U8433 (N_8433,N_8268,N_8279);
or U8434 (N_8434,N_8375,N_8316);
and U8435 (N_8435,N_8288,N_8275);
or U8436 (N_8436,N_8373,N_8337);
and U8437 (N_8437,N_8336,N_8266);
nand U8438 (N_8438,N_8308,N_8363);
nand U8439 (N_8439,N_8394,N_8277);
or U8440 (N_8440,N_8328,N_8378);
nand U8441 (N_8441,N_8204,N_8391);
or U8442 (N_8442,N_8330,N_8384);
nand U8443 (N_8443,N_8380,N_8309);
or U8444 (N_8444,N_8239,N_8344);
or U8445 (N_8445,N_8359,N_8364);
nand U8446 (N_8446,N_8343,N_8254);
or U8447 (N_8447,N_8251,N_8236);
and U8448 (N_8448,N_8205,N_8318);
nand U8449 (N_8449,N_8272,N_8300);
nor U8450 (N_8450,N_8255,N_8323);
nand U8451 (N_8451,N_8368,N_8289);
nand U8452 (N_8452,N_8214,N_8286);
nand U8453 (N_8453,N_8260,N_8327);
and U8454 (N_8454,N_8370,N_8297);
nand U8455 (N_8455,N_8348,N_8225);
or U8456 (N_8456,N_8201,N_8209);
nor U8457 (N_8457,N_8213,N_8219);
nand U8458 (N_8458,N_8215,N_8274);
and U8459 (N_8459,N_8216,N_8273);
nor U8460 (N_8460,N_8267,N_8347);
or U8461 (N_8461,N_8287,N_8346);
xor U8462 (N_8462,N_8256,N_8230);
and U8463 (N_8463,N_8257,N_8357);
and U8464 (N_8464,N_8261,N_8292);
and U8465 (N_8465,N_8367,N_8320);
and U8466 (N_8466,N_8226,N_8240);
and U8467 (N_8467,N_8366,N_8229);
or U8468 (N_8468,N_8293,N_8283);
or U8469 (N_8469,N_8218,N_8386);
or U8470 (N_8470,N_8264,N_8371);
nor U8471 (N_8471,N_8342,N_8302);
nor U8472 (N_8472,N_8356,N_8291);
nor U8473 (N_8473,N_8314,N_8233);
nor U8474 (N_8474,N_8227,N_8207);
or U8475 (N_8475,N_8281,N_8258);
and U8476 (N_8476,N_8242,N_8249);
nor U8477 (N_8477,N_8369,N_8224);
nor U8478 (N_8478,N_8276,N_8306);
xor U8479 (N_8479,N_8247,N_8203);
and U8480 (N_8480,N_8294,N_8338);
or U8481 (N_8481,N_8307,N_8221);
or U8482 (N_8482,N_8335,N_8312);
or U8483 (N_8483,N_8319,N_8299);
or U8484 (N_8484,N_8311,N_8202);
or U8485 (N_8485,N_8355,N_8358);
and U8486 (N_8486,N_8341,N_8200);
nor U8487 (N_8487,N_8326,N_8351);
nand U8488 (N_8488,N_8208,N_8252);
or U8489 (N_8489,N_8360,N_8284);
and U8490 (N_8490,N_8222,N_8379);
nand U8491 (N_8491,N_8395,N_8269);
nand U8492 (N_8492,N_8237,N_8399);
or U8493 (N_8493,N_8271,N_8296);
nand U8494 (N_8494,N_8253,N_8350);
or U8495 (N_8495,N_8250,N_8340);
nand U8496 (N_8496,N_8234,N_8278);
and U8497 (N_8497,N_8265,N_8333);
or U8498 (N_8498,N_8365,N_8361);
and U8499 (N_8499,N_8349,N_8280);
nor U8500 (N_8500,N_8274,N_8251);
or U8501 (N_8501,N_8249,N_8301);
nand U8502 (N_8502,N_8301,N_8278);
and U8503 (N_8503,N_8271,N_8382);
and U8504 (N_8504,N_8273,N_8395);
xor U8505 (N_8505,N_8290,N_8293);
nand U8506 (N_8506,N_8227,N_8283);
nand U8507 (N_8507,N_8281,N_8221);
or U8508 (N_8508,N_8320,N_8201);
or U8509 (N_8509,N_8222,N_8360);
nor U8510 (N_8510,N_8227,N_8206);
nor U8511 (N_8511,N_8231,N_8313);
or U8512 (N_8512,N_8378,N_8290);
and U8513 (N_8513,N_8338,N_8385);
nor U8514 (N_8514,N_8269,N_8378);
and U8515 (N_8515,N_8365,N_8320);
nand U8516 (N_8516,N_8206,N_8278);
nor U8517 (N_8517,N_8261,N_8242);
nand U8518 (N_8518,N_8297,N_8391);
nand U8519 (N_8519,N_8294,N_8249);
and U8520 (N_8520,N_8388,N_8217);
or U8521 (N_8521,N_8383,N_8231);
nor U8522 (N_8522,N_8283,N_8364);
and U8523 (N_8523,N_8351,N_8331);
nand U8524 (N_8524,N_8263,N_8278);
nor U8525 (N_8525,N_8316,N_8243);
and U8526 (N_8526,N_8295,N_8219);
xor U8527 (N_8527,N_8216,N_8221);
or U8528 (N_8528,N_8280,N_8371);
nand U8529 (N_8529,N_8393,N_8363);
nor U8530 (N_8530,N_8356,N_8229);
nand U8531 (N_8531,N_8330,N_8210);
or U8532 (N_8532,N_8306,N_8328);
or U8533 (N_8533,N_8324,N_8246);
nand U8534 (N_8534,N_8373,N_8281);
and U8535 (N_8535,N_8386,N_8383);
nand U8536 (N_8536,N_8212,N_8252);
nand U8537 (N_8537,N_8327,N_8377);
or U8538 (N_8538,N_8386,N_8348);
nor U8539 (N_8539,N_8286,N_8362);
nor U8540 (N_8540,N_8309,N_8391);
xor U8541 (N_8541,N_8249,N_8303);
nor U8542 (N_8542,N_8320,N_8324);
nand U8543 (N_8543,N_8222,N_8349);
or U8544 (N_8544,N_8393,N_8257);
nand U8545 (N_8545,N_8292,N_8364);
nor U8546 (N_8546,N_8259,N_8327);
and U8547 (N_8547,N_8395,N_8303);
nor U8548 (N_8548,N_8382,N_8398);
and U8549 (N_8549,N_8379,N_8209);
nor U8550 (N_8550,N_8247,N_8375);
or U8551 (N_8551,N_8320,N_8368);
or U8552 (N_8552,N_8219,N_8234);
and U8553 (N_8553,N_8241,N_8269);
xor U8554 (N_8554,N_8324,N_8348);
or U8555 (N_8555,N_8373,N_8322);
xnor U8556 (N_8556,N_8205,N_8346);
nor U8557 (N_8557,N_8317,N_8386);
nor U8558 (N_8558,N_8303,N_8279);
and U8559 (N_8559,N_8312,N_8377);
xnor U8560 (N_8560,N_8343,N_8298);
nor U8561 (N_8561,N_8231,N_8217);
nand U8562 (N_8562,N_8331,N_8263);
and U8563 (N_8563,N_8323,N_8247);
xor U8564 (N_8564,N_8204,N_8308);
nand U8565 (N_8565,N_8300,N_8271);
xor U8566 (N_8566,N_8377,N_8361);
nor U8567 (N_8567,N_8209,N_8322);
and U8568 (N_8568,N_8256,N_8235);
or U8569 (N_8569,N_8222,N_8257);
or U8570 (N_8570,N_8271,N_8359);
nor U8571 (N_8571,N_8207,N_8388);
and U8572 (N_8572,N_8202,N_8347);
or U8573 (N_8573,N_8376,N_8384);
nor U8574 (N_8574,N_8253,N_8396);
or U8575 (N_8575,N_8265,N_8271);
nand U8576 (N_8576,N_8283,N_8260);
nand U8577 (N_8577,N_8357,N_8245);
xnor U8578 (N_8578,N_8399,N_8381);
nor U8579 (N_8579,N_8316,N_8269);
or U8580 (N_8580,N_8234,N_8360);
or U8581 (N_8581,N_8228,N_8336);
or U8582 (N_8582,N_8232,N_8225);
and U8583 (N_8583,N_8247,N_8250);
and U8584 (N_8584,N_8369,N_8394);
nor U8585 (N_8585,N_8396,N_8271);
xnor U8586 (N_8586,N_8351,N_8210);
xor U8587 (N_8587,N_8328,N_8284);
xnor U8588 (N_8588,N_8273,N_8364);
or U8589 (N_8589,N_8298,N_8280);
and U8590 (N_8590,N_8225,N_8392);
nor U8591 (N_8591,N_8204,N_8338);
nor U8592 (N_8592,N_8267,N_8212);
nor U8593 (N_8593,N_8341,N_8238);
or U8594 (N_8594,N_8359,N_8366);
and U8595 (N_8595,N_8263,N_8231);
or U8596 (N_8596,N_8338,N_8354);
nor U8597 (N_8597,N_8398,N_8321);
nor U8598 (N_8598,N_8277,N_8243);
nand U8599 (N_8599,N_8253,N_8255);
nand U8600 (N_8600,N_8466,N_8539);
nand U8601 (N_8601,N_8527,N_8549);
and U8602 (N_8602,N_8495,N_8427);
nand U8603 (N_8603,N_8405,N_8449);
nand U8604 (N_8604,N_8580,N_8410);
nor U8605 (N_8605,N_8534,N_8591);
nor U8606 (N_8606,N_8494,N_8576);
or U8607 (N_8607,N_8447,N_8548);
xor U8608 (N_8608,N_8503,N_8565);
or U8609 (N_8609,N_8438,N_8516);
nor U8610 (N_8610,N_8493,N_8560);
nand U8611 (N_8611,N_8451,N_8513);
nor U8612 (N_8612,N_8543,N_8412);
and U8613 (N_8613,N_8409,N_8448);
and U8614 (N_8614,N_8597,N_8505);
nor U8615 (N_8615,N_8423,N_8538);
nand U8616 (N_8616,N_8568,N_8426);
and U8617 (N_8617,N_8564,N_8434);
and U8618 (N_8618,N_8422,N_8402);
nor U8619 (N_8619,N_8478,N_8462);
nand U8620 (N_8620,N_8441,N_8429);
nor U8621 (N_8621,N_8418,N_8574);
and U8622 (N_8622,N_8444,N_8452);
or U8623 (N_8623,N_8512,N_8443);
or U8624 (N_8624,N_8558,N_8545);
nor U8625 (N_8625,N_8599,N_8431);
or U8626 (N_8626,N_8453,N_8459);
and U8627 (N_8627,N_8509,N_8463);
or U8628 (N_8628,N_8585,N_8562);
nand U8629 (N_8629,N_8544,N_8592);
or U8630 (N_8630,N_8432,N_8595);
nor U8631 (N_8631,N_8456,N_8598);
nor U8632 (N_8632,N_8581,N_8587);
and U8633 (N_8633,N_8589,N_8472);
nand U8634 (N_8634,N_8570,N_8556);
nor U8635 (N_8635,N_8442,N_8572);
nand U8636 (N_8636,N_8465,N_8579);
nor U8637 (N_8637,N_8460,N_8566);
or U8638 (N_8638,N_8501,N_8473);
and U8639 (N_8639,N_8553,N_8490);
or U8640 (N_8640,N_8497,N_8520);
or U8641 (N_8641,N_8486,N_8455);
nor U8642 (N_8642,N_8590,N_8425);
nand U8643 (N_8643,N_8530,N_8559);
and U8644 (N_8644,N_8525,N_8415);
nor U8645 (N_8645,N_8540,N_8414);
or U8646 (N_8646,N_8511,N_8502);
or U8647 (N_8647,N_8420,N_8521);
nand U8648 (N_8648,N_8467,N_8489);
nand U8649 (N_8649,N_8428,N_8535);
or U8650 (N_8650,N_8424,N_8471);
nand U8651 (N_8651,N_8468,N_8541);
or U8652 (N_8652,N_8474,N_8557);
and U8653 (N_8653,N_8546,N_8496);
nor U8654 (N_8654,N_8523,N_8584);
nand U8655 (N_8655,N_8536,N_8481);
nor U8656 (N_8656,N_8485,N_8488);
nor U8657 (N_8657,N_8404,N_8437);
and U8658 (N_8658,N_8407,N_8419);
nor U8659 (N_8659,N_8533,N_8479);
nor U8660 (N_8660,N_8596,N_8406);
nor U8661 (N_8661,N_8561,N_8573);
nand U8662 (N_8662,N_8586,N_8484);
nand U8663 (N_8663,N_8400,N_8436);
or U8664 (N_8664,N_8480,N_8524);
nand U8665 (N_8665,N_8499,N_8475);
nor U8666 (N_8666,N_8517,N_8445);
nand U8667 (N_8667,N_8551,N_8594);
nand U8668 (N_8668,N_8550,N_8450);
and U8669 (N_8669,N_8408,N_8498);
nor U8670 (N_8670,N_8518,N_8440);
and U8671 (N_8671,N_8542,N_8582);
nor U8672 (N_8672,N_8457,N_8492);
and U8673 (N_8673,N_8529,N_8411);
or U8674 (N_8674,N_8433,N_8401);
nor U8675 (N_8675,N_8403,N_8464);
nor U8676 (N_8676,N_8417,N_8476);
nand U8677 (N_8677,N_8416,N_8430);
and U8678 (N_8678,N_8507,N_8446);
xor U8679 (N_8679,N_8528,N_8577);
and U8680 (N_8680,N_8413,N_8515);
and U8681 (N_8681,N_8563,N_8458);
or U8682 (N_8682,N_8555,N_8439);
or U8683 (N_8683,N_8593,N_8519);
nand U8684 (N_8684,N_8575,N_8526);
nand U8685 (N_8685,N_8537,N_8491);
nand U8686 (N_8686,N_8547,N_8487);
and U8687 (N_8687,N_8421,N_8552);
or U8688 (N_8688,N_8500,N_8435);
xnor U8689 (N_8689,N_8510,N_8583);
and U8690 (N_8690,N_8571,N_8567);
nor U8691 (N_8691,N_8514,N_8554);
and U8692 (N_8692,N_8461,N_8477);
nor U8693 (N_8693,N_8470,N_8532);
and U8694 (N_8694,N_8506,N_8578);
nor U8695 (N_8695,N_8482,N_8588);
and U8696 (N_8696,N_8483,N_8504);
nand U8697 (N_8697,N_8569,N_8469);
nor U8698 (N_8698,N_8454,N_8508);
and U8699 (N_8699,N_8522,N_8531);
nor U8700 (N_8700,N_8553,N_8536);
nor U8701 (N_8701,N_8438,N_8424);
xnor U8702 (N_8702,N_8561,N_8483);
and U8703 (N_8703,N_8514,N_8461);
and U8704 (N_8704,N_8425,N_8441);
or U8705 (N_8705,N_8453,N_8559);
or U8706 (N_8706,N_8488,N_8439);
or U8707 (N_8707,N_8458,N_8400);
nor U8708 (N_8708,N_8545,N_8444);
nand U8709 (N_8709,N_8464,N_8538);
nor U8710 (N_8710,N_8556,N_8597);
nor U8711 (N_8711,N_8409,N_8487);
or U8712 (N_8712,N_8569,N_8471);
nand U8713 (N_8713,N_8437,N_8594);
or U8714 (N_8714,N_8515,N_8494);
nand U8715 (N_8715,N_8440,N_8510);
and U8716 (N_8716,N_8413,N_8565);
xor U8717 (N_8717,N_8565,N_8421);
nand U8718 (N_8718,N_8427,N_8468);
nand U8719 (N_8719,N_8534,N_8497);
nand U8720 (N_8720,N_8492,N_8581);
or U8721 (N_8721,N_8433,N_8442);
or U8722 (N_8722,N_8497,N_8473);
or U8723 (N_8723,N_8541,N_8402);
xor U8724 (N_8724,N_8463,N_8595);
xor U8725 (N_8725,N_8441,N_8498);
and U8726 (N_8726,N_8592,N_8453);
nand U8727 (N_8727,N_8528,N_8551);
nand U8728 (N_8728,N_8418,N_8441);
nor U8729 (N_8729,N_8513,N_8405);
nand U8730 (N_8730,N_8406,N_8585);
and U8731 (N_8731,N_8530,N_8416);
nand U8732 (N_8732,N_8580,N_8555);
and U8733 (N_8733,N_8473,N_8410);
nor U8734 (N_8734,N_8524,N_8572);
xnor U8735 (N_8735,N_8488,N_8508);
and U8736 (N_8736,N_8599,N_8548);
or U8737 (N_8737,N_8589,N_8460);
and U8738 (N_8738,N_8422,N_8566);
nor U8739 (N_8739,N_8582,N_8432);
or U8740 (N_8740,N_8594,N_8417);
and U8741 (N_8741,N_8403,N_8515);
nor U8742 (N_8742,N_8472,N_8543);
and U8743 (N_8743,N_8581,N_8467);
or U8744 (N_8744,N_8428,N_8536);
or U8745 (N_8745,N_8533,N_8424);
or U8746 (N_8746,N_8512,N_8508);
nor U8747 (N_8747,N_8527,N_8577);
nand U8748 (N_8748,N_8546,N_8512);
nor U8749 (N_8749,N_8472,N_8490);
xor U8750 (N_8750,N_8451,N_8476);
nand U8751 (N_8751,N_8405,N_8540);
nand U8752 (N_8752,N_8402,N_8452);
and U8753 (N_8753,N_8598,N_8481);
nand U8754 (N_8754,N_8529,N_8447);
nand U8755 (N_8755,N_8465,N_8420);
or U8756 (N_8756,N_8598,N_8589);
nor U8757 (N_8757,N_8532,N_8579);
and U8758 (N_8758,N_8471,N_8472);
and U8759 (N_8759,N_8592,N_8474);
nand U8760 (N_8760,N_8508,N_8505);
and U8761 (N_8761,N_8440,N_8454);
nand U8762 (N_8762,N_8417,N_8475);
nand U8763 (N_8763,N_8466,N_8412);
and U8764 (N_8764,N_8425,N_8583);
nor U8765 (N_8765,N_8451,N_8430);
or U8766 (N_8766,N_8471,N_8481);
and U8767 (N_8767,N_8575,N_8426);
nor U8768 (N_8768,N_8432,N_8556);
or U8769 (N_8769,N_8438,N_8556);
nand U8770 (N_8770,N_8546,N_8455);
or U8771 (N_8771,N_8440,N_8412);
or U8772 (N_8772,N_8460,N_8405);
nand U8773 (N_8773,N_8421,N_8562);
nand U8774 (N_8774,N_8549,N_8427);
or U8775 (N_8775,N_8511,N_8418);
and U8776 (N_8776,N_8582,N_8458);
nor U8777 (N_8777,N_8509,N_8593);
nand U8778 (N_8778,N_8594,N_8599);
nand U8779 (N_8779,N_8530,N_8460);
nor U8780 (N_8780,N_8530,N_8476);
nand U8781 (N_8781,N_8434,N_8536);
and U8782 (N_8782,N_8455,N_8469);
and U8783 (N_8783,N_8430,N_8565);
nand U8784 (N_8784,N_8418,N_8461);
nand U8785 (N_8785,N_8527,N_8429);
or U8786 (N_8786,N_8404,N_8522);
nand U8787 (N_8787,N_8429,N_8594);
and U8788 (N_8788,N_8462,N_8490);
nor U8789 (N_8789,N_8567,N_8502);
nor U8790 (N_8790,N_8435,N_8401);
and U8791 (N_8791,N_8445,N_8430);
nor U8792 (N_8792,N_8596,N_8525);
nor U8793 (N_8793,N_8449,N_8571);
nand U8794 (N_8794,N_8476,N_8487);
or U8795 (N_8795,N_8483,N_8458);
and U8796 (N_8796,N_8569,N_8581);
and U8797 (N_8797,N_8588,N_8507);
nor U8798 (N_8798,N_8436,N_8572);
nand U8799 (N_8799,N_8475,N_8542);
and U8800 (N_8800,N_8701,N_8727);
nand U8801 (N_8801,N_8610,N_8744);
nand U8802 (N_8802,N_8723,N_8757);
nand U8803 (N_8803,N_8605,N_8709);
nor U8804 (N_8804,N_8663,N_8661);
and U8805 (N_8805,N_8720,N_8759);
nor U8806 (N_8806,N_8785,N_8674);
nand U8807 (N_8807,N_8717,N_8637);
nor U8808 (N_8808,N_8747,N_8707);
nand U8809 (N_8809,N_8774,N_8602);
nand U8810 (N_8810,N_8629,N_8725);
or U8811 (N_8811,N_8606,N_8765);
nand U8812 (N_8812,N_8746,N_8703);
nand U8813 (N_8813,N_8776,N_8706);
nor U8814 (N_8814,N_8694,N_8611);
and U8815 (N_8815,N_8754,N_8688);
nor U8816 (N_8816,N_8787,N_8702);
and U8817 (N_8817,N_8639,N_8645);
nor U8818 (N_8818,N_8761,N_8788);
nor U8819 (N_8819,N_8786,N_8685);
nor U8820 (N_8820,N_8671,N_8609);
nand U8821 (N_8821,N_8714,N_8771);
or U8822 (N_8822,N_8737,N_8648);
or U8823 (N_8823,N_8656,N_8697);
and U8824 (N_8824,N_8781,N_8740);
xor U8825 (N_8825,N_8768,N_8753);
nand U8826 (N_8826,N_8796,N_8735);
nor U8827 (N_8827,N_8751,N_8724);
nor U8828 (N_8828,N_8764,N_8794);
and U8829 (N_8829,N_8658,N_8732);
or U8830 (N_8830,N_8615,N_8626);
nand U8831 (N_8831,N_8687,N_8792);
nand U8832 (N_8832,N_8614,N_8722);
nand U8833 (N_8833,N_8670,N_8651);
xor U8834 (N_8834,N_8635,N_8642);
or U8835 (N_8835,N_8716,N_8782);
and U8836 (N_8836,N_8721,N_8621);
nand U8837 (N_8837,N_8742,N_8649);
or U8838 (N_8838,N_8601,N_8719);
or U8839 (N_8839,N_8631,N_8692);
and U8840 (N_8840,N_8691,N_8627);
nand U8841 (N_8841,N_8767,N_8750);
or U8842 (N_8842,N_8666,N_8779);
nand U8843 (N_8843,N_8681,N_8693);
nor U8844 (N_8844,N_8608,N_8680);
xor U8845 (N_8845,N_8676,N_8791);
or U8846 (N_8846,N_8797,N_8736);
nand U8847 (N_8847,N_8769,N_8780);
nor U8848 (N_8848,N_8755,N_8738);
and U8849 (N_8849,N_8654,N_8600);
xor U8850 (N_8850,N_8726,N_8766);
nand U8851 (N_8851,N_8728,N_8662);
nand U8852 (N_8852,N_8660,N_8798);
or U8853 (N_8853,N_8778,N_8657);
and U8854 (N_8854,N_8730,N_8665);
xor U8855 (N_8855,N_8760,N_8695);
nor U8856 (N_8856,N_8650,N_8777);
xnor U8857 (N_8857,N_8700,N_8603);
nand U8858 (N_8858,N_8604,N_8679);
and U8859 (N_8859,N_8667,N_8734);
or U8860 (N_8860,N_8718,N_8655);
or U8861 (N_8861,N_8644,N_8628);
or U8862 (N_8862,N_8741,N_8756);
nor U8863 (N_8863,N_8748,N_8715);
and U8864 (N_8864,N_8638,N_8773);
or U8865 (N_8865,N_8618,N_8624);
nand U8866 (N_8866,N_8607,N_8731);
or U8867 (N_8867,N_8711,N_8683);
and U8868 (N_8868,N_8659,N_8708);
nand U8869 (N_8869,N_8641,N_8617);
or U8870 (N_8870,N_8619,N_8699);
nand U8871 (N_8871,N_8673,N_8682);
or U8872 (N_8872,N_8646,N_8770);
or U8873 (N_8873,N_8678,N_8672);
nand U8874 (N_8874,N_8668,N_8799);
nand U8875 (N_8875,N_8643,N_8647);
nor U8876 (N_8876,N_8784,N_8743);
nor U8877 (N_8877,N_8783,N_8795);
and U8878 (N_8878,N_8775,N_8653);
and U8879 (N_8879,N_8762,N_8632);
or U8880 (N_8880,N_8636,N_8675);
nand U8881 (N_8881,N_8669,N_8704);
nor U8882 (N_8882,N_8739,N_8652);
and U8883 (N_8883,N_8623,N_8745);
and U8884 (N_8884,N_8640,N_8758);
or U8885 (N_8885,N_8625,N_8763);
or U8886 (N_8886,N_8705,N_8664);
nand U8887 (N_8887,N_8616,N_8749);
and U8888 (N_8888,N_8712,N_8622);
nand U8889 (N_8889,N_8634,N_8613);
nor U8890 (N_8890,N_8713,N_8698);
nor U8891 (N_8891,N_8686,N_8690);
and U8892 (N_8892,N_8789,N_8684);
nor U8893 (N_8893,N_8677,N_8630);
nand U8894 (N_8894,N_8752,N_8612);
or U8895 (N_8895,N_8710,N_8790);
nand U8896 (N_8896,N_8689,N_8620);
nand U8897 (N_8897,N_8772,N_8729);
or U8898 (N_8898,N_8696,N_8633);
or U8899 (N_8899,N_8733,N_8793);
nand U8900 (N_8900,N_8723,N_8683);
and U8901 (N_8901,N_8755,N_8661);
nand U8902 (N_8902,N_8601,N_8625);
nor U8903 (N_8903,N_8733,N_8725);
and U8904 (N_8904,N_8773,N_8616);
nor U8905 (N_8905,N_8765,N_8635);
nor U8906 (N_8906,N_8667,N_8648);
xnor U8907 (N_8907,N_8691,N_8738);
nor U8908 (N_8908,N_8755,N_8679);
nand U8909 (N_8909,N_8638,N_8780);
nand U8910 (N_8910,N_8608,N_8709);
nor U8911 (N_8911,N_8791,N_8772);
and U8912 (N_8912,N_8627,N_8652);
nor U8913 (N_8913,N_8789,N_8760);
nor U8914 (N_8914,N_8755,N_8715);
nor U8915 (N_8915,N_8652,N_8768);
nand U8916 (N_8916,N_8680,N_8686);
or U8917 (N_8917,N_8731,N_8768);
nor U8918 (N_8918,N_8711,N_8695);
and U8919 (N_8919,N_8710,N_8701);
nand U8920 (N_8920,N_8757,N_8694);
and U8921 (N_8921,N_8674,N_8617);
or U8922 (N_8922,N_8773,N_8615);
nor U8923 (N_8923,N_8644,N_8710);
and U8924 (N_8924,N_8714,N_8717);
xor U8925 (N_8925,N_8632,N_8735);
and U8926 (N_8926,N_8646,N_8687);
nand U8927 (N_8927,N_8787,N_8713);
xnor U8928 (N_8928,N_8719,N_8672);
nand U8929 (N_8929,N_8717,N_8773);
nand U8930 (N_8930,N_8753,N_8614);
or U8931 (N_8931,N_8741,N_8686);
and U8932 (N_8932,N_8667,N_8769);
or U8933 (N_8933,N_8647,N_8725);
or U8934 (N_8934,N_8685,N_8725);
and U8935 (N_8935,N_8790,N_8602);
and U8936 (N_8936,N_8758,N_8653);
or U8937 (N_8937,N_8625,N_8757);
and U8938 (N_8938,N_8601,N_8682);
or U8939 (N_8939,N_8773,N_8623);
and U8940 (N_8940,N_8674,N_8677);
or U8941 (N_8941,N_8723,N_8744);
nand U8942 (N_8942,N_8752,N_8650);
and U8943 (N_8943,N_8772,N_8787);
nand U8944 (N_8944,N_8655,N_8794);
and U8945 (N_8945,N_8716,N_8713);
or U8946 (N_8946,N_8717,N_8667);
and U8947 (N_8947,N_8724,N_8621);
and U8948 (N_8948,N_8686,N_8718);
nor U8949 (N_8949,N_8755,N_8635);
and U8950 (N_8950,N_8780,N_8653);
and U8951 (N_8951,N_8613,N_8729);
nand U8952 (N_8952,N_8779,N_8726);
or U8953 (N_8953,N_8769,N_8725);
nand U8954 (N_8954,N_8609,N_8643);
or U8955 (N_8955,N_8742,N_8793);
nor U8956 (N_8956,N_8615,N_8736);
or U8957 (N_8957,N_8786,N_8778);
and U8958 (N_8958,N_8740,N_8611);
xor U8959 (N_8959,N_8656,N_8729);
or U8960 (N_8960,N_8782,N_8662);
nor U8961 (N_8961,N_8745,N_8754);
or U8962 (N_8962,N_8665,N_8673);
nor U8963 (N_8963,N_8643,N_8779);
nand U8964 (N_8964,N_8638,N_8757);
nand U8965 (N_8965,N_8682,N_8614);
or U8966 (N_8966,N_8711,N_8693);
nand U8967 (N_8967,N_8668,N_8781);
or U8968 (N_8968,N_8749,N_8688);
or U8969 (N_8969,N_8742,N_8779);
nor U8970 (N_8970,N_8626,N_8604);
nor U8971 (N_8971,N_8644,N_8739);
nor U8972 (N_8972,N_8782,N_8703);
nor U8973 (N_8973,N_8711,N_8616);
or U8974 (N_8974,N_8627,N_8745);
and U8975 (N_8975,N_8685,N_8611);
nor U8976 (N_8976,N_8768,N_8666);
and U8977 (N_8977,N_8727,N_8613);
nor U8978 (N_8978,N_8612,N_8700);
nor U8979 (N_8979,N_8606,N_8699);
or U8980 (N_8980,N_8630,N_8665);
and U8981 (N_8981,N_8620,N_8608);
and U8982 (N_8982,N_8722,N_8782);
or U8983 (N_8983,N_8647,N_8787);
and U8984 (N_8984,N_8658,N_8674);
and U8985 (N_8985,N_8744,N_8618);
nor U8986 (N_8986,N_8610,N_8798);
or U8987 (N_8987,N_8733,N_8695);
and U8988 (N_8988,N_8699,N_8703);
nor U8989 (N_8989,N_8727,N_8666);
nor U8990 (N_8990,N_8799,N_8724);
nand U8991 (N_8991,N_8691,N_8752);
nor U8992 (N_8992,N_8795,N_8657);
or U8993 (N_8993,N_8629,N_8616);
and U8994 (N_8994,N_8605,N_8799);
or U8995 (N_8995,N_8676,N_8705);
and U8996 (N_8996,N_8622,N_8710);
and U8997 (N_8997,N_8668,N_8612);
nand U8998 (N_8998,N_8701,N_8602);
nand U8999 (N_8999,N_8700,N_8678);
nand U9000 (N_9000,N_8858,N_8902);
nor U9001 (N_9001,N_8997,N_8826);
or U9002 (N_9002,N_8815,N_8832);
nand U9003 (N_9003,N_8831,N_8991);
or U9004 (N_9004,N_8942,N_8953);
or U9005 (N_9005,N_8967,N_8844);
and U9006 (N_9006,N_8913,N_8899);
nor U9007 (N_9007,N_8947,N_8896);
or U9008 (N_9008,N_8936,N_8876);
nand U9009 (N_9009,N_8834,N_8983);
nand U9010 (N_9010,N_8952,N_8962);
nand U9011 (N_9011,N_8880,N_8929);
or U9012 (N_9012,N_8860,N_8809);
nor U9013 (N_9013,N_8872,N_8937);
xor U9014 (N_9014,N_8986,N_8999);
nor U9015 (N_9015,N_8990,N_8811);
or U9016 (N_9016,N_8973,N_8909);
or U9017 (N_9017,N_8919,N_8971);
or U9018 (N_9018,N_8810,N_8804);
nor U9019 (N_9019,N_8821,N_8931);
and U9020 (N_9020,N_8923,N_8958);
and U9021 (N_9021,N_8998,N_8987);
or U9022 (N_9022,N_8842,N_8857);
nand U9023 (N_9023,N_8892,N_8894);
nor U9024 (N_9024,N_8977,N_8945);
nor U9025 (N_9025,N_8814,N_8928);
or U9026 (N_9026,N_8824,N_8841);
or U9027 (N_9027,N_8819,N_8914);
nand U9028 (N_9028,N_8989,N_8884);
nand U9029 (N_9029,N_8870,N_8907);
and U9030 (N_9030,N_8963,N_8956);
xor U9031 (N_9031,N_8935,N_8954);
and U9032 (N_9032,N_8968,N_8996);
nor U9033 (N_9033,N_8966,N_8807);
nor U9034 (N_9034,N_8843,N_8806);
or U9035 (N_9035,N_8949,N_8915);
and U9036 (N_9036,N_8897,N_8964);
nand U9037 (N_9037,N_8845,N_8934);
nand U9038 (N_9038,N_8818,N_8846);
nand U9039 (N_9039,N_8978,N_8995);
nor U9040 (N_9040,N_8893,N_8836);
and U9041 (N_9041,N_8839,N_8885);
or U9042 (N_9042,N_8813,N_8946);
nand U9043 (N_9043,N_8925,N_8980);
or U9044 (N_9044,N_8833,N_8984);
or U9045 (N_9045,N_8840,N_8822);
nor U9046 (N_9046,N_8829,N_8837);
and U9047 (N_9047,N_8911,N_8861);
nand U9048 (N_9048,N_8873,N_8854);
nor U9049 (N_9049,N_8904,N_8835);
nand U9050 (N_9050,N_8939,N_8865);
nor U9051 (N_9051,N_8901,N_8969);
and U9052 (N_9052,N_8887,N_8874);
nor U9053 (N_9053,N_8976,N_8848);
and U9054 (N_9054,N_8888,N_8906);
nand U9055 (N_9055,N_8869,N_8916);
nor U9056 (N_9056,N_8993,N_8917);
nor U9057 (N_9057,N_8940,N_8941);
nor U9058 (N_9058,N_8805,N_8932);
or U9059 (N_9059,N_8988,N_8875);
and U9060 (N_9060,N_8817,N_8852);
nor U9061 (N_9061,N_8982,N_8801);
nor U9062 (N_9062,N_8985,N_8827);
nand U9063 (N_9063,N_8910,N_8957);
nor U9064 (N_9064,N_8802,N_8981);
and U9065 (N_9065,N_8820,N_8992);
and U9066 (N_9066,N_8828,N_8961);
xor U9067 (N_9067,N_8927,N_8849);
nor U9068 (N_9068,N_8933,N_8859);
nor U9069 (N_9069,N_8900,N_8830);
or U9070 (N_9070,N_8944,N_8803);
nand U9071 (N_9071,N_8863,N_8851);
nor U9072 (N_9072,N_8808,N_8951);
or U9073 (N_9073,N_8847,N_8979);
and U9074 (N_9074,N_8879,N_8898);
and U9075 (N_9075,N_8959,N_8889);
nor U9076 (N_9076,N_8867,N_8890);
and U9077 (N_9077,N_8882,N_8930);
and U9078 (N_9078,N_8853,N_8838);
or U9079 (N_9079,N_8943,N_8955);
nor U9080 (N_9080,N_8823,N_8970);
or U9081 (N_9081,N_8866,N_8877);
nor U9082 (N_9082,N_8800,N_8926);
or U9083 (N_9083,N_8871,N_8965);
nor U9084 (N_9084,N_8856,N_8881);
nor U9085 (N_9085,N_8950,N_8924);
nand U9086 (N_9086,N_8972,N_8908);
nor U9087 (N_9087,N_8868,N_8886);
nor U9088 (N_9088,N_8864,N_8975);
nand U9089 (N_9089,N_8974,N_8883);
nor U9090 (N_9090,N_8921,N_8903);
or U9091 (N_9091,N_8918,N_8912);
and U9092 (N_9092,N_8938,N_8862);
or U9093 (N_9093,N_8895,N_8850);
nand U9094 (N_9094,N_8878,N_8948);
nor U9095 (N_9095,N_8812,N_8960);
and U9096 (N_9096,N_8922,N_8920);
or U9097 (N_9097,N_8994,N_8825);
nor U9098 (N_9098,N_8905,N_8816);
nand U9099 (N_9099,N_8891,N_8855);
nor U9100 (N_9100,N_8921,N_8995);
nor U9101 (N_9101,N_8995,N_8824);
and U9102 (N_9102,N_8978,N_8833);
or U9103 (N_9103,N_8973,N_8836);
nand U9104 (N_9104,N_8875,N_8817);
and U9105 (N_9105,N_8846,N_8954);
nor U9106 (N_9106,N_8836,N_8981);
nor U9107 (N_9107,N_8850,N_8817);
nand U9108 (N_9108,N_8843,N_8998);
nand U9109 (N_9109,N_8879,N_8930);
nor U9110 (N_9110,N_8821,N_8918);
nor U9111 (N_9111,N_8986,N_8971);
or U9112 (N_9112,N_8852,N_8864);
nand U9113 (N_9113,N_8965,N_8914);
and U9114 (N_9114,N_8986,N_8871);
nor U9115 (N_9115,N_8834,N_8876);
and U9116 (N_9116,N_8828,N_8956);
nor U9117 (N_9117,N_8840,N_8883);
nand U9118 (N_9118,N_8936,N_8934);
or U9119 (N_9119,N_8927,N_8839);
nor U9120 (N_9120,N_8962,N_8904);
nand U9121 (N_9121,N_8886,N_8904);
and U9122 (N_9122,N_8811,N_8968);
nor U9123 (N_9123,N_8946,N_8842);
nand U9124 (N_9124,N_8979,N_8877);
nor U9125 (N_9125,N_8856,N_8861);
nand U9126 (N_9126,N_8962,N_8895);
and U9127 (N_9127,N_8819,N_8849);
nor U9128 (N_9128,N_8963,N_8998);
or U9129 (N_9129,N_8992,N_8915);
or U9130 (N_9130,N_8874,N_8855);
nand U9131 (N_9131,N_8933,N_8956);
or U9132 (N_9132,N_8924,N_8922);
nor U9133 (N_9133,N_8889,N_8864);
xnor U9134 (N_9134,N_8966,N_8986);
and U9135 (N_9135,N_8897,N_8862);
or U9136 (N_9136,N_8851,N_8945);
nand U9137 (N_9137,N_8993,N_8978);
or U9138 (N_9138,N_8992,N_8908);
xor U9139 (N_9139,N_8881,N_8802);
nor U9140 (N_9140,N_8850,N_8931);
nor U9141 (N_9141,N_8946,N_8989);
nor U9142 (N_9142,N_8951,N_8969);
or U9143 (N_9143,N_8811,N_8985);
nand U9144 (N_9144,N_8891,N_8955);
and U9145 (N_9145,N_8906,N_8921);
nand U9146 (N_9146,N_8944,N_8925);
or U9147 (N_9147,N_8932,N_8802);
or U9148 (N_9148,N_8804,N_8965);
or U9149 (N_9149,N_8967,N_8831);
nand U9150 (N_9150,N_8895,N_8873);
or U9151 (N_9151,N_8935,N_8962);
or U9152 (N_9152,N_8945,N_8890);
or U9153 (N_9153,N_8920,N_8835);
xnor U9154 (N_9154,N_8870,N_8830);
or U9155 (N_9155,N_8987,N_8862);
or U9156 (N_9156,N_8858,N_8933);
nand U9157 (N_9157,N_8948,N_8983);
or U9158 (N_9158,N_8839,N_8965);
and U9159 (N_9159,N_8989,N_8963);
and U9160 (N_9160,N_8832,N_8963);
nand U9161 (N_9161,N_8883,N_8871);
nor U9162 (N_9162,N_8907,N_8978);
and U9163 (N_9163,N_8900,N_8953);
nand U9164 (N_9164,N_8931,N_8944);
or U9165 (N_9165,N_8839,N_8920);
or U9166 (N_9166,N_8834,N_8839);
and U9167 (N_9167,N_8880,N_8915);
nand U9168 (N_9168,N_8980,N_8813);
nor U9169 (N_9169,N_8942,N_8945);
nor U9170 (N_9170,N_8910,N_8876);
nand U9171 (N_9171,N_8951,N_8913);
or U9172 (N_9172,N_8984,N_8956);
nand U9173 (N_9173,N_8988,N_8842);
or U9174 (N_9174,N_8964,N_8880);
nor U9175 (N_9175,N_8931,N_8858);
or U9176 (N_9176,N_8999,N_8892);
nand U9177 (N_9177,N_8992,N_8926);
or U9178 (N_9178,N_8841,N_8951);
nor U9179 (N_9179,N_8905,N_8909);
and U9180 (N_9180,N_8988,N_8898);
and U9181 (N_9181,N_8955,N_8828);
nor U9182 (N_9182,N_8909,N_8806);
and U9183 (N_9183,N_8887,N_8810);
or U9184 (N_9184,N_8850,N_8858);
and U9185 (N_9185,N_8928,N_8819);
or U9186 (N_9186,N_8876,N_8850);
and U9187 (N_9187,N_8998,N_8839);
nor U9188 (N_9188,N_8831,N_8943);
and U9189 (N_9189,N_8803,N_8842);
nand U9190 (N_9190,N_8966,N_8907);
or U9191 (N_9191,N_8925,N_8856);
nand U9192 (N_9192,N_8810,N_8865);
or U9193 (N_9193,N_8949,N_8860);
nor U9194 (N_9194,N_8958,N_8867);
nand U9195 (N_9195,N_8802,N_8991);
nand U9196 (N_9196,N_8997,N_8856);
nand U9197 (N_9197,N_8875,N_8872);
nor U9198 (N_9198,N_8900,N_8838);
and U9199 (N_9199,N_8988,N_8814);
nor U9200 (N_9200,N_9145,N_9038);
or U9201 (N_9201,N_9045,N_9049);
nand U9202 (N_9202,N_9101,N_9099);
nor U9203 (N_9203,N_9081,N_9040);
and U9204 (N_9204,N_9136,N_9021);
nand U9205 (N_9205,N_9139,N_9193);
nand U9206 (N_9206,N_9025,N_9152);
and U9207 (N_9207,N_9134,N_9196);
nand U9208 (N_9208,N_9010,N_9148);
nand U9209 (N_9209,N_9110,N_9030);
or U9210 (N_9210,N_9187,N_9020);
and U9211 (N_9211,N_9022,N_9177);
nand U9212 (N_9212,N_9032,N_9009);
or U9213 (N_9213,N_9113,N_9090);
nor U9214 (N_9214,N_9005,N_9097);
or U9215 (N_9215,N_9056,N_9012);
nor U9216 (N_9216,N_9072,N_9117);
or U9217 (N_9217,N_9067,N_9132);
nand U9218 (N_9218,N_9190,N_9141);
or U9219 (N_9219,N_9183,N_9195);
and U9220 (N_9220,N_9171,N_9131);
or U9221 (N_9221,N_9035,N_9100);
nor U9222 (N_9222,N_9052,N_9173);
nor U9223 (N_9223,N_9167,N_9017);
nand U9224 (N_9224,N_9197,N_9087);
nor U9225 (N_9225,N_9170,N_9163);
or U9226 (N_9226,N_9119,N_9156);
nand U9227 (N_9227,N_9175,N_9103);
nand U9228 (N_9228,N_9165,N_9000);
or U9229 (N_9229,N_9188,N_9065);
and U9230 (N_9230,N_9185,N_9064);
nor U9231 (N_9231,N_9184,N_9044);
and U9232 (N_9232,N_9161,N_9077);
or U9233 (N_9233,N_9003,N_9172);
nor U9234 (N_9234,N_9026,N_9125);
nor U9235 (N_9235,N_9155,N_9169);
or U9236 (N_9236,N_9106,N_9143);
nor U9237 (N_9237,N_9055,N_9133);
or U9238 (N_9238,N_9191,N_9098);
nand U9239 (N_9239,N_9094,N_9023);
or U9240 (N_9240,N_9138,N_9014);
nor U9241 (N_9241,N_9118,N_9011);
nor U9242 (N_9242,N_9123,N_9179);
nand U9243 (N_9243,N_9178,N_9150);
nand U9244 (N_9244,N_9089,N_9018);
nor U9245 (N_9245,N_9114,N_9047);
xor U9246 (N_9246,N_9007,N_9120);
or U9247 (N_9247,N_9181,N_9121);
nor U9248 (N_9248,N_9192,N_9015);
nand U9249 (N_9249,N_9080,N_9037);
nor U9250 (N_9250,N_9084,N_9111);
and U9251 (N_9251,N_9053,N_9043);
or U9252 (N_9252,N_9137,N_9095);
nor U9253 (N_9253,N_9008,N_9069);
nor U9254 (N_9254,N_9142,N_9158);
nand U9255 (N_9255,N_9058,N_9042);
nand U9256 (N_9256,N_9186,N_9063);
and U9257 (N_9257,N_9078,N_9149);
nor U9258 (N_9258,N_9130,N_9024);
or U9259 (N_9259,N_9092,N_9076);
and U9260 (N_9260,N_9088,N_9073);
or U9261 (N_9261,N_9066,N_9093);
nand U9262 (N_9262,N_9168,N_9105);
nor U9263 (N_9263,N_9109,N_9027);
and U9264 (N_9264,N_9129,N_9016);
nand U9265 (N_9265,N_9002,N_9050);
and U9266 (N_9266,N_9061,N_9147);
nand U9267 (N_9267,N_9194,N_9198);
and U9268 (N_9268,N_9199,N_9128);
and U9269 (N_9269,N_9075,N_9001);
and U9270 (N_9270,N_9104,N_9115);
and U9271 (N_9271,N_9126,N_9127);
nand U9272 (N_9272,N_9096,N_9028);
or U9273 (N_9273,N_9059,N_9144);
nand U9274 (N_9274,N_9057,N_9102);
nand U9275 (N_9275,N_9176,N_9160);
xor U9276 (N_9276,N_9082,N_9054);
nor U9277 (N_9277,N_9085,N_9029);
and U9278 (N_9278,N_9004,N_9180);
nand U9279 (N_9279,N_9070,N_9046);
and U9280 (N_9280,N_9039,N_9013);
and U9281 (N_9281,N_9033,N_9135);
and U9282 (N_9282,N_9051,N_9157);
and U9283 (N_9283,N_9034,N_9112);
and U9284 (N_9284,N_9124,N_9060);
and U9285 (N_9285,N_9108,N_9182);
or U9286 (N_9286,N_9159,N_9174);
xor U9287 (N_9287,N_9086,N_9122);
or U9288 (N_9288,N_9079,N_9041);
or U9289 (N_9289,N_9006,N_9151);
nor U9290 (N_9290,N_9074,N_9031);
nand U9291 (N_9291,N_9116,N_9107);
and U9292 (N_9292,N_9154,N_9189);
nand U9293 (N_9293,N_9166,N_9062);
and U9294 (N_9294,N_9068,N_9146);
and U9295 (N_9295,N_9164,N_9036);
or U9296 (N_9296,N_9153,N_9083);
or U9297 (N_9297,N_9162,N_9048);
or U9298 (N_9298,N_9091,N_9019);
nand U9299 (N_9299,N_9140,N_9071);
nor U9300 (N_9300,N_9050,N_9172);
or U9301 (N_9301,N_9050,N_9182);
nor U9302 (N_9302,N_9079,N_9110);
and U9303 (N_9303,N_9109,N_9107);
nor U9304 (N_9304,N_9001,N_9194);
and U9305 (N_9305,N_9148,N_9017);
and U9306 (N_9306,N_9190,N_9169);
and U9307 (N_9307,N_9094,N_9138);
nor U9308 (N_9308,N_9020,N_9024);
nand U9309 (N_9309,N_9185,N_9157);
nand U9310 (N_9310,N_9179,N_9158);
or U9311 (N_9311,N_9006,N_9094);
or U9312 (N_9312,N_9019,N_9016);
and U9313 (N_9313,N_9144,N_9102);
nand U9314 (N_9314,N_9126,N_9088);
nand U9315 (N_9315,N_9086,N_9013);
nand U9316 (N_9316,N_9174,N_9091);
nand U9317 (N_9317,N_9007,N_9182);
nand U9318 (N_9318,N_9129,N_9149);
nand U9319 (N_9319,N_9157,N_9011);
nand U9320 (N_9320,N_9180,N_9143);
nor U9321 (N_9321,N_9043,N_9122);
nand U9322 (N_9322,N_9010,N_9026);
and U9323 (N_9323,N_9030,N_9073);
nor U9324 (N_9324,N_9096,N_9159);
nand U9325 (N_9325,N_9165,N_9063);
or U9326 (N_9326,N_9163,N_9124);
or U9327 (N_9327,N_9021,N_9119);
and U9328 (N_9328,N_9034,N_9170);
nand U9329 (N_9329,N_9008,N_9190);
nor U9330 (N_9330,N_9127,N_9130);
nand U9331 (N_9331,N_9101,N_9102);
or U9332 (N_9332,N_9138,N_9130);
and U9333 (N_9333,N_9181,N_9177);
or U9334 (N_9334,N_9062,N_9054);
or U9335 (N_9335,N_9071,N_9109);
or U9336 (N_9336,N_9038,N_9027);
and U9337 (N_9337,N_9132,N_9051);
or U9338 (N_9338,N_9110,N_9037);
and U9339 (N_9339,N_9098,N_9037);
or U9340 (N_9340,N_9073,N_9070);
nor U9341 (N_9341,N_9024,N_9070);
and U9342 (N_9342,N_9056,N_9172);
or U9343 (N_9343,N_9021,N_9025);
nand U9344 (N_9344,N_9088,N_9033);
nand U9345 (N_9345,N_9052,N_9101);
nor U9346 (N_9346,N_9134,N_9072);
nand U9347 (N_9347,N_9019,N_9151);
nand U9348 (N_9348,N_9008,N_9136);
nor U9349 (N_9349,N_9163,N_9067);
nor U9350 (N_9350,N_9192,N_9194);
and U9351 (N_9351,N_9022,N_9025);
nand U9352 (N_9352,N_9002,N_9176);
and U9353 (N_9353,N_9085,N_9030);
nand U9354 (N_9354,N_9152,N_9195);
nor U9355 (N_9355,N_9010,N_9104);
xnor U9356 (N_9356,N_9030,N_9170);
or U9357 (N_9357,N_9125,N_9160);
nor U9358 (N_9358,N_9067,N_9085);
nand U9359 (N_9359,N_9192,N_9172);
nand U9360 (N_9360,N_9093,N_9114);
and U9361 (N_9361,N_9145,N_9124);
nor U9362 (N_9362,N_9193,N_9168);
xnor U9363 (N_9363,N_9055,N_9094);
or U9364 (N_9364,N_9082,N_9145);
nand U9365 (N_9365,N_9125,N_9176);
nand U9366 (N_9366,N_9057,N_9014);
and U9367 (N_9367,N_9156,N_9007);
or U9368 (N_9368,N_9041,N_9046);
nand U9369 (N_9369,N_9062,N_9120);
nand U9370 (N_9370,N_9153,N_9114);
and U9371 (N_9371,N_9088,N_9110);
xnor U9372 (N_9372,N_9089,N_9034);
nor U9373 (N_9373,N_9164,N_9075);
and U9374 (N_9374,N_9110,N_9180);
nor U9375 (N_9375,N_9008,N_9092);
nor U9376 (N_9376,N_9177,N_9103);
nor U9377 (N_9377,N_9195,N_9176);
and U9378 (N_9378,N_9123,N_9051);
and U9379 (N_9379,N_9112,N_9092);
nor U9380 (N_9380,N_9037,N_9009);
nor U9381 (N_9381,N_9104,N_9047);
and U9382 (N_9382,N_9166,N_9026);
nor U9383 (N_9383,N_9146,N_9042);
xor U9384 (N_9384,N_9167,N_9126);
nor U9385 (N_9385,N_9173,N_9050);
nand U9386 (N_9386,N_9175,N_9196);
nand U9387 (N_9387,N_9135,N_9024);
nor U9388 (N_9388,N_9113,N_9083);
and U9389 (N_9389,N_9062,N_9004);
nand U9390 (N_9390,N_9191,N_9102);
or U9391 (N_9391,N_9114,N_9052);
nor U9392 (N_9392,N_9053,N_9054);
nand U9393 (N_9393,N_9092,N_9074);
xor U9394 (N_9394,N_9143,N_9035);
and U9395 (N_9395,N_9071,N_9105);
and U9396 (N_9396,N_9053,N_9000);
nor U9397 (N_9397,N_9130,N_9143);
or U9398 (N_9398,N_9133,N_9168);
nand U9399 (N_9399,N_9155,N_9127);
nor U9400 (N_9400,N_9294,N_9398);
nand U9401 (N_9401,N_9222,N_9220);
and U9402 (N_9402,N_9373,N_9314);
and U9403 (N_9403,N_9315,N_9282);
or U9404 (N_9404,N_9232,N_9321);
and U9405 (N_9405,N_9208,N_9370);
nand U9406 (N_9406,N_9359,N_9387);
and U9407 (N_9407,N_9317,N_9245);
nand U9408 (N_9408,N_9356,N_9345);
and U9409 (N_9409,N_9286,N_9348);
and U9410 (N_9410,N_9312,N_9216);
nor U9411 (N_9411,N_9349,N_9293);
nor U9412 (N_9412,N_9327,N_9251);
nor U9413 (N_9413,N_9334,N_9207);
nand U9414 (N_9414,N_9297,N_9254);
and U9415 (N_9415,N_9238,N_9290);
nand U9416 (N_9416,N_9304,N_9278);
and U9417 (N_9417,N_9385,N_9380);
nand U9418 (N_9418,N_9206,N_9397);
nor U9419 (N_9419,N_9256,N_9341);
nand U9420 (N_9420,N_9376,N_9319);
nand U9421 (N_9421,N_9227,N_9284);
nor U9422 (N_9422,N_9234,N_9242);
and U9423 (N_9423,N_9332,N_9263);
nor U9424 (N_9424,N_9275,N_9323);
nor U9425 (N_9425,N_9379,N_9338);
and U9426 (N_9426,N_9382,N_9210);
nor U9427 (N_9427,N_9330,N_9392);
nor U9428 (N_9428,N_9240,N_9307);
nor U9429 (N_9429,N_9374,N_9299);
and U9430 (N_9430,N_9257,N_9394);
or U9431 (N_9431,N_9368,N_9311);
and U9432 (N_9432,N_9389,N_9364);
xnor U9433 (N_9433,N_9260,N_9252);
nor U9434 (N_9434,N_9288,N_9310);
nand U9435 (N_9435,N_9289,N_9237);
or U9436 (N_9436,N_9270,N_9276);
and U9437 (N_9437,N_9246,N_9331);
nor U9438 (N_9438,N_9262,N_9201);
or U9439 (N_9439,N_9233,N_9375);
and U9440 (N_9440,N_9365,N_9213);
and U9441 (N_9441,N_9243,N_9280);
or U9442 (N_9442,N_9378,N_9308);
and U9443 (N_9443,N_9306,N_9265);
or U9444 (N_9444,N_9325,N_9274);
or U9445 (N_9445,N_9360,N_9381);
and U9446 (N_9446,N_9230,N_9247);
nand U9447 (N_9447,N_9258,N_9393);
or U9448 (N_9448,N_9309,N_9287);
nand U9449 (N_9449,N_9209,N_9384);
nor U9450 (N_9450,N_9253,N_9200);
nor U9451 (N_9451,N_9295,N_9204);
nor U9452 (N_9452,N_9283,N_9215);
or U9453 (N_9453,N_9322,N_9344);
or U9454 (N_9454,N_9313,N_9231);
and U9455 (N_9455,N_9221,N_9371);
nor U9456 (N_9456,N_9250,N_9343);
nand U9457 (N_9457,N_9214,N_9386);
or U9458 (N_9458,N_9390,N_9355);
nor U9459 (N_9459,N_9303,N_9369);
nand U9460 (N_9460,N_9347,N_9277);
nor U9461 (N_9461,N_9346,N_9249);
or U9462 (N_9462,N_9320,N_9268);
nor U9463 (N_9463,N_9261,N_9357);
or U9464 (N_9464,N_9372,N_9267);
nand U9465 (N_9465,N_9302,N_9285);
nand U9466 (N_9466,N_9351,N_9329);
xor U9467 (N_9467,N_9391,N_9211);
or U9468 (N_9468,N_9363,N_9395);
nor U9469 (N_9469,N_9361,N_9342);
nand U9470 (N_9470,N_9273,N_9255);
and U9471 (N_9471,N_9305,N_9383);
nor U9472 (N_9472,N_9229,N_9248);
or U9473 (N_9473,N_9236,N_9203);
and U9474 (N_9474,N_9358,N_9228);
and U9475 (N_9475,N_9367,N_9225);
nand U9476 (N_9476,N_9339,N_9350);
or U9477 (N_9477,N_9366,N_9354);
nand U9478 (N_9478,N_9281,N_9336);
or U9479 (N_9479,N_9396,N_9388);
or U9480 (N_9480,N_9296,N_9340);
or U9481 (N_9481,N_9352,N_9266);
or U9482 (N_9482,N_9300,N_9205);
nor U9483 (N_9483,N_9218,N_9241);
and U9484 (N_9484,N_9292,N_9272);
and U9485 (N_9485,N_9337,N_9316);
nor U9486 (N_9486,N_9271,N_9326);
and U9487 (N_9487,N_9377,N_9333);
or U9488 (N_9488,N_9224,N_9235);
nand U9489 (N_9489,N_9202,N_9362);
or U9490 (N_9490,N_9328,N_9324);
nand U9491 (N_9491,N_9279,N_9335);
nand U9492 (N_9492,N_9212,N_9217);
nand U9493 (N_9493,N_9226,N_9244);
or U9494 (N_9494,N_9269,N_9223);
nor U9495 (N_9495,N_9291,N_9318);
or U9496 (N_9496,N_9259,N_9301);
nand U9497 (N_9497,N_9298,N_9399);
nand U9498 (N_9498,N_9353,N_9239);
or U9499 (N_9499,N_9264,N_9219);
or U9500 (N_9500,N_9314,N_9384);
xnor U9501 (N_9501,N_9346,N_9356);
or U9502 (N_9502,N_9379,N_9311);
nor U9503 (N_9503,N_9307,N_9294);
and U9504 (N_9504,N_9225,N_9355);
or U9505 (N_9505,N_9317,N_9371);
nand U9506 (N_9506,N_9335,N_9336);
nand U9507 (N_9507,N_9386,N_9218);
and U9508 (N_9508,N_9278,N_9336);
or U9509 (N_9509,N_9276,N_9332);
nor U9510 (N_9510,N_9215,N_9394);
nand U9511 (N_9511,N_9363,N_9200);
nand U9512 (N_9512,N_9382,N_9262);
nor U9513 (N_9513,N_9355,N_9327);
xor U9514 (N_9514,N_9271,N_9361);
or U9515 (N_9515,N_9257,N_9341);
and U9516 (N_9516,N_9264,N_9276);
and U9517 (N_9517,N_9360,N_9391);
nand U9518 (N_9518,N_9329,N_9299);
nand U9519 (N_9519,N_9347,N_9359);
xor U9520 (N_9520,N_9322,N_9310);
nand U9521 (N_9521,N_9258,N_9368);
or U9522 (N_9522,N_9241,N_9393);
and U9523 (N_9523,N_9344,N_9348);
and U9524 (N_9524,N_9339,N_9363);
and U9525 (N_9525,N_9237,N_9292);
and U9526 (N_9526,N_9363,N_9336);
nor U9527 (N_9527,N_9331,N_9205);
nand U9528 (N_9528,N_9253,N_9212);
or U9529 (N_9529,N_9254,N_9273);
nor U9530 (N_9530,N_9266,N_9294);
nand U9531 (N_9531,N_9301,N_9374);
nand U9532 (N_9532,N_9342,N_9277);
nand U9533 (N_9533,N_9255,N_9301);
and U9534 (N_9534,N_9367,N_9248);
nand U9535 (N_9535,N_9370,N_9336);
or U9536 (N_9536,N_9312,N_9330);
and U9537 (N_9537,N_9201,N_9270);
nand U9538 (N_9538,N_9340,N_9245);
nor U9539 (N_9539,N_9363,N_9399);
or U9540 (N_9540,N_9308,N_9270);
nor U9541 (N_9541,N_9383,N_9281);
or U9542 (N_9542,N_9281,N_9355);
or U9543 (N_9543,N_9337,N_9213);
and U9544 (N_9544,N_9212,N_9329);
and U9545 (N_9545,N_9263,N_9334);
nor U9546 (N_9546,N_9360,N_9367);
nand U9547 (N_9547,N_9253,N_9226);
nand U9548 (N_9548,N_9347,N_9257);
nand U9549 (N_9549,N_9308,N_9282);
and U9550 (N_9550,N_9377,N_9237);
nand U9551 (N_9551,N_9362,N_9262);
nand U9552 (N_9552,N_9210,N_9394);
nand U9553 (N_9553,N_9356,N_9387);
nor U9554 (N_9554,N_9338,N_9294);
nand U9555 (N_9555,N_9387,N_9342);
or U9556 (N_9556,N_9275,N_9290);
and U9557 (N_9557,N_9250,N_9336);
nor U9558 (N_9558,N_9235,N_9334);
and U9559 (N_9559,N_9368,N_9215);
and U9560 (N_9560,N_9228,N_9260);
nor U9561 (N_9561,N_9370,N_9381);
xnor U9562 (N_9562,N_9301,N_9235);
xor U9563 (N_9563,N_9320,N_9228);
or U9564 (N_9564,N_9241,N_9317);
nor U9565 (N_9565,N_9278,N_9321);
nand U9566 (N_9566,N_9238,N_9227);
nand U9567 (N_9567,N_9280,N_9246);
nor U9568 (N_9568,N_9367,N_9372);
nor U9569 (N_9569,N_9357,N_9241);
or U9570 (N_9570,N_9254,N_9315);
and U9571 (N_9571,N_9300,N_9332);
nand U9572 (N_9572,N_9315,N_9224);
or U9573 (N_9573,N_9223,N_9216);
nor U9574 (N_9574,N_9349,N_9232);
nor U9575 (N_9575,N_9210,N_9327);
xnor U9576 (N_9576,N_9277,N_9380);
nor U9577 (N_9577,N_9241,N_9219);
nor U9578 (N_9578,N_9297,N_9267);
nor U9579 (N_9579,N_9285,N_9332);
nand U9580 (N_9580,N_9247,N_9212);
and U9581 (N_9581,N_9261,N_9398);
nand U9582 (N_9582,N_9240,N_9248);
nand U9583 (N_9583,N_9231,N_9371);
and U9584 (N_9584,N_9225,N_9325);
nand U9585 (N_9585,N_9322,N_9319);
nand U9586 (N_9586,N_9208,N_9271);
and U9587 (N_9587,N_9257,N_9250);
nor U9588 (N_9588,N_9230,N_9223);
nand U9589 (N_9589,N_9320,N_9235);
and U9590 (N_9590,N_9257,N_9264);
nor U9591 (N_9591,N_9376,N_9346);
nand U9592 (N_9592,N_9357,N_9385);
and U9593 (N_9593,N_9295,N_9378);
nand U9594 (N_9594,N_9222,N_9329);
nor U9595 (N_9595,N_9204,N_9376);
and U9596 (N_9596,N_9390,N_9209);
and U9597 (N_9597,N_9224,N_9258);
nand U9598 (N_9598,N_9288,N_9298);
and U9599 (N_9599,N_9245,N_9227);
and U9600 (N_9600,N_9427,N_9408);
nand U9601 (N_9601,N_9453,N_9403);
nand U9602 (N_9602,N_9588,N_9545);
and U9603 (N_9603,N_9401,N_9548);
or U9604 (N_9604,N_9552,N_9535);
and U9605 (N_9605,N_9565,N_9541);
or U9606 (N_9606,N_9508,N_9580);
and U9607 (N_9607,N_9446,N_9435);
and U9608 (N_9608,N_9564,N_9524);
nor U9609 (N_9609,N_9411,N_9512);
or U9610 (N_9610,N_9533,N_9520);
or U9611 (N_9611,N_9470,N_9450);
and U9612 (N_9612,N_9546,N_9417);
nor U9613 (N_9613,N_9487,N_9581);
and U9614 (N_9614,N_9591,N_9424);
nand U9615 (N_9615,N_9447,N_9542);
or U9616 (N_9616,N_9493,N_9439);
nand U9617 (N_9617,N_9437,N_9418);
nand U9618 (N_9618,N_9404,N_9509);
nor U9619 (N_9619,N_9505,N_9454);
nand U9620 (N_9620,N_9534,N_9544);
or U9621 (N_9621,N_9459,N_9400);
and U9622 (N_9622,N_9444,N_9563);
nand U9623 (N_9623,N_9500,N_9557);
nand U9624 (N_9624,N_9472,N_9519);
nand U9625 (N_9625,N_9516,N_9525);
nor U9626 (N_9626,N_9539,N_9592);
and U9627 (N_9627,N_9443,N_9458);
nand U9628 (N_9628,N_9478,N_9589);
or U9629 (N_9629,N_9419,N_9596);
and U9630 (N_9630,N_9477,N_9497);
nand U9631 (N_9631,N_9407,N_9576);
or U9632 (N_9632,N_9464,N_9573);
xnor U9633 (N_9633,N_9568,N_9415);
or U9634 (N_9634,N_9503,N_9599);
nand U9635 (N_9635,N_9468,N_9521);
or U9636 (N_9636,N_9507,N_9584);
nor U9637 (N_9637,N_9562,N_9440);
nor U9638 (N_9638,N_9558,N_9593);
nand U9639 (N_9639,N_9486,N_9597);
and U9640 (N_9640,N_9550,N_9441);
and U9641 (N_9641,N_9528,N_9587);
nand U9642 (N_9642,N_9531,N_9574);
nor U9643 (N_9643,N_9577,N_9506);
and U9644 (N_9644,N_9554,N_9504);
nor U9645 (N_9645,N_9479,N_9549);
or U9646 (N_9646,N_9526,N_9421);
or U9647 (N_9647,N_9551,N_9571);
or U9648 (N_9648,N_9514,N_9469);
nand U9649 (N_9649,N_9585,N_9536);
nand U9650 (N_9650,N_9572,N_9561);
xnor U9651 (N_9651,N_9569,N_9511);
nand U9652 (N_9652,N_9537,N_9476);
nor U9653 (N_9653,N_9583,N_9434);
or U9654 (N_9654,N_9595,N_9433);
nor U9655 (N_9655,N_9490,N_9452);
nor U9656 (N_9656,N_9465,N_9513);
nor U9657 (N_9657,N_9494,N_9501);
nand U9658 (N_9658,N_9466,N_9455);
and U9659 (N_9659,N_9429,N_9474);
or U9660 (N_9660,N_9567,N_9570);
and U9661 (N_9661,N_9560,N_9538);
nand U9662 (N_9662,N_9532,N_9559);
nand U9663 (N_9663,N_9405,N_9436);
nor U9664 (N_9664,N_9423,N_9522);
nand U9665 (N_9665,N_9518,N_9484);
nor U9666 (N_9666,N_9471,N_9547);
nand U9667 (N_9667,N_9412,N_9461);
nand U9668 (N_9668,N_9496,N_9566);
and U9669 (N_9669,N_9426,N_9523);
or U9670 (N_9670,N_9438,N_9579);
nand U9671 (N_9671,N_9556,N_9515);
or U9672 (N_9672,N_9488,N_9481);
nand U9673 (N_9673,N_9492,N_9463);
or U9674 (N_9674,N_9510,N_9406);
nor U9675 (N_9675,N_9430,N_9485);
or U9676 (N_9676,N_9594,N_9451);
nand U9677 (N_9677,N_9530,N_9482);
and U9678 (N_9678,N_9483,N_9491);
or U9679 (N_9679,N_9457,N_9499);
or U9680 (N_9680,N_9428,N_9460);
nor U9681 (N_9681,N_9420,N_9527);
nor U9682 (N_9682,N_9432,N_9475);
and U9683 (N_9683,N_9467,N_9489);
nand U9684 (N_9684,N_9582,N_9578);
nand U9685 (N_9685,N_9456,N_9473);
and U9686 (N_9686,N_9495,N_9555);
nor U9687 (N_9687,N_9529,N_9431);
nor U9688 (N_9688,N_9517,N_9553);
and U9689 (N_9689,N_9449,N_9586);
nand U9690 (N_9690,N_9413,N_9575);
or U9691 (N_9691,N_9402,N_9498);
nand U9692 (N_9692,N_9409,N_9425);
and U9693 (N_9693,N_9442,N_9543);
or U9694 (N_9694,N_9462,N_9540);
nand U9695 (N_9695,N_9445,N_9416);
and U9696 (N_9696,N_9598,N_9422);
and U9697 (N_9697,N_9448,N_9410);
or U9698 (N_9698,N_9414,N_9590);
and U9699 (N_9699,N_9480,N_9502);
nor U9700 (N_9700,N_9476,N_9459);
or U9701 (N_9701,N_9447,N_9424);
nand U9702 (N_9702,N_9592,N_9436);
and U9703 (N_9703,N_9533,N_9456);
nand U9704 (N_9704,N_9466,N_9596);
or U9705 (N_9705,N_9539,N_9443);
and U9706 (N_9706,N_9516,N_9520);
and U9707 (N_9707,N_9456,N_9416);
and U9708 (N_9708,N_9439,N_9575);
or U9709 (N_9709,N_9495,N_9419);
and U9710 (N_9710,N_9475,N_9520);
nand U9711 (N_9711,N_9422,N_9414);
and U9712 (N_9712,N_9514,N_9429);
and U9713 (N_9713,N_9452,N_9480);
nand U9714 (N_9714,N_9503,N_9546);
and U9715 (N_9715,N_9508,N_9465);
nand U9716 (N_9716,N_9465,N_9569);
or U9717 (N_9717,N_9433,N_9417);
nand U9718 (N_9718,N_9481,N_9495);
or U9719 (N_9719,N_9502,N_9416);
nand U9720 (N_9720,N_9581,N_9594);
nand U9721 (N_9721,N_9568,N_9477);
nor U9722 (N_9722,N_9447,N_9531);
or U9723 (N_9723,N_9429,N_9540);
or U9724 (N_9724,N_9577,N_9412);
nor U9725 (N_9725,N_9519,N_9543);
and U9726 (N_9726,N_9466,N_9584);
and U9727 (N_9727,N_9418,N_9431);
nor U9728 (N_9728,N_9553,N_9447);
or U9729 (N_9729,N_9489,N_9492);
nand U9730 (N_9730,N_9575,N_9598);
and U9731 (N_9731,N_9599,N_9548);
nor U9732 (N_9732,N_9560,N_9580);
nor U9733 (N_9733,N_9483,N_9439);
and U9734 (N_9734,N_9543,N_9516);
nor U9735 (N_9735,N_9569,N_9563);
nor U9736 (N_9736,N_9405,N_9404);
nor U9737 (N_9737,N_9445,N_9471);
or U9738 (N_9738,N_9560,N_9483);
and U9739 (N_9739,N_9498,N_9454);
nand U9740 (N_9740,N_9574,N_9543);
and U9741 (N_9741,N_9567,N_9582);
nand U9742 (N_9742,N_9512,N_9469);
or U9743 (N_9743,N_9404,N_9431);
and U9744 (N_9744,N_9501,N_9469);
or U9745 (N_9745,N_9494,N_9495);
and U9746 (N_9746,N_9518,N_9412);
nand U9747 (N_9747,N_9553,N_9485);
nand U9748 (N_9748,N_9406,N_9558);
nor U9749 (N_9749,N_9491,N_9572);
or U9750 (N_9750,N_9461,N_9515);
and U9751 (N_9751,N_9416,N_9585);
or U9752 (N_9752,N_9550,N_9443);
nor U9753 (N_9753,N_9585,N_9519);
nand U9754 (N_9754,N_9533,N_9450);
or U9755 (N_9755,N_9481,N_9466);
nor U9756 (N_9756,N_9534,N_9513);
nand U9757 (N_9757,N_9476,N_9506);
nand U9758 (N_9758,N_9542,N_9562);
or U9759 (N_9759,N_9541,N_9475);
nand U9760 (N_9760,N_9471,N_9489);
nor U9761 (N_9761,N_9536,N_9582);
or U9762 (N_9762,N_9557,N_9424);
nand U9763 (N_9763,N_9468,N_9462);
nor U9764 (N_9764,N_9508,N_9563);
and U9765 (N_9765,N_9444,N_9560);
nand U9766 (N_9766,N_9493,N_9457);
nor U9767 (N_9767,N_9527,N_9498);
nor U9768 (N_9768,N_9495,N_9590);
nand U9769 (N_9769,N_9479,N_9570);
xnor U9770 (N_9770,N_9509,N_9497);
nor U9771 (N_9771,N_9466,N_9527);
nand U9772 (N_9772,N_9426,N_9538);
nor U9773 (N_9773,N_9541,N_9496);
nand U9774 (N_9774,N_9423,N_9460);
and U9775 (N_9775,N_9539,N_9489);
nand U9776 (N_9776,N_9558,N_9408);
and U9777 (N_9777,N_9482,N_9526);
nor U9778 (N_9778,N_9491,N_9432);
nor U9779 (N_9779,N_9598,N_9408);
and U9780 (N_9780,N_9568,N_9485);
nor U9781 (N_9781,N_9409,N_9489);
nand U9782 (N_9782,N_9427,N_9465);
nor U9783 (N_9783,N_9597,N_9535);
or U9784 (N_9784,N_9469,N_9549);
nor U9785 (N_9785,N_9597,N_9488);
nor U9786 (N_9786,N_9525,N_9532);
nand U9787 (N_9787,N_9431,N_9540);
nand U9788 (N_9788,N_9446,N_9419);
or U9789 (N_9789,N_9513,N_9529);
or U9790 (N_9790,N_9499,N_9430);
or U9791 (N_9791,N_9508,N_9499);
and U9792 (N_9792,N_9420,N_9490);
nand U9793 (N_9793,N_9456,N_9516);
nor U9794 (N_9794,N_9514,N_9585);
nor U9795 (N_9795,N_9592,N_9484);
nor U9796 (N_9796,N_9456,N_9565);
or U9797 (N_9797,N_9435,N_9545);
and U9798 (N_9798,N_9556,N_9577);
and U9799 (N_9799,N_9562,N_9494);
or U9800 (N_9800,N_9612,N_9687);
nor U9801 (N_9801,N_9792,N_9636);
or U9802 (N_9802,N_9775,N_9610);
nor U9803 (N_9803,N_9797,N_9694);
and U9804 (N_9804,N_9691,N_9648);
nand U9805 (N_9805,N_9733,N_9679);
and U9806 (N_9806,N_9712,N_9731);
and U9807 (N_9807,N_9601,N_9608);
and U9808 (N_9808,N_9696,N_9647);
or U9809 (N_9809,N_9642,N_9618);
nor U9810 (N_9810,N_9690,N_9663);
nand U9811 (N_9811,N_9695,N_9665);
or U9812 (N_9812,N_9768,N_9613);
or U9813 (N_9813,N_9641,N_9660);
and U9814 (N_9814,N_9614,N_9686);
or U9815 (N_9815,N_9786,N_9796);
and U9816 (N_9816,N_9734,N_9682);
and U9817 (N_9817,N_9701,N_9623);
and U9818 (N_9818,N_9709,N_9729);
and U9819 (N_9819,N_9738,N_9782);
and U9820 (N_9820,N_9619,N_9727);
nand U9821 (N_9821,N_9671,N_9676);
or U9822 (N_9822,N_9788,N_9675);
or U9823 (N_9823,N_9726,N_9674);
and U9824 (N_9824,N_9749,N_9684);
or U9825 (N_9825,N_9743,N_9718);
or U9826 (N_9826,N_9627,N_9669);
nand U9827 (N_9827,N_9774,N_9736);
nor U9828 (N_9828,N_9715,N_9628);
and U9829 (N_9829,N_9781,N_9748);
or U9830 (N_9830,N_9711,N_9760);
nor U9831 (N_9831,N_9725,N_9794);
or U9832 (N_9832,N_9629,N_9741);
or U9833 (N_9833,N_9672,N_9637);
or U9834 (N_9834,N_9755,N_9777);
and U9835 (N_9835,N_9615,N_9710);
and U9836 (N_9836,N_9763,N_9606);
and U9837 (N_9837,N_9773,N_9721);
nand U9838 (N_9838,N_9708,N_9722);
and U9839 (N_9839,N_9693,N_9752);
xor U9840 (N_9840,N_9659,N_9759);
or U9841 (N_9841,N_9699,N_9651);
nand U9842 (N_9842,N_9724,N_9622);
nand U9843 (N_9843,N_9621,N_9657);
or U9844 (N_9844,N_9717,N_9704);
nor U9845 (N_9845,N_9791,N_9634);
nor U9846 (N_9846,N_9790,N_9680);
nand U9847 (N_9847,N_9626,N_9624);
nor U9848 (N_9848,N_9751,N_9631);
or U9849 (N_9849,N_9678,N_9728);
and U9850 (N_9850,N_9661,N_9716);
nor U9851 (N_9851,N_9744,N_9778);
or U9852 (N_9852,N_9700,N_9737);
nand U9853 (N_9853,N_9654,N_9772);
nor U9854 (N_9854,N_9666,N_9756);
or U9855 (N_9855,N_9799,N_9653);
nand U9856 (N_9856,N_9732,N_9625);
and U9857 (N_9857,N_9767,N_9633);
or U9858 (N_9858,N_9713,N_9750);
nor U9859 (N_9859,N_9753,N_9706);
or U9860 (N_9860,N_9698,N_9643);
nor U9861 (N_9861,N_9662,N_9673);
and U9862 (N_9862,N_9692,N_9705);
and U9863 (N_9863,N_9620,N_9635);
or U9864 (N_9864,N_9783,N_9605);
or U9865 (N_9865,N_9658,N_9764);
and U9866 (N_9866,N_9779,N_9639);
or U9867 (N_9867,N_9603,N_9638);
nor U9868 (N_9868,N_9681,N_9747);
nand U9869 (N_9869,N_9688,N_9604);
nand U9870 (N_9870,N_9702,N_9632);
xnor U9871 (N_9871,N_9703,N_9739);
nor U9872 (N_9872,N_9668,N_9766);
nor U9873 (N_9873,N_9609,N_9785);
and U9874 (N_9874,N_9611,N_9630);
and U9875 (N_9875,N_9765,N_9670);
or U9876 (N_9876,N_9697,N_9602);
and U9877 (N_9877,N_9740,N_9607);
nand U9878 (N_9878,N_9650,N_9689);
nor U9879 (N_9879,N_9600,N_9616);
nand U9880 (N_9880,N_9719,N_9769);
and U9881 (N_9881,N_9746,N_9758);
or U9882 (N_9882,N_9655,N_9664);
or U9883 (N_9883,N_9720,N_9714);
nand U9884 (N_9884,N_9735,N_9780);
nand U9885 (N_9885,N_9645,N_9730);
nand U9886 (N_9886,N_9644,N_9770);
nor U9887 (N_9887,N_9795,N_9617);
nand U9888 (N_9888,N_9667,N_9656);
nor U9889 (N_9889,N_9640,N_9776);
xor U9890 (N_9890,N_9793,N_9784);
nor U9891 (N_9891,N_9754,N_9652);
or U9892 (N_9892,N_9745,N_9798);
and U9893 (N_9893,N_9762,N_9757);
nand U9894 (N_9894,N_9789,N_9683);
or U9895 (N_9895,N_9649,N_9761);
xnor U9896 (N_9896,N_9771,N_9707);
and U9897 (N_9897,N_9742,N_9723);
nand U9898 (N_9898,N_9646,N_9677);
and U9899 (N_9899,N_9685,N_9787);
or U9900 (N_9900,N_9694,N_9764);
and U9901 (N_9901,N_9699,N_9659);
or U9902 (N_9902,N_9779,N_9791);
nor U9903 (N_9903,N_9782,N_9699);
nand U9904 (N_9904,N_9790,N_9725);
or U9905 (N_9905,N_9644,N_9716);
nand U9906 (N_9906,N_9726,N_9666);
or U9907 (N_9907,N_9708,N_9682);
and U9908 (N_9908,N_9752,N_9751);
nand U9909 (N_9909,N_9731,N_9747);
nand U9910 (N_9910,N_9607,N_9616);
nand U9911 (N_9911,N_9628,N_9730);
or U9912 (N_9912,N_9700,N_9719);
nand U9913 (N_9913,N_9782,N_9600);
and U9914 (N_9914,N_9718,N_9714);
and U9915 (N_9915,N_9654,N_9727);
nand U9916 (N_9916,N_9747,N_9655);
or U9917 (N_9917,N_9745,N_9797);
nand U9918 (N_9918,N_9786,N_9637);
or U9919 (N_9919,N_9688,N_9783);
nor U9920 (N_9920,N_9759,N_9771);
nor U9921 (N_9921,N_9636,N_9618);
and U9922 (N_9922,N_9629,N_9603);
and U9923 (N_9923,N_9766,N_9640);
nor U9924 (N_9924,N_9703,N_9602);
and U9925 (N_9925,N_9635,N_9712);
nand U9926 (N_9926,N_9654,N_9780);
nor U9927 (N_9927,N_9691,N_9658);
nor U9928 (N_9928,N_9603,N_9730);
and U9929 (N_9929,N_9768,N_9621);
nand U9930 (N_9930,N_9768,N_9763);
nand U9931 (N_9931,N_9773,N_9795);
or U9932 (N_9932,N_9677,N_9658);
or U9933 (N_9933,N_9653,N_9795);
nand U9934 (N_9934,N_9784,N_9627);
or U9935 (N_9935,N_9724,N_9717);
nor U9936 (N_9936,N_9639,N_9629);
nor U9937 (N_9937,N_9780,N_9604);
and U9938 (N_9938,N_9764,N_9668);
and U9939 (N_9939,N_9795,N_9606);
or U9940 (N_9940,N_9736,N_9675);
and U9941 (N_9941,N_9612,N_9614);
or U9942 (N_9942,N_9667,N_9621);
nor U9943 (N_9943,N_9601,N_9640);
nor U9944 (N_9944,N_9715,N_9663);
nor U9945 (N_9945,N_9750,N_9669);
and U9946 (N_9946,N_9786,N_9622);
and U9947 (N_9947,N_9704,N_9649);
or U9948 (N_9948,N_9631,N_9795);
nor U9949 (N_9949,N_9673,N_9601);
nor U9950 (N_9950,N_9735,N_9688);
and U9951 (N_9951,N_9775,N_9685);
or U9952 (N_9952,N_9698,N_9616);
and U9953 (N_9953,N_9678,N_9744);
nor U9954 (N_9954,N_9741,N_9731);
nand U9955 (N_9955,N_9627,N_9750);
and U9956 (N_9956,N_9754,N_9713);
and U9957 (N_9957,N_9601,N_9686);
nand U9958 (N_9958,N_9708,N_9678);
nor U9959 (N_9959,N_9764,N_9659);
nand U9960 (N_9960,N_9670,N_9749);
or U9961 (N_9961,N_9731,N_9636);
or U9962 (N_9962,N_9636,N_9611);
nor U9963 (N_9963,N_9696,N_9616);
and U9964 (N_9964,N_9616,N_9651);
nand U9965 (N_9965,N_9666,N_9702);
or U9966 (N_9966,N_9601,N_9688);
and U9967 (N_9967,N_9627,N_9609);
and U9968 (N_9968,N_9628,N_9603);
nor U9969 (N_9969,N_9683,N_9741);
nand U9970 (N_9970,N_9770,N_9642);
or U9971 (N_9971,N_9623,N_9705);
and U9972 (N_9972,N_9622,N_9694);
and U9973 (N_9973,N_9715,N_9664);
and U9974 (N_9974,N_9719,N_9690);
or U9975 (N_9975,N_9731,N_9766);
xnor U9976 (N_9976,N_9643,N_9770);
nand U9977 (N_9977,N_9651,N_9691);
nand U9978 (N_9978,N_9786,N_9696);
or U9979 (N_9979,N_9733,N_9741);
or U9980 (N_9980,N_9657,N_9617);
and U9981 (N_9981,N_9629,N_9790);
or U9982 (N_9982,N_9773,N_9779);
nand U9983 (N_9983,N_9603,N_9733);
nand U9984 (N_9984,N_9757,N_9743);
nor U9985 (N_9985,N_9677,N_9634);
nand U9986 (N_9986,N_9741,N_9781);
and U9987 (N_9987,N_9691,N_9789);
nand U9988 (N_9988,N_9689,N_9687);
or U9989 (N_9989,N_9605,N_9769);
nand U9990 (N_9990,N_9793,N_9758);
and U9991 (N_9991,N_9634,N_9705);
nand U9992 (N_9992,N_9721,N_9729);
nand U9993 (N_9993,N_9653,N_9678);
nor U9994 (N_9994,N_9668,N_9648);
or U9995 (N_9995,N_9626,N_9731);
nor U9996 (N_9996,N_9760,N_9734);
nor U9997 (N_9997,N_9719,N_9612);
or U9998 (N_9998,N_9757,N_9707);
nor U9999 (N_9999,N_9728,N_9786);
and UO_0 (O_0,N_9815,N_9951);
xor UO_1 (O_1,N_9976,N_9995);
and UO_2 (O_2,N_9836,N_9828);
nand UO_3 (O_3,N_9873,N_9946);
and UO_4 (O_4,N_9997,N_9880);
xor UO_5 (O_5,N_9914,N_9849);
or UO_6 (O_6,N_9904,N_9970);
or UO_7 (O_7,N_9982,N_9850);
and UO_8 (O_8,N_9906,N_9994);
and UO_9 (O_9,N_9800,N_9972);
or UO_10 (O_10,N_9943,N_9838);
and UO_11 (O_11,N_9882,N_9969);
or UO_12 (O_12,N_9813,N_9931);
or UO_13 (O_13,N_9826,N_9909);
nor UO_14 (O_14,N_9876,N_9854);
or UO_15 (O_15,N_9855,N_9894);
or UO_16 (O_16,N_9934,N_9954);
nand UO_17 (O_17,N_9979,N_9936);
and UO_18 (O_18,N_9846,N_9991);
and UO_19 (O_19,N_9809,N_9806);
or UO_20 (O_20,N_9844,N_9958);
nor UO_21 (O_21,N_9928,N_9810);
or UO_22 (O_22,N_9864,N_9926);
nor UO_23 (O_23,N_9948,N_9912);
nor UO_24 (O_24,N_9861,N_9808);
nor UO_25 (O_25,N_9987,N_9992);
and UO_26 (O_26,N_9811,N_9922);
nor UO_27 (O_27,N_9971,N_9973);
nand UO_28 (O_28,N_9801,N_9899);
nand UO_29 (O_29,N_9887,N_9860);
and UO_30 (O_30,N_9897,N_9890);
nand UO_31 (O_31,N_9974,N_9905);
and UO_32 (O_32,N_9888,N_9817);
nand UO_33 (O_33,N_9881,N_9956);
and UO_34 (O_34,N_9919,N_9960);
and UO_35 (O_35,N_9869,N_9944);
and UO_36 (O_36,N_9925,N_9840);
nand UO_37 (O_37,N_9959,N_9862);
nor UO_38 (O_38,N_9940,N_9927);
and UO_39 (O_39,N_9975,N_9879);
nor UO_40 (O_40,N_9865,N_9872);
nor UO_41 (O_41,N_9984,N_9834);
or UO_42 (O_42,N_9823,N_9859);
or UO_43 (O_43,N_9981,N_9939);
nor UO_44 (O_44,N_9896,N_9805);
nand UO_45 (O_45,N_9961,N_9918);
nand UO_46 (O_46,N_9833,N_9977);
or UO_47 (O_47,N_9884,N_9952);
nor UO_48 (O_48,N_9938,N_9988);
or UO_49 (O_49,N_9907,N_9929);
or UO_50 (O_50,N_9875,N_9820);
nor UO_51 (O_51,N_9845,N_9878);
and UO_52 (O_52,N_9967,N_9920);
nor UO_53 (O_53,N_9804,N_9924);
nor UO_54 (O_54,N_9963,N_9807);
nor UO_55 (O_55,N_9910,N_9932);
nand UO_56 (O_56,N_9812,N_9983);
xor UO_57 (O_57,N_9978,N_9852);
nand UO_58 (O_58,N_9841,N_9893);
nor UO_59 (O_59,N_9930,N_9892);
nor UO_60 (O_60,N_9913,N_9911);
nand UO_61 (O_61,N_9824,N_9993);
or UO_62 (O_62,N_9903,N_9877);
nor UO_63 (O_63,N_9957,N_9945);
nor UO_64 (O_64,N_9863,N_9830);
xnor UO_65 (O_65,N_9821,N_9853);
nor UO_66 (O_66,N_9898,N_9868);
and UO_67 (O_67,N_9842,N_9871);
nand UO_68 (O_68,N_9949,N_9942);
or UO_69 (O_69,N_9858,N_9816);
and UO_70 (O_70,N_9999,N_9870);
and UO_71 (O_71,N_9856,N_9902);
or UO_72 (O_72,N_9802,N_9891);
nor UO_73 (O_73,N_9851,N_9953);
nand UO_74 (O_74,N_9990,N_9966);
nor UO_75 (O_75,N_9921,N_9827);
nor UO_76 (O_76,N_9829,N_9916);
and UO_77 (O_77,N_9835,N_9883);
nor UO_78 (O_78,N_9937,N_9915);
or UO_79 (O_79,N_9825,N_9989);
nor UO_80 (O_80,N_9814,N_9822);
or UO_81 (O_81,N_9941,N_9950);
nand UO_82 (O_82,N_9962,N_9908);
and UO_83 (O_83,N_9980,N_9947);
nand UO_84 (O_84,N_9839,N_9933);
xor UO_85 (O_85,N_9857,N_9843);
and UO_86 (O_86,N_9923,N_9831);
nor UO_87 (O_87,N_9889,N_9886);
and UO_88 (O_88,N_9885,N_9985);
nand UO_89 (O_89,N_9900,N_9819);
nand UO_90 (O_90,N_9818,N_9895);
or UO_91 (O_91,N_9955,N_9986);
nor UO_92 (O_92,N_9803,N_9901);
nand UO_93 (O_93,N_9866,N_9968);
or UO_94 (O_94,N_9998,N_9996);
nand UO_95 (O_95,N_9847,N_9935);
and UO_96 (O_96,N_9867,N_9848);
and UO_97 (O_97,N_9917,N_9874);
nor UO_98 (O_98,N_9964,N_9832);
nand UO_99 (O_99,N_9965,N_9837);
nand UO_100 (O_100,N_9914,N_9984);
nor UO_101 (O_101,N_9800,N_9999);
and UO_102 (O_102,N_9965,N_9961);
nor UO_103 (O_103,N_9993,N_9815);
or UO_104 (O_104,N_9945,N_9843);
or UO_105 (O_105,N_9962,N_9889);
nand UO_106 (O_106,N_9873,N_9824);
or UO_107 (O_107,N_9907,N_9935);
nor UO_108 (O_108,N_9941,N_9905);
nor UO_109 (O_109,N_9982,N_9967);
and UO_110 (O_110,N_9995,N_9862);
nor UO_111 (O_111,N_9996,N_9948);
xnor UO_112 (O_112,N_9862,N_9957);
nor UO_113 (O_113,N_9824,N_9958);
nor UO_114 (O_114,N_9862,N_9922);
and UO_115 (O_115,N_9805,N_9903);
and UO_116 (O_116,N_9924,N_9892);
and UO_117 (O_117,N_9890,N_9837);
nand UO_118 (O_118,N_9953,N_9952);
and UO_119 (O_119,N_9872,N_9903);
or UO_120 (O_120,N_9835,N_9828);
nand UO_121 (O_121,N_9818,N_9888);
nand UO_122 (O_122,N_9980,N_9808);
or UO_123 (O_123,N_9889,N_9815);
nor UO_124 (O_124,N_9994,N_9862);
and UO_125 (O_125,N_9810,N_9989);
nand UO_126 (O_126,N_9993,N_9957);
or UO_127 (O_127,N_9978,N_9877);
and UO_128 (O_128,N_9977,N_9880);
nand UO_129 (O_129,N_9820,N_9862);
or UO_130 (O_130,N_9885,N_9892);
or UO_131 (O_131,N_9803,N_9989);
nor UO_132 (O_132,N_9873,N_9871);
nand UO_133 (O_133,N_9930,N_9937);
nand UO_134 (O_134,N_9914,N_9890);
nor UO_135 (O_135,N_9867,N_9939);
or UO_136 (O_136,N_9957,N_9974);
nand UO_137 (O_137,N_9968,N_9816);
nor UO_138 (O_138,N_9935,N_9889);
nor UO_139 (O_139,N_9825,N_9940);
and UO_140 (O_140,N_9847,N_9984);
or UO_141 (O_141,N_9829,N_9967);
nand UO_142 (O_142,N_9941,N_9991);
nand UO_143 (O_143,N_9847,N_9943);
nand UO_144 (O_144,N_9861,N_9848);
nor UO_145 (O_145,N_9944,N_9949);
nor UO_146 (O_146,N_9991,N_9966);
and UO_147 (O_147,N_9927,N_9954);
xnor UO_148 (O_148,N_9893,N_9844);
nor UO_149 (O_149,N_9902,N_9849);
or UO_150 (O_150,N_9860,N_9835);
or UO_151 (O_151,N_9851,N_9954);
nor UO_152 (O_152,N_9973,N_9858);
or UO_153 (O_153,N_9882,N_9806);
or UO_154 (O_154,N_9937,N_9875);
and UO_155 (O_155,N_9838,N_9999);
nand UO_156 (O_156,N_9803,N_9948);
nor UO_157 (O_157,N_9823,N_9830);
or UO_158 (O_158,N_9812,N_9889);
xnor UO_159 (O_159,N_9824,N_9834);
or UO_160 (O_160,N_9948,N_9888);
nand UO_161 (O_161,N_9961,N_9868);
xor UO_162 (O_162,N_9966,N_9862);
nand UO_163 (O_163,N_9891,N_9922);
nand UO_164 (O_164,N_9831,N_9857);
or UO_165 (O_165,N_9942,N_9899);
or UO_166 (O_166,N_9865,N_9880);
and UO_167 (O_167,N_9820,N_9863);
and UO_168 (O_168,N_9990,N_9841);
or UO_169 (O_169,N_9880,N_9817);
nand UO_170 (O_170,N_9890,N_9980);
nand UO_171 (O_171,N_9803,N_9982);
nor UO_172 (O_172,N_9880,N_9915);
nand UO_173 (O_173,N_9905,N_9961);
and UO_174 (O_174,N_9974,N_9915);
or UO_175 (O_175,N_9950,N_9904);
or UO_176 (O_176,N_9810,N_9930);
nor UO_177 (O_177,N_9857,N_9919);
nor UO_178 (O_178,N_9849,N_9860);
nand UO_179 (O_179,N_9814,N_9859);
nor UO_180 (O_180,N_9837,N_9921);
nand UO_181 (O_181,N_9809,N_9922);
nand UO_182 (O_182,N_9959,N_9993);
nor UO_183 (O_183,N_9813,N_9875);
or UO_184 (O_184,N_9862,N_9945);
nand UO_185 (O_185,N_9969,N_9817);
nand UO_186 (O_186,N_9919,N_9980);
nor UO_187 (O_187,N_9892,N_9901);
and UO_188 (O_188,N_9804,N_9889);
nor UO_189 (O_189,N_9842,N_9880);
and UO_190 (O_190,N_9945,N_9877);
or UO_191 (O_191,N_9879,N_9991);
and UO_192 (O_192,N_9961,N_9848);
or UO_193 (O_193,N_9849,N_9819);
and UO_194 (O_194,N_9813,N_9854);
xnor UO_195 (O_195,N_9958,N_9965);
nand UO_196 (O_196,N_9960,N_9883);
nand UO_197 (O_197,N_9933,N_9823);
nand UO_198 (O_198,N_9910,N_9907);
or UO_199 (O_199,N_9905,N_9833);
or UO_200 (O_200,N_9891,N_9969);
and UO_201 (O_201,N_9897,N_9926);
nor UO_202 (O_202,N_9986,N_9821);
or UO_203 (O_203,N_9973,N_9918);
nor UO_204 (O_204,N_9997,N_9834);
and UO_205 (O_205,N_9837,N_9809);
nor UO_206 (O_206,N_9930,N_9875);
or UO_207 (O_207,N_9949,N_9977);
or UO_208 (O_208,N_9904,N_9808);
nor UO_209 (O_209,N_9872,N_9923);
nor UO_210 (O_210,N_9912,N_9856);
and UO_211 (O_211,N_9962,N_9927);
nor UO_212 (O_212,N_9997,N_9816);
or UO_213 (O_213,N_9971,N_9891);
nand UO_214 (O_214,N_9810,N_9905);
and UO_215 (O_215,N_9860,N_9905);
nand UO_216 (O_216,N_9875,N_9851);
nand UO_217 (O_217,N_9809,N_9820);
nand UO_218 (O_218,N_9836,N_9904);
or UO_219 (O_219,N_9827,N_9803);
and UO_220 (O_220,N_9894,N_9963);
nor UO_221 (O_221,N_9999,N_9848);
nor UO_222 (O_222,N_9813,N_9852);
nor UO_223 (O_223,N_9954,N_9979);
nand UO_224 (O_224,N_9982,N_9971);
nor UO_225 (O_225,N_9915,N_9990);
and UO_226 (O_226,N_9846,N_9830);
nand UO_227 (O_227,N_9934,N_9811);
and UO_228 (O_228,N_9804,N_9819);
or UO_229 (O_229,N_9924,N_9930);
and UO_230 (O_230,N_9820,N_9963);
nand UO_231 (O_231,N_9884,N_9957);
xnor UO_232 (O_232,N_9930,N_9910);
nor UO_233 (O_233,N_9992,N_9838);
or UO_234 (O_234,N_9911,N_9847);
and UO_235 (O_235,N_9885,N_9949);
nand UO_236 (O_236,N_9818,N_9900);
nand UO_237 (O_237,N_9835,N_9960);
nor UO_238 (O_238,N_9854,N_9945);
and UO_239 (O_239,N_9971,N_9821);
or UO_240 (O_240,N_9968,N_9817);
nor UO_241 (O_241,N_9937,N_9840);
nor UO_242 (O_242,N_9821,N_9894);
nor UO_243 (O_243,N_9949,N_9846);
nor UO_244 (O_244,N_9811,N_9821);
xor UO_245 (O_245,N_9967,N_9844);
or UO_246 (O_246,N_9830,N_9974);
nand UO_247 (O_247,N_9814,N_9804);
nor UO_248 (O_248,N_9898,N_9953);
and UO_249 (O_249,N_9981,N_9938);
nor UO_250 (O_250,N_9908,N_9864);
xor UO_251 (O_251,N_9886,N_9847);
or UO_252 (O_252,N_9827,N_9984);
or UO_253 (O_253,N_9811,N_9924);
xnor UO_254 (O_254,N_9971,N_9913);
nor UO_255 (O_255,N_9953,N_9838);
nor UO_256 (O_256,N_9924,N_9832);
nor UO_257 (O_257,N_9899,N_9863);
and UO_258 (O_258,N_9985,N_9976);
xor UO_259 (O_259,N_9960,N_9841);
or UO_260 (O_260,N_9846,N_9994);
nand UO_261 (O_261,N_9852,N_9985);
and UO_262 (O_262,N_9985,N_9804);
and UO_263 (O_263,N_9986,N_9914);
nand UO_264 (O_264,N_9952,N_9849);
nor UO_265 (O_265,N_9881,N_9992);
or UO_266 (O_266,N_9932,N_9859);
nand UO_267 (O_267,N_9870,N_9927);
or UO_268 (O_268,N_9891,N_9872);
or UO_269 (O_269,N_9839,N_9842);
and UO_270 (O_270,N_9951,N_9845);
or UO_271 (O_271,N_9952,N_9987);
and UO_272 (O_272,N_9956,N_9897);
nand UO_273 (O_273,N_9899,N_9814);
and UO_274 (O_274,N_9877,N_9813);
or UO_275 (O_275,N_9920,N_9844);
or UO_276 (O_276,N_9822,N_9908);
or UO_277 (O_277,N_9914,N_9944);
or UO_278 (O_278,N_9869,N_9835);
nor UO_279 (O_279,N_9921,N_9807);
or UO_280 (O_280,N_9913,N_9826);
nor UO_281 (O_281,N_9924,N_9870);
or UO_282 (O_282,N_9911,N_9925);
nor UO_283 (O_283,N_9856,N_9808);
or UO_284 (O_284,N_9955,N_9894);
and UO_285 (O_285,N_9912,N_9946);
or UO_286 (O_286,N_9837,N_9882);
and UO_287 (O_287,N_9915,N_9900);
and UO_288 (O_288,N_9907,N_9871);
nand UO_289 (O_289,N_9808,N_9990);
nor UO_290 (O_290,N_9994,N_9896);
nor UO_291 (O_291,N_9904,N_9819);
nand UO_292 (O_292,N_9850,N_9998);
nor UO_293 (O_293,N_9847,N_9975);
nor UO_294 (O_294,N_9815,N_9978);
nor UO_295 (O_295,N_9912,N_9873);
nor UO_296 (O_296,N_9949,N_9921);
nor UO_297 (O_297,N_9836,N_9883);
nor UO_298 (O_298,N_9904,N_9999);
nor UO_299 (O_299,N_9955,N_9962);
nand UO_300 (O_300,N_9913,N_9903);
nor UO_301 (O_301,N_9888,N_9901);
nor UO_302 (O_302,N_9810,N_9870);
nor UO_303 (O_303,N_9971,N_9938);
nor UO_304 (O_304,N_9957,N_9983);
nand UO_305 (O_305,N_9921,N_9897);
nor UO_306 (O_306,N_9879,N_9995);
and UO_307 (O_307,N_9805,N_9954);
or UO_308 (O_308,N_9959,N_9870);
nor UO_309 (O_309,N_9995,N_9892);
and UO_310 (O_310,N_9867,N_9841);
nand UO_311 (O_311,N_9836,N_9832);
nand UO_312 (O_312,N_9868,N_9949);
and UO_313 (O_313,N_9808,N_9988);
or UO_314 (O_314,N_9927,N_9894);
nor UO_315 (O_315,N_9918,N_9958);
or UO_316 (O_316,N_9995,N_9951);
nor UO_317 (O_317,N_9929,N_9998);
or UO_318 (O_318,N_9936,N_9900);
and UO_319 (O_319,N_9805,N_9905);
nand UO_320 (O_320,N_9843,N_9954);
or UO_321 (O_321,N_9945,N_9964);
and UO_322 (O_322,N_9932,N_9984);
or UO_323 (O_323,N_9848,N_9990);
nand UO_324 (O_324,N_9837,N_9845);
nor UO_325 (O_325,N_9839,N_9948);
nand UO_326 (O_326,N_9826,N_9811);
nand UO_327 (O_327,N_9991,N_9909);
nand UO_328 (O_328,N_9997,N_9961);
or UO_329 (O_329,N_9849,N_9969);
xnor UO_330 (O_330,N_9890,N_9954);
or UO_331 (O_331,N_9884,N_9979);
nand UO_332 (O_332,N_9816,N_9809);
or UO_333 (O_333,N_9991,N_9999);
nor UO_334 (O_334,N_9947,N_9895);
or UO_335 (O_335,N_9963,N_9844);
nand UO_336 (O_336,N_9862,N_9993);
nand UO_337 (O_337,N_9868,N_9843);
nor UO_338 (O_338,N_9880,N_9954);
and UO_339 (O_339,N_9938,N_9850);
nand UO_340 (O_340,N_9838,N_9991);
and UO_341 (O_341,N_9956,N_9958);
nor UO_342 (O_342,N_9895,N_9905);
nor UO_343 (O_343,N_9861,N_9805);
or UO_344 (O_344,N_9847,N_9928);
xor UO_345 (O_345,N_9920,N_9888);
and UO_346 (O_346,N_9835,N_9966);
or UO_347 (O_347,N_9946,N_9981);
xnor UO_348 (O_348,N_9822,N_9943);
nand UO_349 (O_349,N_9962,N_9963);
nor UO_350 (O_350,N_9934,N_9921);
nor UO_351 (O_351,N_9961,N_9914);
nor UO_352 (O_352,N_9909,N_9872);
and UO_353 (O_353,N_9913,N_9988);
nand UO_354 (O_354,N_9847,N_9858);
nand UO_355 (O_355,N_9804,N_9975);
nand UO_356 (O_356,N_9874,N_9994);
nor UO_357 (O_357,N_9884,N_9833);
nor UO_358 (O_358,N_9990,N_9912);
or UO_359 (O_359,N_9941,N_9958);
xor UO_360 (O_360,N_9917,N_9973);
and UO_361 (O_361,N_9981,N_9977);
nand UO_362 (O_362,N_9856,N_9847);
nor UO_363 (O_363,N_9869,N_9901);
nor UO_364 (O_364,N_9809,N_9848);
nor UO_365 (O_365,N_9930,N_9981);
or UO_366 (O_366,N_9976,N_9906);
nand UO_367 (O_367,N_9832,N_9850);
and UO_368 (O_368,N_9970,N_9987);
nor UO_369 (O_369,N_9955,N_9875);
nor UO_370 (O_370,N_9886,N_9942);
nor UO_371 (O_371,N_9951,N_9959);
nor UO_372 (O_372,N_9971,N_9978);
nand UO_373 (O_373,N_9991,N_9865);
and UO_374 (O_374,N_9909,N_9910);
nand UO_375 (O_375,N_9905,N_9925);
nor UO_376 (O_376,N_9842,N_9833);
nand UO_377 (O_377,N_9864,N_9893);
or UO_378 (O_378,N_9923,N_9827);
nand UO_379 (O_379,N_9821,N_9891);
nor UO_380 (O_380,N_9928,N_9949);
nand UO_381 (O_381,N_9902,N_9904);
and UO_382 (O_382,N_9997,N_9991);
nand UO_383 (O_383,N_9859,N_9868);
or UO_384 (O_384,N_9989,N_9929);
nor UO_385 (O_385,N_9864,N_9886);
and UO_386 (O_386,N_9958,N_9815);
and UO_387 (O_387,N_9927,N_9878);
nand UO_388 (O_388,N_9957,N_9817);
nand UO_389 (O_389,N_9807,N_9907);
nand UO_390 (O_390,N_9863,N_9894);
or UO_391 (O_391,N_9926,N_9975);
and UO_392 (O_392,N_9832,N_9993);
and UO_393 (O_393,N_9909,N_9883);
nand UO_394 (O_394,N_9927,N_9935);
or UO_395 (O_395,N_9838,N_9841);
nand UO_396 (O_396,N_9970,N_9912);
nor UO_397 (O_397,N_9809,N_9805);
nor UO_398 (O_398,N_9990,N_9868);
and UO_399 (O_399,N_9809,N_9985);
or UO_400 (O_400,N_9953,N_9802);
and UO_401 (O_401,N_9849,N_9927);
nand UO_402 (O_402,N_9886,N_9922);
and UO_403 (O_403,N_9915,N_9884);
and UO_404 (O_404,N_9871,N_9852);
nand UO_405 (O_405,N_9991,N_9978);
nor UO_406 (O_406,N_9915,N_9857);
nor UO_407 (O_407,N_9934,N_9998);
and UO_408 (O_408,N_9929,N_9873);
nand UO_409 (O_409,N_9858,N_9818);
xor UO_410 (O_410,N_9810,N_9836);
nand UO_411 (O_411,N_9912,N_9892);
and UO_412 (O_412,N_9992,N_9813);
or UO_413 (O_413,N_9983,N_9888);
nand UO_414 (O_414,N_9956,N_9948);
nand UO_415 (O_415,N_9950,N_9987);
nor UO_416 (O_416,N_9960,N_9980);
and UO_417 (O_417,N_9958,N_9922);
and UO_418 (O_418,N_9934,N_9924);
and UO_419 (O_419,N_9971,N_9844);
nand UO_420 (O_420,N_9965,N_9840);
and UO_421 (O_421,N_9954,N_9882);
nor UO_422 (O_422,N_9861,N_9954);
nor UO_423 (O_423,N_9871,N_9918);
or UO_424 (O_424,N_9965,N_9841);
nor UO_425 (O_425,N_9906,N_9850);
xnor UO_426 (O_426,N_9912,N_9919);
and UO_427 (O_427,N_9860,N_9926);
and UO_428 (O_428,N_9911,N_9805);
or UO_429 (O_429,N_9807,N_9895);
nor UO_430 (O_430,N_9995,N_9898);
nor UO_431 (O_431,N_9928,N_9975);
xnor UO_432 (O_432,N_9973,N_9809);
nor UO_433 (O_433,N_9943,N_9895);
nand UO_434 (O_434,N_9910,N_9938);
or UO_435 (O_435,N_9929,N_9843);
and UO_436 (O_436,N_9943,N_9913);
nor UO_437 (O_437,N_9948,N_9940);
nor UO_438 (O_438,N_9975,N_9905);
and UO_439 (O_439,N_9896,N_9821);
nand UO_440 (O_440,N_9804,N_9918);
or UO_441 (O_441,N_9947,N_9937);
nand UO_442 (O_442,N_9801,N_9850);
nor UO_443 (O_443,N_9992,N_9866);
nand UO_444 (O_444,N_9921,N_9998);
or UO_445 (O_445,N_9936,N_9912);
nor UO_446 (O_446,N_9868,N_9808);
nor UO_447 (O_447,N_9892,N_9988);
or UO_448 (O_448,N_9939,N_9936);
xnor UO_449 (O_449,N_9828,N_9897);
or UO_450 (O_450,N_9963,N_9990);
nor UO_451 (O_451,N_9892,N_9944);
xnor UO_452 (O_452,N_9835,N_9844);
nor UO_453 (O_453,N_9982,N_9880);
nor UO_454 (O_454,N_9806,N_9801);
nand UO_455 (O_455,N_9934,N_9863);
or UO_456 (O_456,N_9986,N_9872);
or UO_457 (O_457,N_9906,N_9833);
or UO_458 (O_458,N_9933,N_9927);
or UO_459 (O_459,N_9839,N_9941);
and UO_460 (O_460,N_9949,N_9833);
nor UO_461 (O_461,N_9940,N_9955);
or UO_462 (O_462,N_9855,N_9999);
nand UO_463 (O_463,N_9835,N_9980);
or UO_464 (O_464,N_9860,N_9985);
nor UO_465 (O_465,N_9872,N_9949);
and UO_466 (O_466,N_9877,N_9859);
or UO_467 (O_467,N_9980,N_9987);
nor UO_468 (O_468,N_9948,N_9876);
nand UO_469 (O_469,N_9983,N_9844);
or UO_470 (O_470,N_9866,N_9817);
nand UO_471 (O_471,N_9811,N_9810);
or UO_472 (O_472,N_9977,N_9901);
nor UO_473 (O_473,N_9865,N_9833);
nor UO_474 (O_474,N_9857,N_9852);
nand UO_475 (O_475,N_9865,N_9974);
or UO_476 (O_476,N_9827,N_9862);
nand UO_477 (O_477,N_9939,N_9884);
and UO_478 (O_478,N_9858,N_9900);
and UO_479 (O_479,N_9880,N_9862);
nand UO_480 (O_480,N_9858,N_9944);
nand UO_481 (O_481,N_9980,N_9868);
xnor UO_482 (O_482,N_9993,N_9855);
nand UO_483 (O_483,N_9852,N_9925);
or UO_484 (O_484,N_9898,N_9971);
and UO_485 (O_485,N_9920,N_9976);
or UO_486 (O_486,N_9837,N_9941);
nand UO_487 (O_487,N_9839,N_9814);
and UO_488 (O_488,N_9935,N_9894);
nor UO_489 (O_489,N_9938,N_9871);
and UO_490 (O_490,N_9865,N_9973);
and UO_491 (O_491,N_9806,N_9802);
nand UO_492 (O_492,N_9993,N_9891);
and UO_493 (O_493,N_9843,N_9836);
and UO_494 (O_494,N_9884,N_9875);
nand UO_495 (O_495,N_9864,N_9994);
and UO_496 (O_496,N_9880,N_9854);
nor UO_497 (O_497,N_9938,N_9806);
nand UO_498 (O_498,N_9864,N_9925);
nor UO_499 (O_499,N_9841,N_9921);
xor UO_500 (O_500,N_9861,N_9935);
or UO_501 (O_501,N_9809,N_9932);
nand UO_502 (O_502,N_9970,N_9881);
and UO_503 (O_503,N_9972,N_9965);
nand UO_504 (O_504,N_9987,N_9976);
nor UO_505 (O_505,N_9849,N_9984);
nor UO_506 (O_506,N_9956,N_9844);
or UO_507 (O_507,N_9986,N_9800);
and UO_508 (O_508,N_9932,N_9835);
or UO_509 (O_509,N_9921,N_9858);
or UO_510 (O_510,N_9981,N_9819);
and UO_511 (O_511,N_9865,N_9901);
nand UO_512 (O_512,N_9918,N_9954);
nor UO_513 (O_513,N_9836,N_9884);
and UO_514 (O_514,N_9849,N_9876);
nor UO_515 (O_515,N_9834,N_9961);
nor UO_516 (O_516,N_9995,N_9833);
nor UO_517 (O_517,N_9925,N_9942);
xnor UO_518 (O_518,N_9975,N_9992);
nor UO_519 (O_519,N_9924,N_9891);
nor UO_520 (O_520,N_9902,N_9888);
nand UO_521 (O_521,N_9967,N_9928);
nor UO_522 (O_522,N_9976,N_9813);
or UO_523 (O_523,N_9926,N_9939);
or UO_524 (O_524,N_9800,N_9838);
nor UO_525 (O_525,N_9917,N_9994);
nor UO_526 (O_526,N_9883,N_9868);
nor UO_527 (O_527,N_9872,N_9811);
nand UO_528 (O_528,N_9992,N_9921);
and UO_529 (O_529,N_9868,N_9872);
nor UO_530 (O_530,N_9869,N_9839);
or UO_531 (O_531,N_9826,N_9815);
or UO_532 (O_532,N_9809,N_9845);
and UO_533 (O_533,N_9894,N_9800);
nand UO_534 (O_534,N_9920,N_9953);
and UO_535 (O_535,N_9906,N_9889);
nand UO_536 (O_536,N_9858,N_9848);
nor UO_537 (O_537,N_9845,N_9938);
xor UO_538 (O_538,N_9846,N_9936);
or UO_539 (O_539,N_9978,N_9965);
nand UO_540 (O_540,N_9999,N_9805);
nand UO_541 (O_541,N_9888,N_9841);
or UO_542 (O_542,N_9953,N_9955);
nor UO_543 (O_543,N_9990,N_9911);
nand UO_544 (O_544,N_9950,N_9864);
nand UO_545 (O_545,N_9988,N_9915);
and UO_546 (O_546,N_9977,N_9808);
nand UO_547 (O_547,N_9950,N_9893);
nor UO_548 (O_548,N_9846,N_9857);
and UO_549 (O_549,N_9849,N_9936);
nor UO_550 (O_550,N_9975,N_9890);
and UO_551 (O_551,N_9809,N_9928);
nor UO_552 (O_552,N_9839,N_9962);
or UO_553 (O_553,N_9992,N_9935);
or UO_554 (O_554,N_9828,N_9842);
and UO_555 (O_555,N_9927,N_9934);
nand UO_556 (O_556,N_9897,N_9905);
nand UO_557 (O_557,N_9858,N_9831);
nand UO_558 (O_558,N_9999,N_9907);
nand UO_559 (O_559,N_9834,N_9833);
nand UO_560 (O_560,N_9835,N_9976);
and UO_561 (O_561,N_9857,N_9803);
nor UO_562 (O_562,N_9864,N_9960);
nor UO_563 (O_563,N_9843,N_9988);
or UO_564 (O_564,N_9856,N_9995);
nand UO_565 (O_565,N_9849,N_9967);
nand UO_566 (O_566,N_9988,N_9865);
and UO_567 (O_567,N_9815,N_9899);
or UO_568 (O_568,N_9858,N_9903);
or UO_569 (O_569,N_9877,N_9816);
nor UO_570 (O_570,N_9965,N_9823);
nor UO_571 (O_571,N_9862,N_9963);
xnor UO_572 (O_572,N_9802,N_9981);
or UO_573 (O_573,N_9979,N_9815);
nor UO_574 (O_574,N_9994,N_9949);
and UO_575 (O_575,N_9814,N_9853);
and UO_576 (O_576,N_9853,N_9935);
nor UO_577 (O_577,N_9962,N_9815);
nor UO_578 (O_578,N_9899,N_9983);
and UO_579 (O_579,N_9818,N_9873);
xnor UO_580 (O_580,N_9828,N_9996);
nand UO_581 (O_581,N_9901,N_9926);
nor UO_582 (O_582,N_9867,N_9958);
nand UO_583 (O_583,N_9930,N_9908);
or UO_584 (O_584,N_9874,N_9877);
or UO_585 (O_585,N_9814,N_9978);
and UO_586 (O_586,N_9861,N_9929);
and UO_587 (O_587,N_9946,N_9935);
nor UO_588 (O_588,N_9924,N_9833);
or UO_589 (O_589,N_9848,N_9869);
or UO_590 (O_590,N_9841,N_9830);
and UO_591 (O_591,N_9907,N_9909);
and UO_592 (O_592,N_9841,N_9832);
xnor UO_593 (O_593,N_9835,N_9878);
or UO_594 (O_594,N_9912,N_9929);
or UO_595 (O_595,N_9806,N_9934);
nor UO_596 (O_596,N_9949,N_9869);
nor UO_597 (O_597,N_9944,N_9956);
or UO_598 (O_598,N_9990,N_9962);
or UO_599 (O_599,N_9814,N_9826);
and UO_600 (O_600,N_9929,N_9961);
nand UO_601 (O_601,N_9843,N_9989);
nor UO_602 (O_602,N_9846,N_9952);
nor UO_603 (O_603,N_9934,N_9853);
or UO_604 (O_604,N_9907,N_9947);
nand UO_605 (O_605,N_9876,N_9992);
nand UO_606 (O_606,N_9927,N_9908);
or UO_607 (O_607,N_9945,N_9894);
and UO_608 (O_608,N_9914,N_9823);
or UO_609 (O_609,N_9829,N_9979);
nand UO_610 (O_610,N_9972,N_9924);
or UO_611 (O_611,N_9818,N_9979);
and UO_612 (O_612,N_9950,N_9927);
nand UO_613 (O_613,N_9802,N_9912);
and UO_614 (O_614,N_9809,N_9959);
nand UO_615 (O_615,N_9931,N_9901);
and UO_616 (O_616,N_9935,N_9822);
nand UO_617 (O_617,N_9993,N_9987);
and UO_618 (O_618,N_9928,N_9833);
nand UO_619 (O_619,N_9917,N_9859);
nor UO_620 (O_620,N_9936,N_9864);
nand UO_621 (O_621,N_9956,N_9834);
nand UO_622 (O_622,N_9952,N_9861);
or UO_623 (O_623,N_9934,N_9928);
nor UO_624 (O_624,N_9923,N_9919);
nor UO_625 (O_625,N_9818,N_9954);
and UO_626 (O_626,N_9944,N_9843);
and UO_627 (O_627,N_9874,N_9949);
nor UO_628 (O_628,N_9843,N_9948);
nor UO_629 (O_629,N_9962,N_9937);
nand UO_630 (O_630,N_9985,N_9891);
nand UO_631 (O_631,N_9853,N_9830);
nor UO_632 (O_632,N_9826,N_9898);
and UO_633 (O_633,N_9929,N_9801);
nand UO_634 (O_634,N_9812,N_9841);
nor UO_635 (O_635,N_9895,N_9872);
and UO_636 (O_636,N_9975,N_9996);
and UO_637 (O_637,N_9892,N_9877);
nand UO_638 (O_638,N_9943,N_9940);
and UO_639 (O_639,N_9948,N_9869);
nand UO_640 (O_640,N_9954,N_9959);
and UO_641 (O_641,N_9836,N_9805);
or UO_642 (O_642,N_9913,N_9802);
nand UO_643 (O_643,N_9950,N_9914);
xor UO_644 (O_644,N_9819,N_9844);
nor UO_645 (O_645,N_9804,N_9870);
nor UO_646 (O_646,N_9963,N_9913);
nor UO_647 (O_647,N_9915,N_9817);
xnor UO_648 (O_648,N_9904,N_9942);
nand UO_649 (O_649,N_9868,N_9979);
nor UO_650 (O_650,N_9920,N_9902);
nand UO_651 (O_651,N_9867,N_9901);
nor UO_652 (O_652,N_9944,N_9931);
or UO_653 (O_653,N_9955,N_9978);
or UO_654 (O_654,N_9895,N_9900);
or UO_655 (O_655,N_9964,N_9825);
or UO_656 (O_656,N_9871,N_9919);
nor UO_657 (O_657,N_9929,N_9958);
nand UO_658 (O_658,N_9835,N_9848);
nand UO_659 (O_659,N_9963,N_9930);
and UO_660 (O_660,N_9802,N_9840);
and UO_661 (O_661,N_9973,N_9902);
nand UO_662 (O_662,N_9946,N_9836);
or UO_663 (O_663,N_9819,N_9956);
and UO_664 (O_664,N_9972,N_9955);
nor UO_665 (O_665,N_9938,N_9830);
and UO_666 (O_666,N_9936,N_9960);
or UO_667 (O_667,N_9958,N_9972);
nand UO_668 (O_668,N_9864,N_9907);
and UO_669 (O_669,N_9914,N_9877);
and UO_670 (O_670,N_9939,N_9901);
nand UO_671 (O_671,N_9815,N_9956);
or UO_672 (O_672,N_9996,N_9856);
nand UO_673 (O_673,N_9822,N_9833);
nand UO_674 (O_674,N_9970,N_9908);
or UO_675 (O_675,N_9980,N_9992);
or UO_676 (O_676,N_9909,N_9853);
nor UO_677 (O_677,N_9941,N_9800);
and UO_678 (O_678,N_9839,N_9884);
xor UO_679 (O_679,N_9973,N_9985);
and UO_680 (O_680,N_9814,N_9842);
nand UO_681 (O_681,N_9896,N_9800);
and UO_682 (O_682,N_9892,N_9931);
nand UO_683 (O_683,N_9984,N_9898);
nor UO_684 (O_684,N_9940,N_9915);
and UO_685 (O_685,N_9918,N_9939);
nor UO_686 (O_686,N_9987,N_9945);
nor UO_687 (O_687,N_9883,N_9911);
nand UO_688 (O_688,N_9869,N_9956);
and UO_689 (O_689,N_9910,N_9860);
and UO_690 (O_690,N_9856,N_9878);
nand UO_691 (O_691,N_9828,N_9856);
nand UO_692 (O_692,N_9936,N_9859);
or UO_693 (O_693,N_9893,N_9908);
nor UO_694 (O_694,N_9809,N_9941);
nand UO_695 (O_695,N_9851,N_9929);
and UO_696 (O_696,N_9920,N_9968);
and UO_697 (O_697,N_9866,N_9924);
nor UO_698 (O_698,N_9913,N_9901);
nand UO_699 (O_699,N_9929,N_9879);
or UO_700 (O_700,N_9879,N_9923);
or UO_701 (O_701,N_9940,N_9899);
and UO_702 (O_702,N_9993,N_9894);
or UO_703 (O_703,N_9846,N_9931);
nor UO_704 (O_704,N_9820,N_9851);
nand UO_705 (O_705,N_9853,N_9833);
nand UO_706 (O_706,N_9874,N_9961);
nand UO_707 (O_707,N_9830,N_9918);
nand UO_708 (O_708,N_9806,N_9907);
nand UO_709 (O_709,N_9968,N_9880);
and UO_710 (O_710,N_9840,N_9899);
or UO_711 (O_711,N_9916,N_9875);
nor UO_712 (O_712,N_9922,N_9898);
xor UO_713 (O_713,N_9829,N_9923);
and UO_714 (O_714,N_9932,N_9836);
nor UO_715 (O_715,N_9820,N_9925);
nor UO_716 (O_716,N_9978,N_9824);
and UO_717 (O_717,N_9829,N_9886);
nor UO_718 (O_718,N_9922,N_9837);
or UO_719 (O_719,N_9848,N_9828);
nand UO_720 (O_720,N_9880,N_9929);
nand UO_721 (O_721,N_9940,N_9958);
or UO_722 (O_722,N_9902,N_9929);
nor UO_723 (O_723,N_9842,N_9931);
nor UO_724 (O_724,N_9865,N_9821);
or UO_725 (O_725,N_9899,N_9848);
or UO_726 (O_726,N_9801,N_9852);
and UO_727 (O_727,N_9956,N_9826);
and UO_728 (O_728,N_9972,N_9808);
nor UO_729 (O_729,N_9962,N_9924);
and UO_730 (O_730,N_9957,N_9848);
nor UO_731 (O_731,N_9901,N_9915);
nand UO_732 (O_732,N_9989,N_9913);
nor UO_733 (O_733,N_9947,N_9880);
nor UO_734 (O_734,N_9876,N_9902);
and UO_735 (O_735,N_9925,N_9822);
xnor UO_736 (O_736,N_9963,N_9980);
nor UO_737 (O_737,N_9860,N_9919);
nor UO_738 (O_738,N_9986,N_9888);
nor UO_739 (O_739,N_9989,N_9924);
and UO_740 (O_740,N_9960,N_9944);
and UO_741 (O_741,N_9944,N_9975);
nand UO_742 (O_742,N_9852,N_9835);
nor UO_743 (O_743,N_9853,N_9932);
nor UO_744 (O_744,N_9925,N_9998);
nor UO_745 (O_745,N_9910,N_9835);
nor UO_746 (O_746,N_9913,N_9812);
and UO_747 (O_747,N_9844,N_9884);
nand UO_748 (O_748,N_9911,N_9955);
nor UO_749 (O_749,N_9953,N_9948);
or UO_750 (O_750,N_9809,N_9961);
nor UO_751 (O_751,N_9818,N_9907);
nand UO_752 (O_752,N_9841,N_9991);
nor UO_753 (O_753,N_9939,N_9825);
nand UO_754 (O_754,N_9939,N_9995);
nand UO_755 (O_755,N_9884,N_9895);
and UO_756 (O_756,N_9922,N_9895);
and UO_757 (O_757,N_9943,N_9954);
or UO_758 (O_758,N_9841,N_9878);
and UO_759 (O_759,N_9853,N_9855);
and UO_760 (O_760,N_9811,N_9979);
and UO_761 (O_761,N_9982,N_9818);
nand UO_762 (O_762,N_9964,N_9907);
and UO_763 (O_763,N_9912,N_9915);
and UO_764 (O_764,N_9861,N_9976);
and UO_765 (O_765,N_9814,N_9996);
and UO_766 (O_766,N_9968,N_9898);
nor UO_767 (O_767,N_9868,N_9993);
nor UO_768 (O_768,N_9843,N_9862);
nand UO_769 (O_769,N_9947,N_9913);
or UO_770 (O_770,N_9941,N_9988);
nand UO_771 (O_771,N_9917,N_9883);
and UO_772 (O_772,N_9812,N_9884);
nor UO_773 (O_773,N_9877,N_9975);
or UO_774 (O_774,N_9909,N_9824);
or UO_775 (O_775,N_9931,N_9847);
or UO_776 (O_776,N_9918,N_9808);
nor UO_777 (O_777,N_9960,N_9837);
and UO_778 (O_778,N_9997,N_9933);
or UO_779 (O_779,N_9974,N_9939);
nor UO_780 (O_780,N_9879,N_9822);
and UO_781 (O_781,N_9949,N_9889);
and UO_782 (O_782,N_9893,N_9895);
nand UO_783 (O_783,N_9902,N_9928);
nand UO_784 (O_784,N_9802,N_9883);
and UO_785 (O_785,N_9810,N_9849);
or UO_786 (O_786,N_9921,N_9848);
nand UO_787 (O_787,N_9832,N_9847);
or UO_788 (O_788,N_9882,N_9824);
and UO_789 (O_789,N_9800,N_9815);
and UO_790 (O_790,N_9821,N_9854);
nor UO_791 (O_791,N_9855,N_9968);
and UO_792 (O_792,N_9938,N_9939);
and UO_793 (O_793,N_9884,N_9874);
and UO_794 (O_794,N_9801,N_9985);
or UO_795 (O_795,N_9836,N_9927);
nand UO_796 (O_796,N_9958,N_9899);
nand UO_797 (O_797,N_9959,N_9880);
xnor UO_798 (O_798,N_9921,N_9945);
nand UO_799 (O_799,N_9953,N_9907);
nor UO_800 (O_800,N_9949,N_9941);
or UO_801 (O_801,N_9959,N_9905);
nor UO_802 (O_802,N_9903,N_9841);
nor UO_803 (O_803,N_9842,N_9947);
and UO_804 (O_804,N_9818,N_9880);
and UO_805 (O_805,N_9803,N_9887);
nor UO_806 (O_806,N_9879,N_9934);
nand UO_807 (O_807,N_9962,N_9851);
nor UO_808 (O_808,N_9817,N_9951);
or UO_809 (O_809,N_9858,N_9862);
nor UO_810 (O_810,N_9965,N_9993);
and UO_811 (O_811,N_9898,N_9990);
nand UO_812 (O_812,N_9879,N_9830);
or UO_813 (O_813,N_9892,N_9896);
nand UO_814 (O_814,N_9992,N_9904);
or UO_815 (O_815,N_9839,N_9953);
or UO_816 (O_816,N_9971,N_9860);
nor UO_817 (O_817,N_9927,N_9994);
and UO_818 (O_818,N_9872,N_9975);
or UO_819 (O_819,N_9964,N_9864);
and UO_820 (O_820,N_9982,N_9957);
nand UO_821 (O_821,N_9931,N_9862);
nor UO_822 (O_822,N_9929,N_9825);
and UO_823 (O_823,N_9953,N_9888);
or UO_824 (O_824,N_9993,N_9954);
or UO_825 (O_825,N_9815,N_9808);
or UO_826 (O_826,N_9811,N_9997);
or UO_827 (O_827,N_9841,N_9882);
or UO_828 (O_828,N_9836,N_9980);
nand UO_829 (O_829,N_9895,N_9959);
nor UO_830 (O_830,N_9945,N_9913);
nand UO_831 (O_831,N_9974,N_9963);
and UO_832 (O_832,N_9935,N_9893);
or UO_833 (O_833,N_9945,N_9870);
nor UO_834 (O_834,N_9962,N_9857);
nor UO_835 (O_835,N_9964,N_9893);
or UO_836 (O_836,N_9890,N_9928);
nor UO_837 (O_837,N_9815,N_9989);
and UO_838 (O_838,N_9965,N_9800);
or UO_839 (O_839,N_9806,N_9980);
nand UO_840 (O_840,N_9870,N_9828);
and UO_841 (O_841,N_9946,N_9928);
nor UO_842 (O_842,N_9947,N_9958);
nand UO_843 (O_843,N_9809,N_9938);
and UO_844 (O_844,N_9910,N_9933);
nand UO_845 (O_845,N_9910,N_9916);
nand UO_846 (O_846,N_9820,N_9984);
and UO_847 (O_847,N_9807,N_9919);
or UO_848 (O_848,N_9980,N_9955);
and UO_849 (O_849,N_9966,N_9974);
or UO_850 (O_850,N_9888,N_9801);
nor UO_851 (O_851,N_9974,N_9962);
and UO_852 (O_852,N_9846,N_9805);
nand UO_853 (O_853,N_9869,N_9926);
or UO_854 (O_854,N_9975,N_9895);
and UO_855 (O_855,N_9938,N_9929);
and UO_856 (O_856,N_9929,N_9980);
or UO_857 (O_857,N_9858,N_9896);
or UO_858 (O_858,N_9885,N_9990);
or UO_859 (O_859,N_9859,N_9804);
nor UO_860 (O_860,N_9947,N_9915);
or UO_861 (O_861,N_9930,N_9934);
nor UO_862 (O_862,N_9863,N_9840);
nor UO_863 (O_863,N_9879,N_9961);
and UO_864 (O_864,N_9823,N_9957);
or UO_865 (O_865,N_9884,N_9811);
nor UO_866 (O_866,N_9948,N_9983);
or UO_867 (O_867,N_9833,N_9969);
nand UO_868 (O_868,N_9916,N_9893);
nor UO_869 (O_869,N_9889,N_9977);
nor UO_870 (O_870,N_9892,N_9937);
nand UO_871 (O_871,N_9835,N_9988);
nor UO_872 (O_872,N_9828,N_9909);
or UO_873 (O_873,N_9817,N_9814);
or UO_874 (O_874,N_9995,N_9930);
nor UO_875 (O_875,N_9951,N_9886);
nand UO_876 (O_876,N_9864,N_9824);
or UO_877 (O_877,N_9874,N_9950);
or UO_878 (O_878,N_9958,N_9862);
or UO_879 (O_879,N_9909,N_9829);
nand UO_880 (O_880,N_9891,N_9833);
and UO_881 (O_881,N_9966,N_9945);
nand UO_882 (O_882,N_9980,N_9990);
nor UO_883 (O_883,N_9959,N_9929);
and UO_884 (O_884,N_9834,N_9854);
or UO_885 (O_885,N_9969,N_9988);
xnor UO_886 (O_886,N_9802,N_9808);
and UO_887 (O_887,N_9995,N_9830);
nor UO_888 (O_888,N_9854,N_9810);
and UO_889 (O_889,N_9817,N_9872);
and UO_890 (O_890,N_9919,N_9990);
nand UO_891 (O_891,N_9800,N_9886);
xnor UO_892 (O_892,N_9887,N_9921);
and UO_893 (O_893,N_9973,N_9805);
nand UO_894 (O_894,N_9849,N_9922);
nand UO_895 (O_895,N_9869,N_9838);
or UO_896 (O_896,N_9927,N_9848);
nand UO_897 (O_897,N_9944,N_9875);
or UO_898 (O_898,N_9851,N_9857);
or UO_899 (O_899,N_9867,N_9998);
nor UO_900 (O_900,N_9983,N_9945);
or UO_901 (O_901,N_9825,N_9871);
or UO_902 (O_902,N_9935,N_9998);
and UO_903 (O_903,N_9891,N_9967);
nor UO_904 (O_904,N_9905,N_9915);
or UO_905 (O_905,N_9886,N_9822);
nand UO_906 (O_906,N_9988,N_9922);
nand UO_907 (O_907,N_9934,N_9877);
and UO_908 (O_908,N_9973,N_9907);
or UO_909 (O_909,N_9884,N_9860);
nor UO_910 (O_910,N_9947,N_9892);
xor UO_911 (O_911,N_9965,N_9944);
and UO_912 (O_912,N_9844,N_9842);
nand UO_913 (O_913,N_9863,N_9904);
and UO_914 (O_914,N_9997,N_9989);
nand UO_915 (O_915,N_9993,N_9827);
nor UO_916 (O_916,N_9975,N_9875);
nand UO_917 (O_917,N_9821,N_9824);
and UO_918 (O_918,N_9920,N_9850);
and UO_919 (O_919,N_9916,N_9982);
and UO_920 (O_920,N_9821,N_9875);
nor UO_921 (O_921,N_9889,N_9898);
nor UO_922 (O_922,N_9804,N_9945);
nand UO_923 (O_923,N_9922,N_9833);
or UO_924 (O_924,N_9841,N_9897);
and UO_925 (O_925,N_9966,N_9853);
nand UO_926 (O_926,N_9858,N_9828);
or UO_927 (O_927,N_9937,N_9925);
and UO_928 (O_928,N_9853,N_9878);
and UO_929 (O_929,N_9876,N_9817);
or UO_930 (O_930,N_9814,N_9868);
or UO_931 (O_931,N_9846,N_9954);
nand UO_932 (O_932,N_9883,N_9916);
nor UO_933 (O_933,N_9895,N_9913);
nor UO_934 (O_934,N_9914,N_9802);
nor UO_935 (O_935,N_9953,N_9962);
or UO_936 (O_936,N_9993,N_9882);
and UO_937 (O_937,N_9845,N_9958);
and UO_938 (O_938,N_9919,N_9916);
or UO_939 (O_939,N_9930,N_9876);
nor UO_940 (O_940,N_9803,N_9825);
xnor UO_941 (O_941,N_9805,N_9952);
and UO_942 (O_942,N_9831,N_9819);
and UO_943 (O_943,N_9951,N_9870);
or UO_944 (O_944,N_9847,N_9925);
nand UO_945 (O_945,N_9946,N_9809);
or UO_946 (O_946,N_9923,N_9873);
nand UO_947 (O_947,N_9955,N_9952);
or UO_948 (O_948,N_9804,N_9891);
and UO_949 (O_949,N_9946,N_9992);
nor UO_950 (O_950,N_9805,N_9942);
and UO_951 (O_951,N_9958,N_9928);
nor UO_952 (O_952,N_9865,N_9832);
nor UO_953 (O_953,N_9947,N_9935);
or UO_954 (O_954,N_9882,N_9913);
and UO_955 (O_955,N_9897,N_9886);
nor UO_956 (O_956,N_9810,N_9900);
and UO_957 (O_957,N_9874,N_9954);
nand UO_958 (O_958,N_9925,N_9967);
nand UO_959 (O_959,N_9950,N_9881);
or UO_960 (O_960,N_9890,N_9867);
nand UO_961 (O_961,N_9988,N_9897);
and UO_962 (O_962,N_9953,N_9980);
nor UO_963 (O_963,N_9862,N_9898);
and UO_964 (O_964,N_9885,N_9821);
nor UO_965 (O_965,N_9959,N_9974);
and UO_966 (O_966,N_9963,N_9970);
or UO_967 (O_967,N_9849,N_9847);
and UO_968 (O_968,N_9992,N_9909);
and UO_969 (O_969,N_9868,N_9829);
nand UO_970 (O_970,N_9897,N_9867);
nor UO_971 (O_971,N_9823,N_9921);
and UO_972 (O_972,N_9989,N_9922);
nand UO_973 (O_973,N_9909,N_9804);
or UO_974 (O_974,N_9999,N_9928);
xor UO_975 (O_975,N_9946,N_9993);
nor UO_976 (O_976,N_9985,N_9858);
and UO_977 (O_977,N_9946,N_9879);
nand UO_978 (O_978,N_9995,N_9907);
and UO_979 (O_979,N_9997,N_9883);
nor UO_980 (O_980,N_9873,N_9825);
and UO_981 (O_981,N_9879,N_9907);
nor UO_982 (O_982,N_9817,N_9950);
or UO_983 (O_983,N_9816,N_9987);
nor UO_984 (O_984,N_9972,N_9930);
or UO_985 (O_985,N_9991,N_9913);
nor UO_986 (O_986,N_9811,N_9818);
or UO_987 (O_987,N_9911,N_9996);
and UO_988 (O_988,N_9898,N_9815);
nor UO_989 (O_989,N_9861,N_9869);
nor UO_990 (O_990,N_9963,N_9999);
nor UO_991 (O_991,N_9834,N_9999);
nand UO_992 (O_992,N_9802,N_9816);
or UO_993 (O_993,N_9809,N_9919);
and UO_994 (O_994,N_9848,N_9806);
and UO_995 (O_995,N_9956,N_9804);
or UO_996 (O_996,N_9813,N_9941);
and UO_997 (O_997,N_9970,N_9988);
nor UO_998 (O_998,N_9980,N_9803);
nand UO_999 (O_999,N_9871,N_9940);
nor UO_1000 (O_1000,N_9914,N_9972);
nand UO_1001 (O_1001,N_9887,N_9964);
or UO_1002 (O_1002,N_9932,N_9904);
nand UO_1003 (O_1003,N_9845,N_9810);
nand UO_1004 (O_1004,N_9994,N_9866);
or UO_1005 (O_1005,N_9975,N_9823);
or UO_1006 (O_1006,N_9941,N_9919);
or UO_1007 (O_1007,N_9875,N_9908);
nor UO_1008 (O_1008,N_9876,N_9814);
nand UO_1009 (O_1009,N_9827,N_9864);
nor UO_1010 (O_1010,N_9880,N_9805);
or UO_1011 (O_1011,N_9947,N_9847);
and UO_1012 (O_1012,N_9892,N_9934);
and UO_1013 (O_1013,N_9827,N_9896);
nand UO_1014 (O_1014,N_9962,N_9920);
nor UO_1015 (O_1015,N_9838,N_9916);
and UO_1016 (O_1016,N_9991,N_9924);
nand UO_1017 (O_1017,N_9968,N_9970);
nand UO_1018 (O_1018,N_9853,N_9865);
nand UO_1019 (O_1019,N_9901,N_9982);
nand UO_1020 (O_1020,N_9888,N_9874);
nor UO_1021 (O_1021,N_9907,N_9882);
nand UO_1022 (O_1022,N_9881,N_9920);
nand UO_1023 (O_1023,N_9988,N_9997);
and UO_1024 (O_1024,N_9927,N_9963);
nor UO_1025 (O_1025,N_9826,N_9998);
and UO_1026 (O_1026,N_9882,N_9981);
nand UO_1027 (O_1027,N_9932,N_9911);
nor UO_1028 (O_1028,N_9931,N_9907);
or UO_1029 (O_1029,N_9814,N_9844);
or UO_1030 (O_1030,N_9940,N_9811);
nor UO_1031 (O_1031,N_9985,N_9926);
or UO_1032 (O_1032,N_9808,N_9862);
nor UO_1033 (O_1033,N_9969,N_9929);
and UO_1034 (O_1034,N_9924,N_9834);
and UO_1035 (O_1035,N_9926,N_9927);
and UO_1036 (O_1036,N_9893,N_9942);
and UO_1037 (O_1037,N_9845,N_9821);
and UO_1038 (O_1038,N_9861,N_9881);
and UO_1039 (O_1039,N_9963,N_9971);
nor UO_1040 (O_1040,N_9811,N_9854);
and UO_1041 (O_1041,N_9806,N_9954);
or UO_1042 (O_1042,N_9886,N_9987);
nand UO_1043 (O_1043,N_9818,N_9884);
nand UO_1044 (O_1044,N_9925,N_9952);
xnor UO_1045 (O_1045,N_9997,N_9945);
and UO_1046 (O_1046,N_9961,N_9902);
xor UO_1047 (O_1047,N_9816,N_9813);
xor UO_1048 (O_1048,N_9921,N_9970);
nor UO_1049 (O_1049,N_9841,N_9975);
nand UO_1050 (O_1050,N_9850,N_9954);
and UO_1051 (O_1051,N_9898,N_9974);
nand UO_1052 (O_1052,N_9866,N_9996);
nand UO_1053 (O_1053,N_9968,N_9913);
and UO_1054 (O_1054,N_9843,N_9899);
and UO_1055 (O_1055,N_9867,N_9926);
nor UO_1056 (O_1056,N_9816,N_9984);
nand UO_1057 (O_1057,N_9926,N_9934);
or UO_1058 (O_1058,N_9874,N_9835);
nor UO_1059 (O_1059,N_9823,N_9846);
and UO_1060 (O_1060,N_9829,N_9880);
nor UO_1061 (O_1061,N_9996,N_9961);
or UO_1062 (O_1062,N_9899,N_9873);
xor UO_1063 (O_1063,N_9934,N_9801);
or UO_1064 (O_1064,N_9847,N_9912);
and UO_1065 (O_1065,N_9937,N_9982);
nand UO_1066 (O_1066,N_9956,N_9846);
and UO_1067 (O_1067,N_9956,N_9902);
or UO_1068 (O_1068,N_9885,N_9903);
or UO_1069 (O_1069,N_9821,N_9830);
or UO_1070 (O_1070,N_9897,N_9949);
nor UO_1071 (O_1071,N_9980,N_9911);
or UO_1072 (O_1072,N_9826,N_9920);
nand UO_1073 (O_1073,N_9985,N_9965);
or UO_1074 (O_1074,N_9885,N_9809);
and UO_1075 (O_1075,N_9968,N_9953);
nor UO_1076 (O_1076,N_9863,N_9887);
nand UO_1077 (O_1077,N_9837,N_9883);
and UO_1078 (O_1078,N_9923,N_9987);
or UO_1079 (O_1079,N_9820,N_9917);
nand UO_1080 (O_1080,N_9834,N_9938);
nand UO_1081 (O_1081,N_9917,N_9980);
nor UO_1082 (O_1082,N_9953,N_9923);
nand UO_1083 (O_1083,N_9913,N_9864);
nand UO_1084 (O_1084,N_9862,N_9934);
and UO_1085 (O_1085,N_9968,N_9977);
nor UO_1086 (O_1086,N_9908,N_9847);
nand UO_1087 (O_1087,N_9900,N_9982);
and UO_1088 (O_1088,N_9872,N_9878);
and UO_1089 (O_1089,N_9899,N_9909);
nor UO_1090 (O_1090,N_9941,N_9955);
nor UO_1091 (O_1091,N_9848,N_9840);
nor UO_1092 (O_1092,N_9955,N_9989);
nor UO_1093 (O_1093,N_9997,N_9868);
and UO_1094 (O_1094,N_9904,N_9993);
or UO_1095 (O_1095,N_9991,N_9895);
or UO_1096 (O_1096,N_9963,N_9996);
and UO_1097 (O_1097,N_9924,N_9914);
and UO_1098 (O_1098,N_9891,N_9815);
and UO_1099 (O_1099,N_9820,N_9918);
nand UO_1100 (O_1100,N_9854,N_9907);
or UO_1101 (O_1101,N_9855,N_9949);
nor UO_1102 (O_1102,N_9965,N_9896);
nor UO_1103 (O_1103,N_9945,N_9861);
xor UO_1104 (O_1104,N_9871,N_9931);
nand UO_1105 (O_1105,N_9864,N_9859);
or UO_1106 (O_1106,N_9852,N_9856);
and UO_1107 (O_1107,N_9937,N_9851);
or UO_1108 (O_1108,N_9884,N_9919);
nor UO_1109 (O_1109,N_9878,N_9829);
nor UO_1110 (O_1110,N_9984,N_9975);
or UO_1111 (O_1111,N_9881,N_9876);
nor UO_1112 (O_1112,N_9942,N_9936);
and UO_1113 (O_1113,N_9882,N_9893);
nand UO_1114 (O_1114,N_9900,N_9825);
and UO_1115 (O_1115,N_9948,N_9998);
or UO_1116 (O_1116,N_9851,N_9909);
and UO_1117 (O_1117,N_9975,N_9888);
or UO_1118 (O_1118,N_9868,N_9857);
or UO_1119 (O_1119,N_9920,N_9988);
and UO_1120 (O_1120,N_9937,N_9849);
or UO_1121 (O_1121,N_9928,N_9832);
or UO_1122 (O_1122,N_9929,N_9977);
nand UO_1123 (O_1123,N_9868,N_9957);
and UO_1124 (O_1124,N_9970,N_9883);
nand UO_1125 (O_1125,N_9838,N_9980);
and UO_1126 (O_1126,N_9814,N_9885);
or UO_1127 (O_1127,N_9903,N_9812);
or UO_1128 (O_1128,N_9913,N_9868);
nand UO_1129 (O_1129,N_9864,N_9986);
and UO_1130 (O_1130,N_9905,N_9987);
or UO_1131 (O_1131,N_9964,N_9962);
nand UO_1132 (O_1132,N_9958,N_9876);
nand UO_1133 (O_1133,N_9962,N_9996);
or UO_1134 (O_1134,N_9871,N_9905);
nor UO_1135 (O_1135,N_9925,N_9803);
nor UO_1136 (O_1136,N_9911,N_9864);
nand UO_1137 (O_1137,N_9901,N_9995);
nor UO_1138 (O_1138,N_9949,N_9912);
and UO_1139 (O_1139,N_9837,N_9830);
and UO_1140 (O_1140,N_9894,N_9943);
and UO_1141 (O_1141,N_9984,N_9996);
nor UO_1142 (O_1142,N_9978,N_9808);
or UO_1143 (O_1143,N_9930,N_9849);
nand UO_1144 (O_1144,N_9818,N_9862);
nor UO_1145 (O_1145,N_9811,N_9909);
and UO_1146 (O_1146,N_9861,N_9913);
or UO_1147 (O_1147,N_9848,N_9838);
nor UO_1148 (O_1148,N_9916,N_9897);
nor UO_1149 (O_1149,N_9825,N_9828);
and UO_1150 (O_1150,N_9864,N_9866);
or UO_1151 (O_1151,N_9963,N_9888);
nand UO_1152 (O_1152,N_9977,N_9904);
and UO_1153 (O_1153,N_9810,N_9812);
or UO_1154 (O_1154,N_9918,N_9849);
xnor UO_1155 (O_1155,N_9845,N_9866);
nand UO_1156 (O_1156,N_9998,N_9887);
and UO_1157 (O_1157,N_9873,N_9843);
nand UO_1158 (O_1158,N_9951,N_9812);
nand UO_1159 (O_1159,N_9889,N_9989);
nor UO_1160 (O_1160,N_9818,N_9814);
nand UO_1161 (O_1161,N_9830,N_9920);
or UO_1162 (O_1162,N_9913,N_9917);
or UO_1163 (O_1163,N_9891,N_9998);
nand UO_1164 (O_1164,N_9883,N_9889);
and UO_1165 (O_1165,N_9869,N_9995);
nand UO_1166 (O_1166,N_9997,N_9976);
xor UO_1167 (O_1167,N_9976,N_9927);
xor UO_1168 (O_1168,N_9977,N_9937);
or UO_1169 (O_1169,N_9802,N_9829);
and UO_1170 (O_1170,N_9823,N_9877);
nor UO_1171 (O_1171,N_9981,N_9828);
and UO_1172 (O_1172,N_9916,N_9822);
or UO_1173 (O_1173,N_9845,N_9968);
nor UO_1174 (O_1174,N_9847,N_9837);
nor UO_1175 (O_1175,N_9959,N_9942);
and UO_1176 (O_1176,N_9946,N_9887);
nand UO_1177 (O_1177,N_9916,N_9997);
nand UO_1178 (O_1178,N_9924,N_9973);
nor UO_1179 (O_1179,N_9983,N_9866);
nand UO_1180 (O_1180,N_9933,N_9881);
nand UO_1181 (O_1181,N_9936,N_9917);
xor UO_1182 (O_1182,N_9882,N_9921);
nor UO_1183 (O_1183,N_9829,N_9876);
and UO_1184 (O_1184,N_9914,N_9912);
and UO_1185 (O_1185,N_9949,N_9816);
or UO_1186 (O_1186,N_9885,N_9904);
and UO_1187 (O_1187,N_9959,N_9941);
nand UO_1188 (O_1188,N_9942,N_9846);
or UO_1189 (O_1189,N_9853,N_9902);
nand UO_1190 (O_1190,N_9993,N_9897);
nand UO_1191 (O_1191,N_9989,N_9953);
and UO_1192 (O_1192,N_9842,N_9987);
nand UO_1193 (O_1193,N_9876,N_9952);
or UO_1194 (O_1194,N_9872,N_9938);
nor UO_1195 (O_1195,N_9874,N_9804);
and UO_1196 (O_1196,N_9934,N_9980);
nor UO_1197 (O_1197,N_9992,N_9890);
nand UO_1198 (O_1198,N_9947,N_9908);
nand UO_1199 (O_1199,N_9890,N_9831);
or UO_1200 (O_1200,N_9842,N_9989);
nand UO_1201 (O_1201,N_9817,N_9811);
xor UO_1202 (O_1202,N_9841,N_9855);
and UO_1203 (O_1203,N_9916,N_9943);
or UO_1204 (O_1204,N_9903,N_9935);
or UO_1205 (O_1205,N_9807,N_9955);
or UO_1206 (O_1206,N_9845,N_9976);
and UO_1207 (O_1207,N_9962,N_9940);
or UO_1208 (O_1208,N_9976,N_9984);
nand UO_1209 (O_1209,N_9903,N_9880);
and UO_1210 (O_1210,N_9860,N_9871);
xnor UO_1211 (O_1211,N_9872,N_9977);
nand UO_1212 (O_1212,N_9815,N_9812);
nor UO_1213 (O_1213,N_9833,N_9813);
xor UO_1214 (O_1214,N_9981,N_9890);
and UO_1215 (O_1215,N_9926,N_9873);
nand UO_1216 (O_1216,N_9823,N_9827);
or UO_1217 (O_1217,N_9912,N_9901);
and UO_1218 (O_1218,N_9831,N_9827);
or UO_1219 (O_1219,N_9942,N_9879);
nor UO_1220 (O_1220,N_9855,N_9935);
and UO_1221 (O_1221,N_9947,N_9939);
or UO_1222 (O_1222,N_9967,N_9812);
nor UO_1223 (O_1223,N_9834,N_9838);
nor UO_1224 (O_1224,N_9952,N_9856);
and UO_1225 (O_1225,N_9849,N_9908);
and UO_1226 (O_1226,N_9832,N_9837);
or UO_1227 (O_1227,N_9927,N_9867);
xnor UO_1228 (O_1228,N_9894,N_9862);
nor UO_1229 (O_1229,N_9887,N_9983);
and UO_1230 (O_1230,N_9890,N_9990);
nor UO_1231 (O_1231,N_9859,N_9860);
nor UO_1232 (O_1232,N_9919,N_9945);
nand UO_1233 (O_1233,N_9941,N_9821);
or UO_1234 (O_1234,N_9813,N_9983);
nand UO_1235 (O_1235,N_9911,N_9947);
nand UO_1236 (O_1236,N_9964,N_9987);
or UO_1237 (O_1237,N_9968,N_9818);
and UO_1238 (O_1238,N_9847,N_9872);
and UO_1239 (O_1239,N_9988,N_9929);
and UO_1240 (O_1240,N_9971,N_9868);
nor UO_1241 (O_1241,N_9866,N_9883);
nand UO_1242 (O_1242,N_9875,N_9891);
or UO_1243 (O_1243,N_9837,N_9954);
or UO_1244 (O_1244,N_9904,N_9923);
xor UO_1245 (O_1245,N_9843,N_9983);
nor UO_1246 (O_1246,N_9913,N_9870);
or UO_1247 (O_1247,N_9802,N_9898);
nand UO_1248 (O_1248,N_9923,N_9983);
and UO_1249 (O_1249,N_9979,N_9826);
and UO_1250 (O_1250,N_9953,N_9905);
and UO_1251 (O_1251,N_9994,N_9829);
nor UO_1252 (O_1252,N_9819,N_9965);
and UO_1253 (O_1253,N_9925,N_9935);
or UO_1254 (O_1254,N_9909,N_9916);
xnor UO_1255 (O_1255,N_9820,N_9985);
and UO_1256 (O_1256,N_9807,N_9856);
and UO_1257 (O_1257,N_9871,N_9976);
and UO_1258 (O_1258,N_9915,N_9927);
and UO_1259 (O_1259,N_9809,N_9986);
or UO_1260 (O_1260,N_9980,N_9821);
or UO_1261 (O_1261,N_9844,N_9982);
nand UO_1262 (O_1262,N_9862,N_9883);
and UO_1263 (O_1263,N_9933,N_9906);
and UO_1264 (O_1264,N_9930,N_9835);
nor UO_1265 (O_1265,N_9828,N_9820);
or UO_1266 (O_1266,N_9912,N_9893);
nor UO_1267 (O_1267,N_9851,N_9862);
nor UO_1268 (O_1268,N_9867,N_9842);
and UO_1269 (O_1269,N_9986,N_9973);
nand UO_1270 (O_1270,N_9883,N_9826);
nand UO_1271 (O_1271,N_9851,N_9978);
or UO_1272 (O_1272,N_9810,N_9833);
or UO_1273 (O_1273,N_9829,N_9977);
or UO_1274 (O_1274,N_9972,N_9944);
nand UO_1275 (O_1275,N_9825,N_9977);
nand UO_1276 (O_1276,N_9899,N_9866);
and UO_1277 (O_1277,N_9802,N_9892);
or UO_1278 (O_1278,N_9873,N_9882);
and UO_1279 (O_1279,N_9996,N_9999);
nor UO_1280 (O_1280,N_9970,N_9854);
nand UO_1281 (O_1281,N_9813,N_9982);
or UO_1282 (O_1282,N_9833,N_9987);
nand UO_1283 (O_1283,N_9965,N_9943);
nor UO_1284 (O_1284,N_9834,N_9804);
nand UO_1285 (O_1285,N_9805,N_9853);
nor UO_1286 (O_1286,N_9802,N_9927);
nor UO_1287 (O_1287,N_9867,N_9831);
nor UO_1288 (O_1288,N_9813,N_9978);
or UO_1289 (O_1289,N_9995,N_9929);
or UO_1290 (O_1290,N_9947,N_9945);
or UO_1291 (O_1291,N_9893,N_9918);
nor UO_1292 (O_1292,N_9875,N_9939);
or UO_1293 (O_1293,N_9958,N_9841);
and UO_1294 (O_1294,N_9819,N_9829);
and UO_1295 (O_1295,N_9921,N_9862);
xor UO_1296 (O_1296,N_9954,N_9855);
xnor UO_1297 (O_1297,N_9842,N_9855);
nand UO_1298 (O_1298,N_9987,N_9852);
nand UO_1299 (O_1299,N_9843,N_9925);
and UO_1300 (O_1300,N_9873,N_9969);
nand UO_1301 (O_1301,N_9863,N_9935);
nor UO_1302 (O_1302,N_9940,N_9892);
nand UO_1303 (O_1303,N_9857,N_9982);
nand UO_1304 (O_1304,N_9800,N_9996);
xor UO_1305 (O_1305,N_9841,N_9800);
or UO_1306 (O_1306,N_9971,N_9849);
or UO_1307 (O_1307,N_9999,N_9888);
and UO_1308 (O_1308,N_9870,N_9807);
nor UO_1309 (O_1309,N_9881,N_9888);
nor UO_1310 (O_1310,N_9954,N_9886);
nor UO_1311 (O_1311,N_9947,N_9874);
or UO_1312 (O_1312,N_9852,N_9943);
nand UO_1313 (O_1313,N_9843,N_9898);
nand UO_1314 (O_1314,N_9989,N_9944);
nand UO_1315 (O_1315,N_9914,N_9967);
or UO_1316 (O_1316,N_9853,N_9952);
nor UO_1317 (O_1317,N_9864,N_9852);
xor UO_1318 (O_1318,N_9913,N_9878);
nand UO_1319 (O_1319,N_9903,N_9813);
nand UO_1320 (O_1320,N_9817,N_9927);
or UO_1321 (O_1321,N_9829,N_9928);
nor UO_1322 (O_1322,N_9861,N_9855);
and UO_1323 (O_1323,N_9969,N_9811);
and UO_1324 (O_1324,N_9986,N_9917);
and UO_1325 (O_1325,N_9894,N_9930);
or UO_1326 (O_1326,N_9923,N_9897);
nor UO_1327 (O_1327,N_9971,N_9806);
and UO_1328 (O_1328,N_9995,N_9936);
nor UO_1329 (O_1329,N_9872,N_9941);
nand UO_1330 (O_1330,N_9814,N_9813);
nand UO_1331 (O_1331,N_9801,N_9884);
and UO_1332 (O_1332,N_9873,N_9990);
or UO_1333 (O_1333,N_9875,N_9847);
and UO_1334 (O_1334,N_9923,N_9988);
and UO_1335 (O_1335,N_9878,N_9866);
nand UO_1336 (O_1336,N_9813,N_9858);
nand UO_1337 (O_1337,N_9852,N_9809);
and UO_1338 (O_1338,N_9928,N_9918);
or UO_1339 (O_1339,N_9885,N_9802);
nand UO_1340 (O_1340,N_9813,N_9914);
nand UO_1341 (O_1341,N_9841,N_9834);
xnor UO_1342 (O_1342,N_9984,N_9895);
and UO_1343 (O_1343,N_9922,N_9906);
or UO_1344 (O_1344,N_9966,N_9918);
and UO_1345 (O_1345,N_9995,N_9935);
nand UO_1346 (O_1346,N_9898,N_9959);
or UO_1347 (O_1347,N_9945,N_9832);
nand UO_1348 (O_1348,N_9945,N_9816);
or UO_1349 (O_1349,N_9938,N_9986);
and UO_1350 (O_1350,N_9961,N_9877);
and UO_1351 (O_1351,N_9928,N_9821);
nor UO_1352 (O_1352,N_9964,N_9997);
and UO_1353 (O_1353,N_9986,N_9855);
xnor UO_1354 (O_1354,N_9813,N_9850);
nand UO_1355 (O_1355,N_9977,N_9946);
or UO_1356 (O_1356,N_9844,N_9940);
xnor UO_1357 (O_1357,N_9910,N_9838);
or UO_1358 (O_1358,N_9978,N_9984);
nor UO_1359 (O_1359,N_9808,N_9840);
nor UO_1360 (O_1360,N_9865,N_9954);
nand UO_1361 (O_1361,N_9921,N_9879);
and UO_1362 (O_1362,N_9816,N_9955);
and UO_1363 (O_1363,N_9875,N_9819);
nand UO_1364 (O_1364,N_9805,N_9817);
and UO_1365 (O_1365,N_9990,N_9937);
nor UO_1366 (O_1366,N_9809,N_9879);
and UO_1367 (O_1367,N_9803,N_9828);
and UO_1368 (O_1368,N_9870,N_9917);
or UO_1369 (O_1369,N_9926,N_9937);
nand UO_1370 (O_1370,N_9845,N_9944);
nor UO_1371 (O_1371,N_9839,N_9878);
nand UO_1372 (O_1372,N_9874,N_9808);
xor UO_1373 (O_1373,N_9877,N_9883);
nor UO_1374 (O_1374,N_9962,N_9807);
or UO_1375 (O_1375,N_9963,N_9854);
and UO_1376 (O_1376,N_9916,N_9872);
nor UO_1377 (O_1377,N_9970,N_9849);
and UO_1378 (O_1378,N_9882,N_9869);
xor UO_1379 (O_1379,N_9815,N_9892);
nand UO_1380 (O_1380,N_9909,N_9944);
and UO_1381 (O_1381,N_9906,N_9836);
and UO_1382 (O_1382,N_9946,N_9824);
and UO_1383 (O_1383,N_9836,N_9887);
nand UO_1384 (O_1384,N_9882,N_9804);
nand UO_1385 (O_1385,N_9966,N_9984);
or UO_1386 (O_1386,N_9954,N_9829);
and UO_1387 (O_1387,N_9864,N_9831);
or UO_1388 (O_1388,N_9987,N_9826);
and UO_1389 (O_1389,N_9942,N_9990);
nand UO_1390 (O_1390,N_9818,N_9859);
and UO_1391 (O_1391,N_9999,N_9837);
nand UO_1392 (O_1392,N_9918,N_9881);
nor UO_1393 (O_1393,N_9994,N_9986);
nand UO_1394 (O_1394,N_9853,N_9835);
nor UO_1395 (O_1395,N_9846,N_9966);
and UO_1396 (O_1396,N_9909,N_9888);
nand UO_1397 (O_1397,N_9824,N_9899);
nor UO_1398 (O_1398,N_9975,N_9950);
nor UO_1399 (O_1399,N_9827,N_9893);
nor UO_1400 (O_1400,N_9879,N_9863);
nor UO_1401 (O_1401,N_9937,N_9883);
or UO_1402 (O_1402,N_9961,N_9859);
nor UO_1403 (O_1403,N_9909,N_9932);
nand UO_1404 (O_1404,N_9923,N_9865);
nor UO_1405 (O_1405,N_9988,N_9802);
and UO_1406 (O_1406,N_9847,N_9807);
or UO_1407 (O_1407,N_9921,N_9972);
or UO_1408 (O_1408,N_9915,N_9963);
nand UO_1409 (O_1409,N_9883,N_9894);
or UO_1410 (O_1410,N_9911,N_9848);
or UO_1411 (O_1411,N_9817,N_9825);
and UO_1412 (O_1412,N_9898,N_9822);
or UO_1413 (O_1413,N_9893,N_9973);
and UO_1414 (O_1414,N_9831,N_9873);
nor UO_1415 (O_1415,N_9838,N_9810);
nand UO_1416 (O_1416,N_9811,N_9989);
and UO_1417 (O_1417,N_9928,N_9803);
nand UO_1418 (O_1418,N_9871,N_9950);
and UO_1419 (O_1419,N_9834,N_9821);
nor UO_1420 (O_1420,N_9839,N_9833);
or UO_1421 (O_1421,N_9958,N_9905);
and UO_1422 (O_1422,N_9800,N_9831);
or UO_1423 (O_1423,N_9836,N_9912);
nor UO_1424 (O_1424,N_9891,N_9958);
or UO_1425 (O_1425,N_9844,N_9987);
xnor UO_1426 (O_1426,N_9879,N_9982);
nand UO_1427 (O_1427,N_9919,N_9821);
nor UO_1428 (O_1428,N_9865,N_9937);
and UO_1429 (O_1429,N_9978,N_9840);
and UO_1430 (O_1430,N_9830,N_9965);
nand UO_1431 (O_1431,N_9939,N_9826);
nand UO_1432 (O_1432,N_9968,N_9933);
nand UO_1433 (O_1433,N_9807,N_9995);
nor UO_1434 (O_1434,N_9823,N_9834);
or UO_1435 (O_1435,N_9863,N_9846);
nor UO_1436 (O_1436,N_9892,N_9874);
nand UO_1437 (O_1437,N_9804,N_9978);
nand UO_1438 (O_1438,N_9840,N_9818);
and UO_1439 (O_1439,N_9831,N_9946);
and UO_1440 (O_1440,N_9918,N_9964);
nor UO_1441 (O_1441,N_9933,N_9959);
nor UO_1442 (O_1442,N_9969,N_9800);
xnor UO_1443 (O_1443,N_9888,N_9857);
or UO_1444 (O_1444,N_9999,N_9844);
and UO_1445 (O_1445,N_9915,N_9838);
nand UO_1446 (O_1446,N_9815,N_9857);
or UO_1447 (O_1447,N_9850,N_9900);
and UO_1448 (O_1448,N_9834,N_9992);
nor UO_1449 (O_1449,N_9931,N_9837);
and UO_1450 (O_1450,N_9905,N_9982);
and UO_1451 (O_1451,N_9897,N_9807);
nand UO_1452 (O_1452,N_9823,N_9913);
nand UO_1453 (O_1453,N_9926,N_9865);
nor UO_1454 (O_1454,N_9969,N_9960);
nand UO_1455 (O_1455,N_9858,N_9877);
nand UO_1456 (O_1456,N_9802,N_9972);
nand UO_1457 (O_1457,N_9958,N_9977);
nor UO_1458 (O_1458,N_9851,N_9987);
nand UO_1459 (O_1459,N_9854,N_9886);
or UO_1460 (O_1460,N_9840,N_9909);
nand UO_1461 (O_1461,N_9871,N_9975);
nor UO_1462 (O_1462,N_9912,N_9825);
and UO_1463 (O_1463,N_9881,N_9997);
and UO_1464 (O_1464,N_9907,N_9870);
or UO_1465 (O_1465,N_9919,N_9834);
nor UO_1466 (O_1466,N_9911,N_9854);
nand UO_1467 (O_1467,N_9847,N_9981);
and UO_1468 (O_1468,N_9803,N_9862);
or UO_1469 (O_1469,N_9997,N_9980);
nor UO_1470 (O_1470,N_9981,N_9873);
nand UO_1471 (O_1471,N_9871,N_9943);
nand UO_1472 (O_1472,N_9815,N_9914);
nand UO_1473 (O_1473,N_9855,N_9972);
or UO_1474 (O_1474,N_9910,N_9804);
and UO_1475 (O_1475,N_9977,N_9849);
nand UO_1476 (O_1476,N_9861,N_9965);
or UO_1477 (O_1477,N_9856,N_9875);
or UO_1478 (O_1478,N_9802,N_9852);
and UO_1479 (O_1479,N_9919,N_9872);
xor UO_1480 (O_1480,N_9944,N_9841);
nor UO_1481 (O_1481,N_9846,N_9943);
nor UO_1482 (O_1482,N_9948,N_9823);
nor UO_1483 (O_1483,N_9823,N_9956);
nand UO_1484 (O_1484,N_9921,N_9918);
nand UO_1485 (O_1485,N_9925,N_9987);
and UO_1486 (O_1486,N_9967,N_9824);
and UO_1487 (O_1487,N_9849,N_9954);
and UO_1488 (O_1488,N_9880,N_9833);
and UO_1489 (O_1489,N_9940,N_9867);
and UO_1490 (O_1490,N_9965,N_9992);
and UO_1491 (O_1491,N_9830,N_9989);
or UO_1492 (O_1492,N_9932,N_9965);
and UO_1493 (O_1493,N_9910,N_9969);
nand UO_1494 (O_1494,N_9831,N_9984);
and UO_1495 (O_1495,N_9875,N_9869);
and UO_1496 (O_1496,N_9823,N_9818);
and UO_1497 (O_1497,N_9986,N_9830);
or UO_1498 (O_1498,N_9850,N_9931);
nand UO_1499 (O_1499,N_9841,N_9986);
endmodule