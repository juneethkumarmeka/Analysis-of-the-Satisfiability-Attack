module basic_750_5000_1000_5_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
xor U0 (N_0,In_86,In_427);
nor U1 (N_1,In_501,In_554);
nor U2 (N_2,In_34,In_289);
nand U3 (N_3,In_516,In_735);
or U4 (N_4,In_649,In_471);
or U5 (N_5,In_416,In_212);
and U6 (N_6,In_737,In_312);
nor U7 (N_7,In_8,In_321);
or U8 (N_8,In_472,In_716);
nor U9 (N_9,In_221,In_238);
or U10 (N_10,In_378,In_461);
or U11 (N_11,In_698,In_147);
xnor U12 (N_12,In_275,In_139);
nor U13 (N_13,In_409,In_180);
and U14 (N_14,In_459,In_30);
and U15 (N_15,In_647,In_656);
nand U16 (N_16,In_567,In_385);
and U17 (N_17,In_497,In_413);
xor U18 (N_18,In_182,In_343);
nand U19 (N_19,In_534,In_125);
xnor U20 (N_20,In_133,In_600);
nor U21 (N_21,In_184,In_106);
nand U22 (N_22,In_678,In_127);
xor U23 (N_23,In_327,In_470);
nand U24 (N_24,In_187,In_85);
nor U25 (N_25,In_183,In_732);
nand U26 (N_26,In_415,In_157);
or U27 (N_27,In_529,In_671);
and U28 (N_28,In_742,In_120);
and U29 (N_29,In_224,In_483);
nor U30 (N_30,In_746,In_488);
and U31 (N_31,In_336,In_747);
xnor U32 (N_32,In_91,In_654);
and U33 (N_33,In_718,In_577);
nand U34 (N_34,In_54,In_196);
nand U35 (N_35,In_103,In_560);
xnor U36 (N_36,In_39,In_69);
nor U37 (N_37,In_94,In_709);
nand U38 (N_38,In_513,In_298);
nor U39 (N_39,In_191,In_435);
and U40 (N_40,In_198,In_725);
nand U41 (N_41,In_525,In_363);
and U42 (N_42,In_229,In_290);
or U43 (N_43,In_154,In_220);
xnor U44 (N_44,In_53,In_268);
nand U45 (N_45,In_116,In_694);
xnor U46 (N_46,In_434,In_580);
nand U47 (N_47,In_587,In_482);
nor U48 (N_48,In_79,In_708);
nand U49 (N_49,In_401,In_429);
and U50 (N_50,In_419,In_328);
and U51 (N_51,In_551,In_109);
and U52 (N_52,In_391,In_546);
nand U53 (N_53,In_699,In_121);
nand U54 (N_54,In_168,In_355);
nor U55 (N_55,In_710,In_216);
xor U56 (N_56,In_98,In_447);
nand U57 (N_57,In_2,In_7);
nor U58 (N_58,In_178,In_72);
xor U59 (N_59,In_228,In_703);
or U60 (N_60,In_644,In_274);
and U61 (N_61,In_349,In_602);
xor U62 (N_62,In_372,In_80);
and U63 (N_63,In_662,In_451);
nor U64 (N_64,In_160,In_190);
nor U65 (N_65,In_402,In_392);
or U66 (N_66,In_235,In_666);
and U67 (N_67,In_324,In_664);
and U68 (N_68,In_421,In_464);
or U69 (N_69,In_663,In_672);
or U70 (N_70,In_232,In_337);
xnor U71 (N_71,In_27,In_712);
xnor U72 (N_72,In_47,In_576);
or U73 (N_73,In_117,In_338);
xor U74 (N_74,In_4,In_548);
nor U75 (N_75,In_440,In_35);
nand U76 (N_76,In_146,In_454);
xnor U77 (N_77,In_405,In_367);
or U78 (N_78,In_730,In_153);
nand U79 (N_79,In_628,In_215);
nand U80 (N_80,In_445,In_45);
nand U81 (N_81,In_37,In_325);
nor U82 (N_82,In_633,In_75);
or U83 (N_83,In_261,In_417);
or U84 (N_84,In_186,In_60);
nand U85 (N_85,In_340,In_739);
xor U86 (N_86,In_585,In_295);
nor U87 (N_87,In_31,In_642);
and U88 (N_88,In_137,In_700);
xor U89 (N_89,In_502,In_179);
nor U90 (N_90,In_403,In_744);
or U91 (N_91,In_498,In_255);
and U92 (N_92,In_462,In_715);
nand U93 (N_93,In_0,In_517);
or U94 (N_94,In_350,In_272);
or U95 (N_95,In_219,In_748);
or U96 (N_96,In_676,In_118);
xor U97 (N_97,In_729,In_648);
nand U98 (N_98,In_252,In_704);
nor U99 (N_99,In_582,In_62);
nor U100 (N_100,In_727,In_315);
and U101 (N_101,In_277,In_428);
xor U102 (N_102,In_404,In_493);
or U103 (N_103,In_563,In_561);
or U104 (N_104,In_209,In_724);
nor U105 (N_105,In_575,In_618);
nor U106 (N_106,In_193,In_568);
nor U107 (N_107,In_697,In_134);
or U108 (N_108,In_129,In_185);
xor U109 (N_109,In_282,In_384);
or U110 (N_110,In_344,In_559);
nand U111 (N_111,In_100,In_484);
or U112 (N_112,In_197,In_16);
nand U113 (N_113,In_266,In_506);
and U114 (N_114,In_669,In_19);
nor U115 (N_115,In_307,In_379);
nand U116 (N_116,In_641,In_164);
nor U117 (N_117,In_466,In_36);
and U118 (N_118,In_695,In_140);
nor U119 (N_119,In_84,In_584);
xnor U120 (N_120,In_627,In_713);
nand U121 (N_121,In_523,In_302);
or U122 (N_122,In_696,In_562);
and U123 (N_123,In_13,In_308);
nand U124 (N_124,In_591,In_607);
xnor U125 (N_125,In_115,In_78);
nand U126 (N_126,In_592,In_539);
nand U127 (N_127,In_364,In_543);
or U128 (N_128,In_284,In_21);
and U129 (N_129,In_393,In_144);
nand U130 (N_130,In_174,In_108);
or U131 (N_131,In_331,In_566);
nand U132 (N_132,In_319,In_262);
xnor U133 (N_133,In_531,In_354);
and U134 (N_134,In_387,In_496);
xnor U135 (N_135,In_468,In_122);
nor U136 (N_136,In_32,In_524);
nor U137 (N_137,In_204,In_356);
nand U138 (N_138,In_227,In_389);
and U139 (N_139,In_638,In_136);
xor U140 (N_140,In_291,In_565);
xnor U141 (N_141,In_104,In_233);
nor U142 (N_142,In_621,In_256);
xor U143 (N_143,In_583,In_130);
or U144 (N_144,In_503,In_43);
and U145 (N_145,In_128,In_423);
xnor U146 (N_146,In_432,In_612);
or U147 (N_147,In_51,In_194);
or U148 (N_148,In_446,In_126);
and U149 (N_149,In_249,In_200);
xor U150 (N_150,In_481,In_303);
nor U151 (N_151,In_689,In_226);
nor U152 (N_152,In_711,In_728);
and U153 (N_153,In_95,In_661);
and U154 (N_154,In_195,In_571);
and U155 (N_155,In_465,In_717);
xnor U156 (N_156,In_203,In_489);
nand U157 (N_157,In_131,In_223);
nor U158 (N_158,In_519,In_682);
and U159 (N_159,In_217,In_486);
or U160 (N_160,In_151,In_145);
and U161 (N_161,In_407,In_453);
nand U162 (N_162,In_11,In_259);
nor U163 (N_163,In_476,In_335);
or U164 (N_164,In_492,In_515);
xnor U165 (N_165,In_723,In_141);
xor U166 (N_166,In_613,In_646);
xor U167 (N_167,In_681,In_594);
nand U168 (N_168,In_317,In_736);
nand U169 (N_169,In_260,In_480);
xor U170 (N_170,In_586,In_635);
nand U171 (N_171,In_225,In_541);
xnor U172 (N_172,In_376,In_509);
or U173 (N_173,In_165,In_706);
nor U174 (N_174,In_251,In_280);
and U175 (N_175,In_522,In_161);
xor U176 (N_176,In_683,In_70);
nor U177 (N_177,In_33,In_166);
nand U178 (N_178,In_458,In_74);
and U179 (N_179,In_601,In_691);
nor U180 (N_180,In_278,In_383);
nor U181 (N_181,In_510,In_107);
nand U182 (N_182,In_386,In_236);
and U183 (N_183,In_538,In_469);
nor U184 (N_184,In_172,In_639);
nand U185 (N_185,In_645,In_443);
nand U186 (N_186,In_526,In_514);
nand U187 (N_187,In_520,In_660);
and U188 (N_188,In_499,In_684);
xnor U189 (N_189,In_50,In_6);
and U190 (N_190,In_597,In_412);
and U191 (N_191,In_345,In_623);
and U192 (N_192,In_143,In_617);
and U193 (N_193,In_270,In_436);
nand U194 (N_194,In_29,In_692);
nand U195 (N_195,In_20,In_213);
nand U196 (N_196,In_640,In_605);
nor U197 (N_197,In_205,In_102);
nor U198 (N_198,In_439,In_540);
nor U199 (N_199,In_388,In_579);
xnor U200 (N_200,In_474,In_420);
xor U201 (N_201,In_686,In_679);
nor U202 (N_202,In_398,In_201);
nand U203 (N_203,In_83,In_555);
or U204 (N_204,In_377,In_248);
nand U205 (N_205,In_693,In_169);
xor U206 (N_206,In_242,In_521);
and U207 (N_207,In_487,In_422);
and U208 (N_208,In_52,In_171);
nand U209 (N_209,In_593,In_473);
or U210 (N_210,In_158,In_622);
and U211 (N_211,In_92,In_655);
and U212 (N_212,In_301,In_347);
nor U213 (N_213,In_76,In_5);
or U214 (N_214,In_680,In_722);
or U215 (N_215,In_370,In_89);
nor U216 (N_216,In_258,In_668);
or U217 (N_217,In_1,In_437);
xnor U218 (N_218,In_619,In_279);
xor U219 (N_219,In_490,In_537);
xnor U220 (N_220,In_606,In_558);
and U221 (N_221,In_518,In_188);
or U222 (N_222,In_626,In_3);
and U223 (N_223,In_310,In_332);
or U224 (N_224,In_374,In_265);
nand U225 (N_225,In_170,In_346);
nand U226 (N_226,In_293,In_142);
or U227 (N_227,In_615,In_323);
and U228 (N_228,In_112,In_24);
nand U229 (N_229,In_296,In_101);
or U230 (N_230,In_64,In_463);
xnor U231 (N_231,In_749,In_659);
and U232 (N_232,In_477,In_285);
or U233 (N_233,In_743,In_528);
nor U234 (N_234,In_556,In_105);
nand U235 (N_235,In_316,In_65);
and U236 (N_236,In_675,In_239);
and U237 (N_237,In_589,In_500);
nor U238 (N_238,In_382,In_342);
xnor U239 (N_239,In_48,In_424);
nor U240 (N_240,In_15,In_93);
and U241 (N_241,In_214,In_527);
nand U242 (N_242,In_721,In_495);
xnor U243 (N_243,In_348,In_17);
nor U244 (N_244,In_467,In_550);
nor U245 (N_245,In_38,In_114);
and U246 (N_246,In_267,In_569);
or U247 (N_247,In_66,In_629);
or U248 (N_248,In_599,In_400);
nor U249 (N_249,In_365,In_720);
or U250 (N_250,In_394,In_44);
or U251 (N_251,In_734,In_155);
xor U252 (N_252,In_287,In_673);
nand U253 (N_253,In_42,In_243);
nor U254 (N_254,In_138,In_449);
or U255 (N_255,In_726,In_369);
and U256 (N_256,In_22,In_59);
xor U257 (N_257,In_552,In_269);
and U258 (N_258,In_254,In_381);
nand U259 (N_259,In_81,In_14);
nand U260 (N_260,In_478,In_741);
nand U261 (N_261,In_333,In_82);
and U262 (N_262,In_23,In_536);
xor U263 (N_263,In_351,In_281);
xnor U264 (N_264,In_677,In_740);
xor U265 (N_265,In_246,In_148);
xor U266 (N_266,In_111,In_110);
and U267 (N_267,In_123,In_653);
xnor U268 (N_268,In_244,In_590);
nor U269 (N_269,In_485,In_192);
nor U270 (N_270,In_177,In_12);
nand U271 (N_271,In_442,In_444);
nor U272 (N_272,In_334,In_207);
or U273 (N_273,In_124,In_595);
nand U274 (N_274,In_479,In_610);
nor U275 (N_275,In_399,In_330);
or U276 (N_276,In_18,In_557);
xnor U277 (N_277,In_175,In_208);
nor U278 (N_278,In_250,In_373);
and U279 (N_279,In_222,In_341);
or U280 (N_280,In_634,In_264);
and U281 (N_281,In_339,In_156);
and U282 (N_282,In_58,In_455);
xnor U283 (N_283,In_701,In_230);
and U284 (N_284,In_326,In_652);
nor U285 (N_285,In_438,In_410);
nor U286 (N_286,In_674,In_288);
and U287 (N_287,In_90,In_452);
nand U288 (N_288,In_359,In_670);
nand U289 (N_289,In_320,In_357);
or U290 (N_290,In_685,In_719);
and U291 (N_291,In_234,In_322);
or U292 (N_292,In_532,In_237);
or U293 (N_293,In_631,In_283);
or U294 (N_294,In_304,In_530);
and U295 (N_295,In_202,In_505);
nand U296 (N_296,In_624,In_549);
nand U297 (N_297,In_276,In_176);
xor U298 (N_298,In_667,In_651);
xnor U299 (N_299,In_688,In_426);
nor U300 (N_300,In_297,In_56);
nor U301 (N_301,In_533,In_306);
and U302 (N_302,In_637,In_611);
nor U303 (N_303,In_564,In_430);
nand U304 (N_304,In_163,In_71);
or U305 (N_305,In_97,In_57);
or U306 (N_306,In_657,In_504);
xor U307 (N_307,In_494,In_665);
xnor U308 (N_308,In_457,In_574);
xor U309 (N_309,In_545,In_245);
or U310 (N_310,In_167,In_544);
xor U311 (N_311,In_313,In_41);
xor U312 (N_312,In_181,In_702);
xnor U313 (N_313,In_67,In_10);
xor U314 (N_314,In_311,In_425);
or U315 (N_315,In_77,In_433);
and U316 (N_316,In_643,In_358);
or U317 (N_317,In_596,In_448);
nor U318 (N_318,In_352,In_189);
nand U319 (N_319,In_247,In_28);
or U320 (N_320,In_218,In_26);
and U321 (N_321,In_570,In_650);
nor U322 (N_322,In_63,In_211);
xor U323 (N_323,In_271,In_714);
nand U324 (N_324,In_632,In_636);
nand U325 (N_325,In_73,In_286);
and U326 (N_326,In_511,In_294);
xor U327 (N_327,In_578,In_368);
and U328 (N_328,In_508,In_309);
nor U329 (N_329,In_396,In_707);
nor U330 (N_330,In_61,In_231);
and U331 (N_331,In_292,In_553);
nor U332 (N_332,In_273,In_49);
or U333 (N_333,In_507,In_96);
xnor U334 (N_334,In_406,In_609);
or U335 (N_335,In_257,In_305);
and U336 (N_336,In_603,In_119);
nand U337 (N_337,In_512,In_608);
xnor U338 (N_338,In_152,In_397);
or U339 (N_339,In_241,In_371);
and U340 (N_340,In_441,In_40);
nand U341 (N_341,In_572,In_690);
nand U342 (N_342,In_210,In_598);
nand U343 (N_343,In_705,In_206);
xor U344 (N_344,In_616,In_25);
and U345 (N_345,In_68,In_87);
and U346 (N_346,In_361,In_460);
xor U347 (N_347,In_588,In_614);
nor U348 (N_348,In_625,In_687);
xor U349 (N_349,In_159,In_450);
xor U350 (N_350,In_547,In_581);
or U351 (N_351,In_314,In_132);
or U352 (N_352,In_149,In_173);
nand U353 (N_353,In_380,In_733);
or U354 (N_354,In_573,In_620);
or U355 (N_355,In_150,In_731);
nor U356 (N_356,In_431,In_113);
nand U357 (N_357,In_390,In_658);
and U358 (N_358,In_395,In_375);
nor U359 (N_359,In_362,In_162);
xor U360 (N_360,In_630,In_240);
nand U361 (N_361,In_99,In_408);
and U362 (N_362,In_263,In_360);
nand U363 (N_363,In_88,In_135);
nor U364 (N_364,In_414,In_329);
nor U365 (N_365,In_542,In_411);
and U366 (N_366,In_491,In_738);
and U367 (N_367,In_353,In_300);
and U368 (N_368,In_55,In_366);
nand U369 (N_369,In_535,In_604);
nand U370 (N_370,In_199,In_299);
or U371 (N_371,In_9,In_253);
and U372 (N_372,In_318,In_418);
nor U373 (N_373,In_475,In_456);
nor U374 (N_374,In_46,In_745);
xor U375 (N_375,In_99,In_591);
nand U376 (N_376,In_649,In_127);
nand U377 (N_377,In_444,In_149);
or U378 (N_378,In_148,In_729);
nor U379 (N_379,In_239,In_203);
nand U380 (N_380,In_371,In_179);
xor U381 (N_381,In_179,In_581);
xnor U382 (N_382,In_236,In_397);
nor U383 (N_383,In_256,In_691);
or U384 (N_384,In_666,In_653);
or U385 (N_385,In_673,In_280);
nand U386 (N_386,In_541,In_599);
or U387 (N_387,In_482,In_109);
or U388 (N_388,In_481,In_665);
xnor U389 (N_389,In_117,In_132);
nand U390 (N_390,In_749,In_282);
nand U391 (N_391,In_112,In_437);
or U392 (N_392,In_229,In_20);
nor U393 (N_393,In_206,In_136);
and U394 (N_394,In_607,In_662);
nand U395 (N_395,In_75,In_697);
or U396 (N_396,In_687,In_194);
nor U397 (N_397,In_436,In_310);
xor U398 (N_398,In_640,In_93);
nor U399 (N_399,In_129,In_498);
and U400 (N_400,In_34,In_525);
or U401 (N_401,In_428,In_601);
nand U402 (N_402,In_696,In_449);
nand U403 (N_403,In_572,In_433);
or U404 (N_404,In_669,In_499);
nor U405 (N_405,In_609,In_628);
nand U406 (N_406,In_475,In_497);
or U407 (N_407,In_48,In_607);
nor U408 (N_408,In_91,In_469);
xnor U409 (N_409,In_714,In_656);
or U410 (N_410,In_678,In_331);
nand U411 (N_411,In_308,In_292);
xnor U412 (N_412,In_255,In_133);
or U413 (N_413,In_616,In_454);
nand U414 (N_414,In_490,In_527);
or U415 (N_415,In_611,In_37);
and U416 (N_416,In_342,In_266);
nand U417 (N_417,In_431,In_441);
nor U418 (N_418,In_647,In_717);
nor U419 (N_419,In_333,In_466);
xor U420 (N_420,In_326,In_507);
nor U421 (N_421,In_285,In_588);
xnor U422 (N_422,In_430,In_356);
nand U423 (N_423,In_546,In_305);
nand U424 (N_424,In_725,In_561);
nor U425 (N_425,In_742,In_636);
nand U426 (N_426,In_437,In_9);
and U427 (N_427,In_503,In_280);
xor U428 (N_428,In_637,In_727);
and U429 (N_429,In_387,In_541);
xnor U430 (N_430,In_547,In_735);
or U431 (N_431,In_505,In_734);
and U432 (N_432,In_31,In_719);
or U433 (N_433,In_108,In_535);
xnor U434 (N_434,In_213,In_161);
nand U435 (N_435,In_251,In_691);
and U436 (N_436,In_253,In_670);
or U437 (N_437,In_112,In_588);
xnor U438 (N_438,In_12,In_171);
nand U439 (N_439,In_534,In_571);
or U440 (N_440,In_547,In_214);
and U441 (N_441,In_711,In_431);
nor U442 (N_442,In_568,In_98);
xor U443 (N_443,In_327,In_726);
nand U444 (N_444,In_121,In_448);
nor U445 (N_445,In_253,In_638);
and U446 (N_446,In_134,In_457);
xnor U447 (N_447,In_706,In_381);
xor U448 (N_448,In_497,In_503);
and U449 (N_449,In_104,In_47);
xnor U450 (N_450,In_644,In_431);
nor U451 (N_451,In_587,In_668);
xor U452 (N_452,In_678,In_236);
and U453 (N_453,In_108,In_702);
xor U454 (N_454,In_607,In_656);
and U455 (N_455,In_71,In_279);
and U456 (N_456,In_532,In_286);
xor U457 (N_457,In_11,In_229);
xnor U458 (N_458,In_608,In_738);
or U459 (N_459,In_540,In_244);
nor U460 (N_460,In_688,In_220);
xnor U461 (N_461,In_332,In_299);
xnor U462 (N_462,In_223,In_599);
and U463 (N_463,In_412,In_502);
and U464 (N_464,In_731,In_509);
and U465 (N_465,In_537,In_686);
and U466 (N_466,In_472,In_325);
and U467 (N_467,In_346,In_629);
xor U468 (N_468,In_205,In_498);
nand U469 (N_469,In_356,In_95);
and U470 (N_470,In_383,In_228);
and U471 (N_471,In_660,In_393);
or U472 (N_472,In_724,In_162);
and U473 (N_473,In_379,In_4);
and U474 (N_474,In_353,In_20);
xnor U475 (N_475,In_44,In_100);
nand U476 (N_476,In_427,In_264);
nand U477 (N_477,In_223,In_735);
or U478 (N_478,In_367,In_649);
nor U479 (N_479,In_76,In_678);
or U480 (N_480,In_589,In_708);
and U481 (N_481,In_634,In_72);
xor U482 (N_482,In_264,In_60);
and U483 (N_483,In_28,In_141);
nor U484 (N_484,In_191,In_66);
nor U485 (N_485,In_602,In_388);
or U486 (N_486,In_639,In_196);
and U487 (N_487,In_192,In_274);
and U488 (N_488,In_512,In_516);
nor U489 (N_489,In_276,In_112);
or U490 (N_490,In_507,In_296);
nand U491 (N_491,In_580,In_334);
and U492 (N_492,In_62,In_5);
and U493 (N_493,In_190,In_548);
xnor U494 (N_494,In_618,In_46);
xor U495 (N_495,In_14,In_470);
nand U496 (N_496,In_168,In_685);
nand U497 (N_497,In_511,In_11);
or U498 (N_498,In_184,In_84);
nand U499 (N_499,In_32,In_189);
and U500 (N_500,In_136,In_568);
nand U501 (N_501,In_341,In_123);
and U502 (N_502,In_581,In_487);
nand U503 (N_503,In_626,In_454);
xnor U504 (N_504,In_212,In_247);
nand U505 (N_505,In_336,In_743);
xnor U506 (N_506,In_523,In_251);
nor U507 (N_507,In_146,In_605);
nor U508 (N_508,In_253,In_531);
xnor U509 (N_509,In_717,In_163);
or U510 (N_510,In_467,In_659);
nand U511 (N_511,In_732,In_209);
or U512 (N_512,In_580,In_7);
nor U513 (N_513,In_70,In_128);
xor U514 (N_514,In_50,In_287);
nor U515 (N_515,In_91,In_643);
xor U516 (N_516,In_161,In_618);
or U517 (N_517,In_315,In_61);
nor U518 (N_518,In_360,In_306);
nand U519 (N_519,In_205,In_173);
xor U520 (N_520,In_697,In_239);
and U521 (N_521,In_652,In_195);
nor U522 (N_522,In_318,In_607);
xor U523 (N_523,In_648,In_719);
or U524 (N_524,In_110,In_108);
xnor U525 (N_525,In_627,In_342);
nand U526 (N_526,In_612,In_694);
and U527 (N_527,In_355,In_170);
nor U528 (N_528,In_423,In_96);
and U529 (N_529,In_583,In_339);
nor U530 (N_530,In_247,In_259);
xor U531 (N_531,In_409,In_205);
and U532 (N_532,In_680,In_736);
xnor U533 (N_533,In_656,In_696);
xor U534 (N_534,In_576,In_261);
nor U535 (N_535,In_342,In_497);
and U536 (N_536,In_389,In_417);
nand U537 (N_537,In_44,In_527);
nor U538 (N_538,In_168,In_481);
or U539 (N_539,In_695,In_591);
and U540 (N_540,In_320,In_682);
xor U541 (N_541,In_87,In_359);
nand U542 (N_542,In_134,In_277);
or U543 (N_543,In_631,In_700);
xnor U544 (N_544,In_407,In_509);
nand U545 (N_545,In_247,In_80);
nand U546 (N_546,In_361,In_319);
or U547 (N_547,In_446,In_209);
nor U548 (N_548,In_741,In_172);
and U549 (N_549,In_204,In_526);
or U550 (N_550,In_375,In_327);
nor U551 (N_551,In_472,In_118);
nor U552 (N_552,In_664,In_373);
or U553 (N_553,In_296,In_494);
nor U554 (N_554,In_636,In_495);
nor U555 (N_555,In_354,In_630);
nand U556 (N_556,In_440,In_139);
nor U557 (N_557,In_422,In_642);
nand U558 (N_558,In_358,In_270);
nor U559 (N_559,In_330,In_309);
nor U560 (N_560,In_541,In_379);
nand U561 (N_561,In_627,In_500);
xor U562 (N_562,In_365,In_502);
nand U563 (N_563,In_253,In_197);
and U564 (N_564,In_156,In_47);
xnor U565 (N_565,In_586,In_139);
and U566 (N_566,In_201,In_180);
and U567 (N_567,In_387,In_663);
nor U568 (N_568,In_373,In_186);
nand U569 (N_569,In_449,In_594);
nor U570 (N_570,In_190,In_668);
nor U571 (N_571,In_170,In_267);
nor U572 (N_572,In_294,In_166);
xnor U573 (N_573,In_189,In_307);
xnor U574 (N_574,In_731,In_61);
nand U575 (N_575,In_232,In_687);
nand U576 (N_576,In_312,In_491);
xnor U577 (N_577,In_444,In_658);
or U578 (N_578,In_496,In_422);
nor U579 (N_579,In_675,In_548);
or U580 (N_580,In_219,In_661);
or U581 (N_581,In_50,In_229);
xor U582 (N_582,In_663,In_28);
xnor U583 (N_583,In_745,In_597);
or U584 (N_584,In_705,In_741);
or U585 (N_585,In_295,In_577);
or U586 (N_586,In_209,In_203);
nand U587 (N_587,In_361,In_186);
and U588 (N_588,In_107,In_196);
or U589 (N_589,In_8,In_631);
nand U590 (N_590,In_685,In_588);
xor U591 (N_591,In_210,In_168);
nand U592 (N_592,In_728,In_442);
nand U593 (N_593,In_30,In_120);
nor U594 (N_594,In_251,In_78);
nor U595 (N_595,In_574,In_202);
nand U596 (N_596,In_298,In_52);
xor U597 (N_597,In_321,In_576);
nor U598 (N_598,In_681,In_415);
or U599 (N_599,In_736,In_281);
nand U600 (N_600,In_52,In_267);
xnor U601 (N_601,In_423,In_133);
and U602 (N_602,In_579,In_348);
or U603 (N_603,In_731,In_598);
nor U604 (N_604,In_622,In_613);
xnor U605 (N_605,In_558,In_356);
xnor U606 (N_606,In_344,In_706);
or U607 (N_607,In_696,In_96);
nor U608 (N_608,In_484,In_194);
and U609 (N_609,In_158,In_254);
nand U610 (N_610,In_404,In_303);
or U611 (N_611,In_425,In_39);
nand U612 (N_612,In_598,In_73);
xor U613 (N_613,In_731,In_661);
or U614 (N_614,In_277,In_187);
or U615 (N_615,In_153,In_447);
and U616 (N_616,In_744,In_31);
nor U617 (N_617,In_733,In_302);
nor U618 (N_618,In_420,In_432);
nand U619 (N_619,In_704,In_489);
nand U620 (N_620,In_70,In_380);
and U621 (N_621,In_450,In_612);
and U622 (N_622,In_746,In_77);
nand U623 (N_623,In_226,In_666);
nor U624 (N_624,In_75,In_638);
nand U625 (N_625,In_305,In_72);
nand U626 (N_626,In_743,In_191);
or U627 (N_627,In_508,In_593);
nand U628 (N_628,In_642,In_583);
and U629 (N_629,In_292,In_255);
nand U630 (N_630,In_636,In_497);
xor U631 (N_631,In_180,In_326);
nand U632 (N_632,In_192,In_546);
nor U633 (N_633,In_655,In_154);
nor U634 (N_634,In_681,In_534);
or U635 (N_635,In_250,In_439);
or U636 (N_636,In_267,In_16);
nor U637 (N_637,In_46,In_326);
nor U638 (N_638,In_297,In_709);
xnor U639 (N_639,In_265,In_248);
nor U640 (N_640,In_287,In_381);
nor U641 (N_641,In_628,In_503);
nand U642 (N_642,In_361,In_363);
and U643 (N_643,In_325,In_385);
and U644 (N_644,In_488,In_330);
nand U645 (N_645,In_107,In_595);
nor U646 (N_646,In_166,In_342);
xnor U647 (N_647,In_197,In_307);
and U648 (N_648,In_132,In_71);
xnor U649 (N_649,In_530,In_396);
nor U650 (N_650,In_482,In_390);
xnor U651 (N_651,In_486,In_516);
or U652 (N_652,In_640,In_135);
nor U653 (N_653,In_185,In_650);
nor U654 (N_654,In_87,In_423);
nand U655 (N_655,In_252,In_127);
nand U656 (N_656,In_32,In_43);
nor U657 (N_657,In_198,In_280);
nor U658 (N_658,In_333,In_493);
or U659 (N_659,In_703,In_43);
nor U660 (N_660,In_557,In_273);
xor U661 (N_661,In_314,In_180);
nand U662 (N_662,In_629,In_437);
nand U663 (N_663,In_480,In_155);
xor U664 (N_664,In_646,In_268);
xnor U665 (N_665,In_229,In_184);
nor U666 (N_666,In_432,In_8);
xnor U667 (N_667,In_607,In_261);
xnor U668 (N_668,In_555,In_237);
nor U669 (N_669,In_446,In_517);
and U670 (N_670,In_225,In_388);
and U671 (N_671,In_679,In_607);
nor U672 (N_672,In_716,In_497);
or U673 (N_673,In_461,In_681);
or U674 (N_674,In_578,In_373);
nand U675 (N_675,In_525,In_135);
nand U676 (N_676,In_630,In_670);
xnor U677 (N_677,In_345,In_411);
or U678 (N_678,In_300,In_458);
and U679 (N_679,In_486,In_374);
or U680 (N_680,In_203,In_518);
nor U681 (N_681,In_440,In_239);
xor U682 (N_682,In_51,In_209);
nor U683 (N_683,In_137,In_458);
and U684 (N_684,In_574,In_442);
or U685 (N_685,In_172,In_235);
nand U686 (N_686,In_12,In_548);
nor U687 (N_687,In_366,In_90);
nor U688 (N_688,In_196,In_47);
xnor U689 (N_689,In_379,In_69);
nand U690 (N_690,In_561,In_457);
nand U691 (N_691,In_394,In_524);
nand U692 (N_692,In_167,In_268);
and U693 (N_693,In_562,In_447);
or U694 (N_694,In_313,In_708);
xnor U695 (N_695,In_428,In_659);
nand U696 (N_696,In_201,In_627);
xnor U697 (N_697,In_378,In_28);
and U698 (N_698,In_228,In_375);
or U699 (N_699,In_692,In_172);
xor U700 (N_700,In_71,In_631);
and U701 (N_701,In_636,In_432);
nand U702 (N_702,In_701,In_623);
and U703 (N_703,In_726,In_250);
or U704 (N_704,In_517,In_501);
or U705 (N_705,In_89,In_658);
xor U706 (N_706,In_316,In_199);
nand U707 (N_707,In_548,In_78);
or U708 (N_708,In_667,In_253);
nand U709 (N_709,In_634,In_397);
xor U710 (N_710,In_97,In_690);
nor U711 (N_711,In_428,In_570);
and U712 (N_712,In_11,In_121);
nand U713 (N_713,In_141,In_590);
nand U714 (N_714,In_408,In_182);
and U715 (N_715,In_616,In_473);
nor U716 (N_716,In_36,In_153);
and U717 (N_717,In_61,In_203);
xnor U718 (N_718,In_110,In_545);
or U719 (N_719,In_504,In_483);
xor U720 (N_720,In_317,In_600);
xnor U721 (N_721,In_85,In_596);
nor U722 (N_722,In_117,In_226);
and U723 (N_723,In_57,In_540);
nand U724 (N_724,In_470,In_329);
xor U725 (N_725,In_554,In_140);
xnor U726 (N_726,In_110,In_732);
or U727 (N_727,In_393,In_403);
and U728 (N_728,In_264,In_337);
nor U729 (N_729,In_512,In_409);
and U730 (N_730,In_514,In_283);
and U731 (N_731,In_453,In_478);
nand U732 (N_732,In_216,In_222);
nor U733 (N_733,In_305,In_335);
and U734 (N_734,In_548,In_215);
xor U735 (N_735,In_93,In_380);
nand U736 (N_736,In_123,In_626);
xor U737 (N_737,In_572,In_627);
and U738 (N_738,In_48,In_71);
xor U739 (N_739,In_249,In_687);
xnor U740 (N_740,In_567,In_465);
xnor U741 (N_741,In_465,In_133);
nand U742 (N_742,In_23,In_222);
xor U743 (N_743,In_669,In_613);
xor U744 (N_744,In_361,In_539);
nor U745 (N_745,In_245,In_547);
nor U746 (N_746,In_406,In_115);
nor U747 (N_747,In_218,In_689);
nor U748 (N_748,In_577,In_430);
and U749 (N_749,In_15,In_515);
nand U750 (N_750,In_419,In_454);
and U751 (N_751,In_269,In_161);
xor U752 (N_752,In_364,In_98);
and U753 (N_753,In_574,In_220);
and U754 (N_754,In_97,In_511);
and U755 (N_755,In_335,In_393);
nand U756 (N_756,In_59,In_483);
or U757 (N_757,In_480,In_439);
nor U758 (N_758,In_86,In_432);
and U759 (N_759,In_610,In_266);
or U760 (N_760,In_500,In_101);
or U761 (N_761,In_692,In_289);
and U762 (N_762,In_513,In_539);
nand U763 (N_763,In_564,In_278);
and U764 (N_764,In_572,In_357);
xor U765 (N_765,In_21,In_2);
or U766 (N_766,In_248,In_576);
or U767 (N_767,In_486,In_276);
or U768 (N_768,In_375,In_546);
and U769 (N_769,In_539,In_716);
and U770 (N_770,In_17,In_234);
and U771 (N_771,In_453,In_622);
xor U772 (N_772,In_603,In_739);
nor U773 (N_773,In_82,In_91);
nor U774 (N_774,In_430,In_601);
nand U775 (N_775,In_201,In_253);
xnor U776 (N_776,In_75,In_27);
nor U777 (N_777,In_400,In_77);
or U778 (N_778,In_223,In_312);
xnor U779 (N_779,In_384,In_219);
nor U780 (N_780,In_254,In_532);
nor U781 (N_781,In_532,In_361);
nand U782 (N_782,In_250,In_358);
xnor U783 (N_783,In_297,In_80);
nor U784 (N_784,In_687,In_121);
nand U785 (N_785,In_111,In_441);
and U786 (N_786,In_542,In_661);
and U787 (N_787,In_246,In_570);
and U788 (N_788,In_65,In_610);
nand U789 (N_789,In_100,In_686);
or U790 (N_790,In_405,In_591);
xor U791 (N_791,In_378,In_300);
and U792 (N_792,In_125,In_307);
nand U793 (N_793,In_581,In_208);
nand U794 (N_794,In_545,In_153);
and U795 (N_795,In_333,In_563);
xnor U796 (N_796,In_313,In_290);
xnor U797 (N_797,In_358,In_729);
nand U798 (N_798,In_65,In_490);
nand U799 (N_799,In_9,In_211);
nand U800 (N_800,In_80,In_701);
or U801 (N_801,In_349,In_352);
nand U802 (N_802,In_671,In_528);
and U803 (N_803,In_290,In_590);
nand U804 (N_804,In_225,In_737);
xnor U805 (N_805,In_640,In_736);
nor U806 (N_806,In_187,In_119);
xnor U807 (N_807,In_165,In_462);
nor U808 (N_808,In_90,In_201);
nand U809 (N_809,In_140,In_317);
nor U810 (N_810,In_77,In_219);
nor U811 (N_811,In_431,In_82);
and U812 (N_812,In_15,In_242);
nand U813 (N_813,In_179,In_455);
and U814 (N_814,In_571,In_280);
nor U815 (N_815,In_185,In_735);
xnor U816 (N_816,In_659,In_158);
nand U817 (N_817,In_385,In_679);
nand U818 (N_818,In_619,In_320);
and U819 (N_819,In_651,In_569);
or U820 (N_820,In_311,In_699);
or U821 (N_821,In_323,In_70);
xor U822 (N_822,In_221,In_675);
or U823 (N_823,In_244,In_640);
nor U824 (N_824,In_158,In_157);
nor U825 (N_825,In_164,In_420);
nor U826 (N_826,In_191,In_688);
xor U827 (N_827,In_41,In_555);
xor U828 (N_828,In_193,In_502);
xnor U829 (N_829,In_662,In_651);
nor U830 (N_830,In_72,In_607);
or U831 (N_831,In_618,In_434);
or U832 (N_832,In_218,In_462);
or U833 (N_833,In_635,In_3);
nand U834 (N_834,In_79,In_381);
xor U835 (N_835,In_305,In_378);
or U836 (N_836,In_386,In_736);
nor U837 (N_837,In_132,In_181);
or U838 (N_838,In_238,In_383);
nor U839 (N_839,In_583,In_80);
or U840 (N_840,In_471,In_382);
nor U841 (N_841,In_691,In_288);
nand U842 (N_842,In_320,In_351);
nor U843 (N_843,In_538,In_651);
and U844 (N_844,In_39,In_313);
and U845 (N_845,In_321,In_504);
and U846 (N_846,In_495,In_731);
and U847 (N_847,In_722,In_303);
or U848 (N_848,In_224,In_227);
nor U849 (N_849,In_576,In_499);
xnor U850 (N_850,In_615,In_240);
or U851 (N_851,In_662,In_444);
or U852 (N_852,In_707,In_164);
and U853 (N_853,In_489,In_406);
nand U854 (N_854,In_511,In_266);
and U855 (N_855,In_186,In_457);
nand U856 (N_856,In_170,In_407);
nor U857 (N_857,In_94,In_379);
xor U858 (N_858,In_281,In_323);
and U859 (N_859,In_466,In_271);
nor U860 (N_860,In_320,In_379);
and U861 (N_861,In_233,In_325);
and U862 (N_862,In_105,In_637);
nor U863 (N_863,In_680,In_720);
nand U864 (N_864,In_571,In_82);
and U865 (N_865,In_567,In_191);
nand U866 (N_866,In_458,In_79);
xnor U867 (N_867,In_502,In_178);
and U868 (N_868,In_473,In_748);
xor U869 (N_869,In_535,In_509);
nor U870 (N_870,In_111,In_398);
or U871 (N_871,In_487,In_301);
xnor U872 (N_872,In_673,In_400);
or U873 (N_873,In_716,In_234);
or U874 (N_874,In_642,In_270);
nand U875 (N_875,In_707,In_49);
or U876 (N_876,In_515,In_352);
or U877 (N_877,In_673,In_277);
and U878 (N_878,In_0,In_143);
nor U879 (N_879,In_196,In_65);
and U880 (N_880,In_232,In_434);
nand U881 (N_881,In_701,In_596);
xor U882 (N_882,In_61,In_232);
or U883 (N_883,In_638,In_315);
nand U884 (N_884,In_431,In_223);
nor U885 (N_885,In_124,In_572);
nand U886 (N_886,In_657,In_649);
nand U887 (N_887,In_184,In_36);
nor U888 (N_888,In_377,In_492);
or U889 (N_889,In_595,In_273);
nand U890 (N_890,In_541,In_742);
or U891 (N_891,In_159,In_520);
or U892 (N_892,In_116,In_18);
nand U893 (N_893,In_237,In_745);
or U894 (N_894,In_304,In_687);
nor U895 (N_895,In_474,In_636);
nor U896 (N_896,In_446,In_571);
or U897 (N_897,In_350,In_319);
or U898 (N_898,In_140,In_28);
or U899 (N_899,In_706,In_136);
xnor U900 (N_900,In_192,In_87);
nor U901 (N_901,In_477,In_219);
nand U902 (N_902,In_665,In_474);
nor U903 (N_903,In_705,In_292);
or U904 (N_904,In_714,In_90);
nor U905 (N_905,In_314,In_718);
nand U906 (N_906,In_46,In_703);
or U907 (N_907,In_337,In_524);
or U908 (N_908,In_311,In_683);
nand U909 (N_909,In_372,In_557);
and U910 (N_910,In_13,In_97);
or U911 (N_911,In_346,In_532);
xor U912 (N_912,In_693,In_647);
or U913 (N_913,In_28,In_603);
and U914 (N_914,In_345,In_733);
and U915 (N_915,In_650,In_116);
and U916 (N_916,In_161,In_425);
or U917 (N_917,In_341,In_266);
nand U918 (N_918,In_596,In_722);
and U919 (N_919,In_464,In_213);
and U920 (N_920,In_51,In_734);
nor U921 (N_921,In_79,In_298);
nor U922 (N_922,In_72,In_81);
and U923 (N_923,In_499,In_593);
xor U924 (N_924,In_142,In_370);
nor U925 (N_925,In_506,In_53);
or U926 (N_926,In_32,In_656);
nor U927 (N_927,In_423,In_35);
nor U928 (N_928,In_432,In_253);
nand U929 (N_929,In_659,In_105);
nand U930 (N_930,In_352,In_37);
or U931 (N_931,In_434,In_520);
xor U932 (N_932,In_657,In_635);
or U933 (N_933,In_47,In_74);
and U934 (N_934,In_570,In_476);
and U935 (N_935,In_418,In_293);
and U936 (N_936,In_535,In_267);
nor U937 (N_937,In_168,In_139);
nor U938 (N_938,In_246,In_263);
nor U939 (N_939,In_236,In_163);
nor U940 (N_940,In_701,In_529);
nand U941 (N_941,In_84,In_182);
and U942 (N_942,In_107,In_441);
nor U943 (N_943,In_125,In_475);
xor U944 (N_944,In_463,In_562);
or U945 (N_945,In_716,In_586);
nor U946 (N_946,In_147,In_221);
nor U947 (N_947,In_463,In_40);
or U948 (N_948,In_2,In_632);
xor U949 (N_949,In_22,In_109);
or U950 (N_950,In_252,In_446);
nand U951 (N_951,In_610,In_200);
or U952 (N_952,In_487,In_268);
xnor U953 (N_953,In_140,In_118);
nor U954 (N_954,In_167,In_77);
or U955 (N_955,In_324,In_14);
and U956 (N_956,In_574,In_593);
nor U957 (N_957,In_195,In_723);
xnor U958 (N_958,In_134,In_338);
or U959 (N_959,In_445,In_300);
or U960 (N_960,In_51,In_742);
nand U961 (N_961,In_589,In_487);
nor U962 (N_962,In_334,In_84);
nand U963 (N_963,In_705,In_359);
nand U964 (N_964,In_532,In_503);
xnor U965 (N_965,In_95,In_158);
nor U966 (N_966,In_71,In_519);
nor U967 (N_967,In_197,In_418);
and U968 (N_968,In_519,In_332);
xnor U969 (N_969,In_127,In_504);
nor U970 (N_970,In_396,In_390);
nand U971 (N_971,In_273,In_153);
or U972 (N_972,In_34,In_195);
nand U973 (N_973,In_413,In_189);
xnor U974 (N_974,In_173,In_326);
nand U975 (N_975,In_186,In_631);
nor U976 (N_976,In_465,In_40);
or U977 (N_977,In_605,In_8);
or U978 (N_978,In_196,In_367);
nand U979 (N_979,In_572,In_553);
or U980 (N_980,In_2,In_732);
and U981 (N_981,In_454,In_204);
nand U982 (N_982,In_578,In_575);
nand U983 (N_983,In_162,In_527);
xor U984 (N_984,In_469,In_21);
or U985 (N_985,In_329,In_535);
and U986 (N_986,In_684,In_579);
and U987 (N_987,In_178,In_149);
xnor U988 (N_988,In_55,In_241);
or U989 (N_989,In_313,In_501);
xnor U990 (N_990,In_412,In_426);
xnor U991 (N_991,In_540,In_492);
and U992 (N_992,In_296,In_497);
nand U993 (N_993,In_162,In_498);
xor U994 (N_994,In_305,In_386);
nor U995 (N_995,In_127,In_616);
nor U996 (N_996,In_116,In_220);
xnor U997 (N_997,In_173,In_614);
nor U998 (N_998,In_464,In_43);
nor U999 (N_999,In_508,In_726);
and U1000 (N_1000,N_857,N_578);
nand U1001 (N_1001,N_950,N_866);
nand U1002 (N_1002,N_860,N_848);
nor U1003 (N_1003,N_703,N_14);
or U1004 (N_1004,N_934,N_689);
nand U1005 (N_1005,N_184,N_981);
nor U1006 (N_1006,N_850,N_448);
and U1007 (N_1007,N_832,N_759);
and U1008 (N_1008,N_326,N_342);
or U1009 (N_1009,N_157,N_491);
nor U1010 (N_1010,N_162,N_956);
nor U1011 (N_1011,N_800,N_944);
or U1012 (N_1012,N_435,N_732);
or U1013 (N_1013,N_922,N_373);
nand U1014 (N_1014,N_280,N_180);
nand U1015 (N_1015,N_138,N_331);
xnor U1016 (N_1016,N_170,N_63);
or U1017 (N_1017,N_838,N_34);
and U1018 (N_1018,N_856,N_243);
or U1019 (N_1019,N_671,N_796);
nand U1020 (N_1020,N_720,N_781);
or U1021 (N_1021,N_707,N_534);
xor U1022 (N_1022,N_805,N_666);
nand U1023 (N_1023,N_196,N_382);
and U1024 (N_1024,N_760,N_190);
xor U1025 (N_1025,N_13,N_388);
or U1026 (N_1026,N_762,N_947);
nand U1027 (N_1027,N_892,N_692);
nand U1028 (N_1028,N_715,N_824);
or U1029 (N_1029,N_94,N_937);
and U1030 (N_1030,N_614,N_723);
and U1031 (N_1031,N_428,N_785);
nand U1032 (N_1032,N_989,N_312);
nor U1033 (N_1033,N_98,N_7);
and U1034 (N_1034,N_545,N_438);
nand U1035 (N_1035,N_230,N_849);
or U1036 (N_1036,N_179,N_322);
nand U1037 (N_1037,N_282,N_885);
nand U1038 (N_1038,N_697,N_275);
nand U1039 (N_1039,N_154,N_651);
nor U1040 (N_1040,N_815,N_175);
and U1041 (N_1041,N_134,N_659);
xnor U1042 (N_1042,N_353,N_470);
nor U1043 (N_1043,N_831,N_35);
xor U1044 (N_1044,N_617,N_683);
nand U1045 (N_1045,N_258,N_276);
and U1046 (N_1046,N_851,N_682);
xor U1047 (N_1047,N_270,N_194);
xor U1048 (N_1048,N_924,N_816);
nor U1049 (N_1049,N_278,N_539);
nor U1050 (N_1050,N_586,N_132);
nor U1051 (N_1051,N_888,N_693);
and U1052 (N_1052,N_57,N_163);
and U1053 (N_1053,N_558,N_395);
or U1054 (N_1054,N_834,N_728);
and U1055 (N_1055,N_262,N_434);
nor U1056 (N_1056,N_630,N_12);
and U1057 (N_1057,N_323,N_488);
or U1058 (N_1058,N_917,N_389);
nor U1059 (N_1059,N_699,N_110);
or U1060 (N_1060,N_891,N_200);
xor U1061 (N_1061,N_199,N_847);
xnor U1062 (N_1062,N_463,N_955);
and U1063 (N_1063,N_468,N_719);
or U1064 (N_1064,N_115,N_637);
and U1065 (N_1065,N_263,N_725);
or U1066 (N_1066,N_487,N_220);
nand U1067 (N_1067,N_537,N_355);
nor U1068 (N_1068,N_321,N_650);
or U1069 (N_1069,N_881,N_293);
nor U1070 (N_1070,N_979,N_198);
and U1071 (N_1071,N_807,N_325);
nor U1072 (N_1072,N_510,N_421);
xor U1073 (N_1073,N_880,N_144);
and U1074 (N_1074,N_764,N_928);
nor U1075 (N_1075,N_563,N_372);
nand U1076 (N_1076,N_155,N_919);
nor U1077 (N_1077,N_392,N_700);
or U1078 (N_1078,N_416,N_381);
and U1079 (N_1079,N_23,N_767);
nor U1080 (N_1080,N_574,N_16);
and U1081 (N_1081,N_73,N_643);
xnor U1082 (N_1082,N_593,N_843);
nor U1083 (N_1083,N_11,N_446);
nor U1084 (N_1084,N_247,N_481);
nor U1085 (N_1085,N_338,N_62);
nand U1086 (N_1086,N_566,N_898);
and U1087 (N_1087,N_511,N_945);
nor U1088 (N_1088,N_791,N_123);
or U1089 (N_1089,N_313,N_384);
or U1090 (N_1090,N_525,N_730);
xnor U1091 (N_1091,N_758,N_902);
or U1092 (N_1092,N_768,N_639);
and U1093 (N_1093,N_973,N_641);
nand U1094 (N_1094,N_610,N_80);
and U1095 (N_1095,N_826,N_647);
or U1096 (N_1096,N_237,N_827);
and U1097 (N_1097,N_646,N_743);
xnor U1098 (N_1098,N_629,N_192);
nor U1099 (N_1099,N_225,N_420);
nor U1100 (N_1100,N_786,N_54);
xor U1101 (N_1101,N_158,N_436);
nand U1102 (N_1102,N_904,N_377);
nor U1103 (N_1103,N_273,N_959);
xnor U1104 (N_1104,N_227,N_32);
and U1105 (N_1105,N_334,N_884);
nor U1106 (N_1106,N_606,N_571);
or U1107 (N_1107,N_980,N_361);
and U1108 (N_1108,N_966,N_588);
nand U1109 (N_1109,N_311,N_479);
nand U1110 (N_1110,N_889,N_560);
nor U1111 (N_1111,N_211,N_212);
nand U1112 (N_1112,N_231,N_242);
nor U1113 (N_1113,N_958,N_665);
nor U1114 (N_1114,N_579,N_315);
xnor U1115 (N_1115,N_925,N_940);
xor U1116 (N_1116,N_971,N_234);
and U1117 (N_1117,N_855,N_741);
and U1118 (N_1118,N_385,N_363);
and U1119 (N_1119,N_718,N_601);
xor U1120 (N_1120,N_969,N_239);
nor U1121 (N_1121,N_336,N_986);
and U1122 (N_1122,N_532,N_267);
or U1123 (N_1123,N_48,N_277);
nand U1124 (N_1124,N_52,N_96);
or U1125 (N_1125,N_508,N_406);
xor U1126 (N_1126,N_489,N_21);
or U1127 (N_1127,N_150,N_79);
and U1128 (N_1128,N_790,N_660);
nor U1129 (N_1129,N_708,N_870);
and U1130 (N_1130,N_688,N_84);
nor U1131 (N_1131,N_260,N_905);
and U1132 (N_1132,N_181,N_77);
or U1133 (N_1133,N_414,N_747);
nor U1134 (N_1134,N_983,N_201);
or U1135 (N_1135,N_871,N_422);
and U1136 (N_1136,N_913,N_256);
or U1137 (N_1137,N_172,N_612);
xnor U1138 (N_1138,N_356,N_36);
xor U1139 (N_1139,N_121,N_946);
or U1140 (N_1140,N_654,N_27);
and U1141 (N_1141,N_24,N_452);
or U1142 (N_1142,N_307,N_66);
xnor U1143 (N_1143,N_426,N_444);
nor U1144 (N_1144,N_920,N_773);
nand U1145 (N_1145,N_254,N_314);
or U1146 (N_1146,N_478,N_100);
nor U1147 (N_1147,N_921,N_352);
xnor U1148 (N_1148,N_357,N_466);
or U1149 (N_1149,N_561,N_923);
or U1150 (N_1150,N_454,N_842);
xnor U1151 (N_1151,N_864,N_521);
nor U1152 (N_1152,N_771,N_85);
xor U1153 (N_1153,N_653,N_543);
xor U1154 (N_1154,N_664,N_555);
nor U1155 (N_1155,N_530,N_792);
or U1156 (N_1156,N_710,N_205);
nand U1157 (N_1157,N_840,N_202);
and U1158 (N_1158,N_61,N_400);
nand U1159 (N_1159,N_104,N_41);
and U1160 (N_1160,N_476,N_717);
xor U1161 (N_1161,N_679,N_109);
and U1162 (N_1162,N_367,N_240);
nor U1163 (N_1163,N_210,N_872);
nor U1164 (N_1164,N_960,N_456);
xnor U1165 (N_1165,N_813,N_365);
and U1166 (N_1166,N_713,N_823);
xnor U1167 (N_1167,N_701,N_462);
and U1168 (N_1168,N_284,N_948);
or U1169 (N_1169,N_592,N_82);
nand U1170 (N_1170,N_497,N_235);
or U1171 (N_1171,N_675,N_59);
or U1172 (N_1172,N_161,N_618);
xnor U1173 (N_1173,N_250,N_982);
or U1174 (N_1174,N_101,N_988);
xor U1175 (N_1175,N_90,N_658);
nand U1176 (N_1176,N_535,N_599);
or U1177 (N_1177,N_129,N_999);
xor U1178 (N_1178,N_663,N_223);
and U1179 (N_1179,N_87,N_895);
nor U1180 (N_1180,N_597,N_569);
and U1181 (N_1181,N_345,N_108);
nand U1182 (N_1182,N_894,N_266);
or U1183 (N_1183,N_89,N_329);
nand U1184 (N_1184,N_442,N_573);
nand U1185 (N_1185,N_246,N_137);
xnor U1186 (N_1186,N_424,N_493);
nand U1187 (N_1187,N_33,N_828);
or U1188 (N_1188,N_327,N_549);
xnor U1189 (N_1189,N_749,N_348);
nor U1190 (N_1190,N_770,N_289);
nand U1191 (N_1191,N_1,N_961);
nor U1192 (N_1192,N_794,N_261);
nand U1193 (N_1193,N_954,N_975);
nor U1194 (N_1194,N_594,N_580);
or U1195 (N_1195,N_241,N_430);
xor U1196 (N_1196,N_590,N_705);
xnor U1197 (N_1197,N_298,N_990);
nand U1198 (N_1198,N_685,N_929);
nor U1199 (N_1199,N_547,N_645);
nand U1200 (N_1200,N_469,N_187);
or U1201 (N_1201,N_711,N_538);
or U1202 (N_1202,N_686,N_425);
nor U1203 (N_1203,N_203,N_145);
nand U1204 (N_1204,N_727,N_712);
or U1205 (N_1205,N_938,N_358);
nor U1206 (N_1206,N_626,N_271);
nand U1207 (N_1207,N_486,N_837);
and U1208 (N_1208,N_97,N_912);
and U1209 (N_1209,N_998,N_964);
nand U1210 (N_1210,N_908,N_795);
xor U1211 (N_1211,N_195,N_787);
xor U1212 (N_1212,N_30,N_903);
nand U1213 (N_1213,N_518,N_118);
and U1214 (N_1214,N_765,N_788);
xor U1215 (N_1215,N_568,N_412);
or U1216 (N_1216,N_789,N_304);
and U1217 (N_1217,N_53,N_106);
or U1218 (N_1218,N_427,N_621);
nor U1219 (N_1219,N_88,N_159);
and U1220 (N_1220,N_253,N_778);
and U1221 (N_1221,N_333,N_402);
xnor U1222 (N_1222,N_25,N_483);
xor U1223 (N_1223,N_405,N_459);
nand U1224 (N_1224,N_825,N_143);
nand U1225 (N_1225,N_836,N_577);
or U1226 (N_1226,N_802,N_776);
and U1227 (N_1227,N_350,N_680);
or U1228 (N_1228,N_429,N_74);
nor U1229 (N_1229,N_15,N_656);
or U1230 (N_1230,N_167,N_523);
nand U1231 (N_1231,N_165,N_480);
nor U1232 (N_1232,N_224,N_985);
and U1233 (N_1233,N_193,N_953);
nor U1234 (N_1234,N_615,N_733);
xor U1235 (N_1235,N_113,N_29);
nor U1236 (N_1236,N_6,N_499);
nor U1237 (N_1237,N_809,N_997);
or U1238 (N_1238,N_572,N_441);
and U1239 (N_1239,N_18,N_642);
xnor U1240 (N_1240,N_835,N_139);
and U1241 (N_1241,N_461,N_166);
and U1242 (N_1242,N_565,N_632);
or U1243 (N_1243,N_620,N_644);
or U1244 (N_1244,N_55,N_761);
and U1245 (N_1245,N_214,N_821);
nor U1246 (N_1246,N_248,N_360);
and U1247 (N_1247,N_337,N_56);
xor U1248 (N_1248,N_8,N_575);
and U1249 (N_1249,N_379,N_957);
and U1250 (N_1250,N_506,N_418);
nor U1251 (N_1251,N_213,N_858);
nand U1252 (N_1252,N_37,N_783);
or U1253 (N_1253,N_745,N_634);
and U1254 (N_1254,N_140,N_542);
xor U1255 (N_1255,N_259,N_882);
xor U1256 (N_1256,N_152,N_351);
or U1257 (N_1257,N_43,N_411);
nand U1258 (N_1258,N_176,N_678);
xor U1259 (N_1259,N_739,N_942);
nor U1260 (N_1260,N_546,N_20);
and U1261 (N_1261,N_359,N_171);
nor U1262 (N_1262,N_527,N_292);
or U1263 (N_1263,N_684,N_513);
nor U1264 (N_1264,N_676,N_591);
nor U1265 (N_1265,N_460,N_736);
xor U1266 (N_1266,N_443,N_726);
and U1267 (N_1267,N_978,N_553);
and U1268 (N_1268,N_817,N_151);
and U1269 (N_1269,N_702,N_433);
xor U1270 (N_1270,N_26,N_368);
nor U1271 (N_1271,N_729,N_375);
nor U1272 (N_1272,N_896,N_657);
nand U1273 (N_1273,N_541,N_288);
xnor U1274 (N_1274,N_440,N_740);
nor U1275 (N_1275,N_906,N_445);
xor U1276 (N_1276,N_987,N_854);
xor U1277 (N_1277,N_9,N_99);
or U1278 (N_1278,N_548,N_965);
nand U1279 (N_1279,N_91,N_907);
or U1280 (N_1280,N_775,N_305);
and U1281 (N_1281,N_387,N_584);
or U1282 (N_1282,N_244,N_124);
and U1283 (N_1283,N_183,N_316);
nor U1284 (N_1284,N_232,N_169);
and U1285 (N_1285,N_559,N_3);
xnor U1286 (N_1286,N_408,N_674);
nor U1287 (N_1287,N_690,N_667);
xor U1288 (N_1288,N_394,N_536);
or U1289 (N_1289,N_627,N_399);
nand U1290 (N_1290,N_482,N_780);
nand U1291 (N_1291,N_886,N_799);
xnor U1292 (N_1292,N_691,N_803);
nand U1293 (N_1293,N_339,N_300);
nor U1294 (N_1294,N_302,N_735);
xor U1295 (N_1295,N_581,N_984);
and U1296 (N_1296,N_128,N_622);
xnor U1297 (N_1297,N_371,N_714);
nand U1298 (N_1298,N_994,N_92);
or U1299 (N_1299,N_931,N_731);
nand U1300 (N_1300,N_233,N_763);
xnor U1301 (N_1301,N_380,N_869);
nand U1302 (N_1302,N_819,N_833);
nor U1303 (N_1303,N_524,N_296);
xor U1304 (N_1304,N_17,N_505);
and U1305 (N_1305,N_301,N_141);
and U1306 (N_1306,N_793,N_127);
nor U1307 (N_1307,N_209,N_133);
nand U1308 (N_1308,N_38,N_533);
and U1309 (N_1309,N_431,N_204);
and U1310 (N_1310,N_142,N_306);
nor U1311 (N_1311,N_228,N_734);
nor U1312 (N_1312,N_933,N_83);
or U1313 (N_1313,N_515,N_75);
or U1314 (N_1314,N_309,N_189);
or U1315 (N_1315,N_766,N_669);
or U1316 (N_1316,N_269,N_107);
or U1317 (N_1317,N_409,N_413);
nand U1318 (N_1318,N_564,N_318);
xnor U1319 (N_1319,N_863,N_50);
and U1320 (N_1320,N_782,N_504);
xor U1321 (N_1321,N_294,N_281);
and U1322 (N_1322,N_512,N_976);
and U1323 (N_1323,N_208,N_619);
and U1324 (N_1324,N_910,N_86);
and U1325 (N_1325,N_81,N_68);
and U1326 (N_1326,N_498,N_774);
nor U1327 (N_1327,N_219,N_485);
xor U1328 (N_1328,N_932,N_393);
and U1329 (N_1329,N_494,N_319);
and U1330 (N_1330,N_191,N_149);
nand U1331 (N_1331,N_875,N_28);
xor U1332 (N_1332,N_297,N_22);
or U1333 (N_1333,N_616,N_814);
or U1334 (N_1334,N_844,N_522);
nor U1335 (N_1335,N_661,N_977);
or U1336 (N_1336,N_467,N_595);
nor U1337 (N_1337,N_188,N_40);
and U1338 (N_1338,N_681,N_598);
or U1339 (N_1339,N_148,N_677);
or U1340 (N_1340,N_335,N_173);
nor U1341 (N_1341,N_818,N_245);
and U1342 (N_1342,N_624,N_829);
or U1343 (N_1343,N_500,N_706);
nor U1344 (N_1344,N_221,N_39);
nor U1345 (N_1345,N_119,N_364);
and U1346 (N_1346,N_197,N_911);
and U1347 (N_1347,N_943,N_502);
and U1348 (N_1348,N_19,N_673);
and U1349 (N_1349,N_517,N_631);
xnor U1350 (N_1350,N_777,N_608);
nand U1351 (N_1351,N_879,N_737);
and U1352 (N_1352,N_804,N_878);
nand U1353 (N_1353,N_70,N_583);
xor U1354 (N_1354,N_520,N_72);
or U1355 (N_1355,N_962,N_628);
xor U1356 (N_1356,N_808,N_635);
and U1357 (N_1357,N_320,N_168);
nand U1358 (N_1358,N_604,N_238);
nor U1359 (N_1359,N_529,N_995);
and U1360 (N_1360,N_963,N_970);
nand U1361 (N_1361,N_2,N_822);
nor U1362 (N_1362,N_528,N_477);
nand U1363 (N_1363,N_410,N_153);
nand U1364 (N_1364,N_640,N_374);
nor U1365 (N_1365,N_274,N_589);
nand U1366 (N_1366,N_285,N_10);
or U1367 (N_1367,N_51,N_146);
and U1368 (N_1368,N_576,N_845);
and U1369 (N_1369,N_865,N_993);
nor U1370 (N_1370,N_694,N_5);
xor U1371 (N_1371,N_102,N_755);
or U1372 (N_1372,N_544,N_974);
and U1373 (N_1373,N_890,N_696);
and U1374 (N_1374,N_362,N_967);
xor U1375 (N_1375,N_972,N_883);
xor U1376 (N_1376,N_936,N_812);
or U1377 (N_1377,N_117,N_229);
nor U1378 (N_1378,N_861,N_797);
nor U1379 (N_1379,N_69,N_396);
and U1380 (N_1380,N_893,N_286);
and U1381 (N_1381,N_397,N_317);
xnor U1382 (N_1382,N_58,N_160);
nand U1383 (N_1383,N_147,N_779);
xor U1384 (N_1384,N_437,N_207);
nor U1385 (N_1385,N_806,N_346);
or U1386 (N_1386,N_876,N_603);
nand U1387 (N_1387,N_432,N_724);
nor U1388 (N_1388,N_217,N_668);
nand U1389 (N_1389,N_670,N_407);
nand U1390 (N_1390,N_332,N_968);
and U1391 (N_1391,N_841,N_746);
nor U1392 (N_1392,N_687,N_449);
nand U1393 (N_1393,N_268,N_655);
or U1394 (N_1394,N_474,N_596);
nor U1395 (N_1395,N_226,N_76);
nor U1396 (N_1396,N_709,N_567);
or U1397 (N_1397,N_447,N_941);
nand U1398 (N_1398,N_704,N_376);
nand U1399 (N_1399,N_215,N_42);
nor U1400 (N_1400,N_695,N_272);
or U1401 (N_1401,N_939,N_114);
or U1402 (N_1402,N_992,N_185);
or U1403 (N_1403,N_453,N_756);
nor U1404 (N_1404,N_607,N_49);
nor U1405 (N_1405,N_31,N_415);
nor U1406 (N_1406,N_265,N_859);
and U1407 (N_1407,N_310,N_283);
or U1408 (N_1408,N_531,N_784);
and U1409 (N_1409,N_417,N_526);
nor U1410 (N_1410,N_926,N_633);
and U1411 (N_1411,N_472,N_811);
xor U1412 (N_1412,N_0,N_330);
and U1413 (N_1413,N_750,N_93);
and U1414 (N_1414,N_909,N_839);
xnor U1415 (N_1415,N_473,N_798);
xnor U1416 (N_1416,N_570,N_439);
nor U1417 (N_1417,N_495,N_308);
or U1418 (N_1418,N_206,N_503);
xnor U1419 (N_1419,N_398,N_949);
and U1420 (N_1420,N_914,N_540);
or U1421 (N_1421,N_501,N_877);
nand U1422 (N_1422,N_514,N_125);
and U1423 (N_1423,N_44,N_550);
and U1424 (N_1424,N_419,N_742);
or U1425 (N_1425,N_722,N_164);
and U1426 (N_1426,N_116,N_873);
or U1427 (N_1427,N_105,N_952);
or U1428 (N_1428,N_457,N_757);
xor U1429 (N_1429,N_874,N_136);
or U1430 (N_1430,N_343,N_178);
and U1431 (N_1431,N_602,N_554);
xnor U1432 (N_1432,N_458,N_383);
nor U1433 (N_1433,N_830,N_901);
nor U1434 (N_1434,N_930,N_662);
nor U1435 (N_1435,N_551,N_174);
or U1436 (N_1436,N_636,N_404);
nand U1437 (N_1437,N_111,N_216);
nand U1438 (N_1438,N_78,N_291);
xor U1439 (N_1439,N_915,N_218);
nand U1440 (N_1440,N_252,N_386);
or U1441 (N_1441,N_744,N_186);
nand U1442 (N_1442,N_279,N_484);
nand U1443 (N_1443,N_853,N_369);
xnor U1444 (N_1444,N_638,N_611);
xnor U1445 (N_1445,N_698,N_585);
nand U1446 (N_1446,N_126,N_465);
nor U1447 (N_1447,N_182,N_716);
and U1448 (N_1448,N_71,N_623);
nor U1449 (N_1449,N_290,N_423);
or U1450 (N_1450,N_347,N_354);
xnor U1451 (N_1451,N_918,N_65);
nand U1452 (N_1452,N_156,N_370);
nand U1453 (N_1453,N_47,N_769);
xor U1454 (N_1454,N_738,N_401);
and U1455 (N_1455,N_609,N_236);
and U1456 (N_1456,N_344,N_600);
nand U1457 (N_1457,N_935,N_341);
nor U1458 (N_1458,N_519,N_112);
xor U1459 (N_1459,N_900,N_868);
or U1460 (N_1460,N_862,N_255);
or U1461 (N_1461,N_130,N_135);
or U1462 (N_1462,N_4,N_852);
nor U1463 (N_1463,N_927,N_67);
nand U1464 (N_1464,N_45,N_328);
or U1465 (N_1465,N_257,N_122);
nand U1466 (N_1466,N_748,N_349);
or U1467 (N_1467,N_672,N_303);
and U1468 (N_1468,N_652,N_587);
nand U1469 (N_1469,N_507,N_492);
xor U1470 (N_1470,N_649,N_801);
nand U1471 (N_1471,N_95,N_772);
xnor U1472 (N_1472,N_562,N_991);
nand U1473 (N_1473,N_496,N_390);
nand U1474 (N_1474,N_120,N_752);
xnor U1475 (N_1475,N_475,N_340);
nor U1476 (N_1476,N_820,N_846);
nand U1477 (N_1477,N_299,N_897);
and U1478 (N_1478,N_324,N_509);
xnor U1479 (N_1479,N_625,N_287);
nand U1480 (N_1480,N_648,N_556);
nand U1481 (N_1481,N_251,N_249);
nand U1482 (N_1482,N_378,N_60);
xor U1483 (N_1483,N_916,N_613);
nand U1484 (N_1484,N_403,N_177);
nor U1485 (N_1485,N_450,N_582);
xor U1486 (N_1486,N_996,N_464);
nand U1487 (N_1487,N_867,N_64);
and U1488 (N_1488,N_899,N_751);
nor U1489 (N_1489,N_887,N_366);
or U1490 (N_1490,N_810,N_552);
nand U1491 (N_1491,N_605,N_951);
nor U1492 (N_1492,N_490,N_131);
nand U1493 (N_1493,N_753,N_103);
or U1494 (N_1494,N_754,N_471);
nand U1495 (N_1495,N_455,N_222);
nor U1496 (N_1496,N_721,N_451);
or U1497 (N_1497,N_264,N_516);
nand U1498 (N_1498,N_295,N_391);
nor U1499 (N_1499,N_46,N_557);
nor U1500 (N_1500,N_645,N_828);
xnor U1501 (N_1501,N_251,N_236);
nor U1502 (N_1502,N_270,N_650);
xnor U1503 (N_1503,N_693,N_108);
nand U1504 (N_1504,N_683,N_158);
and U1505 (N_1505,N_159,N_539);
nor U1506 (N_1506,N_458,N_576);
nor U1507 (N_1507,N_315,N_240);
xnor U1508 (N_1508,N_7,N_205);
or U1509 (N_1509,N_866,N_734);
xnor U1510 (N_1510,N_421,N_64);
or U1511 (N_1511,N_8,N_881);
nor U1512 (N_1512,N_275,N_557);
nor U1513 (N_1513,N_695,N_334);
xnor U1514 (N_1514,N_779,N_580);
xor U1515 (N_1515,N_177,N_284);
nor U1516 (N_1516,N_37,N_163);
and U1517 (N_1517,N_554,N_678);
xor U1518 (N_1518,N_51,N_560);
or U1519 (N_1519,N_123,N_149);
or U1520 (N_1520,N_903,N_819);
xor U1521 (N_1521,N_655,N_507);
nor U1522 (N_1522,N_763,N_239);
and U1523 (N_1523,N_317,N_695);
xnor U1524 (N_1524,N_142,N_950);
nor U1525 (N_1525,N_758,N_667);
nand U1526 (N_1526,N_854,N_176);
nand U1527 (N_1527,N_726,N_632);
nor U1528 (N_1528,N_137,N_910);
nand U1529 (N_1529,N_872,N_96);
nand U1530 (N_1530,N_923,N_368);
and U1531 (N_1531,N_404,N_69);
xnor U1532 (N_1532,N_844,N_785);
nor U1533 (N_1533,N_91,N_724);
nand U1534 (N_1534,N_827,N_677);
xor U1535 (N_1535,N_542,N_216);
xor U1536 (N_1536,N_89,N_855);
or U1537 (N_1537,N_923,N_183);
or U1538 (N_1538,N_796,N_130);
nand U1539 (N_1539,N_283,N_408);
xnor U1540 (N_1540,N_944,N_573);
xnor U1541 (N_1541,N_979,N_297);
nand U1542 (N_1542,N_422,N_324);
nor U1543 (N_1543,N_992,N_216);
or U1544 (N_1544,N_95,N_647);
or U1545 (N_1545,N_615,N_835);
or U1546 (N_1546,N_213,N_34);
nand U1547 (N_1547,N_723,N_118);
and U1548 (N_1548,N_645,N_589);
xor U1549 (N_1549,N_25,N_837);
xor U1550 (N_1550,N_669,N_810);
and U1551 (N_1551,N_351,N_413);
nor U1552 (N_1552,N_27,N_713);
and U1553 (N_1553,N_539,N_5);
nand U1554 (N_1554,N_335,N_149);
xor U1555 (N_1555,N_652,N_446);
nor U1556 (N_1556,N_55,N_874);
nand U1557 (N_1557,N_694,N_78);
nor U1558 (N_1558,N_229,N_305);
nor U1559 (N_1559,N_106,N_127);
xnor U1560 (N_1560,N_397,N_262);
or U1561 (N_1561,N_790,N_122);
nand U1562 (N_1562,N_164,N_313);
nor U1563 (N_1563,N_202,N_721);
xor U1564 (N_1564,N_185,N_627);
and U1565 (N_1565,N_176,N_50);
or U1566 (N_1566,N_691,N_54);
or U1567 (N_1567,N_988,N_761);
xnor U1568 (N_1568,N_835,N_418);
nand U1569 (N_1569,N_277,N_414);
or U1570 (N_1570,N_794,N_317);
or U1571 (N_1571,N_117,N_496);
xnor U1572 (N_1572,N_52,N_103);
and U1573 (N_1573,N_667,N_491);
and U1574 (N_1574,N_541,N_206);
and U1575 (N_1575,N_616,N_447);
or U1576 (N_1576,N_557,N_705);
or U1577 (N_1577,N_60,N_369);
nand U1578 (N_1578,N_0,N_767);
nand U1579 (N_1579,N_421,N_829);
nor U1580 (N_1580,N_841,N_600);
nor U1581 (N_1581,N_394,N_653);
nor U1582 (N_1582,N_478,N_333);
or U1583 (N_1583,N_402,N_552);
xnor U1584 (N_1584,N_267,N_348);
or U1585 (N_1585,N_791,N_327);
nor U1586 (N_1586,N_474,N_377);
nand U1587 (N_1587,N_334,N_814);
and U1588 (N_1588,N_258,N_43);
nand U1589 (N_1589,N_852,N_546);
xnor U1590 (N_1590,N_828,N_842);
xnor U1591 (N_1591,N_462,N_122);
xnor U1592 (N_1592,N_734,N_839);
nor U1593 (N_1593,N_683,N_35);
nor U1594 (N_1594,N_484,N_816);
and U1595 (N_1595,N_72,N_916);
or U1596 (N_1596,N_930,N_924);
xor U1597 (N_1597,N_894,N_110);
or U1598 (N_1598,N_831,N_90);
nand U1599 (N_1599,N_230,N_632);
nand U1600 (N_1600,N_933,N_662);
nor U1601 (N_1601,N_399,N_870);
xor U1602 (N_1602,N_258,N_669);
or U1603 (N_1603,N_536,N_660);
and U1604 (N_1604,N_284,N_142);
nand U1605 (N_1605,N_829,N_970);
nor U1606 (N_1606,N_475,N_769);
xnor U1607 (N_1607,N_652,N_842);
nand U1608 (N_1608,N_533,N_838);
and U1609 (N_1609,N_887,N_845);
or U1610 (N_1610,N_90,N_387);
nand U1611 (N_1611,N_146,N_671);
xnor U1612 (N_1612,N_55,N_897);
nor U1613 (N_1613,N_499,N_247);
or U1614 (N_1614,N_650,N_937);
and U1615 (N_1615,N_774,N_139);
nor U1616 (N_1616,N_407,N_594);
nor U1617 (N_1617,N_606,N_893);
xor U1618 (N_1618,N_163,N_197);
or U1619 (N_1619,N_83,N_43);
or U1620 (N_1620,N_638,N_795);
nand U1621 (N_1621,N_895,N_916);
xnor U1622 (N_1622,N_14,N_460);
xnor U1623 (N_1623,N_157,N_934);
and U1624 (N_1624,N_848,N_344);
nand U1625 (N_1625,N_616,N_565);
nor U1626 (N_1626,N_6,N_741);
xnor U1627 (N_1627,N_559,N_856);
xor U1628 (N_1628,N_293,N_723);
xor U1629 (N_1629,N_917,N_233);
nor U1630 (N_1630,N_701,N_892);
or U1631 (N_1631,N_276,N_645);
nor U1632 (N_1632,N_577,N_943);
nand U1633 (N_1633,N_36,N_282);
or U1634 (N_1634,N_57,N_274);
and U1635 (N_1635,N_761,N_744);
or U1636 (N_1636,N_719,N_565);
nor U1637 (N_1637,N_802,N_376);
and U1638 (N_1638,N_290,N_869);
nor U1639 (N_1639,N_618,N_328);
and U1640 (N_1640,N_123,N_761);
and U1641 (N_1641,N_389,N_734);
and U1642 (N_1642,N_92,N_70);
xor U1643 (N_1643,N_787,N_73);
and U1644 (N_1644,N_110,N_70);
or U1645 (N_1645,N_842,N_500);
or U1646 (N_1646,N_801,N_908);
nor U1647 (N_1647,N_868,N_268);
and U1648 (N_1648,N_865,N_964);
and U1649 (N_1649,N_384,N_289);
nor U1650 (N_1650,N_504,N_365);
nand U1651 (N_1651,N_2,N_141);
and U1652 (N_1652,N_115,N_804);
and U1653 (N_1653,N_240,N_34);
xnor U1654 (N_1654,N_66,N_693);
nor U1655 (N_1655,N_222,N_877);
and U1656 (N_1656,N_400,N_214);
or U1657 (N_1657,N_1,N_362);
nor U1658 (N_1658,N_843,N_994);
or U1659 (N_1659,N_784,N_700);
xnor U1660 (N_1660,N_651,N_996);
xor U1661 (N_1661,N_785,N_290);
nor U1662 (N_1662,N_794,N_386);
and U1663 (N_1663,N_449,N_502);
nor U1664 (N_1664,N_641,N_807);
nor U1665 (N_1665,N_951,N_112);
nand U1666 (N_1666,N_860,N_594);
and U1667 (N_1667,N_196,N_549);
nor U1668 (N_1668,N_146,N_218);
nor U1669 (N_1669,N_755,N_948);
nor U1670 (N_1670,N_832,N_310);
and U1671 (N_1671,N_127,N_792);
xnor U1672 (N_1672,N_700,N_860);
and U1673 (N_1673,N_724,N_504);
or U1674 (N_1674,N_808,N_733);
and U1675 (N_1675,N_549,N_620);
or U1676 (N_1676,N_602,N_630);
or U1677 (N_1677,N_914,N_453);
nor U1678 (N_1678,N_574,N_204);
or U1679 (N_1679,N_653,N_210);
nor U1680 (N_1680,N_907,N_105);
or U1681 (N_1681,N_655,N_621);
nor U1682 (N_1682,N_484,N_480);
xor U1683 (N_1683,N_964,N_168);
or U1684 (N_1684,N_195,N_937);
or U1685 (N_1685,N_382,N_467);
xor U1686 (N_1686,N_203,N_37);
nand U1687 (N_1687,N_776,N_910);
xnor U1688 (N_1688,N_17,N_837);
and U1689 (N_1689,N_249,N_345);
nand U1690 (N_1690,N_300,N_76);
or U1691 (N_1691,N_349,N_24);
or U1692 (N_1692,N_379,N_451);
and U1693 (N_1693,N_558,N_424);
nor U1694 (N_1694,N_453,N_966);
and U1695 (N_1695,N_823,N_138);
or U1696 (N_1696,N_126,N_593);
nor U1697 (N_1697,N_376,N_28);
nor U1698 (N_1698,N_938,N_193);
or U1699 (N_1699,N_22,N_430);
xor U1700 (N_1700,N_912,N_971);
and U1701 (N_1701,N_991,N_980);
nor U1702 (N_1702,N_814,N_155);
nand U1703 (N_1703,N_796,N_495);
nand U1704 (N_1704,N_752,N_1);
and U1705 (N_1705,N_998,N_903);
or U1706 (N_1706,N_62,N_402);
and U1707 (N_1707,N_569,N_957);
nand U1708 (N_1708,N_457,N_904);
nor U1709 (N_1709,N_229,N_700);
nand U1710 (N_1710,N_584,N_853);
nor U1711 (N_1711,N_596,N_189);
nor U1712 (N_1712,N_721,N_750);
xnor U1713 (N_1713,N_399,N_37);
nor U1714 (N_1714,N_276,N_849);
and U1715 (N_1715,N_210,N_102);
nor U1716 (N_1716,N_318,N_75);
and U1717 (N_1717,N_862,N_66);
nand U1718 (N_1718,N_429,N_255);
or U1719 (N_1719,N_126,N_870);
xor U1720 (N_1720,N_803,N_862);
xnor U1721 (N_1721,N_950,N_789);
xor U1722 (N_1722,N_262,N_369);
xnor U1723 (N_1723,N_801,N_285);
nor U1724 (N_1724,N_804,N_651);
and U1725 (N_1725,N_375,N_309);
or U1726 (N_1726,N_851,N_960);
or U1727 (N_1727,N_956,N_102);
nand U1728 (N_1728,N_71,N_160);
or U1729 (N_1729,N_82,N_221);
nor U1730 (N_1730,N_850,N_174);
nor U1731 (N_1731,N_764,N_468);
nand U1732 (N_1732,N_983,N_20);
nand U1733 (N_1733,N_335,N_462);
and U1734 (N_1734,N_895,N_127);
nor U1735 (N_1735,N_225,N_595);
nor U1736 (N_1736,N_30,N_385);
and U1737 (N_1737,N_103,N_693);
nand U1738 (N_1738,N_537,N_434);
and U1739 (N_1739,N_422,N_569);
nor U1740 (N_1740,N_925,N_187);
nor U1741 (N_1741,N_149,N_942);
nor U1742 (N_1742,N_968,N_829);
nor U1743 (N_1743,N_614,N_771);
and U1744 (N_1744,N_140,N_658);
nor U1745 (N_1745,N_188,N_615);
nor U1746 (N_1746,N_881,N_727);
and U1747 (N_1747,N_231,N_782);
nor U1748 (N_1748,N_108,N_898);
xor U1749 (N_1749,N_225,N_19);
nand U1750 (N_1750,N_103,N_48);
xor U1751 (N_1751,N_184,N_534);
nor U1752 (N_1752,N_343,N_797);
or U1753 (N_1753,N_632,N_150);
nor U1754 (N_1754,N_937,N_467);
nand U1755 (N_1755,N_294,N_892);
or U1756 (N_1756,N_760,N_219);
nor U1757 (N_1757,N_733,N_309);
nor U1758 (N_1758,N_229,N_596);
and U1759 (N_1759,N_98,N_158);
xor U1760 (N_1760,N_271,N_309);
xor U1761 (N_1761,N_20,N_111);
or U1762 (N_1762,N_160,N_4);
and U1763 (N_1763,N_639,N_540);
xor U1764 (N_1764,N_66,N_81);
nand U1765 (N_1765,N_196,N_348);
or U1766 (N_1766,N_283,N_277);
nor U1767 (N_1767,N_51,N_50);
or U1768 (N_1768,N_37,N_112);
or U1769 (N_1769,N_500,N_16);
xnor U1770 (N_1770,N_757,N_43);
and U1771 (N_1771,N_70,N_351);
and U1772 (N_1772,N_484,N_9);
xor U1773 (N_1773,N_978,N_144);
or U1774 (N_1774,N_866,N_568);
nand U1775 (N_1775,N_131,N_596);
and U1776 (N_1776,N_635,N_933);
or U1777 (N_1777,N_101,N_765);
and U1778 (N_1778,N_526,N_227);
nor U1779 (N_1779,N_274,N_638);
and U1780 (N_1780,N_615,N_134);
nor U1781 (N_1781,N_285,N_563);
and U1782 (N_1782,N_94,N_391);
nor U1783 (N_1783,N_126,N_777);
nor U1784 (N_1784,N_712,N_304);
xnor U1785 (N_1785,N_124,N_18);
xnor U1786 (N_1786,N_505,N_0);
xnor U1787 (N_1787,N_852,N_414);
nor U1788 (N_1788,N_208,N_231);
nand U1789 (N_1789,N_821,N_11);
and U1790 (N_1790,N_313,N_508);
nor U1791 (N_1791,N_204,N_667);
or U1792 (N_1792,N_815,N_912);
nor U1793 (N_1793,N_505,N_112);
and U1794 (N_1794,N_10,N_229);
and U1795 (N_1795,N_151,N_779);
nor U1796 (N_1796,N_592,N_881);
and U1797 (N_1797,N_65,N_739);
xnor U1798 (N_1798,N_880,N_158);
xnor U1799 (N_1799,N_14,N_999);
nand U1800 (N_1800,N_904,N_459);
nor U1801 (N_1801,N_151,N_355);
and U1802 (N_1802,N_734,N_729);
nor U1803 (N_1803,N_388,N_216);
nand U1804 (N_1804,N_440,N_345);
nand U1805 (N_1805,N_179,N_30);
xor U1806 (N_1806,N_362,N_693);
nand U1807 (N_1807,N_527,N_234);
nand U1808 (N_1808,N_445,N_422);
xor U1809 (N_1809,N_447,N_408);
nand U1810 (N_1810,N_888,N_213);
nand U1811 (N_1811,N_43,N_969);
nand U1812 (N_1812,N_723,N_19);
nor U1813 (N_1813,N_297,N_638);
and U1814 (N_1814,N_534,N_560);
and U1815 (N_1815,N_988,N_360);
or U1816 (N_1816,N_133,N_944);
nor U1817 (N_1817,N_288,N_70);
nor U1818 (N_1818,N_605,N_900);
or U1819 (N_1819,N_35,N_327);
or U1820 (N_1820,N_653,N_209);
nor U1821 (N_1821,N_358,N_577);
nand U1822 (N_1822,N_585,N_499);
nor U1823 (N_1823,N_314,N_802);
nor U1824 (N_1824,N_885,N_347);
nor U1825 (N_1825,N_306,N_578);
or U1826 (N_1826,N_316,N_488);
nor U1827 (N_1827,N_87,N_893);
xor U1828 (N_1828,N_788,N_960);
and U1829 (N_1829,N_539,N_120);
nand U1830 (N_1830,N_338,N_55);
or U1831 (N_1831,N_722,N_777);
xnor U1832 (N_1832,N_209,N_458);
nand U1833 (N_1833,N_799,N_86);
nor U1834 (N_1834,N_639,N_619);
and U1835 (N_1835,N_934,N_902);
or U1836 (N_1836,N_450,N_805);
nand U1837 (N_1837,N_743,N_242);
nor U1838 (N_1838,N_440,N_310);
and U1839 (N_1839,N_779,N_331);
nand U1840 (N_1840,N_515,N_140);
and U1841 (N_1841,N_376,N_385);
xnor U1842 (N_1842,N_90,N_229);
xor U1843 (N_1843,N_350,N_238);
or U1844 (N_1844,N_56,N_973);
nor U1845 (N_1845,N_35,N_533);
and U1846 (N_1846,N_561,N_0);
or U1847 (N_1847,N_705,N_710);
nor U1848 (N_1848,N_86,N_628);
nand U1849 (N_1849,N_723,N_663);
nor U1850 (N_1850,N_551,N_789);
and U1851 (N_1851,N_432,N_995);
xor U1852 (N_1852,N_39,N_741);
nand U1853 (N_1853,N_161,N_240);
nor U1854 (N_1854,N_785,N_951);
xor U1855 (N_1855,N_1,N_112);
nand U1856 (N_1856,N_592,N_650);
or U1857 (N_1857,N_848,N_715);
nand U1858 (N_1858,N_508,N_404);
xor U1859 (N_1859,N_548,N_375);
xnor U1860 (N_1860,N_341,N_175);
nand U1861 (N_1861,N_598,N_461);
or U1862 (N_1862,N_374,N_631);
nor U1863 (N_1863,N_631,N_47);
nand U1864 (N_1864,N_571,N_522);
xor U1865 (N_1865,N_673,N_51);
and U1866 (N_1866,N_360,N_295);
xnor U1867 (N_1867,N_169,N_473);
xnor U1868 (N_1868,N_827,N_979);
nand U1869 (N_1869,N_77,N_115);
or U1870 (N_1870,N_136,N_936);
and U1871 (N_1871,N_972,N_612);
nand U1872 (N_1872,N_268,N_531);
nand U1873 (N_1873,N_403,N_807);
xor U1874 (N_1874,N_912,N_200);
xnor U1875 (N_1875,N_126,N_666);
or U1876 (N_1876,N_919,N_168);
xor U1877 (N_1877,N_841,N_437);
or U1878 (N_1878,N_657,N_518);
or U1879 (N_1879,N_76,N_789);
or U1880 (N_1880,N_203,N_842);
and U1881 (N_1881,N_192,N_678);
nor U1882 (N_1882,N_303,N_410);
nor U1883 (N_1883,N_131,N_330);
or U1884 (N_1884,N_173,N_279);
and U1885 (N_1885,N_811,N_568);
and U1886 (N_1886,N_858,N_552);
nand U1887 (N_1887,N_834,N_500);
nor U1888 (N_1888,N_31,N_80);
and U1889 (N_1889,N_637,N_802);
xnor U1890 (N_1890,N_771,N_697);
and U1891 (N_1891,N_133,N_760);
and U1892 (N_1892,N_663,N_356);
nand U1893 (N_1893,N_941,N_205);
and U1894 (N_1894,N_276,N_349);
nand U1895 (N_1895,N_125,N_824);
xor U1896 (N_1896,N_574,N_933);
and U1897 (N_1897,N_43,N_659);
nand U1898 (N_1898,N_103,N_6);
and U1899 (N_1899,N_232,N_424);
xnor U1900 (N_1900,N_289,N_742);
nor U1901 (N_1901,N_151,N_527);
and U1902 (N_1902,N_671,N_916);
or U1903 (N_1903,N_586,N_669);
or U1904 (N_1904,N_93,N_842);
and U1905 (N_1905,N_575,N_125);
nor U1906 (N_1906,N_98,N_567);
xor U1907 (N_1907,N_617,N_607);
nor U1908 (N_1908,N_675,N_342);
xor U1909 (N_1909,N_481,N_466);
xnor U1910 (N_1910,N_856,N_256);
and U1911 (N_1911,N_214,N_743);
xor U1912 (N_1912,N_981,N_586);
and U1913 (N_1913,N_787,N_114);
and U1914 (N_1914,N_118,N_786);
or U1915 (N_1915,N_930,N_702);
and U1916 (N_1916,N_556,N_124);
xor U1917 (N_1917,N_773,N_901);
and U1918 (N_1918,N_163,N_619);
or U1919 (N_1919,N_328,N_425);
nand U1920 (N_1920,N_622,N_691);
or U1921 (N_1921,N_278,N_400);
xnor U1922 (N_1922,N_883,N_1);
nor U1923 (N_1923,N_281,N_944);
and U1924 (N_1924,N_609,N_528);
xor U1925 (N_1925,N_823,N_601);
xnor U1926 (N_1926,N_473,N_704);
or U1927 (N_1927,N_434,N_362);
nand U1928 (N_1928,N_497,N_795);
nand U1929 (N_1929,N_225,N_953);
or U1930 (N_1930,N_894,N_217);
and U1931 (N_1931,N_652,N_264);
or U1932 (N_1932,N_962,N_879);
nor U1933 (N_1933,N_112,N_355);
and U1934 (N_1934,N_867,N_283);
xnor U1935 (N_1935,N_586,N_501);
and U1936 (N_1936,N_346,N_296);
nand U1937 (N_1937,N_725,N_71);
xnor U1938 (N_1938,N_587,N_968);
and U1939 (N_1939,N_743,N_816);
xnor U1940 (N_1940,N_790,N_368);
or U1941 (N_1941,N_803,N_743);
xnor U1942 (N_1942,N_899,N_281);
or U1943 (N_1943,N_851,N_975);
nor U1944 (N_1944,N_884,N_300);
or U1945 (N_1945,N_483,N_315);
nand U1946 (N_1946,N_670,N_709);
nor U1947 (N_1947,N_168,N_904);
or U1948 (N_1948,N_48,N_453);
or U1949 (N_1949,N_823,N_87);
nor U1950 (N_1950,N_686,N_107);
or U1951 (N_1951,N_964,N_284);
nand U1952 (N_1952,N_777,N_545);
nor U1953 (N_1953,N_576,N_827);
nor U1954 (N_1954,N_56,N_438);
nand U1955 (N_1955,N_203,N_543);
nor U1956 (N_1956,N_798,N_145);
or U1957 (N_1957,N_238,N_760);
or U1958 (N_1958,N_187,N_91);
xor U1959 (N_1959,N_512,N_363);
and U1960 (N_1960,N_374,N_596);
nand U1961 (N_1961,N_785,N_471);
and U1962 (N_1962,N_945,N_667);
or U1963 (N_1963,N_401,N_156);
xor U1964 (N_1964,N_171,N_160);
nor U1965 (N_1965,N_924,N_834);
or U1966 (N_1966,N_517,N_62);
nand U1967 (N_1967,N_317,N_244);
xnor U1968 (N_1968,N_126,N_205);
xnor U1969 (N_1969,N_148,N_658);
nand U1970 (N_1970,N_586,N_369);
and U1971 (N_1971,N_286,N_416);
nor U1972 (N_1972,N_528,N_583);
and U1973 (N_1973,N_842,N_420);
or U1974 (N_1974,N_999,N_988);
nand U1975 (N_1975,N_111,N_297);
nor U1976 (N_1976,N_423,N_218);
nor U1977 (N_1977,N_435,N_633);
nor U1978 (N_1978,N_944,N_400);
or U1979 (N_1979,N_655,N_702);
and U1980 (N_1980,N_100,N_474);
nand U1981 (N_1981,N_323,N_437);
xnor U1982 (N_1982,N_484,N_31);
and U1983 (N_1983,N_438,N_295);
xor U1984 (N_1984,N_795,N_968);
nand U1985 (N_1985,N_440,N_807);
nor U1986 (N_1986,N_318,N_565);
nor U1987 (N_1987,N_53,N_864);
nand U1988 (N_1988,N_641,N_407);
xnor U1989 (N_1989,N_98,N_606);
xor U1990 (N_1990,N_355,N_398);
nor U1991 (N_1991,N_294,N_545);
nand U1992 (N_1992,N_418,N_495);
and U1993 (N_1993,N_926,N_552);
and U1994 (N_1994,N_998,N_716);
and U1995 (N_1995,N_382,N_835);
xor U1996 (N_1996,N_228,N_515);
nand U1997 (N_1997,N_16,N_51);
or U1998 (N_1998,N_155,N_265);
nand U1999 (N_1999,N_10,N_47);
xnor U2000 (N_2000,N_1462,N_1688);
nand U2001 (N_2001,N_1063,N_1079);
xnor U2002 (N_2002,N_1767,N_1625);
xnor U2003 (N_2003,N_1894,N_1518);
xor U2004 (N_2004,N_1008,N_1323);
nand U2005 (N_2005,N_1866,N_1977);
or U2006 (N_2006,N_1312,N_1737);
xor U2007 (N_2007,N_1450,N_1247);
and U2008 (N_2008,N_1050,N_1656);
xor U2009 (N_2009,N_1306,N_1914);
or U2010 (N_2010,N_1933,N_1375);
nand U2011 (N_2011,N_1999,N_1469);
nand U2012 (N_2012,N_1748,N_1562);
nand U2013 (N_2013,N_1700,N_1084);
or U2014 (N_2014,N_1495,N_1074);
xnor U2015 (N_2015,N_1037,N_1416);
nor U2016 (N_2016,N_1046,N_1265);
and U2017 (N_2017,N_1476,N_1376);
or U2018 (N_2018,N_1776,N_1344);
nor U2019 (N_2019,N_1163,N_1338);
nor U2020 (N_2020,N_1153,N_1006);
xor U2021 (N_2021,N_1241,N_1036);
xnor U2022 (N_2022,N_1472,N_1165);
nor U2023 (N_2023,N_1712,N_1387);
xnor U2024 (N_2024,N_1188,N_1978);
and U2025 (N_2025,N_1181,N_1134);
nand U2026 (N_2026,N_1938,N_1807);
or U2027 (N_2027,N_1552,N_1996);
xnor U2028 (N_2028,N_1510,N_1377);
xor U2029 (N_2029,N_1325,N_1105);
xor U2030 (N_2030,N_1584,N_1835);
or U2031 (N_2031,N_1498,N_1603);
nor U2032 (N_2032,N_1794,N_1187);
or U2033 (N_2033,N_1088,N_1734);
nand U2034 (N_2034,N_1072,N_1016);
xnor U2035 (N_2035,N_1659,N_1096);
nor U2036 (N_2036,N_1485,N_1963);
xor U2037 (N_2037,N_1280,N_1919);
and U2038 (N_2038,N_1289,N_1981);
and U2039 (N_2039,N_1151,N_1111);
and U2040 (N_2040,N_1802,N_1693);
nand U2041 (N_2041,N_1002,N_1412);
xor U2042 (N_2042,N_1494,N_1646);
or U2043 (N_2043,N_1129,N_1184);
xor U2044 (N_2044,N_1526,N_1537);
nor U2045 (N_2045,N_1653,N_1649);
or U2046 (N_2046,N_1434,N_1106);
nor U2047 (N_2047,N_1077,N_1374);
xor U2048 (N_2048,N_1137,N_1576);
nand U2049 (N_2049,N_1360,N_1669);
xor U2050 (N_2050,N_1628,N_1217);
or U2051 (N_2051,N_1967,N_1921);
xor U2052 (N_2052,N_1451,N_1073);
nand U2053 (N_2053,N_1590,N_1671);
nor U2054 (N_2054,N_1622,N_1349);
or U2055 (N_2055,N_1270,N_1337);
xor U2056 (N_2056,N_1804,N_1068);
nand U2057 (N_2057,N_1224,N_1186);
and U2058 (N_2058,N_1243,N_1432);
xor U2059 (N_2059,N_1435,N_1883);
and U2060 (N_2060,N_1798,N_1230);
and U2061 (N_2061,N_1054,N_1305);
and U2062 (N_2062,N_1538,N_1439);
xor U2063 (N_2063,N_1309,N_1440);
xnor U2064 (N_2064,N_1682,N_1781);
nand U2065 (N_2065,N_1770,N_1635);
and U2066 (N_2066,N_1095,N_1874);
xor U2067 (N_2067,N_1721,N_1658);
nand U2068 (N_2068,N_1122,N_1460);
or U2069 (N_2069,N_1586,N_1501);
nor U2070 (N_2070,N_1930,N_1028);
nand U2071 (N_2071,N_1665,N_1924);
or U2072 (N_2072,N_1246,N_1250);
nand U2073 (N_2073,N_1346,N_1755);
xor U2074 (N_2074,N_1029,N_1558);
xnor U2075 (N_2075,N_1113,N_1823);
nand U2076 (N_2076,N_1262,N_1971);
xor U2077 (N_2077,N_1190,N_1928);
nor U2078 (N_2078,N_1592,N_1131);
xnor U2079 (N_2079,N_1141,N_1834);
nor U2080 (N_2080,N_1993,N_1396);
or U2081 (N_2081,N_1758,N_1557);
nor U2082 (N_2082,N_1244,N_1275);
xor U2083 (N_2083,N_1140,N_1503);
and U2084 (N_2084,N_1463,N_1814);
nor U2085 (N_2085,N_1411,N_1687);
nor U2086 (N_2086,N_1728,N_1358);
nor U2087 (N_2087,N_1808,N_1752);
xor U2088 (N_2088,N_1848,N_1615);
xor U2089 (N_2089,N_1668,N_1855);
xor U2090 (N_2090,N_1547,N_1984);
nor U2091 (N_2091,N_1828,N_1931);
or U2092 (N_2092,N_1395,N_1525);
xor U2093 (N_2093,N_1708,N_1311);
or U2094 (N_2094,N_1689,N_1602);
nor U2095 (N_2095,N_1629,N_1937);
nor U2096 (N_2096,N_1953,N_1322);
xor U2097 (N_2097,N_1870,N_1057);
nor U2098 (N_2098,N_1284,N_1738);
or U2099 (N_2099,N_1569,N_1044);
xor U2100 (N_2100,N_1817,N_1320);
or U2101 (N_2101,N_1004,N_1561);
nor U2102 (N_2102,N_1594,N_1448);
nor U2103 (N_2103,N_1130,N_1259);
nand U2104 (N_2104,N_1923,N_1836);
xnor U2105 (N_2105,N_1315,N_1643);
nand U2106 (N_2106,N_1031,N_1673);
or U2107 (N_2107,N_1410,N_1988);
nand U2108 (N_2108,N_1211,N_1128);
xor U2109 (N_2109,N_1162,N_1422);
nor U2110 (N_2110,N_1944,N_1098);
nor U2111 (N_2111,N_1570,N_1389);
nor U2112 (N_2112,N_1816,N_1559);
nand U2113 (N_2113,N_1261,N_1221);
xnor U2114 (N_2114,N_1583,N_1127);
or U2115 (N_2115,N_1827,N_1905);
and U2116 (N_2116,N_1651,N_1318);
nor U2117 (N_2117,N_1000,N_1156);
nor U2118 (N_2118,N_1465,N_1852);
or U2119 (N_2119,N_1861,N_1763);
nor U2120 (N_2120,N_1433,N_1936);
nand U2121 (N_2121,N_1343,N_1132);
nor U2122 (N_2122,N_1454,N_1645);
nor U2123 (N_2123,N_1279,N_1269);
xnor U2124 (N_2124,N_1862,N_1932);
nand U2125 (N_2125,N_1509,N_1160);
nor U2126 (N_2126,N_1529,N_1906);
nor U2127 (N_2127,N_1125,N_1427);
or U2128 (N_2128,N_1654,N_1869);
or U2129 (N_2129,N_1588,N_1900);
nor U2130 (N_2130,N_1517,N_1466);
nor U2131 (N_2131,N_1918,N_1973);
and U2132 (N_2132,N_1303,N_1108);
xor U2133 (N_2133,N_1058,N_1324);
and U2134 (N_2134,N_1582,N_1185);
and U2135 (N_2135,N_1220,N_1487);
and U2136 (N_2136,N_1255,N_1753);
or U2137 (N_2137,N_1316,N_1694);
xnor U2138 (N_2138,N_1234,N_1880);
nor U2139 (N_2139,N_1512,N_1745);
and U2140 (N_2140,N_1626,N_1200);
and U2141 (N_2141,N_1496,N_1843);
or U2142 (N_2142,N_1601,N_1053);
nand U2143 (N_2143,N_1075,N_1437);
nand U2144 (N_2144,N_1065,N_1169);
nand U2145 (N_2145,N_1032,N_1692);
nand U2146 (N_2146,N_1296,N_1534);
nand U2147 (N_2147,N_1455,N_1380);
xor U2148 (N_2148,N_1196,N_1639);
and U2149 (N_2149,N_1831,N_1676);
xnor U2150 (N_2150,N_1774,N_1846);
or U2151 (N_2151,N_1373,N_1739);
xnor U2152 (N_2152,N_1722,N_1766);
nor U2153 (N_2153,N_1841,N_1959);
or U2154 (N_2154,N_1307,N_1530);
or U2155 (N_2155,N_1295,N_1922);
or U2156 (N_2156,N_1417,N_1082);
nand U2157 (N_2157,N_1340,N_1236);
and U2158 (N_2158,N_1203,N_1334);
nor U2159 (N_2159,N_1438,N_1772);
nand U2160 (N_2160,N_1458,N_1950);
nor U2161 (N_2161,N_1317,N_1744);
xor U2162 (N_2162,N_1453,N_1667);
nor U2163 (N_2163,N_1741,N_1248);
nand U2164 (N_2164,N_1094,N_1818);
nor U2165 (N_2165,N_1867,N_1449);
or U2166 (N_2166,N_1213,N_1347);
xor U2167 (N_2167,N_1452,N_1017);
and U2168 (N_2168,N_1947,N_1729);
nand U2169 (N_2169,N_1565,N_1837);
or U2170 (N_2170,N_1216,N_1903);
xnor U2171 (N_2171,N_1342,N_1256);
and U2172 (N_2172,N_1064,N_1314);
nand U2173 (N_2173,N_1613,N_1982);
nand U2174 (N_2174,N_1087,N_1274);
or U2175 (N_2175,N_1786,N_1524);
nand U2176 (N_2176,N_1574,N_1158);
nand U2177 (N_2177,N_1563,N_1232);
and U2178 (N_2178,N_1797,N_1251);
xnor U2179 (N_2179,N_1522,N_1975);
nand U2180 (N_2180,N_1235,N_1078);
xnor U2181 (N_2181,N_1424,N_1364);
nor U2182 (N_2182,N_1218,N_1523);
nand U2183 (N_2183,N_1090,N_1281);
and U2184 (N_2184,N_1717,N_1935);
nor U2185 (N_2185,N_1104,N_1779);
xor U2186 (N_2186,N_1383,N_1985);
and U2187 (N_2187,N_1150,N_1803);
or U2188 (N_2188,N_1898,N_1372);
nor U2189 (N_2189,N_1761,N_1182);
or U2190 (N_2190,N_1266,N_1969);
nor U2191 (N_2191,N_1366,N_1033);
nor U2192 (N_2192,N_1927,N_1164);
and U2193 (N_2193,N_1564,N_1484);
xnor U2194 (N_2194,N_1851,N_1701);
and U2195 (N_2195,N_1929,N_1157);
or U2196 (N_2196,N_1277,N_1514);
and U2197 (N_2197,N_1515,N_1597);
and U2198 (N_2198,N_1539,N_1145);
xor U2199 (N_2199,N_1173,N_1020);
nor U2200 (N_2200,N_1093,N_1174);
and U2201 (N_2201,N_1249,N_1979);
and U2202 (N_2202,N_1987,N_1013);
or U2203 (N_2203,N_1854,N_1637);
nand U2204 (N_2204,N_1644,N_1608);
nor U2205 (N_2205,N_1567,N_1675);
xor U2206 (N_2206,N_1391,N_1214);
xor U2207 (N_2207,N_1800,N_1974);
xnor U2208 (N_2208,N_1990,N_1202);
or U2209 (N_2209,N_1352,N_1313);
nand U2210 (N_2210,N_1550,N_1414);
or U2211 (N_2211,N_1055,N_1118);
xnor U2212 (N_2212,N_1775,N_1899);
nor U2213 (N_2213,N_1941,N_1394);
and U2214 (N_2214,N_1952,N_1940);
nor U2215 (N_2215,N_1821,N_1718);
xor U2216 (N_2216,N_1301,N_1014);
or U2217 (N_2217,N_1912,N_1756);
nand U2218 (N_2218,N_1039,N_1664);
nor U2219 (N_2219,N_1691,N_1544);
xor U2220 (N_2220,N_1648,N_1192);
nor U2221 (N_2221,N_1273,N_1201);
and U2222 (N_2222,N_1533,N_1117);
or U2223 (N_2223,N_1473,N_1842);
xnor U2224 (N_2224,N_1853,N_1926);
or U2225 (N_2225,N_1067,N_1003);
or U2226 (N_2226,N_1170,N_1168);
nand U2227 (N_2227,N_1092,N_1822);
xor U2228 (N_2228,N_1685,N_1263);
nor U2229 (N_2229,N_1954,N_1212);
nand U2230 (N_2230,N_1580,N_1351);
nor U2231 (N_2231,N_1009,N_1384);
and U2232 (N_2232,N_1609,N_1404);
nand U2233 (N_2233,N_1983,N_1011);
xnor U2234 (N_2234,N_1155,N_1199);
or U2235 (N_2235,N_1893,N_1840);
or U2236 (N_2236,N_1136,N_1459);
or U2237 (N_2237,N_1471,N_1812);
nand U2238 (N_2238,N_1528,N_1773);
xnor U2239 (N_2239,N_1257,N_1829);
or U2240 (N_2240,N_1399,N_1204);
nand U2241 (N_2241,N_1464,N_1686);
and U2242 (N_2242,N_1430,N_1062);
or U2243 (N_2243,N_1124,N_1707);
nor U2244 (N_2244,N_1120,N_1992);
nor U2245 (N_2245,N_1788,N_1896);
or U2246 (N_2246,N_1830,N_1252);
and U2247 (N_2247,N_1536,N_1619);
or U2248 (N_2248,N_1172,N_1879);
nor U2249 (N_2249,N_1227,N_1504);
nand U2250 (N_2250,N_1995,N_1986);
and U2251 (N_2251,N_1194,N_1461);
or U2252 (N_2252,N_1806,N_1732);
nor U2253 (N_2253,N_1060,N_1371);
xnor U2254 (N_2254,N_1666,N_1429);
and U2255 (N_2255,N_1486,N_1787);
or U2256 (N_2256,N_1606,N_1195);
nor U2257 (N_2257,N_1363,N_1333);
and U2258 (N_2258,N_1397,N_1443);
nor U2259 (N_2259,N_1012,N_1030);
nand U2260 (N_2260,N_1285,N_1703);
nor U2261 (N_2261,N_1386,N_1600);
nor U2262 (N_2262,N_1027,N_1239);
and U2263 (N_2263,N_1059,N_1089);
xor U2264 (N_2264,N_1844,N_1589);
nor U2265 (N_2265,N_1310,N_1962);
nor U2266 (N_2266,N_1976,N_1521);
nand U2267 (N_2267,N_1857,N_1081);
xnor U2268 (N_2268,N_1915,N_1139);
or U2269 (N_2269,N_1785,N_1865);
nor U2270 (N_2270,N_1554,N_1260);
nor U2271 (N_2271,N_1208,N_1636);
xor U2272 (N_2272,N_1237,N_1040);
xnor U2273 (N_2273,N_1596,N_1491);
nor U2274 (N_2274,N_1479,N_1610);
nand U2275 (N_2275,N_1112,N_1946);
or U2276 (N_2276,N_1555,N_1513);
nand U2277 (N_2277,N_1365,N_1901);
nand U2278 (N_2278,N_1850,N_1327);
or U2279 (N_2279,N_1282,N_1791);
xor U2280 (N_2280,N_1875,N_1267);
nor U2281 (N_2281,N_1483,N_1955);
nand U2282 (N_2282,N_1210,N_1661);
nor U2283 (N_2283,N_1041,N_1381);
or U2284 (N_2284,N_1864,N_1329);
and U2285 (N_2285,N_1904,N_1276);
nand U2286 (N_2286,N_1577,N_1206);
nand U2287 (N_2287,N_1705,N_1778);
xor U2288 (N_2288,N_1048,N_1727);
xor U2289 (N_2289,N_1253,N_1332);
and U2290 (N_2290,N_1159,N_1436);
and U2291 (N_2291,N_1726,N_1143);
nor U2292 (N_2292,N_1043,N_1710);
and U2293 (N_2293,N_1294,N_1531);
and U2294 (N_2294,N_1431,N_1650);
or U2295 (N_2295,N_1183,N_1575);
xor U2296 (N_2296,N_1810,N_1768);
xnor U2297 (N_2297,N_1350,N_1070);
xnor U2298 (N_2298,N_1716,N_1750);
xnor U2299 (N_2299,N_1418,N_1478);
or U2300 (N_2300,N_1034,N_1403);
nand U2301 (N_2301,N_1910,N_1860);
or U2302 (N_2302,N_1697,N_1747);
nand U2303 (N_2303,N_1402,N_1598);
or U2304 (N_2304,N_1792,N_1925);
nand U2305 (N_2305,N_1878,N_1240);
nand U2306 (N_2306,N_1630,N_1229);
nor U2307 (N_2307,N_1885,N_1998);
or U2308 (N_2308,N_1578,N_1882);
and U2309 (N_2309,N_1527,N_1488);
nor U2310 (N_2310,N_1623,N_1895);
and U2311 (N_2311,N_1254,N_1392);
xor U2312 (N_2312,N_1551,N_1121);
or U2313 (N_2313,N_1892,N_1298);
nor U2314 (N_2314,N_1069,N_1231);
or U2315 (N_2315,N_1475,N_1456);
xnor U2316 (N_2316,N_1083,N_1945);
nor U2317 (N_2317,N_1742,N_1801);
or U2318 (N_2318,N_1611,N_1783);
and U2319 (N_2319,N_1207,N_1226);
nand U2320 (N_2320,N_1382,N_1233);
and U2321 (N_2321,N_1560,N_1714);
nor U2322 (N_2322,N_1856,N_1467);
nor U2323 (N_2323,N_1711,N_1419);
and U2324 (N_2324,N_1368,N_1110);
and U2325 (N_2325,N_1678,N_1457);
xnor U2326 (N_2326,N_1607,N_1908);
and U2327 (N_2327,N_1022,N_1426);
and U2328 (N_2328,N_1790,N_1328);
or U2329 (N_2329,N_1587,N_1287);
and U2330 (N_2330,N_1683,N_1045);
or U2331 (N_2331,N_1133,N_1178);
nor U2332 (N_2332,N_1171,N_1989);
xnor U2333 (N_2333,N_1949,N_1114);
or U2334 (N_2334,N_1091,N_1390);
nand U2335 (N_2335,N_1780,N_1886);
xor U2336 (N_2336,N_1369,N_1388);
and U2337 (N_2337,N_1638,N_1820);
nor U2338 (N_2338,N_1398,N_1147);
nand U2339 (N_2339,N_1595,N_1167);
or U2340 (N_2340,N_1605,N_1519);
nand U2341 (N_2341,N_1876,N_1264);
nand U2342 (N_2342,N_1796,N_1353);
xor U2343 (N_2343,N_1024,N_1751);
xnor U2344 (N_2344,N_1759,N_1757);
and U2345 (N_2345,N_1920,N_1505);
nor U2346 (N_2346,N_1991,N_1228);
nand U2347 (N_2347,N_1180,N_1754);
nor U2348 (N_2348,N_1470,N_1339);
and U2349 (N_2349,N_1839,N_1420);
nand U2350 (N_2350,N_1061,N_1359);
xor U2351 (N_2351,N_1863,N_1507);
nand U2352 (N_2352,N_1321,N_1965);
and U2353 (N_2353,N_1119,N_1939);
nand U2354 (N_2354,N_1502,N_1152);
nand U2355 (N_2355,N_1425,N_1652);
or U2356 (N_2356,N_1546,N_1720);
nor U2357 (N_2357,N_1764,N_1357);
nand U2358 (N_2358,N_1731,N_1593);
xor U2359 (N_2359,N_1604,N_1428);
nor U2360 (N_2360,N_1957,N_1713);
nor U2361 (N_2361,N_1657,N_1345);
or U2362 (N_2362,N_1367,N_1887);
nor U2363 (N_2363,N_1379,N_1406);
nand U2364 (N_2364,N_1482,N_1934);
xnor U2365 (N_2365,N_1699,N_1733);
nor U2366 (N_2366,N_1408,N_1506);
xor U2367 (N_2367,N_1909,N_1581);
or U2368 (N_2368,N_1847,N_1735);
or U2369 (N_2369,N_1535,N_1618);
and U2370 (N_2370,N_1219,N_1477);
or U2371 (N_2371,N_1662,N_1725);
xnor U2372 (N_2372,N_1508,N_1245);
or U2373 (N_2373,N_1001,N_1005);
nand U2374 (N_2374,N_1166,N_1446);
and U2375 (N_2375,N_1288,N_1026);
nand U2376 (N_2376,N_1579,N_1743);
or U2377 (N_2377,N_1585,N_1149);
nand U2378 (N_2378,N_1268,N_1097);
nor U2379 (N_2379,N_1660,N_1746);
or U2380 (N_2380,N_1647,N_1409);
xnor U2381 (N_2381,N_1489,N_1724);
or U2382 (N_2382,N_1719,N_1330);
and U2383 (N_2383,N_1191,N_1354);
and U2384 (N_2384,N_1293,N_1198);
nor U2385 (N_2385,N_1968,N_1964);
nor U2386 (N_2386,N_1709,N_1080);
nand U2387 (N_2387,N_1789,N_1076);
nor U2388 (N_2388,N_1302,N_1286);
xor U2389 (N_2389,N_1407,N_1331);
xnor U2390 (N_2390,N_1749,N_1445);
nor U2391 (N_2391,N_1010,N_1393);
nor U2392 (N_2392,N_1049,N_1300);
and U2393 (N_2393,N_1341,N_1543);
nand U2394 (N_2394,N_1023,N_1497);
or U2395 (N_2395,N_1385,N_1238);
nand U2396 (N_2396,N_1018,N_1291);
and U2397 (N_2397,N_1102,N_1225);
or U2398 (N_2398,N_1571,N_1481);
nand U2399 (N_2399,N_1499,N_1123);
and U2400 (N_2400,N_1056,N_1566);
and U2401 (N_2401,N_1415,N_1336);
nand U2402 (N_2402,N_1771,N_1702);
nor U2403 (N_2403,N_1642,N_1175);
xor U2404 (N_2404,N_1677,N_1304);
nand U2405 (N_2405,N_1889,N_1897);
nor U2406 (N_2406,N_1553,N_1704);
xor U2407 (N_2407,N_1556,N_1468);
nor U2408 (N_2408,N_1292,N_1299);
nand U2409 (N_2409,N_1826,N_1640);
and U2410 (N_2410,N_1308,N_1051);
or U2411 (N_2411,N_1348,N_1681);
xor U2412 (N_2412,N_1634,N_1811);
nor U2413 (N_2413,N_1760,N_1591);
or U2414 (N_2414,N_1258,N_1126);
xor U2415 (N_2415,N_1911,N_1845);
nand U2416 (N_2416,N_1873,N_1819);
xnor U2417 (N_2417,N_1035,N_1142);
xnor U2418 (N_2418,N_1943,N_1961);
or U2419 (N_2419,N_1684,N_1545);
nand U2420 (N_2420,N_1193,N_1997);
or U2421 (N_2421,N_1474,N_1859);
nand U2422 (N_2422,N_1355,N_1135);
xnor U2423 (N_2423,N_1442,N_1616);
xnor U2424 (N_2424,N_1086,N_1071);
and U2425 (N_2425,N_1913,N_1444);
nand U2426 (N_2426,N_1679,N_1493);
nand U2427 (N_2427,N_1614,N_1272);
or U2428 (N_2428,N_1335,N_1107);
and U2429 (N_2429,N_1215,N_1680);
nor U2430 (N_2430,N_1109,N_1103);
and U2431 (N_2431,N_1189,N_1631);
or U2432 (N_2432,N_1769,N_1401);
or U2433 (N_2433,N_1038,N_1695);
nor U2434 (N_2434,N_1633,N_1101);
and U2435 (N_2435,N_1795,N_1884);
nand U2436 (N_2436,N_1907,N_1066);
and U2437 (N_2437,N_1549,N_1632);
or U2438 (N_2438,N_1917,N_1723);
or U2439 (N_2439,N_1490,N_1881);
or U2440 (N_2440,N_1532,N_1670);
or U2441 (N_2441,N_1793,N_1970);
nand U2442 (N_2442,N_1672,N_1858);
nand U2443 (N_2443,N_1520,N_1916);
or U2444 (N_2444,N_1209,N_1283);
xnor U2445 (N_2445,N_1696,N_1568);
nand U2446 (N_2446,N_1378,N_1815);
or U2447 (N_2447,N_1548,N_1019);
xor U2448 (N_2448,N_1805,N_1813);
and U2449 (N_2449,N_1972,N_1278);
nand U2450 (N_2450,N_1176,N_1223);
xor U2451 (N_2451,N_1115,N_1782);
nand U2452 (N_2452,N_1655,N_1047);
and U2453 (N_2453,N_1480,N_1824);
nor U2454 (N_2454,N_1297,N_1868);
or U2455 (N_2455,N_1612,N_1960);
xor U2456 (N_2456,N_1641,N_1849);
or U2457 (N_2457,N_1441,N_1154);
and U2458 (N_2458,N_1447,N_1617);
and U2459 (N_2459,N_1042,N_1500);
xor U2460 (N_2460,N_1116,N_1951);
and U2461 (N_2461,N_1730,N_1948);
nor U2462 (N_2462,N_1980,N_1326);
nand U2463 (N_2463,N_1765,N_1362);
or U2464 (N_2464,N_1715,N_1966);
nand U2465 (N_2465,N_1624,N_1888);
or U2466 (N_2466,N_1511,N_1177);
or U2467 (N_2467,N_1144,N_1516);
nor U2468 (N_2468,N_1838,N_1148);
nor U2469 (N_2469,N_1572,N_1021);
nor U2470 (N_2470,N_1356,N_1161);
nand U2471 (N_2471,N_1319,N_1958);
or U2472 (N_2472,N_1706,N_1099);
or U2473 (N_2473,N_1492,N_1736);
nor U2474 (N_2474,N_1197,N_1085);
nand U2475 (N_2475,N_1690,N_1956);
nor U2476 (N_2476,N_1242,N_1573);
nor U2477 (N_2477,N_1025,N_1799);
nor U2478 (N_2478,N_1370,N_1890);
nand U2479 (N_2479,N_1413,N_1872);
nor U2480 (N_2480,N_1994,N_1100);
nor U2481 (N_2481,N_1015,N_1421);
nor U2482 (N_2482,N_1271,N_1674);
nand U2483 (N_2483,N_1222,N_1762);
nand U2484 (N_2484,N_1902,N_1621);
nand U2485 (N_2485,N_1809,N_1146);
or U2486 (N_2486,N_1777,N_1627);
nor U2487 (N_2487,N_1361,N_1400);
and U2488 (N_2488,N_1825,N_1620);
nand U2489 (N_2489,N_1179,N_1698);
nand U2490 (N_2490,N_1891,N_1290);
nor U2491 (N_2491,N_1405,N_1052);
nor U2492 (N_2492,N_1540,N_1541);
and U2493 (N_2493,N_1871,N_1007);
xor U2494 (N_2494,N_1663,N_1423);
nand U2495 (N_2495,N_1833,N_1942);
xnor U2496 (N_2496,N_1138,N_1542);
or U2497 (N_2497,N_1205,N_1740);
or U2498 (N_2498,N_1832,N_1784);
xor U2499 (N_2499,N_1877,N_1599);
xnor U2500 (N_2500,N_1289,N_1567);
xor U2501 (N_2501,N_1204,N_1120);
nand U2502 (N_2502,N_1390,N_1380);
nand U2503 (N_2503,N_1731,N_1687);
nand U2504 (N_2504,N_1378,N_1248);
nand U2505 (N_2505,N_1327,N_1919);
or U2506 (N_2506,N_1401,N_1301);
and U2507 (N_2507,N_1975,N_1819);
nand U2508 (N_2508,N_1325,N_1553);
or U2509 (N_2509,N_1757,N_1995);
nor U2510 (N_2510,N_1804,N_1536);
or U2511 (N_2511,N_1644,N_1514);
nand U2512 (N_2512,N_1930,N_1106);
or U2513 (N_2513,N_1421,N_1942);
xor U2514 (N_2514,N_1403,N_1476);
or U2515 (N_2515,N_1485,N_1088);
xnor U2516 (N_2516,N_1109,N_1829);
nor U2517 (N_2517,N_1792,N_1243);
and U2518 (N_2518,N_1442,N_1195);
nand U2519 (N_2519,N_1704,N_1676);
or U2520 (N_2520,N_1217,N_1746);
nand U2521 (N_2521,N_1070,N_1493);
nand U2522 (N_2522,N_1440,N_1679);
and U2523 (N_2523,N_1952,N_1097);
and U2524 (N_2524,N_1212,N_1684);
or U2525 (N_2525,N_1730,N_1613);
nand U2526 (N_2526,N_1046,N_1668);
nand U2527 (N_2527,N_1746,N_1960);
or U2528 (N_2528,N_1606,N_1766);
xor U2529 (N_2529,N_1125,N_1354);
and U2530 (N_2530,N_1609,N_1122);
or U2531 (N_2531,N_1725,N_1461);
or U2532 (N_2532,N_1823,N_1424);
nand U2533 (N_2533,N_1382,N_1319);
xor U2534 (N_2534,N_1722,N_1184);
nor U2535 (N_2535,N_1955,N_1030);
nand U2536 (N_2536,N_1444,N_1910);
and U2537 (N_2537,N_1969,N_1987);
or U2538 (N_2538,N_1575,N_1938);
xor U2539 (N_2539,N_1514,N_1950);
nand U2540 (N_2540,N_1760,N_1716);
xnor U2541 (N_2541,N_1349,N_1368);
xor U2542 (N_2542,N_1327,N_1944);
xnor U2543 (N_2543,N_1684,N_1961);
xnor U2544 (N_2544,N_1676,N_1486);
or U2545 (N_2545,N_1748,N_1822);
and U2546 (N_2546,N_1402,N_1605);
xnor U2547 (N_2547,N_1425,N_1403);
nand U2548 (N_2548,N_1309,N_1464);
nand U2549 (N_2549,N_1308,N_1332);
xor U2550 (N_2550,N_1044,N_1355);
nor U2551 (N_2551,N_1243,N_1558);
and U2552 (N_2552,N_1982,N_1499);
nand U2553 (N_2553,N_1218,N_1143);
or U2554 (N_2554,N_1526,N_1125);
xor U2555 (N_2555,N_1225,N_1604);
xor U2556 (N_2556,N_1675,N_1645);
nand U2557 (N_2557,N_1155,N_1545);
nor U2558 (N_2558,N_1320,N_1923);
or U2559 (N_2559,N_1890,N_1018);
xnor U2560 (N_2560,N_1708,N_1852);
xor U2561 (N_2561,N_1310,N_1872);
and U2562 (N_2562,N_1555,N_1666);
or U2563 (N_2563,N_1293,N_1923);
or U2564 (N_2564,N_1692,N_1613);
nor U2565 (N_2565,N_1230,N_1928);
xnor U2566 (N_2566,N_1108,N_1369);
nor U2567 (N_2567,N_1637,N_1513);
and U2568 (N_2568,N_1894,N_1135);
xor U2569 (N_2569,N_1329,N_1226);
and U2570 (N_2570,N_1951,N_1796);
nor U2571 (N_2571,N_1049,N_1892);
and U2572 (N_2572,N_1114,N_1552);
nor U2573 (N_2573,N_1133,N_1240);
xnor U2574 (N_2574,N_1163,N_1505);
nand U2575 (N_2575,N_1641,N_1793);
and U2576 (N_2576,N_1266,N_1036);
nand U2577 (N_2577,N_1899,N_1519);
or U2578 (N_2578,N_1037,N_1682);
and U2579 (N_2579,N_1439,N_1048);
nand U2580 (N_2580,N_1959,N_1444);
nand U2581 (N_2581,N_1516,N_1013);
nor U2582 (N_2582,N_1784,N_1215);
xor U2583 (N_2583,N_1070,N_1634);
nor U2584 (N_2584,N_1560,N_1387);
or U2585 (N_2585,N_1184,N_1638);
nor U2586 (N_2586,N_1134,N_1557);
nor U2587 (N_2587,N_1708,N_1968);
nor U2588 (N_2588,N_1955,N_1548);
nand U2589 (N_2589,N_1306,N_1558);
xor U2590 (N_2590,N_1168,N_1009);
xnor U2591 (N_2591,N_1402,N_1957);
and U2592 (N_2592,N_1627,N_1618);
nand U2593 (N_2593,N_1871,N_1488);
nor U2594 (N_2594,N_1375,N_1776);
and U2595 (N_2595,N_1933,N_1440);
and U2596 (N_2596,N_1247,N_1043);
and U2597 (N_2597,N_1191,N_1385);
or U2598 (N_2598,N_1594,N_1196);
or U2599 (N_2599,N_1231,N_1764);
or U2600 (N_2600,N_1709,N_1241);
xor U2601 (N_2601,N_1765,N_1517);
nor U2602 (N_2602,N_1959,N_1837);
and U2603 (N_2603,N_1191,N_1257);
nor U2604 (N_2604,N_1353,N_1000);
and U2605 (N_2605,N_1852,N_1035);
or U2606 (N_2606,N_1597,N_1334);
nand U2607 (N_2607,N_1019,N_1049);
or U2608 (N_2608,N_1769,N_1093);
nand U2609 (N_2609,N_1624,N_1365);
nor U2610 (N_2610,N_1009,N_1888);
nor U2611 (N_2611,N_1544,N_1248);
xnor U2612 (N_2612,N_1074,N_1586);
xor U2613 (N_2613,N_1443,N_1983);
nand U2614 (N_2614,N_1445,N_1467);
xor U2615 (N_2615,N_1160,N_1451);
nand U2616 (N_2616,N_1521,N_1379);
nand U2617 (N_2617,N_1678,N_1373);
or U2618 (N_2618,N_1108,N_1037);
and U2619 (N_2619,N_1498,N_1185);
or U2620 (N_2620,N_1961,N_1889);
and U2621 (N_2621,N_1337,N_1024);
nand U2622 (N_2622,N_1101,N_1401);
nand U2623 (N_2623,N_1602,N_1057);
nor U2624 (N_2624,N_1992,N_1732);
and U2625 (N_2625,N_1812,N_1154);
nand U2626 (N_2626,N_1210,N_1728);
nand U2627 (N_2627,N_1781,N_1208);
xnor U2628 (N_2628,N_1561,N_1105);
or U2629 (N_2629,N_1662,N_1606);
and U2630 (N_2630,N_1775,N_1477);
nand U2631 (N_2631,N_1873,N_1182);
or U2632 (N_2632,N_1160,N_1792);
and U2633 (N_2633,N_1032,N_1423);
and U2634 (N_2634,N_1123,N_1071);
and U2635 (N_2635,N_1624,N_1491);
xnor U2636 (N_2636,N_1722,N_1411);
nor U2637 (N_2637,N_1914,N_1414);
nand U2638 (N_2638,N_1581,N_1941);
nor U2639 (N_2639,N_1175,N_1756);
and U2640 (N_2640,N_1711,N_1666);
and U2641 (N_2641,N_1676,N_1891);
or U2642 (N_2642,N_1859,N_1984);
nand U2643 (N_2643,N_1014,N_1127);
nand U2644 (N_2644,N_1035,N_1022);
nand U2645 (N_2645,N_1463,N_1380);
and U2646 (N_2646,N_1296,N_1764);
xnor U2647 (N_2647,N_1861,N_1962);
and U2648 (N_2648,N_1142,N_1499);
nand U2649 (N_2649,N_1074,N_1410);
nor U2650 (N_2650,N_1550,N_1036);
xnor U2651 (N_2651,N_1220,N_1319);
nor U2652 (N_2652,N_1790,N_1296);
and U2653 (N_2653,N_1189,N_1986);
nor U2654 (N_2654,N_1674,N_1344);
nor U2655 (N_2655,N_1158,N_1569);
nand U2656 (N_2656,N_1578,N_1372);
and U2657 (N_2657,N_1718,N_1197);
xnor U2658 (N_2658,N_1406,N_1094);
xnor U2659 (N_2659,N_1999,N_1366);
nor U2660 (N_2660,N_1439,N_1237);
and U2661 (N_2661,N_1190,N_1728);
xnor U2662 (N_2662,N_1750,N_1896);
xor U2663 (N_2663,N_1551,N_1414);
or U2664 (N_2664,N_1452,N_1462);
or U2665 (N_2665,N_1502,N_1840);
nor U2666 (N_2666,N_1279,N_1360);
nor U2667 (N_2667,N_1209,N_1884);
nand U2668 (N_2668,N_1710,N_1874);
nor U2669 (N_2669,N_1189,N_1985);
xnor U2670 (N_2670,N_1488,N_1899);
nand U2671 (N_2671,N_1040,N_1457);
nand U2672 (N_2672,N_1095,N_1525);
and U2673 (N_2673,N_1891,N_1305);
and U2674 (N_2674,N_1556,N_1176);
xor U2675 (N_2675,N_1231,N_1025);
nor U2676 (N_2676,N_1112,N_1754);
nor U2677 (N_2677,N_1967,N_1662);
nand U2678 (N_2678,N_1800,N_1664);
or U2679 (N_2679,N_1486,N_1652);
and U2680 (N_2680,N_1014,N_1213);
or U2681 (N_2681,N_1109,N_1295);
nor U2682 (N_2682,N_1598,N_1169);
nor U2683 (N_2683,N_1372,N_1124);
nor U2684 (N_2684,N_1533,N_1665);
xor U2685 (N_2685,N_1671,N_1195);
nor U2686 (N_2686,N_1298,N_1187);
and U2687 (N_2687,N_1573,N_1308);
nor U2688 (N_2688,N_1627,N_1417);
nand U2689 (N_2689,N_1789,N_1925);
nand U2690 (N_2690,N_1783,N_1725);
and U2691 (N_2691,N_1824,N_1724);
nor U2692 (N_2692,N_1876,N_1752);
or U2693 (N_2693,N_1101,N_1543);
nand U2694 (N_2694,N_1332,N_1097);
or U2695 (N_2695,N_1297,N_1053);
nor U2696 (N_2696,N_1582,N_1533);
nand U2697 (N_2697,N_1429,N_1396);
nand U2698 (N_2698,N_1379,N_1650);
and U2699 (N_2699,N_1054,N_1153);
nor U2700 (N_2700,N_1082,N_1174);
or U2701 (N_2701,N_1096,N_1093);
and U2702 (N_2702,N_1365,N_1906);
nand U2703 (N_2703,N_1874,N_1498);
nor U2704 (N_2704,N_1113,N_1418);
and U2705 (N_2705,N_1660,N_1764);
and U2706 (N_2706,N_1362,N_1646);
nor U2707 (N_2707,N_1786,N_1334);
nand U2708 (N_2708,N_1273,N_1591);
nand U2709 (N_2709,N_1501,N_1635);
and U2710 (N_2710,N_1269,N_1076);
xor U2711 (N_2711,N_1890,N_1204);
and U2712 (N_2712,N_1042,N_1279);
nand U2713 (N_2713,N_1185,N_1020);
and U2714 (N_2714,N_1042,N_1275);
xnor U2715 (N_2715,N_1393,N_1760);
or U2716 (N_2716,N_1881,N_1167);
nor U2717 (N_2717,N_1128,N_1281);
or U2718 (N_2718,N_1152,N_1045);
nand U2719 (N_2719,N_1156,N_1180);
and U2720 (N_2720,N_1923,N_1350);
nor U2721 (N_2721,N_1764,N_1285);
and U2722 (N_2722,N_1680,N_1449);
or U2723 (N_2723,N_1415,N_1186);
or U2724 (N_2724,N_1516,N_1125);
nand U2725 (N_2725,N_1143,N_1790);
nor U2726 (N_2726,N_1573,N_1377);
or U2727 (N_2727,N_1528,N_1480);
nor U2728 (N_2728,N_1408,N_1641);
nand U2729 (N_2729,N_1758,N_1247);
nand U2730 (N_2730,N_1221,N_1245);
nor U2731 (N_2731,N_1687,N_1602);
nand U2732 (N_2732,N_1301,N_1361);
xnor U2733 (N_2733,N_1018,N_1838);
and U2734 (N_2734,N_1585,N_1438);
nor U2735 (N_2735,N_1007,N_1317);
or U2736 (N_2736,N_1216,N_1736);
xnor U2737 (N_2737,N_1394,N_1505);
or U2738 (N_2738,N_1829,N_1094);
or U2739 (N_2739,N_1921,N_1797);
and U2740 (N_2740,N_1998,N_1396);
xnor U2741 (N_2741,N_1474,N_1109);
or U2742 (N_2742,N_1322,N_1744);
nand U2743 (N_2743,N_1433,N_1969);
nand U2744 (N_2744,N_1890,N_1048);
xor U2745 (N_2745,N_1816,N_1865);
or U2746 (N_2746,N_1522,N_1711);
and U2747 (N_2747,N_1547,N_1534);
nand U2748 (N_2748,N_1278,N_1900);
nor U2749 (N_2749,N_1151,N_1030);
nand U2750 (N_2750,N_1422,N_1488);
and U2751 (N_2751,N_1716,N_1363);
xor U2752 (N_2752,N_1220,N_1629);
nor U2753 (N_2753,N_1600,N_1062);
or U2754 (N_2754,N_1116,N_1505);
and U2755 (N_2755,N_1003,N_1689);
and U2756 (N_2756,N_1303,N_1059);
nand U2757 (N_2757,N_1078,N_1526);
or U2758 (N_2758,N_1876,N_1590);
nand U2759 (N_2759,N_1214,N_1550);
or U2760 (N_2760,N_1968,N_1149);
nand U2761 (N_2761,N_1031,N_1581);
nand U2762 (N_2762,N_1090,N_1214);
xor U2763 (N_2763,N_1620,N_1031);
nor U2764 (N_2764,N_1234,N_1525);
or U2765 (N_2765,N_1436,N_1764);
and U2766 (N_2766,N_1313,N_1599);
and U2767 (N_2767,N_1172,N_1385);
nor U2768 (N_2768,N_1622,N_1695);
and U2769 (N_2769,N_1947,N_1168);
xor U2770 (N_2770,N_1426,N_1918);
nand U2771 (N_2771,N_1724,N_1117);
nand U2772 (N_2772,N_1685,N_1977);
nand U2773 (N_2773,N_1313,N_1929);
xnor U2774 (N_2774,N_1503,N_1756);
or U2775 (N_2775,N_1167,N_1467);
nand U2776 (N_2776,N_1891,N_1726);
or U2777 (N_2777,N_1175,N_1904);
and U2778 (N_2778,N_1658,N_1118);
and U2779 (N_2779,N_1416,N_1392);
and U2780 (N_2780,N_1346,N_1287);
xor U2781 (N_2781,N_1674,N_1259);
nand U2782 (N_2782,N_1423,N_1234);
and U2783 (N_2783,N_1435,N_1119);
xnor U2784 (N_2784,N_1574,N_1422);
xnor U2785 (N_2785,N_1004,N_1324);
nor U2786 (N_2786,N_1921,N_1070);
or U2787 (N_2787,N_1725,N_1350);
or U2788 (N_2788,N_1741,N_1200);
nand U2789 (N_2789,N_1399,N_1293);
and U2790 (N_2790,N_1069,N_1978);
xnor U2791 (N_2791,N_1631,N_1826);
and U2792 (N_2792,N_1600,N_1861);
xnor U2793 (N_2793,N_1144,N_1293);
and U2794 (N_2794,N_1846,N_1036);
nand U2795 (N_2795,N_1069,N_1452);
nand U2796 (N_2796,N_1420,N_1231);
nand U2797 (N_2797,N_1718,N_1566);
xor U2798 (N_2798,N_1269,N_1396);
or U2799 (N_2799,N_1761,N_1455);
nand U2800 (N_2800,N_1040,N_1563);
xnor U2801 (N_2801,N_1161,N_1024);
nor U2802 (N_2802,N_1413,N_1142);
and U2803 (N_2803,N_1023,N_1813);
or U2804 (N_2804,N_1510,N_1812);
and U2805 (N_2805,N_1955,N_1629);
or U2806 (N_2806,N_1109,N_1645);
and U2807 (N_2807,N_1801,N_1421);
xor U2808 (N_2808,N_1870,N_1042);
nand U2809 (N_2809,N_1854,N_1397);
nor U2810 (N_2810,N_1690,N_1645);
or U2811 (N_2811,N_1784,N_1700);
and U2812 (N_2812,N_1985,N_1482);
or U2813 (N_2813,N_1350,N_1135);
and U2814 (N_2814,N_1660,N_1851);
xnor U2815 (N_2815,N_1611,N_1125);
or U2816 (N_2816,N_1659,N_1147);
xor U2817 (N_2817,N_1122,N_1236);
xnor U2818 (N_2818,N_1780,N_1963);
xor U2819 (N_2819,N_1870,N_1796);
nand U2820 (N_2820,N_1704,N_1090);
or U2821 (N_2821,N_1926,N_1849);
xor U2822 (N_2822,N_1169,N_1607);
or U2823 (N_2823,N_1518,N_1335);
nand U2824 (N_2824,N_1445,N_1028);
xnor U2825 (N_2825,N_1991,N_1002);
and U2826 (N_2826,N_1702,N_1740);
nor U2827 (N_2827,N_1348,N_1663);
and U2828 (N_2828,N_1222,N_1035);
nand U2829 (N_2829,N_1255,N_1418);
and U2830 (N_2830,N_1978,N_1528);
nor U2831 (N_2831,N_1664,N_1732);
xor U2832 (N_2832,N_1871,N_1235);
nor U2833 (N_2833,N_1042,N_1143);
or U2834 (N_2834,N_1222,N_1570);
xnor U2835 (N_2835,N_1880,N_1850);
xor U2836 (N_2836,N_1403,N_1422);
nor U2837 (N_2837,N_1135,N_1848);
nand U2838 (N_2838,N_1020,N_1101);
xor U2839 (N_2839,N_1952,N_1582);
and U2840 (N_2840,N_1037,N_1177);
and U2841 (N_2841,N_1413,N_1839);
nand U2842 (N_2842,N_1973,N_1380);
xor U2843 (N_2843,N_1449,N_1238);
and U2844 (N_2844,N_1800,N_1386);
and U2845 (N_2845,N_1630,N_1826);
and U2846 (N_2846,N_1653,N_1115);
nand U2847 (N_2847,N_1774,N_1970);
and U2848 (N_2848,N_1705,N_1233);
nor U2849 (N_2849,N_1582,N_1825);
nand U2850 (N_2850,N_1341,N_1967);
nor U2851 (N_2851,N_1585,N_1813);
or U2852 (N_2852,N_1955,N_1168);
nor U2853 (N_2853,N_1160,N_1125);
xnor U2854 (N_2854,N_1797,N_1898);
or U2855 (N_2855,N_1077,N_1784);
and U2856 (N_2856,N_1046,N_1405);
xor U2857 (N_2857,N_1854,N_1446);
xor U2858 (N_2858,N_1688,N_1053);
nand U2859 (N_2859,N_1429,N_1090);
nand U2860 (N_2860,N_1966,N_1423);
or U2861 (N_2861,N_1671,N_1293);
xor U2862 (N_2862,N_1298,N_1897);
nand U2863 (N_2863,N_1583,N_1938);
xor U2864 (N_2864,N_1820,N_1982);
and U2865 (N_2865,N_1244,N_1209);
xor U2866 (N_2866,N_1249,N_1000);
xor U2867 (N_2867,N_1670,N_1867);
nand U2868 (N_2868,N_1806,N_1333);
and U2869 (N_2869,N_1415,N_1759);
xnor U2870 (N_2870,N_1405,N_1287);
or U2871 (N_2871,N_1438,N_1147);
nand U2872 (N_2872,N_1084,N_1382);
or U2873 (N_2873,N_1620,N_1048);
xor U2874 (N_2874,N_1508,N_1800);
nor U2875 (N_2875,N_1128,N_1712);
or U2876 (N_2876,N_1781,N_1182);
or U2877 (N_2877,N_1472,N_1423);
nor U2878 (N_2878,N_1680,N_1987);
and U2879 (N_2879,N_1174,N_1407);
nand U2880 (N_2880,N_1124,N_1363);
nand U2881 (N_2881,N_1751,N_1293);
xnor U2882 (N_2882,N_1521,N_1647);
nand U2883 (N_2883,N_1267,N_1415);
nor U2884 (N_2884,N_1674,N_1632);
or U2885 (N_2885,N_1360,N_1512);
xor U2886 (N_2886,N_1778,N_1747);
nand U2887 (N_2887,N_1562,N_1126);
xnor U2888 (N_2888,N_1771,N_1416);
nor U2889 (N_2889,N_1571,N_1342);
xnor U2890 (N_2890,N_1139,N_1767);
nor U2891 (N_2891,N_1702,N_1133);
nand U2892 (N_2892,N_1160,N_1074);
or U2893 (N_2893,N_1338,N_1518);
or U2894 (N_2894,N_1869,N_1675);
xnor U2895 (N_2895,N_1597,N_1478);
xor U2896 (N_2896,N_1164,N_1405);
or U2897 (N_2897,N_1153,N_1188);
and U2898 (N_2898,N_1739,N_1872);
or U2899 (N_2899,N_1271,N_1366);
nand U2900 (N_2900,N_1163,N_1125);
xnor U2901 (N_2901,N_1407,N_1626);
nor U2902 (N_2902,N_1598,N_1567);
nand U2903 (N_2903,N_1805,N_1985);
or U2904 (N_2904,N_1209,N_1932);
or U2905 (N_2905,N_1936,N_1048);
and U2906 (N_2906,N_1873,N_1032);
or U2907 (N_2907,N_1966,N_1864);
nor U2908 (N_2908,N_1136,N_1048);
nor U2909 (N_2909,N_1602,N_1437);
nor U2910 (N_2910,N_1250,N_1295);
and U2911 (N_2911,N_1933,N_1065);
and U2912 (N_2912,N_1030,N_1767);
or U2913 (N_2913,N_1054,N_1187);
or U2914 (N_2914,N_1559,N_1807);
nand U2915 (N_2915,N_1841,N_1675);
or U2916 (N_2916,N_1488,N_1947);
xor U2917 (N_2917,N_1685,N_1548);
and U2918 (N_2918,N_1702,N_1328);
and U2919 (N_2919,N_1277,N_1084);
and U2920 (N_2920,N_1200,N_1199);
nand U2921 (N_2921,N_1525,N_1061);
nor U2922 (N_2922,N_1754,N_1588);
nor U2923 (N_2923,N_1009,N_1570);
or U2924 (N_2924,N_1591,N_1319);
xnor U2925 (N_2925,N_1611,N_1878);
nor U2926 (N_2926,N_1803,N_1238);
xor U2927 (N_2927,N_1755,N_1158);
and U2928 (N_2928,N_1021,N_1585);
nand U2929 (N_2929,N_1094,N_1139);
or U2930 (N_2930,N_1562,N_1519);
and U2931 (N_2931,N_1183,N_1819);
xor U2932 (N_2932,N_1394,N_1693);
xor U2933 (N_2933,N_1783,N_1001);
nor U2934 (N_2934,N_1694,N_1255);
and U2935 (N_2935,N_1447,N_1663);
xnor U2936 (N_2936,N_1268,N_1455);
nor U2937 (N_2937,N_1426,N_1155);
nor U2938 (N_2938,N_1101,N_1951);
or U2939 (N_2939,N_1148,N_1229);
or U2940 (N_2940,N_1134,N_1198);
xor U2941 (N_2941,N_1114,N_1983);
or U2942 (N_2942,N_1917,N_1876);
nand U2943 (N_2943,N_1487,N_1957);
or U2944 (N_2944,N_1950,N_1671);
xor U2945 (N_2945,N_1539,N_1728);
or U2946 (N_2946,N_1041,N_1607);
nand U2947 (N_2947,N_1735,N_1158);
nor U2948 (N_2948,N_1826,N_1038);
nor U2949 (N_2949,N_1748,N_1409);
xor U2950 (N_2950,N_1145,N_1227);
and U2951 (N_2951,N_1838,N_1849);
or U2952 (N_2952,N_1019,N_1145);
or U2953 (N_2953,N_1322,N_1027);
xor U2954 (N_2954,N_1993,N_1733);
or U2955 (N_2955,N_1899,N_1248);
xnor U2956 (N_2956,N_1521,N_1185);
nand U2957 (N_2957,N_1081,N_1752);
nor U2958 (N_2958,N_1539,N_1247);
nor U2959 (N_2959,N_1099,N_1617);
nor U2960 (N_2960,N_1873,N_1911);
xnor U2961 (N_2961,N_1331,N_1229);
nor U2962 (N_2962,N_1766,N_1167);
nand U2963 (N_2963,N_1566,N_1476);
nand U2964 (N_2964,N_1363,N_1691);
or U2965 (N_2965,N_1791,N_1076);
nor U2966 (N_2966,N_1831,N_1308);
nand U2967 (N_2967,N_1032,N_1743);
nor U2968 (N_2968,N_1368,N_1713);
and U2969 (N_2969,N_1006,N_1355);
xnor U2970 (N_2970,N_1373,N_1555);
or U2971 (N_2971,N_1599,N_1292);
xor U2972 (N_2972,N_1623,N_1691);
xor U2973 (N_2973,N_1290,N_1295);
or U2974 (N_2974,N_1062,N_1826);
and U2975 (N_2975,N_1918,N_1649);
nor U2976 (N_2976,N_1983,N_1514);
or U2977 (N_2977,N_1854,N_1322);
nor U2978 (N_2978,N_1449,N_1703);
nor U2979 (N_2979,N_1980,N_1418);
nand U2980 (N_2980,N_1728,N_1604);
nor U2981 (N_2981,N_1823,N_1548);
or U2982 (N_2982,N_1951,N_1679);
or U2983 (N_2983,N_1871,N_1635);
nand U2984 (N_2984,N_1915,N_1549);
or U2985 (N_2985,N_1777,N_1428);
and U2986 (N_2986,N_1889,N_1493);
or U2987 (N_2987,N_1662,N_1197);
or U2988 (N_2988,N_1487,N_1564);
nor U2989 (N_2989,N_1985,N_1006);
nand U2990 (N_2990,N_1191,N_1249);
or U2991 (N_2991,N_1500,N_1060);
xnor U2992 (N_2992,N_1091,N_1340);
or U2993 (N_2993,N_1307,N_1450);
nand U2994 (N_2994,N_1306,N_1569);
nand U2995 (N_2995,N_1803,N_1302);
nor U2996 (N_2996,N_1931,N_1321);
or U2997 (N_2997,N_1184,N_1527);
nor U2998 (N_2998,N_1701,N_1177);
xor U2999 (N_2999,N_1428,N_1880);
xor U3000 (N_3000,N_2971,N_2411);
nor U3001 (N_3001,N_2355,N_2342);
nand U3002 (N_3002,N_2846,N_2534);
nor U3003 (N_3003,N_2024,N_2906);
nand U3004 (N_3004,N_2339,N_2014);
nand U3005 (N_3005,N_2949,N_2495);
nor U3006 (N_3006,N_2220,N_2958);
xnor U3007 (N_3007,N_2379,N_2380);
nand U3008 (N_3008,N_2117,N_2569);
nor U3009 (N_3009,N_2681,N_2023);
nand U3010 (N_3010,N_2377,N_2278);
or U3011 (N_3011,N_2330,N_2086);
nor U3012 (N_3012,N_2243,N_2490);
nand U3013 (N_3013,N_2494,N_2975);
xor U3014 (N_3014,N_2609,N_2318);
and U3015 (N_3015,N_2749,N_2055);
nor U3016 (N_3016,N_2074,N_2298);
and U3017 (N_3017,N_2670,N_2163);
nand U3018 (N_3018,N_2799,N_2302);
nand U3019 (N_3019,N_2648,N_2112);
xnor U3020 (N_3020,N_2818,N_2015);
nand U3021 (N_3021,N_2463,N_2674);
and U3022 (N_3022,N_2970,N_2802);
and U3023 (N_3023,N_2553,N_2990);
or U3024 (N_3024,N_2868,N_2464);
and U3025 (N_3025,N_2890,N_2424);
xnor U3026 (N_3026,N_2416,N_2502);
xor U3027 (N_3027,N_2735,N_2934);
and U3028 (N_3028,N_2107,N_2049);
or U3029 (N_3029,N_2596,N_2779);
xnor U3030 (N_3030,N_2861,N_2831);
or U3031 (N_3031,N_2085,N_2592);
nand U3032 (N_3032,N_2962,N_2509);
or U3033 (N_3033,N_2331,N_2358);
or U3034 (N_3034,N_2886,N_2199);
xnor U3035 (N_3035,N_2558,N_2179);
or U3036 (N_3036,N_2018,N_2451);
and U3037 (N_3037,N_2485,N_2145);
nor U3038 (N_3038,N_2316,N_2727);
xnor U3039 (N_3039,N_2159,N_2973);
nor U3040 (N_3040,N_2707,N_2041);
or U3041 (N_3041,N_2470,N_2610);
or U3042 (N_3042,N_2757,N_2105);
nand U3043 (N_3043,N_2022,N_2539);
xnor U3044 (N_3044,N_2857,N_2255);
nand U3045 (N_3045,N_2754,N_2497);
and U3046 (N_3046,N_2151,N_2414);
and U3047 (N_3047,N_2081,N_2797);
or U3048 (N_3048,N_2459,N_2170);
nand U3049 (N_3049,N_2439,N_2999);
xor U3050 (N_3050,N_2306,N_2564);
xor U3051 (N_3051,N_2598,N_2139);
nand U3052 (N_3052,N_2031,N_2957);
and U3053 (N_3053,N_2078,N_2121);
or U3054 (N_3054,N_2559,N_2567);
and U3055 (N_3055,N_2373,N_2125);
or U3056 (N_3056,N_2263,N_2311);
nor U3057 (N_3057,N_2165,N_2740);
xnor U3058 (N_3058,N_2104,N_2458);
xor U3059 (N_3059,N_2285,N_2352);
xor U3060 (N_3060,N_2479,N_2501);
or U3061 (N_3061,N_2529,N_2475);
nand U3062 (N_3062,N_2771,N_2437);
or U3063 (N_3063,N_2765,N_2972);
nand U3064 (N_3064,N_2190,N_2192);
nor U3065 (N_3065,N_2325,N_2281);
nand U3066 (N_3066,N_2249,N_2708);
nor U3067 (N_3067,N_2624,N_2301);
xor U3068 (N_3068,N_2425,N_2398);
or U3069 (N_3069,N_2233,N_2578);
nor U3070 (N_3070,N_2634,N_2580);
or U3071 (N_3071,N_2524,N_2985);
or U3072 (N_3072,N_2798,N_2323);
nor U3073 (N_3073,N_2863,N_2732);
and U3074 (N_3074,N_2157,N_2713);
and U3075 (N_3075,N_2853,N_2591);
nand U3076 (N_3076,N_2817,N_2291);
xnor U3077 (N_3077,N_2773,N_2090);
nand U3078 (N_3078,N_2204,N_2620);
nor U3079 (N_3079,N_2296,N_2687);
nor U3080 (N_3080,N_2516,N_2884);
xor U3081 (N_3081,N_2313,N_2824);
nor U3082 (N_3082,N_2743,N_2350);
xnor U3083 (N_3083,N_2914,N_2348);
and U3084 (N_3084,N_2625,N_2694);
or U3085 (N_3085,N_2304,N_2636);
or U3086 (N_3086,N_2734,N_2025);
xnor U3087 (N_3087,N_2261,N_2499);
xor U3088 (N_3088,N_2982,N_2527);
xor U3089 (N_3089,N_2211,N_2770);
xnor U3090 (N_3090,N_2554,N_2341);
xnor U3091 (N_3091,N_2433,N_2334);
or U3092 (N_3092,N_2860,N_2653);
and U3093 (N_3093,N_2231,N_2617);
xnor U3094 (N_3094,N_2756,N_2453);
xnor U3095 (N_3095,N_2717,N_2733);
nand U3096 (N_3096,N_2401,N_2573);
or U3097 (N_3097,N_2080,N_2889);
and U3098 (N_3098,N_2202,N_2088);
nand U3099 (N_3099,N_2655,N_2784);
nand U3100 (N_3100,N_2942,N_2966);
xnor U3101 (N_3101,N_2763,N_2308);
or U3102 (N_3102,N_2536,N_2750);
and U3103 (N_3103,N_2830,N_2801);
xnor U3104 (N_3104,N_2438,N_2388);
nand U3105 (N_3105,N_2994,N_2844);
and U3106 (N_3106,N_2483,N_2372);
nor U3107 (N_3107,N_2703,N_2045);
nor U3108 (N_3108,N_2144,N_2752);
and U3109 (N_3109,N_2978,N_2394);
or U3110 (N_3110,N_2445,N_2476);
nand U3111 (N_3111,N_2943,N_2248);
nor U3112 (N_3112,N_2154,N_2540);
or U3113 (N_3113,N_2371,N_2137);
xnor U3114 (N_3114,N_2809,N_2588);
nor U3115 (N_3115,N_2496,N_2858);
nand U3116 (N_3116,N_2893,N_2661);
nand U3117 (N_3117,N_2859,N_2347);
or U3118 (N_3118,N_2155,N_2603);
nor U3119 (N_3119,N_2198,N_2254);
nand U3120 (N_3120,N_2804,N_2851);
nor U3121 (N_3121,N_2354,N_2531);
or U3122 (N_3122,N_2557,N_2396);
nor U3123 (N_3123,N_2050,N_2829);
or U3124 (N_3124,N_2027,N_2276);
and U3125 (N_3125,N_2864,N_2002);
and U3126 (N_3126,N_2506,N_2127);
and U3127 (N_3127,N_2976,N_2923);
or U3128 (N_3128,N_2639,N_2940);
or U3129 (N_3129,N_2761,N_2512);
nor U3130 (N_3130,N_2718,N_2390);
or U3131 (N_3131,N_2106,N_2087);
nor U3132 (N_3132,N_2028,N_2546);
xor U3133 (N_3133,N_2305,N_2378);
or U3134 (N_3134,N_2442,N_2008);
or U3135 (N_3135,N_2288,N_2217);
nor U3136 (N_3136,N_2412,N_2796);
xnor U3137 (N_3137,N_2650,N_2247);
nand U3138 (N_3138,N_2210,N_2030);
xnor U3139 (N_3139,N_2337,N_2629);
or U3140 (N_3140,N_2549,N_2647);
or U3141 (N_3141,N_2753,N_2520);
nand U3142 (N_3142,N_2669,N_2604);
or U3143 (N_3143,N_2937,N_2375);
nand U3144 (N_3144,N_2699,N_2422);
or U3145 (N_3145,N_2156,N_2852);
nor U3146 (N_3146,N_2939,N_2775);
and U3147 (N_3147,N_2491,N_2432);
or U3148 (N_3148,N_2267,N_2901);
xor U3149 (N_3149,N_2979,N_2026);
nor U3150 (N_3150,N_2374,N_2643);
or U3151 (N_3151,N_2742,N_2399);
nor U3152 (N_3152,N_2309,N_2251);
nor U3153 (N_3153,N_2176,N_2505);
and U3154 (N_3154,N_2187,N_2344);
or U3155 (N_3155,N_2357,N_2938);
or U3156 (N_3156,N_2057,N_2072);
and U3157 (N_3157,N_2040,N_2397);
xnor U3158 (N_3158,N_2663,N_2297);
or U3159 (N_3159,N_2126,N_2046);
nor U3160 (N_3160,N_2984,N_2134);
and U3161 (N_3161,N_2128,N_2327);
and U3162 (N_3162,N_2109,N_2964);
nand U3163 (N_3163,N_2205,N_2519);
and U3164 (N_3164,N_2616,N_2630);
nand U3165 (N_3165,N_2033,N_2284);
or U3166 (N_3166,N_2621,N_2315);
nand U3167 (N_3167,N_2482,N_2132);
or U3168 (N_3168,N_2855,N_2880);
or U3169 (N_3169,N_2043,N_2695);
or U3170 (N_3170,N_2436,N_2869);
and U3171 (N_3171,N_2083,N_2688);
nand U3172 (N_3172,N_2518,N_2336);
nor U3173 (N_3173,N_2787,N_2716);
and U3174 (N_3174,N_2686,N_2129);
nor U3175 (N_3175,N_2961,N_2659);
xor U3176 (N_3176,N_2234,N_2840);
nor U3177 (N_3177,N_2140,N_2228);
or U3178 (N_3178,N_2063,N_2907);
nand U3179 (N_3179,N_2444,N_2206);
nand U3180 (N_3180,N_2474,N_2237);
or U3181 (N_3181,N_2701,N_2381);
nor U3182 (N_3182,N_2715,N_2415);
or U3183 (N_3183,N_2769,N_2785);
nor U3184 (N_3184,N_2574,N_2712);
xnor U3185 (N_3185,N_2486,N_2946);
and U3186 (N_3186,N_2200,N_2929);
nand U3187 (N_3187,N_2434,N_2745);
nor U3188 (N_3188,N_2862,N_2113);
xor U3189 (N_3189,N_2329,N_2720);
xnor U3190 (N_3190,N_2645,N_2235);
nor U3191 (N_3191,N_2816,N_2930);
nand U3192 (N_3192,N_2664,N_2792);
nand U3193 (N_3193,N_2768,N_2423);
nor U3194 (N_3194,N_2841,N_2963);
and U3195 (N_3195,N_2766,N_2098);
xnor U3196 (N_3196,N_2577,N_2881);
xor U3197 (N_3197,N_2418,N_2562);
or U3198 (N_3198,N_2409,N_2294);
xnor U3199 (N_3199,N_2166,N_2469);
nor U3200 (N_3200,N_2216,N_2385);
xor U3201 (N_3201,N_2551,N_2811);
nor U3202 (N_3202,N_2995,N_2061);
nand U3203 (N_3203,N_2266,N_2239);
or U3204 (N_3204,N_2471,N_2956);
or U3205 (N_3205,N_2847,N_2678);
nand U3206 (N_3206,N_2488,N_2510);
nor U3207 (N_3207,N_2910,N_2614);
xor U3208 (N_3208,N_2822,N_2833);
or U3209 (N_3209,N_2478,N_2225);
nand U3210 (N_3210,N_2782,N_2158);
nor U3211 (N_3211,N_2544,N_2921);
xnor U3212 (N_3212,N_2959,N_2102);
or U3213 (N_3213,N_2273,N_2089);
and U3214 (N_3214,N_2264,N_2899);
nor U3215 (N_3215,N_2541,N_2843);
or U3216 (N_3216,N_2036,N_2873);
or U3217 (N_3217,N_2138,N_2032);
and U3218 (N_3218,N_2450,N_2421);
and U3219 (N_3219,N_2133,N_2908);
nor U3220 (N_3220,N_2729,N_2219);
or U3221 (N_3221,N_2571,N_2005);
xnor U3222 (N_3222,N_2891,N_2466);
or U3223 (N_3223,N_2324,N_2062);
nor U3224 (N_3224,N_2806,N_2447);
xor U3225 (N_3225,N_2481,N_2292);
or U3226 (N_3226,N_2250,N_2637);
nor U3227 (N_3227,N_2981,N_2983);
xor U3228 (N_3228,N_2682,N_2079);
or U3229 (N_3229,N_2572,N_2218);
nand U3230 (N_3230,N_2825,N_2110);
nand U3231 (N_3231,N_2673,N_2755);
nor U3232 (N_3232,N_2866,N_2555);
and U3233 (N_3233,N_2455,N_2871);
or U3234 (N_3234,N_2666,N_2736);
xnor U3235 (N_3235,N_2888,N_2191);
nor U3236 (N_3236,N_2149,N_2320);
nor U3237 (N_3237,N_2538,N_2928);
or U3238 (N_3238,N_2513,N_2954);
or U3239 (N_3239,N_2523,N_2094);
and U3240 (N_3240,N_2638,N_2279);
or U3241 (N_3241,N_2627,N_2370);
xor U3242 (N_3242,N_2364,N_2277);
nor U3243 (N_3243,N_2082,N_2178);
nand U3244 (N_3244,N_2556,N_2351);
nand U3245 (N_3245,N_2195,N_2586);
nor U3246 (N_3246,N_2826,N_2006);
and U3247 (N_3247,N_2452,N_2004);
xnor U3248 (N_3248,N_2514,N_2147);
xnor U3249 (N_3249,N_2461,N_2582);
or U3250 (N_3250,N_2737,N_2676);
or U3251 (N_3251,N_2417,N_2389);
and U3252 (N_3252,N_2900,N_2644);
nand U3253 (N_3253,N_2593,N_2987);
nand U3254 (N_3254,N_2842,N_2894);
xor U3255 (N_3255,N_2626,N_2980);
nand U3256 (N_3256,N_2500,N_2376);
nand U3257 (N_3257,N_2876,N_2091);
nor U3258 (N_3258,N_2608,N_2212);
xor U3259 (N_3259,N_2515,N_2084);
xor U3260 (N_3260,N_2188,N_2646);
or U3261 (N_3261,N_2693,N_2196);
and U3262 (N_3262,N_2215,N_2283);
nor U3263 (N_3263,N_2790,N_2017);
or U3264 (N_3264,N_2988,N_2677);
xor U3265 (N_3265,N_2714,N_2056);
nand U3266 (N_3266,N_2965,N_2783);
xnor U3267 (N_3267,N_2902,N_2457);
nor U3268 (N_3268,N_2948,N_2454);
or U3269 (N_3269,N_2810,N_2552);
and U3270 (N_3270,N_2835,N_2680);
nand U3271 (N_3271,N_2635,N_2909);
xor U3272 (N_3272,N_2933,N_2696);
or U3273 (N_3273,N_2116,N_2545);
or U3274 (N_3274,N_2882,N_2530);
nor U3275 (N_3275,N_2435,N_2207);
xnor U3276 (N_3276,N_2384,N_2274);
and U3277 (N_3277,N_2649,N_2492);
xor U3278 (N_3278,N_2001,N_2611);
or U3279 (N_3279,N_2366,N_2996);
nor U3280 (N_3280,N_2685,N_2328);
and U3281 (N_3281,N_2181,N_2124);
nor U3282 (N_3282,N_2382,N_2345);
nand U3283 (N_3283,N_2936,N_2989);
xor U3284 (N_3284,N_2143,N_2054);
xor U3285 (N_3285,N_2526,N_2710);
xnor U3286 (N_3286,N_2628,N_2257);
and U3287 (N_3287,N_2780,N_2473);
and U3288 (N_3288,N_2807,N_2537);
nand U3289 (N_3289,N_2808,N_2340);
xnor U3290 (N_3290,N_2183,N_2722);
or U3291 (N_3291,N_2683,N_2259);
and U3292 (N_3292,N_2226,N_2789);
or U3293 (N_3293,N_2542,N_2402);
xor U3294 (N_3294,N_2854,N_2570);
or U3295 (N_3295,N_2991,N_2993);
and U3296 (N_3296,N_2391,N_2877);
xor U3297 (N_3297,N_2613,N_2214);
nor U3298 (N_3298,N_2066,N_2051);
nor U3299 (N_3299,N_2945,N_2821);
and U3300 (N_3300,N_2172,N_2101);
nor U3301 (N_3301,N_2912,N_2668);
nor U3302 (N_3302,N_2037,N_2997);
nand U3303 (N_3303,N_2905,N_2282);
xnor U3304 (N_3304,N_2813,N_2253);
xnor U3305 (N_3305,N_2977,N_2059);
or U3306 (N_3306,N_2387,N_2606);
or U3307 (N_3307,N_2581,N_2299);
and U3308 (N_3308,N_2468,N_2794);
or U3309 (N_3309,N_2349,N_2815);
xor U3310 (N_3310,N_2590,N_2762);
or U3311 (N_3311,N_2405,N_2230);
and U3312 (N_3312,N_2269,N_2672);
nand U3313 (N_3313,N_2723,N_2922);
or U3314 (N_3314,N_2974,N_2547);
nor U3315 (N_3315,N_2532,N_2788);
xnor U3316 (N_3316,N_2561,N_2772);
or U3317 (N_3317,N_2764,N_2926);
or U3318 (N_3318,N_2020,N_2161);
xor U3319 (N_3319,N_2480,N_2245);
and U3320 (N_3320,N_2640,N_2303);
nor U3321 (N_3321,N_2589,N_2068);
nor U3322 (N_3322,N_2310,N_2652);
nor U3323 (N_3323,N_2335,N_2092);
or U3324 (N_3324,N_2189,N_2227);
xnor U3325 (N_3325,N_2575,N_2223);
xnor U3326 (N_3326,N_2193,N_2268);
xor U3327 (N_3327,N_2924,N_2363);
or U3328 (N_3328,N_2786,N_2413);
or U3329 (N_3329,N_2403,N_2021);
or U3330 (N_3330,N_2706,N_2709);
nand U3331 (N_3331,N_2353,N_2420);
or U3332 (N_3332,N_2393,N_2224);
nand U3333 (N_3333,N_2115,N_2201);
xnor U3334 (N_3334,N_2759,N_2725);
and U3335 (N_3335,N_2849,N_2426);
nor U3336 (N_3336,N_2791,N_2684);
or U3337 (N_3337,N_2493,N_2295);
and U3338 (N_3338,N_2605,N_2838);
and U3339 (N_3339,N_2367,N_2150);
xnor U3340 (N_3340,N_2000,N_2952);
nor U3341 (N_3341,N_2618,N_2579);
xnor U3342 (N_3342,N_2034,N_2845);
or U3343 (N_3343,N_2449,N_2969);
nor U3344 (N_3344,N_2103,N_2428);
xor U3345 (N_3345,N_2690,N_2731);
xnor U3346 (N_3346,N_2152,N_2258);
and U3347 (N_3347,N_2044,N_2213);
nand U3348 (N_3348,N_2111,N_2623);
or U3349 (N_3349,N_2697,N_2728);
or U3350 (N_3350,N_2865,N_2365);
and U3351 (N_3351,N_2186,N_2774);
and U3352 (N_3352,N_2916,N_2878);
or U3353 (N_3353,N_2386,N_2691);
xor U3354 (N_3354,N_2071,N_2872);
or U3355 (N_3355,N_2992,N_2820);
or U3356 (N_3356,N_2711,N_2314);
nand U3357 (N_3357,N_2667,N_2917);
nor U3358 (N_3358,N_2289,N_2748);
and U3359 (N_3359,N_2462,N_2065);
and U3360 (N_3360,N_2960,N_2048);
nor U3361 (N_3361,N_2883,N_2898);
xor U3362 (N_3362,N_2038,N_2108);
and U3363 (N_3363,N_2099,N_2064);
nand U3364 (N_3364,N_2767,N_2585);
or U3365 (N_3365,N_2160,N_2662);
and U3366 (N_3366,N_2035,N_2286);
xor U3367 (N_3367,N_2896,N_2793);
nor U3368 (N_3368,N_2427,N_2070);
nor U3369 (N_3369,N_2332,N_2487);
xor U3370 (N_3370,N_2489,N_2174);
and U3371 (N_3371,N_2832,N_2903);
or U3372 (N_3372,N_2548,N_2760);
nor U3373 (N_3373,N_2343,N_2271);
nand U3374 (N_3374,N_2498,N_2758);
or U3375 (N_3375,N_2229,N_2016);
xnor U3376 (N_3376,N_2317,N_2404);
and U3377 (N_3377,N_2369,N_2067);
or U3378 (N_3378,N_2448,N_2615);
xnor U3379 (N_3379,N_2887,N_2795);
xor U3380 (N_3380,N_2550,N_2925);
nor U3381 (N_3381,N_2197,N_2430);
nor U3382 (N_3382,N_2525,N_2290);
nand U3383 (N_3383,N_2915,N_2511);
or U3384 (N_3384,N_2053,N_2232);
or U3385 (N_3385,N_2911,N_2307);
and U3386 (N_3386,N_2719,N_2955);
nand U3387 (N_3387,N_2777,N_2135);
xor U3388 (N_3388,N_2141,N_2660);
and U3389 (N_3389,N_2913,N_2029);
or U3390 (N_3390,N_2221,N_2503);
nor U3391 (N_3391,N_2507,N_2047);
and U3392 (N_3392,N_2167,N_2892);
and U3393 (N_3393,N_2460,N_2563);
nand U3394 (N_3394,N_2408,N_2814);
nand U3395 (N_3395,N_2180,N_2651);
xnor U3396 (N_3396,N_2293,N_2698);
or U3397 (N_3397,N_2114,N_2184);
and U3398 (N_3398,N_2203,N_2828);
xor U3399 (N_3399,N_2967,N_2075);
nand U3400 (N_3400,N_2885,N_2322);
xor U3401 (N_3401,N_2874,N_2153);
nand U3402 (N_3402,N_2587,N_2130);
and U3403 (N_3403,N_2751,N_2776);
and U3404 (N_3404,N_2656,N_2665);
xor U3405 (N_3405,N_2726,N_2778);
and U3406 (N_3406,N_2222,N_2406);
xor U3407 (N_3407,N_2058,N_2240);
nand U3408 (N_3408,N_2472,N_2671);
and U3409 (N_3409,N_2927,N_2599);
xnor U3410 (N_3410,N_2175,N_2897);
nor U3411 (N_3411,N_2265,N_2280);
or U3412 (N_3412,N_2256,N_2704);
nor U3413 (N_3413,N_2244,N_2602);
or U3414 (N_3414,N_2875,N_2168);
nand U3415 (N_3415,N_2819,N_2568);
or U3416 (N_3416,N_2338,N_2935);
or U3417 (N_3417,N_2007,N_2465);
and U3418 (N_3418,N_2441,N_2392);
or U3419 (N_3419,N_2182,N_2528);
xnor U3420 (N_3420,N_2407,N_2837);
and U3421 (N_3421,N_2275,N_2700);
xnor U3422 (N_3422,N_2042,N_2654);
nor U3423 (N_3423,N_2823,N_2724);
nand U3424 (N_3424,N_2738,N_2093);
nand U3425 (N_3425,N_2333,N_2612);
or U3426 (N_3426,N_2346,N_2504);
and U3427 (N_3427,N_2122,N_2642);
nor U3428 (N_3428,N_2576,N_2262);
nor U3429 (N_3429,N_2919,N_2321);
nor U3430 (N_3430,N_2692,N_2312);
xnor U3431 (N_3431,N_2805,N_2879);
xnor U3432 (N_3432,N_2456,N_2246);
or U3433 (N_3433,N_2300,N_2194);
nor U3434 (N_3434,N_2011,N_2870);
xnor U3435 (N_3435,N_2164,N_2270);
nor U3436 (N_3436,N_2931,N_2739);
or U3437 (N_3437,N_2594,N_2359);
xor U3438 (N_3438,N_2566,N_2010);
nor U3439 (N_3439,N_2951,N_2812);
or U3440 (N_3440,N_2400,N_2443);
and U3441 (N_3441,N_2362,N_2076);
nand U3442 (N_3442,N_2131,N_2136);
or U3443 (N_3443,N_2918,N_2583);
and U3444 (N_3444,N_2721,N_2319);
xor U3445 (N_3445,N_2185,N_2368);
xnor U3446 (N_3446,N_2543,N_2508);
and U3447 (N_3447,N_2920,N_2484);
and U3448 (N_3448,N_2326,N_2741);
or U3449 (N_3449,N_2601,N_2119);
or U3450 (N_3450,N_2009,N_2003);
xor U3451 (N_3451,N_2429,N_2019);
xor U3452 (N_3452,N_2622,N_2827);
and U3453 (N_3453,N_2356,N_2631);
nor U3454 (N_3454,N_2834,N_2632);
and U3455 (N_3455,N_2039,N_2272);
nor U3456 (N_3456,N_2410,N_2361);
xor U3457 (N_3457,N_2702,N_2565);
or U3458 (N_3458,N_2947,N_2953);
and U3459 (N_3459,N_2633,N_2856);
nor U3460 (N_3460,N_2904,N_2998);
nor U3461 (N_3461,N_2123,N_2560);
xnor U3462 (N_3462,N_2162,N_2097);
nor U3463 (N_3463,N_2013,N_2395);
nand U3464 (N_3464,N_2100,N_2836);
and U3465 (N_3465,N_2146,N_2619);
or U3466 (N_3466,N_2177,N_2208);
nand U3467 (N_3467,N_2535,N_2142);
nand U3468 (N_3468,N_2069,N_2944);
and U3469 (N_3469,N_2095,N_2744);
nor U3470 (N_3470,N_2584,N_2120);
nor U3471 (N_3471,N_2209,N_2360);
nand U3472 (N_3472,N_2467,N_2171);
and U3473 (N_3473,N_2746,N_2287);
nor U3474 (N_3474,N_2658,N_2431);
xor U3475 (N_3475,N_2657,N_2730);
xnor U3476 (N_3476,N_2839,N_2522);
nand U3477 (N_3477,N_2533,N_2521);
xnor U3478 (N_3478,N_2607,N_2689);
xnor U3479 (N_3479,N_2950,N_2440);
and U3480 (N_3480,N_2242,N_2867);
or U3481 (N_3481,N_2477,N_2595);
nand U3482 (N_3482,N_2941,N_2173);
nand U3483 (N_3483,N_2241,N_2641);
or U3484 (N_3484,N_2012,N_2597);
nand U3485 (N_3485,N_2600,N_2236);
or U3486 (N_3486,N_2800,N_2968);
nand U3487 (N_3487,N_2260,N_2073);
nor U3488 (N_3488,N_2383,N_2169);
xor U3489 (N_3489,N_2148,N_2803);
xor U3490 (N_3490,N_2679,N_2747);
nand U3491 (N_3491,N_2077,N_2675);
xnor U3492 (N_3492,N_2895,N_2850);
xnor U3493 (N_3493,N_2118,N_2446);
or U3494 (N_3494,N_2419,N_2932);
nor U3495 (N_3495,N_2848,N_2052);
and U3496 (N_3496,N_2705,N_2252);
or U3497 (N_3497,N_2238,N_2060);
nor U3498 (N_3498,N_2781,N_2986);
nor U3499 (N_3499,N_2096,N_2517);
nor U3500 (N_3500,N_2937,N_2348);
nand U3501 (N_3501,N_2367,N_2095);
nand U3502 (N_3502,N_2748,N_2983);
xor U3503 (N_3503,N_2170,N_2224);
and U3504 (N_3504,N_2784,N_2857);
and U3505 (N_3505,N_2670,N_2990);
nand U3506 (N_3506,N_2587,N_2976);
and U3507 (N_3507,N_2835,N_2542);
nand U3508 (N_3508,N_2031,N_2766);
nand U3509 (N_3509,N_2063,N_2827);
and U3510 (N_3510,N_2528,N_2447);
nor U3511 (N_3511,N_2665,N_2808);
nor U3512 (N_3512,N_2547,N_2610);
nor U3513 (N_3513,N_2288,N_2079);
and U3514 (N_3514,N_2621,N_2919);
nand U3515 (N_3515,N_2225,N_2013);
xor U3516 (N_3516,N_2710,N_2882);
nand U3517 (N_3517,N_2270,N_2039);
nor U3518 (N_3518,N_2220,N_2016);
or U3519 (N_3519,N_2768,N_2528);
or U3520 (N_3520,N_2087,N_2029);
nor U3521 (N_3521,N_2877,N_2781);
nor U3522 (N_3522,N_2298,N_2471);
or U3523 (N_3523,N_2006,N_2022);
or U3524 (N_3524,N_2375,N_2920);
and U3525 (N_3525,N_2496,N_2642);
nand U3526 (N_3526,N_2943,N_2244);
nor U3527 (N_3527,N_2219,N_2195);
or U3528 (N_3528,N_2855,N_2603);
or U3529 (N_3529,N_2284,N_2547);
nand U3530 (N_3530,N_2829,N_2002);
or U3531 (N_3531,N_2679,N_2011);
and U3532 (N_3532,N_2212,N_2632);
or U3533 (N_3533,N_2000,N_2028);
nor U3534 (N_3534,N_2338,N_2813);
xor U3535 (N_3535,N_2273,N_2542);
xor U3536 (N_3536,N_2139,N_2741);
or U3537 (N_3537,N_2283,N_2217);
nand U3538 (N_3538,N_2316,N_2656);
nor U3539 (N_3539,N_2775,N_2785);
or U3540 (N_3540,N_2124,N_2154);
nor U3541 (N_3541,N_2135,N_2282);
or U3542 (N_3542,N_2724,N_2920);
xnor U3543 (N_3543,N_2624,N_2586);
or U3544 (N_3544,N_2098,N_2361);
or U3545 (N_3545,N_2695,N_2772);
and U3546 (N_3546,N_2616,N_2045);
xnor U3547 (N_3547,N_2898,N_2994);
or U3548 (N_3548,N_2951,N_2677);
or U3549 (N_3549,N_2319,N_2243);
xor U3550 (N_3550,N_2271,N_2996);
xnor U3551 (N_3551,N_2504,N_2722);
and U3552 (N_3552,N_2495,N_2357);
xnor U3553 (N_3553,N_2270,N_2320);
and U3554 (N_3554,N_2778,N_2140);
nor U3555 (N_3555,N_2113,N_2229);
nand U3556 (N_3556,N_2009,N_2175);
and U3557 (N_3557,N_2686,N_2247);
nor U3558 (N_3558,N_2178,N_2441);
and U3559 (N_3559,N_2065,N_2372);
nor U3560 (N_3560,N_2770,N_2674);
and U3561 (N_3561,N_2485,N_2336);
and U3562 (N_3562,N_2033,N_2261);
or U3563 (N_3563,N_2299,N_2997);
nand U3564 (N_3564,N_2410,N_2528);
and U3565 (N_3565,N_2314,N_2036);
or U3566 (N_3566,N_2718,N_2496);
nor U3567 (N_3567,N_2139,N_2989);
nor U3568 (N_3568,N_2273,N_2210);
nor U3569 (N_3569,N_2734,N_2171);
or U3570 (N_3570,N_2819,N_2913);
nor U3571 (N_3571,N_2448,N_2478);
and U3572 (N_3572,N_2908,N_2553);
nor U3573 (N_3573,N_2239,N_2920);
nand U3574 (N_3574,N_2904,N_2664);
or U3575 (N_3575,N_2262,N_2091);
xnor U3576 (N_3576,N_2216,N_2429);
nand U3577 (N_3577,N_2548,N_2338);
nor U3578 (N_3578,N_2663,N_2182);
nor U3579 (N_3579,N_2173,N_2933);
or U3580 (N_3580,N_2462,N_2374);
or U3581 (N_3581,N_2984,N_2243);
or U3582 (N_3582,N_2445,N_2056);
nand U3583 (N_3583,N_2285,N_2781);
or U3584 (N_3584,N_2576,N_2317);
or U3585 (N_3585,N_2921,N_2851);
xnor U3586 (N_3586,N_2949,N_2428);
nor U3587 (N_3587,N_2381,N_2909);
nor U3588 (N_3588,N_2238,N_2827);
nor U3589 (N_3589,N_2456,N_2882);
nand U3590 (N_3590,N_2873,N_2638);
or U3591 (N_3591,N_2996,N_2589);
and U3592 (N_3592,N_2290,N_2150);
and U3593 (N_3593,N_2647,N_2881);
nor U3594 (N_3594,N_2850,N_2298);
nor U3595 (N_3595,N_2217,N_2420);
nand U3596 (N_3596,N_2346,N_2285);
and U3597 (N_3597,N_2581,N_2010);
xor U3598 (N_3598,N_2180,N_2815);
nand U3599 (N_3599,N_2590,N_2910);
xor U3600 (N_3600,N_2918,N_2639);
nand U3601 (N_3601,N_2730,N_2711);
xnor U3602 (N_3602,N_2611,N_2787);
and U3603 (N_3603,N_2662,N_2089);
and U3604 (N_3604,N_2254,N_2887);
nor U3605 (N_3605,N_2753,N_2103);
nor U3606 (N_3606,N_2995,N_2092);
or U3607 (N_3607,N_2329,N_2681);
nor U3608 (N_3608,N_2319,N_2156);
nand U3609 (N_3609,N_2166,N_2111);
nor U3610 (N_3610,N_2134,N_2171);
nor U3611 (N_3611,N_2010,N_2439);
xor U3612 (N_3612,N_2444,N_2666);
xnor U3613 (N_3613,N_2369,N_2723);
and U3614 (N_3614,N_2126,N_2050);
or U3615 (N_3615,N_2700,N_2973);
or U3616 (N_3616,N_2877,N_2303);
nor U3617 (N_3617,N_2406,N_2319);
xor U3618 (N_3618,N_2384,N_2640);
nor U3619 (N_3619,N_2217,N_2582);
and U3620 (N_3620,N_2792,N_2216);
nor U3621 (N_3621,N_2728,N_2502);
and U3622 (N_3622,N_2248,N_2682);
and U3623 (N_3623,N_2182,N_2744);
nand U3624 (N_3624,N_2197,N_2513);
xnor U3625 (N_3625,N_2286,N_2891);
nand U3626 (N_3626,N_2594,N_2181);
xnor U3627 (N_3627,N_2479,N_2507);
and U3628 (N_3628,N_2448,N_2227);
nor U3629 (N_3629,N_2732,N_2871);
nor U3630 (N_3630,N_2830,N_2763);
nor U3631 (N_3631,N_2812,N_2195);
nor U3632 (N_3632,N_2728,N_2923);
nor U3633 (N_3633,N_2901,N_2864);
nor U3634 (N_3634,N_2114,N_2171);
and U3635 (N_3635,N_2924,N_2495);
and U3636 (N_3636,N_2321,N_2974);
nor U3637 (N_3637,N_2435,N_2760);
nand U3638 (N_3638,N_2466,N_2236);
nor U3639 (N_3639,N_2560,N_2889);
and U3640 (N_3640,N_2708,N_2239);
or U3641 (N_3641,N_2534,N_2978);
or U3642 (N_3642,N_2432,N_2718);
nand U3643 (N_3643,N_2528,N_2717);
nand U3644 (N_3644,N_2633,N_2148);
nor U3645 (N_3645,N_2344,N_2426);
and U3646 (N_3646,N_2857,N_2814);
or U3647 (N_3647,N_2369,N_2070);
nor U3648 (N_3648,N_2824,N_2918);
xnor U3649 (N_3649,N_2534,N_2553);
or U3650 (N_3650,N_2891,N_2437);
and U3651 (N_3651,N_2408,N_2913);
or U3652 (N_3652,N_2090,N_2265);
and U3653 (N_3653,N_2168,N_2183);
xnor U3654 (N_3654,N_2591,N_2497);
nor U3655 (N_3655,N_2683,N_2286);
and U3656 (N_3656,N_2051,N_2884);
or U3657 (N_3657,N_2813,N_2043);
or U3658 (N_3658,N_2463,N_2611);
nand U3659 (N_3659,N_2688,N_2855);
nand U3660 (N_3660,N_2907,N_2449);
xnor U3661 (N_3661,N_2932,N_2831);
nor U3662 (N_3662,N_2526,N_2631);
or U3663 (N_3663,N_2281,N_2509);
xnor U3664 (N_3664,N_2474,N_2546);
nand U3665 (N_3665,N_2072,N_2815);
xor U3666 (N_3666,N_2226,N_2396);
xnor U3667 (N_3667,N_2608,N_2233);
xnor U3668 (N_3668,N_2876,N_2315);
nand U3669 (N_3669,N_2662,N_2585);
xnor U3670 (N_3670,N_2505,N_2080);
xnor U3671 (N_3671,N_2876,N_2965);
xnor U3672 (N_3672,N_2736,N_2285);
or U3673 (N_3673,N_2889,N_2056);
xnor U3674 (N_3674,N_2981,N_2421);
or U3675 (N_3675,N_2618,N_2848);
and U3676 (N_3676,N_2810,N_2694);
nor U3677 (N_3677,N_2673,N_2353);
and U3678 (N_3678,N_2671,N_2055);
nand U3679 (N_3679,N_2870,N_2211);
nor U3680 (N_3680,N_2056,N_2766);
and U3681 (N_3681,N_2412,N_2372);
and U3682 (N_3682,N_2027,N_2704);
xor U3683 (N_3683,N_2813,N_2394);
or U3684 (N_3684,N_2829,N_2198);
and U3685 (N_3685,N_2890,N_2899);
nor U3686 (N_3686,N_2242,N_2002);
or U3687 (N_3687,N_2520,N_2882);
xnor U3688 (N_3688,N_2674,N_2121);
and U3689 (N_3689,N_2923,N_2194);
nand U3690 (N_3690,N_2348,N_2651);
xor U3691 (N_3691,N_2289,N_2027);
nor U3692 (N_3692,N_2883,N_2785);
nor U3693 (N_3693,N_2765,N_2637);
and U3694 (N_3694,N_2183,N_2365);
or U3695 (N_3695,N_2245,N_2835);
nand U3696 (N_3696,N_2104,N_2554);
xor U3697 (N_3697,N_2413,N_2064);
and U3698 (N_3698,N_2411,N_2663);
and U3699 (N_3699,N_2285,N_2707);
xnor U3700 (N_3700,N_2253,N_2867);
nor U3701 (N_3701,N_2121,N_2263);
or U3702 (N_3702,N_2255,N_2050);
nand U3703 (N_3703,N_2597,N_2187);
or U3704 (N_3704,N_2934,N_2801);
or U3705 (N_3705,N_2365,N_2713);
nand U3706 (N_3706,N_2989,N_2595);
xor U3707 (N_3707,N_2172,N_2386);
or U3708 (N_3708,N_2711,N_2988);
nand U3709 (N_3709,N_2375,N_2353);
nor U3710 (N_3710,N_2189,N_2088);
xor U3711 (N_3711,N_2342,N_2873);
and U3712 (N_3712,N_2272,N_2849);
or U3713 (N_3713,N_2267,N_2640);
nand U3714 (N_3714,N_2518,N_2501);
and U3715 (N_3715,N_2012,N_2140);
nor U3716 (N_3716,N_2158,N_2375);
nor U3717 (N_3717,N_2392,N_2904);
xnor U3718 (N_3718,N_2366,N_2522);
or U3719 (N_3719,N_2616,N_2572);
or U3720 (N_3720,N_2728,N_2726);
or U3721 (N_3721,N_2702,N_2650);
xor U3722 (N_3722,N_2496,N_2197);
xnor U3723 (N_3723,N_2607,N_2846);
nand U3724 (N_3724,N_2087,N_2536);
or U3725 (N_3725,N_2705,N_2272);
nand U3726 (N_3726,N_2885,N_2562);
xor U3727 (N_3727,N_2483,N_2024);
or U3728 (N_3728,N_2922,N_2674);
or U3729 (N_3729,N_2758,N_2553);
nor U3730 (N_3730,N_2131,N_2583);
or U3731 (N_3731,N_2023,N_2335);
xnor U3732 (N_3732,N_2586,N_2659);
xnor U3733 (N_3733,N_2842,N_2972);
and U3734 (N_3734,N_2858,N_2499);
or U3735 (N_3735,N_2797,N_2263);
nor U3736 (N_3736,N_2767,N_2928);
nand U3737 (N_3737,N_2383,N_2938);
xnor U3738 (N_3738,N_2408,N_2457);
nor U3739 (N_3739,N_2138,N_2327);
xor U3740 (N_3740,N_2462,N_2846);
nand U3741 (N_3741,N_2491,N_2729);
nand U3742 (N_3742,N_2327,N_2941);
nor U3743 (N_3743,N_2164,N_2109);
xor U3744 (N_3744,N_2868,N_2406);
xor U3745 (N_3745,N_2405,N_2709);
or U3746 (N_3746,N_2618,N_2072);
nand U3747 (N_3747,N_2960,N_2968);
nand U3748 (N_3748,N_2794,N_2388);
nand U3749 (N_3749,N_2886,N_2587);
or U3750 (N_3750,N_2503,N_2230);
and U3751 (N_3751,N_2041,N_2921);
nor U3752 (N_3752,N_2144,N_2271);
nand U3753 (N_3753,N_2772,N_2650);
xor U3754 (N_3754,N_2740,N_2510);
and U3755 (N_3755,N_2977,N_2681);
xor U3756 (N_3756,N_2761,N_2355);
nor U3757 (N_3757,N_2390,N_2532);
xor U3758 (N_3758,N_2780,N_2991);
xnor U3759 (N_3759,N_2101,N_2095);
and U3760 (N_3760,N_2130,N_2137);
or U3761 (N_3761,N_2658,N_2297);
and U3762 (N_3762,N_2288,N_2831);
xnor U3763 (N_3763,N_2514,N_2970);
nand U3764 (N_3764,N_2568,N_2183);
or U3765 (N_3765,N_2179,N_2777);
and U3766 (N_3766,N_2747,N_2217);
and U3767 (N_3767,N_2068,N_2858);
xnor U3768 (N_3768,N_2734,N_2359);
nor U3769 (N_3769,N_2293,N_2327);
nand U3770 (N_3770,N_2981,N_2363);
nor U3771 (N_3771,N_2137,N_2306);
and U3772 (N_3772,N_2235,N_2848);
nand U3773 (N_3773,N_2949,N_2066);
nand U3774 (N_3774,N_2289,N_2640);
nand U3775 (N_3775,N_2101,N_2823);
nor U3776 (N_3776,N_2357,N_2536);
nor U3777 (N_3777,N_2472,N_2085);
and U3778 (N_3778,N_2633,N_2624);
nand U3779 (N_3779,N_2323,N_2392);
and U3780 (N_3780,N_2810,N_2295);
and U3781 (N_3781,N_2397,N_2584);
nor U3782 (N_3782,N_2959,N_2810);
or U3783 (N_3783,N_2595,N_2648);
xor U3784 (N_3784,N_2911,N_2611);
nor U3785 (N_3785,N_2442,N_2537);
and U3786 (N_3786,N_2398,N_2973);
and U3787 (N_3787,N_2358,N_2852);
or U3788 (N_3788,N_2711,N_2792);
or U3789 (N_3789,N_2027,N_2106);
or U3790 (N_3790,N_2379,N_2269);
nand U3791 (N_3791,N_2536,N_2958);
and U3792 (N_3792,N_2701,N_2074);
or U3793 (N_3793,N_2338,N_2897);
nor U3794 (N_3794,N_2835,N_2698);
and U3795 (N_3795,N_2164,N_2362);
xnor U3796 (N_3796,N_2208,N_2617);
or U3797 (N_3797,N_2254,N_2668);
or U3798 (N_3798,N_2476,N_2049);
and U3799 (N_3799,N_2940,N_2472);
nand U3800 (N_3800,N_2879,N_2909);
xnor U3801 (N_3801,N_2438,N_2909);
xnor U3802 (N_3802,N_2939,N_2604);
nor U3803 (N_3803,N_2368,N_2132);
or U3804 (N_3804,N_2973,N_2962);
xor U3805 (N_3805,N_2212,N_2439);
nor U3806 (N_3806,N_2547,N_2542);
and U3807 (N_3807,N_2501,N_2847);
nand U3808 (N_3808,N_2659,N_2170);
nor U3809 (N_3809,N_2107,N_2366);
nand U3810 (N_3810,N_2924,N_2006);
and U3811 (N_3811,N_2241,N_2948);
or U3812 (N_3812,N_2323,N_2565);
or U3813 (N_3813,N_2026,N_2298);
nor U3814 (N_3814,N_2640,N_2551);
nor U3815 (N_3815,N_2873,N_2816);
and U3816 (N_3816,N_2325,N_2130);
and U3817 (N_3817,N_2094,N_2231);
nand U3818 (N_3818,N_2170,N_2615);
and U3819 (N_3819,N_2812,N_2540);
nand U3820 (N_3820,N_2888,N_2832);
nand U3821 (N_3821,N_2090,N_2087);
or U3822 (N_3822,N_2283,N_2438);
xor U3823 (N_3823,N_2287,N_2702);
xor U3824 (N_3824,N_2870,N_2660);
or U3825 (N_3825,N_2633,N_2183);
xor U3826 (N_3826,N_2190,N_2977);
or U3827 (N_3827,N_2936,N_2896);
nor U3828 (N_3828,N_2859,N_2939);
nand U3829 (N_3829,N_2621,N_2423);
nor U3830 (N_3830,N_2917,N_2692);
nand U3831 (N_3831,N_2277,N_2662);
or U3832 (N_3832,N_2117,N_2688);
xor U3833 (N_3833,N_2067,N_2114);
nor U3834 (N_3834,N_2067,N_2886);
xnor U3835 (N_3835,N_2277,N_2856);
xor U3836 (N_3836,N_2214,N_2671);
and U3837 (N_3837,N_2385,N_2833);
nor U3838 (N_3838,N_2650,N_2970);
or U3839 (N_3839,N_2401,N_2230);
xor U3840 (N_3840,N_2217,N_2102);
or U3841 (N_3841,N_2676,N_2079);
xor U3842 (N_3842,N_2061,N_2485);
and U3843 (N_3843,N_2423,N_2940);
nand U3844 (N_3844,N_2352,N_2788);
nand U3845 (N_3845,N_2590,N_2239);
xnor U3846 (N_3846,N_2525,N_2137);
nand U3847 (N_3847,N_2563,N_2077);
and U3848 (N_3848,N_2110,N_2280);
and U3849 (N_3849,N_2975,N_2035);
xor U3850 (N_3850,N_2935,N_2716);
xor U3851 (N_3851,N_2176,N_2320);
nor U3852 (N_3852,N_2346,N_2484);
nor U3853 (N_3853,N_2429,N_2381);
nor U3854 (N_3854,N_2301,N_2660);
or U3855 (N_3855,N_2084,N_2955);
nand U3856 (N_3856,N_2736,N_2396);
xor U3857 (N_3857,N_2729,N_2235);
nor U3858 (N_3858,N_2548,N_2136);
nand U3859 (N_3859,N_2756,N_2636);
nor U3860 (N_3860,N_2534,N_2999);
xor U3861 (N_3861,N_2780,N_2103);
and U3862 (N_3862,N_2553,N_2841);
and U3863 (N_3863,N_2438,N_2855);
nand U3864 (N_3864,N_2252,N_2643);
or U3865 (N_3865,N_2311,N_2406);
xnor U3866 (N_3866,N_2816,N_2349);
xnor U3867 (N_3867,N_2996,N_2088);
xnor U3868 (N_3868,N_2827,N_2355);
or U3869 (N_3869,N_2167,N_2651);
or U3870 (N_3870,N_2163,N_2516);
nor U3871 (N_3871,N_2284,N_2278);
xnor U3872 (N_3872,N_2923,N_2515);
nor U3873 (N_3873,N_2025,N_2973);
and U3874 (N_3874,N_2244,N_2349);
and U3875 (N_3875,N_2462,N_2714);
nand U3876 (N_3876,N_2248,N_2713);
nand U3877 (N_3877,N_2638,N_2843);
nand U3878 (N_3878,N_2330,N_2853);
xor U3879 (N_3879,N_2642,N_2506);
or U3880 (N_3880,N_2458,N_2423);
or U3881 (N_3881,N_2365,N_2740);
and U3882 (N_3882,N_2790,N_2504);
or U3883 (N_3883,N_2637,N_2908);
and U3884 (N_3884,N_2007,N_2533);
xor U3885 (N_3885,N_2330,N_2627);
nor U3886 (N_3886,N_2035,N_2350);
xor U3887 (N_3887,N_2524,N_2978);
nand U3888 (N_3888,N_2774,N_2428);
xor U3889 (N_3889,N_2264,N_2488);
xor U3890 (N_3890,N_2844,N_2513);
nor U3891 (N_3891,N_2800,N_2577);
and U3892 (N_3892,N_2011,N_2368);
xnor U3893 (N_3893,N_2125,N_2301);
and U3894 (N_3894,N_2488,N_2687);
and U3895 (N_3895,N_2678,N_2959);
nor U3896 (N_3896,N_2577,N_2814);
and U3897 (N_3897,N_2506,N_2295);
and U3898 (N_3898,N_2338,N_2788);
and U3899 (N_3899,N_2262,N_2310);
nor U3900 (N_3900,N_2631,N_2942);
and U3901 (N_3901,N_2336,N_2767);
nor U3902 (N_3902,N_2682,N_2214);
and U3903 (N_3903,N_2066,N_2068);
nand U3904 (N_3904,N_2757,N_2223);
and U3905 (N_3905,N_2034,N_2736);
nor U3906 (N_3906,N_2395,N_2759);
nor U3907 (N_3907,N_2092,N_2113);
nand U3908 (N_3908,N_2362,N_2651);
nand U3909 (N_3909,N_2088,N_2091);
or U3910 (N_3910,N_2182,N_2406);
and U3911 (N_3911,N_2250,N_2720);
nor U3912 (N_3912,N_2093,N_2814);
nand U3913 (N_3913,N_2362,N_2436);
and U3914 (N_3914,N_2615,N_2197);
and U3915 (N_3915,N_2606,N_2281);
and U3916 (N_3916,N_2071,N_2647);
nor U3917 (N_3917,N_2429,N_2040);
xor U3918 (N_3918,N_2975,N_2159);
and U3919 (N_3919,N_2512,N_2982);
and U3920 (N_3920,N_2242,N_2518);
nand U3921 (N_3921,N_2787,N_2342);
and U3922 (N_3922,N_2720,N_2240);
nand U3923 (N_3923,N_2961,N_2643);
nor U3924 (N_3924,N_2207,N_2445);
xor U3925 (N_3925,N_2073,N_2862);
nand U3926 (N_3926,N_2043,N_2032);
nand U3927 (N_3927,N_2266,N_2805);
nand U3928 (N_3928,N_2517,N_2886);
xnor U3929 (N_3929,N_2827,N_2993);
xnor U3930 (N_3930,N_2587,N_2599);
nor U3931 (N_3931,N_2967,N_2641);
xor U3932 (N_3932,N_2575,N_2284);
xnor U3933 (N_3933,N_2983,N_2474);
or U3934 (N_3934,N_2673,N_2299);
nor U3935 (N_3935,N_2366,N_2788);
and U3936 (N_3936,N_2562,N_2545);
nand U3937 (N_3937,N_2175,N_2017);
xor U3938 (N_3938,N_2464,N_2646);
nand U3939 (N_3939,N_2330,N_2106);
nand U3940 (N_3940,N_2026,N_2311);
nor U3941 (N_3941,N_2861,N_2834);
and U3942 (N_3942,N_2106,N_2564);
nor U3943 (N_3943,N_2830,N_2678);
and U3944 (N_3944,N_2518,N_2905);
xnor U3945 (N_3945,N_2465,N_2050);
or U3946 (N_3946,N_2372,N_2020);
nor U3947 (N_3947,N_2939,N_2221);
nor U3948 (N_3948,N_2774,N_2448);
xor U3949 (N_3949,N_2434,N_2490);
or U3950 (N_3950,N_2175,N_2117);
nor U3951 (N_3951,N_2269,N_2257);
or U3952 (N_3952,N_2618,N_2958);
or U3953 (N_3953,N_2183,N_2615);
nor U3954 (N_3954,N_2542,N_2272);
nor U3955 (N_3955,N_2557,N_2354);
nand U3956 (N_3956,N_2512,N_2511);
and U3957 (N_3957,N_2776,N_2880);
nor U3958 (N_3958,N_2051,N_2226);
and U3959 (N_3959,N_2809,N_2805);
or U3960 (N_3960,N_2420,N_2404);
and U3961 (N_3961,N_2262,N_2332);
and U3962 (N_3962,N_2670,N_2697);
xor U3963 (N_3963,N_2860,N_2182);
nor U3964 (N_3964,N_2072,N_2194);
or U3965 (N_3965,N_2370,N_2207);
or U3966 (N_3966,N_2296,N_2851);
or U3967 (N_3967,N_2806,N_2495);
nor U3968 (N_3968,N_2835,N_2832);
or U3969 (N_3969,N_2598,N_2581);
nor U3970 (N_3970,N_2110,N_2421);
nor U3971 (N_3971,N_2935,N_2738);
nor U3972 (N_3972,N_2865,N_2740);
xnor U3973 (N_3973,N_2815,N_2296);
and U3974 (N_3974,N_2934,N_2027);
and U3975 (N_3975,N_2819,N_2095);
nor U3976 (N_3976,N_2896,N_2908);
nor U3977 (N_3977,N_2286,N_2136);
and U3978 (N_3978,N_2470,N_2526);
or U3979 (N_3979,N_2916,N_2149);
and U3980 (N_3980,N_2835,N_2028);
or U3981 (N_3981,N_2460,N_2695);
xnor U3982 (N_3982,N_2713,N_2196);
and U3983 (N_3983,N_2275,N_2385);
or U3984 (N_3984,N_2175,N_2821);
nor U3985 (N_3985,N_2345,N_2117);
nor U3986 (N_3986,N_2459,N_2959);
nor U3987 (N_3987,N_2380,N_2935);
nand U3988 (N_3988,N_2285,N_2714);
or U3989 (N_3989,N_2863,N_2534);
xnor U3990 (N_3990,N_2899,N_2056);
nor U3991 (N_3991,N_2944,N_2122);
xnor U3992 (N_3992,N_2026,N_2868);
nor U3993 (N_3993,N_2902,N_2894);
nor U3994 (N_3994,N_2744,N_2501);
nand U3995 (N_3995,N_2977,N_2406);
xnor U3996 (N_3996,N_2758,N_2920);
xor U3997 (N_3997,N_2348,N_2081);
nor U3998 (N_3998,N_2562,N_2079);
nand U3999 (N_3999,N_2736,N_2876);
xnor U4000 (N_4000,N_3665,N_3386);
and U4001 (N_4001,N_3790,N_3146);
nand U4002 (N_4002,N_3644,N_3658);
and U4003 (N_4003,N_3361,N_3450);
or U4004 (N_4004,N_3445,N_3093);
xor U4005 (N_4005,N_3606,N_3229);
nand U4006 (N_4006,N_3461,N_3322);
xor U4007 (N_4007,N_3143,N_3602);
nor U4008 (N_4008,N_3342,N_3954);
or U4009 (N_4009,N_3025,N_3028);
and U4010 (N_4010,N_3203,N_3264);
nand U4011 (N_4011,N_3403,N_3556);
xnor U4012 (N_4012,N_3687,N_3940);
or U4013 (N_4013,N_3615,N_3559);
and U4014 (N_4014,N_3395,N_3111);
and U4015 (N_4015,N_3250,N_3627);
nor U4016 (N_4016,N_3917,N_3145);
xor U4017 (N_4017,N_3127,N_3996);
or U4018 (N_4018,N_3511,N_3712);
nor U4019 (N_4019,N_3955,N_3531);
and U4020 (N_4020,N_3694,N_3743);
and U4021 (N_4021,N_3612,N_3034);
or U4022 (N_4022,N_3488,N_3423);
nor U4023 (N_4023,N_3826,N_3865);
or U4024 (N_4024,N_3630,N_3920);
nor U4025 (N_4025,N_3036,N_3016);
or U4026 (N_4026,N_3001,N_3387);
xnor U4027 (N_4027,N_3498,N_3147);
xor U4028 (N_4028,N_3592,N_3645);
nor U4029 (N_4029,N_3239,N_3906);
nor U4030 (N_4030,N_3839,N_3655);
and U4031 (N_4031,N_3761,N_3447);
or U4032 (N_4032,N_3689,N_3880);
nor U4033 (N_4033,N_3795,N_3750);
or U4034 (N_4034,N_3589,N_3767);
xor U4035 (N_4035,N_3527,N_3174);
nand U4036 (N_4036,N_3378,N_3452);
nor U4037 (N_4037,N_3838,N_3537);
nand U4038 (N_4038,N_3860,N_3693);
xor U4039 (N_4039,N_3169,N_3078);
and U4040 (N_4040,N_3084,N_3613);
nand U4041 (N_4041,N_3079,N_3968);
or U4042 (N_4042,N_3925,N_3811);
nand U4043 (N_4043,N_3916,N_3432);
nor U4044 (N_4044,N_3905,N_3185);
and U4045 (N_4045,N_3998,N_3473);
and U4046 (N_4046,N_3924,N_3439);
nor U4047 (N_4047,N_3942,N_3479);
nand U4048 (N_4048,N_3560,N_3696);
or U4049 (N_4049,N_3047,N_3142);
nor U4050 (N_4050,N_3327,N_3719);
nor U4051 (N_4051,N_3421,N_3818);
nor U4052 (N_4052,N_3113,N_3292);
or U4053 (N_4053,N_3757,N_3549);
nand U4054 (N_4054,N_3262,N_3911);
or U4055 (N_4055,N_3938,N_3813);
and U4056 (N_4056,N_3502,N_3797);
nor U4057 (N_4057,N_3291,N_3434);
nor U4058 (N_4058,N_3414,N_3004);
nor U4059 (N_4059,N_3850,N_3263);
or U4060 (N_4060,N_3637,N_3579);
nor U4061 (N_4061,N_3981,N_3893);
and U4062 (N_4062,N_3503,N_3440);
xor U4063 (N_4063,N_3669,N_3897);
or U4064 (N_4064,N_3334,N_3260);
nand U4065 (N_4065,N_3995,N_3833);
and U4066 (N_4066,N_3989,N_3999);
xor U4067 (N_4067,N_3726,N_3844);
and U4068 (N_4068,N_3883,N_3272);
or U4069 (N_4069,N_3377,N_3934);
nor U4070 (N_4070,N_3889,N_3189);
nor U4071 (N_4071,N_3184,N_3245);
xor U4072 (N_4072,N_3639,N_3216);
or U4073 (N_4073,N_3072,N_3837);
nor U4074 (N_4074,N_3582,N_3345);
nor U4075 (N_4075,N_3504,N_3476);
xor U4076 (N_4076,N_3636,N_3659);
and U4077 (N_4077,N_3483,N_3446);
nand U4078 (N_4078,N_3993,N_3879);
and U4079 (N_4079,N_3755,N_3153);
or U4080 (N_4080,N_3284,N_3633);
and U4081 (N_4081,N_3720,N_3992);
xnor U4082 (N_4082,N_3187,N_3324);
nor U4083 (N_4083,N_3904,N_3902);
nand U4084 (N_4084,N_3033,N_3714);
nand U4085 (N_4085,N_3020,N_3822);
and U4086 (N_4086,N_3759,N_3279);
and U4087 (N_4087,N_3647,N_3769);
or U4088 (N_4088,N_3443,N_3708);
nand U4089 (N_4089,N_3638,N_3182);
nand U4090 (N_4090,N_3186,N_3149);
xor U4091 (N_4091,N_3383,N_3364);
nand U4092 (N_4092,N_3406,N_3908);
or U4093 (N_4093,N_3789,N_3032);
and U4094 (N_4094,N_3832,N_3922);
xnor U4095 (N_4095,N_3201,N_3872);
xnor U4096 (N_4096,N_3990,N_3703);
nand U4097 (N_4097,N_3371,N_3175);
or U4098 (N_4098,N_3429,N_3598);
and U4099 (N_4099,N_3510,N_3027);
nand U4100 (N_4100,N_3303,N_3963);
nor U4101 (N_4101,N_3831,N_3006);
xor U4102 (N_4102,N_3375,N_3901);
nor U4103 (N_4103,N_3877,N_3608);
or U4104 (N_4104,N_3958,N_3609);
nor U4105 (N_4105,N_3578,N_3233);
and U4106 (N_4106,N_3862,N_3148);
nand U4107 (N_4107,N_3629,N_3318);
or U4108 (N_4108,N_3914,N_3382);
or U4109 (N_4109,N_3497,N_3056);
nand U4110 (N_4110,N_3868,N_3120);
xnor U4111 (N_4111,N_3799,N_3086);
or U4112 (N_4112,N_3514,N_3794);
and U4113 (N_4113,N_3209,N_3248);
or U4114 (N_4114,N_3548,N_3017);
or U4115 (N_4115,N_3063,N_3251);
xnor U4116 (N_4116,N_3221,N_3157);
nor U4117 (N_4117,N_3223,N_3426);
nor U4118 (N_4118,N_3709,N_3884);
xnor U4119 (N_4119,N_3624,N_3170);
xnor U4120 (N_4120,N_3165,N_3772);
nand U4121 (N_4121,N_3115,N_3746);
nor U4122 (N_4122,N_3987,N_3700);
xor U4123 (N_4123,N_3254,N_3411);
nand U4124 (N_4124,N_3929,N_3517);
nand U4125 (N_4125,N_3043,N_3711);
or U4126 (N_4126,N_3273,N_3338);
or U4127 (N_4127,N_3129,N_3011);
and U4128 (N_4128,N_3569,N_3845);
xor U4129 (N_4129,N_3379,N_3601);
nor U4130 (N_4130,N_3183,N_3604);
and U4131 (N_4131,N_3941,N_3727);
xnor U4132 (N_4132,N_3951,N_3672);
and U4133 (N_4133,N_3200,N_3753);
and U4134 (N_4134,N_3828,N_3128);
nor U4135 (N_4135,N_3112,N_3923);
xnor U4136 (N_4136,N_3090,N_3685);
and U4137 (N_4137,N_3670,N_3529);
and U4138 (N_4138,N_3437,N_3695);
or U4139 (N_4139,N_3651,N_3910);
or U4140 (N_4140,N_3023,N_3523);
or U4141 (N_4141,N_3349,N_3222);
nor U4142 (N_4142,N_3830,N_3438);
and U4143 (N_4143,N_3247,N_3009);
nand U4144 (N_4144,N_3863,N_3045);
nor U4145 (N_4145,N_3119,N_3053);
nand U4146 (N_4146,N_3050,N_3232);
and U4147 (N_4147,N_3026,N_3648);
xnor U4148 (N_4148,N_3352,N_3874);
or U4149 (N_4149,N_3277,N_3835);
and U4150 (N_4150,N_3758,N_3158);
xnor U4151 (N_4151,N_3354,N_3249);
nor U4152 (N_4152,N_3041,N_3402);
or U4153 (N_4153,N_3763,N_3915);
or U4154 (N_4154,N_3857,N_3280);
nand U4155 (N_4155,N_3163,N_3328);
nand U4156 (N_4156,N_3661,N_3809);
xnor U4157 (N_4157,N_3805,N_3926);
and U4158 (N_4158,N_3180,N_3649);
and U4159 (N_4159,N_3384,N_3887);
and U4160 (N_4160,N_3590,N_3092);
or U4161 (N_4161,N_3405,N_3135);
nand U4162 (N_4162,N_3208,N_3226);
xor U4163 (N_4163,N_3722,N_3238);
xor U4164 (N_4164,N_3583,N_3428);
or U4165 (N_4165,N_3817,N_3586);
and U4166 (N_4166,N_3932,N_3370);
or U4167 (N_4167,N_3984,N_3039);
nor U4168 (N_4168,N_3521,N_3492);
and U4169 (N_4169,N_3010,N_3316);
and U4170 (N_4170,N_3786,N_3357);
or U4171 (N_4171,N_3820,N_3882);
or U4172 (N_4172,N_3089,N_3509);
nand U4173 (N_4173,N_3783,N_3243);
nor U4174 (N_4174,N_3030,N_3935);
and U4175 (N_4175,N_3625,N_3051);
and U4176 (N_4176,N_3731,N_3296);
xnor U4177 (N_4177,N_3031,N_3409);
nand U4178 (N_4178,N_3391,N_3530);
xor U4179 (N_4179,N_3807,N_3875);
xor U4180 (N_4180,N_3946,N_3317);
and U4181 (N_4181,N_3562,N_3132);
xnor U4182 (N_4182,N_3038,N_3528);
nand U4183 (N_4183,N_3224,N_3468);
xnor U4184 (N_4184,N_3507,N_3372);
nor U4185 (N_4185,N_3436,N_3080);
or U4186 (N_4186,N_3048,N_3332);
and U4187 (N_4187,N_3713,N_3765);
or U4188 (N_4188,N_3853,N_3100);
nand U4189 (N_4189,N_3650,N_3538);
or U4190 (N_4190,N_3454,N_3939);
and U4191 (N_4191,N_3131,N_3526);
and U4192 (N_4192,N_3614,N_3546);
nand U4193 (N_4193,N_3305,N_3351);
nand U4194 (N_4194,N_3657,N_3267);
and U4195 (N_4195,N_3485,N_3660);
nand U4196 (N_4196,N_3441,N_3344);
nor U4197 (N_4197,N_3408,N_3197);
nand U4198 (N_4198,N_3557,N_3744);
or U4199 (N_4199,N_3253,N_3044);
or U4200 (N_4200,N_3899,N_3094);
xor U4201 (N_4201,N_3737,N_3340);
and U4202 (N_4202,N_3416,N_3854);
nor U4203 (N_4203,N_3653,N_3717);
xor U4204 (N_4204,N_3302,N_3130);
nor U4205 (N_4205,N_3482,N_3793);
or U4206 (N_4206,N_3550,N_3431);
nand U4207 (N_4207,N_3323,N_3255);
xnor U4208 (N_4208,N_3121,N_3977);
nand U4209 (N_4209,N_3295,N_3155);
or U4210 (N_4210,N_3469,N_3234);
or U4211 (N_4211,N_3894,N_3419);
or U4212 (N_4212,N_3774,N_3240);
and U4213 (N_4213,N_3707,N_3268);
nor U4214 (N_4214,N_3430,N_3088);
and U4215 (N_4215,N_3558,N_3154);
or U4216 (N_4216,N_3739,N_3396);
or U4217 (N_4217,N_3801,N_3500);
or U4218 (N_4218,N_3635,N_3796);
and U4219 (N_4219,N_3029,N_3551);
nand U4220 (N_4220,N_3545,N_3355);
xnor U4221 (N_4221,N_3335,N_3964);
nor U4222 (N_4222,N_3547,N_3435);
xor U4223 (N_4223,N_3478,N_3885);
and U4224 (N_4224,N_3505,N_3288);
nor U4225 (N_4225,N_3881,N_3193);
xor U4226 (N_4226,N_3631,N_3046);
nor U4227 (N_4227,N_3164,N_3433);
nand U4228 (N_4228,N_3580,N_3847);
xor U4229 (N_4229,N_3674,N_3646);
and U4230 (N_4230,N_3936,N_3139);
nor U4231 (N_4231,N_3070,N_3297);
nand U4232 (N_4232,N_3969,N_3591);
xnor U4233 (N_4233,N_3385,N_3871);
xor U4234 (N_4234,N_3227,N_3108);
or U4235 (N_4235,N_3962,N_3365);
or U4236 (N_4236,N_3289,N_3779);
or U4237 (N_4237,N_3778,N_3971);
and U4238 (N_4238,N_3771,N_3073);
xnor U4239 (N_4239,N_3827,N_3716);
nand U4240 (N_4240,N_3159,N_3643);
and U4241 (N_4241,N_3194,N_3252);
nand U4242 (N_4242,N_3195,N_3301);
nor U4243 (N_4243,N_3667,N_3725);
nand U4244 (N_4244,N_3376,N_3561);
xor U4245 (N_4245,N_3161,N_3898);
nand U4246 (N_4246,N_3840,N_3055);
nor U4247 (N_4247,N_3230,N_3098);
and U4248 (N_4248,N_3508,N_3074);
nor U4249 (N_4249,N_3976,N_3015);
nand U4250 (N_4250,N_3870,N_3621);
nand U4251 (N_4251,N_3961,N_3587);
or U4252 (N_4252,N_3160,N_3710);
nor U4253 (N_4253,N_3134,N_3988);
nor U4254 (N_4254,N_3366,N_3652);
nor U4255 (N_4255,N_3718,N_3415);
or U4256 (N_4256,N_3861,N_3616);
nand U4257 (N_4257,N_3196,N_3945);
nor U4258 (N_4258,N_3705,N_3480);
or U4259 (N_4259,N_3347,N_3455);
nand U4260 (N_4260,N_3290,N_3400);
nand U4261 (N_4261,N_3040,N_3848);
nand U4262 (N_4262,N_3486,N_3188);
or U4263 (N_4263,N_3890,N_3677);
xnor U4264 (N_4264,N_3593,N_3067);
nor U4265 (N_4265,N_3325,N_3623);
or U4266 (N_4266,N_3867,N_3059);
nand U4267 (N_4267,N_3540,N_3640);
nor U4268 (N_4268,N_3620,N_3506);
or U4269 (N_4269,N_3581,N_3052);
xnor U4270 (N_4270,N_3764,N_3214);
and U4271 (N_4271,N_3599,N_3541);
nand U4272 (N_4272,N_3049,N_3515);
xor U4273 (N_4273,N_3575,N_3851);
or U4274 (N_4274,N_3019,N_3125);
or U4275 (N_4275,N_3949,N_3204);
nand U4276 (N_4276,N_3064,N_3424);
and U4277 (N_4277,N_3470,N_3662);
or U4278 (N_4278,N_3472,N_3215);
nor U4279 (N_4279,N_3738,N_3320);
nand U4280 (N_4280,N_3261,N_3337);
and U4281 (N_4281,N_3525,N_3002);
nand U4282 (N_4282,N_3389,N_3166);
nand U4283 (N_4283,N_3109,N_3679);
and U4284 (N_4284,N_3736,N_3596);
and U4285 (N_4285,N_3684,N_3594);
and U4286 (N_4286,N_3333,N_3780);
xor U4287 (N_4287,N_3265,N_3212);
nor U4288 (N_4288,N_3381,N_3293);
and U4289 (N_4289,N_3819,N_3133);
or U4290 (N_4290,N_3585,N_3570);
and U4291 (N_4291,N_3751,N_3481);
nand U4292 (N_4292,N_3691,N_3516);
nand U4293 (N_4293,N_3566,N_3256);
and U4294 (N_4294,N_3495,N_3618);
nand U4295 (N_4295,N_3000,N_3137);
nand U4296 (N_4296,N_3276,N_3314);
nor U4297 (N_4297,N_3363,N_3773);
xor U4298 (N_4298,N_3274,N_3307);
nor U4299 (N_4299,N_3855,N_3057);
xor U4300 (N_4300,N_3610,N_3420);
nor U4301 (N_4301,N_3617,N_3448);
and U4302 (N_4302,N_3501,N_3022);
and U4303 (N_4303,N_3791,N_3096);
or U4304 (N_4304,N_3299,N_3933);
nor U4305 (N_4305,N_3206,N_3690);
or U4306 (N_4306,N_3800,N_3810);
or U4307 (N_4307,N_3770,N_3061);
nor U4308 (N_4308,N_3721,N_3417);
xnor U4309 (N_4309,N_3362,N_3663);
xor U4310 (N_4310,N_3422,N_3785);
nand U4311 (N_4311,N_3900,N_3066);
nor U4312 (N_4312,N_3784,N_3595);
nor U4313 (N_4313,N_3058,N_3979);
nand U4314 (N_4314,N_3983,N_3496);
nand U4315 (N_4315,N_3802,N_3336);
nor U4316 (N_4316,N_3171,N_3572);
or U4317 (N_4317,N_3519,N_3427);
nand U4318 (N_4318,N_3686,N_3777);
nand U4319 (N_4319,N_3565,N_3699);
and U4320 (N_4320,N_3823,N_3449);
xor U4321 (N_4321,N_3117,N_3442);
xor U4322 (N_4322,N_3680,N_3309);
nor U4323 (N_4323,N_3458,N_3173);
or U4324 (N_4324,N_3007,N_3972);
nand U4325 (N_4325,N_3841,N_3359);
nor U4326 (N_4326,N_3313,N_3634);
or U4327 (N_4327,N_3607,N_3346);
nor U4328 (N_4328,N_3950,N_3866);
and U4329 (N_4329,N_3281,N_3353);
or U4330 (N_4330,N_3903,N_3285);
xnor U4331 (N_4331,N_3178,N_3733);
and U4332 (N_4332,N_3756,N_3308);
xor U4333 (N_4333,N_3298,N_3054);
xor U4334 (N_4334,N_3682,N_3003);
xor U4335 (N_4335,N_3919,N_3666);
or U4336 (N_4336,N_3846,N_3518);
xnor U4337 (N_4337,N_3312,N_3418);
nor U4338 (N_4338,N_3788,N_3343);
or U4339 (N_4339,N_3013,N_3852);
nand U4340 (N_4340,N_3076,N_3842);
xnor U4341 (N_4341,N_3487,N_3220);
and U4342 (N_4342,N_3018,N_3266);
nor U4343 (N_4343,N_3723,N_3489);
nor U4344 (N_4344,N_3729,N_3404);
nor U4345 (N_4345,N_3329,N_3804);
and U4346 (N_4346,N_3453,N_3918);
xnor U4347 (N_4347,N_3735,N_3388);
or U4348 (N_4348,N_3715,N_3167);
nand U4349 (N_4349,N_3005,N_3896);
xnor U4350 (N_4350,N_3179,N_3543);
nand U4351 (N_4351,N_3787,N_3091);
and U4352 (N_4352,N_3688,N_3869);
xor U4353 (N_4353,N_3948,N_3747);
and U4354 (N_4354,N_3350,N_3563);
or U4355 (N_4355,N_3241,N_3457);
nor U4356 (N_4356,N_3300,N_3218);
and U4357 (N_4357,N_3451,N_3975);
xnor U4358 (N_4358,N_3464,N_3683);
nand U4359 (N_4359,N_3460,N_3664);
xnor U4360 (N_4360,N_3597,N_3225);
nand U4361 (N_4361,N_3973,N_3812);
nand U4362 (N_4362,N_3124,N_3858);
nand U4363 (N_4363,N_3808,N_3270);
xnor U4364 (N_4364,N_3083,N_3490);
nor U4365 (N_4365,N_3339,N_3412);
and U4366 (N_4366,N_3980,N_3675);
or U4367 (N_4367,N_3278,N_3380);
and U4368 (N_4368,N_3271,N_3294);
and U4369 (N_4369,N_3319,N_3927);
xor U4370 (N_4370,N_3207,N_3876);
xor U4371 (N_4371,N_3524,N_3536);
nor U4372 (N_4372,N_3282,N_3012);
and U4373 (N_4373,N_3834,N_3413);
nor U4374 (N_4374,N_3087,N_3697);
and U4375 (N_4375,N_3985,N_3475);
or U4376 (N_4376,N_3678,N_3287);
nor U4377 (N_4377,N_3836,N_3605);
or U4378 (N_4378,N_3762,N_3692);
or U4379 (N_4379,N_3749,N_3199);
xnor U4380 (N_4380,N_3283,N_3732);
nor U4381 (N_4381,N_3728,N_3367);
nand U4382 (N_4382,N_3564,N_3060);
nand U4383 (N_4383,N_3150,N_3702);
or U4384 (N_4384,N_3062,N_3573);
or U4385 (N_4385,N_3105,N_3168);
nand U4386 (N_4386,N_3205,N_3097);
and U4387 (N_4387,N_3895,N_3210);
or U4388 (N_4388,N_3921,N_3095);
nor U4389 (N_4389,N_3390,N_3065);
nor U4390 (N_4390,N_3535,N_3101);
xor U4391 (N_4391,N_3859,N_3397);
nor U4392 (N_4392,N_3956,N_3782);
xnor U4393 (N_4393,N_3520,N_3965);
nor U4394 (N_4394,N_3035,N_3913);
or U4395 (N_4395,N_3068,N_3947);
and U4396 (N_4396,N_3600,N_3997);
nor U4397 (N_4397,N_3474,N_3330);
or U4398 (N_4398,N_3304,N_3588);
and U4399 (N_4399,N_3162,N_3192);
nand U4400 (N_4400,N_3202,N_3775);
or U4401 (N_4401,N_3829,N_3522);
nor U4402 (N_4402,N_3953,N_3966);
nand U4403 (N_4403,N_3994,N_3584);
nor U4404 (N_4404,N_3781,N_3116);
nand U4405 (N_4405,N_3217,N_3491);
nor U4406 (N_4406,N_3331,N_3310);
and U4407 (N_4407,N_3512,N_3748);
and U4408 (N_4408,N_3081,N_3499);
nor U4409 (N_4409,N_3231,N_3311);
or U4410 (N_4410,N_3141,N_3532);
and U4411 (N_4411,N_3176,N_3741);
xor U4412 (N_4412,N_3816,N_3075);
and U4413 (N_4413,N_3156,N_3172);
and U4414 (N_4414,N_3698,N_3246);
nand U4415 (N_4415,N_3856,N_3654);
or U4416 (N_4416,N_3392,N_3024);
nor U4417 (N_4417,N_3542,N_3668);
and U4418 (N_4418,N_3467,N_3766);
xor U4419 (N_4419,N_3211,N_3102);
nor U4420 (N_4420,N_3704,N_3213);
nor U4421 (N_4421,N_3825,N_3394);
nor U4422 (N_4422,N_3959,N_3103);
nand U4423 (N_4423,N_3671,N_3373);
nor U4424 (N_4424,N_3410,N_3348);
or U4425 (N_4425,N_3768,N_3021);
and U4426 (N_4426,N_3803,N_3471);
nor U4427 (N_4427,N_3140,N_3114);
nand U4428 (N_4428,N_3107,N_3151);
nand U4429 (N_4429,N_3356,N_3177);
xnor U4430 (N_4430,N_3909,N_3465);
and U4431 (N_4431,N_3622,N_3891);
xnor U4432 (N_4432,N_3701,N_3071);
nand U4433 (N_4433,N_3513,N_3244);
or U4434 (N_4434,N_3398,N_3306);
and U4435 (N_4435,N_3628,N_3407);
nand U4436 (N_4436,N_3888,N_3912);
xor U4437 (N_4437,N_3494,N_3360);
and U4438 (N_4438,N_3126,N_3967);
nand U4439 (N_4439,N_3673,N_3752);
nor U4440 (N_4440,N_3190,N_3554);
xnor U4441 (N_4441,N_3477,N_3123);
xor U4442 (N_4442,N_3907,N_3534);
nor U4443 (N_4443,N_3886,N_3326);
nor U4444 (N_4444,N_3957,N_3864);
nand U4445 (N_4445,N_3806,N_3815);
or U4446 (N_4446,N_3571,N_3930);
or U4447 (N_4447,N_3776,N_3553);
nand U4448 (N_4448,N_3393,N_3235);
xor U4449 (N_4449,N_3082,N_3136);
nand U4450 (N_4450,N_3960,N_3824);
and U4451 (N_4451,N_3730,N_3228);
xor U4452 (N_4452,N_3237,N_3259);
xor U4453 (N_4453,N_3928,N_3577);
nor U4454 (N_4454,N_3462,N_3974);
nand U4455 (N_4455,N_3152,N_3849);
nand U4456 (N_4456,N_3315,N_3042);
xor U4457 (N_4457,N_3198,N_3118);
xnor U4458 (N_4458,N_3191,N_3986);
or U4459 (N_4459,N_3374,N_3104);
nor U4460 (N_4460,N_3456,N_3878);
nor U4461 (N_4461,N_3037,N_3110);
nor U4462 (N_4462,N_3982,N_3401);
nor U4463 (N_4463,N_3873,N_3574);
xor U4464 (N_4464,N_3568,N_3740);
nor U4465 (N_4465,N_3321,N_3533);
or U4466 (N_4466,N_3341,N_3619);
nand U4467 (N_4467,N_3745,N_3843);
nor U4468 (N_4468,N_3544,N_3085);
nand U4469 (N_4469,N_3632,N_3466);
nor U4470 (N_4470,N_3814,N_3611);
and U4471 (N_4471,N_3425,N_3275);
nor U4472 (N_4472,N_3944,N_3642);
nor U4473 (N_4473,N_3463,N_3742);
nand U4474 (N_4474,N_3991,N_3603);
or U4475 (N_4475,N_3734,N_3943);
nand U4476 (N_4476,N_3952,N_3798);
and U4477 (N_4477,N_3641,N_3931);
nor U4478 (N_4478,N_3181,N_3484);
and U4479 (N_4479,N_3399,N_3724);
nor U4480 (N_4480,N_3369,N_3676);
xor U4481 (N_4481,N_3242,N_3444);
nor U4482 (N_4482,N_3555,N_3269);
nand U4483 (N_4483,N_3937,N_3552);
nor U4484 (N_4484,N_3459,N_3626);
xnor U4485 (N_4485,N_3792,N_3539);
or U4486 (N_4486,N_3077,N_3286);
nor U4487 (N_4487,N_3821,N_3219);
and U4488 (N_4488,N_3970,N_3681);
nor U4489 (N_4489,N_3358,N_3706);
and U4490 (N_4490,N_3258,N_3069);
nor U4491 (N_4491,N_3099,N_3106);
or U4492 (N_4492,N_3008,N_3236);
nand U4493 (N_4493,N_3576,N_3014);
xnor U4494 (N_4494,N_3760,N_3138);
or U4495 (N_4495,N_3368,N_3257);
xnor U4496 (N_4496,N_3493,N_3567);
and U4497 (N_4497,N_3656,N_3978);
nor U4498 (N_4498,N_3892,N_3754);
xnor U4499 (N_4499,N_3144,N_3122);
or U4500 (N_4500,N_3027,N_3148);
and U4501 (N_4501,N_3818,N_3085);
or U4502 (N_4502,N_3933,N_3918);
nand U4503 (N_4503,N_3374,N_3829);
and U4504 (N_4504,N_3197,N_3569);
xnor U4505 (N_4505,N_3464,N_3404);
nand U4506 (N_4506,N_3797,N_3512);
nor U4507 (N_4507,N_3344,N_3345);
nor U4508 (N_4508,N_3871,N_3049);
nand U4509 (N_4509,N_3297,N_3115);
nor U4510 (N_4510,N_3564,N_3375);
and U4511 (N_4511,N_3581,N_3164);
nor U4512 (N_4512,N_3439,N_3397);
and U4513 (N_4513,N_3311,N_3961);
nor U4514 (N_4514,N_3854,N_3246);
xnor U4515 (N_4515,N_3703,N_3686);
nand U4516 (N_4516,N_3569,N_3131);
nor U4517 (N_4517,N_3006,N_3698);
xor U4518 (N_4518,N_3686,N_3413);
xnor U4519 (N_4519,N_3560,N_3600);
or U4520 (N_4520,N_3976,N_3651);
and U4521 (N_4521,N_3325,N_3938);
nand U4522 (N_4522,N_3620,N_3920);
nand U4523 (N_4523,N_3097,N_3638);
xor U4524 (N_4524,N_3542,N_3590);
nand U4525 (N_4525,N_3011,N_3922);
xnor U4526 (N_4526,N_3059,N_3274);
nor U4527 (N_4527,N_3247,N_3256);
and U4528 (N_4528,N_3020,N_3538);
nand U4529 (N_4529,N_3913,N_3365);
or U4530 (N_4530,N_3092,N_3570);
nor U4531 (N_4531,N_3222,N_3962);
nor U4532 (N_4532,N_3945,N_3066);
nand U4533 (N_4533,N_3709,N_3277);
nor U4534 (N_4534,N_3269,N_3400);
or U4535 (N_4535,N_3321,N_3691);
nand U4536 (N_4536,N_3768,N_3904);
or U4537 (N_4537,N_3869,N_3362);
nor U4538 (N_4538,N_3745,N_3174);
and U4539 (N_4539,N_3324,N_3692);
nand U4540 (N_4540,N_3403,N_3342);
or U4541 (N_4541,N_3316,N_3843);
nor U4542 (N_4542,N_3825,N_3729);
and U4543 (N_4543,N_3599,N_3936);
xnor U4544 (N_4544,N_3605,N_3500);
and U4545 (N_4545,N_3425,N_3827);
nand U4546 (N_4546,N_3575,N_3839);
nand U4547 (N_4547,N_3144,N_3929);
nor U4548 (N_4548,N_3757,N_3309);
nand U4549 (N_4549,N_3713,N_3891);
and U4550 (N_4550,N_3942,N_3458);
nand U4551 (N_4551,N_3134,N_3239);
nor U4552 (N_4552,N_3615,N_3093);
or U4553 (N_4553,N_3896,N_3637);
and U4554 (N_4554,N_3105,N_3048);
or U4555 (N_4555,N_3083,N_3507);
or U4556 (N_4556,N_3468,N_3175);
or U4557 (N_4557,N_3624,N_3837);
or U4558 (N_4558,N_3093,N_3810);
xor U4559 (N_4559,N_3878,N_3926);
and U4560 (N_4560,N_3359,N_3776);
nor U4561 (N_4561,N_3861,N_3027);
and U4562 (N_4562,N_3638,N_3992);
nand U4563 (N_4563,N_3969,N_3604);
and U4564 (N_4564,N_3985,N_3006);
nor U4565 (N_4565,N_3567,N_3809);
xnor U4566 (N_4566,N_3138,N_3991);
xor U4567 (N_4567,N_3328,N_3539);
xnor U4568 (N_4568,N_3817,N_3691);
xor U4569 (N_4569,N_3535,N_3321);
nand U4570 (N_4570,N_3855,N_3731);
or U4571 (N_4571,N_3857,N_3395);
and U4572 (N_4572,N_3476,N_3251);
nand U4573 (N_4573,N_3421,N_3560);
or U4574 (N_4574,N_3364,N_3514);
nand U4575 (N_4575,N_3121,N_3927);
nand U4576 (N_4576,N_3370,N_3944);
and U4577 (N_4577,N_3921,N_3738);
nand U4578 (N_4578,N_3222,N_3175);
nand U4579 (N_4579,N_3397,N_3056);
nand U4580 (N_4580,N_3029,N_3465);
or U4581 (N_4581,N_3975,N_3536);
or U4582 (N_4582,N_3863,N_3090);
nand U4583 (N_4583,N_3195,N_3089);
nand U4584 (N_4584,N_3653,N_3894);
nor U4585 (N_4585,N_3582,N_3344);
nand U4586 (N_4586,N_3014,N_3842);
or U4587 (N_4587,N_3623,N_3022);
nor U4588 (N_4588,N_3031,N_3839);
nand U4589 (N_4589,N_3837,N_3138);
and U4590 (N_4590,N_3872,N_3217);
xnor U4591 (N_4591,N_3846,N_3682);
xor U4592 (N_4592,N_3486,N_3656);
and U4593 (N_4593,N_3283,N_3962);
or U4594 (N_4594,N_3417,N_3111);
xnor U4595 (N_4595,N_3562,N_3448);
nor U4596 (N_4596,N_3688,N_3898);
nor U4597 (N_4597,N_3866,N_3184);
nand U4598 (N_4598,N_3566,N_3853);
and U4599 (N_4599,N_3851,N_3273);
xnor U4600 (N_4600,N_3623,N_3084);
nand U4601 (N_4601,N_3337,N_3925);
xor U4602 (N_4602,N_3302,N_3133);
nand U4603 (N_4603,N_3533,N_3306);
xnor U4604 (N_4604,N_3220,N_3474);
or U4605 (N_4605,N_3531,N_3808);
nor U4606 (N_4606,N_3809,N_3187);
nand U4607 (N_4607,N_3428,N_3796);
nor U4608 (N_4608,N_3233,N_3912);
nand U4609 (N_4609,N_3011,N_3024);
and U4610 (N_4610,N_3609,N_3241);
or U4611 (N_4611,N_3631,N_3720);
and U4612 (N_4612,N_3161,N_3050);
or U4613 (N_4613,N_3178,N_3648);
nor U4614 (N_4614,N_3703,N_3389);
and U4615 (N_4615,N_3520,N_3953);
nand U4616 (N_4616,N_3748,N_3216);
nor U4617 (N_4617,N_3292,N_3951);
or U4618 (N_4618,N_3686,N_3272);
nand U4619 (N_4619,N_3726,N_3400);
or U4620 (N_4620,N_3531,N_3039);
or U4621 (N_4621,N_3641,N_3155);
nor U4622 (N_4622,N_3387,N_3153);
nand U4623 (N_4623,N_3885,N_3426);
nand U4624 (N_4624,N_3699,N_3531);
and U4625 (N_4625,N_3342,N_3154);
xnor U4626 (N_4626,N_3146,N_3984);
nor U4627 (N_4627,N_3004,N_3728);
nand U4628 (N_4628,N_3202,N_3369);
xor U4629 (N_4629,N_3168,N_3971);
nand U4630 (N_4630,N_3078,N_3346);
and U4631 (N_4631,N_3363,N_3233);
and U4632 (N_4632,N_3556,N_3830);
and U4633 (N_4633,N_3487,N_3464);
or U4634 (N_4634,N_3717,N_3503);
and U4635 (N_4635,N_3034,N_3302);
or U4636 (N_4636,N_3692,N_3529);
xor U4637 (N_4637,N_3084,N_3491);
and U4638 (N_4638,N_3389,N_3459);
xor U4639 (N_4639,N_3790,N_3830);
and U4640 (N_4640,N_3646,N_3206);
and U4641 (N_4641,N_3559,N_3840);
nand U4642 (N_4642,N_3092,N_3515);
and U4643 (N_4643,N_3051,N_3430);
or U4644 (N_4644,N_3733,N_3421);
nor U4645 (N_4645,N_3077,N_3226);
nand U4646 (N_4646,N_3831,N_3263);
and U4647 (N_4647,N_3210,N_3182);
nor U4648 (N_4648,N_3143,N_3125);
and U4649 (N_4649,N_3946,N_3590);
and U4650 (N_4650,N_3288,N_3534);
xor U4651 (N_4651,N_3344,N_3916);
xor U4652 (N_4652,N_3300,N_3022);
and U4653 (N_4653,N_3076,N_3360);
xnor U4654 (N_4654,N_3137,N_3484);
nor U4655 (N_4655,N_3067,N_3038);
and U4656 (N_4656,N_3548,N_3924);
and U4657 (N_4657,N_3354,N_3408);
or U4658 (N_4658,N_3420,N_3820);
or U4659 (N_4659,N_3556,N_3764);
nand U4660 (N_4660,N_3138,N_3057);
nand U4661 (N_4661,N_3219,N_3807);
or U4662 (N_4662,N_3220,N_3936);
nor U4663 (N_4663,N_3902,N_3135);
xnor U4664 (N_4664,N_3849,N_3877);
nor U4665 (N_4665,N_3296,N_3448);
xnor U4666 (N_4666,N_3091,N_3412);
and U4667 (N_4667,N_3789,N_3713);
or U4668 (N_4668,N_3069,N_3698);
and U4669 (N_4669,N_3016,N_3024);
xor U4670 (N_4670,N_3366,N_3546);
xnor U4671 (N_4671,N_3761,N_3013);
xnor U4672 (N_4672,N_3703,N_3744);
nor U4673 (N_4673,N_3014,N_3698);
nand U4674 (N_4674,N_3614,N_3034);
or U4675 (N_4675,N_3146,N_3662);
and U4676 (N_4676,N_3660,N_3698);
and U4677 (N_4677,N_3154,N_3066);
nor U4678 (N_4678,N_3158,N_3149);
nand U4679 (N_4679,N_3482,N_3687);
or U4680 (N_4680,N_3222,N_3978);
nor U4681 (N_4681,N_3441,N_3110);
or U4682 (N_4682,N_3658,N_3710);
or U4683 (N_4683,N_3500,N_3308);
nor U4684 (N_4684,N_3611,N_3020);
nand U4685 (N_4685,N_3365,N_3230);
nand U4686 (N_4686,N_3647,N_3716);
nand U4687 (N_4687,N_3136,N_3289);
or U4688 (N_4688,N_3073,N_3729);
xor U4689 (N_4689,N_3998,N_3797);
xnor U4690 (N_4690,N_3622,N_3021);
nor U4691 (N_4691,N_3081,N_3621);
nand U4692 (N_4692,N_3279,N_3585);
xnor U4693 (N_4693,N_3109,N_3515);
and U4694 (N_4694,N_3734,N_3132);
nor U4695 (N_4695,N_3237,N_3506);
and U4696 (N_4696,N_3460,N_3981);
xnor U4697 (N_4697,N_3015,N_3016);
nor U4698 (N_4698,N_3821,N_3383);
nor U4699 (N_4699,N_3090,N_3062);
or U4700 (N_4700,N_3889,N_3618);
or U4701 (N_4701,N_3560,N_3212);
nor U4702 (N_4702,N_3426,N_3059);
nor U4703 (N_4703,N_3139,N_3493);
nor U4704 (N_4704,N_3700,N_3694);
xnor U4705 (N_4705,N_3221,N_3233);
and U4706 (N_4706,N_3498,N_3358);
and U4707 (N_4707,N_3371,N_3833);
or U4708 (N_4708,N_3047,N_3597);
and U4709 (N_4709,N_3334,N_3037);
xor U4710 (N_4710,N_3396,N_3200);
and U4711 (N_4711,N_3649,N_3419);
or U4712 (N_4712,N_3933,N_3295);
and U4713 (N_4713,N_3291,N_3365);
xor U4714 (N_4714,N_3528,N_3792);
xor U4715 (N_4715,N_3155,N_3579);
or U4716 (N_4716,N_3403,N_3130);
xor U4717 (N_4717,N_3305,N_3170);
and U4718 (N_4718,N_3780,N_3138);
and U4719 (N_4719,N_3465,N_3370);
xnor U4720 (N_4720,N_3578,N_3063);
nand U4721 (N_4721,N_3462,N_3069);
nand U4722 (N_4722,N_3155,N_3673);
nor U4723 (N_4723,N_3920,N_3704);
or U4724 (N_4724,N_3173,N_3283);
nand U4725 (N_4725,N_3188,N_3501);
xor U4726 (N_4726,N_3318,N_3740);
nand U4727 (N_4727,N_3301,N_3407);
or U4728 (N_4728,N_3346,N_3869);
or U4729 (N_4729,N_3038,N_3306);
and U4730 (N_4730,N_3024,N_3466);
nor U4731 (N_4731,N_3936,N_3282);
nor U4732 (N_4732,N_3885,N_3322);
nor U4733 (N_4733,N_3921,N_3193);
nand U4734 (N_4734,N_3093,N_3627);
and U4735 (N_4735,N_3151,N_3078);
nor U4736 (N_4736,N_3894,N_3760);
or U4737 (N_4737,N_3606,N_3556);
nand U4738 (N_4738,N_3048,N_3453);
xor U4739 (N_4739,N_3756,N_3554);
xor U4740 (N_4740,N_3081,N_3128);
and U4741 (N_4741,N_3054,N_3504);
and U4742 (N_4742,N_3956,N_3824);
nor U4743 (N_4743,N_3341,N_3026);
and U4744 (N_4744,N_3246,N_3580);
xnor U4745 (N_4745,N_3806,N_3996);
nor U4746 (N_4746,N_3444,N_3892);
and U4747 (N_4747,N_3356,N_3609);
or U4748 (N_4748,N_3896,N_3675);
xor U4749 (N_4749,N_3389,N_3306);
xor U4750 (N_4750,N_3510,N_3313);
or U4751 (N_4751,N_3857,N_3220);
xnor U4752 (N_4752,N_3833,N_3108);
xor U4753 (N_4753,N_3570,N_3256);
xor U4754 (N_4754,N_3563,N_3854);
nand U4755 (N_4755,N_3789,N_3605);
or U4756 (N_4756,N_3340,N_3919);
nand U4757 (N_4757,N_3513,N_3645);
nand U4758 (N_4758,N_3844,N_3952);
nor U4759 (N_4759,N_3221,N_3613);
xnor U4760 (N_4760,N_3481,N_3618);
xor U4761 (N_4761,N_3338,N_3994);
and U4762 (N_4762,N_3021,N_3630);
xnor U4763 (N_4763,N_3561,N_3129);
nor U4764 (N_4764,N_3262,N_3980);
and U4765 (N_4765,N_3185,N_3676);
or U4766 (N_4766,N_3850,N_3794);
or U4767 (N_4767,N_3467,N_3830);
xnor U4768 (N_4768,N_3523,N_3873);
or U4769 (N_4769,N_3005,N_3476);
or U4770 (N_4770,N_3823,N_3063);
nor U4771 (N_4771,N_3544,N_3266);
xnor U4772 (N_4772,N_3665,N_3780);
or U4773 (N_4773,N_3354,N_3027);
and U4774 (N_4774,N_3525,N_3818);
nor U4775 (N_4775,N_3193,N_3230);
nor U4776 (N_4776,N_3025,N_3829);
nand U4777 (N_4777,N_3934,N_3209);
nand U4778 (N_4778,N_3015,N_3921);
or U4779 (N_4779,N_3130,N_3754);
or U4780 (N_4780,N_3651,N_3406);
nand U4781 (N_4781,N_3538,N_3273);
nand U4782 (N_4782,N_3607,N_3720);
nor U4783 (N_4783,N_3507,N_3197);
or U4784 (N_4784,N_3566,N_3376);
nor U4785 (N_4785,N_3657,N_3148);
or U4786 (N_4786,N_3424,N_3862);
xnor U4787 (N_4787,N_3954,N_3719);
and U4788 (N_4788,N_3405,N_3472);
xnor U4789 (N_4789,N_3066,N_3104);
and U4790 (N_4790,N_3382,N_3663);
xor U4791 (N_4791,N_3580,N_3571);
nor U4792 (N_4792,N_3645,N_3809);
xor U4793 (N_4793,N_3703,N_3905);
or U4794 (N_4794,N_3136,N_3776);
xnor U4795 (N_4795,N_3099,N_3176);
or U4796 (N_4796,N_3860,N_3474);
nor U4797 (N_4797,N_3194,N_3671);
nand U4798 (N_4798,N_3697,N_3017);
nor U4799 (N_4799,N_3778,N_3353);
or U4800 (N_4800,N_3079,N_3806);
nand U4801 (N_4801,N_3201,N_3149);
and U4802 (N_4802,N_3639,N_3672);
xnor U4803 (N_4803,N_3734,N_3740);
and U4804 (N_4804,N_3923,N_3052);
nor U4805 (N_4805,N_3455,N_3165);
and U4806 (N_4806,N_3141,N_3354);
or U4807 (N_4807,N_3456,N_3443);
or U4808 (N_4808,N_3670,N_3888);
nor U4809 (N_4809,N_3736,N_3592);
nor U4810 (N_4810,N_3881,N_3013);
and U4811 (N_4811,N_3049,N_3615);
and U4812 (N_4812,N_3131,N_3535);
and U4813 (N_4813,N_3736,N_3354);
nor U4814 (N_4814,N_3142,N_3240);
or U4815 (N_4815,N_3484,N_3184);
nor U4816 (N_4816,N_3733,N_3548);
nand U4817 (N_4817,N_3242,N_3690);
nor U4818 (N_4818,N_3221,N_3803);
xor U4819 (N_4819,N_3440,N_3227);
xor U4820 (N_4820,N_3832,N_3489);
xnor U4821 (N_4821,N_3690,N_3949);
or U4822 (N_4822,N_3124,N_3316);
nor U4823 (N_4823,N_3491,N_3034);
xnor U4824 (N_4824,N_3332,N_3402);
or U4825 (N_4825,N_3655,N_3451);
nor U4826 (N_4826,N_3817,N_3372);
and U4827 (N_4827,N_3412,N_3503);
and U4828 (N_4828,N_3026,N_3860);
xor U4829 (N_4829,N_3826,N_3671);
or U4830 (N_4830,N_3970,N_3267);
nand U4831 (N_4831,N_3334,N_3868);
and U4832 (N_4832,N_3430,N_3883);
nor U4833 (N_4833,N_3304,N_3520);
xor U4834 (N_4834,N_3584,N_3918);
and U4835 (N_4835,N_3869,N_3696);
or U4836 (N_4836,N_3120,N_3691);
nand U4837 (N_4837,N_3783,N_3873);
nor U4838 (N_4838,N_3941,N_3870);
or U4839 (N_4839,N_3448,N_3102);
xor U4840 (N_4840,N_3999,N_3327);
or U4841 (N_4841,N_3661,N_3618);
nor U4842 (N_4842,N_3518,N_3018);
nor U4843 (N_4843,N_3860,N_3541);
nor U4844 (N_4844,N_3774,N_3456);
nor U4845 (N_4845,N_3229,N_3395);
and U4846 (N_4846,N_3941,N_3197);
and U4847 (N_4847,N_3713,N_3950);
nand U4848 (N_4848,N_3771,N_3227);
xor U4849 (N_4849,N_3234,N_3163);
or U4850 (N_4850,N_3694,N_3613);
or U4851 (N_4851,N_3553,N_3134);
and U4852 (N_4852,N_3929,N_3613);
xor U4853 (N_4853,N_3183,N_3443);
xor U4854 (N_4854,N_3979,N_3619);
xnor U4855 (N_4855,N_3965,N_3319);
xor U4856 (N_4856,N_3633,N_3146);
or U4857 (N_4857,N_3150,N_3806);
nand U4858 (N_4858,N_3776,N_3847);
xnor U4859 (N_4859,N_3919,N_3990);
or U4860 (N_4860,N_3045,N_3022);
nor U4861 (N_4861,N_3227,N_3501);
or U4862 (N_4862,N_3652,N_3935);
or U4863 (N_4863,N_3152,N_3121);
xor U4864 (N_4864,N_3691,N_3224);
nor U4865 (N_4865,N_3491,N_3088);
nor U4866 (N_4866,N_3562,N_3877);
or U4867 (N_4867,N_3520,N_3473);
xnor U4868 (N_4868,N_3868,N_3631);
and U4869 (N_4869,N_3859,N_3516);
and U4870 (N_4870,N_3783,N_3859);
nand U4871 (N_4871,N_3864,N_3771);
or U4872 (N_4872,N_3350,N_3733);
nand U4873 (N_4873,N_3784,N_3138);
nand U4874 (N_4874,N_3320,N_3151);
nor U4875 (N_4875,N_3983,N_3720);
xor U4876 (N_4876,N_3923,N_3756);
and U4877 (N_4877,N_3327,N_3243);
nand U4878 (N_4878,N_3562,N_3793);
or U4879 (N_4879,N_3623,N_3846);
xnor U4880 (N_4880,N_3255,N_3774);
xor U4881 (N_4881,N_3141,N_3965);
nor U4882 (N_4882,N_3143,N_3336);
nand U4883 (N_4883,N_3667,N_3341);
nor U4884 (N_4884,N_3607,N_3826);
and U4885 (N_4885,N_3803,N_3894);
or U4886 (N_4886,N_3061,N_3320);
and U4887 (N_4887,N_3523,N_3791);
and U4888 (N_4888,N_3582,N_3697);
nand U4889 (N_4889,N_3965,N_3398);
nand U4890 (N_4890,N_3676,N_3510);
and U4891 (N_4891,N_3843,N_3245);
nor U4892 (N_4892,N_3788,N_3637);
nor U4893 (N_4893,N_3309,N_3425);
nand U4894 (N_4894,N_3678,N_3033);
nor U4895 (N_4895,N_3040,N_3321);
nor U4896 (N_4896,N_3937,N_3638);
nor U4897 (N_4897,N_3163,N_3558);
and U4898 (N_4898,N_3685,N_3575);
nand U4899 (N_4899,N_3705,N_3978);
xor U4900 (N_4900,N_3379,N_3892);
nor U4901 (N_4901,N_3450,N_3063);
and U4902 (N_4902,N_3597,N_3965);
or U4903 (N_4903,N_3374,N_3057);
and U4904 (N_4904,N_3229,N_3938);
nand U4905 (N_4905,N_3875,N_3612);
xor U4906 (N_4906,N_3488,N_3858);
or U4907 (N_4907,N_3883,N_3622);
or U4908 (N_4908,N_3646,N_3823);
nor U4909 (N_4909,N_3188,N_3939);
nor U4910 (N_4910,N_3883,N_3315);
xnor U4911 (N_4911,N_3632,N_3958);
nand U4912 (N_4912,N_3036,N_3279);
or U4913 (N_4913,N_3164,N_3218);
xor U4914 (N_4914,N_3436,N_3927);
nand U4915 (N_4915,N_3561,N_3781);
and U4916 (N_4916,N_3687,N_3153);
xor U4917 (N_4917,N_3848,N_3090);
or U4918 (N_4918,N_3554,N_3635);
nand U4919 (N_4919,N_3528,N_3904);
and U4920 (N_4920,N_3806,N_3985);
nand U4921 (N_4921,N_3357,N_3370);
and U4922 (N_4922,N_3224,N_3397);
or U4923 (N_4923,N_3529,N_3153);
xor U4924 (N_4924,N_3680,N_3739);
nand U4925 (N_4925,N_3681,N_3675);
xnor U4926 (N_4926,N_3172,N_3197);
nor U4927 (N_4927,N_3889,N_3215);
xnor U4928 (N_4928,N_3462,N_3871);
nor U4929 (N_4929,N_3040,N_3724);
or U4930 (N_4930,N_3487,N_3735);
or U4931 (N_4931,N_3257,N_3241);
nor U4932 (N_4932,N_3628,N_3707);
or U4933 (N_4933,N_3412,N_3349);
or U4934 (N_4934,N_3176,N_3271);
xor U4935 (N_4935,N_3555,N_3305);
nor U4936 (N_4936,N_3961,N_3929);
and U4937 (N_4937,N_3101,N_3767);
xor U4938 (N_4938,N_3092,N_3149);
and U4939 (N_4939,N_3349,N_3130);
nand U4940 (N_4940,N_3274,N_3815);
nor U4941 (N_4941,N_3895,N_3194);
nor U4942 (N_4942,N_3783,N_3399);
or U4943 (N_4943,N_3158,N_3752);
xnor U4944 (N_4944,N_3038,N_3660);
nand U4945 (N_4945,N_3035,N_3874);
or U4946 (N_4946,N_3100,N_3150);
and U4947 (N_4947,N_3039,N_3176);
or U4948 (N_4948,N_3663,N_3443);
xnor U4949 (N_4949,N_3357,N_3425);
nand U4950 (N_4950,N_3441,N_3340);
xnor U4951 (N_4951,N_3285,N_3648);
and U4952 (N_4952,N_3530,N_3035);
nand U4953 (N_4953,N_3033,N_3974);
and U4954 (N_4954,N_3669,N_3815);
or U4955 (N_4955,N_3072,N_3567);
nor U4956 (N_4956,N_3541,N_3664);
xor U4957 (N_4957,N_3166,N_3779);
and U4958 (N_4958,N_3293,N_3043);
nor U4959 (N_4959,N_3319,N_3486);
or U4960 (N_4960,N_3600,N_3077);
and U4961 (N_4961,N_3555,N_3993);
nand U4962 (N_4962,N_3235,N_3575);
nand U4963 (N_4963,N_3207,N_3306);
xor U4964 (N_4964,N_3157,N_3401);
nor U4965 (N_4965,N_3222,N_3738);
and U4966 (N_4966,N_3267,N_3725);
nand U4967 (N_4967,N_3124,N_3591);
nor U4968 (N_4968,N_3251,N_3156);
nand U4969 (N_4969,N_3465,N_3517);
xor U4970 (N_4970,N_3333,N_3041);
nor U4971 (N_4971,N_3453,N_3012);
or U4972 (N_4972,N_3308,N_3000);
and U4973 (N_4973,N_3332,N_3173);
and U4974 (N_4974,N_3781,N_3598);
nor U4975 (N_4975,N_3509,N_3645);
or U4976 (N_4976,N_3077,N_3953);
or U4977 (N_4977,N_3173,N_3606);
xor U4978 (N_4978,N_3940,N_3700);
nor U4979 (N_4979,N_3366,N_3043);
xnor U4980 (N_4980,N_3681,N_3764);
or U4981 (N_4981,N_3995,N_3075);
nor U4982 (N_4982,N_3973,N_3194);
or U4983 (N_4983,N_3041,N_3837);
or U4984 (N_4984,N_3682,N_3818);
xnor U4985 (N_4985,N_3344,N_3456);
and U4986 (N_4986,N_3576,N_3570);
and U4987 (N_4987,N_3287,N_3402);
nand U4988 (N_4988,N_3585,N_3258);
nor U4989 (N_4989,N_3171,N_3812);
nor U4990 (N_4990,N_3783,N_3368);
and U4991 (N_4991,N_3332,N_3648);
and U4992 (N_4992,N_3758,N_3112);
nor U4993 (N_4993,N_3424,N_3410);
or U4994 (N_4994,N_3716,N_3844);
xor U4995 (N_4995,N_3514,N_3396);
nand U4996 (N_4996,N_3024,N_3490);
and U4997 (N_4997,N_3112,N_3593);
or U4998 (N_4998,N_3881,N_3499);
nand U4999 (N_4999,N_3424,N_3941);
or UO_0 (O_0,N_4528,N_4506);
xnor UO_1 (O_1,N_4573,N_4933);
and UO_2 (O_2,N_4085,N_4433);
or UO_3 (O_3,N_4389,N_4436);
and UO_4 (O_4,N_4668,N_4799);
xor UO_5 (O_5,N_4257,N_4534);
nor UO_6 (O_6,N_4700,N_4677);
and UO_7 (O_7,N_4357,N_4275);
nand UO_8 (O_8,N_4602,N_4443);
nor UO_9 (O_9,N_4122,N_4977);
xor UO_10 (O_10,N_4484,N_4081);
and UO_11 (O_11,N_4398,N_4810);
nor UO_12 (O_12,N_4335,N_4816);
and UO_13 (O_13,N_4806,N_4208);
or UO_14 (O_14,N_4138,N_4464);
nand UO_15 (O_15,N_4059,N_4315);
nor UO_16 (O_16,N_4246,N_4729);
nand UO_17 (O_17,N_4957,N_4211);
xnor UO_18 (O_18,N_4642,N_4260);
or UO_19 (O_19,N_4541,N_4570);
xor UO_20 (O_20,N_4304,N_4886);
nand UO_21 (O_21,N_4838,N_4905);
and UO_22 (O_22,N_4297,N_4007);
or UO_23 (O_23,N_4423,N_4213);
and UO_24 (O_24,N_4497,N_4430);
nor UO_25 (O_25,N_4451,N_4225);
nand UO_26 (O_26,N_4687,N_4409);
nand UO_27 (O_27,N_4117,N_4285);
and UO_28 (O_28,N_4083,N_4148);
or UO_29 (O_29,N_4751,N_4858);
or UO_30 (O_30,N_4281,N_4498);
and UO_31 (O_31,N_4545,N_4851);
or UO_32 (O_32,N_4108,N_4476);
nor UO_33 (O_33,N_4188,N_4600);
and UO_34 (O_34,N_4419,N_4267);
and UO_35 (O_35,N_4948,N_4546);
and UO_36 (O_36,N_4215,N_4292);
nand UO_37 (O_37,N_4701,N_4301);
nand UO_38 (O_38,N_4030,N_4031);
or UO_39 (O_39,N_4171,N_4596);
nor UO_40 (O_40,N_4808,N_4356);
or UO_41 (O_41,N_4716,N_4090);
or UO_42 (O_42,N_4587,N_4462);
or UO_43 (O_43,N_4403,N_4432);
or UO_44 (O_44,N_4441,N_4790);
nand UO_45 (O_45,N_4341,N_4949);
and UO_46 (O_46,N_4204,N_4488);
nor UO_47 (O_47,N_4152,N_4954);
nand UO_48 (O_48,N_4177,N_4008);
and UO_49 (O_49,N_4973,N_4458);
nand UO_50 (O_50,N_4976,N_4683);
nand UO_51 (O_51,N_4864,N_4725);
xnor UO_52 (O_52,N_4053,N_4487);
or UO_53 (O_53,N_4652,N_4503);
nand UO_54 (O_54,N_4351,N_4712);
nor UO_55 (O_55,N_4057,N_4502);
xor UO_56 (O_56,N_4576,N_4040);
nor UO_57 (O_57,N_4704,N_4418);
xnor UO_58 (O_58,N_4453,N_4722);
and UO_59 (O_59,N_4765,N_4468);
or UO_60 (O_60,N_4159,N_4149);
nor UO_61 (O_61,N_4598,N_4906);
and UO_62 (O_62,N_4183,N_4140);
or UO_63 (O_63,N_4003,N_4200);
nor UO_64 (O_64,N_4565,N_4965);
or UO_65 (O_65,N_4147,N_4508);
and UO_66 (O_66,N_4944,N_4477);
or UO_67 (O_67,N_4406,N_4187);
xnor UO_68 (O_68,N_4364,N_4789);
nand UO_69 (O_69,N_4936,N_4524);
nor UO_70 (O_70,N_4029,N_4308);
or UO_71 (O_71,N_4309,N_4220);
nor UO_72 (O_72,N_4656,N_4034);
or UO_73 (O_73,N_4265,N_4532);
xnor UO_74 (O_74,N_4795,N_4313);
nand UO_75 (O_75,N_4161,N_4150);
nor UO_76 (O_76,N_4794,N_4077);
or UO_77 (O_77,N_4037,N_4111);
and UO_78 (O_78,N_4050,N_4793);
or UO_79 (O_79,N_4055,N_4624);
nand UO_80 (O_80,N_4647,N_4619);
nand UO_81 (O_81,N_4785,N_4499);
nor UO_82 (O_82,N_4222,N_4277);
nor UO_83 (O_83,N_4036,N_4852);
nand UO_84 (O_84,N_4123,N_4244);
nand UO_85 (O_85,N_4900,N_4721);
nand UO_86 (O_86,N_4504,N_4256);
nor UO_87 (O_87,N_4153,N_4763);
and UO_88 (O_88,N_4469,N_4828);
or UO_89 (O_89,N_4889,N_4746);
or UO_90 (O_90,N_4294,N_4583);
nor UO_91 (O_91,N_4616,N_4233);
or UO_92 (O_92,N_4110,N_4875);
xnor UO_93 (O_93,N_4466,N_4378);
and UO_94 (O_94,N_4730,N_4412);
nor UO_95 (O_95,N_4100,N_4747);
or UO_96 (O_96,N_4955,N_4132);
or UO_97 (O_97,N_4585,N_4800);
nor UO_98 (O_98,N_4058,N_4359);
and UO_99 (O_99,N_4788,N_4447);
nor UO_100 (O_100,N_4253,N_4556);
and UO_101 (O_101,N_4952,N_4563);
nand UO_102 (O_102,N_4286,N_4971);
nand UO_103 (O_103,N_4329,N_4099);
and UO_104 (O_104,N_4218,N_4792);
xor UO_105 (O_105,N_4066,N_4597);
or UO_106 (O_106,N_4385,N_4612);
and UO_107 (O_107,N_4599,N_4841);
and UO_108 (O_108,N_4494,N_4734);
or UO_109 (O_109,N_4143,N_4630);
xor UO_110 (O_110,N_4996,N_4234);
and UO_111 (O_111,N_4879,N_4925);
xor UO_112 (O_112,N_4743,N_4368);
nand UO_113 (O_113,N_4410,N_4820);
xnor UO_114 (O_114,N_4653,N_4861);
nor UO_115 (O_115,N_4614,N_4766);
nor UO_116 (O_116,N_4891,N_4515);
nand UO_117 (O_117,N_4495,N_4421);
and UO_118 (O_118,N_4089,N_4622);
nand UO_119 (O_119,N_4424,N_4740);
or UO_120 (O_120,N_4843,N_4617);
or UO_121 (O_121,N_4467,N_4779);
nor UO_122 (O_122,N_4103,N_4426);
and UO_123 (O_123,N_4369,N_4849);
or UO_124 (O_124,N_4399,N_4786);
and UO_125 (O_125,N_4860,N_4376);
and UO_126 (O_126,N_4101,N_4978);
or UO_127 (O_127,N_4920,N_4454);
xnor UO_128 (O_128,N_4582,N_4913);
nand UO_129 (O_129,N_4755,N_4829);
nand UO_130 (O_130,N_4017,N_4198);
nor UO_131 (O_131,N_4832,N_4366);
nor UO_132 (O_132,N_4492,N_4073);
and UO_133 (O_133,N_4691,N_4873);
nor UO_134 (O_134,N_4678,N_4427);
or UO_135 (O_135,N_4760,N_4692);
nand UO_136 (O_136,N_4210,N_4555);
xor UO_137 (O_137,N_4529,N_4732);
and UO_138 (O_138,N_4516,N_4380);
or UO_139 (O_139,N_4510,N_4631);
nor UO_140 (O_140,N_4223,N_4295);
or UO_141 (O_141,N_4347,N_4137);
nor UO_142 (O_142,N_4221,N_4240);
nand UO_143 (O_143,N_4390,N_4154);
nand UO_144 (O_144,N_4757,N_4697);
xor UO_145 (O_145,N_4088,N_4848);
xor UO_146 (O_146,N_4553,N_4833);
or UO_147 (O_147,N_4217,N_4823);
nand UO_148 (O_148,N_4394,N_4741);
nand UO_149 (O_149,N_4259,N_4518);
nor UO_150 (O_150,N_4042,N_4658);
xor UO_151 (O_151,N_4781,N_4190);
and UO_152 (O_152,N_4871,N_4916);
nor UO_153 (O_153,N_4770,N_4325);
xor UO_154 (O_154,N_4999,N_4890);
nand UO_155 (O_155,N_4937,N_4715);
nand UO_156 (O_156,N_4056,N_4514);
nand UO_157 (O_157,N_4595,N_4162);
nand UO_158 (O_158,N_4735,N_4919);
or UO_159 (O_159,N_4877,N_4382);
xor UO_160 (O_160,N_4887,N_4374);
xnor UO_161 (O_161,N_4500,N_4588);
xnor UO_162 (O_162,N_4486,N_4431);
nor UO_163 (O_163,N_4513,N_4951);
nor UO_164 (O_164,N_4242,N_4850);
or UO_165 (O_165,N_4826,N_4362);
and UO_166 (O_166,N_4112,N_4386);
nand UO_167 (O_167,N_4191,N_4472);
nand UO_168 (O_168,N_4284,N_4184);
or UO_169 (O_169,N_4186,N_4878);
nand UO_170 (O_170,N_4523,N_4621);
xor UO_171 (O_171,N_4474,N_4736);
and UO_172 (O_172,N_4096,N_4455);
nor UO_173 (O_173,N_4611,N_4011);
nand UO_174 (O_174,N_4530,N_4460);
nor UO_175 (O_175,N_4094,N_4323);
and UO_176 (O_176,N_4839,N_4459);
and UO_177 (O_177,N_4173,N_4146);
nor UO_178 (O_178,N_4870,N_4067);
and UO_179 (O_179,N_4239,N_4927);
or UO_180 (O_180,N_4807,N_4568);
and UO_181 (O_181,N_4899,N_4342);
xnor UO_182 (O_182,N_4991,N_4932);
nand UO_183 (O_183,N_4607,N_4522);
xnor UO_184 (O_184,N_4327,N_4139);
xor UO_185 (O_185,N_4776,N_4646);
nor UO_186 (O_186,N_4194,N_4212);
xor UO_187 (O_187,N_4869,N_4547);
nand UO_188 (O_188,N_4422,N_4535);
nand UO_189 (O_189,N_4288,N_4872);
or UO_190 (O_190,N_4645,N_4482);
nor UO_191 (O_191,N_4511,N_4332);
nand UO_192 (O_192,N_4728,N_4237);
nor UO_193 (O_193,N_4276,N_4046);
xor UO_194 (O_194,N_4783,N_4328);
nor UO_195 (O_195,N_4425,N_4947);
or UO_196 (O_196,N_4798,N_4330);
nor UO_197 (O_197,N_4461,N_4279);
nand UO_198 (O_198,N_4671,N_4192);
or UO_199 (O_199,N_4758,N_4226);
nor UO_200 (O_200,N_4337,N_4501);
nor UO_201 (O_201,N_4026,N_4604);
or UO_202 (O_202,N_4307,N_4033);
and UO_203 (O_203,N_4940,N_4819);
and UO_204 (O_204,N_4505,N_4481);
and UO_205 (O_205,N_4075,N_4102);
and UO_206 (O_206,N_4254,N_4654);
and UO_207 (O_207,N_4322,N_4124);
and UO_208 (O_208,N_4044,N_4980);
nor UO_209 (O_209,N_4303,N_4863);
and UO_210 (O_210,N_4121,N_4283);
or UO_211 (O_211,N_4157,N_4702);
nor UO_212 (O_212,N_4661,N_4338);
nor UO_213 (O_213,N_4274,N_4618);
nand UO_214 (O_214,N_4125,N_4440);
nor UO_215 (O_215,N_4019,N_4216);
nand UO_216 (O_216,N_4623,N_4577);
nand UO_217 (O_217,N_4491,N_4942);
nand UO_218 (O_218,N_4533,N_4723);
xnor UO_219 (O_219,N_4753,N_4012);
or UO_220 (O_220,N_4888,N_4998);
xnor UO_221 (O_221,N_4155,N_4943);
nand UO_222 (O_222,N_4263,N_4857);
and UO_223 (O_223,N_4662,N_4272);
nor UO_224 (O_224,N_4835,N_4560);
nand UO_225 (O_225,N_4252,N_4538);
nor UO_226 (O_226,N_4074,N_4291);
nor UO_227 (O_227,N_4201,N_4854);
or UO_228 (O_228,N_4005,N_4824);
nor UO_229 (O_229,N_4775,N_4749);
and UO_230 (O_230,N_4174,N_4377);
xor UO_231 (O_231,N_4663,N_4639);
and UO_232 (O_232,N_4926,N_4224);
nor UO_233 (O_233,N_4892,N_4293);
and UO_234 (O_234,N_4165,N_4748);
or UO_235 (O_235,N_4797,N_4241);
nand UO_236 (O_236,N_4092,N_4856);
xor UO_237 (O_237,N_4846,N_4710);
nand UO_238 (O_238,N_4950,N_4774);
or UO_239 (O_239,N_4061,N_4685);
nor UO_240 (O_240,N_4446,N_4993);
nand UO_241 (O_241,N_4923,N_4548);
nor UO_242 (O_242,N_4859,N_4724);
nor UO_243 (O_243,N_4444,N_4780);
nor UO_244 (O_244,N_4881,N_4637);
nand UO_245 (O_245,N_4603,N_4756);
or UO_246 (O_246,N_4151,N_4907);
xor UO_247 (O_247,N_4118,N_4842);
and UO_248 (O_248,N_4236,N_4305);
xor UO_249 (O_249,N_4912,N_4214);
nor UO_250 (O_250,N_4674,N_4142);
nand UO_251 (O_251,N_4420,N_4076);
or UO_252 (O_252,N_4115,N_4610);
nor UO_253 (O_253,N_4526,N_4248);
and UO_254 (O_254,N_4428,N_4643);
or UO_255 (O_255,N_4885,N_4694);
nand UO_256 (O_256,N_4311,N_4361);
and UO_257 (O_257,N_4130,N_4627);
or UO_258 (O_258,N_4258,N_4383);
nor UO_259 (O_259,N_4679,N_4733);
and UO_260 (O_260,N_4205,N_4804);
xnor UO_261 (O_261,N_4669,N_4354);
xor UO_262 (O_262,N_4699,N_4365);
or UO_263 (O_263,N_4726,N_4028);
xor UO_264 (O_264,N_4665,N_4401);
xor UO_265 (O_265,N_4967,N_4557);
nand UO_266 (O_266,N_4784,N_4605);
nor UO_267 (O_267,N_4670,N_4994);
and UO_268 (O_268,N_4550,N_4703);
nand UO_269 (O_269,N_4018,N_4648);
nand UO_270 (O_270,N_4986,N_4032);
xnor UO_271 (O_271,N_4634,N_4478);
and UO_272 (O_272,N_4144,N_4915);
or UO_273 (O_273,N_4975,N_4635);
nand UO_274 (O_274,N_4119,N_4371);
nand UO_275 (O_275,N_4025,N_4512);
nand UO_276 (O_276,N_4536,N_4628);
nand UO_277 (O_277,N_4392,N_4827);
and UO_278 (O_278,N_4837,N_4408);
nand UO_279 (O_279,N_4471,N_4475);
and UO_280 (O_280,N_4945,N_4606);
and UO_281 (O_281,N_4717,N_4992);
nor UO_282 (O_282,N_4961,N_4754);
nor UO_283 (O_283,N_4625,N_4742);
xor UO_284 (O_284,N_4960,N_4349);
and UO_285 (O_285,N_4413,N_4688);
or UO_286 (O_286,N_4641,N_4353);
or UO_287 (O_287,N_4189,N_4179);
nand UO_288 (O_288,N_4979,N_4352);
nand UO_289 (O_289,N_4387,N_4289);
xnor UO_290 (O_290,N_4358,N_4015);
nor UO_291 (O_291,N_4882,N_4613);
and UO_292 (O_292,N_4185,N_4227);
or UO_293 (O_293,N_4417,N_4039);
nand UO_294 (O_294,N_4116,N_4230);
nand UO_295 (O_295,N_4867,N_4711);
or UO_296 (O_296,N_4935,N_4038);
nor UO_297 (O_297,N_4862,N_4840);
nand UO_298 (O_298,N_4544,N_4633);
nor UO_299 (O_299,N_4164,N_4300);
nor UO_300 (O_300,N_4035,N_4109);
nor UO_301 (O_301,N_4537,N_4752);
and UO_302 (O_302,N_4280,N_4868);
or UO_303 (O_303,N_4578,N_4166);
nand UO_304 (O_304,N_4709,N_4782);
xor UO_305 (O_305,N_4902,N_4209);
nand UO_306 (O_306,N_4070,N_4391);
nor UO_307 (O_307,N_4238,N_4714);
nand UO_308 (O_308,N_4517,N_4176);
and UO_309 (O_309,N_4567,N_4251);
and UO_310 (O_310,N_4608,N_4707);
nand UO_311 (O_311,N_4589,N_4219);
and UO_312 (O_312,N_4168,N_4069);
and UO_313 (O_313,N_4340,N_4009);
nor UO_314 (O_314,N_4956,N_4813);
or UO_315 (O_315,N_4689,N_4590);
xnor UO_316 (O_316,N_4917,N_4296);
xor UO_317 (O_317,N_4983,N_4355);
or UO_318 (O_318,N_4527,N_4796);
nor UO_319 (O_319,N_4897,N_4145);
or UO_320 (O_320,N_4771,N_4360);
or UO_321 (O_321,N_4594,N_4698);
nand UO_322 (O_322,N_4918,N_4249);
nor UO_323 (O_323,N_4640,N_4317);
nand UO_324 (O_324,N_4812,N_4175);
nand UO_325 (O_325,N_4021,N_4375);
or UO_326 (O_326,N_4762,N_4135);
nor UO_327 (O_327,N_4480,N_4080);
xnor UO_328 (O_328,N_4414,N_4520);
nand UO_329 (O_329,N_4566,N_4001);
nand UO_330 (O_330,N_4024,N_4438);
and UO_331 (O_331,N_4865,N_4946);
nor UO_332 (O_332,N_4196,N_4180);
nand UO_333 (O_333,N_4235,N_4924);
nand UO_334 (O_334,N_4914,N_4203);
nand UO_335 (O_335,N_4802,N_4395);
or UO_336 (O_336,N_4591,N_4120);
or UO_337 (O_337,N_4803,N_4764);
xnor UO_338 (O_338,N_4318,N_4134);
nor UO_339 (O_339,N_4586,N_4326);
and UO_340 (O_340,N_4078,N_4767);
nand UO_341 (O_341,N_4930,N_4127);
and UO_342 (O_342,N_4903,N_4172);
or UO_343 (O_343,N_4310,N_4601);
xnor UO_344 (O_344,N_4014,N_4680);
or UO_345 (O_345,N_4853,N_4681);
nor UO_346 (O_346,N_4638,N_4809);
and UO_347 (O_347,N_4731,N_4266);
and UO_348 (O_348,N_4104,N_4562);
nand UO_349 (O_349,N_4934,N_4896);
nand UO_350 (O_350,N_4396,N_4273);
and UO_351 (O_351,N_4745,N_4054);
xor UO_352 (O_352,N_4539,N_4106);
xor UO_353 (O_353,N_4199,N_4027);
or UO_354 (O_354,N_4004,N_4182);
nor UO_355 (O_355,N_4348,N_4525);
nand UO_356 (O_356,N_4884,N_4049);
and UO_357 (O_357,N_4169,N_4068);
nor UO_358 (O_358,N_4675,N_4987);
and UO_359 (O_359,N_4928,N_4921);
xor UO_360 (O_360,N_4082,N_4690);
xnor UO_361 (O_361,N_4060,N_4232);
nand UO_362 (O_362,N_4834,N_4363);
nand UO_363 (O_363,N_4345,N_4370);
or UO_364 (O_364,N_4811,N_4708);
xor UO_365 (O_365,N_4156,N_4023);
and UO_366 (O_366,N_4552,N_4306);
or UO_367 (O_367,N_4620,N_4962);
xor UO_368 (O_368,N_4470,N_4333);
and UO_369 (O_369,N_4270,N_4572);
xnor UO_370 (O_370,N_4302,N_4298);
nor UO_371 (O_371,N_4052,N_4672);
and UO_372 (O_372,N_4282,N_4133);
nor UO_373 (O_373,N_4346,N_4195);
nand UO_374 (O_374,N_4831,N_4020);
nor UO_375 (O_375,N_4415,N_4372);
or UO_376 (O_376,N_4434,N_4490);
or UO_377 (O_377,N_4316,N_4483);
nor UO_378 (O_378,N_4178,N_4696);
or UO_379 (O_379,N_4435,N_4990);
xnor UO_380 (O_380,N_4904,N_4079);
and UO_381 (O_381,N_4404,N_4207);
xnor UO_382 (O_382,N_4579,N_4988);
and UO_383 (O_383,N_4876,N_4778);
nand UO_384 (O_384,N_4072,N_4787);
nor UO_385 (O_385,N_4047,N_4874);
xor UO_386 (O_386,N_4657,N_4667);
or UO_387 (O_387,N_4429,N_4844);
xnor UO_388 (O_388,N_4400,N_4750);
and UO_389 (O_389,N_4416,N_4002);
and UO_390 (O_390,N_4048,N_4695);
or UO_391 (O_391,N_4367,N_4982);
and UO_392 (O_392,N_4922,N_4334);
nand UO_393 (O_393,N_4437,N_4064);
or UO_394 (O_394,N_4158,N_4738);
nor UO_395 (O_395,N_4706,N_4448);
nand UO_396 (O_396,N_4693,N_4964);
nand UO_397 (O_397,N_4041,N_4910);
xnor UO_398 (O_398,N_4895,N_4939);
and UO_399 (O_399,N_4243,N_4564);
nand UO_400 (O_400,N_4593,N_4814);
and UO_401 (O_401,N_4379,N_4449);
nand UO_402 (O_402,N_4006,N_4972);
or UO_403 (O_403,N_4581,N_4063);
nand UO_404 (O_404,N_4373,N_4941);
or UO_405 (O_405,N_4262,N_4013);
nand UO_406 (O_406,N_4197,N_4575);
nand UO_407 (O_407,N_4247,N_4493);
xor UO_408 (O_408,N_4384,N_4336);
xor UO_409 (O_409,N_4397,N_4727);
nor UO_410 (O_410,N_4393,N_4821);
and UO_411 (O_411,N_4769,N_4312);
xor UO_412 (O_412,N_4084,N_4507);
or UO_413 (O_413,N_4496,N_4388);
nand UO_414 (O_414,N_4901,N_4911);
nor UO_415 (O_415,N_4845,N_4626);
or UO_416 (O_416,N_4772,N_4676);
or UO_417 (O_417,N_4989,N_4022);
or UO_418 (O_418,N_4445,N_4193);
and UO_419 (O_419,N_4580,N_4319);
or UO_420 (O_420,N_4561,N_4719);
or UO_421 (O_421,N_4651,N_4981);
xnor UO_422 (O_422,N_4549,N_4531);
nor UO_423 (O_423,N_4268,N_4091);
and UO_424 (O_424,N_4855,N_4202);
nor UO_425 (O_425,N_4128,N_4953);
nand UO_426 (O_426,N_4473,N_4229);
or UO_427 (O_427,N_4167,N_4314);
nor UO_428 (O_428,N_4344,N_4290);
nand UO_429 (O_429,N_4655,N_4439);
nor UO_430 (O_430,N_4777,N_4271);
xor UO_431 (O_431,N_4574,N_4737);
nand UO_432 (O_432,N_4450,N_4381);
nor UO_433 (O_433,N_4105,N_4720);
and UO_434 (O_434,N_4847,N_4609);
nor UO_435 (O_435,N_4402,N_4995);
nor UO_436 (O_436,N_4181,N_4584);
or UO_437 (O_437,N_4686,N_4984);
or UO_438 (O_438,N_4929,N_4098);
and UO_439 (O_439,N_4883,N_4087);
and UO_440 (O_440,N_4815,N_4664);
nand UO_441 (O_441,N_4016,N_4261);
or UO_442 (O_442,N_4825,N_4485);
and UO_443 (O_443,N_4543,N_4136);
and UO_444 (O_444,N_4343,N_4465);
and UO_445 (O_445,N_4320,N_4893);
nand UO_446 (O_446,N_4107,N_4131);
nand UO_447 (O_447,N_4997,N_4666);
or UO_448 (O_448,N_4559,N_4615);
and UO_449 (O_449,N_4231,N_4264);
nor UO_450 (O_450,N_4718,N_4830);
nor UO_451 (O_451,N_4489,N_4065);
nor UO_452 (O_452,N_4350,N_4966);
nor UO_453 (O_453,N_4959,N_4452);
xnor UO_454 (O_454,N_4908,N_4636);
nand UO_455 (O_455,N_4970,N_4114);
nand UO_456 (O_456,N_4705,N_4457);
nor UO_457 (O_457,N_4000,N_4278);
nand UO_458 (O_458,N_4673,N_4554);
xnor UO_459 (O_459,N_4660,N_4010);
nor UO_460 (O_460,N_4245,N_4521);
nand UO_461 (O_461,N_4713,N_4969);
nor UO_462 (O_462,N_4045,N_4909);
nor UO_463 (O_463,N_4773,N_4632);
nor UO_464 (O_464,N_4097,N_4228);
and UO_465 (O_465,N_4801,N_4126);
nor UO_466 (O_466,N_4093,N_4836);
xnor UO_467 (O_467,N_4805,N_4509);
nand UO_468 (O_468,N_4958,N_4963);
nand UO_469 (O_469,N_4931,N_4129);
nor UO_470 (O_470,N_4250,N_4974);
nor UO_471 (O_471,N_4880,N_4062);
or UO_472 (O_472,N_4086,N_4411);
xor UO_473 (O_473,N_4141,N_4650);
or UO_474 (O_474,N_4405,N_4744);
xor UO_475 (O_475,N_4170,N_4761);
or UO_476 (O_476,N_4324,N_4968);
nand UO_477 (O_477,N_4463,N_4659);
nand UO_478 (O_478,N_4649,N_4866);
nand UO_479 (O_479,N_4321,N_4206);
and UO_480 (O_480,N_4822,N_4095);
and UO_481 (O_481,N_4818,N_4331);
nand UO_482 (O_482,N_4043,N_4071);
and UO_483 (O_483,N_4479,N_4519);
and UO_484 (O_484,N_4569,N_4898);
or UO_485 (O_485,N_4985,N_4540);
nand UO_486 (O_486,N_4629,N_4791);
nor UO_487 (O_487,N_4759,N_4644);
xnor UO_488 (O_488,N_4542,N_4299);
nor UO_489 (O_489,N_4160,N_4739);
nand UO_490 (O_490,N_4817,N_4938);
and UO_491 (O_491,N_4551,N_4255);
or UO_492 (O_492,N_4768,N_4051);
and UO_493 (O_493,N_4113,N_4269);
xor UO_494 (O_494,N_4682,N_4684);
and UO_495 (O_495,N_4407,N_4571);
nand UO_496 (O_496,N_4339,N_4592);
nand UO_497 (O_497,N_4558,N_4163);
xnor UO_498 (O_498,N_4442,N_4894);
nor UO_499 (O_499,N_4456,N_4287);
or UO_500 (O_500,N_4981,N_4509);
or UO_501 (O_501,N_4861,N_4759);
and UO_502 (O_502,N_4810,N_4296);
nand UO_503 (O_503,N_4793,N_4085);
xnor UO_504 (O_504,N_4744,N_4977);
or UO_505 (O_505,N_4063,N_4722);
xnor UO_506 (O_506,N_4243,N_4344);
nand UO_507 (O_507,N_4638,N_4375);
or UO_508 (O_508,N_4756,N_4186);
or UO_509 (O_509,N_4874,N_4316);
xor UO_510 (O_510,N_4027,N_4896);
xnor UO_511 (O_511,N_4250,N_4756);
or UO_512 (O_512,N_4662,N_4932);
and UO_513 (O_513,N_4840,N_4064);
or UO_514 (O_514,N_4910,N_4616);
or UO_515 (O_515,N_4774,N_4829);
nor UO_516 (O_516,N_4561,N_4930);
and UO_517 (O_517,N_4416,N_4266);
nor UO_518 (O_518,N_4291,N_4893);
and UO_519 (O_519,N_4506,N_4208);
nand UO_520 (O_520,N_4680,N_4771);
and UO_521 (O_521,N_4407,N_4866);
or UO_522 (O_522,N_4384,N_4359);
or UO_523 (O_523,N_4258,N_4991);
and UO_524 (O_524,N_4884,N_4433);
or UO_525 (O_525,N_4267,N_4532);
nor UO_526 (O_526,N_4892,N_4101);
nand UO_527 (O_527,N_4138,N_4144);
or UO_528 (O_528,N_4254,N_4441);
and UO_529 (O_529,N_4311,N_4316);
nor UO_530 (O_530,N_4195,N_4813);
nand UO_531 (O_531,N_4830,N_4277);
or UO_532 (O_532,N_4959,N_4140);
nor UO_533 (O_533,N_4615,N_4312);
or UO_534 (O_534,N_4515,N_4900);
nand UO_535 (O_535,N_4624,N_4217);
and UO_536 (O_536,N_4353,N_4476);
and UO_537 (O_537,N_4366,N_4289);
and UO_538 (O_538,N_4249,N_4648);
or UO_539 (O_539,N_4349,N_4771);
and UO_540 (O_540,N_4942,N_4368);
or UO_541 (O_541,N_4015,N_4786);
or UO_542 (O_542,N_4569,N_4182);
xor UO_543 (O_543,N_4714,N_4177);
nand UO_544 (O_544,N_4959,N_4935);
or UO_545 (O_545,N_4288,N_4004);
xnor UO_546 (O_546,N_4434,N_4211);
or UO_547 (O_547,N_4618,N_4689);
or UO_548 (O_548,N_4125,N_4599);
nand UO_549 (O_549,N_4636,N_4779);
nand UO_550 (O_550,N_4478,N_4374);
nor UO_551 (O_551,N_4459,N_4108);
and UO_552 (O_552,N_4263,N_4296);
nor UO_553 (O_553,N_4460,N_4279);
and UO_554 (O_554,N_4633,N_4990);
nand UO_555 (O_555,N_4664,N_4471);
nor UO_556 (O_556,N_4965,N_4579);
nor UO_557 (O_557,N_4067,N_4615);
and UO_558 (O_558,N_4161,N_4462);
and UO_559 (O_559,N_4532,N_4597);
or UO_560 (O_560,N_4475,N_4094);
or UO_561 (O_561,N_4133,N_4053);
nor UO_562 (O_562,N_4738,N_4947);
xnor UO_563 (O_563,N_4922,N_4902);
nand UO_564 (O_564,N_4424,N_4653);
xor UO_565 (O_565,N_4368,N_4690);
and UO_566 (O_566,N_4544,N_4258);
nor UO_567 (O_567,N_4508,N_4100);
nand UO_568 (O_568,N_4593,N_4709);
nor UO_569 (O_569,N_4209,N_4105);
xor UO_570 (O_570,N_4123,N_4545);
nand UO_571 (O_571,N_4812,N_4727);
xnor UO_572 (O_572,N_4758,N_4494);
xor UO_573 (O_573,N_4566,N_4486);
nand UO_574 (O_574,N_4440,N_4772);
or UO_575 (O_575,N_4728,N_4981);
xor UO_576 (O_576,N_4439,N_4544);
xor UO_577 (O_577,N_4706,N_4447);
nand UO_578 (O_578,N_4039,N_4159);
nor UO_579 (O_579,N_4339,N_4902);
and UO_580 (O_580,N_4135,N_4242);
or UO_581 (O_581,N_4601,N_4881);
and UO_582 (O_582,N_4490,N_4766);
nor UO_583 (O_583,N_4055,N_4367);
or UO_584 (O_584,N_4990,N_4809);
nand UO_585 (O_585,N_4768,N_4978);
and UO_586 (O_586,N_4242,N_4154);
or UO_587 (O_587,N_4516,N_4056);
nand UO_588 (O_588,N_4172,N_4432);
xor UO_589 (O_589,N_4772,N_4312);
nor UO_590 (O_590,N_4266,N_4106);
or UO_591 (O_591,N_4755,N_4936);
nor UO_592 (O_592,N_4301,N_4319);
or UO_593 (O_593,N_4963,N_4657);
nor UO_594 (O_594,N_4568,N_4957);
nor UO_595 (O_595,N_4269,N_4574);
xnor UO_596 (O_596,N_4303,N_4120);
and UO_597 (O_597,N_4612,N_4835);
and UO_598 (O_598,N_4412,N_4380);
nand UO_599 (O_599,N_4191,N_4347);
nand UO_600 (O_600,N_4889,N_4118);
xnor UO_601 (O_601,N_4636,N_4669);
and UO_602 (O_602,N_4486,N_4306);
or UO_603 (O_603,N_4851,N_4751);
or UO_604 (O_604,N_4581,N_4283);
or UO_605 (O_605,N_4295,N_4975);
and UO_606 (O_606,N_4841,N_4611);
xnor UO_607 (O_607,N_4675,N_4965);
nor UO_608 (O_608,N_4122,N_4028);
and UO_609 (O_609,N_4344,N_4426);
nor UO_610 (O_610,N_4196,N_4833);
nor UO_611 (O_611,N_4642,N_4533);
or UO_612 (O_612,N_4555,N_4960);
or UO_613 (O_613,N_4931,N_4825);
nand UO_614 (O_614,N_4581,N_4913);
or UO_615 (O_615,N_4429,N_4369);
nand UO_616 (O_616,N_4435,N_4465);
nand UO_617 (O_617,N_4075,N_4908);
and UO_618 (O_618,N_4843,N_4702);
nand UO_619 (O_619,N_4942,N_4541);
xor UO_620 (O_620,N_4614,N_4241);
nand UO_621 (O_621,N_4276,N_4264);
nand UO_622 (O_622,N_4435,N_4039);
xor UO_623 (O_623,N_4531,N_4134);
and UO_624 (O_624,N_4422,N_4632);
nand UO_625 (O_625,N_4751,N_4657);
and UO_626 (O_626,N_4594,N_4149);
nor UO_627 (O_627,N_4207,N_4547);
or UO_628 (O_628,N_4735,N_4235);
nor UO_629 (O_629,N_4807,N_4118);
xor UO_630 (O_630,N_4720,N_4245);
or UO_631 (O_631,N_4507,N_4101);
xnor UO_632 (O_632,N_4234,N_4905);
nor UO_633 (O_633,N_4410,N_4153);
nor UO_634 (O_634,N_4435,N_4261);
xor UO_635 (O_635,N_4110,N_4105);
or UO_636 (O_636,N_4743,N_4313);
xnor UO_637 (O_637,N_4769,N_4946);
xnor UO_638 (O_638,N_4526,N_4066);
or UO_639 (O_639,N_4085,N_4504);
nand UO_640 (O_640,N_4386,N_4865);
nand UO_641 (O_641,N_4794,N_4502);
and UO_642 (O_642,N_4294,N_4089);
or UO_643 (O_643,N_4044,N_4274);
nor UO_644 (O_644,N_4854,N_4110);
xor UO_645 (O_645,N_4272,N_4082);
xnor UO_646 (O_646,N_4285,N_4690);
xnor UO_647 (O_647,N_4196,N_4822);
xnor UO_648 (O_648,N_4388,N_4961);
nand UO_649 (O_649,N_4462,N_4742);
or UO_650 (O_650,N_4474,N_4085);
nor UO_651 (O_651,N_4001,N_4950);
and UO_652 (O_652,N_4012,N_4067);
or UO_653 (O_653,N_4784,N_4596);
or UO_654 (O_654,N_4025,N_4259);
or UO_655 (O_655,N_4347,N_4484);
or UO_656 (O_656,N_4175,N_4724);
or UO_657 (O_657,N_4106,N_4502);
xnor UO_658 (O_658,N_4513,N_4202);
and UO_659 (O_659,N_4797,N_4308);
nand UO_660 (O_660,N_4867,N_4899);
nand UO_661 (O_661,N_4562,N_4869);
and UO_662 (O_662,N_4449,N_4801);
and UO_663 (O_663,N_4602,N_4652);
nand UO_664 (O_664,N_4066,N_4724);
nor UO_665 (O_665,N_4588,N_4294);
nor UO_666 (O_666,N_4905,N_4367);
nand UO_667 (O_667,N_4751,N_4913);
or UO_668 (O_668,N_4948,N_4296);
or UO_669 (O_669,N_4339,N_4813);
xnor UO_670 (O_670,N_4173,N_4468);
nor UO_671 (O_671,N_4537,N_4901);
nand UO_672 (O_672,N_4863,N_4807);
and UO_673 (O_673,N_4913,N_4562);
and UO_674 (O_674,N_4586,N_4282);
nor UO_675 (O_675,N_4874,N_4716);
nor UO_676 (O_676,N_4227,N_4496);
and UO_677 (O_677,N_4716,N_4695);
xnor UO_678 (O_678,N_4269,N_4850);
nand UO_679 (O_679,N_4394,N_4917);
or UO_680 (O_680,N_4477,N_4027);
or UO_681 (O_681,N_4385,N_4330);
nor UO_682 (O_682,N_4893,N_4925);
xnor UO_683 (O_683,N_4527,N_4386);
xnor UO_684 (O_684,N_4145,N_4455);
nor UO_685 (O_685,N_4245,N_4545);
nor UO_686 (O_686,N_4110,N_4686);
xor UO_687 (O_687,N_4489,N_4581);
or UO_688 (O_688,N_4355,N_4338);
nand UO_689 (O_689,N_4066,N_4365);
nor UO_690 (O_690,N_4149,N_4426);
or UO_691 (O_691,N_4477,N_4965);
and UO_692 (O_692,N_4412,N_4145);
nor UO_693 (O_693,N_4298,N_4003);
or UO_694 (O_694,N_4268,N_4740);
or UO_695 (O_695,N_4144,N_4514);
nor UO_696 (O_696,N_4782,N_4050);
nor UO_697 (O_697,N_4728,N_4421);
xnor UO_698 (O_698,N_4491,N_4944);
nand UO_699 (O_699,N_4276,N_4921);
nor UO_700 (O_700,N_4011,N_4723);
nor UO_701 (O_701,N_4205,N_4499);
or UO_702 (O_702,N_4293,N_4672);
nor UO_703 (O_703,N_4972,N_4063);
xnor UO_704 (O_704,N_4243,N_4247);
nand UO_705 (O_705,N_4129,N_4688);
or UO_706 (O_706,N_4207,N_4202);
nand UO_707 (O_707,N_4393,N_4971);
and UO_708 (O_708,N_4882,N_4881);
nor UO_709 (O_709,N_4129,N_4512);
xor UO_710 (O_710,N_4358,N_4451);
and UO_711 (O_711,N_4117,N_4345);
or UO_712 (O_712,N_4769,N_4060);
nor UO_713 (O_713,N_4952,N_4491);
and UO_714 (O_714,N_4979,N_4008);
nand UO_715 (O_715,N_4632,N_4687);
xnor UO_716 (O_716,N_4072,N_4949);
or UO_717 (O_717,N_4640,N_4901);
xor UO_718 (O_718,N_4212,N_4939);
or UO_719 (O_719,N_4888,N_4690);
or UO_720 (O_720,N_4568,N_4327);
xor UO_721 (O_721,N_4565,N_4282);
or UO_722 (O_722,N_4250,N_4622);
nand UO_723 (O_723,N_4690,N_4584);
nor UO_724 (O_724,N_4023,N_4872);
nor UO_725 (O_725,N_4516,N_4587);
nand UO_726 (O_726,N_4221,N_4329);
nand UO_727 (O_727,N_4497,N_4390);
or UO_728 (O_728,N_4427,N_4106);
nor UO_729 (O_729,N_4743,N_4816);
nand UO_730 (O_730,N_4496,N_4328);
xor UO_731 (O_731,N_4357,N_4407);
xnor UO_732 (O_732,N_4436,N_4047);
nor UO_733 (O_733,N_4981,N_4234);
or UO_734 (O_734,N_4343,N_4943);
xor UO_735 (O_735,N_4099,N_4953);
or UO_736 (O_736,N_4349,N_4356);
nor UO_737 (O_737,N_4906,N_4148);
xor UO_738 (O_738,N_4240,N_4510);
and UO_739 (O_739,N_4584,N_4886);
nand UO_740 (O_740,N_4849,N_4051);
nand UO_741 (O_741,N_4860,N_4505);
or UO_742 (O_742,N_4152,N_4752);
nor UO_743 (O_743,N_4064,N_4876);
and UO_744 (O_744,N_4203,N_4521);
or UO_745 (O_745,N_4779,N_4198);
or UO_746 (O_746,N_4260,N_4118);
nand UO_747 (O_747,N_4373,N_4049);
nor UO_748 (O_748,N_4172,N_4758);
nor UO_749 (O_749,N_4079,N_4322);
nand UO_750 (O_750,N_4405,N_4474);
or UO_751 (O_751,N_4341,N_4125);
xor UO_752 (O_752,N_4157,N_4907);
xor UO_753 (O_753,N_4355,N_4200);
and UO_754 (O_754,N_4016,N_4473);
nand UO_755 (O_755,N_4389,N_4046);
or UO_756 (O_756,N_4555,N_4141);
nor UO_757 (O_757,N_4592,N_4703);
and UO_758 (O_758,N_4355,N_4088);
or UO_759 (O_759,N_4770,N_4653);
nand UO_760 (O_760,N_4864,N_4577);
and UO_761 (O_761,N_4177,N_4715);
xor UO_762 (O_762,N_4104,N_4401);
xor UO_763 (O_763,N_4663,N_4123);
xor UO_764 (O_764,N_4436,N_4384);
xor UO_765 (O_765,N_4903,N_4780);
nor UO_766 (O_766,N_4867,N_4169);
or UO_767 (O_767,N_4221,N_4778);
nor UO_768 (O_768,N_4219,N_4652);
and UO_769 (O_769,N_4204,N_4391);
nor UO_770 (O_770,N_4230,N_4562);
and UO_771 (O_771,N_4276,N_4226);
and UO_772 (O_772,N_4885,N_4611);
nand UO_773 (O_773,N_4280,N_4953);
or UO_774 (O_774,N_4528,N_4778);
or UO_775 (O_775,N_4786,N_4325);
nand UO_776 (O_776,N_4089,N_4480);
and UO_777 (O_777,N_4504,N_4221);
xnor UO_778 (O_778,N_4719,N_4926);
nand UO_779 (O_779,N_4467,N_4837);
nand UO_780 (O_780,N_4813,N_4061);
and UO_781 (O_781,N_4944,N_4283);
xor UO_782 (O_782,N_4314,N_4387);
or UO_783 (O_783,N_4456,N_4794);
xnor UO_784 (O_784,N_4097,N_4111);
or UO_785 (O_785,N_4594,N_4972);
nand UO_786 (O_786,N_4226,N_4774);
and UO_787 (O_787,N_4236,N_4343);
and UO_788 (O_788,N_4366,N_4241);
or UO_789 (O_789,N_4077,N_4614);
and UO_790 (O_790,N_4313,N_4315);
nor UO_791 (O_791,N_4833,N_4708);
nand UO_792 (O_792,N_4291,N_4922);
nand UO_793 (O_793,N_4482,N_4797);
xor UO_794 (O_794,N_4651,N_4082);
xnor UO_795 (O_795,N_4509,N_4420);
nand UO_796 (O_796,N_4979,N_4737);
xor UO_797 (O_797,N_4795,N_4984);
nand UO_798 (O_798,N_4540,N_4629);
or UO_799 (O_799,N_4491,N_4878);
nor UO_800 (O_800,N_4829,N_4669);
or UO_801 (O_801,N_4523,N_4301);
nand UO_802 (O_802,N_4461,N_4377);
and UO_803 (O_803,N_4245,N_4469);
nor UO_804 (O_804,N_4574,N_4556);
and UO_805 (O_805,N_4136,N_4088);
nor UO_806 (O_806,N_4239,N_4796);
or UO_807 (O_807,N_4209,N_4401);
nor UO_808 (O_808,N_4027,N_4928);
nand UO_809 (O_809,N_4882,N_4091);
nor UO_810 (O_810,N_4418,N_4429);
or UO_811 (O_811,N_4688,N_4332);
nor UO_812 (O_812,N_4000,N_4838);
nand UO_813 (O_813,N_4678,N_4211);
and UO_814 (O_814,N_4485,N_4578);
nand UO_815 (O_815,N_4160,N_4773);
or UO_816 (O_816,N_4997,N_4555);
nand UO_817 (O_817,N_4052,N_4746);
nand UO_818 (O_818,N_4150,N_4519);
xor UO_819 (O_819,N_4128,N_4482);
xnor UO_820 (O_820,N_4690,N_4845);
and UO_821 (O_821,N_4970,N_4094);
or UO_822 (O_822,N_4316,N_4985);
xnor UO_823 (O_823,N_4617,N_4958);
nor UO_824 (O_824,N_4332,N_4856);
or UO_825 (O_825,N_4675,N_4806);
xor UO_826 (O_826,N_4954,N_4390);
or UO_827 (O_827,N_4612,N_4053);
nand UO_828 (O_828,N_4244,N_4610);
or UO_829 (O_829,N_4509,N_4987);
nand UO_830 (O_830,N_4940,N_4439);
nor UO_831 (O_831,N_4673,N_4729);
nor UO_832 (O_832,N_4417,N_4477);
nor UO_833 (O_833,N_4717,N_4476);
xor UO_834 (O_834,N_4948,N_4705);
nand UO_835 (O_835,N_4201,N_4851);
or UO_836 (O_836,N_4686,N_4412);
xor UO_837 (O_837,N_4970,N_4112);
xor UO_838 (O_838,N_4855,N_4500);
or UO_839 (O_839,N_4633,N_4185);
or UO_840 (O_840,N_4091,N_4659);
nor UO_841 (O_841,N_4495,N_4622);
nor UO_842 (O_842,N_4177,N_4596);
xnor UO_843 (O_843,N_4368,N_4270);
nand UO_844 (O_844,N_4369,N_4557);
or UO_845 (O_845,N_4896,N_4877);
nor UO_846 (O_846,N_4178,N_4518);
nor UO_847 (O_847,N_4309,N_4384);
and UO_848 (O_848,N_4728,N_4922);
nor UO_849 (O_849,N_4560,N_4484);
and UO_850 (O_850,N_4537,N_4203);
or UO_851 (O_851,N_4866,N_4206);
nand UO_852 (O_852,N_4137,N_4449);
nand UO_853 (O_853,N_4391,N_4626);
or UO_854 (O_854,N_4673,N_4007);
nor UO_855 (O_855,N_4572,N_4294);
and UO_856 (O_856,N_4107,N_4366);
and UO_857 (O_857,N_4175,N_4096);
nand UO_858 (O_858,N_4307,N_4955);
or UO_859 (O_859,N_4360,N_4866);
nand UO_860 (O_860,N_4719,N_4676);
and UO_861 (O_861,N_4089,N_4129);
and UO_862 (O_862,N_4539,N_4713);
nand UO_863 (O_863,N_4157,N_4229);
nor UO_864 (O_864,N_4855,N_4260);
or UO_865 (O_865,N_4471,N_4631);
nand UO_866 (O_866,N_4484,N_4190);
and UO_867 (O_867,N_4837,N_4501);
and UO_868 (O_868,N_4135,N_4834);
and UO_869 (O_869,N_4621,N_4639);
nand UO_870 (O_870,N_4095,N_4774);
xnor UO_871 (O_871,N_4735,N_4952);
or UO_872 (O_872,N_4671,N_4960);
and UO_873 (O_873,N_4468,N_4370);
xnor UO_874 (O_874,N_4868,N_4413);
nor UO_875 (O_875,N_4891,N_4070);
xnor UO_876 (O_876,N_4506,N_4809);
nor UO_877 (O_877,N_4006,N_4795);
and UO_878 (O_878,N_4630,N_4416);
xnor UO_879 (O_879,N_4235,N_4124);
nor UO_880 (O_880,N_4820,N_4531);
nand UO_881 (O_881,N_4995,N_4710);
nor UO_882 (O_882,N_4038,N_4202);
or UO_883 (O_883,N_4651,N_4097);
or UO_884 (O_884,N_4696,N_4800);
nand UO_885 (O_885,N_4209,N_4095);
xor UO_886 (O_886,N_4459,N_4593);
nand UO_887 (O_887,N_4916,N_4778);
nand UO_888 (O_888,N_4244,N_4155);
or UO_889 (O_889,N_4535,N_4289);
and UO_890 (O_890,N_4795,N_4206);
xnor UO_891 (O_891,N_4552,N_4961);
and UO_892 (O_892,N_4623,N_4649);
or UO_893 (O_893,N_4344,N_4588);
nor UO_894 (O_894,N_4968,N_4392);
nor UO_895 (O_895,N_4709,N_4015);
or UO_896 (O_896,N_4411,N_4467);
xnor UO_897 (O_897,N_4600,N_4957);
and UO_898 (O_898,N_4544,N_4967);
nor UO_899 (O_899,N_4710,N_4890);
or UO_900 (O_900,N_4321,N_4765);
and UO_901 (O_901,N_4458,N_4138);
nor UO_902 (O_902,N_4668,N_4159);
or UO_903 (O_903,N_4368,N_4566);
or UO_904 (O_904,N_4713,N_4952);
xor UO_905 (O_905,N_4992,N_4390);
nor UO_906 (O_906,N_4564,N_4960);
nor UO_907 (O_907,N_4761,N_4221);
nand UO_908 (O_908,N_4499,N_4037);
xor UO_909 (O_909,N_4513,N_4536);
nand UO_910 (O_910,N_4010,N_4026);
nand UO_911 (O_911,N_4718,N_4635);
or UO_912 (O_912,N_4559,N_4076);
nand UO_913 (O_913,N_4661,N_4401);
and UO_914 (O_914,N_4783,N_4021);
nand UO_915 (O_915,N_4404,N_4065);
or UO_916 (O_916,N_4488,N_4957);
and UO_917 (O_917,N_4301,N_4637);
or UO_918 (O_918,N_4082,N_4511);
nand UO_919 (O_919,N_4078,N_4737);
and UO_920 (O_920,N_4148,N_4062);
and UO_921 (O_921,N_4989,N_4305);
nor UO_922 (O_922,N_4543,N_4626);
or UO_923 (O_923,N_4768,N_4116);
or UO_924 (O_924,N_4063,N_4040);
and UO_925 (O_925,N_4530,N_4664);
nand UO_926 (O_926,N_4894,N_4627);
and UO_927 (O_927,N_4353,N_4485);
nor UO_928 (O_928,N_4477,N_4422);
or UO_929 (O_929,N_4186,N_4301);
nand UO_930 (O_930,N_4828,N_4653);
nand UO_931 (O_931,N_4848,N_4649);
and UO_932 (O_932,N_4253,N_4295);
and UO_933 (O_933,N_4365,N_4714);
or UO_934 (O_934,N_4219,N_4985);
xor UO_935 (O_935,N_4371,N_4164);
xor UO_936 (O_936,N_4916,N_4518);
nand UO_937 (O_937,N_4696,N_4095);
and UO_938 (O_938,N_4966,N_4516);
nor UO_939 (O_939,N_4367,N_4045);
or UO_940 (O_940,N_4564,N_4709);
nand UO_941 (O_941,N_4028,N_4377);
xor UO_942 (O_942,N_4957,N_4788);
nand UO_943 (O_943,N_4373,N_4491);
xor UO_944 (O_944,N_4421,N_4263);
and UO_945 (O_945,N_4480,N_4609);
nor UO_946 (O_946,N_4823,N_4211);
xor UO_947 (O_947,N_4348,N_4550);
xor UO_948 (O_948,N_4557,N_4639);
or UO_949 (O_949,N_4656,N_4425);
and UO_950 (O_950,N_4140,N_4623);
nand UO_951 (O_951,N_4169,N_4854);
xnor UO_952 (O_952,N_4036,N_4971);
xor UO_953 (O_953,N_4725,N_4110);
nand UO_954 (O_954,N_4625,N_4141);
nand UO_955 (O_955,N_4001,N_4690);
nand UO_956 (O_956,N_4814,N_4220);
nand UO_957 (O_957,N_4544,N_4385);
and UO_958 (O_958,N_4095,N_4826);
and UO_959 (O_959,N_4755,N_4681);
nor UO_960 (O_960,N_4538,N_4113);
xnor UO_961 (O_961,N_4691,N_4409);
xor UO_962 (O_962,N_4684,N_4867);
nor UO_963 (O_963,N_4677,N_4612);
xor UO_964 (O_964,N_4612,N_4315);
xnor UO_965 (O_965,N_4165,N_4879);
nand UO_966 (O_966,N_4625,N_4404);
nand UO_967 (O_967,N_4206,N_4500);
and UO_968 (O_968,N_4865,N_4157);
and UO_969 (O_969,N_4685,N_4150);
and UO_970 (O_970,N_4735,N_4305);
or UO_971 (O_971,N_4447,N_4608);
nand UO_972 (O_972,N_4240,N_4210);
xor UO_973 (O_973,N_4512,N_4137);
xnor UO_974 (O_974,N_4598,N_4982);
nor UO_975 (O_975,N_4781,N_4088);
or UO_976 (O_976,N_4196,N_4656);
or UO_977 (O_977,N_4676,N_4154);
xnor UO_978 (O_978,N_4563,N_4456);
and UO_979 (O_979,N_4326,N_4219);
and UO_980 (O_980,N_4504,N_4721);
xor UO_981 (O_981,N_4601,N_4584);
xnor UO_982 (O_982,N_4883,N_4899);
and UO_983 (O_983,N_4679,N_4986);
xnor UO_984 (O_984,N_4577,N_4874);
xnor UO_985 (O_985,N_4638,N_4468);
and UO_986 (O_986,N_4859,N_4758);
nor UO_987 (O_987,N_4028,N_4318);
nand UO_988 (O_988,N_4108,N_4551);
xnor UO_989 (O_989,N_4550,N_4564);
nor UO_990 (O_990,N_4842,N_4695);
nand UO_991 (O_991,N_4665,N_4577);
and UO_992 (O_992,N_4478,N_4005);
and UO_993 (O_993,N_4601,N_4733);
xnor UO_994 (O_994,N_4089,N_4453);
or UO_995 (O_995,N_4446,N_4996);
or UO_996 (O_996,N_4825,N_4455);
nand UO_997 (O_997,N_4474,N_4813);
or UO_998 (O_998,N_4990,N_4591);
nor UO_999 (O_999,N_4496,N_4275);
endmodule