module basic_2000_20000_2500_4_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_1294,In_907);
or U1 (N_1,In_331,In_1786);
xnor U2 (N_2,In_875,In_1420);
nand U3 (N_3,In_1074,In_58);
xnor U4 (N_4,In_980,In_1261);
or U5 (N_5,In_246,In_874);
nand U6 (N_6,In_1590,In_1660);
nand U7 (N_7,In_98,In_992);
nand U8 (N_8,In_1323,In_1316);
nor U9 (N_9,In_1749,In_193);
nand U10 (N_10,In_1032,In_1206);
nand U11 (N_11,In_1227,In_1827);
nor U12 (N_12,In_1266,In_1679);
or U13 (N_13,In_1961,In_1489);
xor U14 (N_14,In_1665,In_211);
nand U15 (N_15,In_1498,In_1372);
nor U16 (N_16,In_641,In_1578);
and U17 (N_17,In_263,In_1101);
or U18 (N_18,In_779,In_1366);
xor U19 (N_19,In_552,In_1431);
xnor U20 (N_20,In_301,In_1284);
nor U21 (N_21,In_1739,In_1600);
xor U22 (N_22,In_1371,In_274);
nand U23 (N_23,In_987,In_63);
and U24 (N_24,In_476,In_293);
or U25 (N_25,In_1921,In_1088);
nor U26 (N_26,In_738,In_1866);
xnor U27 (N_27,In_966,In_1307);
xnor U28 (N_28,In_818,In_102);
nand U29 (N_29,In_249,In_1621);
xnor U30 (N_30,In_23,In_1963);
or U31 (N_31,In_1280,In_1374);
and U32 (N_32,In_1475,In_1606);
and U33 (N_33,In_1762,In_605);
nand U34 (N_34,In_1017,In_633);
or U35 (N_35,In_783,In_332);
and U36 (N_36,In_1196,In_64);
or U37 (N_37,In_1888,In_1178);
nor U38 (N_38,In_1212,In_453);
and U39 (N_39,In_1730,In_625);
or U40 (N_40,In_1932,In_1253);
nor U41 (N_41,In_1133,In_1235);
nor U42 (N_42,In_1650,In_468);
nand U43 (N_43,In_848,In_1170);
xnor U44 (N_44,In_32,In_1340);
nand U45 (N_45,In_1525,In_1377);
nor U46 (N_46,In_1126,In_640);
xnor U47 (N_47,In_48,In_1423);
nand U48 (N_48,In_1700,In_1260);
and U49 (N_49,In_1887,In_664);
nand U50 (N_50,In_16,In_851);
nand U51 (N_51,In_1444,In_976);
nor U52 (N_52,In_208,In_813);
and U53 (N_53,In_648,In_188);
xor U54 (N_54,In_655,In_921);
xor U55 (N_55,In_799,In_800);
xor U56 (N_56,In_629,In_351);
or U57 (N_57,In_1240,In_380);
nor U58 (N_58,In_1996,In_877);
nand U59 (N_59,In_1817,In_430);
nand U60 (N_60,In_1709,In_1626);
nand U61 (N_61,In_1765,In_755);
xnor U62 (N_62,In_124,In_111);
nand U63 (N_63,In_409,In_1322);
nor U64 (N_64,In_906,In_726);
nor U65 (N_65,In_413,In_1850);
nand U66 (N_66,In_828,In_1465);
nor U67 (N_67,In_137,In_589);
or U68 (N_68,In_775,In_1120);
and U69 (N_69,In_538,In_1347);
or U70 (N_70,In_979,In_1271);
nor U71 (N_71,In_1744,In_1285);
xnor U72 (N_72,In_1649,In_270);
and U73 (N_73,In_682,In_223);
nor U74 (N_74,In_819,In_1622);
xnor U75 (N_75,In_1318,In_962);
or U76 (N_76,In_401,In_1645);
xnor U77 (N_77,In_91,In_765);
xor U78 (N_78,In_1326,In_503);
or U79 (N_79,In_10,In_482);
nor U80 (N_80,In_1695,In_954);
nand U81 (N_81,In_900,In_837);
nand U82 (N_82,In_599,In_403);
xor U83 (N_83,In_789,In_1259);
and U84 (N_84,In_1757,In_1310);
xor U85 (N_85,In_168,In_1335);
nand U86 (N_86,In_559,In_917);
or U87 (N_87,In_1497,In_1092);
nor U88 (N_88,In_592,In_317);
xor U89 (N_89,In_548,In_1012);
nor U90 (N_90,In_1780,In_1009);
nand U91 (N_91,In_1189,In_1130);
nand U92 (N_92,In_1636,In_26);
nor U93 (N_93,In_514,In_347);
xor U94 (N_94,In_1474,In_1816);
nor U95 (N_95,In_1179,In_1478);
or U96 (N_96,In_441,In_835);
xnor U97 (N_97,In_700,In_1927);
xnor U98 (N_98,In_522,In_77);
nand U99 (N_99,In_849,In_1561);
and U100 (N_100,In_702,In_1495);
nor U101 (N_101,In_623,In_880);
or U102 (N_102,In_677,In_1492);
xor U103 (N_103,In_1223,In_1777);
and U104 (N_104,In_881,In_923);
or U105 (N_105,In_8,In_1069);
and U106 (N_106,In_1646,In_1380);
nand U107 (N_107,In_661,In_1736);
nand U108 (N_108,In_1060,In_613);
and U109 (N_109,In_1291,In_89);
xor U110 (N_110,In_1354,In_221);
xor U111 (N_111,In_894,In_1230);
nand U112 (N_112,In_822,In_771);
and U113 (N_113,In_20,In_1019);
and U114 (N_114,In_1885,In_1163);
nor U115 (N_115,In_387,In_255);
or U116 (N_116,In_216,In_951);
nand U117 (N_117,In_425,In_689);
xnor U118 (N_118,In_1997,In_1990);
nand U119 (N_119,In_1985,In_1428);
nor U120 (N_120,In_65,In_373);
and U121 (N_121,In_1583,In_1238);
xor U122 (N_122,In_564,In_1720);
and U123 (N_123,In_694,In_967);
nand U124 (N_124,In_997,In_1175);
nand U125 (N_125,In_395,In_1875);
nor U126 (N_126,In_408,In_486);
or U127 (N_127,In_1246,In_1115);
and U128 (N_128,In_1950,In_1205);
nand U129 (N_129,In_1570,In_247);
xnor U130 (N_130,In_1837,In_398);
or U131 (N_131,In_1878,In_250);
or U132 (N_132,In_109,In_70);
and U133 (N_133,In_1719,In_1615);
or U134 (N_134,In_1422,In_1022);
xor U135 (N_135,In_33,In_596);
or U136 (N_136,In_970,In_687);
nand U137 (N_137,In_119,In_1696);
xnor U138 (N_138,In_1249,In_1233);
and U139 (N_139,In_154,In_899);
and U140 (N_140,In_138,In_575);
nand U141 (N_141,In_1286,In_1991);
and U142 (N_142,In_519,In_1384);
nor U143 (N_143,In_722,In_750);
nor U144 (N_144,In_1864,In_782);
nand U145 (N_145,In_934,In_1586);
nand U146 (N_146,In_686,In_684);
xor U147 (N_147,In_649,In_1232);
and U148 (N_148,In_658,In_806);
nand U149 (N_149,In_815,In_359);
and U150 (N_150,In_535,In_1891);
xnor U151 (N_151,In_161,In_846);
nand U152 (N_152,In_158,In_1694);
nor U153 (N_153,In_1998,In_1360);
nor U154 (N_154,In_298,In_415);
nand U155 (N_155,In_929,In_1097);
xnor U156 (N_156,In_1566,In_745);
or U157 (N_157,In_1013,In_1752);
nand U158 (N_158,In_474,In_1016);
nand U159 (N_159,In_787,In_1499);
nand U160 (N_160,In_136,In_1358);
nand U161 (N_161,In_1794,In_1364);
nand U162 (N_162,In_1569,In_478);
nor U163 (N_163,In_1349,In_713);
and U164 (N_164,In_1607,In_1329);
nand U165 (N_165,In_878,In_1802);
nand U166 (N_166,In_525,In_256);
nand U167 (N_167,In_133,In_1003);
or U168 (N_168,In_1063,In_1493);
and U169 (N_169,In_635,In_43);
nor U170 (N_170,In_791,In_852);
nor U171 (N_171,In_614,In_1244);
nor U172 (N_172,In_467,In_1822);
nor U173 (N_173,In_200,In_1530);
nor U174 (N_174,In_1397,In_1139);
nand U175 (N_175,In_1943,In_1741);
nor U176 (N_176,In_1832,In_1596);
nand U177 (N_177,In_245,In_273);
and U178 (N_178,In_475,In_736);
nor U179 (N_179,In_1215,In_438);
and U180 (N_180,In_1664,In_1764);
nand U181 (N_181,In_1024,In_816);
nand U182 (N_182,In_1432,In_1018);
and U183 (N_183,In_455,In_469);
or U184 (N_184,In_219,In_636);
nand U185 (N_185,In_61,In_854);
nor U186 (N_186,In_587,In_1041);
xnor U187 (N_187,In_499,In_1880);
or U188 (N_188,In_885,In_1871);
xnor U189 (N_189,In_845,In_508);
and U190 (N_190,In_350,In_740);
and U191 (N_191,In_424,In_1838);
and U192 (N_192,In_1166,In_4);
and U193 (N_193,In_318,In_1964);
xnor U194 (N_194,In_1930,In_225);
nand U195 (N_195,In_1523,In_1356);
and U196 (N_196,In_404,In_264);
nand U197 (N_197,In_435,In_1225);
nor U198 (N_198,In_1574,In_214);
and U199 (N_199,In_1750,In_1419);
xor U200 (N_200,In_1064,In_608);
xor U201 (N_201,In_22,In_1840);
and U202 (N_202,In_416,In_1278);
xor U203 (N_203,In_1447,In_1920);
nand U204 (N_204,In_1551,In_14);
and U205 (N_205,In_1121,In_155);
or U206 (N_206,In_1256,In_1197);
nand U207 (N_207,In_1071,In_1629);
xnor U208 (N_208,In_1542,In_1538);
or U209 (N_209,In_1528,In_1234);
and U210 (N_210,In_1929,In_1751);
nand U211 (N_211,In_598,In_427);
xor U212 (N_212,In_458,In_284);
xor U213 (N_213,In_184,In_66);
nor U214 (N_214,In_1782,In_1303);
xor U215 (N_215,In_1090,In_1490);
or U216 (N_216,In_1213,In_1521);
or U217 (N_217,In_309,In_744);
and U218 (N_218,In_733,In_1876);
nor U219 (N_219,In_500,In_1911);
nand U220 (N_220,In_1575,In_606);
xor U221 (N_221,In_910,In_1468);
xnor U222 (N_222,In_774,In_938);
nor U223 (N_223,In_593,In_76);
nor U224 (N_224,In_471,In_166);
nand U225 (N_225,In_114,In_1536);
nand U226 (N_226,In_1339,In_1638);
nor U227 (N_227,In_1870,In_516);
xnor U228 (N_228,In_1216,In_1858);
nand U229 (N_229,In_1915,In_820);
or U230 (N_230,In_1882,In_307);
and U231 (N_231,In_271,In_688);
or U232 (N_232,In_1242,In_39);
and U233 (N_233,In_203,In_377);
nor U234 (N_234,In_1301,In_364);
xor U235 (N_235,In_826,In_639);
nand U236 (N_236,In_382,In_326);
and U237 (N_237,In_1801,In_1763);
or U238 (N_238,In_1772,In_555);
nor U239 (N_239,In_1268,In_1515);
nor U240 (N_240,In_1602,In_487);
nand U241 (N_241,In_1226,In_1524);
nor U242 (N_242,In_37,In_1098);
nor U243 (N_243,In_960,In_266);
xnor U244 (N_244,In_329,In_1006);
xnor U245 (N_245,In_953,In_1691);
nor U246 (N_246,In_620,In_1972);
nor U247 (N_247,In_1288,In_1306);
nor U248 (N_248,In_1556,In_784);
or U249 (N_249,In_652,In_1643);
nor U250 (N_250,In_24,In_805);
nor U251 (N_251,In_95,In_1846);
and U252 (N_252,In_268,In_479);
nand U253 (N_253,In_583,In_62);
or U254 (N_254,In_241,In_780);
and U255 (N_255,In_920,In_753);
or U256 (N_256,In_156,In_28);
nor U257 (N_257,In_619,In_1367);
and U258 (N_258,In_786,In_1657);
xor U259 (N_259,In_563,In_454);
and U260 (N_260,In_1540,In_1174);
or U261 (N_261,In_999,In_141);
and U262 (N_262,In_995,In_916);
xor U263 (N_263,In_1684,In_1237);
nor U264 (N_264,In_1957,In_1129);
xor U265 (N_265,In_855,In_604);
nor U266 (N_266,In_357,In_585);
xnor U267 (N_267,In_84,In_501);
nor U268 (N_268,In_104,In_1066);
nor U269 (N_269,In_1313,In_1409);
or U270 (N_270,In_1193,In_1952);
and U271 (N_271,In_1282,In_927);
or U272 (N_272,In_1106,In_720);
xor U273 (N_273,In_991,In_1290);
nor U274 (N_274,In_776,In_666);
and U275 (N_275,In_1015,In_1031);
or U276 (N_276,In_1481,In_692);
and U277 (N_277,In_346,In_226);
and U278 (N_278,In_1701,In_204);
or U279 (N_279,In_1821,In_343);
or U280 (N_280,In_578,In_1095);
nor U281 (N_281,In_1287,In_1434);
nor U282 (N_282,In_480,In_25);
nand U283 (N_283,In_1597,In_1830);
nand U284 (N_284,In_465,In_1376);
or U285 (N_285,In_1382,In_46);
nor U286 (N_286,In_1818,In_1276);
xor U287 (N_287,In_447,In_1674);
nor U288 (N_288,In_1605,In_561);
or U289 (N_289,In_233,In_647);
nor U290 (N_290,In_565,In_1146);
nand U291 (N_291,In_484,In_134);
nor U292 (N_292,In_729,In_1785);
nand U293 (N_293,In_864,In_1211);
nand U294 (N_294,In_1675,In_1894);
nor U295 (N_295,In_532,In_695);
nand U296 (N_296,In_807,In_312);
and U297 (N_297,In_252,In_665);
nor U298 (N_298,In_234,In_251);
or U299 (N_299,In_1159,In_210);
nor U300 (N_300,In_509,In_344);
nand U301 (N_301,In_1430,In_217);
nor U302 (N_302,In_1753,In_1221);
or U303 (N_303,In_1571,In_1325);
and U304 (N_304,In_383,In_356);
nand U305 (N_305,In_547,In_379);
nand U306 (N_306,In_797,In_1637);
xnor U307 (N_307,In_1317,In_1848);
and U308 (N_308,In_1272,In_1793);
nand U309 (N_309,In_439,In_544);
xnor U310 (N_310,In_182,In_1341);
nand U311 (N_311,In_958,In_618);
nor U312 (N_312,In_1704,In_1375);
and U313 (N_313,In_1729,In_1446);
xor U314 (N_314,In_690,In_1724);
or U315 (N_315,In_902,In_809);
or U316 (N_316,In_1010,In_1172);
or U317 (N_317,In_959,In_393);
nand U318 (N_318,In_1144,In_1761);
xnor U319 (N_319,In_1686,In_1725);
and U320 (N_320,In_785,In_669);
or U321 (N_321,In_1080,In_127);
nor U322 (N_322,In_985,In_1102);
nor U323 (N_323,In_195,In_1297);
nand U324 (N_324,In_1849,In_1845);
nand U325 (N_325,In_1118,In_1595);
xor U326 (N_326,In_616,In_1938);
nor U327 (N_327,In_18,In_798);
or U328 (N_328,In_965,In_1328);
xor U329 (N_329,In_770,In_1164);
xnor U330 (N_330,In_278,In_1081);
nor U331 (N_331,In_178,In_1925);
and U332 (N_332,In_667,In_1342);
and U333 (N_333,In_674,In_1903);
and U334 (N_334,In_1553,In_1760);
xor U335 (N_335,In_705,In_1781);
nor U336 (N_336,In_1184,In_1594);
and U337 (N_337,In_1507,In_1245);
nand U338 (N_338,In_286,In_844);
or U339 (N_339,In_367,In_1379);
nor U340 (N_340,In_1788,In_1418);
xnor U341 (N_341,In_1759,In_248);
nand U342 (N_342,In_378,In_1748);
nand U343 (N_343,In_1699,In_1632);
or U344 (N_344,In_660,In_1416);
nor U345 (N_345,In_400,In_1918);
and U346 (N_346,In_988,In_431);
nand U347 (N_347,In_718,In_473);
or U348 (N_348,In_1554,In_1659);
nor U349 (N_349,In_129,In_507);
xnor U350 (N_350,In_1160,In_1441);
nand U351 (N_351,In_697,In_232);
xnor U352 (N_352,In_524,In_895);
xnor U353 (N_353,In_1350,In_1351);
nand U354 (N_354,In_898,In_536);
or U355 (N_355,In_1200,In_1726);
or U356 (N_356,In_1855,In_1958);
or U357 (N_357,In_601,In_579);
and U358 (N_358,In_1792,In_1154);
or U359 (N_359,In_975,In_983);
or U360 (N_360,In_1337,In_314);
xnor U361 (N_361,In_788,In_1440);
or U362 (N_362,In_1180,In_327);
or U363 (N_363,In_1758,In_1560);
or U364 (N_364,In_1642,In_1204);
or U365 (N_365,In_135,In_108);
and U366 (N_366,In_229,In_1136);
xnor U367 (N_367,In_1731,In_1799);
or U368 (N_368,In_1293,In_1773);
xor U369 (N_369,In_1406,In_434);
or U370 (N_370,In_1262,In_1369);
nand U371 (N_371,In_531,In_1161);
and U372 (N_372,In_1940,In_1345);
or U373 (N_373,In_1517,In_769);
nand U374 (N_374,In_998,In_1820);
xor U375 (N_375,In_1986,In_1045);
and U376 (N_376,In_703,In_1808);
nor U377 (N_377,In_1267,In_1941);
and U378 (N_378,In_550,In_101);
xor U379 (N_379,In_663,In_481);
and U380 (N_380,In_390,In_483);
or U381 (N_381,In_1783,In_489);
and U382 (N_382,In_884,In_172);
or U383 (N_383,In_1833,In_632);
or U384 (N_384,In_372,In_1960);
xor U385 (N_385,In_990,In_723);
and U386 (N_386,In_915,In_1733);
or U387 (N_387,In_982,In_1128);
and U388 (N_388,In_176,In_1085);
xor U389 (N_389,In_754,In_57);
xor U390 (N_390,In_748,In_812);
nor U391 (N_391,In_238,In_1913);
and U392 (N_392,In_44,In_1754);
and U393 (N_393,In_594,In_1047);
or U394 (N_394,In_1001,In_192);
nor U395 (N_395,In_1623,In_1086);
and U396 (N_396,In_305,In_423);
and U397 (N_397,In_1207,In_1791);
nand U398 (N_398,In_85,In_186);
or U399 (N_399,In_612,In_1900);
nor U400 (N_400,In_376,In_1896);
nand U401 (N_401,In_180,In_1076);
nor U402 (N_402,In_206,In_181);
and U403 (N_403,In_1770,In_1302);
xnor U404 (N_404,In_1969,In_1411);
and U405 (N_405,In_257,In_803);
nand U406 (N_406,In_103,In_1362);
and U407 (N_407,In_227,In_1873);
nor U408 (N_408,In_603,In_1250);
and U409 (N_409,In_1452,In_1743);
or U410 (N_410,In_228,In_1933);
and U411 (N_411,In_628,In_950);
xor U412 (N_412,In_126,In_558);
nor U413 (N_413,In_654,In_529);
nand U414 (N_414,In_1651,In_1722);
and U415 (N_415,In_928,In_1689);
or U416 (N_416,In_1334,In_1644);
and U417 (N_417,In_1040,In_1055);
nand U418 (N_418,In_831,In_1740);
nand U419 (N_419,In_808,In_100);
nand U420 (N_420,In_1368,In_607);
or U421 (N_421,In_869,In_656);
or U422 (N_422,In_1068,In_1218);
xnor U423 (N_423,In_1039,In_1321);
nand U424 (N_424,In_146,In_1070);
nor U425 (N_425,In_1835,In_1779);
nor U426 (N_426,In_678,In_173);
or U427 (N_427,In_1198,In_1811);
xor U428 (N_428,In_1862,In_1916);
and U429 (N_429,In_450,In_1989);
and U430 (N_430,In_597,In_87);
nor U431 (N_431,In_128,In_511);
and U432 (N_432,In_1581,In_1968);
nand U433 (N_433,In_1292,In_1756);
nand U434 (N_434,In_42,In_1265);
nand U435 (N_435,In_724,In_1470);
or U436 (N_436,In_1949,In_1077);
nand U437 (N_437,In_1094,In_940);
and U438 (N_438,In_93,In_1455);
and U439 (N_439,In_92,In_1111);
nand U440 (N_440,In_1673,In_876);
or U441 (N_441,In_231,In_1955);
nor U442 (N_442,In_913,In_1124);
and U443 (N_443,In_361,In_420);
or U444 (N_444,In_13,In_236);
nand U445 (N_445,In_1580,In_767);
and U446 (N_446,In_762,In_737);
xnor U447 (N_447,In_1361,In_1812);
nand U448 (N_448,In_1370,In_502);
nand U449 (N_449,In_650,In_417);
or U450 (N_450,In_1014,In_242);
xnor U451 (N_451,In_1710,In_222);
nor U452 (N_452,In_1588,In_1591);
xnor U453 (N_453,In_1683,In_1826);
or U454 (N_454,In_325,In_1735);
nand U455 (N_455,In_1831,In_841);
nor U456 (N_456,In_570,In_569);
nor U457 (N_457,In_1251,In_1252);
xnor U458 (N_458,In_1403,In_568);
nor U459 (N_459,In_586,In_793);
nor U460 (N_460,In_717,In_1935);
nor U461 (N_461,In_763,In_488);
xnor U462 (N_462,In_340,In_1201);
nand U463 (N_463,In_595,In_81);
xnor U464 (N_464,In_294,In_237);
xor U465 (N_465,In_1073,In_761);
and U466 (N_466,In_1775,In_964);
nand U467 (N_467,In_1718,In_691);
or U468 (N_468,In_1987,In_1119);
xnor U469 (N_469,In_456,In_1836);
xnor U470 (N_470,In_1687,In_1712);
and U471 (N_471,In_1867,In_1608);
xor U472 (N_472,In_349,In_396);
and U473 (N_473,In_646,In_285);
nor U474 (N_474,In_671,In_1723);
or U475 (N_475,In_1413,In_125);
and U476 (N_476,In_442,In_1004);
and U477 (N_477,In_40,In_337);
and U478 (N_478,In_392,In_348);
and U479 (N_479,In_177,In_291);
xor U480 (N_480,In_735,In_839);
nor U481 (N_481,In_981,In_1967);
nand U482 (N_482,In_572,In_457);
and U483 (N_483,In_253,In_1283);
and U484 (N_484,In_159,In_421);
xor U485 (N_485,In_152,In_1059);
xor U486 (N_486,In_922,In_130);
xnor U487 (N_487,In_97,In_429);
xnor U488 (N_488,In_528,In_283);
xnor U489 (N_489,In_715,In_1378);
and U490 (N_490,In_1884,In_261);
xnor U491 (N_491,In_1148,In_773);
xor U492 (N_492,In_1662,In_9);
and U493 (N_493,In_1036,In_1614);
xor U494 (N_494,In_1589,In_918);
nor U495 (N_495,In_375,In_428);
nor U496 (N_496,In_86,In_1666);
nand U497 (N_497,In_1108,In_644);
or U498 (N_498,In_1093,In_1053);
nor U499 (N_499,In_1389,In_67);
nand U500 (N_500,In_521,In_470);
nand U501 (N_501,In_1473,In_930);
xnor U502 (N_502,In_602,In_626);
nand U503 (N_503,In_662,In_443);
xnor U504 (N_504,In_123,In_1550);
xnor U505 (N_505,In_302,In_562);
xnor U506 (N_506,In_1346,In_1533);
or U507 (N_507,In_1769,In_451);
or U508 (N_508,In_1125,In_355);
nand U509 (N_509,In_1522,In_352);
or U510 (N_510,In_165,In_573);
and U511 (N_511,In_861,In_198);
and U512 (N_512,In_292,In_1937);
xor U513 (N_513,In_1320,In_1096);
and U514 (N_514,In_1167,In_1860);
nand U515 (N_515,In_0,In_941);
or U516 (N_516,In_1585,In_795);
and U517 (N_517,In_259,In_267);
xnor U518 (N_518,In_1815,In_197);
xor U519 (N_519,In_1995,In_1304);
nor U520 (N_520,In_1789,In_1050);
nand U521 (N_521,In_1156,In_194);
nor U522 (N_522,In_1083,In_1439);
or U523 (N_523,In_106,In_1652);
and U524 (N_524,In_1191,In_1412);
nand U525 (N_525,In_1388,In_1856);
xnor U526 (N_526,In_1582,In_533);
nor U527 (N_527,In_1451,In_850);
and U528 (N_528,In_1796,In_1844);
nor U529 (N_529,In_461,In_118);
and U530 (N_530,In_746,In_727);
nand U531 (N_531,In_362,In_1670);
nor U532 (N_532,In_1627,In_1424);
xor U533 (N_533,In_49,In_1567);
nor U534 (N_534,In_407,In_1435);
or U535 (N_535,In_183,In_1678);
nor U536 (N_536,In_804,In_433);
xnor U537 (N_537,In_1464,In_1979);
xnor U538 (N_538,In_1661,In_1910);
and U539 (N_539,In_1897,In_1934);
nand U540 (N_540,In_1618,In_1518);
xnor U541 (N_541,In_1526,In_1755);
xor U542 (N_542,In_1421,In_269);
and U543 (N_543,In_1186,In_973);
nand U544 (N_544,In_840,In_244);
or U545 (N_545,In_446,In_1892);
nand U546 (N_546,In_749,In_1203);
or U547 (N_547,In_75,In_1877);
nor U548 (N_548,In_139,In_1800);
and U549 (N_549,In_1577,In_437);
and U550 (N_550,In_764,In_1711);
and U551 (N_551,In_1559,In_1273);
and U552 (N_552,In_696,In_925);
or U553 (N_553,In_504,In_1488);
nor U554 (N_554,In_1224,In_1270);
xor U555 (N_555,In_1633,In_1568);
xnor U556 (N_556,In_890,In_693);
nand U557 (N_557,In_313,In_1208);
or U558 (N_558,In_1620,In_1889);
or U559 (N_559,In_1264,In_766);
or U560 (N_560,In_310,In_1084);
nor U561 (N_561,In_1572,In_1062);
or U562 (N_562,In_1183,In_584);
xor U563 (N_563,In_833,In_834);
nand U564 (N_564,In_1564,In_472);
and U565 (N_565,In_1655,In_460);
nor U566 (N_566,In_1131,In_1854);
xnor U567 (N_567,In_747,In_218);
nor U568 (N_568,In_1007,In_1734);
and U569 (N_569,In_59,In_1828);
nor U570 (N_570,In_74,In_1698);
xor U571 (N_571,In_865,In_1680);
nand U572 (N_572,In_69,In_147);
nor U573 (N_573,In_105,In_385);
nand U574 (N_574,In_1365,In_1945);
nand U575 (N_575,In_1625,In_896);
nor U576 (N_576,In_1391,In_1486);
nor U577 (N_577,In_289,In_73);
xor U578 (N_578,In_631,In_1399);
xor U579 (N_579,In_540,In_339);
nor U580 (N_580,In_1467,In_512);
or U581 (N_581,In_1162,In_1281);
nand U582 (N_582,In_741,In_1947);
and U583 (N_583,In_1634,In_1026);
and U584 (N_584,In_704,In_919);
and U585 (N_585,In_1681,In_1052);
nand U586 (N_586,In_235,In_1951);
and U587 (N_587,In_926,In_1914);
and U588 (N_588,In_1177,In_153);
xor U589 (N_589,In_1513,In_5);
and U590 (N_590,In_1336,In_1813);
or U591 (N_591,In_381,In_1023);
and U592 (N_592,In_162,In_1476);
nand U593 (N_593,In_1803,In_1936);
xor U594 (N_594,In_871,In_1510);
nand U595 (N_595,In_1445,In_113);
nand U596 (N_596,In_622,In_1274);
and U597 (N_597,In_937,In_1693);
nand U598 (N_598,In_94,In_174);
or U599 (N_599,In_1219,In_449);
and U600 (N_600,In_12,In_879);
nand U601 (N_601,In_388,In_1715);
nor U602 (N_602,In_832,In_904);
xor U603 (N_603,In_335,In_11);
or U604 (N_604,In_353,In_1458);
nor U605 (N_605,In_1565,In_1959);
or U606 (N_606,In_1314,In_330);
nor U607 (N_607,In_1299,In_1134);
nand U608 (N_608,In_1484,In_1705);
or U609 (N_609,In_21,In_1976);
or U610 (N_610,In_627,In_1954);
and U611 (N_611,In_1117,In_88);
xor U612 (N_612,In_402,In_1295);
nand U613 (N_613,In_1429,In_1737);
nor U614 (N_614,In_319,In_79);
nor U615 (N_615,In_977,In_143);
or U616 (N_616,In_448,In_1112);
and U617 (N_617,In_1671,In_254);
or U618 (N_618,In_265,In_334);
and U619 (N_619,In_1002,In_240);
nor U620 (N_620,In_1992,In_949);
nor U621 (N_621,In_1459,In_887);
xor U622 (N_622,In_426,In_1381);
nor U623 (N_623,In_751,In_1535);
nand U624 (N_624,In_1438,In_545);
nand U625 (N_625,In_870,In_1054);
or U626 (N_626,In_1509,In_897);
and U627 (N_627,In_419,In_1942);
and U628 (N_628,In_824,In_1214);
xnor U629 (N_629,In_1044,In_1400);
xnor U630 (N_630,In_78,In_17);
nand U631 (N_631,In_1145,In_701);
nand U632 (N_632,In_955,In_706);
nand U633 (N_633,In_498,In_1469);
xnor U634 (N_634,In_1814,In_802);
nor U635 (N_635,In_1309,In_31);
and U636 (N_636,In_187,In_1974);
and U637 (N_637,In_1137,In_659);
xnor U638 (N_638,In_827,In_50);
nor U639 (N_639,In_1008,In_277);
or U640 (N_640,In_1617,In_946);
nor U641 (N_641,In_760,In_132);
and U642 (N_642,In_157,In_260);
nor U643 (N_643,In_1669,In_574);
nand U644 (N_644,In_1312,In_1548);
nor U645 (N_645,In_1898,In_903);
nor U646 (N_646,In_675,In_1573);
xnor U647 (N_647,In_1386,In_1437);
and U648 (N_648,In_175,In_1289);
xnor U649 (N_649,In_888,In_445);
nand U650 (N_650,In_969,In_1078);
nand U651 (N_651,In_944,In_956);
or U652 (N_652,In_709,In_948);
and U653 (N_653,In_1395,In_1427);
xnor U654 (N_654,In_1917,In_1601);
xor U655 (N_655,In_1984,In_1795);
xnor U656 (N_656,In_145,In_207);
xor U657 (N_657,In_1426,In_7);
xor U658 (N_658,In_1338,In_149);
or U659 (N_659,In_1784,In_170);
nand U660 (N_660,In_933,In_931);
and U661 (N_661,In_1819,In_1480);
and U662 (N_662,In_645,In_1113);
nand U663 (N_663,In_1776,In_942);
nor U664 (N_664,In_1544,In_642);
nor U665 (N_665,In_1869,In_1520);
and U666 (N_666,In_363,In_1220);
nand U667 (N_667,In_1639,In_873);
nor U668 (N_668,In_1043,In_1408);
xnor U669 (N_669,In_374,In_1534);
nor U670 (N_670,In_1727,In_1853);
and U671 (N_671,In_1449,In_144);
and U672 (N_672,In_1332,In_1682);
or U673 (N_673,In_637,In_1169);
and U674 (N_674,In_463,In_1188);
nand U675 (N_675,In_1308,In_338);
xor U676 (N_676,In_1020,In_1980);
or U677 (N_677,In_35,In_117);
or U678 (N_678,In_1872,In_676);
xor U679 (N_679,In_202,In_1448);
nand U680 (N_680,In_296,In_201);
xnor U681 (N_681,In_526,In_1414);
xor U682 (N_682,In_1058,In_1410);
xor U683 (N_683,In_557,In_757);
or U684 (N_684,In_384,In_1082);
xnor U685 (N_685,In_576,In_1692);
nand U686 (N_686,In_397,In_1353);
nand U687 (N_687,In_1067,In_936);
nor U688 (N_688,In_1311,In_1944);
or U689 (N_689,In_112,In_772);
nand U690 (N_690,In_342,In_120);
nor U691 (N_691,In_778,In_892);
xnor U692 (N_692,In_1257,In_1158);
nor U693 (N_693,In_1516,In_1697);
nor U694 (N_694,In_205,In_1787);
or U695 (N_695,In_1552,In_406);
and U696 (N_696,In_710,In_1658);
nor U697 (N_697,In_306,In_634);
and U698 (N_698,In_336,In_1810);
nor U699 (N_699,In_389,In_615);
xnor U700 (N_700,In_1150,In_1025);
and U701 (N_701,In_685,In_1883);
and U702 (N_702,In_169,In_345);
xnor U703 (N_703,In_282,In_1804);
nand U704 (N_704,In_1141,In_276);
nand U705 (N_705,In_1502,In_792);
xnor U706 (N_706,In_1239,In_1168);
xor U707 (N_707,In_1072,In_752);
or U708 (N_708,In_82,In_1797);
nor U709 (N_709,In_768,In_1155);
or U710 (N_710,In_1593,In_1127);
or U711 (N_711,In_1457,In_1182);
xor U712 (N_712,In_1210,In_370);
nand U713 (N_713,In_279,In_150);
xnor U714 (N_714,In_1988,In_1579);
xnor U715 (N_715,In_107,In_1685);
and U716 (N_716,In_1373,In_817);
or U717 (N_717,In_1359,In_847);
nand U718 (N_718,In_1647,In_707);
xor U719 (N_719,In_554,In_1541);
xor U720 (N_720,In_1713,In_1305);
or U721 (N_721,In_1654,In_1558);
nand U722 (N_722,In_1901,In_258);
nand U723 (N_723,In_1089,In_886);
nand U724 (N_724,In_600,In_611);
nand U725 (N_725,In_304,In_1456);
and U726 (N_726,In_1908,In_679);
nor U727 (N_727,In_1048,In_1405);
xnor U728 (N_728,In_734,In_272);
or U729 (N_729,In_1463,In_1923);
nor U730 (N_730,In_866,In_3);
xnor U731 (N_731,In_1185,In_411);
xnor U732 (N_732,In_1363,In_324);
nor U733 (N_733,In_1742,In_1890);
or U734 (N_734,In_1505,In_1254);
or U735 (N_735,In_1433,In_1919);
or U736 (N_736,In_1970,In_730);
xnor U737 (N_737,In_189,In_220);
or U738 (N_738,In_1909,In_1975);
or U739 (N_739,In_1506,In_588);
xor U740 (N_740,In_1417,In_1983);
and U741 (N_741,In_51,In_1151);
or U742 (N_742,In_287,In_1543);
xnor U743 (N_743,In_1904,In_321);
nand U744 (N_744,In_1255,In_151);
and U745 (N_745,In_1839,In_1928);
and U746 (N_746,In_963,In_1404);
or U747 (N_747,In_1592,In_1157);
xnor U748 (N_748,In_1631,In_1333);
nand U749 (N_749,In_1863,In_1051);
and U750 (N_750,In_630,In_539);
nand U751 (N_751,In_790,In_1107);
and U752 (N_752,In_1135,In_191);
and U753 (N_753,In_829,In_1030);
or U754 (N_754,In_905,In_1981);
or U755 (N_755,In_368,In_96);
and U756 (N_756,In_45,In_1676);
xnor U757 (N_757,In_683,In_1181);
xnor U758 (N_758,In_1217,In_224);
or U759 (N_759,In_323,In_399);
or U760 (N_760,In_1190,In_1202);
or U761 (N_761,In_68,In_1688);
xnor U762 (N_762,In_1028,In_1407);
nor U763 (N_763,In_164,In_1153);
or U764 (N_764,In_856,In_994);
or U765 (N_765,In_1962,In_315);
xnor U766 (N_766,In_1708,In_1330);
xor U767 (N_767,In_1613,In_167);
nor U768 (N_768,In_670,In_891);
nor U769 (N_769,In_496,In_796);
xor U770 (N_770,In_1993,In_947);
nor U771 (N_771,In_580,In_1099);
and U772 (N_772,In_41,In_590);
or U773 (N_773,In_386,In_551);
and U774 (N_774,In_621,In_867);
or U775 (N_775,In_262,In_1471);
and U776 (N_776,In_1612,In_1466);
and U777 (N_777,In_978,In_699);
nand U778 (N_778,In_163,In_1355);
xor U779 (N_779,In_440,In_1398);
or U780 (N_780,In_743,In_1263);
and U781 (N_781,In_1462,In_843);
xor U782 (N_782,In_1707,In_914);
and U783 (N_783,In_1401,In_1531);
nand U784 (N_784,In_369,In_582);
xnor U785 (N_785,In_1357,In_160);
and U786 (N_786,In_1668,In_1717);
xor U787 (N_787,In_883,In_1532);
nor U788 (N_788,In_290,In_945);
nand U789 (N_789,In_464,In_1243);
nor U790 (N_790,In_90,In_1442);
or U791 (N_791,In_1176,In_1640);
nor U792 (N_792,In_1545,In_1971);
or U793 (N_793,In_725,In_1079);
xnor U794 (N_794,In_901,In_581);
nand U795 (N_795,In_638,In_1491);
and U796 (N_796,In_872,In_55);
and U797 (N_797,In_280,In_1352);
nand U798 (N_798,In_1624,In_996);
xor U799 (N_799,In_2,In_794);
nand U800 (N_800,In_541,In_1109);
xnor U801 (N_801,In_311,In_1847);
or U802 (N_802,In_1843,In_1461);
nor U803 (N_803,In_1663,In_1809);
nor U804 (N_804,In_1149,In_560);
and U805 (N_805,In_657,In_957);
and U806 (N_806,In_1194,In_1033);
xnor U807 (N_807,In_1774,In_1690);
xnor U808 (N_808,In_1824,In_1123);
xor U809 (N_809,In_989,In_288);
xnor U810 (N_810,In_148,In_80);
or U811 (N_811,In_1324,In_1104);
nor U812 (N_812,In_1460,In_801);
and U813 (N_813,In_412,In_1881);
nand U814 (N_814,In_209,In_366);
nand U815 (N_815,In_1344,In_1977);
or U816 (N_816,In_1778,In_986);
and U817 (N_817,In_320,In_1173);
and U818 (N_818,In_1738,In_1142);
or U819 (N_819,In_1834,In_492);
nor U820 (N_820,In_1825,In_485);
nor U821 (N_821,In_1746,In_1056);
and U822 (N_822,In_728,In_299);
nor U823 (N_823,In_1049,In_830);
nand U824 (N_824,In_1842,In_1648);
nor U825 (N_825,In_935,In_230);
or U826 (N_826,In_1767,In_1672);
nor U827 (N_827,In_1728,In_295);
and U828 (N_828,In_961,In_459);
nor U829 (N_829,In_527,In_1503);
nor U830 (N_830,In_1511,In_523);
xnor U831 (N_831,In_1483,In_56);
xnor U832 (N_832,In_239,In_781);
nor U833 (N_833,In_1087,In_1500);
and U834 (N_834,In_1630,In_836);
or U835 (N_835,In_1514,In_515);
and U836 (N_836,In_1857,In_6);
xor U837 (N_837,In_1105,In_1529);
nor U838 (N_838,In_422,In_971);
nor U839 (N_839,In_882,In_1653);
nor U840 (N_840,In_506,In_1005);
and U841 (N_841,In_1771,In_1436);
or U842 (N_842,In_1851,In_1229);
and U843 (N_843,In_436,In_1065);
nand U844 (N_844,In_1946,In_1383);
or U845 (N_845,In_1319,In_825);
nand U846 (N_846,In_1861,In_122);
nand U847 (N_847,In_1209,In_517);
and U848 (N_848,In_571,In_1035);
and U849 (N_849,In_549,In_811);
or U850 (N_850,In_60,In_1393);
nor U851 (N_851,In_1899,In_212);
nor U852 (N_852,In_477,In_1766);
or U853 (N_853,In_974,In_322);
and U854 (N_854,In_140,In_889);
and U855 (N_855,In_1171,In_566);
nand U856 (N_856,In_30,In_1994);
xor U857 (N_857,In_1598,In_1485);
or U858 (N_858,In_1103,In_1027);
nand U859 (N_859,In_1034,In_1635);
and U860 (N_860,In_1279,In_673);
nand U861 (N_861,In_1790,In_542);
xnor U862 (N_862,In_1716,In_1343);
nand U863 (N_863,In_303,In_952);
nor U864 (N_864,In_1527,In_71);
nand U865 (N_865,In_853,In_495);
and U866 (N_866,In_1392,In_1110);
or U867 (N_867,In_1895,In_414);
nand U868 (N_868,In_1300,In_513);
nand U869 (N_869,In_1275,In_1114);
nor U870 (N_870,In_1396,In_719);
nand U871 (N_871,In_1496,In_643);
nand U872 (N_872,In_553,In_1798);
and U873 (N_873,In_171,In_1494);
and U874 (N_874,In_1037,In_651);
xor U875 (N_875,In_1745,In_567);
or U876 (N_876,In_52,In_142);
nand U877 (N_877,In_1982,In_281);
nand U878 (N_878,In_297,In_29);
xnor U879 (N_879,In_712,In_1805);
and U880 (N_880,In_1893,In_328);
xor U881 (N_881,In_196,In_698);
nand U882 (N_882,In_756,In_862);
or U883 (N_883,In_1721,In_1487);
nand U884 (N_884,In_47,In_1390);
or U885 (N_885,In_1236,In_518);
or U886 (N_886,In_1823,In_810);
and U887 (N_887,In_777,In_1584);
nand U888 (N_888,In_1100,In_1902);
and U889 (N_889,In_1482,In_1331);
nor U890 (N_890,In_1348,In_534);
xor U891 (N_891,In_742,In_681);
or U892 (N_892,In_617,In_863);
nand U893 (N_893,In_1702,In_1926);
and U894 (N_894,In_939,In_1852);
and U895 (N_895,In_714,In_1057);
and U896 (N_896,In_15,In_1562);
nor U897 (N_897,In_1187,In_1879);
xnor U898 (N_898,In_371,In_185);
and U899 (N_899,In_1222,In_1905);
nor U900 (N_900,In_653,In_1922);
or U901 (N_901,In_530,In_1479);
nand U902 (N_902,In_731,In_1924);
nand U903 (N_903,In_1258,In_1000);
or U904 (N_904,In_1703,In_1610);
nand U905 (N_905,In_1611,In_1387);
xor U906 (N_906,In_1931,In_391);
xor U907 (N_907,In_624,In_721);
and U908 (N_908,In_972,In_1277);
and U909 (N_909,In_275,In_1656);
and U910 (N_910,In_1841,In_1886);
and U911 (N_911,In_1199,In_1956);
and U912 (N_912,In_1609,In_1038);
xnor U913 (N_913,In_546,In_1091);
or U914 (N_914,In_1508,In_466);
and U915 (N_915,In_711,In_308);
or U916 (N_916,In_1604,In_497);
or U917 (N_917,In_1966,In_444);
or U918 (N_918,In_1402,In_1512);
xor U919 (N_919,In_1599,In_868);
and U920 (N_920,In_556,In_1999);
or U921 (N_921,In_1138,In_53);
and U922 (N_922,In_1677,In_859);
nor U923 (N_923,In_432,In_823);
xor U924 (N_924,In_1859,In_452);
nor U925 (N_925,In_1046,In_38);
and U926 (N_926,In_493,In_1667);
nor U927 (N_927,In_1587,In_893);
nor U928 (N_928,In_716,In_1563);
and U929 (N_929,In_908,In_1327);
xor U930 (N_930,In_909,In_1143);
xnor U931 (N_931,In_1912,In_1537);
or U932 (N_932,In_1385,In_1865);
xnor U933 (N_933,In_1147,In_1122);
xor U934 (N_934,In_1116,In_213);
or U935 (N_935,In_54,In_1603);
and U936 (N_936,In_1075,In_1714);
nand U937 (N_937,In_732,In_1747);
nand U938 (N_938,In_672,In_609);
xor U939 (N_939,In_520,In_1501);
nor U940 (N_940,In_842,In_510);
or U941 (N_941,In_708,In_34);
and U942 (N_942,In_758,In_912);
and U943 (N_943,In_543,In_1906);
xnor U944 (N_944,In_1247,In_1425);
xnor U945 (N_945,In_1152,In_1195);
xor U946 (N_946,In_1042,In_1868);
nor U947 (N_947,In_739,In_668);
or U948 (N_948,In_418,In_1978);
nand U949 (N_949,In_72,In_1539);
or U950 (N_950,In_360,In_1298);
or U951 (N_951,In_759,In_1472);
nor U952 (N_952,In_1,In_1965);
xor U953 (N_953,In_131,In_341);
nand U954 (N_954,In_1450,In_858);
and U955 (N_955,In_968,In_333);
xnor U956 (N_956,In_110,In_115);
nor U957 (N_957,In_1829,In_1248);
and U958 (N_958,In_1807,In_860);
or U959 (N_959,In_116,In_680);
or U960 (N_960,In_1555,In_358);
xor U961 (N_961,In_1454,In_1619);
xnor U962 (N_962,In_610,In_490);
and U963 (N_963,In_410,In_1394);
or U964 (N_964,In_1029,In_1021);
xnor U965 (N_965,In_1948,In_1231);
and U966 (N_966,In_1504,In_354);
and U967 (N_967,In_190,In_316);
nand U968 (N_968,In_932,In_300);
and U969 (N_969,In_591,In_984);
and U970 (N_970,In_1547,In_1557);
and U971 (N_971,In_857,In_1241);
nand U972 (N_972,In_494,In_1140);
xnor U973 (N_973,In_943,In_243);
and U974 (N_974,In_814,In_365);
xnor U975 (N_975,In_215,In_1296);
nor U976 (N_976,In_1706,In_1061);
nor U977 (N_977,In_1907,In_1228);
nor U978 (N_978,In_1415,In_1192);
xnor U979 (N_979,In_1315,In_1616);
nand U980 (N_980,In_27,In_1269);
nand U981 (N_981,In_838,In_1546);
nand U982 (N_982,In_821,In_1939);
and U983 (N_983,In_1519,In_179);
or U984 (N_984,In_1477,In_505);
nor U985 (N_985,In_911,In_394);
nor U986 (N_986,In_924,In_1443);
nand U987 (N_987,In_36,In_1732);
and U988 (N_988,In_121,In_83);
xor U989 (N_989,In_577,In_1973);
nor U990 (N_990,In_1132,In_1768);
or U991 (N_991,In_993,In_1453);
nand U992 (N_992,In_99,In_1806);
or U993 (N_993,In_405,In_1011);
nand U994 (N_994,In_1628,In_19);
nor U995 (N_995,In_491,In_1953);
xnor U996 (N_996,In_1165,In_1576);
xor U997 (N_997,In_1641,In_462);
xnor U998 (N_998,In_537,In_1549);
nand U999 (N_999,In_199,In_1874);
xnor U1000 (N_1000,In_1427,In_1716);
xor U1001 (N_1001,In_587,In_1074);
nor U1002 (N_1002,In_797,In_160);
nor U1003 (N_1003,In_1565,In_453);
xnor U1004 (N_1004,In_1568,In_1024);
xnor U1005 (N_1005,In_53,In_753);
nand U1006 (N_1006,In_3,In_36);
and U1007 (N_1007,In_1543,In_148);
or U1008 (N_1008,In_410,In_435);
and U1009 (N_1009,In_252,In_1104);
nand U1010 (N_1010,In_987,In_1198);
nor U1011 (N_1011,In_562,In_213);
nor U1012 (N_1012,In_1018,In_1714);
nand U1013 (N_1013,In_783,In_1513);
or U1014 (N_1014,In_151,In_612);
and U1015 (N_1015,In_1000,In_501);
nand U1016 (N_1016,In_556,In_793);
and U1017 (N_1017,In_1383,In_911);
nand U1018 (N_1018,In_1033,In_890);
and U1019 (N_1019,In_1291,In_1297);
or U1020 (N_1020,In_1324,In_678);
nor U1021 (N_1021,In_1681,In_231);
or U1022 (N_1022,In_1488,In_1492);
nor U1023 (N_1023,In_477,In_907);
and U1024 (N_1024,In_1137,In_1670);
and U1025 (N_1025,In_1336,In_345);
or U1026 (N_1026,In_1312,In_1034);
or U1027 (N_1027,In_1112,In_1626);
and U1028 (N_1028,In_1991,In_452);
or U1029 (N_1029,In_157,In_1497);
nand U1030 (N_1030,In_1009,In_1373);
or U1031 (N_1031,In_487,In_1733);
nand U1032 (N_1032,In_926,In_1339);
and U1033 (N_1033,In_956,In_1190);
nor U1034 (N_1034,In_879,In_1692);
and U1035 (N_1035,In_692,In_463);
nand U1036 (N_1036,In_108,In_1911);
and U1037 (N_1037,In_1623,In_1511);
or U1038 (N_1038,In_1110,In_1442);
and U1039 (N_1039,In_1135,In_1141);
and U1040 (N_1040,In_1787,In_1289);
nand U1041 (N_1041,In_876,In_923);
or U1042 (N_1042,In_461,In_1480);
xnor U1043 (N_1043,In_1587,In_1536);
and U1044 (N_1044,In_1544,In_387);
xnor U1045 (N_1045,In_812,In_1544);
and U1046 (N_1046,In_796,In_787);
and U1047 (N_1047,In_1583,In_388);
xor U1048 (N_1048,In_1466,In_491);
xnor U1049 (N_1049,In_1021,In_1016);
nor U1050 (N_1050,In_756,In_1426);
nand U1051 (N_1051,In_1114,In_953);
nand U1052 (N_1052,In_1057,In_153);
nand U1053 (N_1053,In_998,In_1744);
or U1054 (N_1054,In_395,In_490);
nor U1055 (N_1055,In_1235,In_1694);
or U1056 (N_1056,In_971,In_1598);
xor U1057 (N_1057,In_1669,In_1066);
and U1058 (N_1058,In_1876,In_189);
or U1059 (N_1059,In_1640,In_1306);
and U1060 (N_1060,In_886,In_659);
and U1061 (N_1061,In_1820,In_159);
and U1062 (N_1062,In_1712,In_1328);
xor U1063 (N_1063,In_1266,In_1543);
or U1064 (N_1064,In_50,In_851);
nand U1065 (N_1065,In_883,In_188);
and U1066 (N_1066,In_1585,In_1693);
xor U1067 (N_1067,In_772,In_53);
nand U1068 (N_1068,In_450,In_1291);
nand U1069 (N_1069,In_1890,In_507);
nor U1070 (N_1070,In_1812,In_778);
and U1071 (N_1071,In_303,In_1171);
xor U1072 (N_1072,In_24,In_1011);
xnor U1073 (N_1073,In_934,In_1781);
xor U1074 (N_1074,In_1037,In_1280);
nor U1075 (N_1075,In_1002,In_1046);
and U1076 (N_1076,In_27,In_410);
nor U1077 (N_1077,In_471,In_1354);
and U1078 (N_1078,In_978,In_1918);
and U1079 (N_1079,In_285,In_481);
xnor U1080 (N_1080,In_1421,In_17);
xnor U1081 (N_1081,In_909,In_1983);
nor U1082 (N_1082,In_1973,In_703);
or U1083 (N_1083,In_1681,In_289);
nor U1084 (N_1084,In_1893,In_208);
nand U1085 (N_1085,In_1622,In_1601);
or U1086 (N_1086,In_826,In_921);
nor U1087 (N_1087,In_209,In_713);
or U1088 (N_1088,In_242,In_986);
nor U1089 (N_1089,In_787,In_0);
or U1090 (N_1090,In_1158,In_1467);
or U1091 (N_1091,In_1902,In_774);
nor U1092 (N_1092,In_1770,In_2);
xor U1093 (N_1093,In_987,In_261);
nand U1094 (N_1094,In_1303,In_1020);
nand U1095 (N_1095,In_1739,In_1738);
nand U1096 (N_1096,In_471,In_1312);
and U1097 (N_1097,In_1026,In_335);
nor U1098 (N_1098,In_327,In_170);
or U1099 (N_1099,In_224,In_1413);
xnor U1100 (N_1100,In_780,In_422);
and U1101 (N_1101,In_348,In_225);
xor U1102 (N_1102,In_154,In_1270);
or U1103 (N_1103,In_752,In_1877);
nand U1104 (N_1104,In_1690,In_1904);
or U1105 (N_1105,In_613,In_1760);
xor U1106 (N_1106,In_1640,In_427);
nor U1107 (N_1107,In_1463,In_389);
nand U1108 (N_1108,In_1311,In_1612);
nand U1109 (N_1109,In_598,In_1081);
nor U1110 (N_1110,In_1637,In_1302);
or U1111 (N_1111,In_1556,In_1486);
or U1112 (N_1112,In_535,In_33);
nand U1113 (N_1113,In_1068,In_1145);
and U1114 (N_1114,In_1524,In_1507);
nand U1115 (N_1115,In_980,In_1605);
xnor U1116 (N_1116,In_1874,In_994);
nor U1117 (N_1117,In_651,In_1643);
nor U1118 (N_1118,In_679,In_114);
nor U1119 (N_1119,In_162,In_232);
nor U1120 (N_1120,In_442,In_885);
and U1121 (N_1121,In_283,In_1746);
xor U1122 (N_1122,In_1291,In_168);
xor U1123 (N_1123,In_103,In_1823);
and U1124 (N_1124,In_721,In_1674);
nand U1125 (N_1125,In_1439,In_1685);
nor U1126 (N_1126,In_1121,In_600);
xor U1127 (N_1127,In_809,In_1120);
nor U1128 (N_1128,In_944,In_1852);
or U1129 (N_1129,In_864,In_932);
and U1130 (N_1130,In_1868,In_484);
nand U1131 (N_1131,In_267,In_1533);
and U1132 (N_1132,In_768,In_267);
and U1133 (N_1133,In_364,In_276);
and U1134 (N_1134,In_816,In_972);
nand U1135 (N_1135,In_130,In_1700);
xor U1136 (N_1136,In_1727,In_1509);
nand U1137 (N_1137,In_470,In_1628);
or U1138 (N_1138,In_1953,In_761);
nor U1139 (N_1139,In_1759,In_727);
or U1140 (N_1140,In_878,In_1050);
nand U1141 (N_1141,In_792,In_1088);
xnor U1142 (N_1142,In_581,In_1169);
nor U1143 (N_1143,In_599,In_1047);
and U1144 (N_1144,In_1337,In_771);
xor U1145 (N_1145,In_70,In_525);
nor U1146 (N_1146,In_1516,In_800);
or U1147 (N_1147,In_1132,In_1270);
nand U1148 (N_1148,In_1903,In_190);
nor U1149 (N_1149,In_1882,In_696);
xor U1150 (N_1150,In_1047,In_1062);
xor U1151 (N_1151,In_843,In_1504);
or U1152 (N_1152,In_1094,In_1453);
and U1153 (N_1153,In_1771,In_1619);
or U1154 (N_1154,In_1563,In_55);
or U1155 (N_1155,In_366,In_385);
and U1156 (N_1156,In_1727,In_1537);
xor U1157 (N_1157,In_884,In_881);
and U1158 (N_1158,In_681,In_562);
nor U1159 (N_1159,In_1780,In_1299);
or U1160 (N_1160,In_1049,In_971);
or U1161 (N_1161,In_1790,In_92);
or U1162 (N_1162,In_899,In_980);
nand U1163 (N_1163,In_1638,In_1965);
nand U1164 (N_1164,In_1538,In_1893);
or U1165 (N_1165,In_1414,In_1219);
and U1166 (N_1166,In_749,In_786);
nand U1167 (N_1167,In_606,In_1025);
nor U1168 (N_1168,In_1551,In_1279);
nor U1169 (N_1169,In_1053,In_195);
or U1170 (N_1170,In_1344,In_1041);
nand U1171 (N_1171,In_507,In_1680);
xnor U1172 (N_1172,In_741,In_1266);
or U1173 (N_1173,In_1069,In_1126);
or U1174 (N_1174,In_1729,In_1141);
xnor U1175 (N_1175,In_1347,In_496);
nor U1176 (N_1176,In_1429,In_922);
or U1177 (N_1177,In_1506,In_1109);
nand U1178 (N_1178,In_667,In_118);
and U1179 (N_1179,In_1614,In_1472);
or U1180 (N_1180,In_1447,In_1831);
or U1181 (N_1181,In_405,In_1086);
or U1182 (N_1182,In_1127,In_656);
or U1183 (N_1183,In_44,In_265);
nor U1184 (N_1184,In_1725,In_617);
nor U1185 (N_1185,In_1202,In_1421);
xor U1186 (N_1186,In_280,In_1829);
and U1187 (N_1187,In_950,In_925);
or U1188 (N_1188,In_1647,In_1666);
nand U1189 (N_1189,In_1273,In_1255);
xnor U1190 (N_1190,In_1237,In_965);
nor U1191 (N_1191,In_711,In_653);
or U1192 (N_1192,In_465,In_944);
xnor U1193 (N_1193,In_961,In_833);
xor U1194 (N_1194,In_326,In_1585);
nor U1195 (N_1195,In_1990,In_1538);
or U1196 (N_1196,In_1781,In_35);
xnor U1197 (N_1197,In_1389,In_201);
and U1198 (N_1198,In_46,In_1708);
xnor U1199 (N_1199,In_1650,In_783);
nand U1200 (N_1200,In_651,In_116);
and U1201 (N_1201,In_1046,In_192);
xnor U1202 (N_1202,In_1620,In_1502);
and U1203 (N_1203,In_1350,In_1032);
and U1204 (N_1204,In_195,In_1469);
nor U1205 (N_1205,In_598,In_408);
nor U1206 (N_1206,In_874,In_181);
and U1207 (N_1207,In_718,In_134);
nor U1208 (N_1208,In_967,In_1603);
nand U1209 (N_1209,In_947,In_414);
or U1210 (N_1210,In_1171,In_945);
or U1211 (N_1211,In_1344,In_13);
and U1212 (N_1212,In_1279,In_1918);
xnor U1213 (N_1213,In_1451,In_33);
or U1214 (N_1214,In_378,In_547);
xor U1215 (N_1215,In_1478,In_675);
or U1216 (N_1216,In_1778,In_574);
and U1217 (N_1217,In_894,In_1296);
nand U1218 (N_1218,In_542,In_1102);
and U1219 (N_1219,In_1626,In_1468);
and U1220 (N_1220,In_1751,In_755);
xnor U1221 (N_1221,In_1408,In_1390);
or U1222 (N_1222,In_389,In_19);
nor U1223 (N_1223,In_72,In_227);
and U1224 (N_1224,In_91,In_975);
nor U1225 (N_1225,In_1720,In_510);
nor U1226 (N_1226,In_1202,In_1229);
nor U1227 (N_1227,In_1905,In_618);
or U1228 (N_1228,In_1339,In_1886);
xnor U1229 (N_1229,In_838,In_125);
or U1230 (N_1230,In_260,In_488);
and U1231 (N_1231,In_1983,In_663);
nand U1232 (N_1232,In_1527,In_193);
and U1233 (N_1233,In_1658,In_1772);
or U1234 (N_1234,In_1527,In_1875);
xor U1235 (N_1235,In_1126,In_1900);
nand U1236 (N_1236,In_735,In_1002);
xnor U1237 (N_1237,In_1772,In_743);
nor U1238 (N_1238,In_1093,In_848);
nor U1239 (N_1239,In_671,In_1247);
nand U1240 (N_1240,In_82,In_697);
or U1241 (N_1241,In_142,In_1083);
and U1242 (N_1242,In_565,In_1435);
or U1243 (N_1243,In_704,In_595);
xor U1244 (N_1244,In_1484,In_1463);
nor U1245 (N_1245,In_1638,In_1959);
xnor U1246 (N_1246,In_1384,In_820);
and U1247 (N_1247,In_1303,In_403);
and U1248 (N_1248,In_1180,In_1843);
xor U1249 (N_1249,In_1253,In_885);
or U1250 (N_1250,In_1313,In_970);
nand U1251 (N_1251,In_871,In_1123);
nand U1252 (N_1252,In_1268,In_323);
or U1253 (N_1253,In_1744,In_430);
or U1254 (N_1254,In_1417,In_755);
xnor U1255 (N_1255,In_200,In_520);
xnor U1256 (N_1256,In_329,In_1487);
and U1257 (N_1257,In_1104,In_1107);
or U1258 (N_1258,In_314,In_567);
or U1259 (N_1259,In_462,In_977);
nor U1260 (N_1260,In_1502,In_271);
and U1261 (N_1261,In_160,In_159);
and U1262 (N_1262,In_971,In_1298);
xor U1263 (N_1263,In_447,In_1960);
nor U1264 (N_1264,In_1988,In_483);
or U1265 (N_1265,In_949,In_1259);
and U1266 (N_1266,In_806,In_313);
and U1267 (N_1267,In_1162,In_1218);
nor U1268 (N_1268,In_1307,In_1919);
nand U1269 (N_1269,In_501,In_300);
xnor U1270 (N_1270,In_1178,In_1123);
or U1271 (N_1271,In_1180,In_1553);
and U1272 (N_1272,In_1869,In_956);
nor U1273 (N_1273,In_1504,In_33);
and U1274 (N_1274,In_315,In_1710);
nand U1275 (N_1275,In_1553,In_1555);
and U1276 (N_1276,In_1321,In_436);
or U1277 (N_1277,In_735,In_471);
or U1278 (N_1278,In_1264,In_924);
nand U1279 (N_1279,In_1311,In_160);
xnor U1280 (N_1280,In_646,In_1809);
nor U1281 (N_1281,In_1938,In_1154);
nor U1282 (N_1282,In_1319,In_1141);
and U1283 (N_1283,In_601,In_19);
xnor U1284 (N_1284,In_540,In_782);
nand U1285 (N_1285,In_653,In_987);
nand U1286 (N_1286,In_1006,In_1117);
nand U1287 (N_1287,In_1228,In_1174);
xor U1288 (N_1288,In_48,In_671);
and U1289 (N_1289,In_654,In_1823);
or U1290 (N_1290,In_1945,In_46);
nand U1291 (N_1291,In_1929,In_1791);
and U1292 (N_1292,In_1461,In_810);
xor U1293 (N_1293,In_1635,In_1004);
nand U1294 (N_1294,In_1466,In_827);
or U1295 (N_1295,In_1398,In_390);
or U1296 (N_1296,In_1576,In_678);
nor U1297 (N_1297,In_1327,In_308);
or U1298 (N_1298,In_1857,In_899);
nor U1299 (N_1299,In_900,In_1619);
xor U1300 (N_1300,In_32,In_524);
xnor U1301 (N_1301,In_1968,In_501);
and U1302 (N_1302,In_933,In_1440);
nor U1303 (N_1303,In_1090,In_1475);
and U1304 (N_1304,In_1756,In_413);
nand U1305 (N_1305,In_200,In_1729);
or U1306 (N_1306,In_72,In_1351);
nor U1307 (N_1307,In_721,In_96);
xor U1308 (N_1308,In_843,In_1125);
nor U1309 (N_1309,In_1231,In_1190);
nor U1310 (N_1310,In_458,In_1719);
nand U1311 (N_1311,In_1083,In_322);
xnor U1312 (N_1312,In_1685,In_770);
nand U1313 (N_1313,In_1237,In_820);
xnor U1314 (N_1314,In_537,In_1389);
and U1315 (N_1315,In_1511,In_250);
and U1316 (N_1316,In_1489,In_599);
nor U1317 (N_1317,In_609,In_125);
or U1318 (N_1318,In_568,In_1683);
nor U1319 (N_1319,In_174,In_998);
nand U1320 (N_1320,In_708,In_1822);
or U1321 (N_1321,In_1356,In_1983);
nand U1322 (N_1322,In_451,In_1299);
xnor U1323 (N_1323,In_1971,In_434);
xor U1324 (N_1324,In_1199,In_1213);
and U1325 (N_1325,In_3,In_1711);
xor U1326 (N_1326,In_1522,In_1295);
nand U1327 (N_1327,In_1679,In_630);
nand U1328 (N_1328,In_1436,In_575);
and U1329 (N_1329,In_1282,In_247);
and U1330 (N_1330,In_1761,In_187);
nand U1331 (N_1331,In_757,In_471);
xnor U1332 (N_1332,In_1836,In_1702);
nor U1333 (N_1333,In_1076,In_1522);
xor U1334 (N_1334,In_1573,In_1414);
xor U1335 (N_1335,In_1515,In_1433);
nand U1336 (N_1336,In_1900,In_1072);
xnor U1337 (N_1337,In_1458,In_1084);
nand U1338 (N_1338,In_919,In_621);
or U1339 (N_1339,In_1628,In_814);
and U1340 (N_1340,In_616,In_1000);
nand U1341 (N_1341,In_977,In_1489);
xor U1342 (N_1342,In_1439,In_8);
or U1343 (N_1343,In_819,In_161);
nor U1344 (N_1344,In_12,In_1400);
nand U1345 (N_1345,In_1947,In_118);
nand U1346 (N_1346,In_87,In_1289);
nand U1347 (N_1347,In_1350,In_1741);
nand U1348 (N_1348,In_870,In_1322);
nor U1349 (N_1349,In_1939,In_1123);
nand U1350 (N_1350,In_1106,In_1341);
nor U1351 (N_1351,In_1100,In_1343);
nor U1352 (N_1352,In_344,In_251);
or U1353 (N_1353,In_1888,In_1771);
and U1354 (N_1354,In_416,In_179);
nor U1355 (N_1355,In_1444,In_136);
xor U1356 (N_1356,In_987,In_929);
or U1357 (N_1357,In_741,In_710);
or U1358 (N_1358,In_907,In_880);
nor U1359 (N_1359,In_1438,In_798);
xnor U1360 (N_1360,In_878,In_1003);
nor U1361 (N_1361,In_728,In_302);
nor U1362 (N_1362,In_1714,In_760);
nand U1363 (N_1363,In_327,In_136);
or U1364 (N_1364,In_143,In_1006);
and U1365 (N_1365,In_1375,In_1382);
nand U1366 (N_1366,In_1127,In_313);
or U1367 (N_1367,In_496,In_301);
or U1368 (N_1368,In_579,In_461);
nand U1369 (N_1369,In_942,In_1075);
nand U1370 (N_1370,In_923,In_1631);
nor U1371 (N_1371,In_596,In_748);
nor U1372 (N_1372,In_641,In_1538);
nand U1373 (N_1373,In_1748,In_1216);
and U1374 (N_1374,In_1254,In_788);
xnor U1375 (N_1375,In_407,In_1771);
and U1376 (N_1376,In_739,In_649);
and U1377 (N_1377,In_292,In_39);
and U1378 (N_1378,In_783,In_1923);
and U1379 (N_1379,In_496,In_1624);
nand U1380 (N_1380,In_1306,In_486);
nand U1381 (N_1381,In_808,In_1371);
nor U1382 (N_1382,In_196,In_1044);
nand U1383 (N_1383,In_512,In_1140);
nor U1384 (N_1384,In_1256,In_557);
xnor U1385 (N_1385,In_1395,In_277);
and U1386 (N_1386,In_1670,In_1545);
nor U1387 (N_1387,In_1079,In_796);
nor U1388 (N_1388,In_1634,In_277);
nor U1389 (N_1389,In_316,In_1945);
nor U1390 (N_1390,In_1395,In_1713);
nor U1391 (N_1391,In_470,In_574);
xor U1392 (N_1392,In_1543,In_1219);
or U1393 (N_1393,In_851,In_361);
nor U1394 (N_1394,In_1069,In_368);
or U1395 (N_1395,In_981,In_1726);
nor U1396 (N_1396,In_783,In_1574);
and U1397 (N_1397,In_47,In_1582);
nand U1398 (N_1398,In_699,In_1370);
and U1399 (N_1399,In_1580,In_1145);
and U1400 (N_1400,In_1147,In_739);
nand U1401 (N_1401,In_1928,In_151);
or U1402 (N_1402,In_162,In_760);
nand U1403 (N_1403,In_1278,In_1462);
xnor U1404 (N_1404,In_912,In_1341);
xnor U1405 (N_1405,In_626,In_890);
and U1406 (N_1406,In_19,In_1920);
nor U1407 (N_1407,In_914,In_527);
and U1408 (N_1408,In_1870,In_1959);
nand U1409 (N_1409,In_190,In_1319);
nand U1410 (N_1410,In_268,In_1086);
xor U1411 (N_1411,In_1469,In_1960);
xor U1412 (N_1412,In_889,In_1904);
nor U1413 (N_1413,In_334,In_1695);
nor U1414 (N_1414,In_1124,In_194);
nand U1415 (N_1415,In_1300,In_549);
nand U1416 (N_1416,In_613,In_369);
nand U1417 (N_1417,In_89,In_1969);
or U1418 (N_1418,In_533,In_1480);
xnor U1419 (N_1419,In_863,In_1412);
and U1420 (N_1420,In_1325,In_1086);
nand U1421 (N_1421,In_1404,In_853);
nand U1422 (N_1422,In_199,In_557);
nand U1423 (N_1423,In_1099,In_184);
and U1424 (N_1424,In_1152,In_426);
nor U1425 (N_1425,In_105,In_1792);
and U1426 (N_1426,In_1005,In_959);
xnor U1427 (N_1427,In_1803,In_820);
nor U1428 (N_1428,In_1705,In_178);
nand U1429 (N_1429,In_1477,In_1439);
xor U1430 (N_1430,In_1206,In_1735);
nand U1431 (N_1431,In_1244,In_1700);
xor U1432 (N_1432,In_1500,In_110);
and U1433 (N_1433,In_1142,In_42);
and U1434 (N_1434,In_1899,In_1494);
or U1435 (N_1435,In_1165,In_1544);
and U1436 (N_1436,In_1844,In_1352);
nor U1437 (N_1437,In_1698,In_71);
or U1438 (N_1438,In_444,In_1413);
xor U1439 (N_1439,In_1497,In_1769);
nand U1440 (N_1440,In_1399,In_1302);
xnor U1441 (N_1441,In_1310,In_1657);
nand U1442 (N_1442,In_325,In_626);
and U1443 (N_1443,In_893,In_1428);
or U1444 (N_1444,In_308,In_1947);
nor U1445 (N_1445,In_429,In_929);
nand U1446 (N_1446,In_1939,In_348);
xor U1447 (N_1447,In_934,In_471);
or U1448 (N_1448,In_1617,In_987);
nor U1449 (N_1449,In_1048,In_1228);
nand U1450 (N_1450,In_353,In_972);
xnor U1451 (N_1451,In_777,In_960);
and U1452 (N_1452,In_1219,In_238);
nor U1453 (N_1453,In_48,In_1084);
xnor U1454 (N_1454,In_1220,In_390);
or U1455 (N_1455,In_1230,In_473);
xor U1456 (N_1456,In_1111,In_1346);
nor U1457 (N_1457,In_1474,In_1311);
xnor U1458 (N_1458,In_1441,In_1973);
and U1459 (N_1459,In_194,In_1023);
and U1460 (N_1460,In_1533,In_1691);
or U1461 (N_1461,In_299,In_1794);
or U1462 (N_1462,In_877,In_784);
xor U1463 (N_1463,In_740,In_693);
and U1464 (N_1464,In_1463,In_883);
and U1465 (N_1465,In_958,In_1955);
nor U1466 (N_1466,In_1150,In_1752);
nor U1467 (N_1467,In_1752,In_1184);
nand U1468 (N_1468,In_88,In_1176);
or U1469 (N_1469,In_1515,In_1825);
xnor U1470 (N_1470,In_126,In_431);
or U1471 (N_1471,In_1507,In_1607);
xor U1472 (N_1472,In_1180,In_1608);
nor U1473 (N_1473,In_1410,In_1625);
or U1474 (N_1474,In_535,In_728);
or U1475 (N_1475,In_1651,In_582);
or U1476 (N_1476,In_1550,In_1679);
or U1477 (N_1477,In_1482,In_220);
nor U1478 (N_1478,In_1316,In_139);
and U1479 (N_1479,In_1931,In_318);
nor U1480 (N_1480,In_665,In_342);
and U1481 (N_1481,In_6,In_407);
nand U1482 (N_1482,In_1193,In_733);
or U1483 (N_1483,In_244,In_1272);
and U1484 (N_1484,In_1015,In_464);
nor U1485 (N_1485,In_281,In_835);
nor U1486 (N_1486,In_490,In_172);
xor U1487 (N_1487,In_1498,In_627);
nor U1488 (N_1488,In_701,In_1217);
xnor U1489 (N_1489,In_1961,In_409);
and U1490 (N_1490,In_134,In_1093);
and U1491 (N_1491,In_410,In_1372);
or U1492 (N_1492,In_1773,In_1210);
xnor U1493 (N_1493,In_1916,In_1061);
nor U1494 (N_1494,In_334,In_1556);
or U1495 (N_1495,In_1972,In_161);
xnor U1496 (N_1496,In_1077,In_527);
or U1497 (N_1497,In_1882,In_1597);
or U1498 (N_1498,In_1275,In_343);
nor U1499 (N_1499,In_1916,In_384);
or U1500 (N_1500,In_274,In_411);
or U1501 (N_1501,In_1128,In_998);
nand U1502 (N_1502,In_1259,In_1383);
nand U1503 (N_1503,In_1483,In_394);
nor U1504 (N_1504,In_629,In_775);
xnor U1505 (N_1505,In_1487,In_478);
and U1506 (N_1506,In_533,In_108);
xnor U1507 (N_1507,In_316,In_1305);
and U1508 (N_1508,In_140,In_1044);
or U1509 (N_1509,In_1335,In_1985);
nand U1510 (N_1510,In_1999,In_1685);
or U1511 (N_1511,In_1178,In_1959);
nor U1512 (N_1512,In_865,In_826);
or U1513 (N_1513,In_618,In_1340);
or U1514 (N_1514,In_1733,In_1633);
nand U1515 (N_1515,In_1088,In_983);
or U1516 (N_1516,In_1052,In_1385);
or U1517 (N_1517,In_931,In_893);
nor U1518 (N_1518,In_608,In_1364);
and U1519 (N_1519,In_68,In_1473);
and U1520 (N_1520,In_582,In_268);
and U1521 (N_1521,In_1024,In_129);
xor U1522 (N_1522,In_1249,In_999);
or U1523 (N_1523,In_1055,In_1220);
and U1524 (N_1524,In_1465,In_793);
or U1525 (N_1525,In_495,In_1983);
nand U1526 (N_1526,In_1764,In_1852);
xor U1527 (N_1527,In_27,In_1308);
or U1528 (N_1528,In_1432,In_1940);
or U1529 (N_1529,In_1729,In_1841);
nand U1530 (N_1530,In_128,In_1592);
and U1531 (N_1531,In_1316,In_1312);
nor U1532 (N_1532,In_391,In_1604);
or U1533 (N_1533,In_835,In_1091);
nand U1534 (N_1534,In_435,In_1328);
or U1535 (N_1535,In_800,In_819);
nand U1536 (N_1536,In_698,In_1036);
or U1537 (N_1537,In_1941,In_1469);
or U1538 (N_1538,In_127,In_1951);
nand U1539 (N_1539,In_989,In_1444);
or U1540 (N_1540,In_1060,In_1756);
xor U1541 (N_1541,In_1088,In_1021);
nor U1542 (N_1542,In_851,In_698);
xnor U1543 (N_1543,In_1782,In_452);
or U1544 (N_1544,In_547,In_1419);
xor U1545 (N_1545,In_535,In_1333);
nand U1546 (N_1546,In_1041,In_1347);
or U1547 (N_1547,In_1820,In_948);
xor U1548 (N_1548,In_1636,In_1645);
nor U1549 (N_1549,In_280,In_1023);
nand U1550 (N_1550,In_1201,In_287);
xnor U1551 (N_1551,In_1891,In_1158);
or U1552 (N_1552,In_450,In_1290);
nand U1553 (N_1553,In_371,In_968);
xor U1554 (N_1554,In_1229,In_857);
nand U1555 (N_1555,In_919,In_1325);
or U1556 (N_1556,In_460,In_895);
nor U1557 (N_1557,In_1534,In_1266);
and U1558 (N_1558,In_1755,In_500);
nand U1559 (N_1559,In_495,In_1124);
nor U1560 (N_1560,In_1525,In_595);
and U1561 (N_1561,In_673,In_488);
nor U1562 (N_1562,In_974,In_1509);
and U1563 (N_1563,In_359,In_1697);
nor U1564 (N_1564,In_316,In_1067);
and U1565 (N_1565,In_1976,In_846);
nor U1566 (N_1566,In_95,In_454);
or U1567 (N_1567,In_885,In_1409);
xnor U1568 (N_1568,In_1915,In_260);
and U1569 (N_1569,In_613,In_638);
or U1570 (N_1570,In_1567,In_1257);
nand U1571 (N_1571,In_1547,In_76);
xnor U1572 (N_1572,In_1410,In_106);
xnor U1573 (N_1573,In_561,In_1153);
and U1574 (N_1574,In_826,In_1902);
or U1575 (N_1575,In_715,In_1453);
nand U1576 (N_1576,In_853,In_622);
nor U1577 (N_1577,In_69,In_290);
and U1578 (N_1578,In_1529,In_1950);
nand U1579 (N_1579,In_1445,In_1855);
and U1580 (N_1580,In_909,In_703);
xor U1581 (N_1581,In_1393,In_1722);
nor U1582 (N_1582,In_121,In_404);
xor U1583 (N_1583,In_1749,In_1900);
nor U1584 (N_1584,In_328,In_905);
and U1585 (N_1585,In_265,In_1853);
or U1586 (N_1586,In_1468,In_358);
or U1587 (N_1587,In_580,In_184);
nand U1588 (N_1588,In_1048,In_342);
and U1589 (N_1589,In_747,In_819);
xnor U1590 (N_1590,In_1062,In_175);
xor U1591 (N_1591,In_374,In_491);
xor U1592 (N_1592,In_1113,In_1664);
nor U1593 (N_1593,In_918,In_1638);
nor U1594 (N_1594,In_1937,In_767);
xor U1595 (N_1595,In_570,In_1006);
or U1596 (N_1596,In_801,In_203);
xor U1597 (N_1597,In_1810,In_1602);
nor U1598 (N_1598,In_1721,In_851);
nor U1599 (N_1599,In_1521,In_1268);
nor U1600 (N_1600,In_1625,In_1012);
nor U1601 (N_1601,In_1852,In_464);
nand U1602 (N_1602,In_564,In_1425);
and U1603 (N_1603,In_563,In_1755);
nor U1604 (N_1604,In_658,In_1373);
and U1605 (N_1605,In_1708,In_1188);
nand U1606 (N_1606,In_1136,In_1886);
nand U1607 (N_1607,In_1634,In_390);
and U1608 (N_1608,In_1006,In_606);
nor U1609 (N_1609,In_1598,In_1413);
nor U1610 (N_1610,In_1954,In_805);
nand U1611 (N_1611,In_1881,In_1099);
and U1612 (N_1612,In_614,In_1786);
nor U1613 (N_1613,In_1688,In_66);
or U1614 (N_1614,In_1340,In_584);
and U1615 (N_1615,In_1324,In_830);
nor U1616 (N_1616,In_1085,In_28);
or U1617 (N_1617,In_1659,In_914);
and U1618 (N_1618,In_818,In_895);
and U1619 (N_1619,In_1735,In_1556);
or U1620 (N_1620,In_1490,In_1710);
xnor U1621 (N_1621,In_408,In_1450);
xnor U1622 (N_1622,In_1728,In_617);
or U1623 (N_1623,In_1784,In_1577);
xor U1624 (N_1624,In_820,In_1690);
nand U1625 (N_1625,In_1103,In_787);
nor U1626 (N_1626,In_1993,In_321);
nand U1627 (N_1627,In_1766,In_354);
nor U1628 (N_1628,In_1464,In_838);
and U1629 (N_1629,In_1988,In_358);
xor U1630 (N_1630,In_1089,In_1838);
and U1631 (N_1631,In_1630,In_781);
xor U1632 (N_1632,In_1566,In_969);
or U1633 (N_1633,In_87,In_1861);
nor U1634 (N_1634,In_465,In_1402);
nand U1635 (N_1635,In_119,In_1976);
or U1636 (N_1636,In_520,In_467);
nor U1637 (N_1637,In_1925,In_1987);
or U1638 (N_1638,In_1307,In_1955);
and U1639 (N_1639,In_518,In_1217);
nand U1640 (N_1640,In_1970,In_104);
xnor U1641 (N_1641,In_836,In_1709);
and U1642 (N_1642,In_1888,In_1784);
and U1643 (N_1643,In_1815,In_271);
and U1644 (N_1644,In_471,In_1628);
and U1645 (N_1645,In_1902,In_252);
nor U1646 (N_1646,In_1251,In_610);
nor U1647 (N_1647,In_1975,In_1538);
nor U1648 (N_1648,In_1007,In_9);
nor U1649 (N_1649,In_804,In_191);
nand U1650 (N_1650,In_1494,In_213);
xnor U1651 (N_1651,In_913,In_377);
or U1652 (N_1652,In_246,In_898);
nand U1653 (N_1653,In_1585,In_1011);
or U1654 (N_1654,In_1543,In_150);
and U1655 (N_1655,In_1642,In_826);
or U1656 (N_1656,In_186,In_1618);
nand U1657 (N_1657,In_1573,In_1282);
nor U1658 (N_1658,In_131,In_692);
xor U1659 (N_1659,In_493,In_331);
xor U1660 (N_1660,In_891,In_800);
nor U1661 (N_1661,In_268,In_991);
xor U1662 (N_1662,In_1701,In_1996);
nor U1663 (N_1663,In_230,In_918);
xnor U1664 (N_1664,In_1699,In_1297);
nand U1665 (N_1665,In_1774,In_1723);
and U1666 (N_1666,In_337,In_1496);
and U1667 (N_1667,In_688,In_329);
and U1668 (N_1668,In_239,In_1782);
xor U1669 (N_1669,In_976,In_171);
nor U1670 (N_1670,In_880,In_583);
nand U1671 (N_1671,In_391,In_1662);
nand U1672 (N_1672,In_1342,In_398);
and U1673 (N_1673,In_1368,In_1973);
xor U1674 (N_1674,In_1733,In_143);
nor U1675 (N_1675,In_1529,In_927);
xnor U1676 (N_1676,In_1337,In_1516);
nor U1677 (N_1677,In_921,In_1911);
nor U1678 (N_1678,In_487,In_1709);
nor U1679 (N_1679,In_596,In_1340);
and U1680 (N_1680,In_517,In_871);
or U1681 (N_1681,In_311,In_546);
and U1682 (N_1682,In_741,In_850);
xor U1683 (N_1683,In_1094,In_1384);
nand U1684 (N_1684,In_1145,In_139);
xor U1685 (N_1685,In_343,In_566);
or U1686 (N_1686,In_1478,In_642);
or U1687 (N_1687,In_1100,In_737);
xnor U1688 (N_1688,In_1147,In_1581);
nand U1689 (N_1689,In_134,In_1409);
or U1690 (N_1690,In_1788,In_1482);
nand U1691 (N_1691,In_1415,In_774);
nand U1692 (N_1692,In_561,In_1861);
nor U1693 (N_1693,In_1268,In_1058);
xnor U1694 (N_1694,In_1949,In_452);
and U1695 (N_1695,In_67,In_1339);
nand U1696 (N_1696,In_1652,In_1671);
nand U1697 (N_1697,In_1562,In_1958);
or U1698 (N_1698,In_63,In_377);
and U1699 (N_1699,In_1905,In_1805);
xnor U1700 (N_1700,In_481,In_766);
and U1701 (N_1701,In_1730,In_721);
and U1702 (N_1702,In_46,In_1848);
xor U1703 (N_1703,In_1806,In_177);
nand U1704 (N_1704,In_968,In_158);
nand U1705 (N_1705,In_1112,In_1463);
nor U1706 (N_1706,In_1186,In_297);
nand U1707 (N_1707,In_1659,In_1169);
xor U1708 (N_1708,In_356,In_1845);
and U1709 (N_1709,In_1500,In_1969);
nor U1710 (N_1710,In_586,In_1809);
nor U1711 (N_1711,In_822,In_1041);
nand U1712 (N_1712,In_788,In_204);
and U1713 (N_1713,In_1890,In_1736);
nor U1714 (N_1714,In_884,In_93);
or U1715 (N_1715,In_411,In_1911);
nor U1716 (N_1716,In_873,In_1547);
nand U1717 (N_1717,In_765,In_982);
nand U1718 (N_1718,In_376,In_1730);
or U1719 (N_1719,In_714,In_99);
xnor U1720 (N_1720,In_1184,In_1716);
xnor U1721 (N_1721,In_1819,In_574);
nor U1722 (N_1722,In_1376,In_1419);
nor U1723 (N_1723,In_1607,In_976);
xnor U1724 (N_1724,In_949,In_555);
nor U1725 (N_1725,In_1528,In_108);
nor U1726 (N_1726,In_1854,In_1819);
nor U1727 (N_1727,In_271,In_952);
and U1728 (N_1728,In_31,In_1085);
or U1729 (N_1729,In_1647,In_1367);
or U1730 (N_1730,In_1582,In_1750);
and U1731 (N_1731,In_122,In_32);
nand U1732 (N_1732,In_1950,In_182);
nand U1733 (N_1733,In_1431,In_1639);
nand U1734 (N_1734,In_561,In_160);
and U1735 (N_1735,In_338,In_1638);
xor U1736 (N_1736,In_1218,In_613);
nor U1737 (N_1737,In_1788,In_397);
xnor U1738 (N_1738,In_1815,In_1759);
and U1739 (N_1739,In_533,In_746);
nand U1740 (N_1740,In_1738,In_218);
xor U1741 (N_1741,In_955,In_83);
nand U1742 (N_1742,In_1336,In_1130);
and U1743 (N_1743,In_448,In_613);
or U1744 (N_1744,In_200,In_362);
nor U1745 (N_1745,In_86,In_584);
and U1746 (N_1746,In_1792,In_1408);
or U1747 (N_1747,In_1952,In_1359);
nor U1748 (N_1748,In_1178,In_1446);
or U1749 (N_1749,In_639,In_1671);
nand U1750 (N_1750,In_1929,In_1602);
nor U1751 (N_1751,In_687,In_1938);
nor U1752 (N_1752,In_1396,In_1359);
xnor U1753 (N_1753,In_1216,In_1706);
xnor U1754 (N_1754,In_871,In_124);
xor U1755 (N_1755,In_233,In_225);
xnor U1756 (N_1756,In_161,In_1653);
xnor U1757 (N_1757,In_1631,In_865);
and U1758 (N_1758,In_1224,In_1320);
and U1759 (N_1759,In_1664,In_1073);
or U1760 (N_1760,In_611,In_1719);
xor U1761 (N_1761,In_772,In_82);
nand U1762 (N_1762,In_143,In_460);
nor U1763 (N_1763,In_1947,In_1055);
and U1764 (N_1764,In_1075,In_1480);
nor U1765 (N_1765,In_1242,In_1945);
and U1766 (N_1766,In_331,In_659);
xnor U1767 (N_1767,In_956,In_359);
xnor U1768 (N_1768,In_1877,In_318);
nand U1769 (N_1769,In_1485,In_3);
nor U1770 (N_1770,In_1156,In_1763);
nor U1771 (N_1771,In_1509,In_1440);
or U1772 (N_1772,In_1893,In_20);
or U1773 (N_1773,In_942,In_475);
xnor U1774 (N_1774,In_304,In_707);
or U1775 (N_1775,In_406,In_224);
and U1776 (N_1776,In_1643,In_1761);
and U1777 (N_1777,In_197,In_1526);
nand U1778 (N_1778,In_1842,In_682);
nand U1779 (N_1779,In_111,In_1912);
nand U1780 (N_1780,In_1492,In_1140);
nor U1781 (N_1781,In_1798,In_1939);
and U1782 (N_1782,In_727,In_1557);
or U1783 (N_1783,In_814,In_1036);
or U1784 (N_1784,In_1196,In_849);
or U1785 (N_1785,In_1492,In_1502);
nor U1786 (N_1786,In_590,In_957);
xor U1787 (N_1787,In_1731,In_1428);
nor U1788 (N_1788,In_1369,In_1245);
or U1789 (N_1789,In_1731,In_504);
nand U1790 (N_1790,In_1656,In_1868);
or U1791 (N_1791,In_774,In_660);
nand U1792 (N_1792,In_1941,In_1614);
or U1793 (N_1793,In_257,In_1123);
nand U1794 (N_1794,In_83,In_1841);
nor U1795 (N_1795,In_605,In_1473);
nand U1796 (N_1796,In_1,In_1214);
nor U1797 (N_1797,In_1300,In_71);
and U1798 (N_1798,In_975,In_651);
xor U1799 (N_1799,In_841,In_1665);
nor U1800 (N_1800,In_600,In_576);
nand U1801 (N_1801,In_434,In_1479);
and U1802 (N_1802,In_1203,In_1136);
xor U1803 (N_1803,In_1715,In_1881);
xor U1804 (N_1804,In_182,In_144);
and U1805 (N_1805,In_1036,In_1812);
and U1806 (N_1806,In_541,In_1364);
and U1807 (N_1807,In_449,In_1580);
and U1808 (N_1808,In_851,In_1919);
and U1809 (N_1809,In_699,In_1805);
xnor U1810 (N_1810,In_51,In_1878);
nor U1811 (N_1811,In_1921,In_1908);
and U1812 (N_1812,In_396,In_418);
xor U1813 (N_1813,In_1009,In_845);
nor U1814 (N_1814,In_1823,In_1862);
nor U1815 (N_1815,In_1711,In_70);
nand U1816 (N_1816,In_1898,In_979);
and U1817 (N_1817,In_878,In_178);
or U1818 (N_1818,In_87,In_71);
nand U1819 (N_1819,In_1818,In_708);
xor U1820 (N_1820,In_1162,In_640);
or U1821 (N_1821,In_672,In_1099);
xnor U1822 (N_1822,In_1751,In_1668);
or U1823 (N_1823,In_1265,In_513);
nor U1824 (N_1824,In_1223,In_1331);
and U1825 (N_1825,In_1982,In_1230);
xnor U1826 (N_1826,In_23,In_1838);
nand U1827 (N_1827,In_821,In_202);
or U1828 (N_1828,In_858,In_733);
or U1829 (N_1829,In_1297,In_1604);
or U1830 (N_1830,In_1656,In_1877);
nand U1831 (N_1831,In_478,In_358);
and U1832 (N_1832,In_1258,In_1610);
or U1833 (N_1833,In_395,In_1457);
nor U1834 (N_1834,In_1533,In_686);
nor U1835 (N_1835,In_976,In_478);
xor U1836 (N_1836,In_15,In_1358);
or U1837 (N_1837,In_201,In_1405);
nand U1838 (N_1838,In_739,In_501);
or U1839 (N_1839,In_1044,In_1344);
nand U1840 (N_1840,In_1315,In_1847);
xnor U1841 (N_1841,In_1052,In_1321);
xnor U1842 (N_1842,In_1938,In_1425);
nor U1843 (N_1843,In_194,In_1426);
or U1844 (N_1844,In_1648,In_291);
nand U1845 (N_1845,In_515,In_655);
xor U1846 (N_1846,In_507,In_937);
nor U1847 (N_1847,In_1686,In_1988);
and U1848 (N_1848,In_1894,In_562);
or U1849 (N_1849,In_937,In_954);
xnor U1850 (N_1850,In_726,In_1983);
or U1851 (N_1851,In_850,In_954);
or U1852 (N_1852,In_1837,In_979);
and U1853 (N_1853,In_718,In_1733);
xnor U1854 (N_1854,In_208,In_1734);
and U1855 (N_1855,In_1773,In_1715);
nand U1856 (N_1856,In_1259,In_313);
and U1857 (N_1857,In_1492,In_1516);
or U1858 (N_1858,In_240,In_1227);
xor U1859 (N_1859,In_1791,In_1056);
xnor U1860 (N_1860,In_1445,In_805);
xnor U1861 (N_1861,In_1664,In_577);
and U1862 (N_1862,In_476,In_960);
and U1863 (N_1863,In_1541,In_1148);
or U1864 (N_1864,In_1890,In_1028);
nand U1865 (N_1865,In_596,In_1020);
nand U1866 (N_1866,In_76,In_389);
nor U1867 (N_1867,In_1215,In_439);
nor U1868 (N_1868,In_1401,In_458);
nor U1869 (N_1869,In_325,In_304);
nand U1870 (N_1870,In_673,In_550);
nand U1871 (N_1871,In_202,In_1995);
xor U1872 (N_1872,In_884,In_1855);
nor U1873 (N_1873,In_517,In_228);
and U1874 (N_1874,In_1967,In_285);
nor U1875 (N_1875,In_199,In_1796);
nand U1876 (N_1876,In_1858,In_11);
and U1877 (N_1877,In_92,In_300);
nand U1878 (N_1878,In_52,In_1364);
xnor U1879 (N_1879,In_539,In_18);
or U1880 (N_1880,In_1145,In_1276);
xor U1881 (N_1881,In_204,In_1708);
xnor U1882 (N_1882,In_1502,In_949);
nor U1883 (N_1883,In_1926,In_1386);
xor U1884 (N_1884,In_1245,In_1525);
nor U1885 (N_1885,In_1793,In_1470);
nor U1886 (N_1886,In_1497,In_1816);
nand U1887 (N_1887,In_4,In_1118);
xor U1888 (N_1888,In_183,In_1720);
xor U1889 (N_1889,In_37,In_1064);
or U1890 (N_1890,In_1165,In_1994);
and U1891 (N_1891,In_531,In_313);
or U1892 (N_1892,In_906,In_444);
xnor U1893 (N_1893,In_76,In_414);
nor U1894 (N_1894,In_635,In_5);
or U1895 (N_1895,In_943,In_1812);
nand U1896 (N_1896,In_1250,In_1674);
or U1897 (N_1897,In_1392,In_1190);
nor U1898 (N_1898,In_1054,In_404);
or U1899 (N_1899,In_1230,In_651);
xnor U1900 (N_1900,In_566,In_1438);
nand U1901 (N_1901,In_1836,In_414);
nand U1902 (N_1902,In_678,In_1558);
nand U1903 (N_1903,In_251,In_869);
or U1904 (N_1904,In_1745,In_672);
nand U1905 (N_1905,In_1854,In_73);
nor U1906 (N_1906,In_62,In_504);
and U1907 (N_1907,In_1985,In_1003);
xor U1908 (N_1908,In_1298,In_1059);
and U1909 (N_1909,In_1848,In_1469);
or U1910 (N_1910,In_1028,In_661);
nor U1911 (N_1911,In_1528,In_603);
and U1912 (N_1912,In_1016,In_988);
nor U1913 (N_1913,In_723,In_1258);
nand U1914 (N_1914,In_359,In_545);
xor U1915 (N_1915,In_958,In_179);
nand U1916 (N_1916,In_607,In_1971);
or U1917 (N_1917,In_1893,In_1530);
or U1918 (N_1918,In_1030,In_170);
xor U1919 (N_1919,In_853,In_320);
nor U1920 (N_1920,In_581,In_305);
nor U1921 (N_1921,In_1179,In_932);
xnor U1922 (N_1922,In_1469,In_1873);
xor U1923 (N_1923,In_1672,In_1402);
nor U1924 (N_1924,In_955,In_654);
nand U1925 (N_1925,In_969,In_1827);
nand U1926 (N_1926,In_1025,In_390);
nand U1927 (N_1927,In_765,In_129);
nor U1928 (N_1928,In_1619,In_1465);
xnor U1929 (N_1929,In_813,In_1345);
and U1930 (N_1930,In_350,In_1017);
or U1931 (N_1931,In_1130,In_1201);
or U1932 (N_1932,In_1811,In_1847);
xor U1933 (N_1933,In_1815,In_476);
or U1934 (N_1934,In_1252,In_900);
nand U1935 (N_1935,In_507,In_159);
and U1936 (N_1936,In_506,In_1980);
and U1937 (N_1937,In_1879,In_1473);
nor U1938 (N_1938,In_929,In_1782);
xor U1939 (N_1939,In_1337,In_1933);
or U1940 (N_1940,In_1853,In_1047);
or U1941 (N_1941,In_885,In_19);
xor U1942 (N_1942,In_1385,In_1604);
or U1943 (N_1943,In_849,In_1854);
nor U1944 (N_1944,In_1563,In_1778);
and U1945 (N_1945,In_1595,In_1650);
and U1946 (N_1946,In_1430,In_1506);
and U1947 (N_1947,In_1521,In_517);
or U1948 (N_1948,In_80,In_1232);
nor U1949 (N_1949,In_697,In_859);
xnor U1950 (N_1950,In_688,In_657);
and U1951 (N_1951,In_1781,In_1164);
nand U1952 (N_1952,In_1099,In_1127);
xor U1953 (N_1953,In_118,In_1963);
nor U1954 (N_1954,In_242,In_729);
nor U1955 (N_1955,In_394,In_1385);
and U1956 (N_1956,In_362,In_747);
xnor U1957 (N_1957,In_872,In_1065);
or U1958 (N_1958,In_1464,In_21);
or U1959 (N_1959,In_773,In_1470);
nand U1960 (N_1960,In_746,In_1731);
xor U1961 (N_1961,In_868,In_1488);
xor U1962 (N_1962,In_1972,In_1410);
and U1963 (N_1963,In_1682,In_1249);
nand U1964 (N_1964,In_1851,In_43);
nand U1965 (N_1965,In_1594,In_1204);
or U1966 (N_1966,In_731,In_408);
nor U1967 (N_1967,In_406,In_675);
nand U1968 (N_1968,In_1097,In_1707);
or U1969 (N_1969,In_308,In_518);
and U1970 (N_1970,In_1139,In_663);
nor U1971 (N_1971,In_1184,In_1168);
or U1972 (N_1972,In_1623,In_631);
nand U1973 (N_1973,In_1385,In_1694);
nor U1974 (N_1974,In_741,In_988);
and U1975 (N_1975,In_1651,In_1232);
nor U1976 (N_1976,In_1908,In_293);
or U1977 (N_1977,In_1904,In_237);
or U1978 (N_1978,In_1218,In_1314);
nor U1979 (N_1979,In_702,In_1680);
nor U1980 (N_1980,In_685,In_401);
and U1981 (N_1981,In_384,In_1256);
and U1982 (N_1982,In_821,In_1231);
nor U1983 (N_1983,In_1245,In_248);
and U1984 (N_1984,In_1470,In_1579);
or U1985 (N_1985,In_1334,In_235);
nand U1986 (N_1986,In_122,In_1911);
or U1987 (N_1987,In_551,In_1870);
or U1988 (N_1988,In_822,In_1464);
or U1989 (N_1989,In_661,In_1670);
nor U1990 (N_1990,In_1018,In_376);
or U1991 (N_1991,In_435,In_129);
nand U1992 (N_1992,In_1739,In_556);
or U1993 (N_1993,In_42,In_1038);
xnor U1994 (N_1994,In_765,In_975);
xnor U1995 (N_1995,In_1009,In_1069);
nor U1996 (N_1996,In_711,In_1230);
or U1997 (N_1997,In_237,In_861);
nand U1998 (N_1998,In_1867,In_1925);
nor U1999 (N_1999,In_790,In_1435);
nor U2000 (N_2000,In_222,In_29);
and U2001 (N_2001,In_877,In_1658);
or U2002 (N_2002,In_990,In_649);
nor U2003 (N_2003,In_681,In_1613);
or U2004 (N_2004,In_1582,In_539);
or U2005 (N_2005,In_954,In_1543);
or U2006 (N_2006,In_260,In_1087);
nor U2007 (N_2007,In_185,In_27);
nor U2008 (N_2008,In_680,In_228);
xor U2009 (N_2009,In_1418,In_1587);
nand U2010 (N_2010,In_136,In_196);
or U2011 (N_2011,In_1438,In_1638);
or U2012 (N_2012,In_236,In_1163);
nand U2013 (N_2013,In_976,In_1493);
or U2014 (N_2014,In_485,In_1926);
xnor U2015 (N_2015,In_1376,In_666);
and U2016 (N_2016,In_1862,In_1144);
xnor U2017 (N_2017,In_226,In_398);
or U2018 (N_2018,In_394,In_661);
nand U2019 (N_2019,In_367,In_740);
nor U2020 (N_2020,In_1085,In_1217);
xnor U2021 (N_2021,In_1859,In_1324);
and U2022 (N_2022,In_1072,In_323);
and U2023 (N_2023,In_650,In_281);
nand U2024 (N_2024,In_1395,In_1877);
nor U2025 (N_2025,In_689,In_1375);
nand U2026 (N_2026,In_134,In_212);
nand U2027 (N_2027,In_1381,In_558);
nand U2028 (N_2028,In_762,In_1864);
xor U2029 (N_2029,In_1716,In_1036);
or U2030 (N_2030,In_824,In_1973);
and U2031 (N_2031,In_1021,In_231);
nand U2032 (N_2032,In_1522,In_328);
nor U2033 (N_2033,In_1913,In_34);
and U2034 (N_2034,In_1630,In_909);
nand U2035 (N_2035,In_835,In_1050);
nand U2036 (N_2036,In_337,In_520);
nor U2037 (N_2037,In_1174,In_1240);
nor U2038 (N_2038,In_637,In_886);
or U2039 (N_2039,In_1060,In_629);
nor U2040 (N_2040,In_1516,In_1223);
xor U2041 (N_2041,In_327,In_1744);
and U2042 (N_2042,In_1115,In_1341);
or U2043 (N_2043,In_1279,In_1667);
nand U2044 (N_2044,In_883,In_805);
xor U2045 (N_2045,In_53,In_1516);
nor U2046 (N_2046,In_1990,In_1039);
nand U2047 (N_2047,In_697,In_736);
xor U2048 (N_2048,In_215,In_219);
and U2049 (N_2049,In_235,In_502);
nand U2050 (N_2050,In_485,In_415);
and U2051 (N_2051,In_1517,In_1560);
xor U2052 (N_2052,In_166,In_85);
or U2053 (N_2053,In_483,In_131);
or U2054 (N_2054,In_793,In_137);
and U2055 (N_2055,In_247,In_1586);
nor U2056 (N_2056,In_600,In_1716);
xor U2057 (N_2057,In_425,In_1438);
nor U2058 (N_2058,In_109,In_440);
nand U2059 (N_2059,In_684,In_1378);
or U2060 (N_2060,In_117,In_1178);
xor U2061 (N_2061,In_1451,In_152);
and U2062 (N_2062,In_1115,In_811);
nand U2063 (N_2063,In_1980,In_1067);
nand U2064 (N_2064,In_245,In_916);
xor U2065 (N_2065,In_909,In_44);
and U2066 (N_2066,In_801,In_711);
or U2067 (N_2067,In_798,In_1005);
and U2068 (N_2068,In_904,In_241);
nor U2069 (N_2069,In_1992,In_327);
and U2070 (N_2070,In_1669,In_1213);
and U2071 (N_2071,In_1561,In_1598);
xnor U2072 (N_2072,In_321,In_1670);
nor U2073 (N_2073,In_1218,In_244);
nor U2074 (N_2074,In_916,In_1775);
nor U2075 (N_2075,In_339,In_1907);
nand U2076 (N_2076,In_729,In_1908);
or U2077 (N_2077,In_905,In_899);
nor U2078 (N_2078,In_1785,In_90);
xor U2079 (N_2079,In_1689,In_493);
nor U2080 (N_2080,In_643,In_101);
or U2081 (N_2081,In_345,In_1393);
nor U2082 (N_2082,In_1705,In_548);
nand U2083 (N_2083,In_866,In_315);
xor U2084 (N_2084,In_103,In_1262);
xor U2085 (N_2085,In_162,In_1679);
and U2086 (N_2086,In_1701,In_1624);
and U2087 (N_2087,In_1675,In_1609);
and U2088 (N_2088,In_1777,In_41);
and U2089 (N_2089,In_1921,In_26);
xnor U2090 (N_2090,In_510,In_1434);
and U2091 (N_2091,In_319,In_1963);
and U2092 (N_2092,In_198,In_263);
xnor U2093 (N_2093,In_705,In_1017);
nand U2094 (N_2094,In_78,In_1044);
xor U2095 (N_2095,In_293,In_1550);
or U2096 (N_2096,In_41,In_1078);
nand U2097 (N_2097,In_209,In_138);
nor U2098 (N_2098,In_1505,In_520);
and U2099 (N_2099,In_1848,In_1287);
xnor U2100 (N_2100,In_1662,In_1677);
xnor U2101 (N_2101,In_78,In_1431);
xor U2102 (N_2102,In_1338,In_584);
nor U2103 (N_2103,In_846,In_1187);
or U2104 (N_2104,In_1281,In_759);
or U2105 (N_2105,In_259,In_761);
nand U2106 (N_2106,In_974,In_1064);
or U2107 (N_2107,In_1741,In_672);
and U2108 (N_2108,In_1871,In_1459);
nand U2109 (N_2109,In_999,In_1437);
or U2110 (N_2110,In_1050,In_1561);
or U2111 (N_2111,In_1962,In_1190);
xnor U2112 (N_2112,In_1685,In_1780);
and U2113 (N_2113,In_1649,In_421);
xor U2114 (N_2114,In_1572,In_987);
nand U2115 (N_2115,In_259,In_1239);
and U2116 (N_2116,In_693,In_666);
xor U2117 (N_2117,In_1363,In_683);
nand U2118 (N_2118,In_1314,In_749);
nor U2119 (N_2119,In_776,In_302);
or U2120 (N_2120,In_1416,In_49);
and U2121 (N_2121,In_1308,In_766);
and U2122 (N_2122,In_798,In_1452);
xnor U2123 (N_2123,In_1850,In_1778);
xor U2124 (N_2124,In_148,In_756);
nor U2125 (N_2125,In_1962,In_1608);
xor U2126 (N_2126,In_1800,In_738);
nor U2127 (N_2127,In_276,In_1886);
nand U2128 (N_2128,In_1028,In_1355);
xnor U2129 (N_2129,In_1351,In_355);
nor U2130 (N_2130,In_1841,In_1309);
nand U2131 (N_2131,In_488,In_444);
and U2132 (N_2132,In_459,In_66);
and U2133 (N_2133,In_1553,In_227);
or U2134 (N_2134,In_1723,In_1957);
nor U2135 (N_2135,In_1178,In_696);
nor U2136 (N_2136,In_1010,In_454);
xnor U2137 (N_2137,In_485,In_1252);
and U2138 (N_2138,In_1909,In_1451);
or U2139 (N_2139,In_285,In_782);
nor U2140 (N_2140,In_1455,In_1593);
nor U2141 (N_2141,In_656,In_1371);
xnor U2142 (N_2142,In_1367,In_170);
nor U2143 (N_2143,In_539,In_1472);
and U2144 (N_2144,In_926,In_1266);
or U2145 (N_2145,In_810,In_1345);
xnor U2146 (N_2146,In_133,In_1956);
or U2147 (N_2147,In_1955,In_1239);
nor U2148 (N_2148,In_430,In_152);
nor U2149 (N_2149,In_284,In_234);
nor U2150 (N_2150,In_1018,In_1396);
xnor U2151 (N_2151,In_1333,In_1112);
xnor U2152 (N_2152,In_1918,In_429);
nor U2153 (N_2153,In_620,In_1722);
xnor U2154 (N_2154,In_411,In_517);
or U2155 (N_2155,In_1753,In_1144);
nand U2156 (N_2156,In_271,In_1112);
and U2157 (N_2157,In_1025,In_288);
or U2158 (N_2158,In_1363,In_1689);
xor U2159 (N_2159,In_1965,In_971);
xnor U2160 (N_2160,In_1185,In_174);
and U2161 (N_2161,In_189,In_639);
nand U2162 (N_2162,In_6,In_754);
xor U2163 (N_2163,In_1383,In_1626);
xnor U2164 (N_2164,In_202,In_789);
nand U2165 (N_2165,In_573,In_1786);
and U2166 (N_2166,In_472,In_226);
nor U2167 (N_2167,In_904,In_1324);
nor U2168 (N_2168,In_1545,In_1480);
nand U2169 (N_2169,In_1536,In_920);
or U2170 (N_2170,In_169,In_1511);
xor U2171 (N_2171,In_1338,In_249);
or U2172 (N_2172,In_345,In_1737);
nand U2173 (N_2173,In_581,In_1938);
xnor U2174 (N_2174,In_1971,In_319);
or U2175 (N_2175,In_249,In_1509);
nor U2176 (N_2176,In_772,In_974);
and U2177 (N_2177,In_438,In_1428);
and U2178 (N_2178,In_1084,In_1879);
xnor U2179 (N_2179,In_1681,In_103);
or U2180 (N_2180,In_324,In_131);
and U2181 (N_2181,In_1526,In_1420);
and U2182 (N_2182,In_167,In_688);
nand U2183 (N_2183,In_1322,In_8);
xnor U2184 (N_2184,In_1480,In_653);
and U2185 (N_2185,In_86,In_1982);
nor U2186 (N_2186,In_858,In_1334);
xnor U2187 (N_2187,In_783,In_1763);
or U2188 (N_2188,In_1222,In_1649);
nand U2189 (N_2189,In_521,In_223);
xor U2190 (N_2190,In_1246,In_365);
xor U2191 (N_2191,In_628,In_373);
nand U2192 (N_2192,In_1196,In_1831);
and U2193 (N_2193,In_679,In_823);
nor U2194 (N_2194,In_1658,In_1890);
xnor U2195 (N_2195,In_588,In_1461);
nand U2196 (N_2196,In_185,In_742);
xnor U2197 (N_2197,In_141,In_1687);
xnor U2198 (N_2198,In_549,In_953);
xor U2199 (N_2199,In_1716,In_1474);
nand U2200 (N_2200,In_140,In_1217);
xnor U2201 (N_2201,In_1344,In_408);
nand U2202 (N_2202,In_842,In_113);
xor U2203 (N_2203,In_1366,In_540);
nor U2204 (N_2204,In_132,In_1259);
nor U2205 (N_2205,In_232,In_1271);
nor U2206 (N_2206,In_220,In_1970);
nor U2207 (N_2207,In_285,In_1725);
or U2208 (N_2208,In_1308,In_1885);
xnor U2209 (N_2209,In_509,In_1953);
xnor U2210 (N_2210,In_600,In_663);
or U2211 (N_2211,In_372,In_1454);
and U2212 (N_2212,In_759,In_184);
or U2213 (N_2213,In_920,In_19);
nor U2214 (N_2214,In_1097,In_438);
nor U2215 (N_2215,In_1529,In_24);
nor U2216 (N_2216,In_141,In_1360);
nor U2217 (N_2217,In_414,In_1547);
and U2218 (N_2218,In_1516,In_179);
xnor U2219 (N_2219,In_1307,In_115);
nand U2220 (N_2220,In_1677,In_450);
or U2221 (N_2221,In_425,In_1976);
nand U2222 (N_2222,In_1309,In_1685);
xnor U2223 (N_2223,In_1200,In_1834);
or U2224 (N_2224,In_920,In_60);
xor U2225 (N_2225,In_522,In_1451);
xnor U2226 (N_2226,In_32,In_1367);
and U2227 (N_2227,In_1181,In_1894);
nor U2228 (N_2228,In_1351,In_1672);
or U2229 (N_2229,In_1285,In_239);
xnor U2230 (N_2230,In_1573,In_1401);
xor U2231 (N_2231,In_596,In_650);
nor U2232 (N_2232,In_1835,In_1106);
and U2233 (N_2233,In_1790,In_58);
or U2234 (N_2234,In_1622,In_1112);
xor U2235 (N_2235,In_1571,In_448);
nand U2236 (N_2236,In_1769,In_303);
nand U2237 (N_2237,In_31,In_917);
nand U2238 (N_2238,In_1233,In_1383);
nor U2239 (N_2239,In_489,In_797);
nor U2240 (N_2240,In_630,In_5);
xnor U2241 (N_2241,In_1293,In_1278);
or U2242 (N_2242,In_1646,In_689);
and U2243 (N_2243,In_1440,In_1839);
nor U2244 (N_2244,In_1029,In_1424);
xor U2245 (N_2245,In_1864,In_135);
nand U2246 (N_2246,In_1938,In_1012);
nand U2247 (N_2247,In_936,In_266);
nor U2248 (N_2248,In_787,In_764);
and U2249 (N_2249,In_391,In_1582);
nor U2250 (N_2250,In_65,In_1313);
xnor U2251 (N_2251,In_989,In_1778);
nand U2252 (N_2252,In_1021,In_1870);
or U2253 (N_2253,In_1850,In_1955);
xnor U2254 (N_2254,In_1117,In_654);
xnor U2255 (N_2255,In_1098,In_1545);
and U2256 (N_2256,In_513,In_332);
or U2257 (N_2257,In_1255,In_1303);
xor U2258 (N_2258,In_1625,In_1573);
nand U2259 (N_2259,In_1135,In_1812);
and U2260 (N_2260,In_103,In_765);
xor U2261 (N_2261,In_1654,In_1514);
xor U2262 (N_2262,In_1310,In_91);
xor U2263 (N_2263,In_160,In_1281);
xnor U2264 (N_2264,In_416,In_898);
xor U2265 (N_2265,In_1369,In_996);
nor U2266 (N_2266,In_1313,In_1622);
or U2267 (N_2267,In_782,In_541);
and U2268 (N_2268,In_1549,In_1022);
xor U2269 (N_2269,In_229,In_1032);
nor U2270 (N_2270,In_1168,In_622);
or U2271 (N_2271,In_1449,In_130);
xor U2272 (N_2272,In_982,In_1414);
and U2273 (N_2273,In_721,In_478);
nor U2274 (N_2274,In_1930,In_166);
xnor U2275 (N_2275,In_1116,In_1582);
nand U2276 (N_2276,In_1092,In_1357);
nor U2277 (N_2277,In_848,In_1882);
xor U2278 (N_2278,In_490,In_1771);
xnor U2279 (N_2279,In_505,In_550);
nand U2280 (N_2280,In_1508,In_1114);
and U2281 (N_2281,In_329,In_0);
nand U2282 (N_2282,In_1381,In_162);
or U2283 (N_2283,In_1911,In_364);
xnor U2284 (N_2284,In_1676,In_366);
and U2285 (N_2285,In_214,In_262);
nand U2286 (N_2286,In_784,In_1219);
xnor U2287 (N_2287,In_373,In_525);
or U2288 (N_2288,In_757,In_1472);
and U2289 (N_2289,In_769,In_210);
xnor U2290 (N_2290,In_540,In_1329);
nand U2291 (N_2291,In_41,In_1260);
and U2292 (N_2292,In_1711,In_1197);
and U2293 (N_2293,In_1418,In_825);
or U2294 (N_2294,In_631,In_1443);
and U2295 (N_2295,In_736,In_1964);
xnor U2296 (N_2296,In_1479,In_1937);
nor U2297 (N_2297,In_1636,In_1734);
and U2298 (N_2298,In_83,In_369);
nor U2299 (N_2299,In_1778,In_1634);
or U2300 (N_2300,In_1993,In_539);
and U2301 (N_2301,In_1817,In_1845);
and U2302 (N_2302,In_1536,In_28);
nand U2303 (N_2303,In_1681,In_266);
and U2304 (N_2304,In_859,In_1324);
or U2305 (N_2305,In_595,In_1704);
xnor U2306 (N_2306,In_32,In_304);
nor U2307 (N_2307,In_1199,In_1958);
xor U2308 (N_2308,In_451,In_780);
and U2309 (N_2309,In_994,In_1997);
nand U2310 (N_2310,In_1026,In_1027);
or U2311 (N_2311,In_1585,In_1251);
and U2312 (N_2312,In_857,In_567);
or U2313 (N_2313,In_727,In_198);
and U2314 (N_2314,In_101,In_25);
nand U2315 (N_2315,In_1341,In_1117);
nand U2316 (N_2316,In_1119,In_1652);
nand U2317 (N_2317,In_795,In_862);
xor U2318 (N_2318,In_1480,In_1586);
and U2319 (N_2319,In_1537,In_899);
or U2320 (N_2320,In_1587,In_1530);
nor U2321 (N_2321,In_1990,In_1244);
nand U2322 (N_2322,In_1111,In_1130);
nand U2323 (N_2323,In_59,In_595);
xnor U2324 (N_2324,In_184,In_1864);
nor U2325 (N_2325,In_500,In_349);
xor U2326 (N_2326,In_1093,In_1279);
nand U2327 (N_2327,In_226,In_497);
or U2328 (N_2328,In_792,In_1887);
nor U2329 (N_2329,In_1350,In_1733);
and U2330 (N_2330,In_47,In_727);
or U2331 (N_2331,In_1279,In_1737);
or U2332 (N_2332,In_1607,In_200);
or U2333 (N_2333,In_932,In_1076);
xnor U2334 (N_2334,In_1634,In_646);
xor U2335 (N_2335,In_37,In_713);
nor U2336 (N_2336,In_1497,In_1749);
nand U2337 (N_2337,In_544,In_1457);
or U2338 (N_2338,In_1178,In_484);
nor U2339 (N_2339,In_1391,In_1788);
or U2340 (N_2340,In_1881,In_1208);
nor U2341 (N_2341,In_423,In_177);
or U2342 (N_2342,In_1902,In_463);
or U2343 (N_2343,In_90,In_788);
xor U2344 (N_2344,In_913,In_325);
nand U2345 (N_2345,In_575,In_1068);
nand U2346 (N_2346,In_357,In_805);
xor U2347 (N_2347,In_1957,In_1326);
xor U2348 (N_2348,In_380,In_198);
nor U2349 (N_2349,In_970,In_880);
and U2350 (N_2350,In_1775,In_1172);
xnor U2351 (N_2351,In_1111,In_1769);
nand U2352 (N_2352,In_1607,In_1876);
nor U2353 (N_2353,In_902,In_1425);
nand U2354 (N_2354,In_1689,In_525);
and U2355 (N_2355,In_763,In_1185);
or U2356 (N_2356,In_1248,In_1502);
xnor U2357 (N_2357,In_1496,In_1695);
nand U2358 (N_2358,In_1578,In_1912);
and U2359 (N_2359,In_1261,In_1952);
nor U2360 (N_2360,In_324,In_25);
xor U2361 (N_2361,In_1465,In_890);
nor U2362 (N_2362,In_1001,In_970);
nor U2363 (N_2363,In_1311,In_251);
nor U2364 (N_2364,In_342,In_1677);
and U2365 (N_2365,In_874,In_529);
nor U2366 (N_2366,In_149,In_1439);
nand U2367 (N_2367,In_610,In_1092);
xor U2368 (N_2368,In_1675,In_1657);
and U2369 (N_2369,In_1914,In_391);
or U2370 (N_2370,In_1468,In_100);
nor U2371 (N_2371,In_313,In_660);
nor U2372 (N_2372,In_1340,In_1669);
or U2373 (N_2373,In_351,In_181);
xnor U2374 (N_2374,In_97,In_599);
or U2375 (N_2375,In_1423,In_1683);
nand U2376 (N_2376,In_1566,In_374);
or U2377 (N_2377,In_1108,In_1694);
or U2378 (N_2378,In_943,In_1526);
xnor U2379 (N_2379,In_556,In_619);
and U2380 (N_2380,In_1219,In_1618);
nand U2381 (N_2381,In_27,In_272);
nand U2382 (N_2382,In_553,In_912);
xor U2383 (N_2383,In_1945,In_1226);
and U2384 (N_2384,In_1367,In_145);
and U2385 (N_2385,In_148,In_238);
nand U2386 (N_2386,In_540,In_1620);
and U2387 (N_2387,In_542,In_1978);
or U2388 (N_2388,In_499,In_30);
nor U2389 (N_2389,In_1981,In_1726);
and U2390 (N_2390,In_267,In_1829);
nand U2391 (N_2391,In_1444,In_1562);
nand U2392 (N_2392,In_222,In_1379);
xnor U2393 (N_2393,In_1846,In_58);
and U2394 (N_2394,In_1892,In_236);
or U2395 (N_2395,In_1571,In_1422);
nand U2396 (N_2396,In_1219,In_1361);
and U2397 (N_2397,In_1372,In_1941);
xor U2398 (N_2398,In_1974,In_1017);
nand U2399 (N_2399,In_1817,In_1519);
or U2400 (N_2400,In_1278,In_1621);
nand U2401 (N_2401,In_115,In_1040);
nor U2402 (N_2402,In_961,In_761);
xnor U2403 (N_2403,In_1171,In_1310);
and U2404 (N_2404,In_1211,In_874);
or U2405 (N_2405,In_1246,In_1020);
xnor U2406 (N_2406,In_834,In_286);
and U2407 (N_2407,In_727,In_1643);
nor U2408 (N_2408,In_1293,In_1663);
and U2409 (N_2409,In_15,In_69);
nor U2410 (N_2410,In_384,In_943);
xnor U2411 (N_2411,In_316,In_311);
xor U2412 (N_2412,In_576,In_341);
xor U2413 (N_2413,In_1305,In_539);
xor U2414 (N_2414,In_6,In_268);
nor U2415 (N_2415,In_1380,In_1582);
xnor U2416 (N_2416,In_35,In_89);
xnor U2417 (N_2417,In_1893,In_3);
nand U2418 (N_2418,In_220,In_1943);
and U2419 (N_2419,In_1710,In_1773);
nor U2420 (N_2420,In_1584,In_94);
xor U2421 (N_2421,In_1058,In_1575);
and U2422 (N_2422,In_1584,In_1913);
xor U2423 (N_2423,In_512,In_1846);
xor U2424 (N_2424,In_974,In_1438);
or U2425 (N_2425,In_1024,In_840);
xnor U2426 (N_2426,In_1840,In_1711);
xor U2427 (N_2427,In_850,In_1169);
and U2428 (N_2428,In_888,In_1695);
xor U2429 (N_2429,In_733,In_1843);
and U2430 (N_2430,In_1895,In_1807);
nand U2431 (N_2431,In_984,In_1930);
xor U2432 (N_2432,In_1589,In_243);
or U2433 (N_2433,In_223,In_905);
xor U2434 (N_2434,In_1912,In_1813);
or U2435 (N_2435,In_1340,In_1099);
xor U2436 (N_2436,In_167,In_1473);
nand U2437 (N_2437,In_1539,In_1179);
nand U2438 (N_2438,In_1749,In_819);
nor U2439 (N_2439,In_1827,In_92);
nand U2440 (N_2440,In_1404,In_1158);
nor U2441 (N_2441,In_948,In_1000);
nand U2442 (N_2442,In_831,In_636);
nor U2443 (N_2443,In_1179,In_1263);
xnor U2444 (N_2444,In_1044,In_1548);
nand U2445 (N_2445,In_1208,In_1395);
and U2446 (N_2446,In_1403,In_1078);
xnor U2447 (N_2447,In_1621,In_717);
or U2448 (N_2448,In_240,In_511);
xnor U2449 (N_2449,In_233,In_756);
nor U2450 (N_2450,In_1168,In_630);
or U2451 (N_2451,In_236,In_835);
and U2452 (N_2452,In_1337,In_167);
nand U2453 (N_2453,In_303,In_930);
or U2454 (N_2454,In_1463,In_1678);
or U2455 (N_2455,In_874,In_883);
or U2456 (N_2456,In_662,In_3);
or U2457 (N_2457,In_239,In_1185);
and U2458 (N_2458,In_1668,In_1079);
or U2459 (N_2459,In_1630,In_713);
or U2460 (N_2460,In_1090,In_1790);
and U2461 (N_2461,In_1350,In_1711);
nand U2462 (N_2462,In_1340,In_1835);
and U2463 (N_2463,In_852,In_391);
and U2464 (N_2464,In_903,In_916);
nor U2465 (N_2465,In_1074,In_1349);
or U2466 (N_2466,In_654,In_1407);
nor U2467 (N_2467,In_580,In_1747);
nor U2468 (N_2468,In_189,In_1229);
nand U2469 (N_2469,In_1112,In_194);
nand U2470 (N_2470,In_1490,In_1604);
and U2471 (N_2471,In_445,In_1728);
or U2472 (N_2472,In_392,In_1958);
and U2473 (N_2473,In_292,In_1667);
and U2474 (N_2474,In_206,In_1697);
or U2475 (N_2475,In_1748,In_927);
xnor U2476 (N_2476,In_1237,In_1769);
nand U2477 (N_2477,In_1855,In_252);
nor U2478 (N_2478,In_1966,In_866);
or U2479 (N_2479,In_1647,In_1675);
and U2480 (N_2480,In_988,In_249);
nand U2481 (N_2481,In_1996,In_969);
or U2482 (N_2482,In_274,In_188);
nand U2483 (N_2483,In_927,In_1681);
and U2484 (N_2484,In_1571,In_368);
nand U2485 (N_2485,In_1883,In_366);
nor U2486 (N_2486,In_1004,In_1105);
and U2487 (N_2487,In_1322,In_1225);
and U2488 (N_2488,In_751,In_244);
nor U2489 (N_2489,In_881,In_1154);
xor U2490 (N_2490,In_1396,In_1413);
or U2491 (N_2491,In_1345,In_1323);
nand U2492 (N_2492,In_808,In_1091);
nor U2493 (N_2493,In_1024,In_722);
and U2494 (N_2494,In_1546,In_172);
xor U2495 (N_2495,In_1710,In_47);
nand U2496 (N_2496,In_1139,In_208);
nor U2497 (N_2497,In_11,In_893);
nand U2498 (N_2498,In_1898,In_234);
nor U2499 (N_2499,In_659,In_1515);
nand U2500 (N_2500,In_446,In_835);
nor U2501 (N_2501,In_494,In_956);
xnor U2502 (N_2502,In_191,In_96);
xor U2503 (N_2503,In_978,In_972);
and U2504 (N_2504,In_611,In_200);
xor U2505 (N_2505,In_1971,In_1196);
xnor U2506 (N_2506,In_1299,In_1241);
and U2507 (N_2507,In_687,In_436);
xor U2508 (N_2508,In_1050,In_201);
or U2509 (N_2509,In_880,In_1532);
and U2510 (N_2510,In_250,In_1106);
xor U2511 (N_2511,In_53,In_1282);
or U2512 (N_2512,In_130,In_160);
nor U2513 (N_2513,In_624,In_52);
nand U2514 (N_2514,In_952,In_330);
and U2515 (N_2515,In_4,In_1838);
nor U2516 (N_2516,In_1625,In_1511);
or U2517 (N_2517,In_1675,In_1157);
xnor U2518 (N_2518,In_172,In_384);
and U2519 (N_2519,In_1210,In_1351);
and U2520 (N_2520,In_443,In_1332);
xnor U2521 (N_2521,In_961,In_1130);
xor U2522 (N_2522,In_1668,In_648);
xnor U2523 (N_2523,In_48,In_657);
and U2524 (N_2524,In_376,In_1223);
or U2525 (N_2525,In_1321,In_223);
nand U2526 (N_2526,In_968,In_1269);
xor U2527 (N_2527,In_286,In_1369);
xnor U2528 (N_2528,In_1534,In_1354);
xor U2529 (N_2529,In_1828,In_1059);
or U2530 (N_2530,In_1767,In_307);
nand U2531 (N_2531,In_1100,In_1146);
or U2532 (N_2532,In_295,In_1858);
nor U2533 (N_2533,In_1382,In_578);
xnor U2534 (N_2534,In_1255,In_179);
nand U2535 (N_2535,In_772,In_1287);
and U2536 (N_2536,In_480,In_1693);
xor U2537 (N_2537,In_1280,In_1555);
nand U2538 (N_2538,In_1924,In_466);
or U2539 (N_2539,In_660,In_46);
and U2540 (N_2540,In_1610,In_546);
or U2541 (N_2541,In_151,In_1953);
or U2542 (N_2542,In_1244,In_1001);
nand U2543 (N_2543,In_1871,In_243);
xor U2544 (N_2544,In_1739,In_1581);
or U2545 (N_2545,In_1377,In_111);
xor U2546 (N_2546,In_734,In_1234);
or U2547 (N_2547,In_1894,In_1658);
or U2548 (N_2548,In_893,In_1891);
nand U2549 (N_2549,In_36,In_1180);
and U2550 (N_2550,In_880,In_484);
or U2551 (N_2551,In_960,In_588);
nand U2552 (N_2552,In_9,In_540);
xnor U2553 (N_2553,In_198,In_1973);
and U2554 (N_2554,In_1803,In_612);
nor U2555 (N_2555,In_1234,In_170);
xnor U2556 (N_2556,In_24,In_1286);
and U2557 (N_2557,In_547,In_517);
xor U2558 (N_2558,In_316,In_258);
or U2559 (N_2559,In_1169,In_499);
and U2560 (N_2560,In_5,In_550);
or U2561 (N_2561,In_1784,In_1543);
xnor U2562 (N_2562,In_55,In_1173);
nor U2563 (N_2563,In_1762,In_767);
nand U2564 (N_2564,In_1421,In_421);
nor U2565 (N_2565,In_419,In_92);
nor U2566 (N_2566,In_816,In_86);
nor U2567 (N_2567,In_856,In_1413);
or U2568 (N_2568,In_536,In_666);
nor U2569 (N_2569,In_207,In_1283);
and U2570 (N_2570,In_1045,In_765);
or U2571 (N_2571,In_1987,In_655);
nor U2572 (N_2572,In_1180,In_1933);
and U2573 (N_2573,In_1907,In_744);
xor U2574 (N_2574,In_1581,In_1079);
nand U2575 (N_2575,In_705,In_1921);
nor U2576 (N_2576,In_1799,In_244);
and U2577 (N_2577,In_968,In_624);
or U2578 (N_2578,In_1169,In_1203);
and U2579 (N_2579,In_638,In_821);
and U2580 (N_2580,In_259,In_960);
nor U2581 (N_2581,In_1654,In_1141);
nand U2582 (N_2582,In_1816,In_1920);
or U2583 (N_2583,In_109,In_792);
xnor U2584 (N_2584,In_924,In_361);
and U2585 (N_2585,In_1239,In_16);
nand U2586 (N_2586,In_1145,In_1365);
or U2587 (N_2587,In_1926,In_1863);
xor U2588 (N_2588,In_991,In_1269);
nand U2589 (N_2589,In_1081,In_947);
nand U2590 (N_2590,In_1593,In_1414);
or U2591 (N_2591,In_766,In_273);
or U2592 (N_2592,In_591,In_1477);
xnor U2593 (N_2593,In_481,In_1494);
nand U2594 (N_2594,In_1501,In_1885);
xnor U2595 (N_2595,In_220,In_756);
nor U2596 (N_2596,In_1801,In_112);
nand U2597 (N_2597,In_1248,In_1019);
xor U2598 (N_2598,In_517,In_1566);
or U2599 (N_2599,In_499,In_967);
and U2600 (N_2600,In_817,In_97);
nor U2601 (N_2601,In_707,In_309);
and U2602 (N_2602,In_885,In_1495);
or U2603 (N_2603,In_1331,In_1487);
nand U2604 (N_2604,In_1723,In_1254);
and U2605 (N_2605,In_603,In_666);
or U2606 (N_2606,In_350,In_1296);
nand U2607 (N_2607,In_405,In_1027);
xor U2608 (N_2608,In_1219,In_1506);
nand U2609 (N_2609,In_305,In_169);
and U2610 (N_2610,In_40,In_1987);
nand U2611 (N_2611,In_409,In_728);
nand U2612 (N_2612,In_1649,In_1941);
nor U2613 (N_2613,In_1062,In_626);
xor U2614 (N_2614,In_1816,In_212);
and U2615 (N_2615,In_1957,In_97);
or U2616 (N_2616,In_1058,In_1119);
and U2617 (N_2617,In_360,In_1022);
nand U2618 (N_2618,In_296,In_1559);
nand U2619 (N_2619,In_1387,In_1008);
nor U2620 (N_2620,In_550,In_1191);
or U2621 (N_2621,In_1384,In_590);
nor U2622 (N_2622,In_348,In_1941);
nor U2623 (N_2623,In_565,In_140);
nand U2624 (N_2624,In_1450,In_1272);
nand U2625 (N_2625,In_1229,In_1858);
and U2626 (N_2626,In_1638,In_605);
and U2627 (N_2627,In_1295,In_744);
xnor U2628 (N_2628,In_1582,In_1710);
or U2629 (N_2629,In_1243,In_183);
or U2630 (N_2630,In_22,In_1502);
nor U2631 (N_2631,In_235,In_53);
nand U2632 (N_2632,In_1844,In_806);
nand U2633 (N_2633,In_318,In_867);
nor U2634 (N_2634,In_1589,In_5);
and U2635 (N_2635,In_1209,In_1755);
nor U2636 (N_2636,In_1301,In_1560);
nand U2637 (N_2637,In_1670,In_189);
xnor U2638 (N_2638,In_1984,In_1544);
nor U2639 (N_2639,In_1805,In_916);
nand U2640 (N_2640,In_1520,In_1791);
nor U2641 (N_2641,In_535,In_935);
or U2642 (N_2642,In_1107,In_1718);
nand U2643 (N_2643,In_148,In_1944);
or U2644 (N_2644,In_964,In_521);
and U2645 (N_2645,In_1819,In_747);
nand U2646 (N_2646,In_1644,In_1123);
xor U2647 (N_2647,In_208,In_32);
and U2648 (N_2648,In_1829,In_886);
nand U2649 (N_2649,In_226,In_360);
and U2650 (N_2650,In_1886,In_1158);
nor U2651 (N_2651,In_1650,In_878);
and U2652 (N_2652,In_1899,In_1100);
xnor U2653 (N_2653,In_1717,In_112);
xor U2654 (N_2654,In_1078,In_1590);
nand U2655 (N_2655,In_848,In_65);
xor U2656 (N_2656,In_1323,In_738);
or U2657 (N_2657,In_140,In_932);
nor U2658 (N_2658,In_75,In_1042);
and U2659 (N_2659,In_1620,In_1531);
xor U2660 (N_2660,In_1718,In_249);
or U2661 (N_2661,In_981,In_1727);
or U2662 (N_2662,In_1292,In_908);
nand U2663 (N_2663,In_1003,In_427);
nor U2664 (N_2664,In_1514,In_1067);
nor U2665 (N_2665,In_423,In_596);
nor U2666 (N_2666,In_1727,In_1651);
or U2667 (N_2667,In_1561,In_399);
xor U2668 (N_2668,In_1417,In_1779);
xnor U2669 (N_2669,In_1402,In_600);
and U2670 (N_2670,In_1407,In_420);
nand U2671 (N_2671,In_1670,In_1374);
nor U2672 (N_2672,In_510,In_1354);
or U2673 (N_2673,In_1625,In_7);
xor U2674 (N_2674,In_464,In_1039);
xor U2675 (N_2675,In_687,In_1070);
and U2676 (N_2676,In_1199,In_177);
and U2677 (N_2677,In_199,In_899);
nor U2678 (N_2678,In_92,In_588);
xnor U2679 (N_2679,In_764,In_102);
xnor U2680 (N_2680,In_569,In_1777);
nor U2681 (N_2681,In_217,In_1196);
and U2682 (N_2682,In_447,In_515);
nor U2683 (N_2683,In_1928,In_526);
and U2684 (N_2684,In_644,In_1619);
nor U2685 (N_2685,In_1501,In_1844);
xor U2686 (N_2686,In_1073,In_515);
and U2687 (N_2687,In_1400,In_963);
nor U2688 (N_2688,In_1596,In_666);
nor U2689 (N_2689,In_125,In_699);
nor U2690 (N_2690,In_129,In_1108);
or U2691 (N_2691,In_1733,In_1446);
nor U2692 (N_2692,In_1009,In_996);
or U2693 (N_2693,In_890,In_1998);
nand U2694 (N_2694,In_309,In_623);
nor U2695 (N_2695,In_1378,In_753);
and U2696 (N_2696,In_934,In_159);
nor U2697 (N_2697,In_1581,In_740);
nand U2698 (N_2698,In_637,In_432);
xnor U2699 (N_2699,In_1758,In_735);
and U2700 (N_2700,In_720,In_117);
nand U2701 (N_2701,In_753,In_1925);
xnor U2702 (N_2702,In_1216,In_370);
and U2703 (N_2703,In_713,In_402);
nand U2704 (N_2704,In_945,In_1989);
xnor U2705 (N_2705,In_1128,In_374);
xor U2706 (N_2706,In_114,In_261);
and U2707 (N_2707,In_1028,In_1998);
or U2708 (N_2708,In_844,In_889);
xor U2709 (N_2709,In_1077,In_368);
or U2710 (N_2710,In_1285,In_734);
and U2711 (N_2711,In_160,In_1453);
nor U2712 (N_2712,In_146,In_1470);
or U2713 (N_2713,In_171,In_210);
nand U2714 (N_2714,In_1262,In_1520);
xor U2715 (N_2715,In_653,In_1783);
nor U2716 (N_2716,In_266,In_1238);
or U2717 (N_2717,In_1295,In_716);
or U2718 (N_2718,In_1419,In_463);
or U2719 (N_2719,In_1089,In_1153);
nor U2720 (N_2720,In_716,In_1192);
or U2721 (N_2721,In_1630,In_1002);
nor U2722 (N_2722,In_1743,In_1642);
xor U2723 (N_2723,In_1797,In_742);
xnor U2724 (N_2724,In_699,In_847);
xor U2725 (N_2725,In_236,In_111);
xor U2726 (N_2726,In_1604,In_1891);
or U2727 (N_2727,In_1503,In_1326);
or U2728 (N_2728,In_1503,In_1802);
or U2729 (N_2729,In_279,In_181);
and U2730 (N_2730,In_1000,In_1122);
or U2731 (N_2731,In_1079,In_1854);
nand U2732 (N_2732,In_464,In_1323);
or U2733 (N_2733,In_848,In_183);
or U2734 (N_2734,In_1086,In_1825);
or U2735 (N_2735,In_1003,In_925);
xor U2736 (N_2736,In_1906,In_1025);
nor U2737 (N_2737,In_1212,In_584);
nor U2738 (N_2738,In_1717,In_1672);
xnor U2739 (N_2739,In_75,In_46);
or U2740 (N_2740,In_117,In_1937);
and U2741 (N_2741,In_371,In_268);
or U2742 (N_2742,In_522,In_1033);
nand U2743 (N_2743,In_677,In_1126);
xnor U2744 (N_2744,In_1921,In_736);
or U2745 (N_2745,In_543,In_1124);
nand U2746 (N_2746,In_1701,In_1904);
or U2747 (N_2747,In_1520,In_1959);
xor U2748 (N_2748,In_1830,In_1900);
nor U2749 (N_2749,In_345,In_606);
xnor U2750 (N_2750,In_622,In_1561);
nand U2751 (N_2751,In_1010,In_1685);
nor U2752 (N_2752,In_882,In_99);
nand U2753 (N_2753,In_910,In_1508);
or U2754 (N_2754,In_571,In_1007);
and U2755 (N_2755,In_1172,In_1965);
nand U2756 (N_2756,In_1264,In_232);
nor U2757 (N_2757,In_1485,In_305);
xnor U2758 (N_2758,In_1335,In_311);
xor U2759 (N_2759,In_321,In_678);
xor U2760 (N_2760,In_1637,In_132);
nand U2761 (N_2761,In_1527,In_1359);
and U2762 (N_2762,In_595,In_559);
or U2763 (N_2763,In_943,In_403);
xor U2764 (N_2764,In_1658,In_531);
nor U2765 (N_2765,In_697,In_1479);
and U2766 (N_2766,In_1038,In_1774);
and U2767 (N_2767,In_680,In_1199);
nor U2768 (N_2768,In_1811,In_281);
nand U2769 (N_2769,In_151,In_855);
and U2770 (N_2770,In_85,In_1216);
and U2771 (N_2771,In_367,In_811);
xnor U2772 (N_2772,In_1581,In_1790);
xnor U2773 (N_2773,In_939,In_787);
or U2774 (N_2774,In_85,In_737);
and U2775 (N_2775,In_1260,In_381);
nand U2776 (N_2776,In_1533,In_1420);
xor U2777 (N_2777,In_547,In_449);
nor U2778 (N_2778,In_1952,In_1933);
or U2779 (N_2779,In_1498,In_1445);
or U2780 (N_2780,In_735,In_990);
xor U2781 (N_2781,In_399,In_1785);
nor U2782 (N_2782,In_1852,In_1343);
xnor U2783 (N_2783,In_1372,In_1931);
xnor U2784 (N_2784,In_17,In_105);
or U2785 (N_2785,In_824,In_1767);
xnor U2786 (N_2786,In_152,In_1308);
xnor U2787 (N_2787,In_705,In_1146);
nor U2788 (N_2788,In_1075,In_1905);
xnor U2789 (N_2789,In_23,In_215);
nand U2790 (N_2790,In_766,In_122);
nand U2791 (N_2791,In_666,In_239);
nand U2792 (N_2792,In_555,In_1879);
and U2793 (N_2793,In_363,In_1097);
xnor U2794 (N_2794,In_604,In_195);
and U2795 (N_2795,In_1592,In_1376);
nand U2796 (N_2796,In_1011,In_830);
nor U2797 (N_2797,In_232,In_862);
or U2798 (N_2798,In_631,In_592);
xor U2799 (N_2799,In_1307,In_1474);
and U2800 (N_2800,In_138,In_914);
nand U2801 (N_2801,In_334,In_1093);
xnor U2802 (N_2802,In_337,In_823);
xor U2803 (N_2803,In_1352,In_393);
nand U2804 (N_2804,In_1970,In_625);
nand U2805 (N_2805,In_601,In_1339);
or U2806 (N_2806,In_1413,In_1524);
xor U2807 (N_2807,In_8,In_1294);
and U2808 (N_2808,In_555,In_1526);
nor U2809 (N_2809,In_1861,In_859);
or U2810 (N_2810,In_1889,In_734);
nand U2811 (N_2811,In_523,In_476);
nand U2812 (N_2812,In_765,In_1531);
xnor U2813 (N_2813,In_1716,In_1165);
nand U2814 (N_2814,In_483,In_1672);
xor U2815 (N_2815,In_1625,In_613);
nand U2816 (N_2816,In_1295,In_1247);
or U2817 (N_2817,In_16,In_541);
nand U2818 (N_2818,In_810,In_1696);
nor U2819 (N_2819,In_1899,In_844);
nand U2820 (N_2820,In_769,In_1266);
or U2821 (N_2821,In_65,In_706);
xor U2822 (N_2822,In_1014,In_1194);
or U2823 (N_2823,In_1206,In_155);
and U2824 (N_2824,In_1158,In_442);
or U2825 (N_2825,In_587,In_1403);
nor U2826 (N_2826,In_63,In_744);
or U2827 (N_2827,In_1236,In_1733);
or U2828 (N_2828,In_714,In_992);
nand U2829 (N_2829,In_711,In_770);
nand U2830 (N_2830,In_394,In_813);
and U2831 (N_2831,In_744,In_1112);
and U2832 (N_2832,In_270,In_1669);
xor U2833 (N_2833,In_1055,In_1336);
nand U2834 (N_2834,In_310,In_657);
nand U2835 (N_2835,In_1762,In_802);
nor U2836 (N_2836,In_1485,In_542);
xnor U2837 (N_2837,In_1619,In_1488);
or U2838 (N_2838,In_1279,In_161);
or U2839 (N_2839,In_1011,In_1795);
or U2840 (N_2840,In_1964,In_1798);
and U2841 (N_2841,In_1757,In_400);
and U2842 (N_2842,In_1742,In_468);
xnor U2843 (N_2843,In_1834,In_1693);
xnor U2844 (N_2844,In_730,In_758);
and U2845 (N_2845,In_107,In_137);
and U2846 (N_2846,In_1768,In_1056);
xnor U2847 (N_2847,In_1321,In_947);
nand U2848 (N_2848,In_751,In_1052);
and U2849 (N_2849,In_700,In_1079);
or U2850 (N_2850,In_1636,In_861);
or U2851 (N_2851,In_1072,In_1096);
nand U2852 (N_2852,In_1301,In_640);
or U2853 (N_2853,In_475,In_1150);
nor U2854 (N_2854,In_362,In_1950);
nor U2855 (N_2855,In_1453,In_1561);
and U2856 (N_2856,In_405,In_95);
nor U2857 (N_2857,In_827,In_1515);
nor U2858 (N_2858,In_296,In_1192);
nand U2859 (N_2859,In_371,In_1359);
or U2860 (N_2860,In_1633,In_287);
and U2861 (N_2861,In_641,In_1192);
and U2862 (N_2862,In_344,In_219);
nand U2863 (N_2863,In_592,In_1349);
and U2864 (N_2864,In_940,In_809);
nand U2865 (N_2865,In_844,In_1077);
xor U2866 (N_2866,In_1508,In_333);
nor U2867 (N_2867,In_174,In_244);
nand U2868 (N_2868,In_939,In_1452);
or U2869 (N_2869,In_788,In_1019);
or U2870 (N_2870,In_701,In_1692);
nor U2871 (N_2871,In_1001,In_666);
xor U2872 (N_2872,In_1124,In_1633);
or U2873 (N_2873,In_72,In_1869);
nand U2874 (N_2874,In_990,In_598);
and U2875 (N_2875,In_1133,In_1372);
nand U2876 (N_2876,In_144,In_638);
nand U2877 (N_2877,In_1373,In_1231);
and U2878 (N_2878,In_561,In_76);
xor U2879 (N_2879,In_1959,In_1773);
or U2880 (N_2880,In_991,In_1416);
xor U2881 (N_2881,In_1209,In_164);
and U2882 (N_2882,In_1570,In_922);
or U2883 (N_2883,In_1601,In_359);
nor U2884 (N_2884,In_1091,In_1725);
or U2885 (N_2885,In_1981,In_1303);
xor U2886 (N_2886,In_304,In_1582);
or U2887 (N_2887,In_94,In_140);
and U2888 (N_2888,In_213,In_451);
xnor U2889 (N_2889,In_542,In_1036);
and U2890 (N_2890,In_1826,In_1601);
nor U2891 (N_2891,In_1616,In_1550);
xnor U2892 (N_2892,In_297,In_1827);
nand U2893 (N_2893,In_1578,In_418);
nor U2894 (N_2894,In_1930,In_706);
nor U2895 (N_2895,In_1203,In_1759);
xnor U2896 (N_2896,In_1955,In_934);
or U2897 (N_2897,In_848,In_57);
nand U2898 (N_2898,In_918,In_1229);
nor U2899 (N_2899,In_578,In_146);
and U2900 (N_2900,In_1179,In_682);
and U2901 (N_2901,In_361,In_772);
nor U2902 (N_2902,In_982,In_679);
nand U2903 (N_2903,In_712,In_1374);
xnor U2904 (N_2904,In_45,In_1847);
nor U2905 (N_2905,In_368,In_355);
xor U2906 (N_2906,In_915,In_980);
nor U2907 (N_2907,In_1189,In_1429);
and U2908 (N_2908,In_1410,In_213);
xnor U2909 (N_2909,In_1909,In_1002);
nand U2910 (N_2910,In_1841,In_1663);
and U2911 (N_2911,In_164,In_1670);
xnor U2912 (N_2912,In_1503,In_110);
and U2913 (N_2913,In_301,In_533);
nand U2914 (N_2914,In_1695,In_1063);
xor U2915 (N_2915,In_461,In_1610);
nor U2916 (N_2916,In_818,In_253);
nor U2917 (N_2917,In_761,In_1279);
nand U2918 (N_2918,In_9,In_1341);
nor U2919 (N_2919,In_1074,In_1890);
and U2920 (N_2920,In_1061,In_1248);
or U2921 (N_2921,In_675,In_818);
or U2922 (N_2922,In_1579,In_1006);
nand U2923 (N_2923,In_1892,In_158);
and U2924 (N_2924,In_856,In_323);
nor U2925 (N_2925,In_1007,In_1090);
nand U2926 (N_2926,In_12,In_1373);
and U2927 (N_2927,In_1550,In_577);
or U2928 (N_2928,In_1065,In_1489);
and U2929 (N_2929,In_602,In_811);
nor U2930 (N_2930,In_114,In_644);
nor U2931 (N_2931,In_1154,In_1898);
and U2932 (N_2932,In_1256,In_1115);
xor U2933 (N_2933,In_1845,In_1061);
or U2934 (N_2934,In_1991,In_1037);
and U2935 (N_2935,In_1784,In_85);
or U2936 (N_2936,In_832,In_1142);
nand U2937 (N_2937,In_568,In_1398);
nor U2938 (N_2938,In_1005,In_1648);
and U2939 (N_2939,In_387,In_1322);
nand U2940 (N_2940,In_326,In_908);
nand U2941 (N_2941,In_151,In_1511);
xnor U2942 (N_2942,In_675,In_1340);
and U2943 (N_2943,In_487,In_272);
or U2944 (N_2944,In_78,In_1722);
xnor U2945 (N_2945,In_1755,In_658);
and U2946 (N_2946,In_1045,In_744);
xor U2947 (N_2947,In_556,In_942);
nor U2948 (N_2948,In_101,In_1039);
and U2949 (N_2949,In_693,In_903);
nor U2950 (N_2950,In_331,In_1540);
nor U2951 (N_2951,In_487,In_248);
or U2952 (N_2952,In_379,In_1543);
nand U2953 (N_2953,In_766,In_640);
or U2954 (N_2954,In_803,In_420);
nand U2955 (N_2955,In_958,In_1856);
or U2956 (N_2956,In_933,In_1162);
nor U2957 (N_2957,In_1609,In_64);
nand U2958 (N_2958,In_1644,In_320);
nand U2959 (N_2959,In_1585,In_443);
xnor U2960 (N_2960,In_467,In_1530);
nor U2961 (N_2961,In_34,In_869);
xor U2962 (N_2962,In_110,In_521);
nor U2963 (N_2963,In_1156,In_566);
nor U2964 (N_2964,In_692,In_1313);
or U2965 (N_2965,In_110,In_222);
and U2966 (N_2966,In_1120,In_1650);
or U2967 (N_2967,In_523,In_360);
or U2968 (N_2968,In_1044,In_1028);
or U2969 (N_2969,In_1806,In_158);
nor U2970 (N_2970,In_233,In_2);
nor U2971 (N_2971,In_368,In_1884);
nand U2972 (N_2972,In_1638,In_1003);
and U2973 (N_2973,In_948,In_668);
xnor U2974 (N_2974,In_42,In_997);
and U2975 (N_2975,In_244,In_42);
xor U2976 (N_2976,In_1535,In_156);
and U2977 (N_2977,In_1651,In_966);
and U2978 (N_2978,In_768,In_1193);
and U2979 (N_2979,In_400,In_1059);
and U2980 (N_2980,In_732,In_491);
nand U2981 (N_2981,In_1483,In_1743);
or U2982 (N_2982,In_1465,In_918);
xnor U2983 (N_2983,In_902,In_371);
or U2984 (N_2984,In_561,In_479);
xnor U2985 (N_2985,In_1817,In_658);
or U2986 (N_2986,In_1273,In_1122);
xnor U2987 (N_2987,In_1331,In_1551);
nor U2988 (N_2988,In_104,In_673);
and U2989 (N_2989,In_845,In_1187);
nor U2990 (N_2990,In_196,In_1298);
nand U2991 (N_2991,In_1552,In_1818);
xor U2992 (N_2992,In_1411,In_1294);
xor U2993 (N_2993,In_784,In_306);
and U2994 (N_2994,In_1621,In_876);
and U2995 (N_2995,In_884,In_920);
and U2996 (N_2996,In_80,In_1424);
or U2997 (N_2997,In_1867,In_647);
xnor U2998 (N_2998,In_82,In_1828);
nor U2999 (N_2999,In_1259,In_926);
nand U3000 (N_3000,In_548,In_631);
nor U3001 (N_3001,In_1307,In_1643);
nor U3002 (N_3002,In_227,In_1412);
nand U3003 (N_3003,In_1847,In_1892);
nor U3004 (N_3004,In_908,In_915);
or U3005 (N_3005,In_278,In_248);
or U3006 (N_3006,In_1943,In_612);
nor U3007 (N_3007,In_788,In_1731);
nand U3008 (N_3008,In_323,In_523);
and U3009 (N_3009,In_1693,In_1901);
nor U3010 (N_3010,In_651,In_1571);
nand U3011 (N_3011,In_887,In_731);
and U3012 (N_3012,In_513,In_981);
and U3013 (N_3013,In_1456,In_1024);
nor U3014 (N_3014,In_26,In_1928);
nor U3015 (N_3015,In_130,In_271);
and U3016 (N_3016,In_706,In_174);
or U3017 (N_3017,In_1722,In_331);
or U3018 (N_3018,In_67,In_1289);
nand U3019 (N_3019,In_1146,In_778);
nand U3020 (N_3020,In_910,In_1525);
nor U3021 (N_3021,In_393,In_1430);
nand U3022 (N_3022,In_1691,In_1360);
and U3023 (N_3023,In_1571,In_92);
or U3024 (N_3024,In_901,In_1366);
xor U3025 (N_3025,In_1803,In_401);
and U3026 (N_3026,In_500,In_71);
xnor U3027 (N_3027,In_1671,In_325);
and U3028 (N_3028,In_787,In_90);
nand U3029 (N_3029,In_1283,In_586);
or U3030 (N_3030,In_648,In_1200);
xnor U3031 (N_3031,In_1386,In_1832);
nor U3032 (N_3032,In_65,In_1603);
xnor U3033 (N_3033,In_1689,In_1315);
xor U3034 (N_3034,In_18,In_1723);
and U3035 (N_3035,In_1392,In_1800);
xor U3036 (N_3036,In_1399,In_1216);
and U3037 (N_3037,In_1478,In_1286);
nand U3038 (N_3038,In_258,In_1895);
xor U3039 (N_3039,In_1070,In_1402);
xor U3040 (N_3040,In_819,In_1840);
or U3041 (N_3041,In_1413,In_506);
nand U3042 (N_3042,In_1703,In_1013);
nor U3043 (N_3043,In_570,In_1754);
and U3044 (N_3044,In_1000,In_558);
nand U3045 (N_3045,In_1855,In_1906);
nor U3046 (N_3046,In_1577,In_1931);
nor U3047 (N_3047,In_23,In_1676);
xor U3048 (N_3048,In_993,In_1830);
nand U3049 (N_3049,In_1277,In_1746);
nand U3050 (N_3050,In_1581,In_250);
and U3051 (N_3051,In_1003,In_1441);
nand U3052 (N_3052,In_1072,In_1835);
nor U3053 (N_3053,In_920,In_1226);
nor U3054 (N_3054,In_1204,In_1106);
nor U3055 (N_3055,In_827,In_218);
and U3056 (N_3056,In_1406,In_601);
xnor U3057 (N_3057,In_549,In_1927);
and U3058 (N_3058,In_258,In_1989);
xor U3059 (N_3059,In_689,In_886);
nor U3060 (N_3060,In_1980,In_1455);
and U3061 (N_3061,In_222,In_505);
nor U3062 (N_3062,In_756,In_1471);
xor U3063 (N_3063,In_1409,In_1167);
or U3064 (N_3064,In_1491,In_358);
and U3065 (N_3065,In_230,In_623);
or U3066 (N_3066,In_1465,In_289);
nor U3067 (N_3067,In_275,In_609);
nor U3068 (N_3068,In_1243,In_1049);
xnor U3069 (N_3069,In_1845,In_1515);
xnor U3070 (N_3070,In_1543,In_1867);
xor U3071 (N_3071,In_115,In_1695);
xnor U3072 (N_3072,In_1465,In_1053);
nor U3073 (N_3073,In_1564,In_68);
xor U3074 (N_3074,In_850,In_322);
xnor U3075 (N_3075,In_1233,In_1457);
xnor U3076 (N_3076,In_801,In_926);
nand U3077 (N_3077,In_816,In_1046);
nand U3078 (N_3078,In_844,In_395);
or U3079 (N_3079,In_1299,In_159);
nor U3080 (N_3080,In_67,In_1224);
and U3081 (N_3081,In_1713,In_247);
or U3082 (N_3082,In_1670,In_939);
and U3083 (N_3083,In_202,In_234);
xor U3084 (N_3084,In_230,In_1023);
or U3085 (N_3085,In_409,In_1531);
nor U3086 (N_3086,In_917,In_868);
and U3087 (N_3087,In_847,In_1058);
nor U3088 (N_3088,In_722,In_1657);
and U3089 (N_3089,In_864,In_1672);
or U3090 (N_3090,In_278,In_801);
or U3091 (N_3091,In_286,In_1753);
or U3092 (N_3092,In_652,In_1874);
nand U3093 (N_3093,In_1687,In_1627);
nand U3094 (N_3094,In_580,In_706);
nor U3095 (N_3095,In_173,In_446);
nor U3096 (N_3096,In_1724,In_45);
and U3097 (N_3097,In_117,In_890);
or U3098 (N_3098,In_899,In_1275);
nand U3099 (N_3099,In_1628,In_490);
xnor U3100 (N_3100,In_1716,In_45);
and U3101 (N_3101,In_1604,In_389);
nand U3102 (N_3102,In_766,In_1135);
or U3103 (N_3103,In_949,In_1273);
xnor U3104 (N_3104,In_778,In_296);
nand U3105 (N_3105,In_474,In_646);
nand U3106 (N_3106,In_1862,In_1544);
or U3107 (N_3107,In_438,In_403);
or U3108 (N_3108,In_1334,In_1820);
and U3109 (N_3109,In_1184,In_249);
xnor U3110 (N_3110,In_1020,In_997);
xor U3111 (N_3111,In_1894,In_1013);
or U3112 (N_3112,In_1044,In_869);
or U3113 (N_3113,In_896,In_1662);
or U3114 (N_3114,In_164,In_1015);
xnor U3115 (N_3115,In_1146,In_1720);
or U3116 (N_3116,In_1839,In_721);
nor U3117 (N_3117,In_1490,In_592);
nand U3118 (N_3118,In_59,In_526);
or U3119 (N_3119,In_833,In_308);
or U3120 (N_3120,In_985,In_1266);
nor U3121 (N_3121,In_741,In_445);
and U3122 (N_3122,In_821,In_567);
nand U3123 (N_3123,In_123,In_344);
nor U3124 (N_3124,In_1148,In_993);
and U3125 (N_3125,In_1814,In_1685);
nor U3126 (N_3126,In_185,In_702);
nor U3127 (N_3127,In_1525,In_1917);
nor U3128 (N_3128,In_627,In_1501);
or U3129 (N_3129,In_917,In_411);
and U3130 (N_3130,In_942,In_851);
nor U3131 (N_3131,In_599,In_589);
or U3132 (N_3132,In_859,In_1278);
or U3133 (N_3133,In_230,In_1989);
xor U3134 (N_3134,In_455,In_604);
nand U3135 (N_3135,In_1289,In_140);
and U3136 (N_3136,In_682,In_513);
xnor U3137 (N_3137,In_917,In_1258);
nor U3138 (N_3138,In_681,In_1978);
nor U3139 (N_3139,In_278,In_81);
and U3140 (N_3140,In_1222,In_1763);
nand U3141 (N_3141,In_1884,In_1504);
nand U3142 (N_3142,In_1363,In_538);
nor U3143 (N_3143,In_1303,In_264);
or U3144 (N_3144,In_1195,In_796);
xor U3145 (N_3145,In_1196,In_1885);
nand U3146 (N_3146,In_758,In_760);
and U3147 (N_3147,In_1921,In_8);
and U3148 (N_3148,In_1262,In_287);
nand U3149 (N_3149,In_706,In_1387);
nand U3150 (N_3150,In_1343,In_991);
or U3151 (N_3151,In_1659,In_89);
nand U3152 (N_3152,In_715,In_1767);
nand U3153 (N_3153,In_1444,In_1800);
or U3154 (N_3154,In_1659,In_348);
xor U3155 (N_3155,In_433,In_777);
nor U3156 (N_3156,In_1245,In_1754);
or U3157 (N_3157,In_1500,In_1357);
nor U3158 (N_3158,In_943,In_937);
nor U3159 (N_3159,In_1369,In_1515);
or U3160 (N_3160,In_1959,In_1329);
xor U3161 (N_3161,In_210,In_442);
and U3162 (N_3162,In_607,In_1626);
or U3163 (N_3163,In_1778,In_1953);
or U3164 (N_3164,In_899,In_362);
nand U3165 (N_3165,In_1435,In_561);
and U3166 (N_3166,In_867,In_910);
and U3167 (N_3167,In_1573,In_955);
xnor U3168 (N_3168,In_829,In_216);
xor U3169 (N_3169,In_202,In_1147);
and U3170 (N_3170,In_107,In_1677);
nor U3171 (N_3171,In_840,In_1805);
xnor U3172 (N_3172,In_1524,In_1908);
nand U3173 (N_3173,In_734,In_4);
nand U3174 (N_3174,In_1125,In_70);
xor U3175 (N_3175,In_1364,In_1705);
and U3176 (N_3176,In_569,In_698);
nor U3177 (N_3177,In_731,In_929);
or U3178 (N_3178,In_1038,In_1349);
nand U3179 (N_3179,In_1292,In_1477);
and U3180 (N_3180,In_689,In_533);
nand U3181 (N_3181,In_627,In_46);
nand U3182 (N_3182,In_1421,In_706);
or U3183 (N_3183,In_1816,In_117);
and U3184 (N_3184,In_1345,In_1723);
or U3185 (N_3185,In_774,In_51);
nand U3186 (N_3186,In_1080,In_375);
nor U3187 (N_3187,In_768,In_575);
xnor U3188 (N_3188,In_317,In_1620);
or U3189 (N_3189,In_163,In_1493);
nand U3190 (N_3190,In_710,In_1218);
xnor U3191 (N_3191,In_848,In_1789);
nor U3192 (N_3192,In_9,In_1796);
and U3193 (N_3193,In_126,In_1815);
and U3194 (N_3194,In_1249,In_1123);
nor U3195 (N_3195,In_252,In_1253);
and U3196 (N_3196,In_1838,In_1244);
xor U3197 (N_3197,In_1520,In_629);
or U3198 (N_3198,In_1385,In_1677);
nor U3199 (N_3199,In_133,In_479);
and U3200 (N_3200,In_1932,In_639);
xnor U3201 (N_3201,In_1843,In_1858);
or U3202 (N_3202,In_541,In_1629);
nand U3203 (N_3203,In_312,In_1281);
nand U3204 (N_3204,In_1612,In_1256);
nand U3205 (N_3205,In_1721,In_367);
or U3206 (N_3206,In_234,In_1451);
and U3207 (N_3207,In_1561,In_1906);
xnor U3208 (N_3208,In_336,In_387);
and U3209 (N_3209,In_1856,In_533);
or U3210 (N_3210,In_394,In_1676);
nor U3211 (N_3211,In_1941,In_405);
nand U3212 (N_3212,In_745,In_1338);
xnor U3213 (N_3213,In_1520,In_1864);
or U3214 (N_3214,In_723,In_582);
nor U3215 (N_3215,In_1761,In_312);
nand U3216 (N_3216,In_1298,In_791);
nor U3217 (N_3217,In_1795,In_818);
and U3218 (N_3218,In_613,In_1312);
and U3219 (N_3219,In_1447,In_261);
and U3220 (N_3220,In_1191,In_695);
nand U3221 (N_3221,In_549,In_1683);
nand U3222 (N_3222,In_1651,In_879);
and U3223 (N_3223,In_63,In_1934);
and U3224 (N_3224,In_1711,In_780);
nand U3225 (N_3225,In_1256,In_516);
nand U3226 (N_3226,In_781,In_58);
nor U3227 (N_3227,In_1466,In_1390);
nor U3228 (N_3228,In_1792,In_1504);
or U3229 (N_3229,In_1337,In_554);
and U3230 (N_3230,In_489,In_761);
nor U3231 (N_3231,In_1240,In_431);
or U3232 (N_3232,In_323,In_1813);
nand U3233 (N_3233,In_488,In_1152);
xnor U3234 (N_3234,In_1838,In_910);
nand U3235 (N_3235,In_1909,In_1275);
or U3236 (N_3236,In_1570,In_1925);
xnor U3237 (N_3237,In_304,In_60);
nor U3238 (N_3238,In_418,In_568);
and U3239 (N_3239,In_1007,In_1103);
xor U3240 (N_3240,In_1759,In_1945);
and U3241 (N_3241,In_1515,In_252);
and U3242 (N_3242,In_1453,In_1102);
nor U3243 (N_3243,In_1121,In_1749);
nand U3244 (N_3244,In_1420,In_1238);
nand U3245 (N_3245,In_1503,In_1978);
or U3246 (N_3246,In_1372,In_973);
xnor U3247 (N_3247,In_456,In_1965);
and U3248 (N_3248,In_1039,In_916);
and U3249 (N_3249,In_408,In_467);
nand U3250 (N_3250,In_195,In_1982);
and U3251 (N_3251,In_1718,In_1300);
nand U3252 (N_3252,In_1297,In_1857);
or U3253 (N_3253,In_659,In_324);
nand U3254 (N_3254,In_211,In_918);
xnor U3255 (N_3255,In_892,In_1020);
or U3256 (N_3256,In_732,In_207);
nor U3257 (N_3257,In_1840,In_796);
nand U3258 (N_3258,In_1166,In_1176);
or U3259 (N_3259,In_418,In_1324);
xor U3260 (N_3260,In_1012,In_1142);
and U3261 (N_3261,In_419,In_1636);
nand U3262 (N_3262,In_41,In_983);
and U3263 (N_3263,In_1774,In_1119);
or U3264 (N_3264,In_124,In_1380);
or U3265 (N_3265,In_1266,In_324);
xor U3266 (N_3266,In_664,In_920);
or U3267 (N_3267,In_881,In_98);
or U3268 (N_3268,In_16,In_1575);
nor U3269 (N_3269,In_1576,In_1046);
and U3270 (N_3270,In_1231,In_248);
and U3271 (N_3271,In_261,In_1876);
and U3272 (N_3272,In_1147,In_1903);
nor U3273 (N_3273,In_641,In_666);
or U3274 (N_3274,In_312,In_1907);
or U3275 (N_3275,In_1248,In_671);
nor U3276 (N_3276,In_103,In_519);
xnor U3277 (N_3277,In_1366,In_546);
nor U3278 (N_3278,In_1081,In_1918);
and U3279 (N_3279,In_1640,In_1396);
xor U3280 (N_3280,In_441,In_1954);
xnor U3281 (N_3281,In_203,In_1544);
xnor U3282 (N_3282,In_628,In_1967);
nand U3283 (N_3283,In_584,In_485);
and U3284 (N_3284,In_288,In_153);
and U3285 (N_3285,In_142,In_577);
or U3286 (N_3286,In_1134,In_795);
and U3287 (N_3287,In_1048,In_1152);
and U3288 (N_3288,In_307,In_733);
nor U3289 (N_3289,In_1055,In_1642);
nand U3290 (N_3290,In_1888,In_754);
nor U3291 (N_3291,In_1849,In_733);
xor U3292 (N_3292,In_706,In_78);
nand U3293 (N_3293,In_596,In_85);
nand U3294 (N_3294,In_1227,In_1952);
nor U3295 (N_3295,In_897,In_1667);
and U3296 (N_3296,In_427,In_718);
or U3297 (N_3297,In_711,In_203);
or U3298 (N_3298,In_1497,In_1847);
and U3299 (N_3299,In_610,In_1716);
or U3300 (N_3300,In_1393,In_896);
xnor U3301 (N_3301,In_1138,In_199);
nor U3302 (N_3302,In_1598,In_606);
xnor U3303 (N_3303,In_1039,In_1240);
and U3304 (N_3304,In_936,In_1739);
or U3305 (N_3305,In_1925,In_522);
and U3306 (N_3306,In_496,In_122);
xnor U3307 (N_3307,In_1777,In_635);
nand U3308 (N_3308,In_1174,In_229);
xnor U3309 (N_3309,In_1983,In_215);
and U3310 (N_3310,In_1263,In_1707);
nand U3311 (N_3311,In_1832,In_1874);
and U3312 (N_3312,In_1001,In_26);
or U3313 (N_3313,In_116,In_1274);
xor U3314 (N_3314,In_1001,In_57);
nand U3315 (N_3315,In_630,In_1333);
or U3316 (N_3316,In_1750,In_1779);
or U3317 (N_3317,In_753,In_1095);
xor U3318 (N_3318,In_1951,In_223);
and U3319 (N_3319,In_401,In_863);
and U3320 (N_3320,In_1148,In_1039);
or U3321 (N_3321,In_1554,In_461);
xnor U3322 (N_3322,In_1781,In_347);
nand U3323 (N_3323,In_728,In_551);
or U3324 (N_3324,In_645,In_1931);
xor U3325 (N_3325,In_1469,In_1840);
and U3326 (N_3326,In_682,In_1361);
nor U3327 (N_3327,In_1589,In_1693);
nor U3328 (N_3328,In_504,In_34);
xnor U3329 (N_3329,In_277,In_907);
or U3330 (N_3330,In_481,In_1212);
nor U3331 (N_3331,In_746,In_1072);
nor U3332 (N_3332,In_982,In_1419);
and U3333 (N_3333,In_146,In_1372);
nor U3334 (N_3334,In_266,In_1082);
nand U3335 (N_3335,In_713,In_554);
and U3336 (N_3336,In_1367,In_517);
xor U3337 (N_3337,In_1128,In_903);
nand U3338 (N_3338,In_1875,In_886);
and U3339 (N_3339,In_623,In_1515);
nand U3340 (N_3340,In_120,In_95);
and U3341 (N_3341,In_1654,In_509);
and U3342 (N_3342,In_1138,In_1952);
nor U3343 (N_3343,In_1513,In_1440);
or U3344 (N_3344,In_1357,In_1663);
xor U3345 (N_3345,In_1811,In_552);
nand U3346 (N_3346,In_1236,In_805);
or U3347 (N_3347,In_1337,In_279);
nor U3348 (N_3348,In_1474,In_1525);
or U3349 (N_3349,In_1446,In_1138);
nor U3350 (N_3350,In_1099,In_1012);
nand U3351 (N_3351,In_1187,In_849);
nand U3352 (N_3352,In_1461,In_471);
or U3353 (N_3353,In_1710,In_1154);
or U3354 (N_3354,In_1886,In_352);
nor U3355 (N_3355,In_1146,In_722);
nor U3356 (N_3356,In_204,In_539);
nand U3357 (N_3357,In_1705,In_1004);
and U3358 (N_3358,In_404,In_1935);
nor U3359 (N_3359,In_1682,In_275);
nor U3360 (N_3360,In_502,In_224);
or U3361 (N_3361,In_468,In_981);
nor U3362 (N_3362,In_456,In_283);
and U3363 (N_3363,In_465,In_517);
and U3364 (N_3364,In_629,In_1833);
or U3365 (N_3365,In_1683,In_422);
nand U3366 (N_3366,In_934,In_1271);
and U3367 (N_3367,In_377,In_1175);
xnor U3368 (N_3368,In_620,In_160);
nor U3369 (N_3369,In_1803,In_1137);
and U3370 (N_3370,In_1610,In_850);
xor U3371 (N_3371,In_1918,In_715);
nand U3372 (N_3372,In_791,In_415);
xor U3373 (N_3373,In_1035,In_171);
nand U3374 (N_3374,In_1945,In_1990);
and U3375 (N_3375,In_1909,In_1102);
xnor U3376 (N_3376,In_1355,In_95);
and U3377 (N_3377,In_1887,In_1917);
or U3378 (N_3378,In_1641,In_660);
and U3379 (N_3379,In_27,In_299);
or U3380 (N_3380,In_683,In_739);
nor U3381 (N_3381,In_1625,In_10);
or U3382 (N_3382,In_111,In_1767);
xnor U3383 (N_3383,In_1422,In_1781);
or U3384 (N_3384,In_212,In_1883);
nor U3385 (N_3385,In_33,In_1229);
and U3386 (N_3386,In_831,In_454);
and U3387 (N_3387,In_107,In_1673);
nor U3388 (N_3388,In_75,In_1769);
and U3389 (N_3389,In_387,In_1404);
and U3390 (N_3390,In_869,In_420);
or U3391 (N_3391,In_1652,In_636);
nand U3392 (N_3392,In_1180,In_1243);
and U3393 (N_3393,In_929,In_1439);
and U3394 (N_3394,In_1208,In_120);
nand U3395 (N_3395,In_1034,In_472);
or U3396 (N_3396,In_89,In_1252);
nor U3397 (N_3397,In_405,In_621);
nand U3398 (N_3398,In_616,In_1332);
nand U3399 (N_3399,In_928,In_945);
nor U3400 (N_3400,In_1125,In_1190);
and U3401 (N_3401,In_1497,In_1915);
nor U3402 (N_3402,In_1907,In_841);
or U3403 (N_3403,In_680,In_1412);
or U3404 (N_3404,In_977,In_1018);
or U3405 (N_3405,In_1135,In_239);
xor U3406 (N_3406,In_1750,In_1840);
or U3407 (N_3407,In_1072,In_218);
and U3408 (N_3408,In_1784,In_636);
xnor U3409 (N_3409,In_78,In_601);
xor U3410 (N_3410,In_865,In_6);
or U3411 (N_3411,In_589,In_1238);
or U3412 (N_3412,In_1833,In_1220);
or U3413 (N_3413,In_163,In_149);
or U3414 (N_3414,In_85,In_1587);
or U3415 (N_3415,In_1936,In_61);
nor U3416 (N_3416,In_1748,In_213);
and U3417 (N_3417,In_736,In_975);
nand U3418 (N_3418,In_1703,In_620);
xnor U3419 (N_3419,In_1449,In_332);
or U3420 (N_3420,In_1580,In_1380);
xor U3421 (N_3421,In_1851,In_181);
xnor U3422 (N_3422,In_1877,In_473);
nor U3423 (N_3423,In_1512,In_382);
xnor U3424 (N_3424,In_9,In_624);
or U3425 (N_3425,In_1402,In_1964);
nor U3426 (N_3426,In_1804,In_188);
nor U3427 (N_3427,In_104,In_1561);
nand U3428 (N_3428,In_513,In_548);
nor U3429 (N_3429,In_1150,In_1210);
nand U3430 (N_3430,In_1079,In_1769);
and U3431 (N_3431,In_1775,In_326);
nor U3432 (N_3432,In_560,In_108);
and U3433 (N_3433,In_14,In_35);
nand U3434 (N_3434,In_693,In_788);
nand U3435 (N_3435,In_408,In_522);
xor U3436 (N_3436,In_385,In_278);
nor U3437 (N_3437,In_1474,In_696);
nand U3438 (N_3438,In_326,In_1704);
nor U3439 (N_3439,In_1659,In_742);
or U3440 (N_3440,In_596,In_613);
nor U3441 (N_3441,In_439,In_1975);
or U3442 (N_3442,In_842,In_1154);
xor U3443 (N_3443,In_424,In_201);
or U3444 (N_3444,In_1758,In_192);
or U3445 (N_3445,In_532,In_1759);
xnor U3446 (N_3446,In_747,In_648);
xor U3447 (N_3447,In_935,In_1117);
nand U3448 (N_3448,In_1168,In_1206);
xnor U3449 (N_3449,In_1735,In_1407);
nand U3450 (N_3450,In_165,In_544);
xnor U3451 (N_3451,In_517,In_854);
xor U3452 (N_3452,In_1735,In_625);
xor U3453 (N_3453,In_1477,In_31);
and U3454 (N_3454,In_1716,In_1873);
xnor U3455 (N_3455,In_130,In_1962);
xnor U3456 (N_3456,In_1288,In_966);
and U3457 (N_3457,In_1319,In_41);
and U3458 (N_3458,In_1185,In_186);
and U3459 (N_3459,In_590,In_49);
or U3460 (N_3460,In_1831,In_1281);
and U3461 (N_3461,In_352,In_209);
nor U3462 (N_3462,In_1761,In_1740);
nand U3463 (N_3463,In_887,In_1929);
nor U3464 (N_3464,In_1775,In_1456);
or U3465 (N_3465,In_190,In_405);
nand U3466 (N_3466,In_635,In_1879);
xnor U3467 (N_3467,In_1938,In_1088);
nor U3468 (N_3468,In_598,In_448);
xor U3469 (N_3469,In_959,In_1108);
nor U3470 (N_3470,In_720,In_1668);
xnor U3471 (N_3471,In_508,In_798);
nor U3472 (N_3472,In_1280,In_595);
or U3473 (N_3473,In_133,In_102);
or U3474 (N_3474,In_1600,In_544);
or U3475 (N_3475,In_1611,In_921);
or U3476 (N_3476,In_364,In_1393);
or U3477 (N_3477,In_1151,In_577);
or U3478 (N_3478,In_1503,In_60);
nor U3479 (N_3479,In_1070,In_904);
nand U3480 (N_3480,In_1125,In_81);
nor U3481 (N_3481,In_1884,In_1026);
and U3482 (N_3482,In_217,In_1904);
nor U3483 (N_3483,In_15,In_104);
nor U3484 (N_3484,In_893,In_1394);
or U3485 (N_3485,In_802,In_183);
nor U3486 (N_3486,In_646,In_449);
nand U3487 (N_3487,In_1773,In_798);
or U3488 (N_3488,In_321,In_1899);
xor U3489 (N_3489,In_447,In_1556);
and U3490 (N_3490,In_1811,In_1392);
xnor U3491 (N_3491,In_447,In_588);
xnor U3492 (N_3492,In_657,In_69);
nor U3493 (N_3493,In_112,In_767);
nand U3494 (N_3494,In_904,In_420);
or U3495 (N_3495,In_1288,In_1399);
xor U3496 (N_3496,In_1436,In_541);
nand U3497 (N_3497,In_1598,In_1299);
or U3498 (N_3498,In_1850,In_1528);
nor U3499 (N_3499,In_204,In_767);
nor U3500 (N_3500,In_1621,In_1632);
nor U3501 (N_3501,In_906,In_64);
and U3502 (N_3502,In_319,In_1714);
nor U3503 (N_3503,In_1925,In_1184);
nor U3504 (N_3504,In_1695,In_1519);
nor U3505 (N_3505,In_1609,In_257);
nand U3506 (N_3506,In_981,In_1695);
xor U3507 (N_3507,In_447,In_1646);
nor U3508 (N_3508,In_1968,In_699);
and U3509 (N_3509,In_1017,In_347);
nor U3510 (N_3510,In_701,In_1141);
nand U3511 (N_3511,In_963,In_987);
nor U3512 (N_3512,In_346,In_501);
nand U3513 (N_3513,In_12,In_1016);
and U3514 (N_3514,In_216,In_1139);
xnor U3515 (N_3515,In_82,In_1247);
xor U3516 (N_3516,In_933,In_1099);
nand U3517 (N_3517,In_1836,In_683);
xor U3518 (N_3518,In_961,In_623);
or U3519 (N_3519,In_1316,In_383);
xnor U3520 (N_3520,In_1461,In_337);
and U3521 (N_3521,In_1041,In_958);
or U3522 (N_3522,In_1449,In_1392);
nand U3523 (N_3523,In_418,In_1206);
nor U3524 (N_3524,In_1488,In_1310);
or U3525 (N_3525,In_1848,In_1668);
nand U3526 (N_3526,In_1723,In_958);
xor U3527 (N_3527,In_341,In_1041);
nor U3528 (N_3528,In_912,In_96);
or U3529 (N_3529,In_1751,In_1225);
xor U3530 (N_3530,In_1954,In_1345);
and U3531 (N_3531,In_1308,In_256);
xnor U3532 (N_3532,In_437,In_781);
nand U3533 (N_3533,In_412,In_1457);
nor U3534 (N_3534,In_1289,In_1210);
nand U3535 (N_3535,In_1620,In_989);
or U3536 (N_3536,In_474,In_1678);
nand U3537 (N_3537,In_765,In_576);
and U3538 (N_3538,In_1557,In_644);
or U3539 (N_3539,In_1461,In_218);
nor U3540 (N_3540,In_271,In_1920);
xnor U3541 (N_3541,In_1224,In_196);
nor U3542 (N_3542,In_946,In_204);
nand U3543 (N_3543,In_991,In_101);
or U3544 (N_3544,In_1857,In_165);
xnor U3545 (N_3545,In_879,In_1142);
and U3546 (N_3546,In_1068,In_55);
xnor U3547 (N_3547,In_546,In_366);
and U3548 (N_3548,In_13,In_27);
and U3549 (N_3549,In_1390,In_706);
and U3550 (N_3550,In_961,In_516);
xnor U3551 (N_3551,In_1434,In_1975);
and U3552 (N_3552,In_1499,In_1301);
and U3553 (N_3553,In_926,In_916);
xor U3554 (N_3554,In_1124,In_555);
and U3555 (N_3555,In_1594,In_1704);
nor U3556 (N_3556,In_292,In_1466);
or U3557 (N_3557,In_36,In_1027);
nand U3558 (N_3558,In_1591,In_300);
xnor U3559 (N_3559,In_133,In_561);
or U3560 (N_3560,In_278,In_277);
nor U3561 (N_3561,In_1266,In_1488);
or U3562 (N_3562,In_1587,In_388);
and U3563 (N_3563,In_613,In_1146);
nor U3564 (N_3564,In_968,In_532);
and U3565 (N_3565,In_244,In_1539);
nand U3566 (N_3566,In_367,In_713);
xnor U3567 (N_3567,In_189,In_1992);
xor U3568 (N_3568,In_712,In_478);
nand U3569 (N_3569,In_273,In_831);
xor U3570 (N_3570,In_1300,In_1159);
nand U3571 (N_3571,In_78,In_558);
nor U3572 (N_3572,In_1509,In_1450);
xnor U3573 (N_3573,In_1331,In_1386);
xor U3574 (N_3574,In_279,In_515);
or U3575 (N_3575,In_720,In_233);
xnor U3576 (N_3576,In_1883,In_234);
xor U3577 (N_3577,In_1648,In_1123);
nor U3578 (N_3578,In_104,In_1949);
xor U3579 (N_3579,In_1105,In_141);
nand U3580 (N_3580,In_1930,In_1573);
xnor U3581 (N_3581,In_1637,In_464);
xor U3582 (N_3582,In_519,In_1160);
nand U3583 (N_3583,In_465,In_1870);
and U3584 (N_3584,In_919,In_856);
xor U3585 (N_3585,In_91,In_1227);
nand U3586 (N_3586,In_1218,In_682);
xor U3587 (N_3587,In_1040,In_672);
nand U3588 (N_3588,In_1591,In_846);
nor U3589 (N_3589,In_389,In_883);
nor U3590 (N_3590,In_943,In_970);
nand U3591 (N_3591,In_637,In_835);
nand U3592 (N_3592,In_1792,In_1330);
and U3593 (N_3593,In_742,In_1724);
and U3594 (N_3594,In_1606,In_1511);
nand U3595 (N_3595,In_1885,In_1);
or U3596 (N_3596,In_117,In_670);
nand U3597 (N_3597,In_1734,In_124);
xnor U3598 (N_3598,In_433,In_1218);
xnor U3599 (N_3599,In_491,In_1508);
and U3600 (N_3600,In_1883,In_210);
nor U3601 (N_3601,In_1784,In_1781);
and U3602 (N_3602,In_230,In_1315);
xnor U3603 (N_3603,In_79,In_1753);
nor U3604 (N_3604,In_1244,In_1012);
and U3605 (N_3605,In_321,In_1574);
and U3606 (N_3606,In_278,In_1954);
xnor U3607 (N_3607,In_1801,In_737);
xnor U3608 (N_3608,In_310,In_1643);
xnor U3609 (N_3609,In_1408,In_1055);
or U3610 (N_3610,In_846,In_343);
nand U3611 (N_3611,In_34,In_169);
or U3612 (N_3612,In_134,In_141);
or U3613 (N_3613,In_1268,In_1440);
or U3614 (N_3614,In_488,In_868);
xnor U3615 (N_3615,In_1105,In_401);
xor U3616 (N_3616,In_1544,In_659);
xnor U3617 (N_3617,In_21,In_1079);
and U3618 (N_3618,In_1986,In_299);
or U3619 (N_3619,In_1607,In_960);
or U3620 (N_3620,In_1148,In_244);
or U3621 (N_3621,In_788,In_1620);
and U3622 (N_3622,In_1386,In_1341);
xnor U3623 (N_3623,In_681,In_199);
nand U3624 (N_3624,In_1608,In_851);
xor U3625 (N_3625,In_834,In_1117);
or U3626 (N_3626,In_924,In_1370);
xor U3627 (N_3627,In_509,In_1038);
and U3628 (N_3628,In_1787,In_1020);
and U3629 (N_3629,In_9,In_1307);
or U3630 (N_3630,In_425,In_126);
nor U3631 (N_3631,In_1771,In_613);
and U3632 (N_3632,In_188,In_60);
xnor U3633 (N_3633,In_1381,In_1643);
nand U3634 (N_3634,In_1205,In_659);
xnor U3635 (N_3635,In_842,In_599);
or U3636 (N_3636,In_1844,In_1370);
and U3637 (N_3637,In_1150,In_1079);
or U3638 (N_3638,In_1629,In_1612);
or U3639 (N_3639,In_828,In_1908);
xnor U3640 (N_3640,In_81,In_1002);
xnor U3641 (N_3641,In_1327,In_1150);
nor U3642 (N_3642,In_1734,In_1464);
xor U3643 (N_3643,In_106,In_1992);
and U3644 (N_3644,In_531,In_216);
or U3645 (N_3645,In_1203,In_1449);
or U3646 (N_3646,In_1136,In_1749);
xor U3647 (N_3647,In_849,In_1158);
nand U3648 (N_3648,In_209,In_622);
xnor U3649 (N_3649,In_1951,In_801);
nand U3650 (N_3650,In_1514,In_766);
or U3651 (N_3651,In_738,In_1236);
and U3652 (N_3652,In_712,In_1571);
xnor U3653 (N_3653,In_1779,In_898);
xnor U3654 (N_3654,In_1494,In_1890);
nor U3655 (N_3655,In_272,In_1462);
xor U3656 (N_3656,In_1610,In_149);
and U3657 (N_3657,In_1155,In_952);
and U3658 (N_3658,In_1073,In_682);
nand U3659 (N_3659,In_1123,In_1109);
or U3660 (N_3660,In_550,In_121);
nand U3661 (N_3661,In_1605,In_1352);
nand U3662 (N_3662,In_591,In_492);
or U3663 (N_3663,In_877,In_406);
nor U3664 (N_3664,In_109,In_1906);
nor U3665 (N_3665,In_135,In_720);
and U3666 (N_3666,In_938,In_1878);
nor U3667 (N_3667,In_1432,In_1325);
nor U3668 (N_3668,In_323,In_1166);
xnor U3669 (N_3669,In_679,In_534);
and U3670 (N_3670,In_718,In_1668);
xnor U3671 (N_3671,In_1629,In_1881);
xor U3672 (N_3672,In_1040,In_698);
nor U3673 (N_3673,In_925,In_839);
xor U3674 (N_3674,In_478,In_1557);
xnor U3675 (N_3675,In_599,In_1219);
nor U3676 (N_3676,In_1173,In_1755);
nand U3677 (N_3677,In_1993,In_1612);
or U3678 (N_3678,In_511,In_894);
or U3679 (N_3679,In_348,In_1204);
nand U3680 (N_3680,In_1650,In_1630);
and U3681 (N_3681,In_935,In_1949);
or U3682 (N_3682,In_1022,In_1726);
nor U3683 (N_3683,In_1203,In_948);
nor U3684 (N_3684,In_476,In_749);
or U3685 (N_3685,In_1684,In_1712);
nor U3686 (N_3686,In_1543,In_1599);
nand U3687 (N_3687,In_1255,In_415);
nand U3688 (N_3688,In_61,In_609);
nor U3689 (N_3689,In_1003,In_575);
nand U3690 (N_3690,In_471,In_1074);
and U3691 (N_3691,In_117,In_1278);
or U3692 (N_3692,In_372,In_404);
nand U3693 (N_3693,In_796,In_302);
and U3694 (N_3694,In_942,In_1051);
or U3695 (N_3695,In_1419,In_97);
nor U3696 (N_3696,In_268,In_732);
and U3697 (N_3697,In_1074,In_1143);
or U3698 (N_3698,In_317,In_1321);
nor U3699 (N_3699,In_76,In_956);
nor U3700 (N_3700,In_1235,In_1490);
nand U3701 (N_3701,In_479,In_1607);
nor U3702 (N_3702,In_1091,In_1078);
xnor U3703 (N_3703,In_1989,In_324);
nor U3704 (N_3704,In_1375,In_847);
or U3705 (N_3705,In_610,In_525);
or U3706 (N_3706,In_1534,In_272);
and U3707 (N_3707,In_1777,In_1259);
xor U3708 (N_3708,In_492,In_287);
nand U3709 (N_3709,In_284,In_1927);
nor U3710 (N_3710,In_1319,In_145);
nor U3711 (N_3711,In_1011,In_1791);
xor U3712 (N_3712,In_1088,In_441);
and U3713 (N_3713,In_1522,In_446);
nor U3714 (N_3714,In_1504,In_36);
nor U3715 (N_3715,In_757,In_109);
xnor U3716 (N_3716,In_1033,In_353);
nand U3717 (N_3717,In_303,In_814);
xnor U3718 (N_3718,In_648,In_694);
nand U3719 (N_3719,In_805,In_562);
or U3720 (N_3720,In_386,In_1265);
or U3721 (N_3721,In_1424,In_1556);
nand U3722 (N_3722,In_1452,In_631);
nor U3723 (N_3723,In_1753,In_525);
nand U3724 (N_3724,In_118,In_426);
nor U3725 (N_3725,In_1557,In_511);
or U3726 (N_3726,In_1578,In_1528);
xnor U3727 (N_3727,In_1217,In_401);
and U3728 (N_3728,In_690,In_1021);
nand U3729 (N_3729,In_1308,In_692);
and U3730 (N_3730,In_1642,In_1113);
xnor U3731 (N_3731,In_881,In_1621);
nand U3732 (N_3732,In_1522,In_624);
and U3733 (N_3733,In_1873,In_59);
nor U3734 (N_3734,In_138,In_604);
xor U3735 (N_3735,In_1308,In_634);
or U3736 (N_3736,In_643,In_1929);
nor U3737 (N_3737,In_469,In_672);
nand U3738 (N_3738,In_515,In_1384);
or U3739 (N_3739,In_1119,In_1559);
nand U3740 (N_3740,In_1603,In_423);
xor U3741 (N_3741,In_708,In_1827);
xor U3742 (N_3742,In_1943,In_1272);
nor U3743 (N_3743,In_47,In_1640);
and U3744 (N_3744,In_1771,In_238);
nor U3745 (N_3745,In_1889,In_722);
xnor U3746 (N_3746,In_1944,In_1524);
nand U3747 (N_3747,In_363,In_335);
nor U3748 (N_3748,In_298,In_1411);
nand U3749 (N_3749,In_1697,In_425);
and U3750 (N_3750,In_664,In_788);
or U3751 (N_3751,In_869,In_1445);
xor U3752 (N_3752,In_737,In_1876);
and U3753 (N_3753,In_283,In_1446);
nor U3754 (N_3754,In_1723,In_694);
nor U3755 (N_3755,In_235,In_1761);
or U3756 (N_3756,In_1989,In_1534);
xor U3757 (N_3757,In_1151,In_1572);
or U3758 (N_3758,In_100,In_120);
xor U3759 (N_3759,In_1166,In_1577);
and U3760 (N_3760,In_347,In_308);
or U3761 (N_3761,In_1893,In_335);
or U3762 (N_3762,In_1674,In_1298);
nor U3763 (N_3763,In_1593,In_1347);
and U3764 (N_3764,In_37,In_112);
xor U3765 (N_3765,In_1478,In_267);
nand U3766 (N_3766,In_1842,In_385);
or U3767 (N_3767,In_1104,In_1808);
and U3768 (N_3768,In_477,In_1904);
nor U3769 (N_3769,In_981,In_266);
nor U3770 (N_3770,In_906,In_1565);
nand U3771 (N_3771,In_1287,In_281);
nor U3772 (N_3772,In_819,In_855);
nand U3773 (N_3773,In_649,In_1837);
or U3774 (N_3774,In_612,In_1396);
nand U3775 (N_3775,In_873,In_323);
xnor U3776 (N_3776,In_1316,In_458);
nor U3777 (N_3777,In_910,In_269);
xnor U3778 (N_3778,In_1161,In_875);
or U3779 (N_3779,In_1731,In_568);
nand U3780 (N_3780,In_1091,In_1442);
nand U3781 (N_3781,In_524,In_143);
or U3782 (N_3782,In_1910,In_672);
nor U3783 (N_3783,In_1182,In_1728);
and U3784 (N_3784,In_19,In_1916);
nand U3785 (N_3785,In_1532,In_1269);
xor U3786 (N_3786,In_1119,In_430);
nor U3787 (N_3787,In_1018,In_459);
or U3788 (N_3788,In_1842,In_466);
nand U3789 (N_3789,In_1336,In_875);
and U3790 (N_3790,In_887,In_403);
xor U3791 (N_3791,In_1531,In_1839);
or U3792 (N_3792,In_594,In_1727);
nand U3793 (N_3793,In_1552,In_1010);
nor U3794 (N_3794,In_1679,In_460);
or U3795 (N_3795,In_925,In_995);
nand U3796 (N_3796,In_1964,In_1733);
nand U3797 (N_3797,In_1258,In_308);
and U3798 (N_3798,In_183,In_984);
xor U3799 (N_3799,In_972,In_1125);
or U3800 (N_3800,In_1113,In_1002);
nand U3801 (N_3801,In_1577,In_1494);
nor U3802 (N_3802,In_1859,In_1412);
nor U3803 (N_3803,In_1883,In_11);
nand U3804 (N_3804,In_1380,In_936);
or U3805 (N_3805,In_160,In_44);
nor U3806 (N_3806,In_1422,In_1163);
xor U3807 (N_3807,In_836,In_705);
xnor U3808 (N_3808,In_159,In_643);
xnor U3809 (N_3809,In_1169,In_1247);
or U3810 (N_3810,In_1555,In_736);
xnor U3811 (N_3811,In_1201,In_1088);
xnor U3812 (N_3812,In_642,In_378);
xnor U3813 (N_3813,In_1,In_1367);
or U3814 (N_3814,In_488,In_1769);
nand U3815 (N_3815,In_1227,In_1470);
or U3816 (N_3816,In_1807,In_1444);
nand U3817 (N_3817,In_667,In_655);
xnor U3818 (N_3818,In_1558,In_149);
nand U3819 (N_3819,In_1790,In_1529);
nand U3820 (N_3820,In_1801,In_1381);
xor U3821 (N_3821,In_291,In_408);
nand U3822 (N_3822,In_825,In_1141);
xnor U3823 (N_3823,In_1642,In_100);
nand U3824 (N_3824,In_359,In_1765);
xnor U3825 (N_3825,In_1062,In_1175);
nor U3826 (N_3826,In_693,In_993);
and U3827 (N_3827,In_611,In_166);
and U3828 (N_3828,In_1988,In_1797);
nand U3829 (N_3829,In_168,In_436);
or U3830 (N_3830,In_1989,In_263);
or U3831 (N_3831,In_827,In_224);
and U3832 (N_3832,In_281,In_375);
or U3833 (N_3833,In_896,In_1916);
nand U3834 (N_3834,In_620,In_1699);
nand U3835 (N_3835,In_1156,In_934);
nor U3836 (N_3836,In_1598,In_600);
xnor U3837 (N_3837,In_1880,In_4);
and U3838 (N_3838,In_1053,In_1417);
nor U3839 (N_3839,In_1340,In_1545);
nand U3840 (N_3840,In_982,In_642);
or U3841 (N_3841,In_1816,In_1767);
nand U3842 (N_3842,In_631,In_564);
and U3843 (N_3843,In_940,In_127);
or U3844 (N_3844,In_112,In_758);
and U3845 (N_3845,In_476,In_288);
nor U3846 (N_3846,In_711,In_1464);
xnor U3847 (N_3847,In_1295,In_405);
xnor U3848 (N_3848,In_1412,In_977);
and U3849 (N_3849,In_1170,In_750);
nor U3850 (N_3850,In_1398,In_238);
nand U3851 (N_3851,In_907,In_591);
or U3852 (N_3852,In_797,In_1468);
xor U3853 (N_3853,In_1890,In_1258);
and U3854 (N_3854,In_1052,In_37);
or U3855 (N_3855,In_1709,In_576);
nor U3856 (N_3856,In_1955,In_1330);
xnor U3857 (N_3857,In_1315,In_1809);
or U3858 (N_3858,In_1206,In_689);
or U3859 (N_3859,In_711,In_310);
nor U3860 (N_3860,In_1441,In_1317);
nand U3861 (N_3861,In_520,In_658);
nor U3862 (N_3862,In_1813,In_1402);
nor U3863 (N_3863,In_731,In_1406);
xnor U3864 (N_3864,In_1224,In_1765);
nor U3865 (N_3865,In_614,In_75);
xnor U3866 (N_3866,In_1908,In_568);
nor U3867 (N_3867,In_693,In_790);
nor U3868 (N_3868,In_83,In_1155);
or U3869 (N_3869,In_1513,In_1845);
or U3870 (N_3870,In_1250,In_615);
and U3871 (N_3871,In_1833,In_1313);
or U3872 (N_3872,In_1045,In_508);
or U3873 (N_3873,In_1040,In_779);
nor U3874 (N_3874,In_1392,In_1635);
nor U3875 (N_3875,In_340,In_740);
nand U3876 (N_3876,In_1341,In_815);
nor U3877 (N_3877,In_1105,In_1483);
or U3878 (N_3878,In_1633,In_1381);
and U3879 (N_3879,In_194,In_787);
nand U3880 (N_3880,In_416,In_63);
xnor U3881 (N_3881,In_721,In_1570);
or U3882 (N_3882,In_353,In_812);
and U3883 (N_3883,In_440,In_277);
nor U3884 (N_3884,In_770,In_1488);
nand U3885 (N_3885,In_1246,In_1121);
or U3886 (N_3886,In_817,In_1697);
xnor U3887 (N_3887,In_464,In_273);
and U3888 (N_3888,In_453,In_1863);
and U3889 (N_3889,In_1838,In_605);
and U3890 (N_3890,In_170,In_1368);
or U3891 (N_3891,In_458,In_1786);
or U3892 (N_3892,In_900,In_556);
or U3893 (N_3893,In_655,In_225);
and U3894 (N_3894,In_1653,In_1554);
and U3895 (N_3895,In_793,In_46);
and U3896 (N_3896,In_177,In_52);
xor U3897 (N_3897,In_1681,In_71);
or U3898 (N_3898,In_7,In_328);
and U3899 (N_3899,In_1379,In_1614);
nor U3900 (N_3900,In_985,In_210);
xor U3901 (N_3901,In_608,In_844);
nand U3902 (N_3902,In_1653,In_993);
nand U3903 (N_3903,In_1685,In_774);
or U3904 (N_3904,In_1766,In_1674);
or U3905 (N_3905,In_1116,In_176);
nand U3906 (N_3906,In_1899,In_609);
and U3907 (N_3907,In_1389,In_1235);
nand U3908 (N_3908,In_1458,In_503);
nand U3909 (N_3909,In_1041,In_583);
and U3910 (N_3910,In_857,In_1589);
xor U3911 (N_3911,In_1735,In_1606);
xor U3912 (N_3912,In_1621,In_1374);
nand U3913 (N_3913,In_532,In_1735);
xnor U3914 (N_3914,In_1280,In_1044);
nor U3915 (N_3915,In_1794,In_1979);
and U3916 (N_3916,In_1167,In_925);
xnor U3917 (N_3917,In_327,In_245);
xnor U3918 (N_3918,In_448,In_1748);
or U3919 (N_3919,In_222,In_746);
nand U3920 (N_3920,In_166,In_1018);
xor U3921 (N_3921,In_872,In_639);
and U3922 (N_3922,In_696,In_1039);
nand U3923 (N_3923,In_1813,In_1481);
nor U3924 (N_3924,In_146,In_1767);
or U3925 (N_3925,In_874,In_870);
nor U3926 (N_3926,In_1984,In_340);
and U3927 (N_3927,In_268,In_1343);
and U3928 (N_3928,In_1822,In_544);
xor U3929 (N_3929,In_885,In_80);
nand U3930 (N_3930,In_696,In_1906);
or U3931 (N_3931,In_1320,In_1318);
nor U3932 (N_3932,In_1944,In_427);
and U3933 (N_3933,In_1949,In_1807);
and U3934 (N_3934,In_433,In_1349);
nand U3935 (N_3935,In_467,In_1027);
nor U3936 (N_3936,In_126,In_1884);
nand U3937 (N_3937,In_1873,In_1218);
or U3938 (N_3938,In_727,In_1942);
and U3939 (N_3939,In_800,In_238);
nor U3940 (N_3940,In_1710,In_241);
nor U3941 (N_3941,In_1354,In_942);
and U3942 (N_3942,In_1989,In_672);
xnor U3943 (N_3943,In_1552,In_1524);
nor U3944 (N_3944,In_1417,In_1142);
and U3945 (N_3945,In_859,In_736);
xnor U3946 (N_3946,In_704,In_1264);
or U3947 (N_3947,In_1106,In_220);
nor U3948 (N_3948,In_474,In_797);
nor U3949 (N_3949,In_1566,In_1294);
and U3950 (N_3950,In_1607,In_523);
or U3951 (N_3951,In_1558,In_0);
xor U3952 (N_3952,In_1435,In_1716);
and U3953 (N_3953,In_736,In_939);
nor U3954 (N_3954,In_1191,In_416);
and U3955 (N_3955,In_82,In_849);
or U3956 (N_3956,In_36,In_544);
and U3957 (N_3957,In_1611,In_68);
nand U3958 (N_3958,In_644,In_322);
nand U3959 (N_3959,In_254,In_1542);
nand U3960 (N_3960,In_1503,In_1133);
or U3961 (N_3961,In_486,In_1802);
nand U3962 (N_3962,In_1869,In_890);
nand U3963 (N_3963,In_488,In_56);
xor U3964 (N_3964,In_1106,In_135);
or U3965 (N_3965,In_1093,In_1851);
or U3966 (N_3966,In_280,In_1730);
or U3967 (N_3967,In_115,In_31);
or U3968 (N_3968,In_1579,In_1493);
xnor U3969 (N_3969,In_1806,In_1261);
and U3970 (N_3970,In_557,In_679);
nor U3971 (N_3971,In_643,In_413);
xnor U3972 (N_3972,In_538,In_1515);
nor U3973 (N_3973,In_1351,In_1009);
nor U3974 (N_3974,In_966,In_964);
nor U3975 (N_3975,In_1430,In_387);
nand U3976 (N_3976,In_1252,In_958);
and U3977 (N_3977,In_202,In_1903);
or U3978 (N_3978,In_996,In_822);
or U3979 (N_3979,In_1696,In_1986);
nand U3980 (N_3980,In_715,In_509);
xor U3981 (N_3981,In_499,In_1921);
nand U3982 (N_3982,In_608,In_1375);
and U3983 (N_3983,In_958,In_472);
xor U3984 (N_3984,In_309,In_206);
and U3985 (N_3985,In_1002,In_13);
xor U3986 (N_3986,In_1404,In_699);
xor U3987 (N_3987,In_1105,In_1766);
nor U3988 (N_3988,In_1938,In_1616);
or U3989 (N_3989,In_397,In_102);
and U3990 (N_3990,In_1230,In_465);
xor U3991 (N_3991,In_288,In_934);
or U3992 (N_3992,In_1755,In_1203);
xor U3993 (N_3993,In_107,In_1087);
or U3994 (N_3994,In_1751,In_1026);
and U3995 (N_3995,In_374,In_1127);
nor U3996 (N_3996,In_1640,In_78);
xnor U3997 (N_3997,In_452,In_1433);
and U3998 (N_3998,In_1260,In_1889);
nand U3999 (N_3999,In_565,In_633);
nand U4000 (N_4000,In_143,In_1736);
nand U4001 (N_4001,In_740,In_86);
and U4002 (N_4002,In_1279,In_1105);
nor U4003 (N_4003,In_1595,In_1235);
nand U4004 (N_4004,In_338,In_931);
xor U4005 (N_4005,In_973,In_840);
xor U4006 (N_4006,In_1352,In_1580);
nor U4007 (N_4007,In_1173,In_1335);
nand U4008 (N_4008,In_1862,In_111);
xor U4009 (N_4009,In_1420,In_1179);
and U4010 (N_4010,In_1082,In_1559);
and U4011 (N_4011,In_1562,In_1081);
and U4012 (N_4012,In_730,In_1825);
xnor U4013 (N_4013,In_1117,In_27);
nand U4014 (N_4014,In_1751,In_1406);
nand U4015 (N_4015,In_1012,In_1888);
xor U4016 (N_4016,In_969,In_840);
nor U4017 (N_4017,In_252,In_1226);
and U4018 (N_4018,In_1362,In_45);
xor U4019 (N_4019,In_1818,In_995);
xor U4020 (N_4020,In_501,In_1210);
nand U4021 (N_4021,In_31,In_1437);
xor U4022 (N_4022,In_41,In_954);
and U4023 (N_4023,In_1033,In_1628);
and U4024 (N_4024,In_776,In_1735);
nor U4025 (N_4025,In_126,In_1717);
nor U4026 (N_4026,In_584,In_332);
nor U4027 (N_4027,In_253,In_1006);
xor U4028 (N_4028,In_1176,In_1281);
nor U4029 (N_4029,In_1953,In_579);
nor U4030 (N_4030,In_461,In_885);
and U4031 (N_4031,In_585,In_286);
or U4032 (N_4032,In_1474,In_1761);
and U4033 (N_4033,In_41,In_501);
nor U4034 (N_4034,In_165,In_726);
and U4035 (N_4035,In_678,In_1207);
and U4036 (N_4036,In_1952,In_1326);
nand U4037 (N_4037,In_232,In_1404);
and U4038 (N_4038,In_168,In_442);
or U4039 (N_4039,In_401,In_1830);
nand U4040 (N_4040,In_230,In_35);
nand U4041 (N_4041,In_101,In_715);
nor U4042 (N_4042,In_841,In_1671);
nand U4043 (N_4043,In_104,In_1324);
and U4044 (N_4044,In_279,In_183);
nand U4045 (N_4045,In_134,In_280);
and U4046 (N_4046,In_959,In_1506);
xor U4047 (N_4047,In_1666,In_498);
or U4048 (N_4048,In_629,In_1431);
and U4049 (N_4049,In_829,In_1756);
and U4050 (N_4050,In_733,In_1536);
and U4051 (N_4051,In_587,In_1340);
or U4052 (N_4052,In_1590,In_409);
and U4053 (N_4053,In_602,In_1112);
and U4054 (N_4054,In_405,In_394);
xor U4055 (N_4055,In_1576,In_1904);
xnor U4056 (N_4056,In_316,In_1149);
xor U4057 (N_4057,In_706,In_855);
xnor U4058 (N_4058,In_1837,In_430);
xnor U4059 (N_4059,In_1691,In_1819);
and U4060 (N_4060,In_1380,In_876);
nand U4061 (N_4061,In_1050,In_642);
nor U4062 (N_4062,In_820,In_1609);
nand U4063 (N_4063,In_446,In_125);
or U4064 (N_4064,In_47,In_1970);
nand U4065 (N_4065,In_1229,In_1097);
xor U4066 (N_4066,In_20,In_56);
nand U4067 (N_4067,In_387,In_918);
xnor U4068 (N_4068,In_502,In_384);
and U4069 (N_4069,In_868,In_957);
nand U4070 (N_4070,In_58,In_1791);
xor U4071 (N_4071,In_910,In_762);
nor U4072 (N_4072,In_1765,In_1602);
and U4073 (N_4073,In_1351,In_1769);
nand U4074 (N_4074,In_1007,In_1182);
and U4075 (N_4075,In_1633,In_1799);
nor U4076 (N_4076,In_335,In_1152);
and U4077 (N_4077,In_1124,In_36);
and U4078 (N_4078,In_489,In_1938);
and U4079 (N_4079,In_1326,In_1117);
xnor U4080 (N_4080,In_1635,In_1256);
or U4081 (N_4081,In_70,In_1117);
or U4082 (N_4082,In_607,In_369);
or U4083 (N_4083,In_991,In_871);
or U4084 (N_4084,In_1403,In_444);
nand U4085 (N_4085,In_1546,In_57);
or U4086 (N_4086,In_635,In_1534);
xnor U4087 (N_4087,In_1983,In_961);
nand U4088 (N_4088,In_1436,In_660);
nor U4089 (N_4089,In_395,In_766);
xnor U4090 (N_4090,In_792,In_994);
and U4091 (N_4091,In_938,In_1290);
or U4092 (N_4092,In_148,In_1888);
or U4093 (N_4093,In_640,In_274);
xor U4094 (N_4094,In_1718,In_103);
xor U4095 (N_4095,In_1834,In_1401);
xor U4096 (N_4096,In_1211,In_876);
and U4097 (N_4097,In_1663,In_41);
nor U4098 (N_4098,In_1763,In_1252);
nor U4099 (N_4099,In_1140,In_87);
nor U4100 (N_4100,In_688,In_1475);
or U4101 (N_4101,In_1916,In_1252);
nand U4102 (N_4102,In_1784,In_1045);
nand U4103 (N_4103,In_306,In_1112);
and U4104 (N_4104,In_1908,In_685);
nand U4105 (N_4105,In_41,In_1396);
xor U4106 (N_4106,In_1135,In_1797);
or U4107 (N_4107,In_203,In_1660);
nand U4108 (N_4108,In_563,In_62);
xor U4109 (N_4109,In_1630,In_1527);
nand U4110 (N_4110,In_217,In_1144);
or U4111 (N_4111,In_1478,In_1403);
nor U4112 (N_4112,In_1981,In_510);
nand U4113 (N_4113,In_727,In_453);
nor U4114 (N_4114,In_201,In_237);
xor U4115 (N_4115,In_1148,In_337);
nor U4116 (N_4116,In_33,In_650);
and U4117 (N_4117,In_623,In_313);
and U4118 (N_4118,In_584,In_293);
and U4119 (N_4119,In_1643,In_1076);
xor U4120 (N_4120,In_1206,In_1265);
xnor U4121 (N_4121,In_1352,In_542);
nor U4122 (N_4122,In_1102,In_541);
xnor U4123 (N_4123,In_1425,In_1730);
or U4124 (N_4124,In_1289,In_1430);
and U4125 (N_4125,In_1093,In_1651);
nor U4126 (N_4126,In_1370,In_176);
nor U4127 (N_4127,In_849,In_185);
or U4128 (N_4128,In_731,In_1968);
nand U4129 (N_4129,In_1849,In_1759);
and U4130 (N_4130,In_1207,In_1894);
nor U4131 (N_4131,In_1152,In_1843);
or U4132 (N_4132,In_218,In_907);
nand U4133 (N_4133,In_638,In_1690);
nor U4134 (N_4134,In_1815,In_541);
nor U4135 (N_4135,In_549,In_20);
or U4136 (N_4136,In_878,In_666);
nor U4137 (N_4137,In_1259,In_1430);
nand U4138 (N_4138,In_537,In_427);
xnor U4139 (N_4139,In_1950,In_1767);
and U4140 (N_4140,In_562,In_1784);
nand U4141 (N_4141,In_499,In_1476);
nor U4142 (N_4142,In_1059,In_714);
xnor U4143 (N_4143,In_1990,In_733);
and U4144 (N_4144,In_1364,In_825);
or U4145 (N_4145,In_1512,In_1919);
or U4146 (N_4146,In_904,In_1759);
and U4147 (N_4147,In_955,In_315);
nor U4148 (N_4148,In_1055,In_1143);
nor U4149 (N_4149,In_345,In_1878);
and U4150 (N_4150,In_1873,In_499);
or U4151 (N_4151,In_365,In_565);
nor U4152 (N_4152,In_201,In_22);
and U4153 (N_4153,In_909,In_1997);
nand U4154 (N_4154,In_1410,In_291);
and U4155 (N_4155,In_1073,In_535);
and U4156 (N_4156,In_845,In_1999);
and U4157 (N_4157,In_1732,In_404);
xor U4158 (N_4158,In_56,In_1574);
or U4159 (N_4159,In_1574,In_756);
xor U4160 (N_4160,In_1975,In_783);
and U4161 (N_4161,In_1917,In_860);
nand U4162 (N_4162,In_1760,In_1468);
nor U4163 (N_4163,In_242,In_472);
and U4164 (N_4164,In_1209,In_938);
and U4165 (N_4165,In_196,In_1594);
xnor U4166 (N_4166,In_1348,In_447);
or U4167 (N_4167,In_1792,In_727);
and U4168 (N_4168,In_87,In_958);
xnor U4169 (N_4169,In_72,In_944);
nand U4170 (N_4170,In_889,In_312);
nand U4171 (N_4171,In_197,In_1061);
nand U4172 (N_4172,In_1979,In_652);
and U4173 (N_4173,In_1599,In_777);
xor U4174 (N_4174,In_1963,In_24);
or U4175 (N_4175,In_87,In_1160);
or U4176 (N_4176,In_392,In_1498);
nand U4177 (N_4177,In_679,In_1932);
or U4178 (N_4178,In_1186,In_1678);
nand U4179 (N_4179,In_397,In_1378);
xnor U4180 (N_4180,In_152,In_1279);
nand U4181 (N_4181,In_496,In_1483);
nor U4182 (N_4182,In_1336,In_338);
nand U4183 (N_4183,In_1387,In_1581);
and U4184 (N_4184,In_933,In_51);
or U4185 (N_4185,In_1046,In_804);
nand U4186 (N_4186,In_86,In_1730);
nand U4187 (N_4187,In_1933,In_823);
and U4188 (N_4188,In_239,In_1605);
nand U4189 (N_4189,In_346,In_1302);
xor U4190 (N_4190,In_1225,In_575);
xor U4191 (N_4191,In_1592,In_1143);
and U4192 (N_4192,In_772,In_110);
and U4193 (N_4193,In_1050,In_1935);
and U4194 (N_4194,In_832,In_1373);
nor U4195 (N_4195,In_1090,In_302);
xnor U4196 (N_4196,In_1475,In_1973);
or U4197 (N_4197,In_503,In_1916);
and U4198 (N_4198,In_1994,In_1757);
xnor U4199 (N_4199,In_262,In_612);
xor U4200 (N_4200,In_1661,In_136);
nor U4201 (N_4201,In_555,In_1673);
or U4202 (N_4202,In_49,In_689);
and U4203 (N_4203,In_1610,In_696);
and U4204 (N_4204,In_602,In_234);
or U4205 (N_4205,In_407,In_190);
nand U4206 (N_4206,In_957,In_1086);
and U4207 (N_4207,In_1574,In_639);
or U4208 (N_4208,In_127,In_1028);
or U4209 (N_4209,In_1437,In_1952);
and U4210 (N_4210,In_1747,In_1138);
and U4211 (N_4211,In_1265,In_1388);
or U4212 (N_4212,In_476,In_1009);
or U4213 (N_4213,In_671,In_674);
nor U4214 (N_4214,In_1906,In_876);
or U4215 (N_4215,In_1369,In_338);
or U4216 (N_4216,In_495,In_300);
xnor U4217 (N_4217,In_1345,In_586);
nand U4218 (N_4218,In_1503,In_209);
nor U4219 (N_4219,In_289,In_1015);
nor U4220 (N_4220,In_1531,In_628);
nand U4221 (N_4221,In_711,In_1543);
nand U4222 (N_4222,In_1057,In_511);
and U4223 (N_4223,In_418,In_206);
or U4224 (N_4224,In_179,In_1543);
or U4225 (N_4225,In_1216,In_378);
nor U4226 (N_4226,In_1142,In_751);
or U4227 (N_4227,In_660,In_865);
nor U4228 (N_4228,In_730,In_514);
nor U4229 (N_4229,In_1754,In_1639);
xnor U4230 (N_4230,In_1079,In_1218);
nor U4231 (N_4231,In_660,In_1818);
xnor U4232 (N_4232,In_1238,In_1553);
xnor U4233 (N_4233,In_1295,In_1681);
nand U4234 (N_4234,In_1296,In_1872);
and U4235 (N_4235,In_1631,In_292);
nand U4236 (N_4236,In_1462,In_1873);
nor U4237 (N_4237,In_425,In_1563);
xor U4238 (N_4238,In_1768,In_1315);
xor U4239 (N_4239,In_1850,In_1844);
xnor U4240 (N_4240,In_1046,In_514);
and U4241 (N_4241,In_1714,In_1098);
nand U4242 (N_4242,In_1744,In_1906);
nand U4243 (N_4243,In_817,In_1258);
xnor U4244 (N_4244,In_314,In_970);
or U4245 (N_4245,In_1846,In_787);
nand U4246 (N_4246,In_52,In_1476);
and U4247 (N_4247,In_1329,In_1700);
nor U4248 (N_4248,In_1381,In_1036);
or U4249 (N_4249,In_1281,In_954);
nand U4250 (N_4250,In_1290,In_1171);
xnor U4251 (N_4251,In_1790,In_86);
xor U4252 (N_4252,In_996,In_826);
nor U4253 (N_4253,In_1906,In_111);
and U4254 (N_4254,In_1777,In_1469);
nand U4255 (N_4255,In_509,In_1537);
or U4256 (N_4256,In_1773,In_1273);
nand U4257 (N_4257,In_1940,In_1896);
nor U4258 (N_4258,In_1417,In_492);
and U4259 (N_4259,In_1803,In_163);
xor U4260 (N_4260,In_1843,In_26);
or U4261 (N_4261,In_32,In_790);
and U4262 (N_4262,In_439,In_1348);
xnor U4263 (N_4263,In_1300,In_1240);
xor U4264 (N_4264,In_1844,In_1037);
nand U4265 (N_4265,In_948,In_1069);
xnor U4266 (N_4266,In_898,In_43);
nand U4267 (N_4267,In_1261,In_183);
nand U4268 (N_4268,In_1907,In_98);
or U4269 (N_4269,In_1364,In_68);
nor U4270 (N_4270,In_832,In_1553);
and U4271 (N_4271,In_1359,In_1354);
xor U4272 (N_4272,In_48,In_1564);
nor U4273 (N_4273,In_565,In_1380);
and U4274 (N_4274,In_60,In_1298);
nand U4275 (N_4275,In_1219,In_1531);
or U4276 (N_4276,In_225,In_464);
xnor U4277 (N_4277,In_1249,In_928);
nand U4278 (N_4278,In_1469,In_1298);
nor U4279 (N_4279,In_900,In_1430);
and U4280 (N_4280,In_1770,In_1683);
or U4281 (N_4281,In_1194,In_538);
nor U4282 (N_4282,In_236,In_20);
nand U4283 (N_4283,In_1102,In_1231);
and U4284 (N_4284,In_422,In_83);
and U4285 (N_4285,In_1634,In_45);
xnor U4286 (N_4286,In_1391,In_46);
nor U4287 (N_4287,In_177,In_1317);
xor U4288 (N_4288,In_1795,In_933);
nor U4289 (N_4289,In_1455,In_358);
or U4290 (N_4290,In_968,In_1812);
and U4291 (N_4291,In_645,In_1347);
nor U4292 (N_4292,In_922,In_902);
xor U4293 (N_4293,In_1911,In_15);
and U4294 (N_4294,In_1489,In_154);
nor U4295 (N_4295,In_1764,In_1144);
nor U4296 (N_4296,In_580,In_1414);
and U4297 (N_4297,In_1922,In_1208);
nand U4298 (N_4298,In_296,In_1034);
and U4299 (N_4299,In_904,In_1817);
nor U4300 (N_4300,In_411,In_1288);
nor U4301 (N_4301,In_786,In_752);
and U4302 (N_4302,In_1159,In_260);
nand U4303 (N_4303,In_1187,In_1429);
nor U4304 (N_4304,In_1521,In_1251);
or U4305 (N_4305,In_1933,In_996);
nand U4306 (N_4306,In_268,In_484);
or U4307 (N_4307,In_1821,In_780);
nand U4308 (N_4308,In_1072,In_863);
or U4309 (N_4309,In_35,In_209);
nand U4310 (N_4310,In_802,In_1091);
and U4311 (N_4311,In_623,In_1059);
or U4312 (N_4312,In_1637,In_186);
nor U4313 (N_4313,In_126,In_1301);
xor U4314 (N_4314,In_19,In_1341);
nand U4315 (N_4315,In_1337,In_1559);
nor U4316 (N_4316,In_787,In_28);
nor U4317 (N_4317,In_551,In_1149);
nand U4318 (N_4318,In_353,In_697);
nand U4319 (N_4319,In_1313,In_768);
xnor U4320 (N_4320,In_754,In_973);
and U4321 (N_4321,In_1291,In_226);
nor U4322 (N_4322,In_1685,In_1437);
nand U4323 (N_4323,In_287,In_1675);
xor U4324 (N_4324,In_1099,In_1731);
nor U4325 (N_4325,In_1259,In_747);
nand U4326 (N_4326,In_1202,In_1666);
or U4327 (N_4327,In_678,In_365);
nor U4328 (N_4328,In_769,In_1453);
xor U4329 (N_4329,In_441,In_490);
xor U4330 (N_4330,In_789,In_1280);
nor U4331 (N_4331,In_1084,In_1466);
nor U4332 (N_4332,In_997,In_739);
and U4333 (N_4333,In_1502,In_759);
xnor U4334 (N_4334,In_1953,In_964);
and U4335 (N_4335,In_891,In_181);
and U4336 (N_4336,In_1864,In_347);
xnor U4337 (N_4337,In_962,In_237);
nand U4338 (N_4338,In_1480,In_1547);
nor U4339 (N_4339,In_1648,In_1704);
or U4340 (N_4340,In_641,In_552);
and U4341 (N_4341,In_394,In_1383);
xor U4342 (N_4342,In_360,In_1025);
nand U4343 (N_4343,In_721,In_174);
and U4344 (N_4344,In_859,In_490);
nand U4345 (N_4345,In_1890,In_1747);
nand U4346 (N_4346,In_471,In_1625);
and U4347 (N_4347,In_1905,In_376);
nand U4348 (N_4348,In_710,In_626);
nand U4349 (N_4349,In_1056,In_1168);
nand U4350 (N_4350,In_1349,In_1677);
nand U4351 (N_4351,In_597,In_145);
nor U4352 (N_4352,In_688,In_1339);
and U4353 (N_4353,In_1070,In_97);
nand U4354 (N_4354,In_520,In_69);
and U4355 (N_4355,In_18,In_868);
nor U4356 (N_4356,In_1649,In_1156);
or U4357 (N_4357,In_838,In_1789);
nor U4358 (N_4358,In_1819,In_81);
xnor U4359 (N_4359,In_923,In_752);
nand U4360 (N_4360,In_448,In_1205);
or U4361 (N_4361,In_171,In_487);
xor U4362 (N_4362,In_1356,In_984);
nand U4363 (N_4363,In_540,In_1726);
and U4364 (N_4364,In_1467,In_1527);
and U4365 (N_4365,In_683,In_1170);
or U4366 (N_4366,In_1426,In_997);
and U4367 (N_4367,In_87,In_425);
nand U4368 (N_4368,In_883,In_444);
or U4369 (N_4369,In_70,In_354);
and U4370 (N_4370,In_28,In_598);
nand U4371 (N_4371,In_762,In_1040);
nand U4372 (N_4372,In_149,In_1172);
or U4373 (N_4373,In_156,In_1695);
xnor U4374 (N_4374,In_1247,In_1960);
nand U4375 (N_4375,In_693,In_747);
nor U4376 (N_4376,In_1578,In_104);
and U4377 (N_4377,In_1311,In_848);
nor U4378 (N_4378,In_533,In_1908);
xor U4379 (N_4379,In_1755,In_623);
xor U4380 (N_4380,In_339,In_1829);
and U4381 (N_4381,In_997,In_734);
or U4382 (N_4382,In_1535,In_633);
nand U4383 (N_4383,In_1571,In_1462);
nor U4384 (N_4384,In_1024,In_1785);
or U4385 (N_4385,In_1342,In_1438);
and U4386 (N_4386,In_1024,In_1075);
or U4387 (N_4387,In_1691,In_627);
nor U4388 (N_4388,In_35,In_838);
and U4389 (N_4389,In_1086,In_1887);
xnor U4390 (N_4390,In_288,In_1827);
nand U4391 (N_4391,In_826,In_895);
nand U4392 (N_4392,In_1132,In_1997);
or U4393 (N_4393,In_951,In_173);
nor U4394 (N_4394,In_1284,In_978);
xnor U4395 (N_4395,In_948,In_1044);
and U4396 (N_4396,In_1219,In_1204);
or U4397 (N_4397,In_1443,In_684);
xnor U4398 (N_4398,In_1436,In_112);
nor U4399 (N_4399,In_851,In_337);
nand U4400 (N_4400,In_336,In_1613);
xor U4401 (N_4401,In_591,In_243);
or U4402 (N_4402,In_455,In_1816);
nor U4403 (N_4403,In_465,In_696);
or U4404 (N_4404,In_1828,In_1039);
and U4405 (N_4405,In_1541,In_1073);
xor U4406 (N_4406,In_679,In_1130);
nand U4407 (N_4407,In_254,In_266);
and U4408 (N_4408,In_1575,In_120);
nor U4409 (N_4409,In_48,In_777);
or U4410 (N_4410,In_354,In_1725);
or U4411 (N_4411,In_626,In_1481);
or U4412 (N_4412,In_928,In_445);
and U4413 (N_4413,In_979,In_720);
xnor U4414 (N_4414,In_1730,In_778);
xor U4415 (N_4415,In_1592,In_1894);
xor U4416 (N_4416,In_1371,In_1964);
nand U4417 (N_4417,In_611,In_345);
nand U4418 (N_4418,In_1357,In_714);
and U4419 (N_4419,In_795,In_581);
xor U4420 (N_4420,In_1218,In_1902);
xor U4421 (N_4421,In_1956,In_125);
xor U4422 (N_4422,In_340,In_896);
or U4423 (N_4423,In_1286,In_110);
xor U4424 (N_4424,In_900,In_271);
and U4425 (N_4425,In_272,In_1087);
nand U4426 (N_4426,In_1071,In_189);
and U4427 (N_4427,In_970,In_1776);
and U4428 (N_4428,In_1186,In_1806);
and U4429 (N_4429,In_201,In_1688);
xnor U4430 (N_4430,In_296,In_657);
nand U4431 (N_4431,In_1174,In_1997);
or U4432 (N_4432,In_828,In_1927);
xor U4433 (N_4433,In_160,In_254);
xor U4434 (N_4434,In_358,In_977);
or U4435 (N_4435,In_1943,In_1562);
nor U4436 (N_4436,In_152,In_658);
xor U4437 (N_4437,In_483,In_1572);
nor U4438 (N_4438,In_1190,In_1221);
nor U4439 (N_4439,In_1168,In_1680);
nor U4440 (N_4440,In_1563,In_1455);
nand U4441 (N_4441,In_1584,In_409);
xor U4442 (N_4442,In_198,In_1071);
nand U4443 (N_4443,In_1042,In_1330);
xor U4444 (N_4444,In_1571,In_644);
and U4445 (N_4445,In_1098,In_185);
nor U4446 (N_4446,In_1029,In_1185);
nor U4447 (N_4447,In_1796,In_1945);
nor U4448 (N_4448,In_540,In_1593);
nand U4449 (N_4449,In_1303,In_1472);
and U4450 (N_4450,In_463,In_1573);
and U4451 (N_4451,In_1151,In_403);
or U4452 (N_4452,In_1742,In_1065);
or U4453 (N_4453,In_466,In_182);
nand U4454 (N_4454,In_1245,In_1079);
nand U4455 (N_4455,In_1345,In_929);
nor U4456 (N_4456,In_313,In_511);
nand U4457 (N_4457,In_936,In_1320);
or U4458 (N_4458,In_1415,In_42);
or U4459 (N_4459,In_768,In_621);
and U4460 (N_4460,In_1812,In_109);
or U4461 (N_4461,In_1434,In_294);
nor U4462 (N_4462,In_1864,In_636);
nor U4463 (N_4463,In_1332,In_45);
and U4464 (N_4464,In_1603,In_1922);
xnor U4465 (N_4465,In_259,In_1817);
or U4466 (N_4466,In_1242,In_1642);
and U4467 (N_4467,In_1013,In_729);
nor U4468 (N_4468,In_116,In_659);
or U4469 (N_4469,In_983,In_681);
nor U4470 (N_4470,In_799,In_768);
or U4471 (N_4471,In_265,In_864);
nand U4472 (N_4472,In_769,In_507);
xnor U4473 (N_4473,In_1369,In_692);
nor U4474 (N_4474,In_1603,In_1126);
and U4475 (N_4475,In_1725,In_409);
xor U4476 (N_4476,In_291,In_1691);
xor U4477 (N_4477,In_135,In_1294);
or U4478 (N_4478,In_1627,In_1214);
and U4479 (N_4479,In_1914,In_57);
or U4480 (N_4480,In_1640,In_647);
nand U4481 (N_4481,In_619,In_659);
xnor U4482 (N_4482,In_378,In_36);
xnor U4483 (N_4483,In_659,In_1499);
or U4484 (N_4484,In_239,In_803);
xor U4485 (N_4485,In_1577,In_479);
nor U4486 (N_4486,In_79,In_1320);
or U4487 (N_4487,In_16,In_845);
xnor U4488 (N_4488,In_342,In_1573);
nand U4489 (N_4489,In_1421,In_1055);
or U4490 (N_4490,In_569,In_683);
or U4491 (N_4491,In_559,In_1776);
nand U4492 (N_4492,In_156,In_1753);
and U4493 (N_4493,In_1573,In_535);
nand U4494 (N_4494,In_306,In_1400);
nand U4495 (N_4495,In_1637,In_501);
and U4496 (N_4496,In_1625,In_1274);
nor U4497 (N_4497,In_1306,In_1496);
nor U4498 (N_4498,In_598,In_1633);
and U4499 (N_4499,In_600,In_827);
or U4500 (N_4500,In_369,In_10);
nand U4501 (N_4501,In_1953,In_840);
and U4502 (N_4502,In_1283,In_56);
nand U4503 (N_4503,In_544,In_513);
xnor U4504 (N_4504,In_1413,In_37);
and U4505 (N_4505,In_830,In_97);
xnor U4506 (N_4506,In_537,In_276);
and U4507 (N_4507,In_49,In_329);
and U4508 (N_4508,In_804,In_1141);
or U4509 (N_4509,In_1022,In_482);
or U4510 (N_4510,In_522,In_1002);
nand U4511 (N_4511,In_945,In_1436);
xnor U4512 (N_4512,In_641,In_233);
or U4513 (N_4513,In_1049,In_888);
or U4514 (N_4514,In_528,In_442);
and U4515 (N_4515,In_790,In_123);
or U4516 (N_4516,In_1063,In_1043);
and U4517 (N_4517,In_403,In_404);
nand U4518 (N_4518,In_1244,In_237);
and U4519 (N_4519,In_1995,In_666);
xnor U4520 (N_4520,In_1281,In_197);
xor U4521 (N_4521,In_1027,In_1936);
xor U4522 (N_4522,In_1161,In_1679);
or U4523 (N_4523,In_1135,In_687);
nand U4524 (N_4524,In_1948,In_1228);
nand U4525 (N_4525,In_1159,In_1883);
xnor U4526 (N_4526,In_1492,In_843);
nand U4527 (N_4527,In_50,In_677);
and U4528 (N_4528,In_299,In_1563);
and U4529 (N_4529,In_228,In_1414);
nand U4530 (N_4530,In_1029,In_52);
nand U4531 (N_4531,In_1786,In_207);
nand U4532 (N_4532,In_1924,In_802);
and U4533 (N_4533,In_1743,In_507);
nor U4534 (N_4534,In_931,In_136);
and U4535 (N_4535,In_1236,In_1951);
nand U4536 (N_4536,In_1928,In_1004);
xnor U4537 (N_4537,In_498,In_1797);
nand U4538 (N_4538,In_730,In_1168);
nor U4539 (N_4539,In_1073,In_1259);
or U4540 (N_4540,In_1658,In_708);
nor U4541 (N_4541,In_238,In_1248);
nor U4542 (N_4542,In_1190,In_974);
xnor U4543 (N_4543,In_1312,In_1424);
and U4544 (N_4544,In_927,In_310);
and U4545 (N_4545,In_456,In_670);
and U4546 (N_4546,In_537,In_1099);
nor U4547 (N_4547,In_257,In_1604);
or U4548 (N_4548,In_423,In_1555);
nor U4549 (N_4549,In_1839,In_366);
nor U4550 (N_4550,In_1605,In_1188);
nand U4551 (N_4551,In_172,In_779);
and U4552 (N_4552,In_365,In_599);
nand U4553 (N_4553,In_1681,In_15);
nand U4554 (N_4554,In_1185,In_1063);
xor U4555 (N_4555,In_1150,In_16);
and U4556 (N_4556,In_611,In_1612);
xnor U4557 (N_4557,In_1426,In_400);
xnor U4558 (N_4558,In_670,In_1198);
or U4559 (N_4559,In_1222,In_722);
or U4560 (N_4560,In_620,In_1170);
nor U4561 (N_4561,In_1040,In_1101);
nand U4562 (N_4562,In_138,In_1176);
or U4563 (N_4563,In_1077,In_1569);
xnor U4564 (N_4564,In_572,In_856);
and U4565 (N_4565,In_259,In_345);
nand U4566 (N_4566,In_83,In_1239);
and U4567 (N_4567,In_1098,In_87);
nor U4568 (N_4568,In_548,In_425);
nor U4569 (N_4569,In_752,In_488);
xnor U4570 (N_4570,In_1372,In_1604);
nor U4571 (N_4571,In_37,In_696);
nand U4572 (N_4572,In_1927,In_948);
nor U4573 (N_4573,In_1030,In_1925);
and U4574 (N_4574,In_991,In_877);
and U4575 (N_4575,In_1666,In_1149);
or U4576 (N_4576,In_516,In_679);
xnor U4577 (N_4577,In_607,In_1217);
xnor U4578 (N_4578,In_760,In_1164);
and U4579 (N_4579,In_1533,In_121);
nor U4580 (N_4580,In_282,In_368);
or U4581 (N_4581,In_828,In_62);
nand U4582 (N_4582,In_967,In_1351);
or U4583 (N_4583,In_1803,In_442);
xor U4584 (N_4584,In_924,In_1859);
and U4585 (N_4585,In_1195,In_1535);
nand U4586 (N_4586,In_1694,In_334);
or U4587 (N_4587,In_1577,In_1410);
or U4588 (N_4588,In_585,In_1719);
or U4589 (N_4589,In_1942,In_1397);
nor U4590 (N_4590,In_1593,In_788);
xnor U4591 (N_4591,In_642,In_486);
xor U4592 (N_4592,In_1794,In_1575);
nor U4593 (N_4593,In_789,In_169);
nor U4594 (N_4594,In_800,In_110);
and U4595 (N_4595,In_1200,In_1213);
or U4596 (N_4596,In_358,In_190);
and U4597 (N_4597,In_1571,In_1752);
nand U4598 (N_4598,In_1285,In_1733);
xor U4599 (N_4599,In_718,In_1456);
nand U4600 (N_4600,In_1972,In_548);
and U4601 (N_4601,In_1963,In_1089);
nor U4602 (N_4602,In_587,In_740);
xnor U4603 (N_4603,In_1879,In_1566);
xnor U4604 (N_4604,In_1093,In_986);
and U4605 (N_4605,In_1223,In_1332);
nand U4606 (N_4606,In_1003,In_837);
nor U4607 (N_4607,In_1249,In_804);
or U4608 (N_4608,In_226,In_1719);
or U4609 (N_4609,In_944,In_1128);
xor U4610 (N_4610,In_963,In_184);
xnor U4611 (N_4611,In_1030,In_9);
xnor U4612 (N_4612,In_1271,In_533);
nand U4613 (N_4613,In_1861,In_1244);
or U4614 (N_4614,In_797,In_1236);
and U4615 (N_4615,In_1470,In_663);
nand U4616 (N_4616,In_1287,In_1181);
and U4617 (N_4617,In_1696,In_519);
and U4618 (N_4618,In_1804,In_1214);
and U4619 (N_4619,In_1700,In_791);
nor U4620 (N_4620,In_1415,In_1493);
nand U4621 (N_4621,In_580,In_1736);
and U4622 (N_4622,In_4,In_393);
and U4623 (N_4623,In_202,In_1418);
or U4624 (N_4624,In_543,In_326);
nor U4625 (N_4625,In_1008,In_1337);
xor U4626 (N_4626,In_1575,In_1179);
nor U4627 (N_4627,In_1172,In_1805);
or U4628 (N_4628,In_890,In_651);
xnor U4629 (N_4629,In_1605,In_1451);
nor U4630 (N_4630,In_1873,In_1846);
or U4631 (N_4631,In_1082,In_854);
xor U4632 (N_4632,In_37,In_584);
and U4633 (N_4633,In_981,In_1754);
nand U4634 (N_4634,In_1513,In_771);
xor U4635 (N_4635,In_1683,In_871);
and U4636 (N_4636,In_879,In_1627);
nor U4637 (N_4637,In_477,In_130);
nor U4638 (N_4638,In_1781,In_1123);
nor U4639 (N_4639,In_1259,In_1356);
nor U4640 (N_4640,In_724,In_753);
nor U4641 (N_4641,In_897,In_894);
xor U4642 (N_4642,In_536,In_1736);
and U4643 (N_4643,In_224,In_28);
nor U4644 (N_4644,In_1364,In_359);
xor U4645 (N_4645,In_1165,In_558);
xor U4646 (N_4646,In_207,In_1082);
and U4647 (N_4647,In_1723,In_152);
nor U4648 (N_4648,In_310,In_1069);
or U4649 (N_4649,In_1037,In_249);
nand U4650 (N_4650,In_1197,In_185);
or U4651 (N_4651,In_241,In_1447);
nor U4652 (N_4652,In_1092,In_729);
nor U4653 (N_4653,In_1274,In_1312);
or U4654 (N_4654,In_287,In_1131);
xnor U4655 (N_4655,In_1424,In_1551);
xor U4656 (N_4656,In_536,In_103);
or U4657 (N_4657,In_322,In_294);
and U4658 (N_4658,In_1002,In_677);
nand U4659 (N_4659,In_1863,In_34);
or U4660 (N_4660,In_1761,In_1165);
or U4661 (N_4661,In_1109,In_1790);
nor U4662 (N_4662,In_1546,In_71);
or U4663 (N_4663,In_34,In_645);
or U4664 (N_4664,In_472,In_1321);
nor U4665 (N_4665,In_1754,In_1565);
and U4666 (N_4666,In_1329,In_66);
nand U4667 (N_4667,In_1801,In_125);
nand U4668 (N_4668,In_756,In_1298);
or U4669 (N_4669,In_1464,In_1627);
or U4670 (N_4670,In_1598,In_1395);
nand U4671 (N_4671,In_158,In_1199);
or U4672 (N_4672,In_453,In_1754);
and U4673 (N_4673,In_1993,In_1668);
xor U4674 (N_4674,In_1359,In_700);
or U4675 (N_4675,In_1916,In_1958);
xnor U4676 (N_4676,In_1128,In_547);
nor U4677 (N_4677,In_1841,In_1982);
and U4678 (N_4678,In_1235,In_1949);
xor U4679 (N_4679,In_902,In_1897);
nor U4680 (N_4680,In_1759,In_1992);
nor U4681 (N_4681,In_1846,In_1168);
or U4682 (N_4682,In_860,In_718);
nand U4683 (N_4683,In_428,In_1267);
or U4684 (N_4684,In_104,In_682);
or U4685 (N_4685,In_559,In_635);
or U4686 (N_4686,In_1971,In_445);
or U4687 (N_4687,In_1286,In_1709);
and U4688 (N_4688,In_797,In_1143);
nor U4689 (N_4689,In_634,In_832);
and U4690 (N_4690,In_52,In_658);
nor U4691 (N_4691,In_1221,In_1301);
or U4692 (N_4692,In_1069,In_917);
and U4693 (N_4693,In_1455,In_776);
nor U4694 (N_4694,In_1420,In_158);
and U4695 (N_4695,In_7,In_1917);
nor U4696 (N_4696,In_480,In_80);
nor U4697 (N_4697,In_1542,In_472);
nor U4698 (N_4698,In_1286,In_713);
and U4699 (N_4699,In_1179,In_1474);
or U4700 (N_4700,In_92,In_585);
or U4701 (N_4701,In_1613,In_1999);
nand U4702 (N_4702,In_577,In_700);
nor U4703 (N_4703,In_700,In_1160);
or U4704 (N_4704,In_288,In_747);
xnor U4705 (N_4705,In_302,In_1151);
nor U4706 (N_4706,In_1872,In_64);
and U4707 (N_4707,In_540,In_617);
or U4708 (N_4708,In_290,In_714);
nor U4709 (N_4709,In_680,In_75);
nand U4710 (N_4710,In_136,In_1958);
nand U4711 (N_4711,In_1853,In_1922);
nand U4712 (N_4712,In_1637,In_1740);
or U4713 (N_4713,In_1795,In_865);
nand U4714 (N_4714,In_1418,In_233);
and U4715 (N_4715,In_639,In_1598);
xnor U4716 (N_4716,In_1585,In_643);
nor U4717 (N_4717,In_1937,In_1844);
nor U4718 (N_4718,In_1658,In_1991);
and U4719 (N_4719,In_701,In_788);
xor U4720 (N_4720,In_1865,In_1160);
and U4721 (N_4721,In_984,In_160);
or U4722 (N_4722,In_497,In_1172);
or U4723 (N_4723,In_1118,In_29);
or U4724 (N_4724,In_1179,In_1317);
nand U4725 (N_4725,In_376,In_1238);
nor U4726 (N_4726,In_606,In_784);
xor U4727 (N_4727,In_423,In_308);
xor U4728 (N_4728,In_1389,In_316);
xnor U4729 (N_4729,In_1027,In_1856);
nand U4730 (N_4730,In_45,In_359);
and U4731 (N_4731,In_125,In_590);
xor U4732 (N_4732,In_939,In_1492);
and U4733 (N_4733,In_1665,In_400);
or U4734 (N_4734,In_1281,In_1898);
nand U4735 (N_4735,In_350,In_1546);
nand U4736 (N_4736,In_304,In_1172);
nand U4737 (N_4737,In_311,In_305);
nor U4738 (N_4738,In_624,In_1707);
and U4739 (N_4739,In_991,In_1384);
or U4740 (N_4740,In_1332,In_602);
xor U4741 (N_4741,In_1119,In_581);
nor U4742 (N_4742,In_1804,In_346);
nor U4743 (N_4743,In_862,In_1078);
or U4744 (N_4744,In_850,In_485);
or U4745 (N_4745,In_1715,In_1169);
and U4746 (N_4746,In_786,In_760);
or U4747 (N_4747,In_172,In_1572);
xor U4748 (N_4748,In_262,In_1586);
xor U4749 (N_4749,In_314,In_208);
or U4750 (N_4750,In_818,In_1457);
xnor U4751 (N_4751,In_1464,In_748);
or U4752 (N_4752,In_1925,In_1132);
or U4753 (N_4753,In_1918,In_196);
xnor U4754 (N_4754,In_1472,In_1144);
nor U4755 (N_4755,In_1507,In_276);
xnor U4756 (N_4756,In_1006,In_542);
or U4757 (N_4757,In_1915,In_1181);
nor U4758 (N_4758,In_1570,In_1061);
xor U4759 (N_4759,In_1296,In_1492);
nor U4760 (N_4760,In_735,In_410);
and U4761 (N_4761,In_1325,In_803);
xor U4762 (N_4762,In_324,In_1281);
nor U4763 (N_4763,In_1145,In_1253);
xor U4764 (N_4764,In_1959,In_1118);
nor U4765 (N_4765,In_1276,In_621);
and U4766 (N_4766,In_1838,In_827);
nand U4767 (N_4767,In_316,In_1083);
nand U4768 (N_4768,In_1262,In_669);
nand U4769 (N_4769,In_401,In_944);
and U4770 (N_4770,In_181,In_1980);
nor U4771 (N_4771,In_1189,In_781);
nor U4772 (N_4772,In_458,In_1938);
nand U4773 (N_4773,In_1994,In_850);
or U4774 (N_4774,In_1132,In_638);
nand U4775 (N_4775,In_1833,In_270);
or U4776 (N_4776,In_135,In_408);
or U4777 (N_4777,In_1936,In_657);
and U4778 (N_4778,In_862,In_482);
nand U4779 (N_4779,In_1085,In_1347);
nand U4780 (N_4780,In_790,In_650);
nand U4781 (N_4781,In_785,In_933);
or U4782 (N_4782,In_414,In_1905);
or U4783 (N_4783,In_1253,In_163);
or U4784 (N_4784,In_897,In_1392);
or U4785 (N_4785,In_645,In_892);
and U4786 (N_4786,In_1193,In_1772);
and U4787 (N_4787,In_1064,In_1763);
and U4788 (N_4788,In_1953,In_1808);
and U4789 (N_4789,In_762,In_1670);
nor U4790 (N_4790,In_423,In_665);
nor U4791 (N_4791,In_1634,In_1888);
nand U4792 (N_4792,In_833,In_109);
or U4793 (N_4793,In_179,In_1569);
nand U4794 (N_4794,In_1265,In_239);
nor U4795 (N_4795,In_402,In_1305);
or U4796 (N_4796,In_681,In_611);
or U4797 (N_4797,In_14,In_1041);
nor U4798 (N_4798,In_1393,In_657);
and U4799 (N_4799,In_1241,In_1338);
xnor U4800 (N_4800,In_960,In_1566);
and U4801 (N_4801,In_33,In_1875);
and U4802 (N_4802,In_1297,In_156);
or U4803 (N_4803,In_1179,In_345);
or U4804 (N_4804,In_261,In_340);
or U4805 (N_4805,In_1056,In_1272);
nor U4806 (N_4806,In_1507,In_467);
and U4807 (N_4807,In_540,In_294);
or U4808 (N_4808,In_1833,In_301);
xor U4809 (N_4809,In_1202,In_808);
and U4810 (N_4810,In_741,In_1601);
xnor U4811 (N_4811,In_887,In_1578);
xor U4812 (N_4812,In_944,In_1602);
nor U4813 (N_4813,In_236,In_1758);
xnor U4814 (N_4814,In_580,In_1339);
nand U4815 (N_4815,In_367,In_1628);
or U4816 (N_4816,In_620,In_797);
nor U4817 (N_4817,In_811,In_680);
or U4818 (N_4818,In_612,In_241);
xnor U4819 (N_4819,In_1654,In_1427);
or U4820 (N_4820,In_1947,In_575);
nor U4821 (N_4821,In_530,In_541);
nand U4822 (N_4822,In_482,In_1817);
or U4823 (N_4823,In_102,In_899);
or U4824 (N_4824,In_1295,In_1734);
nand U4825 (N_4825,In_421,In_977);
nand U4826 (N_4826,In_1127,In_1951);
and U4827 (N_4827,In_1087,In_215);
nor U4828 (N_4828,In_1500,In_1165);
nand U4829 (N_4829,In_857,In_1675);
and U4830 (N_4830,In_1712,In_1277);
xor U4831 (N_4831,In_1652,In_1081);
nand U4832 (N_4832,In_336,In_1302);
nor U4833 (N_4833,In_1470,In_91);
or U4834 (N_4834,In_105,In_727);
xor U4835 (N_4835,In_712,In_1502);
xnor U4836 (N_4836,In_1925,In_1166);
nor U4837 (N_4837,In_534,In_833);
nand U4838 (N_4838,In_1866,In_297);
or U4839 (N_4839,In_1793,In_243);
xor U4840 (N_4840,In_1400,In_1757);
xor U4841 (N_4841,In_1161,In_1194);
nand U4842 (N_4842,In_80,In_510);
xor U4843 (N_4843,In_1729,In_676);
nor U4844 (N_4844,In_763,In_770);
xnor U4845 (N_4845,In_1989,In_1896);
xor U4846 (N_4846,In_1678,In_661);
or U4847 (N_4847,In_1122,In_866);
nand U4848 (N_4848,In_209,In_1711);
xor U4849 (N_4849,In_1377,In_529);
and U4850 (N_4850,In_1352,In_839);
or U4851 (N_4851,In_1290,In_1695);
xor U4852 (N_4852,In_618,In_458);
xor U4853 (N_4853,In_654,In_1619);
xor U4854 (N_4854,In_1113,In_1469);
nand U4855 (N_4855,In_583,In_1951);
nand U4856 (N_4856,In_992,In_1156);
xnor U4857 (N_4857,In_658,In_1929);
nand U4858 (N_4858,In_916,In_1914);
nand U4859 (N_4859,In_1243,In_915);
or U4860 (N_4860,In_140,In_258);
and U4861 (N_4861,In_1014,In_1350);
xor U4862 (N_4862,In_279,In_542);
nor U4863 (N_4863,In_673,In_640);
or U4864 (N_4864,In_824,In_642);
xor U4865 (N_4865,In_1047,In_1798);
or U4866 (N_4866,In_1002,In_371);
nand U4867 (N_4867,In_1498,In_359);
nor U4868 (N_4868,In_1711,In_1504);
nor U4869 (N_4869,In_1149,In_867);
xor U4870 (N_4870,In_993,In_979);
nand U4871 (N_4871,In_1530,In_728);
nand U4872 (N_4872,In_1371,In_1558);
xor U4873 (N_4873,In_506,In_487);
xor U4874 (N_4874,In_60,In_1038);
or U4875 (N_4875,In_672,In_1851);
or U4876 (N_4876,In_542,In_18);
or U4877 (N_4877,In_34,In_131);
or U4878 (N_4878,In_840,In_670);
nor U4879 (N_4879,In_604,In_706);
nand U4880 (N_4880,In_1154,In_508);
xnor U4881 (N_4881,In_1826,In_747);
xnor U4882 (N_4882,In_1902,In_1587);
xnor U4883 (N_4883,In_594,In_1142);
or U4884 (N_4884,In_982,In_1488);
and U4885 (N_4885,In_1056,In_1547);
or U4886 (N_4886,In_676,In_45);
xor U4887 (N_4887,In_1574,In_1086);
nand U4888 (N_4888,In_552,In_1311);
nand U4889 (N_4889,In_2,In_745);
and U4890 (N_4890,In_1503,In_1400);
nor U4891 (N_4891,In_1192,In_289);
or U4892 (N_4892,In_1742,In_1147);
or U4893 (N_4893,In_1621,In_771);
nand U4894 (N_4894,In_1282,In_915);
or U4895 (N_4895,In_756,In_1658);
nand U4896 (N_4896,In_1797,In_821);
nand U4897 (N_4897,In_889,In_1241);
or U4898 (N_4898,In_490,In_1784);
nand U4899 (N_4899,In_747,In_1793);
or U4900 (N_4900,In_1365,In_1239);
nand U4901 (N_4901,In_184,In_1681);
xor U4902 (N_4902,In_1902,In_543);
xnor U4903 (N_4903,In_190,In_252);
nor U4904 (N_4904,In_489,In_535);
nor U4905 (N_4905,In_477,In_1245);
or U4906 (N_4906,In_264,In_738);
xnor U4907 (N_4907,In_1287,In_1888);
nand U4908 (N_4908,In_580,In_396);
or U4909 (N_4909,In_1220,In_1718);
or U4910 (N_4910,In_170,In_582);
and U4911 (N_4911,In_1333,In_1575);
or U4912 (N_4912,In_168,In_429);
nand U4913 (N_4913,In_1918,In_1184);
nor U4914 (N_4914,In_1883,In_749);
nor U4915 (N_4915,In_1948,In_1356);
xor U4916 (N_4916,In_1610,In_1433);
nor U4917 (N_4917,In_900,In_156);
xnor U4918 (N_4918,In_744,In_1830);
and U4919 (N_4919,In_641,In_1373);
or U4920 (N_4920,In_1487,In_1179);
nor U4921 (N_4921,In_942,In_317);
nand U4922 (N_4922,In_790,In_31);
xor U4923 (N_4923,In_876,In_1054);
nand U4924 (N_4924,In_737,In_961);
xor U4925 (N_4925,In_405,In_315);
nor U4926 (N_4926,In_369,In_664);
xnor U4927 (N_4927,In_1390,In_1229);
nand U4928 (N_4928,In_1056,In_92);
nor U4929 (N_4929,In_1054,In_673);
and U4930 (N_4930,In_1832,In_1125);
and U4931 (N_4931,In_247,In_1989);
nand U4932 (N_4932,In_1050,In_776);
nand U4933 (N_4933,In_816,In_1353);
and U4934 (N_4934,In_444,In_816);
nand U4935 (N_4935,In_883,In_1859);
or U4936 (N_4936,In_1125,In_836);
and U4937 (N_4937,In_358,In_98);
nand U4938 (N_4938,In_1805,In_1242);
nand U4939 (N_4939,In_1506,In_1154);
nand U4940 (N_4940,In_1400,In_888);
or U4941 (N_4941,In_1710,In_395);
or U4942 (N_4942,In_53,In_1989);
xor U4943 (N_4943,In_944,In_156);
or U4944 (N_4944,In_977,In_870);
nand U4945 (N_4945,In_1969,In_1359);
and U4946 (N_4946,In_916,In_978);
nor U4947 (N_4947,In_1681,In_1947);
xnor U4948 (N_4948,In_1746,In_1990);
xnor U4949 (N_4949,In_1764,In_787);
nor U4950 (N_4950,In_1759,In_87);
or U4951 (N_4951,In_1177,In_292);
nand U4952 (N_4952,In_440,In_1103);
and U4953 (N_4953,In_623,In_1390);
xor U4954 (N_4954,In_842,In_906);
xor U4955 (N_4955,In_1814,In_1866);
nand U4956 (N_4956,In_972,In_825);
xnor U4957 (N_4957,In_1160,In_1353);
and U4958 (N_4958,In_1190,In_1419);
xor U4959 (N_4959,In_1680,In_1822);
nor U4960 (N_4960,In_1875,In_619);
and U4961 (N_4961,In_223,In_927);
nand U4962 (N_4962,In_357,In_1097);
or U4963 (N_4963,In_1518,In_820);
nand U4964 (N_4964,In_1776,In_1028);
or U4965 (N_4965,In_93,In_1702);
and U4966 (N_4966,In_181,In_108);
nor U4967 (N_4967,In_601,In_349);
or U4968 (N_4968,In_1675,In_1179);
xnor U4969 (N_4969,In_1497,In_1303);
nor U4970 (N_4970,In_848,In_1004);
or U4971 (N_4971,In_1606,In_530);
or U4972 (N_4972,In_1050,In_1642);
nor U4973 (N_4973,In_1790,In_1497);
nand U4974 (N_4974,In_288,In_1089);
and U4975 (N_4975,In_1857,In_1911);
and U4976 (N_4976,In_198,In_467);
or U4977 (N_4977,In_222,In_330);
or U4978 (N_4978,In_798,In_1653);
nand U4979 (N_4979,In_1386,In_261);
and U4980 (N_4980,In_51,In_68);
xor U4981 (N_4981,In_1539,In_1692);
nor U4982 (N_4982,In_1289,In_568);
xor U4983 (N_4983,In_180,In_1627);
and U4984 (N_4984,In_986,In_158);
and U4985 (N_4985,In_1704,In_159);
xor U4986 (N_4986,In_675,In_1183);
xnor U4987 (N_4987,In_472,In_282);
nand U4988 (N_4988,In_584,In_513);
nand U4989 (N_4989,In_1866,In_1759);
nor U4990 (N_4990,In_1304,In_878);
nand U4991 (N_4991,In_535,In_904);
or U4992 (N_4992,In_1211,In_948);
xor U4993 (N_4993,In_446,In_23);
and U4994 (N_4994,In_777,In_1443);
nor U4995 (N_4995,In_904,In_941);
xnor U4996 (N_4996,In_1931,In_1289);
and U4997 (N_4997,In_513,In_1163);
or U4998 (N_4998,In_951,In_505);
nor U4999 (N_4999,In_1790,In_1884);
or U5000 (N_5000,N_4087,N_2423);
or U5001 (N_5001,N_3385,N_2587);
or U5002 (N_5002,N_2835,N_913);
nor U5003 (N_5003,N_4270,N_3080);
xor U5004 (N_5004,N_4838,N_9);
nor U5005 (N_5005,N_2130,N_3061);
nand U5006 (N_5006,N_483,N_1926);
and U5007 (N_5007,N_281,N_1388);
nand U5008 (N_5008,N_1725,N_4013);
xnor U5009 (N_5009,N_3770,N_3811);
nand U5010 (N_5010,N_2115,N_2634);
xor U5011 (N_5011,N_4525,N_43);
nand U5012 (N_5012,N_2348,N_3124);
xor U5013 (N_5013,N_2193,N_664);
nand U5014 (N_5014,N_541,N_4743);
or U5015 (N_5015,N_535,N_3041);
xor U5016 (N_5016,N_1941,N_92);
nand U5017 (N_5017,N_412,N_4551);
or U5018 (N_5018,N_4608,N_4226);
and U5019 (N_5019,N_1030,N_3355);
nand U5020 (N_5020,N_2026,N_2476);
nor U5021 (N_5021,N_4437,N_4362);
and U5022 (N_5022,N_2836,N_2350);
or U5023 (N_5023,N_1986,N_3435);
nand U5024 (N_5024,N_1367,N_1570);
or U5025 (N_5025,N_2894,N_1733);
xnor U5026 (N_5026,N_3219,N_28);
and U5027 (N_5027,N_3945,N_3805);
and U5028 (N_5028,N_4397,N_482);
nand U5029 (N_5029,N_3457,N_3640);
nand U5030 (N_5030,N_4496,N_1089);
and U5031 (N_5031,N_2332,N_2290);
xnor U5032 (N_5032,N_1820,N_3532);
or U5033 (N_5033,N_4317,N_1215);
or U5034 (N_5034,N_4125,N_4550);
or U5035 (N_5035,N_3942,N_764);
nand U5036 (N_5036,N_2777,N_1095);
or U5037 (N_5037,N_2694,N_938);
nor U5038 (N_5038,N_1415,N_4773);
xor U5039 (N_5039,N_3345,N_2722);
or U5040 (N_5040,N_30,N_1689);
nor U5041 (N_5041,N_3315,N_3684);
xnor U5042 (N_5042,N_4053,N_4043);
nand U5043 (N_5043,N_4161,N_3719);
nand U5044 (N_5044,N_2518,N_4670);
xor U5045 (N_5045,N_1723,N_1546);
nand U5046 (N_5046,N_2526,N_4346);
or U5047 (N_5047,N_1746,N_2626);
xor U5048 (N_5048,N_1049,N_3371);
nor U5049 (N_5049,N_4477,N_3224);
or U5050 (N_5050,N_2662,N_1363);
and U5051 (N_5051,N_2843,N_1027);
nand U5052 (N_5052,N_3905,N_3973);
nor U5053 (N_5053,N_1348,N_3341);
and U5054 (N_5054,N_191,N_596);
nor U5055 (N_5055,N_2119,N_1845);
nand U5056 (N_5056,N_2774,N_158);
or U5057 (N_5057,N_4794,N_397);
and U5058 (N_5058,N_1405,N_2454);
or U5059 (N_5059,N_1867,N_3117);
and U5060 (N_5060,N_431,N_1561);
xnor U5061 (N_5061,N_1885,N_474);
nor U5062 (N_5062,N_144,N_4533);
xor U5063 (N_5063,N_1403,N_4997);
nand U5064 (N_5064,N_563,N_62);
nand U5065 (N_5065,N_3577,N_4588);
and U5066 (N_5066,N_4885,N_4776);
or U5067 (N_5067,N_1242,N_3077);
nor U5068 (N_5068,N_4790,N_324);
and U5069 (N_5069,N_4452,N_4425);
nand U5070 (N_5070,N_1001,N_503);
nor U5071 (N_5071,N_651,N_1019);
nor U5072 (N_5072,N_2109,N_125);
and U5073 (N_5073,N_3829,N_3308);
xor U5074 (N_5074,N_215,N_2433);
xor U5075 (N_5075,N_4430,N_340);
xnor U5076 (N_5076,N_2838,N_1855);
nand U5077 (N_5077,N_3575,N_1978);
nor U5078 (N_5078,N_4895,N_3116);
nand U5079 (N_5079,N_136,N_969);
nor U5080 (N_5080,N_4319,N_655);
or U5081 (N_5081,N_3204,N_361);
nand U5082 (N_5082,N_4916,N_511);
nand U5083 (N_5083,N_2315,N_1998);
nor U5084 (N_5084,N_2751,N_2001);
nor U5085 (N_5085,N_1268,N_864);
xnor U5086 (N_5086,N_4047,N_1209);
or U5087 (N_5087,N_4908,N_1518);
or U5088 (N_5088,N_1784,N_4574);
xor U5089 (N_5089,N_4180,N_1204);
or U5090 (N_5090,N_819,N_1525);
and U5091 (N_5091,N_1887,N_3843);
xor U5092 (N_5092,N_2708,N_1603);
or U5093 (N_5093,N_4591,N_3763);
xor U5094 (N_5094,N_2242,N_4386);
xnor U5095 (N_5095,N_430,N_942);
nor U5096 (N_5096,N_3239,N_2444);
or U5097 (N_5097,N_4927,N_755);
or U5098 (N_5098,N_1530,N_3418);
and U5099 (N_5099,N_2707,N_3434);
nand U5100 (N_5100,N_757,N_4489);
nor U5101 (N_5101,N_591,N_4966);
nand U5102 (N_5102,N_1829,N_3853);
or U5103 (N_5103,N_1811,N_3191);
and U5104 (N_5104,N_2912,N_3436);
nor U5105 (N_5105,N_4182,N_76);
nor U5106 (N_5106,N_4157,N_4858);
xor U5107 (N_5107,N_3320,N_1770);
xnor U5108 (N_5108,N_4594,N_2642);
nor U5109 (N_5109,N_3798,N_2314);
xor U5110 (N_5110,N_4914,N_4981);
nor U5111 (N_5111,N_4713,N_2849);
or U5112 (N_5112,N_2091,N_2850);
nand U5113 (N_5113,N_4953,N_3443);
and U5114 (N_5114,N_1282,N_1868);
or U5115 (N_5115,N_3807,N_2061);
nand U5116 (N_5116,N_2337,N_388);
nand U5117 (N_5117,N_4442,N_3503);
nor U5118 (N_5118,N_674,N_1053);
nand U5119 (N_5119,N_649,N_1864);
or U5120 (N_5120,N_4375,N_2171);
nand U5121 (N_5121,N_3878,N_3880);
and U5122 (N_5122,N_387,N_1543);
and U5123 (N_5123,N_3476,N_1915);
and U5124 (N_5124,N_1759,N_1951);
or U5125 (N_5125,N_2724,N_1743);
nor U5126 (N_5126,N_1709,N_2855);
nor U5127 (N_5127,N_604,N_4519);
and U5128 (N_5128,N_4417,N_1526);
or U5129 (N_5129,N_2846,N_337);
nand U5130 (N_5130,N_3721,N_2035);
nand U5131 (N_5131,N_790,N_4706);
nor U5132 (N_5132,N_3502,N_2220);
nor U5133 (N_5133,N_2267,N_4980);
xnor U5134 (N_5134,N_4006,N_4870);
nand U5135 (N_5135,N_2555,N_1054);
or U5136 (N_5136,N_4181,N_533);
nand U5137 (N_5137,N_1647,N_194);
nand U5138 (N_5138,N_2089,N_1732);
or U5139 (N_5139,N_3274,N_4286);
nor U5140 (N_5140,N_3005,N_167);
and U5141 (N_5141,N_2477,N_4612);
nand U5142 (N_5142,N_405,N_3910);
and U5143 (N_5143,N_3466,N_615);
nand U5144 (N_5144,N_3437,N_4145);
or U5145 (N_5145,N_732,N_1226);
xnor U5146 (N_5146,N_2151,N_4038);
nand U5147 (N_5147,N_776,N_4571);
nor U5148 (N_5148,N_3148,N_4129);
and U5149 (N_5149,N_4253,N_1057);
nand U5150 (N_5150,N_3470,N_3304);
or U5151 (N_5151,N_325,N_4617);
nor U5152 (N_5152,N_3190,N_1059);
or U5153 (N_5153,N_1581,N_57);
or U5154 (N_5154,N_235,N_3388);
xor U5155 (N_5155,N_1767,N_2686);
and U5156 (N_5156,N_3255,N_4839);
and U5157 (N_5157,N_4643,N_3967);
or U5158 (N_5158,N_908,N_4341);
and U5159 (N_5159,N_2182,N_2302);
or U5160 (N_5160,N_3100,N_498);
xnor U5161 (N_5161,N_4630,N_61);
nor U5162 (N_5162,N_546,N_2891);
and U5163 (N_5163,N_1630,N_2081);
or U5164 (N_5164,N_3273,N_2823);
or U5165 (N_5165,N_295,N_4788);
nand U5166 (N_5166,N_3481,N_1754);
nor U5167 (N_5167,N_1078,N_813);
nand U5168 (N_5168,N_464,N_1531);
nand U5169 (N_5169,N_839,N_4530);
nor U5170 (N_5170,N_3586,N_3644);
and U5171 (N_5171,N_565,N_401);
xor U5172 (N_5172,N_3562,N_2986);
or U5173 (N_5173,N_3520,N_4616);
or U5174 (N_5174,N_4208,N_2468);
nor U5175 (N_5175,N_1642,N_2558);
nor U5176 (N_5176,N_3695,N_1004);
nor U5177 (N_5177,N_1283,N_2588);
nor U5178 (N_5178,N_1039,N_2647);
nand U5179 (N_5179,N_901,N_582);
nand U5180 (N_5180,N_3073,N_1460);
and U5181 (N_5181,N_2591,N_1555);
nor U5182 (N_5182,N_2692,N_4779);
xnor U5183 (N_5183,N_1838,N_3856);
xor U5184 (N_5184,N_3797,N_4472);
and U5185 (N_5185,N_4158,N_2284);
xor U5186 (N_5186,N_4913,N_1610);
and U5187 (N_5187,N_1175,N_494);
nor U5188 (N_5188,N_3493,N_4810);
nand U5189 (N_5189,N_13,N_74);
or U5190 (N_5190,N_2861,N_2786);
or U5191 (N_5191,N_492,N_4451);
or U5192 (N_5192,N_3143,N_1097);
nor U5193 (N_5193,N_1150,N_4526);
xnor U5194 (N_5194,N_3333,N_303);
nor U5195 (N_5195,N_679,N_748);
nand U5196 (N_5196,N_4026,N_4761);
xor U5197 (N_5197,N_1858,N_1072);
nand U5198 (N_5198,N_3414,N_3523);
or U5199 (N_5199,N_3707,N_3722);
or U5200 (N_5200,N_1520,N_3011);
xnor U5201 (N_5201,N_4712,N_2784);
nand U5202 (N_5202,N_4553,N_1794);
xnor U5203 (N_5203,N_1317,N_2914);
nand U5204 (N_5204,N_4723,N_4032);
xor U5205 (N_5205,N_1933,N_4604);
nor U5206 (N_5206,N_838,N_3901);
nor U5207 (N_5207,N_3934,N_1645);
nand U5208 (N_5208,N_1582,N_4968);
or U5209 (N_5209,N_2699,N_1076);
xor U5210 (N_5210,N_2152,N_402);
or U5211 (N_5211,N_360,N_3761);
nor U5212 (N_5212,N_939,N_1967);
xnor U5213 (N_5213,N_876,N_3076);
or U5214 (N_5214,N_2601,N_2996);
or U5215 (N_5215,N_690,N_1437);
nor U5216 (N_5216,N_2259,N_1098);
nand U5217 (N_5217,N_3576,N_1745);
nand U5218 (N_5218,N_2319,N_2111);
or U5219 (N_5219,N_472,N_522);
xor U5220 (N_5220,N_50,N_2425);
or U5221 (N_5221,N_3758,N_1814);
or U5222 (N_5222,N_1708,N_4466);
xnor U5223 (N_5223,N_3166,N_4056);
nand U5224 (N_5224,N_2866,N_3032);
xor U5225 (N_5225,N_1073,N_4052);
xor U5226 (N_5226,N_2781,N_4900);
and U5227 (N_5227,N_72,N_4391);
nand U5228 (N_5228,N_1239,N_644);
or U5229 (N_5229,N_3969,N_1840);
nor U5230 (N_5230,N_4348,N_185);
nor U5231 (N_5231,N_173,N_4025);
and U5232 (N_5232,N_1693,N_1632);
or U5233 (N_5233,N_4146,N_2999);
xor U5234 (N_5234,N_2131,N_4474);
or U5235 (N_5235,N_1914,N_2192);
and U5236 (N_5236,N_465,N_4255);
xnor U5237 (N_5237,N_2787,N_4349);
and U5238 (N_5238,N_2973,N_237);
and U5239 (N_5239,N_4620,N_2056);
or U5240 (N_5240,N_1261,N_2978);
nand U5241 (N_5241,N_3785,N_4249);
nand U5242 (N_5242,N_4892,N_2103);
or U5243 (N_5243,N_1913,N_3107);
xor U5244 (N_5244,N_4429,N_416);
nand U5245 (N_5245,N_4316,N_1685);
and U5246 (N_5246,N_2712,N_4098);
nand U5247 (N_5247,N_1529,N_1199);
xor U5248 (N_5248,N_317,N_1850);
or U5249 (N_5249,N_1524,N_3213);
nand U5250 (N_5250,N_1222,N_886);
or U5251 (N_5251,N_4971,N_698);
and U5252 (N_5252,N_2434,N_250);
nor U5253 (N_5253,N_2196,N_4393);
and U5254 (N_5254,N_1122,N_4775);
xor U5255 (N_5255,N_259,N_3214);
nand U5256 (N_5256,N_3376,N_484);
nand U5257 (N_5257,N_1198,N_1277);
xnor U5258 (N_5258,N_1975,N_845);
or U5259 (N_5259,N_2253,N_4527);
or U5260 (N_5260,N_2416,N_4521);
nand U5261 (N_5261,N_481,N_4659);
nand U5262 (N_5262,N_460,N_4461);
nor U5263 (N_5263,N_3142,N_4860);
or U5264 (N_5264,N_1126,N_3555);
and U5265 (N_5265,N_2217,N_4201);
nor U5266 (N_5266,N_1756,N_4545);
and U5267 (N_5267,N_666,N_3492);
and U5268 (N_5268,N_1656,N_3459);
xnor U5269 (N_5269,N_4088,N_1139);
nand U5270 (N_5270,N_4213,N_4322);
nand U5271 (N_5271,N_2550,N_1876);
or U5272 (N_5272,N_2236,N_64);
or U5273 (N_5273,N_3625,N_1668);
xnor U5274 (N_5274,N_1965,N_2365);
xor U5275 (N_5275,N_3029,N_4045);
xnor U5276 (N_5276,N_2414,N_129);
nand U5277 (N_5277,N_4911,N_4566);
xnor U5278 (N_5278,N_641,N_396);
or U5279 (N_5279,N_1343,N_1103);
xor U5280 (N_5280,N_2869,N_310);
xnor U5281 (N_5281,N_3623,N_1295);
nor U5282 (N_5282,N_1163,N_599);
xnor U5283 (N_5283,N_3933,N_3280);
nor U5284 (N_5284,N_1451,N_2422);
and U5285 (N_5285,N_3017,N_643);
or U5286 (N_5286,N_2689,N_1187);
xor U5287 (N_5287,N_1003,N_1866);
or U5288 (N_5288,N_584,N_4217);
and U5289 (N_5289,N_3151,N_4347);
nor U5290 (N_5290,N_415,N_2481);
nand U5291 (N_5291,N_138,N_601);
and U5292 (N_5292,N_1022,N_1463);
nand U5293 (N_5293,N_2813,N_3086);
nor U5294 (N_5294,N_2521,N_2922);
and U5295 (N_5295,N_2055,N_1402);
and U5296 (N_5296,N_2616,N_798);
nor U5297 (N_5297,N_2547,N_4721);
or U5298 (N_5298,N_1556,N_1773);
xor U5299 (N_5299,N_103,N_4586);
nor U5300 (N_5300,N_1124,N_1425);
nor U5301 (N_5301,N_1002,N_2198);
and U5302 (N_5302,N_2760,N_2471);
xnor U5303 (N_5303,N_3711,N_2503);
xor U5304 (N_5304,N_4479,N_455);
or U5305 (N_5305,N_2505,N_3067);
and U5306 (N_5306,N_4114,N_3930);
xnor U5307 (N_5307,N_4421,N_1189);
xnor U5308 (N_5308,N_4887,N_4890);
and U5309 (N_5309,N_2445,N_1616);
xnor U5310 (N_5310,N_4613,N_1895);
and U5311 (N_5311,N_858,N_3387);
nand U5312 (N_5312,N_3847,N_3357);
and U5313 (N_5313,N_3679,N_4872);
nor U5314 (N_5314,N_1465,N_52);
xor U5315 (N_5315,N_1406,N_4599);
or U5316 (N_5316,N_831,N_181);
or U5317 (N_5317,N_3705,N_4705);
xor U5318 (N_5318,N_1737,N_2145);
and U5319 (N_5319,N_3757,N_268);
xnor U5320 (N_5320,N_2690,N_3051);
and U5321 (N_5321,N_1266,N_4378);
nor U5322 (N_5322,N_3646,N_1924);
xor U5323 (N_5323,N_4977,N_2679);
xor U5324 (N_5324,N_3920,N_3513);
and U5325 (N_5325,N_3461,N_2752);
nand U5326 (N_5326,N_1633,N_4809);
nand U5327 (N_5327,N_1422,N_2054);
nand U5328 (N_5328,N_1740,N_1516);
nand U5329 (N_5329,N_1532,N_1925);
xor U5330 (N_5330,N_998,N_1155);
nor U5331 (N_5331,N_60,N_283);
and U5332 (N_5332,N_4002,N_1486);
nand U5333 (N_5333,N_4439,N_3449);
and U5334 (N_5334,N_3530,N_4654);
nor U5335 (N_5335,N_1648,N_4500);
nor U5336 (N_5336,N_3423,N_97);
nand U5337 (N_5337,N_4287,N_956);
nand U5338 (N_5338,N_3653,N_4863);
and U5339 (N_5339,N_1397,N_462);
nand U5340 (N_5340,N_1123,N_1815);
and U5341 (N_5341,N_3028,N_2469);
or U5342 (N_5342,N_3702,N_3289);
nand U5343 (N_5343,N_1598,N_4131);
nand U5344 (N_5344,N_274,N_3821);
and U5345 (N_5345,N_2762,N_319);
xnor U5346 (N_5346,N_4112,N_2715);
and U5347 (N_5347,N_721,N_3645);
or U5348 (N_5348,N_1937,N_3656);
and U5349 (N_5349,N_3981,N_3346);
nor U5350 (N_5350,N_2256,N_1612);
and U5351 (N_5351,N_965,N_2807);
nor U5352 (N_5352,N_747,N_807);
nor U5353 (N_5353,N_2596,N_1843);
or U5354 (N_5354,N_442,N_2420);
nor U5355 (N_5355,N_1628,N_3671);
nor U5356 (N_5356,N_769,N_539);
nor U5357 (N_5357,N_4849,N_350);
and U5358 (N_5358,N_3216,N_701);
or U5359 (N_5359,N_4427,N_4751);
xnor U5360 (N_5360,N_3783,N_1835);
nor U5361 (N_5361,N_2143,N_2272);
xnor U5362 (N_5362,N_2254,N_4767);
nor U5363 (N_5363,N_1010,N_2308);
nand U5364 (N_5364,N_1842,N_1712);
nor U5365 (N_5365,N_977,N_266);
nor U5366 (N_5366,N_1786,N_2099);
xnor U5367 (N_5367,N_2878,N_2578);
xnor U5368 (N_5368,N_2400,N_3331);
nand U5369 (N_5369,N_3582,N_1990);
nand U5370 (N_5370,N_2666,N_2525);
nand U5371 (N_5371,N_3053,N_3710);
xnor U5372 (N_5372,N_2517,N_334);
and U5373 (N_5373,N_3339,N_1481);
and U5374 (N_5374,N_1623,N_3515);
and U5375 (N_5375,N_1228,N_1253);
and U5376 (N_5376,N_1025,N_3442);
xor U5377 (N_5377,N_1392,N_104);
and U5378 (N_5378,N_3013,N_621);
or U5379 (N_5379,N_2004,N_1020);
nand U5380 (N_5380,N_1017,N_3293);
and U5381 (N_5381,N_0,N_1901);
xnor U5382 (N_5382,N_3751,N_1651);
or U5383 (N_5383,N_1545,N_1903);
or U5384 (N_5384,N_3337,N_3560);
and U5385 (N_5385,N_2128,N_4110);
and U5386 (N_5386,N_4662,N_26);
nand U5387 (N_5387,N_2357,N_3329);
or U5388 (N_5388,N_3429,N_1075);
and U5389 (N_5389,N_2569,N_1479);
nand U5390 (N_5390,N_713,N_3698);
and U5391 (N_5391,N_4749,N_3902);
or U5392 (N_5392,N_986,N_867);
xnor U5393 (N_5393,N_1900,N_3736);
or U5394 (N_5394,N_801,N_2387);
xor U5395 (N_5395,N_2825,N_3178);
nor U5396 (N_5396,N_3729,N_2801);
or U5397 (N_5397,N_2375,N_2022);
and U5398 (N_5398,N_56,N_4948);
and U5399 (N_5399,N_3595,N_849);
nor U5400 (N_5400,N_1672,N_2120);
and U5401 (N_5401,N_2144,N_121);
and U5402 (N_5402,N_1236,N_4435);
nand U5403 (N_5403,N_4447,N_2757);
nand U5404 (N_5404,N_109,N_3439);
nand U5405 (N_5405,N_1781,N_2952);
and U5406 (N_5406,N_336,N_4066);
xor U5407 (N_5407,N_3034,N_1819);
and U5408 (N_5408,N_3629,N_2168);
nor U5409 (N_5409,N_4083,N_4577);
nand U5410 (N_5410,N_2079,N_1969);
nand U5411 (N_5411,N_4652,N_4564);
or U5412 (N_5412,N_4658,N_1064);
nor U5413 (N_5413,N_4988,N_1874);
xor U5414 (N_5414,N_3179,N_3536);
xnor U5415 (N_5415,N_352,N_2716);
nor U5416 (N_5416,N_2811,N_2135);
xnor U5417 (N_5417,N_3898,N_1775);
nor U5418 (N_5418,N_2816,N_2392);
and U5419 (N_5419,N_4982,N_857);
nor U5420 (N_5420,N_2459,N_654);
and U5421 (N_5421,N_3257,N_67);
nor U5422 (N_5422,N_3683,N_632);
and U5423 (N_5423,N_1580,N_1849);
or U5424 (N_5424,N_214,N_4744);
nor U5425 (N_5425,N_137,N_77);
or U5426 (N_5426,N_1094,N_4507);
or U5427 (N_5427,N_4314,N_2695);
nand U5428 (N_5428,N_3641,N_7);
and U5429 (N_5429,N_3860,N_1687);
nor U5430 (N_5430,N_4709,N_2335);
and U5431 (N_5431,N_3330,N_556);
or U5432 (N_5432,N_2396,N_2824);
xnor U5433 (N_5433,N_4491,N_2141);
and U5434 (N_5434,N_3480,N_4958);
nand U5435 (N_5435,N_3855,N_3411);
nand U5436 (N_5436,N_3496,N_3206);
or U5437 (N_5437,N_3205,N_3535);
xnor U5438 (N_5438,N_2584,N_1145);
xnor U5439 (N_5439,N_3614,N_2613);
nand U5440 (N_5440,N_4089,N_414);
or U5441 (N_5441,N_3174,N_3478);
xnor U5442 (N_5442,N_4768,N_404);
and U5443 (N_5443,N_3830,N_557);
xor U5444 (N_5444,N_1143,N_3064);
nand U5445 (N_5445,N_2020,N_3781);
nand U5446 (N_5446,N_1158,N_3563);
nand U5447 (N_5447,N_909,N_3448);
xnor U5448 (N_5448,N_2687,N_630);
nand U5449 (N_5449,N_3431,N_4311);
or U5450 (N_5450,N_4410,N_631);
xor U5451 (N_5451,N_1440,N_2260);
nor U5452 (N_5452,N_182,N_2472);
or U5453 (N_5453,N_3673,N_410);
nand U5454 (N_5454,N_227,N_90);
or U5455 (N_5455,N_3774,N_2639);
nor U5456 (N_5456,N_151,N_4372);
or U5457 (N_5457,N_855,N_4148);
and U5458 (N_5458,N_1350,N_4504);
and U5459 (N_5459,N_33,N_3170);
xor U5460 (N_5460,N_3324,N_1673);
nor U5461 (N_5461,N_4832,N_2175);
or U5462 (N_5462,N_2565,N_4034);
nor U5463 (N_5463,N_3229,N_131);
or U5464 (N_5464,N_201,N_2998);
and U5465 (N_5465,N_1188,N_1167);
nand U5466 (N_5466,N_988,N_2102);
nor U5467 (N_5467,N_25,N_4626);
and U5468 (N_5468,N_1265,N_2432);
and U5469 (N_5469,N_4358,N_1141);
and U5470 (N_5470,N_1857,N_4937);
and U5471 (N_5471,N_2710,N_2863);
and U5472 (N_5472,N_198,N_459);
nand U5473 (N_5473,N_683,N_2268);
nor U5474 (N_5474,N_257,N_4306);
xor U5475 (N_5475,N_2541,N_510);
nand U5476 (N_5476,N_963,N_4944);
xnor U5477 (N_5477,N_15,N_2147);
and U5478 (N_5478,N_4882,N_2788);
nand U5479 (N_5479,N_3144,N_2017);
or U5480 (N_5480,N_765,N_1861);
nand U5481 (N_5481,N_1551,N_2595);
xor U5482 (N_5482,N_2096,N_3887);
nand U5483 (N_5483,N_1184,N_1621);
and U5484 (N_5484,N_3718,N_2785);
nor U5485 (N_5485,N_1413,N_991);
xor U5486 (N_5486,N_1875,N_937);
or U5487 (N_5487,N_242,N_2614);
nand U5488 (N_5488,N_1462,N_2174);
nor U5489 (N_5489,N_1575,N_1488);
nand U5490 (N_5490,N_4576,N_4587);
or U5491 (N_5491,N_323,N_1583);
and U5492 (N_5492,N_3591,N_2919);
and U5493 (N_5493,N_3579,N_1935);
and U5494 (N_5494,N_68,N_1504);
nor U5495 (N_5495,N_2768,N_1641);
and U5496 (N_5496,N_4414,N_3734);
or U5497 (N_5497,N_4544,N_2435);
nand U5498 (N_5498,N_1663,N_3176);
or U5499 (N_5499,N_2516,N_1506);
nand U5500 (N_5500,N_3771,N_3959);
nor U5501 (N_5501,N_3343,N_200);
nand U5502 (N_5502,N_366,N_24);
xnor U5503 (N_5503,N_4476,N_285);
and U5504 (N_5504,N_284,N_4019);
or U5505 (N_5505,N_1982,N_4669);
xor U5506 (N_5506,N_3940,N_124);
or U5507 (N_5507,N_2191,N_4419);
xnor U5508 (N_5508,N_3160,N_2234);
nor U5509 (N_5509,N_495,N_810);
or U5510 (N_5510,N_4134,N_3351);
xnor U5511 (N_5511,N_3003,N_2053);
and U5512 (N_5512,N_2605,N_2250);
nand U5513 (N_5513,N_3183,N_3222);
nor U5514 (N_5514,N_2510,N_4815);
nor U5515 (N_5515,N_3082,N_4864);
nor U5516 (N_5516,N_3420,N_1063);
nor U5517 (N_5517,N_2833,N_638);
nor U5518 (N_5518,N_3398,N_3927);
xor U5519 (N_5519,N_3688,N_4408);
and U5520 (N_5520,N_466,N_1217);
nand U5521 (N_5521,N_1036,N_3740);
nand U5522 (N_5522,N_3118,N_1498);
or U5523 (N_5523,N_110,N_4869);
and U5524 (N_5524,N_3624,N_394);
xnor U5525 (N_5525,N_229,N_1664);
and U5526 (N_5526,N_620,N_2301);
xor U5527 (N_5527,N_3739,N_2743);
nand U5528 (N_5528,N_3392,N_3592);
nor U5529 (N_5529,N_4581,N_58);
and U5530 (N_5530,N_4797,N_702);
xor U5531 (N_5531,N_2670,N_554);
nor U5532 (N_5532,N_746,N_1503);
nor U5533 (N_5533,N_2502,N_787);
xnor U5534 (N_5534,N_2277,N_4678);
or U5535 (N_5535,N_817,N_293);
nand U5536 (N_5536,N_935,N_949);
nor U5537 (N_5537,N_2625,N_850);
and U5538 (N_5538,N_1591,N_3413);
or U5539 (N_5539,N_1607,N_3567);
or U5540 (N_5540,N_355,N_2534);
nor U5541 (N_5541,N_3716,N_432);
or U5542 (N_5542,N_3991,N_2431);
nor U5543 (N_5543,N_1361,N_3277);
or U5544 (N_5544,N_4122,N_436);
xor U5545 (N_5545,N_2490,N_2876);
nand U5546 (N_5546,N_3680,N_3909);
nand U5547 (N_5547,N_3796,N_3726);
nand U5548 (N_5548,N_2819,N_256);
and U5549 (N_5549,N_2736,N_1917);
or U5550 (N_5550,N_1107,N_3792);
and U5551 (N_5551,N_3382,N_2621);
xnor U5552 (N_5552,N_4628,N_1172);
and U5553 (N_5553,N_2222,N_4693);
or U5554 (N_5554,N_2430,N_4061);
and U5555 (N_5555,N_3676,N_4755);
and U5556 (N_5556,N_753,N_1256);
nor U5557 (N_5557,N_2631,N_1216);
or U5558 (N_5558,N_2489,N_330);
nor U5559 (N_5559,N_2654,N_3596);
or U5560 (N_5560,N_1777,N_1300);
and U5561 (N_5561,N_3831,N_3033);
and U5562 (N_5562,N_204,N_1106);
xnor U5563 (N_5563,N_1860,N_126);
nor U5564 (N_5564,N_3039,N_1267);
and U5565 (N_5565,N_4058,N_3342);
xnor U5566 (N_5566,N_735,N_3960);
or U5567 (N_5567,N_4099,N_3199);
or U5568 (N_5568,N_2466,N_3338);
nand U5569 (N_5569,N_4298,N_426);
or U5570 (N_5570,N_4862,N_3068);
and U5571 (N_5571,N_1194,N_4030);
nor U5572 (N_5572,N_4200,N_2165);
xor U5573 (N_5573,N_2951,N_4499);
and U5574 (N_5574,N_3639,N_4510);
xor U5575 (N_5575,N_4730,N_1905);
nand U5576 (N_5576,N_684,N_3088);
xnor U5577 (N_5577,N_2665,N_1891);
xnor U5578 (N_5578,N_3922,N_2336);
or U5579 (N_5579,N_282,N_2049);
nand U5580 (N_5580,N_2697,N_841);
nor U5581 (N_5581,N_4737,N_2040);
and U5582 (N_5582,N_4187,N_3265);
and U5583 (N_5583,N_1945,N_4851);
nor U5584 (N_5584,N_970,N_3966);
or U5585 (N_5585,N_2372,N_2052);
xor U5586 (N_5586,N_2252,N_2566);
or U5587 (N_5587,N_1297,N_661);
xor U5588 (N_5588,N_4004,N_1542);
nand U5589 (N_5589,N_2457,N_4436);
xnor U5590 (N_5590,N_170,N_47);
nand U5591 (N_5591,N_2470,N_1650);
and U5592 (N_5592,N_716,N_3877);
nor U5593 (N_5593,N_708,N_3074);
and U5594 (N_5594,N_4135,N_3424);
and U5595 (N_5595,N_3799,N_3926);
or U5596 (N_5596,N_4901,N_1475);
xnor U5597 (N_5597,N_4722,N_3544);
or U5598 (N_5598,N_4090,N_4891);
and U5599 (N_5599,N_2064,N_3745);
xnor U5600 (N_5600,N_1159,N_4460);
or U5601 (N_5601,N_2636,N_2772);
nand U5602 (N_5602,N_264,N_4656);
or U5603 (N_5603,N_659,N_3123);
or U5604 (N_5604,N_4528,N_730);
or U5605 (N_5605,N_758,N_4936);
nor U5606 (N_5606,N_1806,N_1494);
and U5607 (N_5607,N_4542,N_5);
or U5608 (N_5608,N_3234,N_1589);
nand U5609 (N_5609,N_4492,N_4536);
or U5610 (N_5610,N_3869,N_315);
and U5611 (N_5611,N_2649,N_800);
and U5612 (N_5612,N_3616,N_2016);
xor U5613 (N_5613,N_626,N_869);
or U5614 (N_5614,N_842,N_1438);
or U5615 (N_5615,N_3801,N_2948);
and U5616 (N_5616,N_2727,N_3093);
xnor U5617 (N_5617,N_4299,N_3728);
xor U5618 (N_5618,N_3814,N_3677);
nand U5619 (N_5619,N_2493,N_1595);
nand U5620 (N_5620,N_3057,N_2546);
or U5621 (N_5621,N_667,N_3662);
nor U5622 (N_5622,N_4018,N_4423);
and U5623 (N_5623,N_3248,N_1971);
xnor U5624 (N_5624,N_3889,N_4784);
nand U5625 (N_5625,N_4711,N_4609);
xnor U5626 (N_5626,N_4303,N_2070);
nor U5627 (N_5627,N_2374,N_3775);
nor U5628 (N_5628,N_1444,N_302);
nor U5629 (N_5629,N_2180,N_4482);
nor U5630 (N_5630,N_4740,N_3950);
nor U5631 (N_5631,N_663,N_4123);
nand U5632 (N_5632,N_4902,N_3670);
or U5633 (N_5633,N_3501,N_4219);
or U5634 (N_5634,N_1210,N_4242);
or U5635 (N_5635,N_3773,N_4331);
nand U5636 (N_5636,N_4363,N_545);
nand U5637 (N_5637,N_1062,N_4789);
xor U5638 (N_5638,N_3506,N_4153);
nand U5639 (N_5639,N_1752,N_3915);
and U5640 (N_5640,N_4277,N_3464);
nor U5641 (N_5641,N_660,N_2610);
and U5642 (N_5642,N_1015,N_1102);
nor U5643 (N_5643,N_1390,N_1567);
xnor U5644 (N_5644,N_1453,N_1372);
nand U5645 (N_5645,N_2644,N_3161);
and U5646 (N_5646,N_4736,N_811);
xnor U5647 (N_5647,N_2840,N_4569);
and U5648 (N_5648,N_3340,N_3512);
nand U5649 (N_5649,N_3169,N_4904);
or U5650 (N_5650,N_2248,N_1890);
nor U5651 (N_5651,N_4385,N_2391);
nand U5652 (N_5652,N_3403,N_3390);
or U5653 (N_5653,N_933,N_1896);
xnor U5654 (N_5654,N_289,N_2497);
nand U5655 (N_5655,N_832,N_3900);
or U5656 (N_5656,N_945,N_3911);
nor U5657 (N_5657,N_647,N_1250);
or U5658 (N_5658,N_3356,N_3894);
or U5659 (N_5659,N_847,N_947);
or U5660 (N_5660,N_915,N_4449);
nand U5661 (N_5661,N_3007,N_2674);
xnor U5662 (N_5662,N_1690,N_2632);
xor U5663 (N_5663,N_878,N_2366);
nand U5664 (N_5664,N_1243,N_1130);
or U5665 (N_5665,N_3181,N_3301);
nand U5666 (N_5666,N_884,N_4484);
nor U5667 (N_5667,N_4538,N_1597);
nand U5668 (N_5668,N_3008,N_978);
and U5669 (N_5669,N_1902,N_1264);
xor U5670 (N_5670,N_4493,N_2559);
xor U5671 (N_5671,N_4610,N_2058);
xnor U5672 (N_5672,N_341,N_3870);
nand U5673 (N_5673,N_1499,N_2602);
nor U5674 (N_5674,N_1544,N_3402);
xnor U5675 (N_5675,N_4109,N_477);
and U5676 (N_5676,N_3899,N_3733);
and U5677 (N_5677,N_2508,N_4402);
or U5678 (N_5678,N_2002,N_1326);
and U5679 (N_5679,N_189,N_3606);
or U5680 (N_5680,N_1493,N_4893);
xnor U5681 (N_5681,N_729,N_4837);
or U5682 (N_5682,N_3583,N_1371);
nand U5683 (N_5683,N_1869,N_203);
and U5684 (N_5684,N_4930,N_3394);
nor U5685 (N_5685,N_3534,N_792);
nand U5686 (N_5686,N_4934,N_4495);
and U5687 (N_5687,N_1149,N_524);
xnor U5688 (N_5688,N_4165,N_1412);
nand U5689 (N_5689,N_3026,N_3238);
xor U5690 (N_5690,N_2795,N_4805);
and U5691 (N_5691,N_3790,N_809);
nor U5692 (N_5692,N_1470,N_1110);
or U5693 (N_5693,N_1823,N_1259);
xnor U5694 (N_5694,N_347,N_433);
or U5695 (N_5695,N_3095,N_1703);
nor U5696 (N_5696,N_907,N_4539);
and U5697 (N_5697,N_3935,N_4563);
nand U5698 (N_5698,N_3727,N_4054);
nand U5699 (N_5699,N_4621,N_4238);
nor U5700 (N_5700,N_4448,N_444);
and U5701 (N_5701,N_4956,N_3044);
nor U5702 (N_5702,N_874,N_3198);
nor U5703 (N_5703,N_1813,N_1791);
nand U5704 (N_5704,N_3322,N_4195);
and U5705 (N_5705,N_1321,N_1325);
or U5706 (N_5706,N_2887,N_2834);
nor U5707 (N_5707,N_3133,N_1093);
and U5708 (N_5708,N_3553,N_1090);
or U5709 (N_5709,N_2815,N_476);
and U5710 (N_5710,N_1452,N_3405);
or U5711 (N_5711,N_625,N_2123);
nor U5712 (N_5712,N_3030,N_2734);
nor U5713 (N_5713,N_2413,N_3747);
nand U5714 (N_5714,N_4697,N_2100);
nor U5715 (N_5715,N_2395,N_2479);
nor U5716 (N_5716,N_544,N_3141);
nand U5717 (N_5717,N_3245,N_2945);
and U5718 (N_5718,N_3070,N_914);
xor U5719 (N_5719,N_3916,N_1278);
nand U5720 (N_5720,N_1286,N_3835);
nand U5721 (N_5721,N_2359,N_140);
xor U5722 (N_5722,N_4861,N_4434);
nand U5723 (N_5723,N_1622,N_3997);
xor U5724 (N_5724,N_2225,N_4585);
xnor U5725 (N_5725,N_1354,N_4830);
nand U5726 (N_5726,N_3743,N_3412);
nor U5727 (N_5727,N_3119,N_1411);
and U5728 (N_5728,N_3021,N_4280);
or U5729 (N_5729,N_1554,N_3284);
nand U5730 (N_5730,N_4672,N_307);
xnor U5731 (N_5731,N_4633,N_3776);
xnor U5732 (N_5732,N_3958,N_4921);
nand U5733 (N_5733,N_1922,N_4124);
and U5734 (N_5734,N_440,N_662);
or U5735 (N_5735,N_834,N_4735);
and U5736 (N_5736,N_1798,N_2536);
nor U5737 (N_5737,N_2381,N_1018);
nor U5738 (N_5738,N_1404,N_3929);
and U5739 (N_5739,N_3804,N_1851);
xor U5740 (N_5740,N_2449,N_881);
xor U5741 (N_5741,N_2126,N_944);
nand U5742 (N_5742,N_311,N_4687);
nand U5743 (N_5743,N_425,N_2025);
and U5744 (N_5744,N_1456,N_294);
xor U5745 (N_5745,N_2465,N_2832);
xnor U5746 (N_5746,N_2890,N_1964);
or U5747 (N_5747,N_575,N_4540);
and U5748 (N_5748,N_3243,N_1302);
or U5749 (N_5749,N_4468,N_4325);
and U5750 (N_5750,N_3789,N_2188);
or U5751 (N_5751,N_560,N_1537);
or U5752 (N_5752,N_1638,N_3613);
nor U5753 (N_5753,N_1557,N_4486);
or U5754 (N_5754,N_2388,N_316);
and U5755 (N_5755,N_1249,N_2748);
nand U5756 (N_5756,N_3965,N_1692);
nor U5757 (N_5757,N_4438,N_2997);
nor U5758 (N_5758,N_4568,N_3720);
nand U5759 (N_5759,N_736,N_4689);
xnor U5760 (N_5760,N_1016,N_1118);
nand U5761 (N_5761,N_3813,N_1197);
xnor U5762 (N_5762,N_3874,N_4817);
nor U5763 (N_5763,N_1445,N_290);
and U5764 (N_5764,N_984,N_338);
xnor U5765 (N_5765,N_4251,N_979);
xnor U5766 (N_5766,N_127,N_2221);
or U5767 (N_5767,N_2275,N_4193);
xnor U5768 (N_5768,N_339,N_4624);
and U5769 (N_5769,N_4879,N_1008);
xor U5770 (N_5770,N_2946,N_4007);
xnor U5771 (N_5771,N_2215,N_4388);
nor U5772 (N_5772,N_1576,N_3686);
nand U5773 (N_5773,N_1579,N_3299);
xor U5774 (N_5774,N_1378,N_4188);
and U5775 (N_5775,N_1340,N_3659);
or U5776 (N_5776,N_3767,N_4204);
nor U5777 (N_5777,N_3842,N_3681);
xor U5778 (N_5778,N_2261,N_2122);
or U5779 (N_5779,N_4638,N_941);
or U5780 (N_5780,N_3187,N_4288);
nand U5781 (N_5781,N_3528,N_2288);
nand U5782 (N_5782,N_2167,N_3578);
or U5783 (N_5783,N_55,N_2691);
nand U5784 (N_5784,N_3895,N_435);
and U5785 (N_5785,N_1047,N_3287);
nor U5786 (N_5786,N_1596,N_2618);
xor U5787 (N_5787,N_1368,N_2138);
nand U5788 (N_5788,N_549,N_3759);
xor U5789 (N_5789,N_2725,N_3924);
xor U5790 (N_5790,N_2829,N_1881);
or U5791 (N_5791,N_1035,N_1337);
nor U5792 (N_5792,N_3527,N_4263);
and U5793 (N_5793,N_3079,N_1783);
or U5794 (N_5794,N_3432,N_1620);
nor U5795 (N_5795,N_1571,N_2065);
and U5796 (N_5796,N_1161,N_2873);
xnor U5797 (N_5797,N_3628,N_3742);
nor U5798 (N_5798,N_3019,N_4967);
or U5799 (N_5799,N_1559,N_2617);
or U5800 (N_5800,N_4963,N_1353);
or U5801 (N_5801,N_923,N_4445);
and U5802 (N_5802,N_3669,N_378);
or U5803 (N_5803,N_1790,N_1751);
or U5804 (N_5804,N_1240,N_2418);
or U5805 (N_5805,N_1590,N_1185);
nor U5806 (N_5806,N_2354,N_1682);
xnor U5807 (N_5807,N_4237,N_4856);
nand U5808 (N_5808,N_120,N_1893);
xnor U5809 (N_5809,N_1844,N_4619);
xnor U5810 (N_5810,N_1789,N_902);
nand U5811 (N_5811,N_1852,N_572);
nor U5812 (N_5812,N_236,N_2028);
and U5813 (N_5813,N_2334,N_3602);
xor U5814 (N_5814,N_46,N_1088);
or U5815 (N_5815,N_705,N_2966);
and U5816 (N_5816,N_4073,N_719);
nand U5817 (N_5817,N_1505,N_779);
xor U5818 (N_5818,N_4985,N_4690);
and U5819 (N_5819,N_4481,N_4300);
nor U5820 (N_5820,N_450,N_1087);
and U5821 (N_5821,N_4411,N_222);
and U5822 (N_5822,N_172,N_2226);
and U5823 (N_5823,N_4235,N_3565);
nand U5824 (N_5824,N_2342,N_3682);
and U5825 (N_5825,N_4745,N_304);
xnor U5826 (N_5826,N_95,N_4261);
and U5827 (N_5827,N_561,N_2330);
and U5828 (N_5828,N_2276,N_1566);
nor U5829 (N_5829,N_368,N_3986);
xor U5830 (N_5830,N_2607,N_2353);
and U5831 (N_5831,N_4868,N_760);
nand U5832 (N_5832,N_1801,N_2299);
xor U5833 (N_5833,N_1448,N_2346);
xnor U5834 (N_5834,N_1995,N_1454);
and U5835 (N_5835,N_2717,N_4698);
and U5836 (N_5836,N_1702,N_4040);
or U5837 (N_5837,N_3025,N_1023);
nor U5838 (N_5838,N_1474,N_2186);
xor U5839 (N_5839,N_2352,N_4546);
nor U5840 (N_5840,N_868,N_83);
xor U5841 (N_5841,N_2044,N_4822);
nand U5842 (N_5842,N_1356,N_4726);
or U5843 (N_5843,N_4174,N_2461);
and U5844 (N_5844,N_3155,N_1058);
and U5845 (N_5845,N_1979,N_1771);
xor U5846 (N_5846,N_4172,N_4912);
or U5847 (N_5847,N_4144,N_1691);
nor U5848 (N_5848,N_216,N_3366);
and U5849 (N_5849,N_1136,N_493);
xnor U5850 (N_5850,N_2940,N_767);
nand U5851 (N_5851,N_990,N_2938);
nor U5852 (N_5852,N_2671,N_3865);
nor U5853 (N_5853,N_210,N_4673);
nand U5854 (N_5854,N_4320,N_3631);
nand U5855 (N_5855,N_871,N_4329);
and U5856 (N_5856,N_2121,N_489);
nor U5857 (N_5857,N_885,N_3651);
xnor U5858 (N_5858,N_362,N_712);
xnor U5859 (N_5859,N_3401,N_1931);
nor U5860 (N_5860,N_919,N_1347);
nor U5861 (N_5861,N_42,N_2498);
nor U5862 (N_5862,N_911,N_4718);
xor U5863 (N_5863,N_3438,N_1886);
nor U5864 (N_5864,N_1700,N_3791);
nand U5865 (N_5865,N_2305,N_1918);
nor U5866 (N_5866,N_826,N_4694);
xnor U5867 (N_5867,N_1152,N_2901);
xnor U5868 (N_5868,N_1067,N_1521);
nor U5869 (N_5869,N_569,N_3168);
and U5870 (N_5870,N_2942,N_2961);
nor U5871 (N_5871,N_3989,N_877);
nor U5872 (N_5872,N_4812,N_1223);
nor U5873 (N_5873,N_4183,N_896);
or U5874 (N_5874,N_3475,N_89);
nand U5875 (N_5875,N_3001,N_3139);
nor U5876 (N_5876,N_3648,N_2746);
and U5877 (N_5877,N_4142,N_786);
or U5878 (N_5878,N_4607,N_1170);
xor U5879 (N_5879,N_4149,N_3200);
nor U5880 (N_5880,N_3888,N_1731);
and U5881 (N_5881,N_2970,N_1833);
and U5882 (N_5882,N_4297,N_4302);
or U5883 (N_5883,N_1082,N_4478);
xnor U5884 (N_5884,N_4108,N_4295);
and U5885 (N_5885,N_2106,N_2513);
xor U5886 (N_5886,N_2892,N_276);
nor U5887 (N_5887,N_2417,N_2057);
or U5888 (N_5888,N_2719,N_2380);
and U5889 (N_5889,N_1889,N_3864);
or U5890 (N_5890,N_4756,N_4367);
nor U5891 (N_5891,N_1536,N_3833);
nand U5892 (N_5892,N_1328,N_731);
nor U5893 (N_5893,N_2295,N_1509);
or U5894 (N_5894,N_3953,N_581);
and U5895 (N_5895,N_4014,N_2447);
xor U5896 (N_5896,N_4383,N_1148);
and U5897 (N_5897,N_1332,N_2628);
xnor U5898 (N_5898,N_955,N_4380);
nand U5899 (N_5899,N_1640,N_1748);
or U5900 (N_5900,N_66,N_3724);
nand U5901 (N_5901,N_1677,N_69);
xnor U5902 (N_5902,N_1074,N_3794);
nand U5903 (N_5903,N_4150,N_2810);
or U5904 (N_5904,N_4192,N_162);
and U5905 (N_5905,N_1084,N_3164);
nor U5906 (N_5906,N_3358,N_1705);
nand U5907 (N_5907,N_4106,N_1879);
xor U5908 (N_5908,N_1480,N_2067);
and U5909 (N_5909,N_4457,N_1911);
xnor U5910 (N_5910,N_4850,N_3539);
and U5911 (N_5911,N_1387,N_3207);
nor U5912 (N_5912,N_3597,N_4688);
or U5913 (N_5913,N_733,N_1179);
or U5914 (N_5914,N_3753,N_1684);
or U5915 (N_5915,N_1573,N_4770);
and U5916 (N_5916,N_1338,N_4096);
nor U5917 (N_5917,N_4947,N_3867);
xnor U5918 (N_5918,N_2769,N_2529);
nand U5919 (N_5919,N_3931,N_1281);
nor U5920 (N_5920,N_4801,N_512);
nand U5921 (N_5921,N_815,N_3550);
nor U5922 (N_5922,N_547,N_598);
and U5923 (N_5923,N_4289,N_872);
xor U5924 (N_5924,N_2895,N_1883);
nor U5925 (N_5925,N_4923,N_1096);
nand U5926 (N_5926,N_875,N_1165);
xor U5927 (N_5927,N_4352,N_4074);
nand U5928 (N_5928,N_1816,N_574);
and U5929 (N_5929,N_177,N_406);
and U5930 (N_5930,N_759,N_1288);
and U5931 (N_5931,N_1502,N_2638);
nor U5932 (N_5932,N_1360,N_4248);
xnor U5933 (N_5933,N_2925,N_288);
nand U5934 (N_5934,N_2556,N_2977);
and U5935 (N_5935,N_3165,N_1882);
and U5936 (N_5936,N_1310,N_4178);
and U5937 (N_5937,N_2473,N_488);
or U5938 (N_5938,N_1201,N_4166);
nand U5939 (N_5939,N_1948,N_4381);
and U5940 (N_5940,N_4351,N_4748);
xnor U5941 (N_5941,N_1963,N_4884);
xnor U5942 (N_5942,N_4704,N_3072);
nand U5943 (N_5943,N_332,N_3225);
nand U5944 (N_5944,N_4044,N_2867);
and U5945 (N_5945,N_169,N_3643);
xnor U5946 (N_5946,N_2586,N_3441);
xnor U5947 (N_5947,N_2797,N_3521);
nor U5948 (N_5948,N_2851,N_1710);
xor U5949 (N_5949,N_3802,N_2105);
xnor U5950 (N_5950,N_4078,N_852);
and U5951 (N_5951,N_2291,N_4312);
and U5952 (N_5952,N_2729,N_4989);
or U5953 (N_5953,N_3035,N_364);
and U5954 (N_5954,N_840,N_3211);
or U5955 (N_5955,N_2920,N_2229);
and U5956 (N_5956,N_3159,N_3760);
xor U5957 (N_5957,N_1308,N_4197);
nor U5958 (N_5958,N_1005,N_1983);
xor U5959 (N_5959,N_1809,N_1846);
nand U5960 (N_5960,N_4095,N_3195);
or U5961 (N_5961,N_1836,N_804);
nand U5962 (N_5962,N_357,N_3717);
nand U5963 (N_5963,N_2376,N_1627);
xnor U5964 (N_5964,N_183,N_682);
xor U5965 (N_5965,N_2037,N_2763);
nand U5966 (N_5966,N_3556,N_1830);
xnor U5967 (N_5967,N_846,N_749);
nand U5968 (N_5968,N_1383,N_3561);
or U5969 (N_5969,N_1810,N_3819);
and U5970 (N_5970,N_1450,N_2176);
or U5971 (N_5971,N_4949,N_4854);
nand U5972 (N_5972,N_4513,N_2251);
xnor U5973 (N_5973,N_417,N_343);
xor U5974 (N_5974,N_1660,N_3630);
and U5975 (N_5975,N_2701,N_4220);
or U5976 (N_5976,N_3611,N_2545);
and U5977 (N_5977,N_1296,N_4919);
nand U5978 (N_5978,N_2663,N_1694);
nand U5979 (N_5979,N_1698,N_2538);
xnor U5980 (N_5980,N_2738,N_2693);
xor U5981 (N_5981,N_2676,N_4759);
and U5982 (N_5982,N_3278,N_3875);
xnor U5983 (N_5983,N_3,N_327);
and U5984 (N_5984,N_2574,N_3456);
xor U5985 (N_5985,N_862,N_3474);
and U5986 (N_5986,N_4206,N_2680);
nand U5987 (N_5987,N_318,N_3552);
nand U5988 (N_5988,N_328,N_624);
and U5989 (N_5989,N_3296,N_1248);
or U5990 (N_5990,N_3125,N_4326);
and U5991 (N_5991,N_1662,N_527);
nor U5992 (N_5992,N_4232,N_4813);
xnor U5993 (N_5993,N_3321,N_2185);
and U5994 (N_5994,N_4342,N_1469);
or U5995 (N_5995,N_4037,N_156);
nand U5996 (N_5996,N_3173,N_2077);
and U5997 (N_5997,N_4853,N_570);
nor U5998 (N_5998,N_2101,N_386);
xnor U5999 (N_5999,N_1029,N_188);
nor U6000 (N_6000,N_2562,N_38);
xnor U6001 (N_6001,N_2886,N_3317);
xnor U6002 (N_6002,N_4243,N_2909);
and U6003 (N_6003,N_2620,N_3419);
and U6004 (N_6004,N_4196,N_1907);
xor U6005 (N_6005,N_954,N_4294);
xnor U6006 (N_6006,N_3518,N_2913);
nor U6007 (N_6007,N_812,N_3097);
xor U6008 (N_6008,N_616,N_79);
xnor U6009 (N_6009,N_4440,N_199);
nand U6010 (N_6010,N_2487,N_4816);
xor U6011 (N_6011,N_3145,N_1626);
xnor U6012 (N_6012,N_3655,N_3533);
xnor U6013 (N_6013,N_4506,N_1606);
or U6014 (N_6014,N_490,N_202);
nand U6015 (N_6015,N_452,N_3319);
nor U6016 (N_6016,N_2113,N_3416);
nor U6017 (N_6017,N_2249,N_3422);
nor U6018 (N_6018,N_63,N_1091);
nand U6019 (N_6019,N_159,N_197);
nand U6020 (N_6020,N_2227,N_3816);
xor U6021 (N_6021,N_657,N_2358);
nand U6022 (N_6022,N_1323,N_4646);
xor U6023 (N_6023,N_2439,N_161);
nor U6024 (N_6024,N_3226,N_4055);
nand U6025 (N_6025,N_3447,N_1208);
or U6026 (N_6026,N_689,N_4842);
nor U6027 (N_6027,N_112,N_2075);
xor U6028 (N_6028,N_3451,N_4184);
or U6029 (N_6029,N_1287,N_724);
and U6030 (N_6030,N_142,N_2911);
xor U6031 (N_6031,N_3952,N_4211);
nand U6032 (N_6032,N_4935,N_2594);
xnor U6033 (N_6033,N_1930,N_1376);
or U6034 (N_6034,N_1138,N_4844);
xnor U6035 (N_6035,N_1683,N_1449);
xor U6036 (N_6036,N_722,N_957);
nand U6037 (N_6037,N_291,N_3499);
nor U6038 (N_6038,N_1635,N_595);
nor U6039 (N_6039,N_418,N_1322);
and U6040 (N_6040,N_3918,N_1237);
nor U6041 (N_6041,N_1056,N_1120);
and U6042 (N_6042,N_4752,N_744);
and U6043 (N_6043,N_1021,N_4580);
or U6044 (N_6044,N_2910,N_4855);
nand U6045 (N_6045,N_2202,N_3004);
nand U6046 (N_6046,N_4834,N_374);
and U6047 (N_6047,N_2818,N_1327);
and U6048 (N_6048,N_14,N_1319);
nand U6049 (N_6049,N_617,N_4806);
and U6050 (N_6050,N_4234,N_3291);
nand U6051 (N_6051,N_3167,N_3668);
or U6052 (N_6052,N_4023,N_1034);
nand U6053 (N_6053,N_4473,N_2187);
and U6054 (N_6054,N_3665,N_1472);
nand U6055 (N_6055,N_2172,N_1961);
or U6056 (N_6056,N_3840,N_4105);
and U6057 (N_6057,N_2223,N_3913);
nand U6058 (N_6058,N_3078,N_1426);
xor U6059 (N_6059,N_3311,N_2362);
nand U6060 (N_6060,N_4077,N_797);
or U6061 (N_6061,N_1496,N_3851);
xnor U6062 (N_6062,N_1292,N_806);
nand U6063 (N_6063,N_711,N_835);
nand U6064 (N_6064,N_398,N_3858);
and U6065 (N_6065,N_791,N_4081);
nor U6066 (N_6066,N_84,N_1517);
xor U6067 (N_6067,N_3465,N_4771);
and U6068 (N_6068,N_171,N_652);
or U6069 (N_6069,N_4596,N_4198);
xnor U6070 (N_6070,N_1817,N_3247);
or U6071 (N_6071,N_4462,N_4772);
xnor U6072 (N_6072,N_4651,N_3545);
nand U6073 (N_6073,N_3795,N_1038);
or U6074 (N_6074,N_958,N_4483);
or U6075 (N_6075,N_4279,N_635);
and U6076 (N_6076,N_4139,N_3227);
or U6077 (N_6077,N_3744,N_1795);
nand U6078 (N_6078,N_1051,N_2405);
nor U6079 (N_6079,N_1834,N_3282);
or U6080 (N_6080,N_4700,N_952);
nor U6081 (N_6081,N_1680,N_4874);
or U6082 (N_6082,N_4623,N_2990);
xor U6083 (N_6083,N_4717,N_1586);
and U6084 (N_6084,N_2072,N_564);
or U6085 (N_6085,N_2640,N_1695);
and U6086 (N_6086,N_4567,N_4962);
and U6087 (N_6087,N_380,N_2675);
and U6088 (N_6088,N_2583,N_420);
xor U6089 (N_6089,N_19,N_4932);
xnor U6090 (N_6090,N_78,N_3635);
nor U6091 (N_6091,N_927,N_3735);
nor U6092 (N_6092,N_4334,N_1510);
nand U6093 (N_6093,N_4209,N_2345);
nand U6094 (N_6094,N_2660,N_3260);
nand U6095 (N_6095,N_1940,N_2589);
nand U6096 (N_6096,N_739,N_31);
and U6097 (N_6097,N_656,N_4308);
nor U6098 (N_6098,N_4267,N_2495);
and U6099 (N_6099,N_2134,N_4920);
nor U6100 (N_6100,N_3379,N_2739);
nand U6101 (N_6101,N_4515,N_3149);
nand U6102 (N_6102,N_3498,N_1131);
and U6103 (N_6103,N_1768,N_3297);
nand U6104 (N_6104,N_2322,N_4366);
or U6105 (N_6105,N_580,N_4811);
or U6106 (N_6106,N_1238,N_2117);
nor U6107 (N_6107,N_164,N_1953);
xnor U6108 (N_6108,N_1374,N_3455);
and U6109 (N_6109,N_1244,N_1293);
nand U6110 (N_6110,N_10,N_1457);
nand U6111 (N_6111,N_2318,N_3850);
xor U6112 (N_6112,N_668,N_3012);
nand U6113 (N_6113,N_1805,N_2453);
and U6114 (N_6114,N_3202,N_2756);
and U6115 (N_6115,N_2831,N_223);
and U6116 (N_6116,N_1381,N_814);
and U6117 (N_6117,N_1441,N_548);
and U6118 (N_6118,N_4750,N_3425);
nor U6119 (N_6119,N_1447,N_1468);
nor U6120 (N_6120,N_4117,N_542);
nor U6121 (N_6121,N_1667,N_3350);
and U6122 (N_6122,N_2306,N_742);
nand U6123 (N_6123,N_1108,N_2575);
nand U6124 (N_6124,N_3620,N_671);
nand U6125 (N_6125,N_4175,N_691);
xor U6126 (N_6126,N_231,N_2499);
and U6127 (N_6127,N_3730,N_4428);
or U6128 (N_6128,N_166,N_728);
nor U6129 (N_6129,N_108,N_4683);
nor U6130 (N_6130,N_4821,N_2401);
xor U6131 (N_6131,N_1055,N_469);
and U6132 (N_6132,N_3570,N_741);
or U6133 (N_6133,N_2957,N_4291);
nand U6134 (N_6134,N_3036,N_3660);
and U6135 (N_6135,N_3326,N_1631);
nor U6136 (N_6136,N_174,N_3917);
nor U6137 (N_6137,N_2947,N_3974);
or U6138 (N_6138,N_329,N_308);
nor U6139 (N_6139,N_3846,N_4327);
nand U6140 (N_6140,N_3992,N_2533);
and U6141 (N_6141,N_3046,N_653);
and U6142 (N_6142,N_32,N_2023);
or U6143 (N_6143,N_2609,N_3162);
and U6144 (N_6144,N_1585,N_1280);
and U6145 (N_6145,N_1988,N_519);
xor U6146 (N_6146,N_3075,N_1936);
or U6147 (N_6147,N_2902,N_1974);
xor U6148 (N_6148,N_4843,N_1760);
nor U6149 (N_6149,N_132,N_1588);
or U6150 (N_6150,N_4852,N_205);
nand U6151 (N_6151,N_3941,N_2872);
nor U6152 (N_6152,N_3943,N_4031);
nand U6153 (N_6153,N_825,N_2941);
nand U6154 (N_6154,N_1324,N_1366);
and U6155 (N_6155,N_1681,N_1658);
xor U6156 (N_6156,N_597,N_1384);
nor U6157 (N_6157,N_3045,N_637);
nand U6158 (N_6158,N_3956,N_1255);
or U6159 (N_6159,N_4648,N_4808);
or U6160 (N_6160,N_2860,N_4845);
and U6161 (N_6161,N_2664,N_4905);
xnor U6162 (N_6162,N_2232,N_1424);
xor U6163 (N_6163,N_413,N_272);
xor U6164 (N_6164,N_3000,N_4780);
nand U6165 (N_6165,N_4009,N_1312);
or U6166 (N_6166,N_70,N_4888);
or U6167 (N_6167,N_1758,N_1919);
nand U6168 (N_6168,N_4353,N_4965);
and U6169 (N_6169,N_4631,N_4455);
xor U6170 (N_6170,N_795,N_1602);
nand U6171 (N_6171,N_4354,N_96);
or U6172 (N_6172,N_1263,N_2316);
or U6173 (N_6173,N_4877,N_4389);
xnor U6174 (N_6174,N_1044,N_3084);
nand U6175 (N_6175,N_1997,N_3381);
nor U6176 (N_6176,N_1032,N_3112);
nor U6177 (N_6177,N_4917,N_606);
xnor U6178 (N_6178,N_2258,N_2355);
and U6179 (N_6179,N_3410,N_1227);
xor U6180 (N_6180,N_1364,N_4582);
xor U6181 (N_6181,N_2590,N_4512);
nor U6182 (N_6182,N_4886,N_3784);
nand U6183 (N_6183,N_3863,N_441);
and U6184 (N_6184,N_403,N_1848);
nor U6185 (N_6185,N_4955,N_1944);
and U6186 (N_6186,N_54,N_1920);
nor U6187 (N_6187,N_3240,N_3175);
or U6188 (N_6188,N_603,N_4974);
or U6189 (N_6189,N_3458,N_2822);
xor U6190 (N_6190,N_1565,N_2809);
nand U6191 (N_6191,N_3332,N_3018);
xor U6192 (N_6192,N_4925,N_2014);
or U6193 (N_6193,N_3177,N_1707);
and U6194 (N_6194,N_816,N_3907);
nor U6195 (N_6195,N_2994,N_3497);
nand U6196 (N_6196,N_1298,N_3006);
nand U6197 (N_6197,N_4065,N_3010);
or U6198 (N_6198,N_726,N_1908);
nor U6199 (N_6199,N_3389,N_2837);
nor U6200 (N_6200,N_1144,N_2407);
nand U6201 (N_6201,N_114,N_1943);
nor U6202 (N_6202,N_2112,N_4156);
nor U6203 (N_6203,N_703,N_3507);
nand U6204 (N_6204,N_4224,N_3307);
nor U6205 (N_6205,N_389,N_4906);
xor U6206 (N_6206,N_4422,N_1615);
or U6207 (N_6207,N_497,N_423);
xor U6208 (N_6208,N_3147,N_1563);
and U6209 (N_6209,N_1999,N_4116);
and U6210 (N_6210,N_2356,N_1704);
xnor U6211 (N_6211,N_122,N_887);
nor U6212 (N_6212,N_3589,N_920);
nor U6213 (N_6213,N_2735,N_725);
nor U6214 (N_6214,N_2643,N_1219);
nor U6215 (N_6215,N_4522,N_356);
or U6216 (N_6216,N_478,N_1977);
nor U6217 (N_6217,N_2820,N_973);
and U6218 (N_6218,N_4641,N_4979);
xor U6219 (N_6219,N_3490,N_1976);
nor U6220 (N_6220,N_2982,N_3109);
nor U6221 (N_6221,N_251,N_486);
and U6222 (N_6222,N_233,N_2782);
xor U6223 (N_6223,N_2544,N_3302);
or U6224 (N_6224,N_3984,N_1183);
or U6225 (N_6225,N_4282,N_4296);
and U6226 (N_6226,N_4441,N_485);
or U6227 (N_6227,N_1400,N_2443);
nand U6228 (N_6228,N_349,N_1959);
nand U6229 (N_6229,N_3043,N_4975);
nand U6230 (N_6230,N_4221,N_2934);
and U6231 (N_6231,N_2969,N_438);
xnor U6232 (N_6232,N_40,N_3834);
or U6233 (N_6233,N_2704,N_467);
or U6234 (N_6234,N_4632,N_3085);
or U6235 (N_6235,N_1807,N_1303);
xnor U6236 (N_6236,N_2183,N_4559);
nor U6237 (N_6237,N_3344,N_220);
or U6238 (N_6238,N_468,N_101);
xnor U6239 (N_6239,N_2496,N_1115);
nand U6240 (N_6240,N_3055,N_3906);
and U6241 (N_6241,N_1114,N_727);
xor U6242 (N_6242,N_263,N_1600);
and U6243 (N_6243,N_4276,N_2195);
or U6244 (N_6244,N_823,N_2108);
xnor U6245 (N_6245,N_2577,N_3096);
nor U6246 (N_6246,N_1624,N_2794);
nor U6247 (N_6247,N_1562,N_2018);
xor U6248 (N_6248,N_3047,N_409);
or U6249 (N_6249,N_1938,N_3525);
nand U6250 (N_6250,N_163,N_3140);
xor U6251 (N_6251,N_2745,N_894);
nor U6252 (N_6252,N_3837,N_4778);
nor U6253 (N_6253,N_4945,N_4404);
xnor U6254 (N_6254,N_353,N_774);
nor U6255 (N_6255,N_4285,N_4757);
xor U6256 (N_6256,N_3754,N_2703);
and U6257 (N_6257,N_2560,N_2024);
nand U6258 (N_6258,N_1989,N_966);
or U6259 (N_6259,N_275,N_1369);
nand U6260 (N_6260,N_1960,N_1169);
or U6261 (N_6261,N_1747,N_3335);
nand U6262 (N_6262,N_1859,N_2297);
nor U6263 (N_6263,N_4614,N_3937);
xor U6264 (N_6264,N_2983,N_859);
nand U6265 (N_6265,N_2765,N_2955);
and U6266 (N_6266,N_4067,N_3485);
nand U6267 (N_6267,N_2331,N_4781);
nor U6268 (N_6268,N_4554,N_2013);
nor U6269 (N_6269,N_4163,N_3373);
and U6270 (N_6270,N_2755,N_2646);
and U6271 (N_6271,N_710,N_4642);
and U6272 (N_6272,N_1957,N_2981);
and U6273 (N_6273,N_1608,N_1129);
or U6274 (N_6274,N_1174,N_905);
xnor U6275 (N_6275,N_3836,N_4051);
xnor U6276 (N_6276,N_1552,N_427);
nand U6277 (N_6277,N_2042,N_3091);
and U6278 (N_6278,N_4433,N_3473);
and U6279 (N_6279,N_2341,N_1564);
or U6280 (N_6280,N_2364,N_2349);
xor U6281 (N_6281,N_3378,N_429);
xnor U6282 (N_6282,N_2451,N_1433);
nand U6283 (N_6283,N_2828,N_4875);
nand U6284 (N_6284,N_213,N_4162);
nand U6285 (N_6285,N_4677,N_777);
xnor U6286 (N_6286,N_3551,N_4130);
or U6287 (N_6287,N_808,N_609);
and U6288 (N_6288,N_2730,N_2930);
or U6289 (N_6289,N_1928,N_3594);
and U6290 (N_6290,N_633,N_4724);
nor U6291 (N_6291,N_16,N_3832);
nand U6292 (N_6292,N_4625,N_219);
or U6293 (N_6293,N_4069,N_880);
nand U6294 (N_6294,N_1593,N_4753);
xnor U6295 (N_6295,N_1611,N_3571);
or U6296 (N_6296,N_321,N_718);
and U6297 (N_6297,N_3657,N_761);
and U6298 (N_6298,N_3131,N_4222);
xnor U6299 (N_6299,N_1766,N_1309);
nand U6300 (N_6300,N_2210,N_322);
nand U6301 (N_6301,N_4731,N_4120);
nor U6302 (N_6302,N_904,N_1720);
nor U6303 (N_6303,N_3605,N_3052);
and U6304 (N_6304,N_2780,N_2791);
nor U6305 (N_6305,N_4880,N_931);
or U6306 (N_6306,N_1419,N_2412);
or U6307 (N_6307,N_3270,N_1211);
or U6308 (N_6308,N_3701,N_3737);
and U6309 (N_6309,N_1186,N_992);
or U6310 (N_6310,N_1803,N_3272);
xor U6311 (N_6311,N_3230,N_238);
and U6312 (N_6312,N_2437,N_82);
nor U6313 (N_6313,N_4871,N_3132);
or U6314 (N_6314,N_2501,N_3647);
nor U6315 (N_6315,N_514,N_2237);
or U6316 (N_6316,N_4747,N_4012);
nor U6317 (N_6317,N_3685,N_4814);
nor U6318 (N_6318,N_4649,N_1587);
nand U6319 (N_6319,N_3872,N_267);
nor U6320 (N_6320,N_3374,N_1947);
nor U6321 (N_6321,N_2280,N_2684);
nor U6322 (N_6322,N_499,N_975);
nand U6323 (N_6323,N_2859,N_1501);
xor U6324 (N_6324,N_2884,N_4938);
nor U6325 (N_6325,N_487,N_4589);
nor U6326 (N_6326,N_2847,N_4939);
xor U6327 (N_6327,N_980,N_1099);
or U6328 (N_6328,N_192,N_3971);
nor U6329 (N_6329,N_3706,N_3352);
and U6330 (N_6330,N_2572,N_4036);
nand U6331 (N_6331,N_2338,N_750);
xor U6332 (N_6332,N_2475,N_4191);
or U6333 (N_6333,N_4524,N_2200);
or U6334 (N_6334,N_2411,N_1459);
xor U6335 (N_6335,N_1769,N_2436);
xor U6336 (N_6336,N_4064,N_379);
xor U6337 (N_6337,N_4359,N_4729);
nand U6338 (N_6338,N_882,N_4301);
nor U6339 (N_6339,N_4993,N_4373);
nand U6340 (N_6340,N_3121,N_34);
or U6341 (N_6341,N_4070,N_2095);
nor U6342 (N_6342,N_244,N_2317);
nand U6343 (N_6343,N_2012,N_3818);
xnor U6344 (N_6344,N_612,N_1666);
nor U6345 (N_6345,N_2184,N_4969);
nor U6346 (N_6346,N_921,N_2585);
or U6347 (N_6347,N_1972,N_3554);
or U6348 (N_6348,N_4523,N_2304);
nor U6349 (N_6349,N_968,N_421);
nor U6350 (N_6350,N_860,N_4138);
xor U6351 (N_6351,N_1153,N_2848);
or U6352 (N_6352,N_3593,N_1985);
or U6353 (N_6353,N_20,N_2906);
nor U6354 (N_6354,N_4597,N_3861);
nand U6355 (N_6355,N_2879,N_1812);
xnor U6356 (N_6356,N_1146,N_1193);
nor U6357 (N_6357,N_2339,N_269);
or U6358 (N_6358,N_212,N_3292);
nand U6359 (N_6359,N_1014,N_3440);
and U6360 (N_6360,N_1251,N_2995);
and U6361 (N_6361,N_4699,N_4370);
and U6362 (N_6362,N_262,N_2862);
or U6363 (N_6363,N_526,N_3996);
and U6364 (N_6364,N_2324,N_1863);
and U6365 (N_6365,N_3081,N_2347);
nor U6366 (N_6366,N_3746,N_2723);
and U6367 (N_6367,N_2452,N_3188);
or U6368 (N_6368,N_2421,N_1764);
or U6369 (N_6369,N_2482,N_1000);
xor U6370 (N_6370,N_738,N_2611);
xnor U6371 (N_6371,N_3483,N_715);
and U6372 (N_6372,N_2127,N_3618);
nor U6373 (N_6373,N_3246,N_737);
and U6374 (N_6374,N_3108,N_4420);
nand U6375 (N_6375,N_4010,N_2792);
nand U6376 (N_6376,N_2323,N_3955);
xor U6377 (N_6377,N_2150,N_2068);
or U6378 (N_6378,N_3349,N_1706);
nand U6379 (N_6379,N_4537,N_3281);
nor U6380 (N_6380,N_2931,N_3254);
nor U6381 (N_6381,N_2003,N_1686);
or U6382 (N_6382,N_3866,N_2404);
and U6383 (N_6383,N_4562,N_3541);
xor U6384 (N_6384,N_2668,N_2060);
xor U6385 (N_6385,N_1872,N_4050);
and U6386 (N_6386,N_2333,N_2773);
xnor U6387 (N_6387,N_3510,N_4746);
nor U6388 (N_6388,N_2889,N_2926);
xor U6389 (N_6389,N_4318,N_3154);
and U6390 (N_6390,N_1200,N_4763);
and U6391 (N_6391,N_1230,N_4829);
xor U6392 (N_6392,N_3923,N_1180);
and U6393 (N_6393,N_3921,N_1697);
xnor U6394 (N_6394,N_296,N_532);
nor U6395 (N_6395,N_3714,N_3393);
nor U6396 (N_6396,N_1052,N_2328);
or U6397 (N_6397,N_3135,N_1490);
and U6398 (N_6398,N_1385,N_1065);
nand U6399 (N_6399,N_4804,N_618);
nand U6400 (N_6400,N_2651,N_1407);
or U6401 (N_6401,N_3193,N_4113);
or U6402 (N_6402,N_4926,N_1304);
xor U6403 (N_6403,N_4456,N_3569);
xnor U6404 (N_6404,N_1678,N_829);
nand U6405 (N_6405,N_1068,N_1522);
nand U6406 (N_6406,N_4022,N_3241);
xnor U6407 (N_6407,N_1568,N_585);
xor U6408 (N_6408,N_1285,N_530);
or U6409 (N_6409,N_306,N_3288);
nor U6410 (N_6410,N_1799,N_3886);
nand U6411 (N_6411,N_1788,N_2230);
and U6412 (N_6412,N_1738,N_118);
and U6413 (N_6413,N_3114,N_4405);
or U6414 (N_6414,N_2084,N_4964);
xnor U6415 (N_6415,N_1643,N_301);
nand U6416 (N_6416,N_796,N_2063);
nand U6417 (N_6417,N_2968,N_2087);
or U6418 (N_6418,N_3709,N_3014);
and U6419 (N_6419,N_2158,N_2747);
or U6420 (N_6420,N_4583,N_2971);
nand U6421 (N_6421,N_2,N_2793);
or U6422 (N_6422,N_4394,N_3251);
nand U6423 (N_6423,N_2678,N_2956);
nor U6424 (N_6424,N_2132,N_3294);
xnor U6425 (N_6425,N_3568,N_383);
xor U6426 (N_6426,N_1,N_3522);
xnor U6427 (N_6427,N_3087,N_1229);
nor U6428 (N_6428,N_2868,N_3990);
nand U6429 (N_6429,N_2904,N_4225);
or U6430 (N_6430,N_4976,N_3212);
or U6431 (N_6431,N_1272,N_411);
nor U6432 (N_6432,N_2173,N_1921);
and U6433 (N_6433,N_4278,N_2742);
or U6434 (N_6434,N_2385,N_2700);
or U6435 (N_6435,N_3223,N_2092);
xor U6436 (N_6436,N_2857,N_2808);
xnor U6437 (N_6437,N_2568,N_3822);
xor U6438 (N_6438,N_491,N_3453);
xnor U6439 (N_6439,N_4432,N_2219);
nand U6440 (N_6440,N_3023,N_4918);
nand U6441 (N_6441,N_4315,N_929);
or U6442 (N_6442,N_1841,N_3982);
nor U6443 (N_6443,N_3661,N_3962);
nand U6444 (N_6444,N_4151,N_2178);
xor U6445 (N_6445,N_4611,N_4275);
or U6446 (N_6446,N_2570,N_3838);
and U6447 (N_6447,N_4846,N_133);
and U6448 (N_6448,N_1140,N_1133);
nor U6449 (N_6449,N_2409,N_2269);
nand U6450 (N_6450,N_3925,N_2897);
or U6451 (N_6451,N_4218,N_4256);
or U6452 (N_6452,N_4060,N_924);
nor U6453 (N_6453,N_1661,N_49);
or U6454 (N_6454,N_4488,N_4141);
and U6455 (N_6455,N_4929,N_3599);
or U6456 (N_6456,N_2672,N_501);
nor U6457 (N_6457,N_2460,N_2567);
and U6458 (N_6458,N_1176,N_2311);
and U6459 (N_6459,N_91,N_4847);
nor U6460 (N_6460,N_1294,N_1260);
and U6461 (N_6461,N_1853,N_558);
xnor U6462 (N_6462,N_1955,N_4340);
or U6463 (N_6463,N_680,N_458);
xnor U6464 (N_6464,N_4384,N_2796);
nand U6465 (N_6465,N_2403,N_4094);
xor U6466 (N_6466,N_3186,N_461);
and U6467 (N_6467,N_3427,N_3452);
nor U6468 (N_6468,N_3772,N_2382);
nand U6469 (N_6469,N_1946,N_1618);
nand U6470 (N_6470,N_4127,N_1527);
nor U6471 (N_6471,N_1671,N_1962);
xor U6472 (N_6472,N_37,N_1147);
nand U6473 (N_6473,N_3094,N_4464);
or U6474 (N_6474,N_2163,N_706);
nand U6475 (N_6475,N_1793,N_2450);
nand U6476 (N_6476,N_4903,N_457);
and U6477 (N_6477,N_2939,N_1688);
nor U6478 (N_6478,N_4392,N_1512);
nand U6479 (N_6479,N_3954,N_995);
nand U6480 (N_6480,N_3415,N_1142);
and U6481 (N_6481,N_1275,N_4412);
xnor U6482 (N_6482,N_3261,N_3372);
xnor U6483 (N_6483,N_1421,N_2537);
xor U6484 (N_6484,N_3983,N_4502);
nor U6485 (N_6485,N_4637,N_422);
nor U6486 (N_6486,N_1206,N_1351);
or U6487 (N_6487,N_2972,N_3634);
xnor U6488 (N_6488,N_4928,N_4661);
xor U6489 (N_6489,N_1987,N_997);
or U6490 (N_6490,N_1012,N_2871);
nand U6491 (N_6491,N_4572,N_1370);
xor U6492 (N_6492,N_4169,N_3627);
nand U6493 (N_6493,N_4645,N_4994);
or U6494 (N_6494,N_3998,N_2580);
and U6495 (N_6495,N_3903,N_1329);
nor U6496 (N_6496,N_1013,N_2208);
or U6497 (N_6497,N_2532,N_3314);
and U6498 (N_6498,N_2714,N_3189);
nand U6499 (N_6499,N_4514,N_2688);
or U6500 (N_6500,N_781,N_2488);
nand U6501 (N_6501,N_309,N_4159);
nand U6502 (N_6502,N_4205,N_4068);
nor U6503 (N_6503,N_1307,N_2085);
and U6504 (N_6504,N_4635,N_1992);
nor U6505 (N_6505,N_4185,N_2702);
nand U6506 (N_6506,N_2507,N_2673);
nor U6507 (N_6507,N_1289,N_3988);
xnor U6508 (N_6508,N_4494,N_385);
nor U6509 (N_6509,N_4259,N_1083);
nor U6510 (N_6510,N_4828,N_3196);
or U6511 (N_6511,N_2991,N_2320);
or U6512 (N_6512,N_2645,N_335);
xor U6513 (N_6513,N_2571,N_4041);
xnor U6514 (N_6514,N_2159,N_1344);
nor U6515 (N_6515,N_534,N_1718);
nand U6516 (N_6516,N_4951,N_4505);
xnor U6517 (N_6517,N_1041,N_4176);
nor U6518 (N_6518,N_2428,N_3336);
nor U6519 (N_6519,N_2371,N_4570);
and U6520 (N_6520,N_2658,N_833);
xor U6521 (N_6521,N_1808,N_1670);
nand U6522 (N_6522,N_2239,N_3203);
nand U6523 (N_6523,N_4076,N_3557);
nor U6524 (N_6524,N_4922,N_4766);
nor U6525 (N_6525,N_2344,N_480);
or U6526 (N_6526,N_3881,N_1439);
xor U6527 (N_6527,N_2711,N_2265);
or U6528 (N_6528,N_4084,N_4848);
xnor U6529 (N_6529,N_3626,N_4071);
nand U6530 (N_6530,N_4998,N_1871);
and U6531 (N_6531,N_723,N_3253);
nor U6532 (N_6532,N_4029,N_479);
or U6533 (N_6533,N_1634,N_3777);
or U6534 (N_6534,N_2090,N_4520);
or U6535 (N_6535,N_1898,N_2927);
nand U6536 (N_6536,N_2698,N_1006);
or U6537 (N_6537,N_4831,N_3573);
or U6538 (N_6538,N_3601,N_827);
nand U6539 (N_6539,N_4085,N_4268);
nand U6540 (N_6540,N_2548,N_2527);
xor U6541 (N_6541,N_1492,N_2029);
nand U6542 (N_6542,N_780,N_2579);
or U6543 (N_6543,N_3690,N_3559);
nor U6544 (N_6544,N_3468,N_2962);
nand U6545 (N_6545,N_2918,N_1753);
nor U6546 (N_6546,N_2965,N_1313);
and U6547 (N_6547,N_1639,N_4682);
and U6548 (N_6548,N_2074,N_3756);
nor U6549 (N_6549,N_3220,N_2800);
nand U6550 (N_6550,N_4991,N_4984);
nand U6551 (N_6551,N_922,N_3538);
and U6552 (N_6552,N_1178,N_555);
and U6553 (N_6553,N_2512,N_3961);
and U6554 (N_6554,N_2542,N_252);
xor U6555 (N_6555,N_148,N_1414);
nand U6556 (N_6556,N_4498,N_2500);
nand U6557 (N_6557,N_4016,N_4458);
or U6558 (N_6558,N_351,N_300);
or U6559 (N_6559,N_2059,N_280);
and U6560 (N_6560,N_4867,N_2462);
nor U6561 (N_6561,N_2924,N_4592);
nand U6562 (N_6562,N_4107,N_951);
and U6563 (N_6563,N_234,N_4137);
xnor U6564 (N_6564,N_4702,N_658);
nand U6565 (N_6565,N_2118,N_1966);
or U6566 (N_6566,N_1779,N_2406);
nand U6567 (N_6567,N_2943,N_3460);
nor U6568 (N_6568,N_2205,N_4942);
and U6569 (N_6569,N_4364,N_3509);
or U6570 (N_6570,N_4203,N_551);
nand U6571 (N_6571,N_3069,N_4760);
nor U6572 (N_6572,N_4894,N_209);
and U6573 (N_6573,N_695,N_3172);
nand U6574 (N_6574,N_4578,N_1578);
or U6575 (N_6575,N_2874,N_4426);
or U6576 (N_6576,N_4179,N_4376);
or U6577 (N_6577,N_1431,N_2511);
xor U6578 (N_6578,N_1391,N_4328);
and U6579 (N_6579,N_1092,N_2817);
nor U6580 (N_6580,N_1316,N_4356);
or U6581 (N_6581,N_2298,N_2842);
nand U6582 (N_6582,N_149,N_614);
nand U6583 (N_6583,N_3598,N_4973);
xnor U6584 (N_6584,N_239,N_4155);
and U6585 (N_6585,N_448,N_3951);
nor U6586 (N_6586,N_4140,N_1513);
nand U6587 (N_6587,N_2898,N_2606);
and U6588 (N_6588,N_4733,N_1396);
or U6589 (N_6589,N_2933,N_1722);
xor U6590 (N_6590,N_553,N_3637);
and U6591 (N_6591,N_4742,N_3652);
and U6592 (N_6592,N_906,N_3494);
xor U6593 (N_6593,N_1780,N_86);
or U6594 (N_6594,N_4668,N_3489);
nand U6595 (N_6595,N_3244,N_1993);
nor U6596 (N_6596,N_1854,N_286);
nand U6597 (N_6597,N_1862,N_1831);
and U6598 (N_6598,N_3428,N_3218);
nor U6599 (N_6599,N_3827,N_4734);
nor U6600 (N_6600,N_1151,N_2564);
or U6601 (N_6601,N_2650,N_2032);
or U6602 (N_6602,N_2681,N_1070);
nor U6603 (N_6603,N_2169,N_610);
nor U6604 (N_6604,N_879,N_646);
xor U6605 (N_6605,N_4335,N_3765);
or U6606 (N_6606,N_4686,N_3258);
or U6607 (N_6607,N_1113,N_1787);
nand U6608 (N_6608,N_2310,N_2093);
and U6609 (N_6609,N_2767,N_3817);
nor U6610 (N_6610,N_3152,N_292);
nand U6611 (N_6611,N_588,N_948);
nor U6612 (N_6612,N_3806,N_3146);
or U6613 (N_6613,N_1646,N_4644);
nor U6614 (N_6614,N_3687,N_4716);
xnor U6615 (N_6615,N_2682,N_3508);
nand U6616 (N_6616,N_4910,N_2097);
and U6617 (N_6617,N_4720,N_2806);
nor U6618 (N_6618,N_1119,N_4719);
xor U6619 (N_6619,N_2094,N_4897);
or U6620 (N_6620,N_2812,N_4560);
xor U6621 (N_6621,N_141,N_4463);
nand U6622 (N_6622,N_2988,N_1906);
nor U6623 (N_6623,N_4836,N_255);
or U6624 (N_6624,N_4454,N_4827);
and U6625 (N_6625,N_2608,N_3328);
nor U6626 (N_6626,N_1377,N_762);
nor U6627 (N_6627,N_3380,N_1339);
or U6628 (N_6628,N_4003,N_2899);
nand U6629 (N_6629,N_694,N_249);
nor U6630 (N_6630,N_2844,N_439);
and U6631 (N_6631,N_3103,N_4337);
nor U6632 (N_6632,N_4008,N_2856);
or U6633 (N_6633,N_928,N_4027);
xnor U6634 (N_6634,N_4758,N_4665);
nor U6635 (N_6635,N_2224,N_3516);
or U6636 (N_6636,N_4015,N_2110);
xnor U6637 (N_6637,N_1870,N_3048);
and U6638 (N_6638,N_2656,N_4680);
nor U6639 (N_6639,N_2935,N_2921);
and U6640 (N_6640,N_1497,N_3786);
nand U6641 (N_6641,N_2573,N_1485);
nor U6642 (N_6642,N_2386,N_2754);
nand U6643 (N_6643,N_1482,N_22);
and U6644 (N_6644,N_4575,N_3469);
xnor U6645 (N_6645,N_1929,N_2228);
and U6646 (N_6646,N_2841,N_2492);
and U6647 (N_6647,N_3099,N_4826);
and U6648 (N_6648,N_3546,N_1299);
nor U6649 (N_6649,N_1744,N_3009);
nand U6650 (N_6650,N_4395,N_2661);
xnor U6651 (N_6651,N_1408,N_2394);
nand U6652 (N_6652,N_2039,N_1420);
and U6653 (N_6653,N_4898,N_3306);
xnor U6654 (N_6654,N_4679,N_4338);
xnor U6655 (N_6655,N_4558,N_3367);
nand U6656 (N_6656,N_73,N_1832);
or U6657 (N_6657,N_4681,N_1942);
nand U6658 (N_6658,N_3808,N_4529);
nor U6659 (N_6659,N_4943,N_1476);
or U6660 (N_6660,N_4387,N_1279);
or U6661 (N_6661,N_4273,N_678);
or U6662 (N_6662,N_3884,N_3908);
or U6663 (N_6663,N_3977,N_434);
or U6664 (N_6664,N_2720,N_4666);
and U6665 (N_6665,N_4543,N_39);
or U6666 (N_6666,N_3163,N_2802);
or U6667 (N_6667,N_4177,N_1897);
or U6668 (N_6668,N_1432,N_1401);
nand U6669 (N_6669,N_2923,N_4782);
and U6670 (N_6670,N_2076,N_2129);
and U6671 (N_6671,N_2137,N_4671);
nand U6672 (N_6672,N_4590,N_2718);
and U6673 (N_6673,N_640,N_348);
xnor U6674 (N_6674,N_1483,N_1724);
xnor U6675 (N_6675,N_3632,N_2845);
or U6676 (N_6676,N_1156,N_1549);
and U6677 (N_6677,N_2936,N_4593);
or U6678 (N_6678,N_4660,N_1358);
or U6679 (N_6679,N_3040,N_3891);
xnor U6680 (N_6680,N_253,N_636);
xnor U6681 (N_6681,N_2034,N_502);
or U6682 (N_6682,N_51,N_1467);
xnor U6683 (N_6683,N_2652,N_2520);
nor U6684 (N_6684,N_1196,N_184);
nor U6685 (N_6685,N_2073,N_1824);
xor U6686 (N_6686,N_2393,N_18);
and U6687 (N_6687,N_2814,N_573);
nand U6688 (N_6688,N_3158,N_4728);
nand U6689 (N_6689,N_2340,N_3505);
xor U6690 (N_6690,N_3787,N_3134);
nand U6691 (N_6691,N_2114,N_3136);
or U6692 (N_6692,N_4199,N_1399);
and U6693 (N_6693,N_391,N_2464);
or U6694 (N_6694,N_3675,N_676);
xnor U6695 (N_6695,N_2062,N_2552);
nand U6696 (N_6696,N_4676,N_4332);
nor U6697 (N_6697,N_1772,N_2031);
and U6698 (N_6698,N_4883,N_2627);
nand U6699 (N_6699,N_1629,N_1665);
nor U6700 (N_6700,N_157,N_2015);
xnor U6701 (N_6701,N_579,N_2619);
or U6702 (N_6702,N_1050,N_1547);
nor U6703 (N_6703,N_3995,N_4033);
nand U6704 (N_6704,N_1714,N_536);
nor U6705 (N_6705,N_3928,N_4889);
xnor U6706 (N_6706,N_1675,N_2170);
nand U6707 (N_6707,N_1676,N_1739);
nand U6708 (N_6708,N_3517,N_206);
and U6709 (N_6709,N_4377,N_4738);
nand U6710 (N_6710,N_2155,N_2071);
nor U6711 (N_6711,N_2139,N_3409);
xor U6712 (N_6712,N_2390,N_4170);
nor U6713 (N_6713,N_699,N_2741);
and U6714 (N_6714,N_4777,N_4876);
xnor U6715 (N_6715,N_2563,N_2485);
xor U6716 (N_6716,N_778,N_299);
or U6717 (N_6717,N_4330,N_507);
and U6718 (N_6718,N_2728,N_1357);
and U6719 (N_6719,N_1669,N_3809);
xor U6720 (N_6720,N_1715,N_75);
xnor U6721 (N_6721,N_2446,N_6);
xor U6722 (N_6722,N_611,N_4024);
nor U6723 (N_6723,N_714,N_3327);
or U6724 (N_6724,N_1290,N_354);
nor U6725 (N_6725,N_248,N_1728);
or U6726 (N_6726,N_2709,N_1112);
or U6727 (N_6727,N_1484,N_3985);
xor U6728 (N_6728,N_3897,N_1932);
or U6729 (N_6729,N_1713,N_2098);
and U6730 (N_6730,N_1429,N_917);
or U6731 (N_6731,N_3725,N_500);
and U6732 (N_6732,N_3604,N_346);
or U6733 (N_6733,N_525,N_2030);
xor U6734 (N_6734,N_1792,N_4361);
and U6735 (N_6735,N_3778,N_4115);
xnor U6736 (N_6736,N_1258,N_4152);
xnor U6737 (N_6737,N_4765,N_1654);
xor U6738 (N_6738,N_4732,N_1826);
nor U6739 (N_6739,N_1717,N_820);
nand U6740 (N_6740,N_4345,N_4792);
xor U6741 (N_6741,N_2885,N_892);
or U6742 (N_6742,N_2916,N_4305);
or U6743 (N_6743,N_2641,N_4896);
nor U6744 (N_6744,N_175,N_2038);
or U6745 (N_6745,N_3658,N_961);
xor U6746 (N_6746,N_3732,N_314);
nand U6747 (N_6747,N_3993,N_4509);
xor U6748 (N_6748,N_4171,N_999);
nand U6749 (N_6749,N_830,N_2798);
nor U6750 (N_6750,N_2046,N_3362);
or U6751 (N_6751,N_153,N_3375);
and U6752 (N_6752,N_2214,N_3779);
nor U6753 (N_6753,N_3904,N_2050);
nor U6754 (N_6754,N_382,N_3197);
xor U6755 (N_6755,N_2531,N_2993);
nand U6756 (N_6756,N_1416,N_2992);
nand U6757 (N_6757,N_4992,N_3113);
or U6758 (N_6758,N_3970,N_628);
nor U6759 (N_6759,N_3217,N_1899);
nor U6760 (N_6760,N_2370,N_2932);
or U6761 (N_6761,N_4878,N_818);
nor U6762 (N_6762,N_673,N_113);
and U6763 (N_6763,N_2778,N_1359);
and U6764 (N_6764,N_4695,N_3065);
and U6765 (N_6765,N_567,N_1427);
or U6766 (N_6766,N_3566,N_1213);
and U6767 (N_6767,N_367,N_2622);
xnor U6768 (N_6768,N_4413,N_1730);
nand U6769 (N_6769,N_3038,N_4675);
xor U6770 (N_6770,N_2351,N_4132);
xor U6771 (N_6771,N_1636,N_3849);
nand U6772 (N_6772,N_4557,N_1168);
nor U6773 (N_6773,N_3564,N_1534);
or U6774 (N_6774,N_789,N_1320);
and U6775 (N_6775,N_2553,N_3050);
nand U6776 (N_6776,N_3233,N_3445);
nor U6777 (N_6777,N_3828,N_528);
nor U6778 (N_6778,N_1085,N_2761);
or U6779 (N_6779,N_2194,N_3975);
nor U6780 (N_6780,N_2426,N_898);
nor U6781 (N_6781,N_2737,N_3269);
or U6782 (N_6782,N_3397,N_3364);
nor U6783 (N_6783,N_1735,N_2088);
nor U6784 (N_6784,N_2799,N_3463);
and U6785 (N_6785,N_1257,N_3890);
xor U6786 (N_6786,N_1701,N_168);
or U6787 (N_6787,N_1981,N_41);
nand U6788 (N_6788,N_2776,N_1519);
or U6789 (N_6789,N_1574,N_4739);
or U6790 (N_6790,N_587,N_1489);
or U6791 (N_6791,N_4147,N_2282);
nor U6792 (N_6792,N_4247,N_36);
nand U6793 (N_6793,N_2974,N_2456);
xnor U6794 (N_6794,N_4465,N_900);
xor U6795 (N_6795,N_2300,N_1314);
xnor U6796 (N_6796,N_4266,N_424);
nand U6797 (N_6797,N_1956,N_4035);
nor U6798 (N_6798,N_1398,N_1318);
xor U6799 (N_6799,N_3885,N_751);
and U6800 (N_6800,N_1984,N_4531);
xnor U6801 (N_6801,N_2289,N_2779);
and U6802 (N_6802,N_4344,N_3590);
nand U6803 (N_6803,N_600,N_3268);
or U6804 (N_6804,N_4691,N_4360);
nor U6805 (N_6805,N_4207,N_1528);
nand U6806 (N_6806,N_3462,N_1233);
nor U6807 (N_6807,N_3249,N_4072);
xor U6808 (N_6808,N_230,N_4534);
xor U6809 (N_6809,N_910,N_2292);
and U6810 (N_6810,N_1040,N_2598);
nor U6811 (N_6811,N_3396,N_959);
and U6812 (N_6812,N_516,N_2048);
xor U6813 (N_6813,N_313,N_65);
and U6814 (N_6814,N_2154,N_2881);
xor U6815 (N_6815,N_1195,N_784);
nand U6816 (N_6816,N_531,N_4961);
nand U6817 (N_6817,N_2543,N_4823);
nor U6818 (N_6818,N_4664,N_2964);
and U6819 (N_6819,N_1033,N_1991);
and U6820 (N_6820,N_375,N_117);
and U6821 (N_6821,N_4246,N_782);
nor U6822 (N_6822,N_1409,N_2427);
or U6823 (N_6823,N_4657,N_1423);
nor U6824 (N_6824,N_1291,N_3237);
xnor U6825 (N_6825,N_130,N_1716);
and U6826 (N_6826,N_2086,N_3609);
xor U6827 (N_6827,N_623,N_123);
nor U6828 (N_6828,N_3755,N_3537);
and U6829 (N_6829,N_2257,N_4290);
nor U6830 (N_6830,N_208,N_3694);
nand U6831 (N_6831,N_2880,N_3228);
nand U6832 (N_6832,N_1652,N_1121);
nor U6833 (N_6833,N_2441,N_4173);
or U6834 (N_6834,N_407,N_987);
nor U6835 (N_6835,N_2648,N_3664);
nor U6836 (N_6836,N_916,N_1166);
xnor U6837 (N_6837,N_2597,N_4369);
and U6838 (N_6838,N_2929,N_4840);
or U6839 (N_6839,N_150,N_1637);
and U6840 (N_6840,N_4223,N_1727);
and U6841 (N_6841,N_2764,N_369);
and U6842 (N_6842,N_953,N_1346);
or U6843 (N_6843,N_4715,N_2066);
nand U6844 (N_6844,N_2153,N_4100);
or U6845 (N_6845,N_4859,N_4467);
nand U6846 (N_6846,N_3271,N_2893);
nor U6847 (N_6847,N_4561,N_4470);
nand U6848 (N_6848,N_2484,N_17);
and U6849 (N_6849,N_2604,N_2166);
xor U6850 (N_6850,N_1954,N_3540);
nand U6851 (N_6851,N_1514,N_3365);
or U6852 (N_6852,N_1434,N_4190);
or U6853 (N_6853,N_1464,N_1711);
or U6854 (N_6854,N_3649,N_3852);
xnor U6855 (N_6855,N_3868,N_4741);
nor U6856 (N_6856,N_2402,N_586);
xor U6857 (N_6857,N_3558,N_3663);
nand U6858 (N_6858,N_629,N_3363);
or U6859 (N_6859,N_2830,N_2104);
nand U6860 (N_6860,N_4532,N_4406);
xnor U6861 (N_6861,N_3697,N_2283);
nor U6862 (N_6862,N_2312,N_993);
nor U6863 (N_6863,N_2019,N_4333);
xnor U6864 (N_6864,N_4075,N_521);
nor U6865 (N_6865,N_87,N_1980);
and U6866 (N_6866,N_3071,N_2361);
and U6867 (N_6867,N_3171,N_4017);
and U6868 (N_6868,N_3689,N_88);
and U6869 (N_6869,N_1625,N_2455);
xor U6870 (N_6870,N_4833,N_4264);
xnor U6871 (N_6871,N_3654,N_3290);
and U6872 (N_6872,N_1442,N_1572);
and U6873 (N_6873,N_3857,N_473);
nor U6874 (N_6874,N_4390,N_2203);
nand U6875 (N_6875,N_1207,N_2615);
xor U6876 (N_6876,N_4485,N_1069);
nor U6877 (N_6877,N_2524,N_4272);
nand U6878 (N_6878,N_2603,N_1436);
nor U6879 (N_6879,N_4118,N_4866);
and U6880 (N_6880,N_4431,N_529);
or U6881 (N_6881,N_4086,N_1331);
and U6882 (N_6882,N_1127,N_3826);
nand U6883 (N_6883,N_2440,N_3444);
xor U6884 (N_6884,N_1458,N_1604);
and U6885 (N_6885,N_3619,N_2989);
or U6886 (N_6886,N_650,N_2612);
or U6887 (N_6887,N_2858,N_803);
nor U6888 (N_6888,N_4398,N_844);
and U6889 (N_6889,N_3608,N_1220);
and U6890 (N_6890,N_4189,N_4703);
or U6891 (N_6891,N_3471,N_4097);
nand U6892 (N_6892,N_3964,N_925);
nand U6893 (N_6893,N_2263,N_4186);
xnor U6894 (N_6894,N_3484,N_3812);
and U6895 (N_6895,N_2535,N_3871);
or U6896 (N_6896,N_4960,N_2581);
and U6897 (N_6897,N_1916,N_4049);
nor U6898 (N_6898,N_639,N_146);
xor U6899 (N_6899,N_2494,N_2281);
nand U6900 (N_6900,N_2033,N_1417);
and U6901 (N_6901,N_1071,N_4453);
xnor U6902 (N_6902,N_3318,N_261);
xor U6903 (N_6903,N_3780,N_2271);
xor U6904 (N_6904,N_1410,N_3844);
and U6905 (N_6905,N_4111,N_3948);
or U6906 (N_6906,N_1101,N_2882);
or U6907 (N_6907,N_4986,N_3377);
nor U6908 (N_6908,N_3395,N_1137);
xnor U6909 (N_6909,N_2069,N_2021);
and U6910 (N_6910,N_245,N_1729);
nor U6911 (N_6911,N_228,N_1511);
or U6912 (N_6912,N_331,N_11);
nor U6913 (N_6913,N_81,N_2733);
and U6914 (N_6914,N_3120,N_3426);
and U6915 (N_6915,N_4692,N_1273);
xnor U6916 (N_6916,N_3215,N_2522);
nor U6917 (N_6917,N_962,N_552);
and U6918 (N_6918,N_4252,N_1225);
or U6919 (N_6919,N_4444,N_3360);
nor U6920 (N_6920,N_3748,N_669);
and U6921 (N_6921,N_4212,N_2854);
nor U6922 (N_6922,N_2307,N_3477);
xnor U6923 (N_6923,N_1105,N_2008);
xnor U6924 (N_6924,N_1171,N_3105);
or U6925 (N_6925,N_2181,N_3042);
nand U6926 (N_6926,N_1653,N_4841);
nor U6927 (N_6927,N_1910,N_4547);
and U6928 (N_6928,N_1837,N_4230);
and U6929 (N_6929,N_1128,N_1066);
and U6930 (N_6930,N_4469,N_665);
or U6931 (N_6931,N_1856,N_1487);
nand U6932 (N_6932,N_3938,N_3548);
nor U6933 (N_6933,N_3488,N_3762);
or U6934 (N_6934,N_4374,N_2706);
nor U6935 (N_6935,N_180,N_861);
or U6936 (N_6936,N_568,N_187);
xor U6937 (N_6937,N_2984,N_471);
nand U6938 (N_6938,N_1892,N_3912);
nand U6939 (N_6939,N_700,N_3310);
or U6940 (N_6940,N_2480,N_772);
or U6941 (N_6941,N_2744,N_3588);
nor U6942 (N_6942,N_1950,N_305);
and U6943 (N_6943,N_707,N_2231);
and U6944 (N_6944,N_3526,N_4480);
and U6945 (N_6945,N_2243,N_828);
nor U6946 (N_6946,N_2623,N_4265);
or U6947 (N_6947,N_3115,N_3309);
and U6948 (N_6948,N_4972,N_4324);
and U6949 (N_6949,N_2201,N_974);
and U6950 (N_6950,N_3713,N_3892);
or U6951 (N_6951,N_2805,N_1389);
xor U6952 (N_6952,N_2360,N_2262);
or U6953 (N_6953,N_1674,N_3361);
and U6954 (N_6954,N_2438,N_3936);
nor U6955 (N_6955,N_4541,N_447);
or U6956 (N_6956,N_4336,N_1839);
nand U6957 (N_6957,N_2669,N_1614);
nand U6958 (N_6958,N_3699,N_3316);
or U6959 (N_6959,N_3692,N_3137);
and U6960 (N_6960,N_3450,N_3472);
nor U6961 (N_6961,N_287,N_342);
xor U6962 (N_6962,N_693,N_4952);
nor U6963 (N_6963,N_4059,N_3300);
nor U6964 (N_6964,N_2713,N_2917);
or U6965 (N_6965,N_4950,N_1380);
and U6966 (N_6966,N_837,N_326);
or U6967 (N_6967,N_4793,N_2161);
nand U6968 (N_6968,N_589,N_2540);
or U6969 (N_6969,N_3914,N_4119);
or U6970 (N_6970,N_4629,N_3825);
and U6971 (N_6971,N_1500,N_2164);
nand U6972 (N_6972,N_3313,N_2483);
and U6973 (N_6973,N_1330,N_1719);
nor U6974 (N_6974,N_504,N_2264);
or U6975 (N_6975,N_152,N_672);
and U6976 (N_6976,N_3285,N_4321);
and U6977 (N_6977,N_2325,N_1061);
nand U6978 (N_6978,N_3235,N_463);
nor U6979 (N_6979,N_3276,N_3127);
nand U6980 (N_6980,N_1080,N_3678);
nor U6981 (N_6981,N_2908,N_605);
and U6982 (N_6982,N_4450,N_359);
nand U6983 (N_6983,N_3693,N_3092);
nor U6984 (N_6984,N_4835,N_926);
and U6985 (N_6985,N_1785,N_4005);
nor U6986 (N_6986,N_2041,N_2758);
and U6987 (N_6987,N_4915,N_4415);
nand U6988 (N_6988,N_4959,N_3882);
nand U6989 (N_6989,N_1592,N_376);
xor U6990 (N_6990,N_3150,N_2384);
nand U6991 (N_6991,N_578,N_1736);
nor U6992 (N_6992,N_2107,N_3089);
nor U6993 (N_6993,N_4650,N_2530);
nand U6994 (N_6994,N_4028,N_107);
xor U6995 (N_6995,N_2125,N_3749);
xor U6996 (N_6996,N_4271,N_2705);
nor U6997 (N_6997,N_273,N_3636);
xnor U6998 (N_6998,N_2036,N_1443);
and U6999 (N_6999,N_1231,N_2593);
nor U7000 (N_7000,N_4517,N_2783);
xnor U7001 (N_7001,N_2329,N_1601);
or U7002 (N_7002,N_4684,N_143);
and U7003 (N_7003,N_2415,N_2883);
nor U7004 (N_7004,N_3873,N_821);
nor U7005 (N_7005,N_1042,N_3421);
xnor U7006 (N_7006,N_1246,N_2156);
nor U7007 (N_7007,N_870,N_4990);
and U7008 (N_7008,N_4214,N_3949);
or U7009 (N_7009,N_363,N_890);
xnor U7010 (N_7010,N_1548,N_4343);
nor U7011 (N_7011,N_226,N_443);
nor U7012 (N_7012,N_688,N_3433);
and U7013 (N_7013,N_2937,N_4443);
and U7014 (N_7014,N_1221,N_232);
xnor U7015 (N_7015,N_373,N_2327);
nand U7016 (N_7016,N_1349,N_196);
nor U7017 (N_7017,N_3932,N_1782);
nand U7018 (N_7018,N_2235,N_4639);
or U7019 (N_7019,N_2309,N_3674);
and U7020 (N_7020,N_2136,N_2116);
nor U7021 (N_7021,N_4685,N_3353);
and U7022 (N_7022,N_1362,N_4824);
and U7023 (N_7023,N_4082,N_720);
and U7024 (N_7024,N_2463,N_2599);
xnor U7025 (N_7025,N_4820,N_3059);
nor U7026 (N_7026,N_3782,N_1154);
or U7027 (N_7027,N_619,N_277);
and U7028 (N_7028,N_4996,N_1173);
and U7029 (N_7029,N_2146,N_4516);
nand U7030 (N_7030,N_836,N_2726);
xnor U7031 (N_7031,N_4262,N_1117);
xnor U7032 (N_7032,N_1135,N_4154);
and U7033 (N_7033,N_93,N_506);
xor U7034 (N_7034,N_4769,N_193);
or U7035 (N_7035,N_4798,N_2189);
nor U7036 (N_7036,N_2852,N_2399);
and U7037 (N_7037,N_4490,N_1696);
nor U7038 (N_7038,N_3295,N_822);
nand U7039 (N_7039,N_1192,N_1026);
nor U7040 (N_7040,N_1045,N_775);
nand U7041 (N_7041,N_2467,N_3621);
xor U7042 (N_7042,N_1345,N_897);
nor U7043 (N_7043,N_4143,N_3370);
and U7044 (N_7044,N_2980,N_3999);
or U7045 (N_7045,N_4987,N_4940);
nor U7046 (N_7046,N_4091,N_3016);
xnor U7047 (N_7047,N_4000,N_4446);
xnor U7048 (N_7048,N_1994,N_437);
or U7049 (N_7049,N_3524,N_1100);
nand U7050 (N_7050,N_2240,N_1086);
nor U7051 (N_7051,N_3236,N_224);
nor U7052 (N_7052,N_3712,N_4079);
and U7053 (N_7053,N_866,N_4245);
and U7054 (N_7054,N_2771,N_2721);
xor U7055 (N_7055,N_622,N_4063);
or U7056 (N_7056,N_1535,N_3369);
and U7057 (N_7057,N_3262,N_1011);
xor U7058 (N_7058,N_2303,N_111);
nand U7059 (N_7059,N_3859,N_1104);
and U7060 (N_7060,N_1335,N_982);
and U7061 (N_7061,N_1473,N_1079);
or U7062 (N_7062,N_1334,N_2246);
nand U7063 (N_7063,N_793,N_2740);
nand U7064 (N_7064,N_4258,N_4274);
and U7065 (N_7065,N_2278,N_4701);
and U7066 (N_7066,N_134,N_3250);
xnor U7067 (N_7067,N_408,N_4102);
nor U7068 (N_7068,N_559,N_3708);
xor U7069 (N_7069,N_3600,N_48);
xnor U7070 (N_7070,N_687,N_802);
xnor U7071 (N_7071,N_4310,N_1679);
xnor U7072 (N_7072,N_3587,N_2953);
nand U7073 (N_7073,N_2491,N_1927);
xor U7074 (N_7074,N_3209,N_2212);
nand U7075 (N_7075,N_696,N_370);
and U7076 (N_7076,N_165,N_2600);
xnor U7077 (N_7077,N_3845,N_3738);
and U7078 (N_7078,N_128,N_3968);
or U7079 (N_7079,N_3939,N_1617);
nor U7080 (N_7080,N_102,N_4605);
xnor U7081 (N_7081,N_1162,N_971);
and U7082 (N_7082,N_2209,N_4039);
nor U7083 (N_7083,N_27,N_419);
nand U7084 (N_7084,N_1877,N_3303);
nor U7085 (N_7085,N_3232,N_4471);
nand U7086 (N_7086,N_2373,N_3633);
or U7087 (N_7087,N_2504,N_930);
or U7088 (N_7088,N_3157,N_3504);
nand U7089 (N_7089,N_4239,N_240);
xnor U7090 (N_7090,N_3946,N_3279);
nand U7091 (N_7091,N_2293,N_2190);
nand U7092 (N_7092,N_4240,N_4909);
and U7093 (N_7093,N_3334,N_4663);
and U7094 (N_7094,N_2888,N_912);
nand U7095 (N_7095,N_4304,N_2865);
and U7096 (N_7096,N_3407,N_2637);
and U7097 (N_7097,N_2731,N_4501);
or U7098 (N_7098,N_1394,N_2753);
nor U7099 (N_7099,N_3325,N_392);
and U7100 (N_7100,N_2448,N_3110);
xnor U7101 (N_7101,N_891,N_246);
nand U7102 (N_7102,N_1234,N_3479);
or U7103 (N_7103,N_3529,N_2667);
nand U7104 (N_7104,N_3201,N_1466);
nor U7105 (N_7105,N_1109,N_3408);
xor U7106 (N_7106,N_1800,N_1560);
and U7107 (N_7107,N_950,N_254);
nand U7108 (N_7108,N_645,N_4459);
nor U7109 (N_7109,N_4714,N_145);
xnor U7110 (N_7110,N_3286,N_4231);
and U7111 (N_7111,N_4057,N_3062);
nand U7112 (N_7112,N_1125,N_3404);
and U7113 (N_7113,N_1134,N_2378);
or U7114 (N_7114,N_3919,N_2279);
xnor U7115 (N_7115,N_4379,N_2657);
and U7116 (N_7116,N_677,N_2474);
and U7117 (N_7117,N_4503,N_4128);
nand U7118 (N_7118,N_1763,N_3883);
nand U7119 (N_7119,N_4819,N_1533);
and U7120 (N_7120,N_1968,N_3815);
or U7121 (N_7121,N_2789,N_4424);
nor U7122 (N_7122,N_2582,N_1952);
xnor U7123 (N_7123,N_4970,N_770);
nor U7124 (N_7124,N_453,N_2255);
xor U7125 (N_7125,N_3283,N_4);
nor U7126 (N_7126,N_4552,N_1028);
nand U7127 (N_7127,N_607,N_520);
nor U7128 (N_7128,N_2635,N_2826);
or U7129 (N_7129,N_3259,N_4603);
and U7130 (N_7130,N_2419,N_517);
xor U7131 (N_7131,N_344,N_2486);
and U7132 (N_7132,N_1726,N_4655);
and U7133 (N_7133,N_4365,N_4606);
and U7134 (N_7134,N_3650,N_2429);
xnor U7135 (N_7135,N_3058,N_2624);
xor U7136 (N_7136,N_2000,N_4548);
nand U7137 (N_7137,N_2199,N_2133);
xor U7138 (N_7138,N_4881,N_4368);
xor U7139 (N_7139,N_2549,N_3024);
and U7140 (N_7140,N_1774,N_4487);
xor U7141 (N_7141,N_449,N_1455);
and U7142 (N_7142,N_4933,N_2557);
xnor U7143 (N_7143,N_1478,N_4595);
nand U7144 (N_7144,N_853,N_23);
nor U7145 (N_7145,N_1262,N_851);
nand U7146 (N_7146,N_4653,N_1797);
or U7147 (N_7147,N_105,N_571);
nor U7148 (N_7148,N_1182,N_1418);
nor U7149 (N_7149,N_3037,N_4194);
nor U7150 (N_7150,N_2285,N_1333);
xor U7151 (N_7151,N_1923,N_154);
and U7152 (N_7152,N_225,N_2976);
nand U7153 (N_7153,N_475,N_1284);
or U7154 (N_7154,N_4400,N_3399);
and U7155 (N_7155,N_1245,N_895);
xor U7156 (N_7156,N_115,N_3354);
or U7157 (N_7157,N_395,N_508);
nand U7158 (N_7158,N_3696,N_566);
or U7159 (N_7159,N_1827,N_377);
xnor U7160 (N_7160,N_2273,N_59);
and U7161 (N_7161,N_4511,N_243);
and U7162 (N_7162,N_4674,N_1742);
nor U7163 (N_7163,N_2875,N_3298);
nor U7164 (N_7164,N_799,N_1828);
and U7165 (N_7165,N_1880,N_1365);
or U7166 (N_7166,N_400,N_2949);
and U7167 (N_7167,N_3194,N_1949);
and U7168 (N_7168,N_3446,N_1190);
xnor U7169 (N_7169,N_270,N_3467);
nand U7170 (N_7170,N_4136,N_4508);
nand U7171 (N_7171,N_3221,N_608);
and U7172 (N_7172,N_3266,N_3622);
and U7173 (N_7173,N_1577,N_3854);
xor U7174 (N_7174,N_1757,N_2528);
nand U7175 (N_7175,N_116,N_2082);
and U7176 (N_7176,N_1395,N_4244);
nand U7177 (N_7177,N_824,N_4228);
nor U7178 (N_7178,N_4269,N_4907);
xnor U7179 (N_7179,N_903,N_4241);
and U7180 (N_7180,N_3106,N_1762);
or U7181 (N_7181,N_2960,N_3607);
and U7182 (N_7182,N_1569,N_4042);
xor U7183 (N_7183,N_2398,N_428);
nand U7184 (N_7184,N_2179,N_4001);
or U7185 (N_7185,N_743,N_4941);
nor U7186 (N_7186,N_1538,N_312);
nor U7187 (N_7187,N_4647,N_1305);
or U7188 (N_7188,N_2750,N_843);
nor U7189 (N_7189,N_2975,N_2377);
nor U7190 (N_7190,N_4168,N_358);
and U7191 (N_7191,N_3750,N_3723);
nor U7192 (N_7192,N_1342,N_4260);
and U7193 (N_7193,N_1649,N_1315);
nand U7194 (N_7194,N_1116,N_4339);
and U7195 (N_7195,N_3700,N_734);
nand U7196 (N_7196,N_4104,N_1644);
xor U7197 (N_7197,N_271,N_2979);
and U7198 (N_7198,N_45,N_1796);
xnor U7199 (N_7199,N_1541,N_1311);
and U7200 (N_7200,N_2296,N_4046);
or U7201 (N_7201,N_3547,N_147);
xor U7202 (N_7202,N_4164,N_2853);
nor U7203 (N_7203,N_278,N_976);
or U7204 (N_7204,N_1912,N_2633);
nand U7205 (N_7205,N_1203,N_2515);
or U7206 (N_7206,N_2149,N_763);
nand U7207 (N_7207,N_3980,N_593);
and U7208 (N_7208,N_446,N_745);
or U7209 (N_7209,N_1379,N_3066);
nor U7210 (N_7210,N_594,N_2047);
nand U7211 (N_7211,N_8,N_1205);
or U7212 (N_7212,N_1157,N_1247);
xnor U7213 (N_7213,N_4250,N_345);
and U7214 (N_7214,N_44,N_936);
xnor U7215 (N_7215,N_3368,N_4899);
or U7216 (N_7216,N_1818,N_3603);
nor U7217 (N_7217,N_3800,N_883);
and U7218 (N_7218,N_211,N_2944);
xor U7219 (N_7219,N_4696,N_4800);
xnor U7220 (N_7220,N_2954,N_865);
nor U7221 (N_7221,N_3987,N_3672);
xnor U7222 (N_7222,N_258,N_972);
xnor U7223 (N_7223,N_4215,N_1778);
and U7224 (N_7224,N_2274,N_3514);
and U7225 (N_7225,N_670,N_3384);
or U7226 (N_7226,N_1584,N_4727);
or U7227 (N_7227,N_4293,N_2078);
or U7228 (N_7228,N_1336,N_1232);
nor U7229 (N_7229,N_3101,N_1958);
or U7230 (N_7230,N_4783,N_1306);
nor U7231 (N_7231,N_2389,N_4535);
nor U7232 (N_7232,N_372,N_2766);
and U7233 (N_7233,N_2363,N_1355);
nand U7234 (N_7234,N_3063,N_675);
nor U7235 (N_7235,N_2458,N_805);
and U7236 (N_7236,N_3242,N_2629);
or U7237 (N_7237,N_523,N_1009);
and U7238 (N_7238,N_709,N_3543);
nor U7239 (N_7239,N_1619,N_3111);
nor U7240 (N_7240,N_1212,N_934);
xor U7241 (N_7241,N_2124,N_692);
and U7242 (N_7242,N_454,N_2592);
nor U7243 (N_7243,N_3585,N_768);
and U7244 (N_7244,N_3182,N_4229);
nor U7245 (N_7245,N_3957,N_1111);
nor U7246 (N_7246,N_3766,N_4710);
or U7247 (N_7247,N_1904,N_854);
and U7248 (N_7248,N_3978,N_2204);
or U7249 (N_7249,N_2514,N_135);
and U7250 (N_7250,N_602,N_260);
and U7251 (N_7251,N_2677,N_1274);
xnor U7252 (N_7252,N_1270,N_4418);
xnor U7253 (N_7253,N_3752,N_1755);
or U7254 (N_7254,N_3638,N_1160);
nor U7255 (N_7255,N_4126,N_3531);
xnor U7256 (N_7256,N_3574,N_754);
or U7257 (N_7257,N_2630,N_4210);
xor U7258 (N_7258,N_888,N_3862);
nand U7259 (N_7259,N_4600,N_393);
xnor U7260 (N_7260,N_3210,N_4708);
and U7261 (N_7261,N_1776,N_4946);
and U7262 (N_7262,N_2367,N_4627);
nor U7263 (N_7263,N_1181,N_2197);
and U7264 (N_7264,N_550,N_3192);
xnor U7265 (N_7265,N_3049,N_1382);
xnor U7266 (N_7266,N_1375,N_2010);
and U7267 (N_7267,N_21,N_4254);
xor U7268 (N_7268,N_1609,N_4802);
and U7269 (N_7269,N_2247,N_2207);
nor U7270 (N_7270,N_3944,N_3741);
xnor U7271 (N_7271,N_4283,N_1802);
xor U7272 (N_7272,N_3022,N_4233);
nand U7273 (N_7273,N_3256,N_4292);
nor U7274 (N_7274,N_2915,N_1878);
and U7275 (N_7275,N_4787,N_1865);
nor U7276 (N_7276,N_515,N_4093);
and U7277 (N_7277,N_3584,N_1765);
nand U7278 (N_7278,N_247,N_681);
nor U7279 (N_7279,N_3793,N_1352);
nand U7280 (N_7280,N_333,N_2749);
and U7281 (N_7281,N_1461,N_3231);
nand U7282 (N_7282,N_4754,N_783);
or U7283 (N_7283,N_1659,N_3002);
or U7284 (N_7284,N_2397,N_3056);
and U7285 (N_7285,N_3130,N_2294);
and U7286 (N_7286,N_4307,N_3715);
xnor U7287 (N_7287,N_1550,N_2162);
and U7288 (N_7288,N_4636,N_4518);
and U7289 (N_7289,N_106,N_1271);
and U7290 (N_7290,N_4236,N_179);
nand U7291 (N_7291,N_1822,N_1393);
nand U7292 (N_7292,N_1218,N_1821);
xor U7293 (N_7293,N_4924,N_2379);
xor U7294 (N_7294,N_4791,N_3572);
nand U7295 (N_7295,N_2759,N_2864);
nand U7296 (N_7296,N_2523,N_456);
nand U7297 (N_7297,N_756,N_2900);
or U7298 (N_7298,N_4160,N_3610);
nand U7299 (N_7299,N_2213,N_634);
nand U7300 (N_7300,N_4556,N_445);
xor U7301 (N_7301,N_3896,N_2313);
nor U7302 (N_7302,N_2245,N_85);
or U7303 (N_7303,N_2160,N_381);
xor U7304 (N_7304,N_1539,N_943);
nor U7305 (N_7305,N_2732,N_80);
xor U7306 (N_7306,N_4323,N_3180);
nor U7307 (N_7307,N_642,N_4873);
nor U7308 (N_7308,N_4774,N_3979);
xnor U7309 (N_7309,N_3054,N_2554);
nand U7310 (N_7310,N_3138,N_1024);
xor U7311 (N_7311,N_1699,N_1430);
xor U7312 (N_7312,N_2266,N_1177);
or U7313 (N_7313,N_4357,N_1750);
xnor U7314 (N_7314,N_3491,N_3015);
nand U7315 (N_7315,N_3495,N_4403);
and U7316 (N_7316,N_3581,N_1031);
nor U7317 (N_7317,N_1594,N_2967);
or U7318 (N_7318,N_996,N_221);
nand U7319 (N_7319,N_592,N_4796);
and U7320 (N_7320,N_1252,N_371);
and U7321 (N_7321,N_1655,N_4764);
nor U7322 (N_7322,N_4121,N_3430);
or U7323 (N_7323,N_577,N_1605);
nand U7324 (N_7324,N_576,N_4257);
nor U7325 (N_7325,N_893,N_1909);
and U7326 (N_7326,N_3386,N_1060);
nand U7327 (N_7327,N_3156,N_4602);
or U7328 (N_7328,N_298,N_2148);
nor U7329 (N_7329,N_4584,N_1007);
and U7330 (N_7330,N_2442,N_562);
and U7331 (N_7331,N_3848,N_3083);
nand U7332 (N_7332,N_2655,N_2506);
or U7333 (N_7333,N_1428,N_540);
nand U7334 (N_7334,N_3824,N_3841);
xnor U7335 (N_7335,N_3839,N_4667);
nand U7336 (N_7336,N_2509,N_863);
xnor U7337 (N_7337,N_1077,N_265);
nand U7338 (N_7338,N_964,N_4555);
nor U7339 (N_7339,N_4707,N_3994);
xor U7340 (N_7340,N_4497,N_3482);
nand U7341 (N_7341,N_2218,N_29);
xor U7342 (N_7342,N_1132,N_2478);
xnor U7343 (N_7343,N_4227,N_3820);
nor U7344 (N_7344,N_4313,N_2383);
nor U7345 (N_7345,N_241,N_3976);
nand U7346 (N_7346,N_509,N_4396);
xor U7347 (N_7347,N_2827,N_4579);
nor U7348 (N_7348,N_4020,N_994);
or U7349 (N_7349,N_4281,N_3153);
nand U7350 (N_7350,N_2659,N_2368);
and U7351 (N_7351,N_190,N_1446);
or U7352 (N_7352,N_1804,N_4103);
or U7353 (N_7353,N_2959,N_3704);
and U7354 (N_7354,N_2343,N_2083);
nor U7355 (N_7355,N_3267,N_2821);
nand U7356 (N_7356,N_3769,N_985);
or U7357 (N_7357,N_1202,N_1043);
or U7358 (N_7358,N_4371,N_1761);
xor U7359 (N_7359,N_4401,N_2027);
nor U7360 (N_7360,N_590,N_2987);
or U7361 (N_7361,N_2683,N_1164);
nand U7362 (N_7362,N_2519,N_3184);
and U7363 (N_7363,N_2005,N_2985);
or U7364 (N_7364,N_1214,N_4634);
xnor U7365 (N_7365,N_3359,N_207);
and U7366 (N_7366,N_1373,N_4807);
or U7367 (N_7367,N_3323,N_2326);
xnor U7368 (N_7368,N_1734,N_3768);
or U7369 (N_7369,N_3098,N_1939);
nor U7370 (N_7370,N_100,N_4399);
xor U7371 (N_7371,N_704,N_4355);
nor U7372 (N_7372,N_2870,N_2539);
nand U7373 (N_7373,N_3126,N_2653);
and U7374 (N_7374,N_2241,N_160);
nor U7375 (N_7375,N_1301,N_3122);
nand U7376 (N_7376,N_4167,N_1081);
or U7377 (N_7377,N_1235,N_94);
or U7378 (N_7378,N_12,N_2051);
nor U7379 (N_7379,N_1191,N_697);
and U7380 (N_7380,N_1276,N_3519);
nor U7381 (N_7381,N_2804,N_856);
xor U7382 (N_7382,N_4284,N_2238);
and U7383 (N_7383,N_3810,N_4786);
nor U7384 (N_7384,N_2551,N_1435);
xnor U7385 (N_7385,N_1934,N_71);
xnor U7386 (N_7386,N_4573,N_1471);
and U7387 (N_7387,N_946,N_1477);
nor U7388 (N_7388,N_3823,N_4101);
and U7389 (N_7389,N_3027,N_4409);
or U7390 (N_7390,N_3104,N_3252);
xor U7391 (N_7391,N_3400,N_613);
nand U7392 (N_7392,N_788,N_2424);
or U7393 (N_7393,N_4825,N_2244);
xnor U7394 (N_7394,N_2369,N_3972);
and U7395 (N_7395,N_3208,N_119);
xnor U7396 (N_7396,N_4954,N_1721);
or U7397 (N_7397,N_3383,N_451);
nand U7398 (N_7398,N_1613,N_4475);
xnor U7399 (N_7399,N_960,N_4785);
nand U7400 (N_7400,N_4622,N_2905);
or U7401 (N_7401,N_2080,N_2408);
or U7402 (N_7402,N_2011,N_2561);
and U7403 (N_7403,N_3487,N_2775);
or U7404 (N_7404,N_1224,N_1825);
nand U7405 (N_7405,N_1254,N_1553);
xnor U7406 (N_7406,N_1491,N_1241);
and U7407 (N_7407,N_1599,N_3102);
xnor U7408 (N_7408,N_279,N_3879);
and U7409 (N_7409,N_4999,N_4978);
nand U7410 (N_7410,N_3947,N_1558);
xnor U7411 (N_7411,N_2206,N_1386);
and U7412 (N_7412,N_3129,N_3876);
nand U7413 (N_7413,N_218,N_4795);
nand U7414 (N_7414,N_4799,N_2287);
or U7415 (N_7415,N_4202,N_2790);
or U7416 (N_7416,N_4601,N_3803);
nand U7417 (N_7417,N_155,N_4762);
nand U7418 (N_7418,N_3667,N_390);
nor U7419 (N_7419,N_940,N_752);
nand U7420 (N_7420,N_3549,N_2157);
nand U7421 (N_7421,N_2877,N_1970);
and U7422 (N_7422,N_2958,N_4957);
and U7423 (N_7423,N_3275,N_53);
and U7424 (N_7424,N_4216,N_4080);
or U7425 (N_7425,N_538,N_186);
or U7426 (N_7426,N_4549,N_1495);
nand U7427 (N_7427,N_4995,N_3486);
xor U7428 (N_7428,N_470,N_4309);
nor U7429 (N_7429,N_3511,N_3617);
or U7430 (N_7430,N_3031,N_685);
nor U7431 (N_7431,N_2950,N_2963);
nor U7432 (N_7432,N_2903,N_1894);
or U7433 (N_7433,N_4598,N_3090);
and U7434 (N_7434,N_1046,N_1873);
xnor U7435 (N_7435,N_1269,N_1508);
nand U7436 (N_7436,N_2233,N_4062);
and U7437 (N_7437,N_648,N_513);
and U7438 (N_7438,N_98,N_4382);
nor U7439 (N_7439,N_3703,N_717);
and U7440 (N_7440,N_3020,N_4803);
nor U7441 (N_7441,N_794,N_2009);
nand U7442 (N_7442,N_2045,N_3731);
nand U7443 (N_7443,N_4011,N_1749);
nand U7444 (N_7444,N_873,N_4725);
or U7445 (N_7445,N_2140,N_4931);
or U7446 (N_7446,N_1507,N_195);
xnor U7447 (N_7447,N_3764,N_1973);
nor U7448 (N_7448,N_4133,N_4865);
or U7449 (N_7449,N_365,N_2211);
or U7450 (N_7450,N_686,N_3185);
xnor U7451 (N_7451,N_2321,N_1540);
nor U7452 (N_7452,N_2907,N_3691);
and U7453 (N_7453,N_297,N_4615);
and U7454 (N_7454,N_899,N_320);
xnor U7455 (N_7455,N_3612,N_1884);
and U7456 (N_7456,N_983,N_3391);
nor U7457 (N_7457,N_3963,N_1741);
nand U7458 (N_7458,N_1888,N_35);
nor U7459 (N_7459,N_3264,N_2043);
and U7460 (N_7460,N_3615,N_848);
nand U7461 (N_7461,N_4983,N_889);
xnor U7462 (N_7462,N_2177,N_3580);
xor U7463 (N_7463,N_543,N_3305);
nand U7464 (N_7464,N_1657,N_3642);
nand U7465 (N_7465,N_505,N_3788);
nand U7466 (N_7466,N_2685,N_399);
and U7467 (N_7467,N_981,N_176);
and U7468 (N_7468,N_4818,N_627);
nand U7469 (N_7469,N_785,N_4092);
xor U7470 (N_7470,N_3263,N_2770);
and U7471 (N_7471,N_2410,N_771);
or U7472 (N_7472,N_3454,N_1523);
xnor U7473 (N_7473,N_2006,N_178);
or U7474 (N_7474,N_3666,N_3500);
and U7475 (N_7475,N_217,N_537);
nand U7476 (N_7476,N_740,N_2696);
nand U7477 (N_7477,N_2007,N_496);
nor U7478 (N_7478,N_1048,N_384);
xnor U7479 (N_7479,N_4048,N_4640);
and U7480 (N_7480,N_4021,N_2286);
nor U7481 (N_7481,N_4618,N_4416);
nor U7482 (N_7482,N_989,N_3406);
nor U7483 (N_7483,N_3417,N_1341);
and U7484 (N_7484,N_4350,N_2839);
and U7485 (N_7485,N_773,N_4857);
and U7486 (N_7486,N_3312,N_139);
nand U7487 (N_7487,N_2803,N_518);
or U7488 (N_7488,N_2270,N_583);
xor U7489 (N_7489,N_918,N_1847);
or U7490 (N_7490,N_1515,N_2142);
nor U7491 (N_7491,N_932,N_3128);
nand U7492 (N_7492,N_2928,N_1037);
xnor U7493 (N_7493,N_3893,N_99);
xnor U7494 (N_7494,N_766,N_2896);
or U7495 (N_7495,N_3348,N_2576);
nand U7496 (N_7496,N_4565,N_3347);
nand U7497 (N_7497,N_3060,N_1996);
xnor U7498 (N_7498,N_967,N_4407);
nor U7499 (N_7499,N_2216,N_3542);
xnor U7500 (N_7500,N_1485,N_4964);
or U7501 (N_7501,N_4556,N_4313);
xor U7502 (N_7502,N_2140,N_1667);
xnor U7503 (N_7503,N_1658,N_437);
and U7504 (N_7504,N_2913,N_4472);
nor U7505 (N_7505,N_3463,N_1225);
and U7506 (N_7506,N_2779,N_4462);
nor U7507 (N_7507,N_1078,N_2650);
nand U7508 (N_7508,N_1371,N_2627);
and U7509 (N_7509,N_4850,N_1923);
nand U7510 (N_7510,N_1979,N_1059);
or U7511 (N_7511,N_394,N_3455);
nand U7512 (N_7512,N_1521,N_2303);
xor U7513 (N_7513,N_2979,N_583);
nor U7514 (N_7514,N_1513,N_2050);
and U7515 (N_7515,N_1388,N_692);
nand U7516 (N_7516,N_3950,N_3967);
nor U7517 (N_7517,N_2848,N_2892);
or U7518 (N_7518,N_1488,N_4770);
nand U7519 (N_7519,N_3113,N_2671);
nor U7520 (N_7520,N_3749,N_2394);
or U7521 (N_7521,N_1558,N_3266);
nand U7522 (N_7522,N_1869,N_4142);
and U7523 (N_7523,N_4714,N_4574);
xor U7524 (N_7524,N_771,N_758);
nor U7525 (N_7525,N_2600,N_4912);
nand U7526 (N_7526,N_1514,N_1548);
or U7527 (N_7527,N_94,N_2357);
or U7528 (N_7528,N_2899,N_2127);
nand U7529 (N_7529,N_1751,N_4883);
nor U7530 (N_7530,N_4143,N_1949);
or U7531 (N_7531,N_1585,N_2004);
nor U7532 (N_7532,N_189,N_1088);
nor U7533 (N_7533,N_1459,N_449);
and U7534 (N_7534,N_3771,N_1815);
and U7535 (N_7535,N_1863,N_2190);
xnor U7536 (N_7536,N_2613,N_3053);
nand U7537 (N_7537,N_4398,N_4222);
nor U7538 (N_7538,N_3680,N_1198);
xor U7539 (N_7539,N_421,N_1807);
nand U7540 (N_7540,N_4029,N_1845);
and U7541 (N_7541,N_1662,N_3894);
nor U7542 (N_7542,N_985,N_526);
nand U7543 (N_7543,N_140,N_3713);
xnor U7544 (N_7544,N_3772,N_1452);
nand U7545 (N_7545,N_99,N_769);
and U7546 (N_7546,N_2071,N_471);
xnor U7547 (N_7547,N_444,N_4688);
or U7548 (N_7548,N_3247,N_1391);
nand U7549 (N_7549,N_2540,N_3198);
and U7550 (N_7550,N_4976,N_2316);
or U7551 (N_7551,N_4044,N_4620);
nand U7552 (N_7552,N_4092,N_255);
and U7553 (N_7553,N_2892,N_4765);
nand U7554 (N_7554,N_3324,N_2083);
nand U7555 (N_7555,N_1547,N_2336);
or U7556 (N_7556,N_1085,N_2501);
nand U7557 (N_7557,N_4168,N_4771);
xor U7558 (N_7558,N_4904,N_1287);
or U7559 (N_7559,N_1183,N_1603);
or U7560 (N_7560,N_3728,N_3017);
nor U7561 (N_7561,N_3245,N_29);
or U7562 (N_7562,N_4961,N_1274);
xnor U7563 (N_7563,N_1746,N_37);
or U7564 (N_7564,N_363,N_3097);
or U7565 (N_7565,N_4948,N_4117);
nand U7566 (N_7566,N_4664,N_3698);
or U7567 (N_7567,N_1530,N_191);
xor U7568 (N_7568,N_1865,N_3738);
or U7569 (N_7569,N_3494,N_158);
and U7570 (N_7570,N_292,N_4676);
and U7571 (N_7571,N_2170,N_3615);
or U7572 (N_7572,N_1456,N_2885);
xnor U7573 (N_7573,N_2682,N_2072);
nor U7574 (N_7574,N_656,N_2282);
nor U7575 (N_7575,N_1459,N_3357);
or U7576 (N_7576,N_648,N_3888);
xnor U7577 (N_7577,N_1594,N_4354);
and U7578 (N_7578,N_1372,N_1741);
and U7579 (N_7579,N_3792,N_417);
nor U7580 (N_7580,N_4412,N_524);
and U7581 (N_7581,N_1631,N_2591);
and U7582 (N_7582,N_3990,N_3185);
xnor U7583 (N_7583,N_3801,N_2996);
nand U7584 (N_7584,N_699,N_4683);
nor U7585 (N_7585,N_3359,N_3499);
or U7586 (N_7586,N_4453,N_3196);
and U7587 (N_7587,N_47,N_4911);
nand U7588 (N_7588,N_227,N_888);
nand U7589 (N_7589,N_2226,N_2036);
and U7590 (N_7590,N_4264,N_3980);
or U7591 (N_7591,N_31,N_4796);
xor U7592 (N_7592,N_1841,N_1264);
or U7593 (N_7593,N_3550,N_794);
nand U7594 (N_7594,N_814,N_1959);
or U7595 (N_7595,N_4788,N_2106);
nand U7596 (N_7596,N_1158,N_3604);
nor U7597 (N_7597,N_760,N_2219);
nand U7598 (N_7598,N_888,N_4342);
nor U7599 (N_7599,N_2586,N_1752);
xnor U7600 (N_7600,N_1963,N_3099);
xnor U7601 (N_7601,N_4146,N_4125);
and U7602 (N_7602,N_4448,N_2108);
xor U7603 (N_7603,N_4931,N_1789);
xor U7604 (N_7604,N_3998,N_545);
or U7605 (N_7605,N_4154,N_3541);
and U7606 (N_7606,N_2262,N_938);
nand U7607 (N_7607,N_4395,N_3149);
nor U7608 (N_7608,N_2665,N_4487);
xor U7609 (N_7609,N_3983,N_1002);
nand U7610 (N_7610,N_2108,N_1542);
nor U7611 (N_7611,N_3201,N_1906);
and U7612 (N_7612,N_2950,N_1495);
nand U7613 (N_7613,N_465,N_3641);
and U7614 (N_7614,N_1075,N_442);
and U7615 (N_7615,N_2987,N_3296);
xor U7616 (N_7616,N_3899,N_3210);
nor U7617 (N_7617,N_4932,N_322);
nor U7618 (N_7618,N_2701,N_167);
nand U7619 (N_7619,N_2878,N_4433);
xor U7620 (N_7620,N_267,N_1030);
nand U7621 (N_7621,N_4983,N_439);
or U7622 (N_7622,N_4034,N_1191);
or U7623 (N_7623,N_3469,N_4137);
xor U7624 (N_7624,N_4767,N_4661);
nor U7625 (N_7625,N_2709,N_338);
xor U7626 (N_7626,N_2013,N_3719);
nor U7627 (N_7627,N_4984,N_4443);
nor U7628 (N_7628,N_4687,N_3919);
and U7629 (N_7629,N_4759,N_4639);
nand U7630 (N_7630,N_2121,N_3969);
and U7631 (N_7631,N_4561,N_591);
nor U7632 (N_7632,N_2332,N_1103);
xnor U7633 (N_7633,N_2994,N_4996);
or U7634 (N_7634,N_2269,N_3982);
nand U7635 (N_7635,N_4670,N_2850);
or U7636 (N_7636,N_3294,N_3186);
and U7637 (N_7637,N_1865,N_1461);
or U7638 (N_7638,N_3415,N_3859);
and U7639 (N_7639,N_4669,N_2755);
xnor U7640 (N_7640,N_839,N_143);
nand U7641 (N_7641,N_2638,N_2087);
or U7642 (N_7642,N_4605,N_671);
nor U7643 (N_7643,N_2226,N_2322);
and U7644 (N_7644,N_506,N_4543);
nor U7645 (N_7645,N_2759,N_4461);
nand U7646 (N_7646,N_3017,N_1513);
or U7647 (N_7647,N_4692,N_3408);
and U7648 (N_7648,N_4510,N_2587);
and U7649 (N_7649,N_1614,N_3519);
or U7650 (N_7650,N_3367,N_4104);
nand U7651 (N_7651,N_3085,N_1850);
xnor U7652 (N_7652,N_863,N_2406);
and U7653 (N_7653,N_269,N_1414);
xnor U7654 (N_7654,N_827,N_1449);
nand U7655 (N_7655,N_4226,N_633);
xor U7656 (N_7656,N_3207,N_1248);
nor U7657 (N_7657,N_3815,N_4788);
xor U7658 (N_7658,N_2703,N_2595);
nand U7659 (N_7659,N_2676,N_1609);
and U7660 (N_7660,N_2358,N_4243);
xnor U7661 (N_7661,N_3278,N_1688);
nand U7662 (N_7662,N_2325,N_1172);
nor U7663 (N_7663,N_242,N_1174);
nor U7664 (N_7664,N_3975,N_4082);
xor U7665 (N_7665,N_2234,N_3157);
or U7666 (N_7666,N_992,N_4738);
and U7667 (N_7667,N_3317,N_1780);
and U7668 (N_7668,N_1434,N_4006);
nor U7669 (N_7669,N_4018,N_4226);
or U7670 (N_7670,N_3412,N_621);
and U7671 (N_7671,N_1764,N_2712);
nand U7672 (N_7672,N_3285,N_3724);
nor U7673 (N_7673,N_2805,N_1473);
xor U7674 (N_7674,N_4062,N_732);
nor U7675 (N_7675,N_634,N_174);
or U7676 (N_7676,N_4173,N_4022);
xnor U7677 (N_7677,N_2761,N_105);
nor U7678 (N_7678,N_730,N_4832);
nand U7679 (N_7679,N_500,N_4109);
xor U7680 (N_7680,N_2711,N_1699);
xnor U7681 (N_7681,N_1556,N_318);
and U7682 (N_7682,N_3614,N_1864);
nor U7683 (N_7683,N_4608,N_3250);
xnor U7684 (N_7684,N_4767,N_482);
xnor U7685 (N_7685,N_3544,N_1992);
and U7686 (N_7686,N_3250,N_3656);
and U7687 (N_7687,N_1265,N_2999);
and U7688 (N_7688,N_3173,N_268);
and U7689 (N_7689,N_4671,N_3840);
or U7690 (N_7690,N_4818,N_4868);
and U7691 (N_7691,N_3956,N_3001);
nor U7692 (N_7692,N_2269,N_188);
nor U7693 (N_7693,N_4639,N_3030);
xnor U7694 (N_7694,N_4106,N_3370);
nor U7695 (N_7695,N_4347,N_1240);
or U7696 (N_7696,N_1610,N_1360);
xor U7697 (N_7697,N_832,N_3596);
xnor U7698 (N_7698,N_4850,N_2623);
and U7699 (N_7699,N_1581,N_2304);
nand U7700 (N_7700,N_561,N_4654);
and U7701 (N_7701,N_749,N_1085);
or U7702 (N_7702,N_828,N_2829);
and U7703 (N_7703,N_2410,N_530);
xnor U7704 (N_7704,N_3355,N_4539);
nor U7705 (N_7705,N_1749,N_455);
nand U7706 (N_7706,N_1463,N_2471);
and U7707 (N_7707,N_4590,N_3715);
xnor U7708 (N_7708,N_3586,N_1639);
xnor U7709 (N_7709,N_4394,N_2412);
nor U7710 (N_7710,N_4672,N_2659);
nor U7711 (N_7711,N_4674,N_105);
and U7712 (N_7712,N_534,N_1269);
and U7713 (N_7713,N_1426,N_738);
nor U7714 (N_7714,N_3957,N_1254);
nor U7715 (N_7715,N_3,N_292);
or U7716 (N_7716,N_1108,N_4995);
and U7717 (N_7717,N_1165,N_2547);
nor U7718 (N_7718,N_4948,N_1919);
xor U7719 (N_7719,N_1780,N_1623);
nand U7720 (N_7720,N_3653,N_570);
and U7721 (N_7721,N_2097,N_346);
xor U7722 (N_7722,N_2092,N_4036);
nand U7723 (N_7723,N_1665,N_4077);
nand U7724 (N_7724,N_3143,N_1401);
xor U7725 (N_7725,N_2204,N_3959);
and U7726 (N_7726,N_1306,N_3699);
and U7727 (N_7727,N_4738,N_4224);
or U7728 (N_7728,N_445,N_912);
xor U7729 (N_7729,N_4176,N_4385);
nand U7730 (N_7730,N_3575,N_3989);
nand U7731 (N_7731,N_4514,N_899);
nand U7732 (N_7732,N_1150,N_2026);
nand U7733 (N_7733,N_71,N_1068);
xor U7734 (N_7734,N_423,N_3355);
nand U7735 (N_7735,N_1844,N_3023);
or U7736 (N_7736,N_560,N_940);
nand U7737 (N_7737,N_122,N_2085);
and U7738 (N_7738,N_2750,N_4176);
nor U7739 (N_7739,N_4496,N_922);
or U7740 (N_7740,N_1810,N_1091);
nor U7741 (N_7741,N_358,N_680);
nand U7742 (N_7742,N_4693,N_4552);
or U7743 (N_7743,N_4465,N_2484);
or U7744 (N_7744,N_2313,N_4835);
nand U7745 (N_7745,N_2924,N_2143);
and U7746 (N_7746,N_1522,N_1217);
and U7747 (N_7747,N_4789,N_4311);
nand U7748 (N_7748,N_2670,N_4175);
nor U7749 (N_7749,N_441,N_4895);
nor U7750 (N_7750,N_1765,N_363);
nor U7751 (N_7751,N_2342,N_4556);
nand U7752 (N_7752,N_1402,N_640);
xnor U7753 (N_7753,N_1634,N_2980);
nor U7754 (N_7754,N_753,N_3903);
xnor U7755 (N_7755,N_233,N_1296);
nor U7756 (N_7756,N_2512,N_4726);
nor U7757 (N_7757,N_4068,N_193);
nor U7758 (N_7758,N_2220,N_1650);
nor U7759 (N_7759,N_2434,N_1786);
and U7760 (N_7760,N_2629,N_4856);
nand U7761 (N_7761,N_3131,N_203);
nor U7762 (N_7762,N_3115,N_4643);
nor U7763 (N_7763,N_4593,N_1181);
nand U7764 (N_7764,N_253,N_4253);
or U7765 (N_7765,N_4861,N_1163);
xor U7766 (N_7766,N_694,N_2618);
and U7767 (N_7767,N_1856,N_4800);
xnor U7768 (N_7768,N_595,N_3377);
and U7769 (N_7769,N_2203,N_4306);
nand U7770 (N_7770,N_3344,N_2185);
nor U7771 (N_7771,N_1387,N_4742);
nor U7772 (N_7772,N_697,N_1972);
xnor U7773 (N_7773,N_2501,N_1445);
nand U7774 (N_7774,N_2125,N_4748);
and U7775 (N_7775,N_2469,N_2180);
nor U7776 (N_7776,N_2735,N_3014);
or U7777 (N_7777,N_3471,N_3920);
or U7778 (N_7778,N_2789,N_2282);
nand U7779 (N_7779,N_3160,N_4643);
and U7780 (N_7780,N_4968,N_4580);
nand U7781 (N_7781,N_8,N_1495);
nand U7782 (N_7782,N_4326,N_1697);
nand U7783 (N_7783,N_3426,N_2414);
nand U7784 (N_7784,N_3527,N_1689);
nand U7785 (N_7785,N_2185,N_491);
or U7786 (N_7786,N_1229,N_1858);
and U7787 (N_7787,N_2738,N_4802);
xor U7788 (N_7788,N_3153,N_387);
nand U7789 (N_7789,N_4946,N_2958);
and U7790 (N_7790,N_708,N_1591);
nand U7791 (N_7791,N_42,N_1940);
xnor U7792 (N_7792,N_4382,N_2558);
and U7793 (N_7793,N_1767,N_3229);
nor U7794 (N_7794,N_4786,N_3355);
nor U7795 (N_7795,N_2395,N_2079);
xnor U7796 (N_7796,N_2217,N_250);
and U7797 (N_7797,N_1471,N_4451);
or U7798 (N_7798,N_545,N_4981);
and U7799 (N_7799,N_784,N_791);
xor U7800 (N_7800,N_2837,N_749);
and U7801 (N_7801,N_1881,N_3847);
xnor U7802 (N_7802,N_1781,N_1929);
nor U7803 (N_7803,N_3796,N_2025);
and U7804 (N_7804,N_4269,N_1674);
and U7805 (N_7805,N_4643,N_569);
nor U7806 (N_7806,N_3492,N_4073);
nor U7807 (N_7807,N_3561,N_214);
or U7808 (N_7808,N_4084,N_925);
nor U7809 (N_7809,N_4329,N_2618);
xnor U7810 (N_7810,N_3727,N_3780);
or U7811 (N_7811,N_3195,N_1815);
nand U7812 (N_7812,N_3235,N_2928);
nand U7813 (N_7813,N_352,N_3514);
and U7814 (N_7814,N_288,N_4617);
nand U7815 (N_7815,N_1540,N_382);
nor U7816 (N_7816,N_1663,N_3371);
and U7817 (N_7817,N_1697,N_286);
and U7818 (N_7818,N_813,N_626);
and U7819 (N_7819,N_514,N_3144);
xor U7820 (N_7820,N_2759,N_4731);
xor U7821 (N_7821,N_3679,N_933);
or U7822 (N_7822,N_787,N_1506);
xor U7823 (N_7823,N_4427,N_3903);
and U7824 (N_7824,N_664,N_342);
nor U7825 (N_7825,N_984,N_4164);
xor U7826 (N_7826,N_2734,N_3947);
or U7827 (N_7827,N_3323,N_1544);
xnor U7828 (N_7828,N_584,N_1467);
xnor U7829 (N_7829,N_2233,N_3985);
and U7830 (N_7830,N_2876,N_1286);
xor U7831 (N_7831,N_40,N_3376);
or U7832 (N_7832,N_4793,N_4879);
nor U7833 (N_7833,N_4047,N_449);
or U7834 (N_7834,N_727,N_3572);
xnor U7835 (N_7835,N_1445,N_4074);
and U7836 (N_7836,N_4452,N_4517);
xnor U7837 (N_7837,N_421,N_1926);
or U7838 (N_7838,N_852,N_2048);
nor U7839 (N_7839,N_1896,N_3636);
or U7840 (N_7840,N_1655,N_1977);
or U7841 (N_7841,N_1786,N_795);
and U7842 (N_7842,N_4094,N_1664);
nor U7843 (N_7843,N_4526,N_2659);
or U7844 (N_7844,N_3624,N_3336);
and U7845 (N_7845,N_4834,N_4343);
or U7846 (N_7846,N_4681,N_2938);
nor U7847 (N_7847,N_2254,N_1260);
and U7848 (N_7848,N_1554,N_4939);
xor U7849 (N_7849,N_1203,N_1724);
xnor U7850 (N_7850,N_138,N_1205);
xor U7851 (N_7851,N_596,N_3581);
xor U7852 (N_7852,N_3573,N_4422);
nand U7853 (N_7853,N_1568,N_2801);
or U7854 (N_7854,N_3988,N_831);
nand U7855 (N_7855,N_3600,N_3703);
xor U7856 (N_7856,N_2477,N_558);
and U7857 (N_7857,N_4430,N_1614);
and U7858 (N_7858,N_672,N_2159);
or U7859 (N_7859,N_3970,N_522);
xor U7860 (N_7860,N_1214,N_48);
and U7861 (N_7861,N_2239,N_2529);
nand U7862 (N_7862,N_4298,N_109);
nand U7863 (N_7863,N_2750,N_4292);
and U7864 (N_7864,N_3372,N_4821);
or U7865 (N_7865,N_2745,N_4081);
or U7866 (N_7866,N_3842,N_3146);
xor U7867 (N_7867,N_947,N_3252);
and U7868 (N_7868,N_4181,N_846);
nor U7869 (N_7869,N_4808,N_1);
xnor U7870 (N_7870,N_465,N_4619);
xnor U7871 (N_7871,N_2774,N_2300);
and U7872 (N_7872,N_2392,N_4331);
or U7873 (N_7873,N_1552,N_4580);
or U7874 (N_7874,N_394,N_1346);
or U7875 (N_7875,N_2171,N_391);
nor U7876 (N_7876,N_903,N_2229);
nand U7877 (N_7877,N_427,N_161);
xnor U7878 (N_7878,N_1146,N_3776);
nor U7879 (N_7879,N_3347,N_2636);
xnor U7880 (N_7880,N_1617,N_940);
xor U7881 (N_7881,N_732,N_253);
xnor U7882 (N_7882,N_2835,N_1671);
nor U7883 (N_7883,N_148,N_2837);
or U7884 (N_7884,N_2960,N_3803);
nand U7885 (N_7885,N_3116,N_81);
nor U7886 (N_7886,N_1091,N_1324);
xor U7887 (N_7887,N_4598,N_3224);
nor U7888 (N_7888,N_920,N_4535);
xor U7889 (N_7889,N_3716,N_1316);
or U7890 (N_7890,N_1324,N_2338);
and U7891 (N_7891,N_4657,N_2849);
nor U7892 (N_7892,N_2290,N_3409);
or U7893 (N_7893,N_1782,N_4330);
nand U7894 (N_7894,N_2263,N_462);
or U7895 (N_7895,N_2307,N_2269);
nand U7896 (N_7896,N_3485,N_846);
nand U7897 (N_7897,N_1399,N_3618);
xor U7898 (N_7898,N_2749,N_164);
nand U7899 (N_7899,N_4034,N_3380);
nand U7900 (N_7900,N_2608,N_3250);
xnor U7901 (N_7901,N_2039,N_592);
nand U7902 (N_7902,N_3642,N_482);
xnor U7903 (N_7903,N_3976,N_1439);
xor U7904 (N_7904,N_263,N_1381);
nor U7905 (N_7905,N_1646,N_4445);
nor U7906 (N_7906,N_1619,N_2359);
nor U7907 (N_7907,N_2473,N_671);
or U7908 (N_7908,N_2337,N_3564);
and U7909 (N_7909,N_2878,N_1403);
xor U7910 (N_7910,N_1889,N_1890);
and U7911 (N_7911,N_1667,N_3820);
or U7912 (N_7912,N_2237,N_370);
xnor U7913 (N_7913,N_2427,N_4477);
xor U7914 (N_7914,N_2814,N_3939);
nor U7915 (N_7915,N_962,N_427);
xnor U7916 (N_7916,N_4980,N_36);
or U7917 (N_7917,N_862,N_3733);
nand U7918 (N_7918,N_2682,N_4745);
or U7919 (N_7919,N_4552,N_2125);
xnor U7920 (N_7920,N_4397,N_2838);
and U7921 (N_7921,N_3005,N_2753);
and U7922 (N_7922,N_634,N_1186);
and U7923 (N_7923,N_793,N_3389);
xor U7924 (N_7924,N_25,N_2281);
and U7925 (N_7925,N_3647,N_2690);
and U7926 (N_7926,N_1982,N_4330);
or U7927 (N_7927,N_135,N_4825);
or U7928 (N_7928,N_4984,N_1370);
nor U7929 (N_7929,N_1961,N_2712);
nor U7930 (N_7930,N_1639,N_2263);
nor U7931 (N_7931,N_2522,N_1342);
nor U7932 (N_7932,N_684,N_1595);
or U7933 (N_7933,N_4243,N_4255);
nand U7934 (N_7934,N_2752,N_3529);
or U7935 (N_7935,N_2104,N_1674);
xnor U7936 (N_7936,N_1268,N_3685);
or U7937 (N_7937,N_1238,N_4843);
and U7938 (N_7938,N_741,N_3011);
nand U7939 (N_7939,N_2675,N_4247);
xnor U7940 (N_7940,N_3756,N_4007);
xnor U7941 (N_7941,N_989,N_359);
xnor U7942 (N_7942,N_439,N_2066);
and U7943 (N_7943,N_2924,N_893);
and U7944 (N_7944,N_1115,N_3610);
or U7945 (N_7945,N_311,N_1862);
and U7946 (N_7946,N_3337,N_2149);
nor U7947 (N_7947,N_3807,N_953);
xnor U7948 (N_7948,N_1938,N_4450);
nor U7949 (N_7949,N_4258,N_3295);
or U7950 (N_7950,N_2204,N_2924);
nor U7951 (N_7951,N_758,N_475);
nor U7952 (N_7952,N_4045,N_2038);
xnor U7953 (N_7953,N_2497,N_2691);
xnor U7954 (N_7954,N_626,N_2468);
and U7955 (N_7955,N_3984,N_491);
and U7956 (N_7956,N_66,N_3298);
and U7957 (N_7957,N_4958,N_1382);
nand U7958 (N_7958,N_3436,N_4243);
nand U7959 (N_7959,N_4067,N_2979);
and U7960 (N_7960,N_4870,N_4264);
nor U7961 (N_7961,N_4273,N_1698);
nor U7962 (N_7962,N_4406,N_3667);
or U7963 (N_7963,N_193,N_3464);
nor U7964 (N_7964,N_448,N_2272);
nand U7965 (N_7965,N_878,N_2475);
and U7966 (N_7966,N_1857,N_2418);
and U7967 (N_7967,N_4419,N_4432);
xnor U7968 (N_7968,N_20,N_2244);
or U7969 (N_7969,N_2688,N_3755);
nand U7970 (N_7970,N_187,N_4516);
nand U7971 (N_7971,N_4918,N_1919);
and U7972 (N_7972,N_428,N_2992);
and U7973 (N_7973,N_1036,N_4219);
nand U7974 (N_7974,N_3543,N_2523);
or U7975 (N_7975,N_2649,N_1792);
and U7976 (N_7976,N_1252,N_3593);
nor U7977 (N_7977,N_759,N_1789);
and U7978 (N_7978,N_1692,N_3002);
nand U7979 (N_7979,N_3994,N_4629);
and U7980 (N_7980,N_2119,N_1226);
nor U7981 (N_7981,N_4448,N_3632);
or U7982 (N_7982,N_4979,N_1735);
or U7983 (N_7983,N_3271,N_1878);
or U7984 (N_7984,N_1757,N_3194);
nor U7985 (N_7985,N_3858,N_1197);
or U7986 (N_7986,N_724,N_3718);
and U7987 (N_7987,N_225,N_1922);
or U7988 (N_7988,N_198,N_443);
or U7989 (N_7989,N_1137,N_1822);
xnor U7990 (N_7990,N_307,N_732);
nor U7991 (N_7991,N_2065,N_4633);
nor U7992 (N_7992,N_1722,N_3113);
nor U7993 (N_7993,N_884,N_1837);
and U7994 (N_7994,N_2751,N_3890);
or U7995 (N_7995,N_4647,N_1877);
xnor U7996 (N_7996,N_266,N_546);
nor U7997 (N_7997,N_3660,N_804);
xnor U7998 (N_7998,N_4474,N_2389);
and U7999 (N_7999,N_8,N_4803);
or U8000 (N_8000,N_1905,N_2141);
nor U8001 (N_8001,N_1043,N_4167);
and U8002 (N_8002,N_1708,N_3016);
nand U8003 (N_8003,N_3317,N_4403);
or U8004 (N_8004,N_4925,N_89);
nand U8005 (N_8005,N_1698,N_3256);
and U8006 (N_8006,N_698,N_4137);
nand U8007 (N_8007,N_4251,N_4300);
nand U8008 (N_8008,N_4535,N_2545);
nor U8009 (N_8009,N_1453,N_4747);
xnor U8010 (N_8010,N_415,N_4055);
nor U8011 (N_8011,N_641,N_1516);
and U8012 (N_8012,N_1168,N_4663);
or U8013 (N_8013,N_2696,N_4983);
nor U8014 (N_8014,N_1848,N_1845);
and U8015 (N_8015,N_902,N_1820);
or U8016 (N_8016,N_1831,N_567);
nor U8017 (N_8017,N_393,N_4702);
nor U8018 (N_8018,N_3257,N_271);
nor U8019 (N_8019,N_4052,N_3601);
nor U8020 (N_8020,N_1786,N_2170);
nor U8021 (N_8021,N_1068,N_2506);
nor U8022 (N_8022,N_4216,N_3147);
or U8023 (N_8023,N_2746,N_1303);
or U8024 (N_8024,N_2925,N_1198);
or U8025 (N_8025,N_1657,N_2594);
or U8026 (N_8026,N_3858,N_2978);
xnor U8027 (N_8027,N_3635,N_4448);
xor U8028 (N_8028,N_198,N_1930);
xnor U8029 (N_8029,N_1461,N_2326);
nand U8030 (N_8030,N_2267,N_2774);
and U8031 (N_8031,N_1738,N_4403);
and U8032 (N_8032,N_156,N_4871);
and U8033 (N_8033,N_4478,N_3679);
and U8034 (N_8034,N_4912,N_3534);
or U8035 (N_8035,N_2925,N_4530);
nor U8036 (N_8036,N_779,N_2970);
nand U8037 (N_8037,N_2566,N_4705);
or U8038 (N_8038,N_2532,N_1704);
nand U8039 (N_8039,N_3828,N_81);
and U8040 (N_8040,N_4585,N_3179);
or U8041 (N_8041,N_2381,N_1123);
nand U8042 (N_8042,N_723,N_1059);
nand U8043 (N_8043,N_4798,N_2822);
nor U8044 (N_8044,N_781,N_202);
nor U8045 (N_8045,N_1270,N_3565);
or U8046 (N_8046,N_3764,N_896);
and U8047 (N_8047,N_3733,N_3495);
or U8048 (N_8048,N_4960,N_3396);
or U8049 (N_8049,N_3196,N_1797);
nand U8050 (N_8050,N_2590,N_90);
nand U8051 (N_8051,N_3477,N_3631);
and U8052 (N_8052,N_1717,N_1246);
nand U8053 (N_8053,N_1972,N_2062);
nand U8054 (N_8054,N_1032,N_202);
and U8055 (N_8055,N_4757,N_4985);
xnor U8056 (N_8056,N_974,N_2366);
nor U8057 (N_8057,N_652,N_940);
nor U8058 (N_8058,N_2578,N_3447);
nor U8059 (N_8059,N_4817,N_1945);
or U8060 (N_8060,N_4990,N_327);
xnor U8061 (N_8061,N_996,N_4262);
nor U8062 (N_8062,N_1448,N_202);
nand U8063 (N_8063,N_3648,N_4035);
and U8064 (N_8064,N_3061,N_2572);
xnor U8065 (N_8065,N_972,N_2398);
xor U8066 (N_8066,N_3464,N_368);
xor U8067 (N_8067,N_3352,N_1010);
or U8068 (N_8068,N_3659,N_2785);
xor U8069 (N_8069,N_981,N_460);
xnor U8070 (N_8070,N_4107,N_4510);
nor U8071 (N_8071,N_3324,N_2723);
or U8072 (N_8072,N_4664,N_963);
nand U8073 (N_8073,N_3854,N_1422);
and U8074 (N_8074,N_3224,N_3584);
and U8075 (N_8075,N_1457,N_3260);
nand U8076 (N_8076,N_249,N_2747);
and U8077 (N_8077,N_3349,N_740);
and U8078 (N_8078,N_162,N_4395);
nand U8079 (N_8079,N_1353,N_2320);
nand U8080 (N_8080,N_701,N_2391);
nand U8081 (N_8081,N_2509,N_2562);
xor U8082 (N_8082,N_3613,N_200);
nand U8083 (N_8083,N_1391,N_1836);
nand U8084 (N_8084,N_5,N_1176);
nand U8085 (N_8085,N_3930,N_853);
and U8086 (N_8086,N_562,N_255);
xor U8087 (N_8087,N_1159,N_2730);
nor U8088 (N_8088,N_4003,N_3708);
and U8089 (N_8089,N_3448,N_2533);
and U8090 (N_8090,N_4482,N_3808);
and U8091 (N_8091,N_4846,N_2059);
xor U8092 (N_8092,N_462,N_2165);
xnor U8093 (N_8093,N_3394,N_3635);
nand U8094 (N_8094,N_3895,N_2048);
xor U8095 (N_8095,N_4361,N_3571);
nand U8096 (N_8096,N_2153,N_590);
xnor U8097 (N_8097,N_2557,N_3246);
xor U8098 (N_8098,N_503,N_3552);
and U8099 (N_8099,N_1210,N_4562);
or U8100 (N_8100,N_3881,N_4342);
nor U8101 (N_8101,N_4633,N_4997);
or U8102 (N_8102,N_1615,N_1055);
and U8103 (N_8103,N_4868,N_2787);
xnor U8104 (N_8104,N_2045,N_4869);
or U8105 (N_8105,N_610,N_3111);
and U8106 (N_8106,N_1215,N_3823);
or U8107 (N_8107,N_557,N_901);
nand U8108 (N_8108,N_2277,N_2983);
or U8109 (N_8109,N_809,N_3177);
and U8110 (N_8110,N_1335,N_2024);
and U8111 (N_8111,N_1718,N_786);
nor U8112 (N_8112,N_1303,N_2282);
and U8113 (N_8113,N_1478,N_2943);
nor U8114 (N_8114,N_1483,N_3563);
xor U8115 (N_8115,N_4011,N_1223);
xor U8116 (N_8116,N_854,N_1489);
xnor U8117 (N_8117,N_4660,N_509);
or U8118 (N_8118,N_3251,N_2692);
xnor U8119 (N_8119,N_4150,N_356);
nand U8120 (N_8120,N_986,N_1696);
or U8121 (N_8121,N_1800,N_3231);
xor U8122 (N_8122,N_2204,N_2947);
and U8123 (N_8123,N_676,N_1462);
nor U8124 (N_8124,N_3290,N_4449);
xor U8125 (N_8125,N_846,N_858);
xnor U8126 (N_8126,N_2042,N_1736);
nor U8127 (N_8127,N_418,N_3449);
nor U8128 (N_8128,N_1984,N_4337);
or U8129 (N_8129,N_2846,N_4630);
xor U8130 (N_8130,N_2388,N_3336);
xnor U8131 (N_8131,N_2329,N_3757);
xor U8132 (N_8132,N_2629,N_1330);
xor U8133 (N_8133,N_2992,N_2094);
nor U8134 (N_8134,N_735,N_4976);
xnor U8135 (N_8135,N_3093,N_2653);
and U8136 (N_8136,N_2268,N_3356);
xor U8137 (N_8137,N_2863,N_3775);
xor U8138 (N_8138,N_2311,N_2895);
or U8139 (N_8139,N_881,N_3241);
or U8140 (N_8140,N_782,N_157);
nor U8141 (N_8141,N_2799,N_2863);
and U8142 (N_8142,N_3357,N_2474);
or U8143 (N_8143,N_4028,N_456);
nor U8144 (N_8144,N_728,N_4365);
and U8145 (N_8145,N_4474,N_607);
xor U8146 (N_8146,N_2342,N_3282);
nor U8147 (N_8147,N_3399,N_2736);
and U8148 (N_8148,N_2898,N_4481);
xor U8149 (N_8149,N_167,N_3879);
nand U8150 (N_8150,N_159,N_3062);
or U8151 (N_8151,N_4391,N_2154);
xor U8152 (N_8152,N_3536,N_2974);
nand U8153 (N_8153,N_1237,N_1302);
xnor U8154 (N_8154,N_3400,N_4460);
xor U8155 (N_8155,N_1866,N_3301);
nor U8156 (N_8156,N_1292,N_3029);
nand U8157 (N_8157,N_4870,N_4782);
or U8158 (N_8158,N_3342,N_4779);
nand U8159 (N_8159,N_2747,N_3397);
xor U8160 (N_8160,N_2195,N_1304);
or U8161 (N_8161,N_4051,N_1008);
and U8162 (N_8162,N_1392,N_1631);
nor U8163 (N_8163,N_1757,N_210);
xnor U8164 (N_8164,N_2892,N_2645);
nand U8165 (N_8165,N_3564,N_2399);
or U8166 (N_8166,N_2175,N_2388);
and U8167 (N_8167,N_894,N_2837);
and U8168 (N_8168,N_763,N_4274);
nand U8169 (N_8169,N_3476,N_1148);
nand U8170 (N_8170,N_3683,N_3331);
nand U8171 (N_8171,N_2691,N_1588);
nand U8172 (N_8172,N_3170,N_3189);
xnor U8173 (N_8173,N_3808,N_1846);
and U8174 (N_8174,N_4065,N_3350);
or U8175 (N_8175,N_4053,N_2072);
nor U8176 (N_8176,N_4076,N_2661);
xnor U8177 (N_8177,N_4146,N_1037);
nand U8178 (N_8178,N_4719,N_3054);
xor U8179 (N_8179,N_4164,N_2817);
or U8180 (N_8180,N_1237,N_4695);
and U8181 (N_8181,N_4699,N_760);
and U8182 (N_8182,N_1331,N_1243);
or U8183 (N_8183,N_4712,N_1992);
nand U8184 (N_8184,N_2973,N_3106);
or U8185 (N_8185,N_1130,N_826);
or U8186 (N_8186,N_1279,N_2027);
nand U8187 (N_8187,N_819,N_4189);
nand U8188 (N_8188,N_4811,N_158);
nand U8189 (N_8189,N_69,N_2105);
and U8190 (N_8190,N_3615,N_2150);
nor U8191 (N_8191,N_4378,N_1831);
or U8192 (N_8192,N_4760,N_3985);
and U8193 (N_8193,N_2800,N_2767);
nor U8194 (N_8194,N_2810,N_1266);
and U8195 (N_8195,N_4283,N_92);
nor U8196 (N_8196,N_3145,N_1247);
nand U8197 (N_8197,N_2523,N_3350);
nor U8198 (N_8198,N_2398,N_4189);
and U8199 (N_8199,N_4593,N_3993);
nand U8200 (N_8200,N_1991,N_4670);
and U8201 (N_8201,N_851,N_996);
or U8202 (N_8202,N_4161,N_1997);
and U8203 (N_8203,N_4799,N_3037);
nor U8204 (N_8204,N_2635,N_2210);
xnor U8205 (N_8205,N_2087,N_3514);
or U8206 (N_8206,N_2361,N_1200);
xor U8207 (N_8207,N_4547,N_430);
xnor U8208 (N_8208,N_2431,N_125);
nor U8209 (N_8209,N_4283,N_4962);
or U8210 (N_8210,N_2918,N_761);
nand U8211 (N_8211,N_826,N_1106);
nor U8212 (N_8212,N_3219,N_1817);
or U8213 (N_8213,N_4282,N_2452);
and U8214 (N_8214,N_553,N_3355);
and U8215 (N_8215,N_3845,N_1548);
or U8216 (N_8216,N_1149,N_4503);
nand U8217 (N_8217,N_4597,N_2009);
nand U8218 (N_8218,N_1413,N_187);
nand U8219 (N_8219,N_1220,N_2894);
and U8220 (N_8220,N_4922,N_1116);
and U8221 (N_8221,N_673,N_3836);
nor U8222 (N_8222,N_3783,N_2388);
xor U8223 (N_8223,N_1334,N_4182);
and U8224 (N_8224,N_4583,N_2729);
xor U8225 (N_8225,N_4160,N_2272);
nor U8226 (N_8226,N_2870,N_1025);
nand U8227 (N_8227,N_3335,N_622);
nor U8228 (N_8228,N_948,N_533);
nor U8229 (N_8229,N_1811,N_2575);
nand U8230 (N_8230,N_4012,N_2186);
nor U8231 (N_8231,N_4381,N_256);
nand U8232 (N_8232,N_3198,N_1749);
xnor U8233 (N_8233,N_3538,N_3364);
or U8234 (N_8234,N_4552,N_3291);
nand U8235 (N_8235,N_1375,N_210);
nor U8236 (N_8236,N_4772,N_1075);
xor U8237 (N_8237,N_3311,N_1691);
or U8238 (N_8238,N_40,N_740);
xor U8239 (N_8239,N_2607,N_3133);
nand U8240 (N_8240,N_1204,N_401);
nand U8241 (N_8241,N_2536,N_1969);
xnor U8242 (N_8242,N_474,N_4630);
and U8243 (N_8243,N_2500,N_4739);
and U8244 (N_8244,N_1256,N_1633);
and U8245 (N_8245,N_354,N_4155);
xnor U8246 (N_8246,N_2000,N_1109);
xor U8247 (N_8247,N_648,N_1943);
and U8248 (N_8248,N_4112,N_4271);
nor U8249 (N_8249,N_1104,N_1800);
and U8250 (N_8250,N_3646,N_3111);
xor U8251 (N_8251,N_4829,N_360);
nand U8252 (N_8252,N_1827,N_4914);
and U8253 (N_8253,N_2046,N_3042);
or U8254 (N_8254,N_3982,N_4725);
nor U8255 (N_8255,N_792,N_3128);
nand U8256 (N_8256,N_3394,N_1173);
nand U8257 (N_8257,N_2034,N_1989);
and U8258 (N_8258,N_511,N_3433);
nand U8259 (N_8259,N_1468,N_4218);
xor U8260 (N_8260,N_4670,N_1071);
nor U8261 (N_8261,N_3590,N_3141);
nand U8262 (N_8262,N_3841,N_4750);
and U8263 (N_8263,N_50,N_685);
xor U8264 (N_8264,N_4724,N_4669);
nand U8265 (N_8265,N_4581,N_78);
xnor U8266 (N_8266,N_1408,N_3133);
nand U8267 (N_8267,N_1804,N_4780);
nand U8268 (N_8268,N_435,N_342);
nand U8269 (N_8269,N_899,N_4909);
nand U8270 (N_8270,N_265,N_1162);
and U8271 (N_8271,N_3383,N_3902);
nor U8272 (N_8272,N_4614,N_3574);
nor U8273 (N_8273,N_1732,N_3635);
or U8274 (N_8274,N_297,N_510);
and U8275 (N_8275,N_1012,N_3762);
and U8276 (N_8276,N_3621,N_2575);
and U8277 (N_8277,N_4072,N_4083);
and U8278 (N_8278,N_3611,N_4463);
or U8279 (N_8279,N_4879,N_3136);
nand U8280 (N_8280,N_3466,N_3056);
nor U8281 (N_8281,N_4848,N_3791);
and U8282 (N_8282,N_4094,N_2148);
or U8283 (N_8283,N_2852,N_1677);
nand U8284 (N_8284,N_1869,N_1094);
nand U8285 (N_8285,N_397,N_3304);
and U8286 (N_8286,N_3281,N_833);
nand U8287 (N_8287,N_3555,N_390);
or U8288 (N_8288,N_707,N_0);
or U8289 (N_8289,N_4264,N_2105);
or U8290 (N_8290,N_4799,N_2770);
xnor U8291 (N_8291,N_4175,N_4939);
xor U8292 (N_8292,N_1050,N_1958);
and U8293 (N_8293,N_638,N_3436);
nand U8294 (N_8294,N_1815,N_1964);
nor U8295 (N_8295,N_208,N_1750);
or U8296 (N_8296,N_1980,N_2324);
xor U8297 (N_8297,N_3011,N_2971);
nand U8298 (N_8298,N_2119,N_4095);
xnor U8299 (N_8299,N_2631,N_1703);
and U8300 (N_8300,N_2118,N_2013);
nand U8301 (N_8301,N_3653,N_4990);
nand U8302 (N_8302,N_906,N_2935);
or U8303 (N_8303,N_4691,N_1348);
nor U8304 (N_8304,N_1287,N_4275);
nand U8305 (N_8305,N_1416,N_4234);
and U8306 (N_8306,N_2899,N_3548);
xnor U8307 (N_8307,N_3376,N_721);
nor U8308 (N_8308,N_2281,N_4817);
or U8309 (N_8309,N_802,N_4858);
and U8310 (N_8310,N_1502,N_2104);
xor U8311 (N_8311,N_1411,N_1441);
and U8312 (N_8312,N_3830,N_3816);
nand U8313 (N_8313,N_2897,N_1534);
xor U8314 (N_8314,N_4427,N_3054);
nand U8315 (N_8315,N_4343,N_973);
and U8316 (N_8316,N_1113,N_796);
and U8317 (N_8317,N_4138,N_678);
or U8318 (N_8318,N_2754,N_1988);
xnor U8319 (N_8319,N_1790,N_282);
nor U8320 (N_8320,N_42,N_4244);
xor U8321 (N_8321,N_4477,N_1208);
nor U8322 (N_8322,N_1804,N_606);
or U8323 (N_8323,N_4266,N_588);
nor U8324 (N_8324,N_3330,N_950);
nor U8325 (N_8325,N_4924,N_1389);
and U8326 (N_8326,N_653,N_4740);
nor U8327 (N_8327,N_4640,N_3454);
nand U8328 (N_8328,N_484,N_1415);
nor U8329 (N_8329,N_929,N_4396);
nor U8330 (N_8330,N_2982,N_4846);
and U8331 (N_8331,N_1208,N_3063);
nand U8332 (N_8332,N_951,N_4037);
nor U8333 (N_8333,N_604,N_4673);
and U8334 (N_8334,N_197,N_2095);
xnor U8335 (N_8335,N_1165,N_4361);
nor U8336 (N_8336,N_747,N_3283);
xnor U8337 (N_8337,N_2339,N_4667);
and U8338 (N_8338,N_964,N_801);
and U8339 (N_8339,N_2824,N_4720);
nor U8340 (N_8340,N_617,N_530);
nor U8341 (N_8341,N_652,N_4141);
and U8342 (N_8342,N_2157,N_4061);
and U8343 (N_8343,N_3429,N_4295);
or U8344 (N_8344,N_2107,N_984);
and U8345 (N_8345,N_2000,N_3015);
nand U8346 (N_8346,N_3335,N_2627);
or U8347 (N_8347,N_2590,N_1271);
nor U8348 (N_8348,N_813,N_945);
nor U8349 (N_8349,N_4080,N_4403);
and U8350 (N_8350,N_2621,N_2483);
xor U8351 (N_8351,N_440,N_2462);
or U8352 (N_8352,N_798,N_4119);
and U8353 (N_8353,N_4526,N_4681);
nand U8354 (N_8354,N_4093,N_3685);
nor U8355 (N_8355,N_3893,N_1938);
xnor U8356 (N_8356,N_4882,N_3730);
nand U8357 (N_8357,N_4823,N_3618);
or U8358 (N_8358,N_3475,N_1233);
and U8359 (N_8359,N_4464,N_1409);
xnor U8360 (N_8360,N_3092,N_604);
or U8361 (N_8361,N_337,N_4083);
and U8362 (N_8362,N_4419,N_280);
and U8363 (N_8363,N_4864,N_2864);
or U8364 (N_8364,N_1246,N_794);
nor U8365 (N_8365,N_61,N_680);
nor U8366 (N_8366,N_2957,N_1785);
nor U8367 (N_8367,N_1479,N_3067);
nand U8368 (N_8368,N_3110,N_1048);
or U8369 (N_8369,N_830,N_4774);
xor U8370 (N_8370,N_324,N_4505);
xnor U8371 (N_8371,N_4839,N_3146);
nor U8372 (N_8372,N_1594,N_3479);
xnor U8373 (N_8373,N_3802,N_3213);
nand U8374 (N_8374,N_3352,N_3247);
or U8375 (N_8375,N_3766,N_1559);
xnor U8376 (N_8376,N_3761,N_791);
xor U8377 (N_8377,N_4131,N_1037);
and U8378 (N_8378,N_3140,N_3970);
nor U8379 (N_8379,N_3149,N_4531);
or U8380 (N_8380,N_2473,N_172);
xnor U8381 (N_8381,N_1452,N_3550);
or U8382 (N_8382,N_4243,N_4839);
xor U8383 (N_8383,N_4018,N_756);
nand U8384 (N_8384,N_1949,N_3801);
xnor U8385 (N_8385,N_1364,N_2411);
or U8386 (N_8386,N_2798,N_3267);
nand U8387 (N_8387,N_3530,N_2960);
and U8388 (N_8388,N_2814,N_1227);
nand U8389 (N_8389,N_4728,N_1059);
nor U8390 (N_8390,N_4012,N_4404);
nand U8391 (N_8391,N_3993,N_4373);
nor U8392 (N_8392,N_3064,N_4728);
or U8393 (N_8393,N_3667,N_4305);
nand U8394 (N_8394,N_4978,N_4104);
nand U8395 (N_8395,N_3896,N_4450);
xor U8396 (N_8396,N_2727,N_2886);
and U8397 (N_8397,N_549,N_4237);
nor U8398 (N_8398,N_1406,N_3545);
nor U8399 (N_8399,N_3105,N_2434);
nor U8400 (N_8400,N_752,N_1759);
nor U8401 (N_8401,N_4465,N_2520);
nor U8402 (N_8402,N_1720,N_783);
xor U8403 (N_8403,N_4857,N_479);
nand U8404 (N_8404,N_1125,N_4221);
nor U8405 (N_8405,N_201,N_715);
nand U8406 (N_8406,N_1489,N_4519);
nand U8407 (N_8407,N_4175,N_3829);
or U8408 (N_8408,N_3071,N_920);
xor U8409 (N_8409,N_1179,N_2372);
or U8410 (N_8410,N_2240,N_2111);
or U8411 (N_8411,N_4513,N_1920);
and U8412 (N_8412,N_3352,N_979);
nor U8413 (N_8413,N_3934,N_1227);
xor U8414 (N_8414,N_3385,N_1204);
and U8415 (N_8415,N_1667,N_2350);
or U8416 (N_8416,N_1446,N_2783);
xor U8417 (N_8417,N_2997,N_2778);
and U8418 (N_8418,N_4149,N_429);
nor U8419 (N_8419,N_401,N_782);
xor U8420 (N_8420,N_4301,N_2782);
xor U8421 (N_8421,N_3105,N_2795);
nor U8422 (N_8422,N_2724,N_4586);
xnor U8423 (N_8423,N_4910,N_160);
xor U8424 (N_8424,N_4882,N_3383);
nor U8425 (N_8425,N_4779,N_2629);
nor U8426 (N_8426,N_2303,N_2942);
xnor U8427 (N_8427,N_4116,N_522);
nor U8428 (N_8428,N_4595,N_4017);
or U8429 (N_8429,N_1241,N_3943);
nand U8430 (N_8430,N_1497,N_3292);
or U8431 (N_8431,N_4406,N_103);
xor U8432 (N_8432,N_3604,N_3350);
and U8433 (N_8433,N_557,N_2155);
nand U8434 (N_8434,N_4749,N_3812);
nor U8435 (N_8435,N_1358,N_449);
nor U8436 (N_8436,N_4852,N_1943);
nor U8437 (N_8437,N_3917,N_1542);
and U8438 (N_8438,N_3629,N_1079);
and U8439 (N_8439,N_3575,N_253);
xor U8440 (N_8440,N_2287,N_396);
or U8441 (N_8441,N_107,N_3492);
or U8442 (N_8442,N_1771,N_21);
nor U8443 (N_8443,N_2347,N_2086);
xnor U8444 (N_8444,N_2324,N_626);
nand U8445 (N_8445,N_1635,N_3961);
and U8446 (N_8446,N_1904,N_879);
and U8447 (N_8447,N_34,N_4873);
nand U8448 (N_8448,N_3370,N_1217);
xnor U8449 (N_8449,N_1446,N_634);
and U8450 (N_8450,N_535,N_3926);
nor U8451 (N_8451,N_2338,N_4430);
and U8452 (N_8452,N_2475,N_2331);
xor U8453 (N_8453,N_4843,N_4807);
nand U8454 (N_8454,N_2940,N_4542);
xor U8455 (N_8455,N_1277,N_1553);
and U8456 (N_8456,N_3255,N_1298);
nor U8457 (N_8457,N_597,N_922);
nor U8458 (N_8458,N_838,N_2455);
nand U8459 (N_8459,N_2631,N_3318);
nor U8460 (N_8460,N_3089,N_1750);
nand U8461 (N_8461,N_2919,N_2343);
nor U8462 (N_8462,N_1161,N_4503);
or U8463 (N_8463,N_3099,N_4244);
nor U8464 (N_8464,N_2855,N_4616);
nand U8465 (N_8465,N_1895,N_4126);
nor U8466 (N_8466,N_2443,N_619);
and U8467 (N_8467,N_1334,N_3013);
nand U8468 (N_8468,N_816,N_718);
nand U8469 (N_8469,N_2693,N_1397);
xnor U8470 (N_8470,N_2514,N_227);
and U8471 (N_8471,N_4913,N_3658);
nor U8472 (N_8472,N_844,N_4026);
xnor U8473 (N_8473,N_2440,N_1251);
xor U8474 (N_8474,N_1082,N_4657);
nand U8475 (N_8475,N_293,N_1055);
nor U8476 (N_8476,N_734,N_2085);
or U8477 (N_8477,N_2468,N_4378);
nand U8478 (N_8478,N_3385,N_4373);
nand U8479 (N_8479,N_1976,N_3759);
or U8480 (N_8480,N_1938,N_840);
nor U8481 (N_8481,N_4169,N_322);
or U8482 (N_8482,N_2079,N_3216);
xor U8483 (N_8483,N_704,N_4305);
or U8484 (N_8484,N_2987,N_1505);
or U8485 (N_8485,N_3381,N_1071);
or U8486 (N_8486,N_705,N_2836);
or U8487 (N_8487,N_4141,N_980);
and U8488 (N_8488,N_2709,N_951);
and U8489 (N_8489,N_4195,N_2500);
nand U8490 (N_8490,N_3776,N_2160);
nand U8491 (N_8491,N_3328,N_2604);
xnor U8492 (N_8492,N_1847,N_2908);
nor U8493 (N_8493,N_42,N_4777);
or U8494 (N_8494,N_4538,N_2973);
nand U8495 (N_8495,N_1551,N_2405);
or U8496 (N_8496,N_463,N_707);
and U8497 (N_8497,N_480,N_4054);
or U8498 (N_8498,N_4721,N_158);
or U8499 (N_8499,N_2884,N_3574);
nor U8500 (N_8500,N_2331,N_2150);
nor U8501 (N_8501,N_3525,N_4453);
xnor U8502 (N_8502,N_3456,N_652);
or U8503 (N_8503,N_4176,N_4331);
xor U8504 (N_8504,N_4042,N_4916);
or U8505 (N_8505,N_3625,N_252);
nand U8506 (N_8506,N_998,N_1945);
xor U8507 (N_8507,N_334,N_3680);
and U8508 (N_8508,N_4400,N_348);
xnor U8509 (N_8509,N_3487,N_2563);
nand U8510 (N_8510,N_2278,N_2571);
nand U8511 (N_8511,N_3331,N_793);
or U8512 (N_8512,N_2104,N_1910);
and U8513 (N_8513,N_95,N_2991);
nand U8514 (N_8514,N_791,N_33);
nor U8515 (N_8515,N_4722,N_2799);
xor U8516 (N_8516,N_4729,N_1278);
xnor U8517 (N_8517,N_1701,N_844);
or U8518 (N_8518,N_829,N_4520);
xor U8519 (N_8519,N_2167,N_912);
nor U8520 (N_8520,N_3179,N_1144);
xnor U8521 (N_8521,N_1660,N_4011);
and U8522 (N_8522,N_42,N_846);
xor U8523 (N_8523,N_438,N_3066);
nor U8524 (N_8524,N_3274,N_3182);
and U8525 (N_8525,N_3774,N_2397);
xnor U8526 (N_8526,N_4299,N_3942);
and U8527 (N_8527,N_4092,N_2452);
xnor U8528 (N_8528,N_2159,N_1396);
xor U8529 (N_8529,N_751,N_2071);
or U8530 (N_8530,N_2518,N_3439);
nor U8531 (N_8531,N_3401,N_3443);
nor U8532 (N_8532,N_3002,N_1468);
and U8533 (N_8533,N_4108,N_2002);
xnor U8534 (N_8534,N_52,N_4079);
nor U8535 (N_8535,N_4166,N_2509);
and U8536 (N_8536,N_3785,N_1829);
nor U8537 (N_8537,N_1792,N_3031);
nor U8538 (N_8538,N_3839,N_3178);
xnor U8539 (N_8539,N_1502,N_3300);
and U8540 (N_8540,N_3939,N_93);
or U8541 (N_8541,N_2804,N_246);
nand U8542 (N_8542,N_2972,N_2268);
nor U8543 (N_8543,N_2875,N_1872);
and U8544 (N_8544,N_1047,N_1193);
xor U8545 (N_8545,N_3890,N_4933);
and U8546 (N_8546,N_996,N_4561);
and U8547 (N_8547,N_988,N_4546);
or U8548 (N_8548,N_2506,N_1584);
nor U8549 (N_8549,N_1565,N_1187);
and U8550 (N_8550,N_1018,N_4799);
nor U8551 (N_8551,N_4174,N_1187);
nand U8552 (N_8552,N_1622,N_4129);
or U8553 (N_8553,N_1937,N_213);
and U8554 (N_8554,N_545,N_1287);
or U8555 (N_8555,N_1612,N_4379);
and U8556 (N_8556,N_171,N_3286);
nor U8557 (N_8557,N_1814,N_2623);
and U8558 (N_8558,N_2187,N_1709);
and U8559 (N_8559,N_2652,N_2513);
or U8560 (N_8560,N_3216,N_1813);
and U8561 (N_8561,N_2531,N_4218);
nand U8562 (N_8562,N_103,N_2997);
nor U8563 (N_8563,N_1741,N_3791);
xor U8564 (N_8564,N_3063,N_318);
or U8565 (N_8565,N_1376,N_3534);
xnor U8566 (N_8566,N_4838,N_3390);
and U8567 (N_8567,N_2548,N_3369);
and U8568 (N_8568,N_4539,N_1138);
or U8569 (N_8569,N_1859,N_742);
or U8570 (N_8570,N_2618,N_4241);
xor U8571 (N_8571,N_1046,N_2137);
or U8572 (N_8572,N_4133,N_1859);
or U8573 (N_8573,N_297,N_4637);
or U8574 (N_8574,N_1748,N_2220);
xor U8575 (N_8575,N_4042,N_1211);
nor U8576 (N_8576,N_1687,N_2044);
nor U8577 (N_8577,N_4382,N_4395);
nor U8578 (N_8578,N_1054,N_1983);
or U8579 (N_8579,N_118,N_673);
xnor U8580 (N_8580,N_391,N_250);
nor U8581 (N_8581,N_1575,N_3162);
and U8582 (N_8582,N_4637,N_3739);
or U8583 (N_8583,N_2506,N_3336);
nor U8584 (N_8584,N_3626,N_4649);
nand U8585 (N_8585,N_3384,N_2400);
or U8586 (N_8586,N_1264,N_2901);
or U8587 (N_8587,N_22,N_1802);
nor U8588 (N_8588,N_108,N_4071);
and U8589 (N_8589,N_63,N_1759);
or U8590 (N_8590,N_4184,N_105);
xor U8591 (N_8591,N_4189,N_791);
nor U8592 (N_8592,N_1406,N_3026);
or U8593 (N_8593,N_193,N_1532);
nor U8594 (N_8594,N_3450,N_4089);
nor U8595 (N_8595,N_415,N_4147);
xnor U8596 (N_8596,N_1725,N_1667);
nor U8597 (N_8597,N_4944,N_4198);
or U8598 (N_8598,N_1199,N_265);
or U8599 (N_8599,N_3340,N_4885);
xor U8600 (N_8600,N_748,N_2294);
nand U8601 (N_8601,N_349,N_1707);
and U8602 (N_8602,N_4009,N_564);
xnor U8603 (N_8603,N_4607,N_1259);
xor U8604 (N_8604,N_738,N_3806);
and U8605 (N_8605,N_4535,N_943);
and U8606 (N_8606,N_3876,N_3912);
nand U8607 (N_8607,N_2646,N_3278);
and U8608 (N_8608,N_2527,N_603);
xor U8609 (N_8609,N_3558,N_1266);
or U8610 (N_8610,N_1419,N_2254);
or U8611 (N_8611,N_3799,N_1060);
or U8612 (N_8612,N_4103,N_3374);
nand U8613 (N_8613,N_205,N_1918);
nor U8614 (N_8614,N_3856,N_4668);
and U8615 (N_8615,N_388,N_4733);
nor U8616 (N_8616,N_4382,N_2703);
nor U8617 (N_8617,N_3495,N_4281);
or U8618 (N_8618,N_1246,N_355);
or U8619 (N_8619,N_3708,N_3017);
nand U8620 (N_8620,N_1852,N_4181);
xnor U8621 (N_8621,N_1470,N_2149);
or U8622 (N_8622,N_2365,N_139);
or U8623 (N_8623,N_359,N_1392);
nand U8624 (N_8624,N_1129,N_4046);
nor U8625 (N_8625,N_4311,N_2249);
xor U8626 (N_8626,N_156,N_3147);
xor U8627 (N_8627,N_1819,N_1);
xor U8628 (N_8628,N_4092,N_3741);
nand U8629 (N_8629,N_1124,N_4756);
and U8630 (N_8630,N_4510,N_4082);
nor U8631 (N_8631,N_3002,N_1709);
nor U8632 (N_8632,N_3263,N_1293);
or U8633 (N_8633,N_2953,N_2022);
nand U8634 (N_8634,N_4094,N_2282);
nand U8635 (N_8635,N_3916,N_4395);
nand U8636 (N_8636,N_4587,N_728);
nand U8637 (N_8637,N_2276,N_4675);
nor U8638 (N_8638,N_226,N_2336);
nand U8639 (N_8639,N_1324,N_4040);
or U8640 (N_8640,N_221,N_3781);
nor U8641 (N_8641,N_3754,N_1217);
nor U8642 (N_8642,N_2938,N_2541);
xor U8643 (N_8643,N_958,N_1843);
nor U8644 (N_8644,N_2836,N_4624);
xnor U8645 (N_8645,N_4413,N_3979);
xor U8646 (N_8646,N_4150,N_886);
xor U8647 (N_8647,N_1343,N_4471);
nor U8648 (N_8648,N_4041,N_1830);
xnor U8649 (N_8649,N_4098,N_324);
and U8650 (N_8650,N_3673,N_45);
or U8651 (N_8651,N_1303,N_3158);
nor U8652 (N_8652,N_34,N_685);
nand U8653 (N_8653,N_1418,N_2631);
xnor U8654 (N_8654,N_3942,N_1028);
nand U8655 (N_8655,N_4902,N_3750);
xor U8656 (N_8656,N_938,N_4864);
xnor U8657 (N_8657,N_3215,N_4076);
nand U8658 (N_8658,N_3782,N_4503);
nor U8659 (N_8659,N_4485,N_3205);
xor U8660 (N_8660,N_1921,N_2320);
nand U8661 (N_8661,N_4996,N_4613);
and U8662 (N_8662,N_2558,N_252);
xnor U8663 (N_8663,N_599,N_517);
or U8664 (N_8664,N_4480,N_2746);
and U8665 (N_8665,N_4073,N_1984);
nor U8666 (N_8666,N_4423,N_3063);
and U8667 (N_8667,N_3093,N_4087);
nand U8668 (N_8668,N_3353,N_657);
nand U8669 (N_8669,N_4465,N_4276);
and U8670 (N_8670,N_3172,N_4507);
xor U8671 (N_8671,N_546,N_2107);
nor U8672 (N_8672,N_2528,N_154);
xnor U8673 (N_8673,N_565,N_3467);
and U8674 (N_8674,N_2788,N_1335);
xor U8675 (N_8675,N_1002,N_29);
nor U8676 (N_8676,N_4543,N_1023);
or U8677 (N_8677,N_2375,N_3955);
or U8678 (N_8678,N_2878,N_2958);
nor U8679 (N_8679,N_233,N_4659);
and U8680 (N_8680,N_4477,N_1600);
nand U8681 (N_8681,N_3245,N_1108);
or U8682 (N_8682,N_4188,N_4665);
nor U8683 (N_8683,N_4525,N_1105);
nor U8684 (N_8684,N_1169,N_2252);
nor U8685 (N_8685,N_3890,N_2517);
nor U8686 (N_8686,N_1221,N_3930);
or U8687 (N_8687,N_4144,N_4246);
and U8688 (N_8688,N_3247,N_4088);
nor U8689 (N_8689,N_2400,N_1176);
nor U8690 (N_8690,N_4965,N_3247);
nand U8691 (N_8691,N_3889,N_1385);
nor U8692 (N_8692,N_1394,N_3051);
xnor U8693 (N_8693,N_600,N_1727);
xnor U8694 (N_8694,N_119,N_3385);
and U8695 (N_8695,N_1867,N_1535);
nand U8696 (N_8696,N_1451,N_4710);
or U8697 (N_8697,N_938,N_4902);
nand U8698 (N_8698,N_4946,N_1896);
and U8699 (N_8699,N_4587,N_3625);
and U8700 (N_8700,N_792,N_4847);
or U8701 (N_8701,N_3605,N_3071);
or U8702 (N_8702,N_80,N_3104);
or U8703 (N_8703,N_2076,N_1903);
xnor U8704 (N_8704,N_1351,N_4507);
xor U8705 (N_8705,N_3018,N_1186);
nor U8706 (N_8706,N_489,N_807);
or U8707 (N_8707,N_3441,N_4889);
or U8708 (N_8708,N_3767,N_3297);
xnor U8709 (N_8709,N_4480,N_3115);
xor U8710 (N_8710,N_2731,N_4533);
xor U8711 (N_8711,N_3749,N_2484);
xor U8712 (N_8712,N_1274,N_200);
nor U8713 (N_8713,N_496,N_4866);
xor U8714 (N_8714,N_4946,N_3617);
or U8715 (N_8715,N_3343,N_2109);
nand U8716 (N_8716,N_1307,N_13);
or U8717 (N_8717,N_2764,N_4158);
nand U8718 (N_8718,N_1023,N_3902);
nor U8719 (N_8719,N_397,N_764);
nand U8720 (N_8720,N_341,N_3775);
or U8721 (N_8721,N_3540,N_4239);
xnor U8722 (N_8722,N_3354,N_484);
and U8723 (N_8723,N_680,N_573);
nand U8724 (N_8724,N_3386,N_4080);
xnor U8725 (N_8725,N_4615,N_513);
xor U8726 (N_8726,N_3915,N_2995);
and U8727 (N_8727,N_2695,N_350);
or U8728 (N_8728,N_159,N_798);
nand U8729 (N_8729,N_4336,N_2589);
nor U8730 (N_8730,N_4685,N_2520);
nand U8731 (N_8731,N_3170,N_4427);
nand U8732 (N_8732,N_1147,N_2726);
nand U8733 (N_8733,N_4576,N_967);
nor U8734 (N_8734,N_3715,N_700);
and U8735 (N_8735,N_3027,N_1807);
xnor U8736 (N_8736,N_537,N_4753);
nor U8737 (N_8737,N_1702,N_4766);
or U8738 (N_8738,N_4129,N_3133);
and U8739 (N_8739,N_2138,N_4063);
xnor U8740 (N_8740,N_1685,N_287);
xor U8741 (N_8741,N_2468,N_1796);
or U8742 (N_8742,N_4042,N_525);
and U8743 (N_8743,N_3120,N_277);
and U8744 (N_8744,N_3623,N_1074);
and U8745 (N_8745,N_2953,N_2568);
nand U8746 (N_8746,N_2682,N_3488);
xnor U8747 (N_8747,N_4398,N_973);
or U8748 (N_8748,N_629,N_1902);
and U8749 (N_8749,N_2710,N_2650);
nor U8750 (N_8750,N_1942,N_4379);
nor U8751 (N_8751,N_569,N_1927);
and U8752 (N_8752,N_1127,N_585);
or U8753 (N_8753,N_1005,N_2153);
or U8754 (N_8754,N_4073,N_2033);
nor U8755 (N_8755,N_4113,N_3699);
nor U8756 (N_8756,N_2811,N_2390);
xnor U8757 (N_8757,N_671,N_3123);
nand U8758 (N_8758,N_1189,N_227);
or U8759 (N_8759,N_4634,N_173);
nand U8760 (N_8760,N_3797,N_3614);
nand U8761 (N_8761,N_4242,N_2563);
xor U8762 (N_8762,N_4286,N_4305);
and U8763 (N_8763,N_3169,N_3559);
nor U8764 (N_8764,N_56,N_1040);
nand U8765 (N_8765,N_1601,N_2901);
and U8766 (N_8766,N_3701,N_884);
or U8767 (N_8767,N_1991,N_1005);
or U8768 (N_8768,N_1746,N_4919);
and U8769 (N_8769,N_210,N_3518);
or U8770 (N_8770,N_4754,N_4044);
and U8771 (N_8771,N_1115,N_2357);
nor U8772 (N_8772,N_413,N_4718);
nand U8773 (N_8773,N_2288,N_2342);
and U8774 (N_8774,N_1281,N_2482);
nand U8775 (N_8775,N_3733,N_4896);
xnor U8776 (N_8776,N_4258,N_666);
xnor U8777 (N_8777,N_1370,N_4335);
xnor U8778 (N_8778,N_3410,N_4402);
or U8779 (N_8779,N_3092,N_4340);
or U8780 (N_8780,N_2234,N_4480);
or U8781 (N_8781,N_3809,N_2155);
nor U8782 (N_8782,N_3037,N_2448);
xor U8783 (N_8783,N_4996,N_4541);
nor U8784 (N_8784,N_1723,N_1324);
xor U8785 (N_8785,N_2745,N_4162);
xor U8786 (N_8786,N_1376,N_2272);
xor U8787 (N_8787,N_1363,N_3341);
xnor U8788 (N_8788,N_4642,N_319);
nand U8789 (N_8789,N_2659,N_2586);
xor U8790 (N_8790,N_464,N_4782);
xnor U8791 (N_8791,N_270,N_2495);
nor U8792 (N_8792,N_237,N_2282);
nor U8793 (N_8793,N_4406,N_2060);
nand U8794 (N_8794,N_247,N_531);
nor U8795 (N_8795,N_1315,N_885);
and U8796 (N_8796,N_1870,N_4654);
xor U8797 (N_8797,N_4339,N_518);
nand U8798 (N_8798,N_2046,N_4464);
nand U8799 (N_8799,N_3873,N_4224);
nand U8800 (N_8800,N_911,N_1512);
nor U8801 (N_8801,N_3116,N_1124);
xnor U8802 (N_8802,N_2181,N_1403);
and U8803 (N_8803,N_4026,N_1732);
nor U8804 (N_8804,N_4539,N_1719);
xnor U8805 (N_8805,N_4216,N_894);
and U8806 (N_8806,N_4946,N_658);
xnor U8807 (N_8807,N_903,N_3333);
and U8808 (N_8808,N_1716,N_3711);
or U8809 (N_8809,N_4799,N_89);
nand U8810 (N_8810,N_3352,N_4);
nor U8811 (N_8811,N_1664,N_163);
nor U8812 (N_8812,N_3393,N_2611);
nor U8813 (N_8813,N_1114,N_59);
or U8814 (N_8814,N_127,N_3922);
nand U8815 (N_8815,N_3515,N_2981);
nor U8816 (N_8816,N_67,N_1512);
xnor U8817 (N_8817,N_2915,N_540);
nor U8818 (N_8818,N_1367,N_3408);
and U8819 (N_8819,N_4767,N_2283);
nor U8820 (N_8820,N_368,N_556);
xor U8821 (N_8821,N_1372,N_2301);
xor U8822 (N_8822,N_4423,N_1988);
or U8823 (N_8823,N_2852,N_3912);
and U8824 (N_8824,N_4974,N_264);
or U8825 (N_8825,N_1570,N_2424);
nand U8826 (N_8826,N_786,N_4401);
or U8827 (N_8827,N_697,N_4191);
nor U8828 (N_8828,N_753,N_2394);
nand U8829 (N_8829,N_2603,N_3091);
nor U8830 (N_8830,N_3494,N_2467);
nor U8831 (N_8831,N_1175,N_1018);
nand U8832 (N_8832,N_3367,N_3401);
or U8833 (N_8833,N_1993,N_4112);
nand U8834 (N_8834,N_2075,N_4301);
nor U8835 (N_8835,N_1613,N_64);
xor U8836 (N_8836,N_2061,N_935);
or U8837 (N_8837,N_3922,N_3735);
xnor U8838 (N_8838,N_1608,N_1038);
nand U8839 (N_8839,N_1398,N_4779);
or U8840 (N_8840,N_4856,N_1679);
and U8841 (N_8841,N_1120,N_2631);
nor U8842 (N_8842,N_783,N_3065);
xnor U8843 (N_8843,N_2267,N_1947);
or U8844 (N_8844,N_872,N_2370);
nand U8845 (N_8845,N_2830,N_2987);
or U8846 (N_8846,N_406,N_1799);
nor U8847 (N_8847,N_2021,N_4614);
xor U8848 (N_8848,N_2643,N_1363);
xnor U8849 (N_8849,N_1168,N_1682);
and U8850 (N_8850,N_1503,N_4495);
xor U8851 (N_8851,N_3016,N_4371);
nand U8852 (N_8852,N_3162,N_4938);
nor U8853 (N_8853,N_2905,N_4697);
nand U8854 (N_8854,N_2043,N_3397);
nor U8855 (N_8855,N_3093,N_7);
xor U8856 (N_8856,N_2435,N_4902);
nand U8857 (N_8857,N_23,N_2435);
nand U8858 (N_8858,N_670,N_263);
and U8859 (N_8859,N_2878,N_246);
or U8860 (N_8860,N_1639,N_4647);
nor U8861 (N_8861,N_2043,N_283);
and U8862 (N_8862,N_3507,N_1444);
and U8863 (N_8863,N_955,N_2568);
nand U8864 (N_8864,N_155,N_3735);
xnor U8865 (N_8865,N_3031,N_4414);
xnor U8866 (N_8866,N_1,N_2904);
nor U8867 (N_8867,N_1296,N_87);
and U8868 (N_8868,N_3373,N_3319);
nor U8869 (N_8869,N_4263,N_4237);
or U8870 (N_8870,N_1730,N_2354);
xnor U8871 (N_8871,N_56,N_1269);
and U8872 (N_8872,N_4253,N_2201);
xor U8873 (N_8873,N_3211,N_3470);
nor U8874 (N_8874,N_3741,N_2418);
and U8875 (N_8875,N_1556,N_2542);
or U8876 (N_8876,N_1507,N_1106);
nand U8877 (N_8877,N_801,N_1275);
and U8878 (N_8878,N_3862,N_36);
nand U8879 (N_8879,N_3178,N_618);
nand U8880 (N_8880,N_839,N_3436);
and U8881 (N_8881,N_75,N_3122);
nand U8882 (N_8882,N_1256,N_977);
and U8883 (N_8883,N_1573,N_7);
nor U8884 (N_8884,N_2440,N_3354);
and U8885 (N_8885,N_1477,N_1355);
nand U8886 (N_8886,N_1430,N_3991);
nand U8887 (N_8887,N_4521,N_972);
xor U8888 (N_8888,N_3810,N_4354);
nor U8889 (N_8889,N_4442,N_680);
and U8890 (N_8890,N_678,N_258);
nor U8891 (N_8891,N_1397,N_4785);
xor U8892 (N_8892,N_3293,N_2848);
xnor U8893 (N_8893,N_3713,N_2248);
nor U8894 (N_8894,N_2858,N_4794);
and U8895 (N_8895,N_3591,N_4702);
xor U8896 (N_8896,N_2280,N_2564);
or U8897 (N_8897,N_1804,N_3177);
xor U8898 (N_8898,N_2110,N_2839);
and U8899 (N_8899,N_1848,N_1509);
nor U8900 (N_8900,N_2289,N_4934);
or U8901 (N_8901,N_3780,N_2303);
nor U8902 (N_8902,N_877,N_4280);
or U8903 (N_8903,N_114,N_1787);
nand U8904 (N_8904,N_237,N_4758);
and U8905 (N_8905,N_28,N_407);
or U8906 (N_8906,N_2817,N_3943);
nand U8907 (N_8907,N_2304,N_3693);
nor U8908 (N_8908,N_760,N_3959);
nand U8909 (N_8909,N_683,N_485);
xnor U8910 (N_8910,N_2697,N_2688);
nand U8911 (N_8911,N_4643,N_488);
xor U8912 (N_8912,N_549,N_3338);
nor U8913 (N_8913,N_3173,N_3159);
nor U8914 (N_8914,N_4281,N_1688);
and U8915 (N_8915,N_3950,N_459);
and U8916 (N_8916,N_3533,N_3989);
or U8917 (N_8917,N_1375,N_1696);
nor U8918 (N_8918,N_2307,N_954);
nor U8919 (N_8919,N_536,N_4384);
xnor U8920 (N_8920,N_3387,N_2395);
xor U8921 (N_8921,N_1818,N_4484);
nor U8922 (N_8922,N_4412,N_1108);
nand U8923 (N_8923,N_236,N_754);
nand U8924 (N_8924,N_4475,N_699);
xor U8925 (N_8925,N_2929,N_1864);
nor U8926 (N_8926,N_615,N_1291);
nor U8927 (N_8927,N_745,N_2018);
or U8928 (N_8928,N_1660,N_4835);
nand U8929 (N_8929,N_3074,N_2180);
nor U8930 (N_8930,N_2078,N_2453);
nand U8931 (N_8931,N_4064,N_2558);
xor U8932 (N_8932,N_219,N_4139);
xor U8933 (N_8933,N_108,N_1561);
nand U8934 (N_8934,N_1750,N_4987);
or U8935 (N_8935,N_788,N_2940);
nand U8936 (N_8936,N_2864,N_2175);
and U8937 (N_8937,N_2219,N_4803);
xnor U8938 (N_8938,N_576,N_4139);
xnor U8939 (N_8939,N_2118,N_4676);
or U8940 (N_8940,N_2231,N_4399);
nor U8941 (N_8941,N_4566,N_1474);
or U8942 (N_8942,N_4145,N_4174);
or U8943 (N_8943,N_2016,N_1069);
xnor U8944 (N_8944,N_4575,N_1991);
or U8945 (N_8945,N_3797,N_559);
nand U8946 (N_8946,N_934,N_715);
and U8947 (N_8947,N_2190,N_3560);
or U8948 (N_8948,N_474,N_3895);
and U8949 (N_8949,N_913,N_1088);
and U8950 (N_8950,N_365,N_1003);
nand U8951 (N_8951,N_1090,N_4990);
or U8952 (N_8952,N_1892,N_4946);
nand U8953 (N_8953,N_638,N_300);
nor U8954 (N_8954,N_2764,N_1423);
nand U8955 (N_8955,N_1098,N_3247);
or U8956 (N_8956,N_4733,N_402);
or U8957 (N_8957,N_1658,N_2019);
and U8958 (N_8958,N_2837,N_1345);
or U8959 (N_8959,N_1730,N_1936);
and U8960 (N_8960,N_3147,N_407);
nor U8961 (N_8961,N_273,N_1590);
nand U8962 (N_8962,N_3972,N_2916);
nand U8963 (N_8963,N_1268,N_4451);
and U8964 (N_8964,N_2248,N_437);
nor U8965 (N_8965,N_905,N_3514);
nand U8966 (N_8966,N_1762,N_689);
xor U8967 (N_8967,N_2225,N_281);
xnor U8968 (N_8968,N_4698,N_4444);
or U8969 (N_8969,N_2728,N_367);
nand U8970 (N_8970,N_1922,N_1011);
or U8971 (N_8971,N_1492,N_1921);
xor U8972 (N_8972,N_3145,N_2188);
or U8973 (N_8973,N_1525,N_4848);
or U8974 (N_8974,N_4494,N_2802);
nand U8975 (N_8975,N_3768,N_3006);
nor U8976 (N_8976,N_3360,N_1113);
nand U8977 (N_8977,N_2550,N_46);
nor U8978 (N_8978,N_3158,N_2111);
nor U8979 (N_8979,N_1144,N_3477);
or U8980 (N_8980,N_15,N_2560);
nand U8981 (N_8981,N_1913,N_3367);
xnor U8982 (N_8982,N_557,N_3077);
and U8983 (N_8983,N_77,N_4920);
and U8984 (N_8984,N_2551,N_1615);
xnor U8985 (N_8985,N_2730,N_4491);
nor U8986 (N_8986,N_4423,N_4791);
nor U8987 (N_8987,N_594,N_4688);
and U8988 (N_8988,N_4803,N_4420);
or U8989 (N_8989,N_713,N_2967);
and U8990 (N_8990,N_1181,N_2097);
xnor U8991 (N_8991,N_4386,N_3250);
nor U8992 (N_8992,N_220,N_686);
nand U8993 (N_8993,N_2527,N_718);
nor U8994 (N_8994,N_39,N_1176);
or U8995 (N_8995,N_2848,N_2714);
or U8996 (N_8996,N_3753,N_1217);
nor U8997 (N_8997,N_725,N_3735);
nand U8998 (N_8998,N_3441,N_1548);
nor U8999 (N_8999,N_322,N_992);
nor U9000 (N_9000,N_2869,N_3930);
and U9001 (N_9001,N_4561,N_633);
or U9002 (N_9002,N_1928,N_2292);
or U9003 (N_9003,N_486,N_1907);
and U9004 (N_9004,N_3818,N_2980);
and U9005 (N_9005,N_4040,N_586);
nand U9006 (N_9006,N_3372,N_1590);
nor U9007 (N_9007,N_3885,N_4841);
nand U9008 (N_9008,N_2617,N_2727);
nor U9009 (N_9009,N_4452,N_2641);
xnor U9010 (N_9010,N_3950,N_272);
nor U9011 (N_9011,N_3541,N_1178);
nand U9012 (N_9012,N_3192,N_2893);
xnor U9013 (N_9013,N_3456,N_4505);
nand U9014 (N_9014,N_3231,N_1310);
nand U9015 (N_9015,N_682,N_1216);
and U9016 (N_9016,N_734,N_1463);
nor U9017 (N_9017,N_4508,N_2408);
xor U9018 (N_9018,N_4237,N_2004);
nand U9019 (N_9019,N_3484,N_2964);
and U9020 (N_9020,N_3073,N_2898);
or U9021 (N_9021,N_3521,N_3090);
nor U9022 (N_9022,N_4533,N_835);
nor U9023 (N_9023,N_3149,N_1539);
and U9024 (N_9024,N_1560,N_3348);
xor U9025 (N_9025,N_4831,N_4328);
xor U9026 (N_9026,N_4879,N_4904);
nand U9027 (N_9027,N_1674,N_3925);
or U9028 (N_9028,N_459,N_3896);
xor U9029 (N_9029,N_649,N_3277);
xnor U9030 (N_9030,N_3880,N_3676);
or U9031 (N_9031,N_2155,N_1029);
xnor U9032 (N_9032,N_675,N_544);
xor U9033 (N_9033,N_1532,N_1644);
nor U9034 (N_9034,N_4406,N_1269);
or U9035 (N_9035,N_2490,N_3941);
or U9036 (N_9036,N_4568,N_443);
or U9037 (N_9037,N_476,N_3036);
and U9038 (N_9038,N_667,N_3881);
nand U9039 (N_9039,N_127,N_4730);
nor U9040 (N_9040,N_4359,N_333);
or U9041 (N_9041,N_232,N_1428);
xnor U9042 (N_9042,N_3151,N_1956);
nand U9043 (N_9043,N_2505,N_993);
xor U9044 (N_9044,N_3162,N_167);
nor U9045 (N_9045,N_1015,N_3837);
and U9046 (N_9046,N_699,N_4306);
and U9047 (N_9047,N_3668,N_1341);
or U9048 (N_9048,N_3526,N_3561);
and U9049 (N_9049,N_2765,N_1384);
nand U9050 (N_9050,N_1140,N_3729);
nor U9051 (N_9051,N_1823,N_1000);
or U9052 (N_9052,N_4655,N_813);
nand U9053 (N_9053,N_3693,N_945);
and U9054 (N_9054,N_4698,N_2211);
and U9055 (N_9055,N_3401,N_2897);
nor U9056 (N_9056,N_4532,N_4759);
and U9057 (N_9057,N_4078,N_2274);
and U9058 (N_9058,N_2563,N_652);
or U9059 (N_9059,N_4783,N_323);
and U9060 (N_9060,N_1288,N_1239);
or U9061 (N_9061,N_1446,N_4818);
and U9062 (N_9062,N_1793,N_948);
nor U9063 (N_9063,N_1364,N_2130);
and U9064 (N_9064,N_541,N_2139);
nand U9065 (N_9065,N_3260,N_3917);
xnor U9066 (N_9066,N_2014,N_2943);
nand U9067 (N_9067,N_3716,N_1266);
or U9068 (N_9068,N_4964,N_3974);
or U9069 (N_9069,N_4766,N_3094);
nor U9070 (N_9070,N_451,N_615);
xnor U9071 (N_9071,N_2654,N_1993);
nor U9072 (N_9072,N_2645,N_2779);
nor U9073 (N_9073,N_3198,N_992);
nand U9074 (N_9074,N_3674,N_4082);
nor U9075 (N_9075,N_386,N_2547);
xnor U9076 (N_9076,N_1172,N_855);
or U9077 (N_9077,N_2401,N_4870);
nor U9078 (N_9078,N_82,N_3100);
nand U9079 (N_9079,N_1851,N_1474);
and U9080 (N_9080,N_4361,N_1595);
xor U9081 (N_9081,N_1766,N_3622);
and U9082 (N_9082,N_195,N_1004);
nand U9083 (N_9083,N_2873,N_474);
nand U9084 (N_9084,N_360,N_2322);
or U9085 (N_9085,N_3064,N_4251);
or U9086 (N_9086,N_4423,N_839);
nand U9087 (N_9087,N_2220,N_4220);
and U9088 (N_9088,N_348,N_52);
xnor U9089 (N_9089,N_1380,N_863);
nand U9090 (N_9090,N_2575,N_131);
nor U9091 (N_9091,N_4172,N_3300);
and U9092 (N_9092,N_3596,N_216);
nand U9093 (N_9093,N_2541,N_374);
xnor U9094 (N_9094,N_2510,N_1862);
or U9095 (N_9095,N_519,N_2833);
or U9096 (N_9096,N_2589,N_3779);
xor U9097 (N_9097,N_3619,N_2482);
or U9098 (N_9098,N_1574,N_1316);
nor U9099 (N_9099,N_4480,N_2707);
xnor U9100 (N_9100,N_2695,N_4147);
nand U9101 (N_9101,N_797,N_601);
nand U9102 (N_9102,N_1759,N_2069);
xnor U9103 (N_9103,N_1106,N_2398);
and U9104 (N_9104,N_1757,N_1720);
xor U9105 (N_9105,N_884,N_705);
nand U9106 (N_9106,N_4200,N_3419);
nor U9107 (N_9107,N_2710,N_3501);
nor U9108 (N_9108,N_2840,N_2061);
or U9109 (N_9109,N_579,N_543);
or U9110 (N_9110,N_436,N_1052);
nand U9111 (N_9111,N_3523,N_738);
xor U9112 (N_9112,N_2868,N_3247);
nand U9113 (N_9113,N_35,N_2567);
or U9114 (N_9114,N_2528,N_3258);
nand U9115 (N_9115,N_391,N_4882);
or U9116 (N_9116,N_1600,N_3032);
nor U9117 (N_9117,N_3593,N_3364);
or U9118 (N_9118,N_3908,N_4915);
xor U9119 (N_9119,N_649,N_2883);
or U9120 (N_9120,N_4943,N_3914);
xnor U9121 (N_9121,N_2112,N_1533);
or U9122 (N_9122,N_2376,N_220);
and U9123 (N_9123,N_612,N_3053);
nand U9124 (N_9124,N_4690,N_3757);
or U9125 (N_9125,N_1415,N_2917);
or U9126 (N_9126,N_1089,N_1567);
xor U9127 (N_9127,N_1913,N_1805);
and U9128 (N_9128,N_1015,N_4716);
or U9129 (N_9129,N_566,N_4697);
nor U9130 (N_9130,N_964,N_3986);
nand U9131 (N_9131,N_3450,N_3124);
or U9132 (N_9132,N_1830,N_1895);
xor U9133 (N_9133,N_3667,N_2759);
nand U9134 (N_9134,N_2692,N_1311);
and U9135 (N_9135,N_2179,N_2962);
or U9136 (N_9136,N_2884,N_4043);
nor U9137 (N_9137,N_1299,N_1749);
or U9138 (N_9138,N_2495,N_3470);
xor U9139 (N_9139,N_2101,N_995);
nor U9140 (N_9140,N_3754,N_3018);
nor U9141 (N_9141,N_175,N_535);
or U9142 (N_9142,N_4820,N_2066);
and U9143 (N_9143,N_3741,N_2411);
nand U9144 (N_9144,N_3625,N_656);
and U9145 (N_9145,N_444,N_1921);
xor U9146 (N_9146,N_3317,N_4781);
xnor U9147 (N_9147,N_2694,N_1995);
nand U9148 (N_9148,N_3974,N_3729);
or U9149 (N_9149,N_1005,N_3581);
nand U9150 (N_9150,N_1077,N_163);
nand U9151 (N_9151,N_2608,N_994);
xor U9152 (N_9152,N_680,N_3299);
xor U9153 (N_9153,N_1696,N_2633);
nor U9154 (N_9154,N_4979,N_1363);
xnor U9155 (N_9155,N_4067,N_918);
and U9156 (N_9156,N_3045,N_4562);
nor U9157 (N_9157,N_2453,N_4172);
nor U9158 (N_9158,N_3773,N_2168);
xor U9159 (N_9159,N_3484,N_1436);
nor U9160 (N_9160,N_4168,N_2711);
and U9161 (N_9161,N_534,N_4704);
nand U9162 (N_9162,N_4594,N_388);
nand U9163 (N_9163,N_1296,N_1117);
nor U9164 (N_9164,N_4142,N_4707);
or U9165 (N_9165,N_4669,N_916);
xnor U9166 (N_9166,N_567,N_4737);
and U9167 (N_9167,N_3700,N_1192);
and U9168 (N_9168,N_4545,N_3478);
nor U9169 (N_9169,N_3191,N_3945);
or U9170 (N_9170,N_333,N_2517);
and U9171 (N_9171,N_4959,N_1191);
and U9172 (N_9172,N_2082,N_321);
and U9173 (N_9173,N_4846,N_4906);
and U9174 (N_9174,N_1565,N_252);
or U9175 (N_9175,N_4875,N_942);
nand U9176 (N_9176,N_3978,N_3344);
nand U9177 (N_9177,N_3599,N_1272);
nand U9178 (N_9178,N_4825,N_4233);
xnor U9179 (N_9179,N_708,N_1342);
nand U9180 (N_9180,N_2154,N_353);
xor U9181 (N_9181,N_569,N_2409);
nand U9182 (N_9182,N_2328,N_272);
nand U9183 (N_9183,N_4089,N_4060);
nor U9184 (N_9184,N_3496,N_2258);
nand U9185 (N_9185,N_1211,N_957);
and U9186 (N_9186,N_1630,N_1984);
xnor U9187 (N_9187,N_1059,N_4172);
nor U9188 (N_9188,N_1684,N_931);
nor U9189 (N_9189,N_4581,N_1315);
and U9190 (N_9190,N_2181,N_3936);
nor U9191 (N_9191,N_1358,N_51);
or U9192 (N_9192,N_544,N_3897);
or U9193 (N_9193,N_1768,N_2831);
or U9194 (N_9194,N_4905,N_3843);
and U9195 (N_9195,N_4886,N_1491);
nand U9196 (N_9196,N_1314,N_2238);
nand U9197 (N_9197,N_456,N_4243);
nor U9198 (N_9198,N_2288,N_340);
nand U9199 (N_9199,N_1477,N_620);
xor U9200 (N_9200,N_2266,N_2222);
nand U9201 (N_9201,N_4231,N_17);
or U9202 (N_9202,N_3446,N_3489);
or U9203 (N_9203,N_1109,N_3331);
and U9204 (N_9204,N_4754,N_2865);
nand U9205 (N_9205,N_3728,N_3992);
and U9206 (N_9206,N_3418,N_2985);
nand U9207 (N_9207,N_1216,N_2291);
or U9208 (N_9208,N_4121,N_307);
nand U9209 (N_9209,N_454,N_4593);
nand U9210 (N_9210,N_1792,N_3747);
nor U9211 (N_9211,N_4753,N_156);
nor U9212 (N_9212,N_1710,N_4952);
nor U9213 (N_9213,N_995,N_509);
or U9214 (N_9214,N_4124,N_4349);
or U9215 (N_9215,N_2405,N_2736);
nand U9216 (N_9216,N_2648,N_2183);
xor U9217 (N_9217,N_3320,N_3860);
and U9218 (N_9218,N_1532,N_4618);
or U9219 (N_9219,N_1242,N_3178);
nand U9220 (N_9220,N_4182,N_2819);
and U9221 (N_9221,N_3875,N_4732);
nor U9222 (N_9222,N_751,N_1600);
or U9223 (N_9223,N_2919,N_1581);
or U9224 (N_9224,N_4296,N_788);
and U9225 (N_9225,N_1391,N_1435);
xnor U9226 (N_9226,N_492,N_4841);
and U9227 (N_9227,N_2688,N_2528);
or U9228 (N_9228,N_1770,N_4030);
nor U9229 (N_9229,N_2753,N_858);
nor U9230 (N_9230,N_4854,N_3708);
nand U9231 (N_9231,N_4940,N_4223);
or U9232 (N_9232,N_1798,N_1585);
nor U9233 (N_9233,N_4607,N_527);
nand U9234 (N_9234,N_4567,N_276);
xnor U9235 (N_9235,N_1033,N_1355);
nand U9236 (N_9236,N_440,N_159);
nand U9237 (N_9237,N_4187,N_2133);
xnor U9238 (N_9238,N_2758,N_2652);
nand U9239 (N_9239,N_3354,N_4564);
nor U9240 (N_9240,N_639,N_1846);
nand U9241 (N_9241,N_3597,N_1262);
and U9242 (N_9242,N_2641,N_4998);
nand U9243 (N_9243,N_225,N_4490);
and U9244 (N_9244,N_1253,N_4473);
and U9245 (N_9245,N_17,N_1784);
nand U9246 (N_9246,N_2633,N_4298);
and U9247 (N_9247,N_3424,N_1022);
or U9248 (N_9248,N_3108,N_3278);
or U9249 (N_9249,N_4396,N_857);
or U9250 (N_9250,N_3062,N_2206);
and U9251 (N_9251,N_3416,N_3392);
or U9252 (N_9252,N_202,N_728);
and U9253 (N_9253,N_23,N_4922);
nor U9254 (N_9254,N_1889,N_456);
and U9255 (N_9255,N_3836,N_3967);
or U9256 (N_9256,N_3142,N_2438);
nor U9257 (N_9257,N_2236,N_3082);
xor U9258 (N_9258,N_1122,N_4353);
or U9259 (N_9259,N_1691,N_2134);
nor U9260 (N_9260,N_842,N_837);
xor U9261 (N_9261,N_2526,N_1976);
and U9262 (N_9262,N_4733,N_1976);
or U9263 (N_9263,N_774,N_380);
or U9264 (N_9264,N_998,N_713);
and U9265 (N_9265,N_2811,N_1430);
nor U9266 (N_9266,N_3003,N_4410);
xnor U9267 (N_9267,N_3017,N_3611);
xor U9268 (N_9268,N_2920,N_1011);
nand U9269 (N_9269,N_3437,N_3559);
xnor U9270 (N_9270,N_887,N_3640);
nand U9271 (N_9271,N_1443,N_4996);
xor U9272 (N_9272,N_1586,N_2035);
and U9273 (N_9273,N_363,N_115);
or U9274 (N_9274,N_3072,N_2372);
or U9275 (N_9275,N_2536,N_4206);
and U9276 (N_9276,N_3978,N_2421);
and U9277 (N_9277,N_1219,N_4561);
and U9278 (N_9278,N_2778,N_1775);
or U9279 (N_9279,N_84,N_4583);
and U9280 (N_9280,N_2296,N_4364);
or U9281 (N_9281,N_4227,N_2521);
nand U9282 (N_9282,N_4190,N_3809);
xor U9283 (N_9283,N_2019,N_3942);
or U9284 (N_9284,N_4205,N_426);
or U9285 (N_9285,N_2858,N_3513);
and U9286 (N_9286,N_3091,N_4713);
nor U9287 (N_9287,N_4850,N_1844);
nand U9288 (N_9288,N_177,N_4595);
nor U9289 (N_9289,N_2049,N_4089);
nand U9290 (N_9290,N_38,N_4957);
nor U9291 (N_9291,N_4460,N_3132);
or U9292 (N_9292,N_1183,N_651);
or U9293 (N_9293,N_2408,N_2011);
nand U9294 (N_9294,N_2081,N_608);
nand U9295 (N_9295,N_2988,N_1029);
nand U9296 (N_9296,N_2873,N_1896);
or U9297 (N_9297,N_3947,N_1434);
nor U9298 (N_9298,N_3595,N_2466);
nand U9299 (N_9299,N_1440,N_463);
and U9300 (N_9300,N_283,N_1802);
nand U9301 (N_9301,N_2267,N_1331);
xor U9302 (N_9302,N_585,N_2484);
or U9303 (N_9303,N_1302,N_3294);
xor U9304 (N_9304,N_1805,N_4533);
and U9305 (N_9305,N_4748,N_4542);
or U9306 (N_9306,N_1432,N_453);
nor U9307 (N_9307,N_249,N_2324);
or U9308 (N_9308,N_2508,N_2519);
and U9309 (N_9309,N_2672,N_2095);
or U9310 (N_9310,N_1071,N_4203);
nand U9311 (N_9311,N_538,N_3467);
and U9312 (N_9312,N_3614,N_0);
nor U9313 (N_9313,N_1943,N_219);
nor U9314 (N_9314,N_2160,N_3502);
nand U9315 (N_9315,N_4453,N_1268);
nand U9316 (N_9316,N_1737,N_3444);
and U9317 (N_9317,N_3786,N_1232);
and U9318 (N_9318,N_4105,N_1618);
nor U9319 (N_9319,N_952,N_3709);
or U9320 (N_9320,N_3868,N_3017);
or U9321 (N_9321,N_2333,N_231);
xnor U9322 (N_9322,N_1909,N_2732);
nand U9323 (N_9323,N_237,N_1010);
nand U9324 (N_9324,N_472,N_2062);
xor U9325 (N_9325,N_1723,N_3031);
and U9326 (N_9326,N_1547,N_2761);
and U9327 (N_9327,N_1935,N_1505);
nor U9328 (N_9328,N_4771,N_4776);
or U9329 (N_9329,N_3631,N_835);
nor U9330 (N_9330,N_1946,N_2583);
nor U9331 (N_9331,N_358,N_1859);
nor U9332 (N_9332,N_612,N_746);
nand U9333 (N_9333,N_684,N_4725);
nor U9334 (N_9334,N_3344,N_4956);
nor U9335 (N_9335,N_1666,N_803);
nor U9336 (N_9336,N_2930,N_1762);
and U9337 (N_9337,N_4382,N_769);
nand U9338 (N_9338,N_3794,N_4450);
or U9339 (N_9339,N_2567,N_2770);
nand U9340 (N_9340,N_2682,N_1793);
and U9341 (N_9341,N_1387,N_3795);
nor U9342 (N_9342,N_150,N_544);
or U9343 (N_9343,N_4403,N_271);
nand U9344 (N_9344,N_1036,N_723);
xnor U9345 (N_9345,N_2806,N_2758);
nand U9346 (N_9346,N_4780,N_3826);
and U9347 (N_9347,N_4560,N_3079);
and U9348 (N_9348,N_235,N_4514);
nand U9349 (N_9349,N_4524,N_2923);
xnor U9350 (N_9350,N_3449,N_3932);
or U9351 (N_9351,N_4706,N_3);
nor U9352 (N_9352,N_721,N_1377);
xor U9353 (N_9353,N_403,N_4797);
nor U9354 (N_9354,N_624,N_1399);
or U9355 (N_9355,N_3984,N_131);
and U9356 (N_9356,N_4177,N_334);
nor U9357 (N_9357,N_4845,N_3714);
nor U9358 (N_9358,N_2694,N_3492);
nand U9359 (N_9359,N_3048,N_2372);
nand U9360 (N_9360,N_510,N_2183);
and U9361 (N_9361,N_3391,N_3462);
nor U9362 (N_9362,N_868,N_1506);
and U9363 (N_9363,N_3360,N_1084);
nor U9364 (N_9364,N_4770,N_3165);
or U9365 (N_9365,N_2690,N_4418);
nand U9366 (N_9366,N_1787,N_4829);
and U9367 (N_9367,N_3933,N_1575);
nor U9368 (N_9368,N_1704,N_2429);
nor U9369 (N_9369,N_538,N_1365);
xnor U9370 (N_9370,N_1468,N_2850);
and U9371 (N_9371,N_153,N_236);
xor U9372 (N_9372,N_2103,N_3699);
nor U9373 (N_9373,N_4175,N_4283);
nand U9374 (N_9374,N_101,N_1303);
xnor U9375 (N_9375,N_3984,N_89);
nand U9376 (N_9376,N_4938,N_1104);
nand U9377 (N_9377,N_1713,N_3723);
xnor U9378 (N_9378,N_1483,N_3543);
xor U9379 (N_9379,N_1012,N_2086);
nand U9380 (N_9380,N_2635,N_77);
and U9381 (N_9381,N_4776,N_2339);
nor U9382 (N_9382,N_139,N_179);
or U9383 (N_9383,N_1208,N_4356);
xnor U9384 (N_9384,N_3430,N_4067);
nor U9385 (N_9385,N_526,N_4962);
nor U9386 (N_9386,N_914,N_2189);
xnor U9387 (N_9387,N_3107,N_3605);
and U9388 (N_9388,N_2928,N_1491);
and U9389 (N_9389,N_754,N_2227);
nand U9390 (N_9390,N_1529,N_2771);
nand U9391 (N_9391,N_4363,N_3906);
or U9392 (N_9392,N_385,N_3049);
or U9393 (N_9393,N_3346,N_980);
nand U9394 (N_9394,N_2395,N_2580);
nor U9395 (N_9395,N_3999,N_4888);
xor U9396 (N_9396,N_763,N_2728);
nor U9397 (N_9397,N_2174,N_1554);
xor U9398 (N_9398,N_66,N_2352);
and U9399 (N_9399,N_1082,N_3709);
and U9400 (N_9400,N_3077,N_4753);
and U9401 (N_9401,N_3445,N_1687);
nand U9402 (N_9402,N_1155,N_1164);
nand U9403 (N_9403,N_3597,N_4698);
nor U9404 (N_9404,N_2045,N_4354);
xor U9405 (N_9405,N_2389,N_4124);
and U9406 (N_9406,N_3641,N_2600);
xor U9407 (N_9407,N_1175,N_141);
nor U9408 (N_9408,N_2800,N_1798);
and U9409 (N_9409,N_4766,N_2174);
and U9410 (N_9410,N_3270,N_1819);
nand U9411 (N_9411,N_3404,N_3328);
or U9412 (N_9412,N_1826,N_4717);
or U9413 (N_9413,N_561,N_1305);
xnor U9414 (N_9414,N_4271,N_2144);
and U9415 (N_9415,N_1204,N_2917);
nor U9416 (N_9416,N_2822,N_1259);
or U9417 (N_9417,N_3528,N_59);
nand U9418 (N_9418,N_3541,N_2272);
or U9419 (N_9419,N_4245,N_1023);
nand U9420 (N_9420,N_2200,N_2623);
xor U9421 (N_9421,N_262,N_4188);
nand U9422 (N_9422,N_974,N_1389);
nor U9423 (N_9423,N_3189,N_4730);
and U9424 (N_9424,N_178,N_3218);
and U9425 (N_9425,N_3496,N_378);
and U9426 (N_9426,N_471,N_684);
xor U9427 (N_9427,N_3162,N_308);
nor U9428 (N_9428,N_4515,N_2564);
nor U9429 (N_9429,N_224,N_3954);
nor U9430 (N_9430,N_4249,N_1849);
nor U9431 (N_9431,N_4409,N_2474);
nand U9432 (N_9432,N_2998,N_1142);
or U9433 (N_9433,N_1439,N_1215);
nand U9434 (N_9434,N_1706,N_4437);
nor U9435 (N_9435,N_4839,N_842);
nand U9436 (N_9436,N_2319,N_1431);
and U9437 (N_9437,N_3879,N_4760);
or U9438 (N_9438,N_1828,N_3027);
nand U9439 (N_9439,N_3612,N_4041);
or U9440 (N_9440,N_68,N_1271);
or U9441 (N_9441,N_3027,N_4781);
and U9442 (N_9442,N_2822,N_1109);
nand U9443 (N_9443,N_372,N_2111);
nand U9444 (N_9444,N_891,N_142);
nand U9445 (N_9445,N_2997,N_3981);
nand U9446 (N_9446,N_3758,N_3717);
nor U9447 (N_9447,N_3492,N_2487);
nand U9448 (N_9448,N_1012,N_2442);
and U9449 (N_9449,N_2614,N_835);
and U9450 (N_9450,N_3401,N_4644);
nand U9451 (N_9451,N_389,N_4059);
nand U9452 (N_9452,N_1741,N_2030);
xor U9453 (N_9453,N_3152,N_2739);
nor U9454 (N_9454,N_3907,N_26);
or U9455 (N_9455,N_4765,N_2685);
or U9456 (N_9456,N_1210,N_2968);
and U9457 (N_9457,N_3334,N_619);
or U9458 (N_9458,N_4370,N_2951);
or U9459 (N_9459,N_2202,N_2115);
nor U9460 (N_9460,N_815,N_4286);
and U9461 (N_9461,N_1852,N_162);
nand U9462 (N_9462,N_4118,N_841);
nor U9463 (N_9463,N_599,N_2563);
and U9464 (N_9464,N_1684,N_3354);
nor U9465 (N_9465,N_3269,N_1692);
and U9466 (N_9466,N_637,N_4165);
and U9467 (N_9467,N_1109,N_3625);
xnor U9468 (N_9468,N_2931,N_3266);
xnor U9469 (N_9469,N_3192,N_2552);
nor U9470 (N_9470,N_1875,N_3478);
nor U9471 (N_9471,N_1630,N_2271);
nor U9472 (N_9472,N_1408,N_1556);
or U9473 (N_9473,N_3926,N_3649);
and U9474 (N_9474,N_3103,N_1913);
or U9475 (N_9475,N_3253,N_1498);
and U9476 (N_9476,N_1889,N_2953);
nand U9477 (N_9477,N_444,N_4400);
xor U9478 (N_9478,N_3126,N_3109);
or U9479 (N_9479,N_2138,N_1705);
and U9480 (N_9480,N_328,N_3303);
or U9481 (N_9481,N_2532,N_1476);
nand U9482 (N_9482,N_936,N_3096);
nand U9483 (N_9483,N_1026,N_1432);
nand U9484 (N_9484,N_1591,N_164);
or U9485 (N_9485,N_1386,N_115);
or U9486 (N_9486,N_1556,N_1509);
and U9487 (N_9487,N_2855,N_2120);
xnor U9488 (N_9488,N_4444,N_625);
xnor U9489 (N_9489,N_3052,N_665);
nor U9490 (N_9490,N_2630,N_3279);
or U9491 (N_9491,N_1506,N_847);
and U9492 (N_9492,N_1076,N_4110);
xnor U9493 (N_9493,N_2555,N_2044);
or U9494 (N_9494,N_4341,N_2880);
nor U9495 (N_9495,N_3600,N_3391);
and U9496 (N_9496,N_2732,N_955);
or U9497 (N_9497,N_3273,N_3418);
or U9498 (N_9498,N_4159,N_973);
and U9499 (N_9499,N_2494,N_4802);
xor U9500 (N_9500,N_383,N_1322);
or U9501 (N_9501,N_1464,N_400);
xor U9502 (N_9502,N_1820,N_2296);
nand U9503 (N_9503,N_2858,N_1736);
or U9504 (N_9504,N_1325,N_2110);
nor U9505 (N_9505,N_2105,N_1851);
nor U9506 (N_9506,N_2380,N_2356);
and U9507 (N_9507,N_4381,N_3010);
nor U9508 (N_9508,N_3201,N_4995);
or U9509 (N_9509,N_2293,N_1983);
nor U9510 (N_9510,N_3421,N_4732);
or U9511 (N_9511,N_3863,N_1684);
and U9512 (N_9512,N_4164,N_2859);
or U9513 (N_9513,N_4671,N_1422);
or U9514 (N_9514,N_3155,N_1564);
xnor U9515 (N_9515,N_3935,N_2967);
or U9516 (N_9516,N_347,N_806);
nand U9517 (N_9517,N_4571,N_2120);
xor U9518 (N_9518,N_4111,N_562);
or U9519 (N_9519,N_3856,N_2990);
or U9520 (N_9520,N_612,N_689);
and U9521 (N_9521,N_1462,N_3473);
nor U9522 (N_9522,N_4098,N_1677);
nor U9523 (N_9523,N_4535,N_2197);
nand U9524 (N_9524,N_2197,N_3229);
nand U9525 (N_9525,N_1069,N_2523);
and U9526 (N_9526,N_548,N_4876);
and U9527 (N_9527,N_3551,N_4458);
nand U9528 (N_9528,N_3069,N_2809);
and U9529 (N_9529,N_4572,N_1745);
nand U9530 (N_9530,N_1124,N_864);
nand U9531 (N_9531,N_3067,N_1590);
nor U9532 (N_9532,N_3807,N_1240);
or U9533 (N_9533,N_4133,N_2220);
nand U9534 (N_9534,N_4859,N_2306);
and U9535 (N_9535,N_3819,N_4013);
or U9536 (N_9536,N_4421,N_3363);
nand U9537 (N_9537,N_744,N_3985);
nor U9538 (N_9538,N_193,N_58);
nand U9539 (N_9539,N_4931,N_3879);
nor U9540 (N_9540,N_3026,N_3199);
and U9541 (N_9541,N_3492,N_794);
xnor U9542 (N_9542,N_1760,N_4033);
or U9543 (N_9543,N_3983,N_3826);
nor U9544 (N_9544,N_1333,N_3832);
or U9545 (N_9545,N_3770,N_1584);
or U9546 (N_9546,N_3547,N_1528);
nor U9547 (N_9547,N_1179,N_4866);
nor U9548 (N_9548,N_3281,N_3760);
nor U9549 (N_9549,N_3887,N_3549);
xor U9550 (N_9550,N_2904,N_3762);
or U9551 (N_9551,N_2578,N_3287);
and U9552 (N_9552,N_3849,N_3502);
and U9553 (N_9553,N_4038,N_2897);
nor U9554 (N_9554,N_652,N_959);
and U9555 (N_9555,N_1316,N_593);
xor U9556 (N_9556,N_1967,N_1438);
and U9557 (N_9557,N_3066,N_1551);
or U9558 (N_9558,N_92,N_2119);
xor U9559 (N_9559,N_2918,N_3918);
xnor U9560 (N_9560,N_2380,N_924);
and U9561 (N_9561,N_3656,N_1240);
nand U9562 (N_9562,N_2944,N_3);
nand U9563 (N_9563,N_522,N_4263);
nand U9564 (N_9564,N_881,N_4663);
or U9565 (N_9565,N_1642,N_2203);
nor U9566 (N_9566,N_2783,N_2490);
or U9567 (N_9567,N_3585,N_2172);
nor U9568 (N_9568,N_1818,N_2727);
nor U9569 (N_9569,N_549,N_3411);
xor U9570 (N_9570,N_4949,N_2150);
nor U9571 (N_9571,N_4469,N_1680);
or U9572 (N_9572,N_4585,N_2815);
and U9573 (N_9573,N_3930,N_1412);
nor U9574 (N_9574,N_3958,N_230);
xor U9575 (N_9575,N_2950,N_2351);
and U9576 (N_9576,N_4289,N_2463);
or U9577 (N_9577,N_4165,N_4095);
nand U9578 (N_9578,N_1520,N_757);
nand U9579 (N_9579,N_1770,N_3364);
xnor U9580 (N_9580,N_1962,N_2331);
and U9581 (N_9581,N_1049,N_369);
or U9582 (N_9582,N_854,N_2381);
and U9583 (N_9583,N_432,N_4805);
nand U9584 (N_9584,N_1057,N_1327);
and U9585 (N_9585,N_4515,N_1652);
and U9586 (N_9586,N_2250,N_1384);
nand U9587 (N_9587,N_3913,N_2756);
nor U9588 (N_9588,N_524,N_4400);
nand U9589 (N_9589,N_2124,N_4446);
or U9590 (N_9590,N_2466,N_3332);
nor U9591 (N_9591,N_3660,N_1309);
nand U9592 (N_9592,N_3528,N_3237);
xnor U9593 (N_9593,N_4370,N_2226);
nand U9594 (N_9594,N_2854,N_2730);
nand U9595 (N_9595,N_2530,N_2099);
and U9596 (N_9596,N_1693,N_4713);
nor U9597 (N_9597,N_1684,N_565);
and U9598 (N_9598,N_875,N_3415);
nor U9599 (N_9599,N_4037,N_736);
or U9600 (N_9600,N_3865,N_2689);
nand U9601 (N_9601,N_3566,N_2677);
xor U9602 (N_9602,N_697,N_2176);
xor U9603 (N_9603,N_585,N_1893);
xnor U9604 (N_9604,N_4422,N_2847);
nand U9605 (N_9605,N_829,N_2154);
and U9606 (N_9606,N_2461,N_2951);
nor U9607 (N_9607,N_3200,N_4853);
nor U9608 (N_9608,N_2391,N_4140);
or U9609 (N_9609,N_1158,N_4470);
or U9610 (N_9610,N_838,N_1000);
or U9611 (N_9611,N_2781,N_3423);
and U9612 (N_9612,N_2353,N_2365);
or U9613 (N_9613,N_683,N_3393);
nand U9614 (N_9614,N_632,N_4860);
xor U9615 (N_9615,N_1508,N_206);
and U9616 (N_9616,N_616,N_4398);
nor U9617 (N_9617,N_3309,N_978);
and U9618 (N_9618,N_4556,N_1868);
nor U9619 (N_9619,N_3561,N_3260);
and U9620 (N_9620,N_3188,N_4515);
and U9621 (N_9621,N_304,N_4907);
nand U9622 (N_9622,N_888,N_1472);
and U9623 (N_9623,N_1884,N_1578);
and U9624 (N_9624,N_3070,N_2784);
and U9625 (N_9625,N_617,N_2664);
nand U9626 (N_9626,N_2568,N_999);
xnor U9627 (N_9627,N_1092,N_4125);
nand U9628 (N_9628,N_48,N_3052);
or U9629 (N_9629,N_3103,N_4372);
or U9630 (N_9630,N_2540,N_2262);
nor U9631 (N_9631,N_1641,N_3965);
or U9632 (N_9632,N_173,N_2376);
nand U9633 (N_9633,N_2274,N_1658);
nand U9634 (N_9634,N_2125,N_3535);
nor U9635 (N_9635,N_2363,N_1839);
xnor U9636 (N_9636,N_926,N_2978);
or U9637 (N_9637,N_1197,N_2131);
xor U9638 (N_9638,N_4139,N_1419);
nor U9639 (N_9639,N_3240,N_794);
nor U9640 (N_9640,N_4665,N_1537);
and U9641 (N_9641,N_201,N_3639);
xnor U9642 (N_9642,N_570,N_2238);
xnor U9643 (N_9643,N_5,N_4647);
nor U9644 (N_9644,N_693,N_2035);
nor U9645 (N_9645,N_2084,N_4259);
xnor U9646 (N_9646,N_2642,N_2200);
nand U9647 (N_9647,N_2906,N_2464);
and U9648 (N_9648,N_1984,N_1247);
xnor U9649 (N_9649,N_893,N_4867);
and U9650 (N_9650,N_345,N_1736);
and U9651 (N_9651,N_3481,N_4408);
nor U9652 (N_9652,N_2310,N_3895);
nand U9653 (N_9653,N_4651,N_3966);
and U9654 (N_9654,N_1818,N_4784);
nand U9655 (N_9655,N_3000,N_570);
xnor U9656 (N_9656,N_2984,N_2256);
xor U9657 (N_9657,N_1060,N_837);
nand U9658 (N_9658,N_4176,N_3069);
xor U9659 (N_9659,N_1430,N_3388);
nor U9660 (N_9660,N_789,N_1936);
nand U9661 (N_9661,N_2443,N_132);
nand U9662 (N_9662,N_3044,N_3719);
xnor U9663 (N_9663,N_2065,N_625);
nand U9664 (N_9664,N_1457,N_1594);
and U9665 (N_9665,N_4376,N_4607);
nand U9666 (N_9666,N_2424,N_97);
or U9667 (N_9667,N_4966,N_2186);
nand U9668 (N_9668,N_3304,N_748);
or U9669 (N_9669,N_944,N_172);
nand U9670 (N_9670,N_821,N_35);
or U9671 (N_9671,N_4792,N_1821);
nand U9672 (N_9672,N_4943,N_1744);
and U9673 (N_9673,N_2900,N_1124);
or U9674 (N_9674,N_1682,N_4231);
and U9675 (N_9675,N_2719,N_3748);
nand U9676 (N_9676,N_4341,N_4827);
nand U9677 (N_9677,N_625,N_2277);
or U9678 (N_9678,N_2457,N_3062);
or U9679 (N_9679,N_3664,N_1416);
and U9680 (N_9680,N_2853,N_253);
nand U9681 (N_9681,N_1262,N_1575);
nor U9682 (N_9682,N_3086,N_4989);
or U9683 (N_9683,N_2671,N_3831);
and U9684 (N_9684,N_4750,N_3340);
nand U9685 (N_9685,N_3825,N_874);
nand U9686 (N_9686,N_3595,N_4913);
xor U9687 (N_9687,N_160,N_3482);
nor U9688 (N_9688,N_3850,N_2827);
nand U9689 (N_9689,N_2557,N_2963);
nand U9690 (N_9690,N_704,N_2948);
nand U9691 (N_9691,N_3577,N_2874);
nand U9692 (N_9692,N_4148,N_2585);
nor U9693 (N_9693,N_2702,N_2427);
nor U9694 (N_9694,N_528,N_2059);
and U9695 (N_9695,N_292,N_1852);
nand U9696 (N_9696,N_1947,N_356);
nor U9697 (N_9697,N_2073,N_2085);
and U9698 (N_9698,N_1062,N_4769);
or U9699 (N_9699,N_3080,N_431);
nand U9700 (N_9700,N_1551,N_2668);
and U9701 (N_9701,N_4073,N_4714);
nor U9702 (N_9702,N_2807,N_3025);
or U9703 (N_9703,N_1476,N_620);
or U9704 (N_9704,N_3360,N_732);
nand U9705 (N_9705,N_1258,N_1385);
and U9706 (N_9706,N_1345,N_1681);
and U9707 (N_9707,N_2179,N_1305);
and U9708 (N_9708,N_3990,N_4331);
xnor U9709 (N_9709,N_2721,N_3207);
or U9710 (N_9710,N_2562,N_2034);
and U9711 (N_9711,N_783,N_3499);
nand U9712 (N_9712,N_90,N_4634);
nor U9713 (N_9713,N_707,N_1367);
nor U9714 (N_9714,N_3520,N_2829);
or U9715 (N_9715,N_1038,N_4659);
xnor U9716 (N_9716,N_2617,N_3303);
xnor U9717 (N_9717,N_3639,N_1648);
and U9718 (N_9718,N_1178,N_2144);
nor U9719 (N_9719,N_2963,N_2143);
or U9720 (N_9720,N_2046,N_4162);
nor U9721 (N_9721,N_4593,N_2594);
nand U9722 (N_9722,N_3870,N_1752);
or U9723 (N_9723,N_2865,N_3336);
nor U9724 (N_9724,N_3940,N_4683);
or U9725 (N_9725,N_1652,N_2343);
xnor U9726 (N_9726,N_4136,N_322);
and U9727 (N_9727,N_3315,N_1454);
or U9728 (N_9728,N_4502,N_1222);
xor U9729 (N_9729,N_3697,N_3024);
nand U9730 (N_9730,N_1473,N_4460);
and U9731 (N_9731,N_4177,N_1257);
and U9732 (N_9732,N_341,N_2609);
nor U9733 (N_9733,N_1969,N_505);
nor U9734 (N_9734,N_2938,N_4383);
nand U9735 (N_9735,N_4213,N_3778);
or U9736 (N_9736,N_1063,N_2950);
nand U9737 (N_9737,N_4457,N_4884);
nand U9738 (N_9738,N_1399,N_2774);
or U9739 (N_9739,N_101,N_330);
nand U9740 (N_9740,N_4714,N_1356);
nor U9741 (N_9741,N_2299,N_3317);
or U9742 (N_9742,N_3406,N_162);
nand U9743 (N_9743,N_3261,N_1027);
or U9744 (N_9744,N_3314,N_419);
nor U9745 (N_9745,N_83,N_3471);
or U9746 (N_9746,N_4580,N_3867);
and U9747 (N_9747,N_494,N_1300);
xnor U9748 (N_9748,N_4529,N_3961);
and U9749 (N_9749,N_3249,N_1333);
nor U9750 (N_9750,N_2782,N_2901);
nand U9751 (N_9751,N_4545,N_4225);
xnor U9752 (N_9752,N_3145,N_2788);
and U9753 (N_9753,N_4609,N_4365);
xor U9754 (N_9754,N_440,N_4195);
nor U9755 (N_9755,N_138,N_4086);
nor U9756 (N_9756,N_1081,N_805);
nand U9757 (N_9757,N_3167,N_3159);
nand U9758 (N_9758,N_4844,N_3219);
nor U9759 (N_9759,N_658,N_2514);
xnor U9760 (N_9760,N_4594,N_1006);
xor U9761 (N_9761,N_10,N_279);
nand U9762 (N_9762,N_2885,N_2911);
xnor U9763 (N_9763,N_4443,N_1667);
nor U9764 (N_9764,N_2413,N_2650);
xor U9765 (N_9765,N_2139,N_2273);
nor U9766 (N_9766,N_529,N_4267);
or U9767 (N_9767,N_2266,N_414);
or U9768 (N_9768,N_3485,N_2941);
nand U9769 (N_9769,N_3380,N_1057);
xnor U9770 (N_9770,N_3627,N_3522);
or U9771 (N_9771,N_3732,N_1429);
nand U9772 (N_9772,N_419,N_4077);
and U9773 (N_9773,N_2112,N_3210);
xnor U9774 (N_9774,N_627,N_2265);
and U9775 (N_9775,N_3444,N_423);
or U9776 (N_9776,N_2682,N_2692);
or U9777 (N_9777,N_2854,N_4374);
and U9778 (N_9778,N_442,N_4731);
xnor U9779 (N_9779,N_256,N_1465);
or U9780 (N_9780,N_4687,N_3201);
nor U9781 (N_9781,N_2072,N_3037);
xnor U9782 (N_9782,N_3734,N_3013);
xor U9783 (N_9783,N_4264,N_1090);
xor U9784 (N_9784,N_2844,N_285);
nor U9785 (N_9785,N_3789,N_4986);
or U9786 (N_9786,N_2146,N_2238);
xnor U9787 (N_9787,N_4388,N_3652);
xnor U9788 (N_9788,N_4248,N_1114);
nand U9789 (N_9789,N_4470,N_1171);
and U9790 (N_9790,N_4695,N_3643);
or U9791 (N_9791,N_4499,N_4013);
or U9792 (N_9792,N_3803,N_647);
xnor U9793 (N_9793,N_3822,N_4553);
nor U9794 (N_9794,N_1034,N_4314);
nor U9795 (N_9795,N_4707,N_4440);
and U9796 (N_9796,N_3292,N_343);
nor U9797 (N_9797,N_900,N_2434);
or U9798 (N_9798,N_33,N_3072);
nand U9799 (N_9799,N_1963,N_4445);
nand U9800 (N_9800,N_1348,N_1674);
nor U9801 (N_9801,N_3254,N_3319);
nand U9802 (N_9802,N_668,N_4075);
or U9803 (N_9803,N_2712,N_4104);
nor U9804 (N_9804,N_4701,N_3658);
and U9805 (N_9805,N_2730,N_2357);
or U9806 (N_9806,N_4264,N_844);
or U9807 (N_9807,N_400,N_2876);
or U9808 (N_9808,N_1811,N_3441);
and U9809 (N_9809,N_3345,N_3875);
nand U9810 (N_9810,N_1523,N_1714);
and U9811 (N_9811,N_1720,N_1249);
or U9812 (N_9812,N_4461,N_4143);
or U9813 (N_9813,N_1829,N_4895);
nor U9814 (N_9814,N_4298,N_4335);
or U9815 (N_9815,N_1035,N_2517);
xnor U9816 (N_9816,N_989,N_423);
nand U9817 (N_9817,N_104,N_955);
or U9818 (N_9818,N_2766,N_2503);
nand U9819 (N_9819,N_4336,N_4430);
or U9820 (N_9820,N_4627,N_4900);
nand U9821 (N_9821,N_3767,N_1747);
nor U9822 (N_9822,N_3531,N_987);
or U9823 (N_9823,N_3834,N_367);
nor U9824 (N_9824,N_2236,N_4565);
and U9825 (N_9825,N_3521,N_1823);
or U9826 (N_9826,N_4840,N_52);
and U9827 (N_9827,N_321,N_1477);
nand U9828 (N_9828,N_2319,N_2091);
xor U9829 (N_9829,N_4117,N_2108);
or U9830 (N_9830,N_3934,N_848);
nor U9831 (N_9831,N_1866,N_1249);
nor U9832 (N_9832,N_2903,N_2763);
or U9833 (N_9833,N_2045,N_2597);
xor U9834 (N_9834,N_3085,N_462);
or U9835 (N_9835,N_3027,N_3655);
or U9836 (N_9836,N_1925,N_66);
nor U9837 (N_9837,N_1864,N_3860);
or U9838 (N_9838,N_3415,N_1141);
xnor U9839 (N_9839,N_2436,N_3210);
nand U9840 (N_9840,N_4534,N_4171);
xnor U9841 (N_9841,N_1134,N_62);
nand U9842 (N_9842,N_319,N_4938);
or U9843 (N_9843,N_135,N_4705);
nand U9844 (N_9844,N_417,N_1297);
nor U9845 (N_9845,N_3123,N_575);
and U9846 (N_9846,N_3309,N_2056);
xor U9847 (N_9847,N_2428,N_1739);
and U9848 (N_9848,N_864,N_3785);
or U9849 (N_9849,N_136,N_1661);
nor U9850 (N_9850,N_4094,N_4109);
xor U9851 (N_9851,N_3280,N_3304);
and U9852 (N_9852,N_855,N_649);
nor U9853 (N_9853,N_4253,N_1702);
nand U9854 (N_9854,N_4980,N_654);
or U9855 (N_9855,N_4411,N_4172);
xnor U9856 (N_9856,N_2101,N_4088);
or U9857 (N_9857,N_3509,N_4241);
nand U9858 (N_9858,N_3700,N_1792);
nand U9859 (N_9859,N_2118,N_2406);
and U9860 (N_9860,N_2654,N_195);
nor U9861 (N_9861,N_3889,N_3450);
nand U9862 (N_9862,N_1004,N_4077);
xnor U9863 (N_9863,N_2303,N_3757);
nor U9864 (N_9864,N_577,N_4134);
nor U9865 (N_9865,N_4089,N_2896);
and U9866 (N_9866,N_2691,N_602);
nor U9867 (N_9867,N_4911,N_2595);
nand U9868 (N_9868,N_2318,N_1856);
and U9869 (N_9869,N_3761,N_2307);
nand U9870 (N_9870,N_4304,N_3299);
nand U9871 (N_9871,N_710,N_3494);
xnor U9872 (N_9872,N_3860,N_1244);
nand U9873 (N_9873,N_3973,N_4025);
xnor U9874 (N_9874,N_3204,N_260);
and U9875 (N_9875,N_517,N_2360);
and U9876 (N_9876,N_3172,N_4394);
nand U9877 (N_9877,N_1427,N_3995);
and U9878 (N_9878,N_71,N_4591);
nor U9879 (N_9879,N_3711,N_3954);
and U9880 (N_9880,N_2734,N_917);
nand U9881 (N_9881,N_4770,N_898);
or U9882 (N_9882,N_3107,N_660);
and U9883 (N_9883,N_907,N_3232);
and U9884 (N_9884,N_4767,N_595);
or U9885 (N_9885,N_2435,N_3950);
nand U9886 (N_9886,N_869,N_2304);
and U9887 (N_9887,N_2062,N_2343);
or U9888 (N_9888,N_235,N_3203);
or U9889 (N_9889,N_4533,N_1204);
nand U9890 (N_9890,N_4725,N_2089);
xor U9891 (N_9891,N_2291,N_1750);
xnor U9892 (N_9892,N_3419,N_654);
and U9893 (N_9893,N_3919,N_1448);
xor U9894 (N_9894,N_905,N_981);
or U9895 (N_9895,N_1123,N_3011);
nand U9896 (N_9896,N_2773,N_4689);
xor U9897 (N_9897,N_994,N_2216);
nand U9898 (N_9898,N_3814,N_4111);
nand U9899 (N_9899,N_2709,N_1805);
xnor U9900 (N_9900,N_3808,N_709);
xor U9901 (N_9901,N_4562,N_3109);
nand U9902 (N_9902,N_2839,N_2120);
or U9903 (N_9903,N_3548,N_1784);
xor U9904 (N_9904,N_683,N_3334);
xor U9905 (N_9905,N_748,N_3292);
and U9906 (N_9906,N_2647,N_638);
and U9907 (N_9907,N_2051,N_84);
nand U9908 (N_9908,N_2670,N_1038);
nand U9909 (N_9909,N_2242,N_3005);
or U9910 (N_9910,N_3329,N_4007);
xnor U9911 (N_9911,N_2994,N_3822);
or U9912 (N_9912,N_224,N_2948);
or U9913 (N_9913,N_3188,N_2572);
and U9914 (N_9914,N_3792,N_813);
nor U9915 (N_9915,N_1130,N_3040);
nand U9916 (N_9916,N_767,N_4818);
and U9917 (N_9917,N_382,N_3415);
xor U9918 (N_9918,N_482,N_2738);
nor U9919 (N_9919,N_4239,N_3599);
xnor U9920 (N_9920,N_3559,N_1004);
nand U9921 (N_9921,N_1453,N_4751);
and U9922 (N_9922,N_2583,N_21);
and U9923 (N_9923,N_473,N_864);
nand U9924 (N_9924,N_1829,N_4885);
nor U9925 (N_9925,N_4120,N_1891);
xor U9926 (N_9926,N_4391,N_1930);
nand U9927 (N_9927,N_77,N_1011);
nand U9928 (N_9928,N_3846,N_74);
xnor U9929 (N_9929,N_2075,N_4801);
or U9930 (N_9930,N_1441,N_4335);
nor U9931 (N_9931,N_3731,N_2800);
and U9932 (N_9932,N_2855,N_3316);
nor U9933 (N_9933,N_1866,N_1683);
nor U9934 (N_9934,N_3853,N_2257);
or U9935 (N_9935,N_4390,N_753);
nor U9936 (N_9936,N_1152,N_2724);
nand U9937 (N_9937,N_4099,N_3031);
nand U9938 (N_9938,N_2349,N_3936);
nand U9939 (N_9939,N_1246,N_3854);
or U9940 (N_9940,N_2146,N_2090);
nand U9941 (N_9941,N_3807,N_572);
xor U9942 (N_9942,N_1140,N_3067);
nand U9943 (N_9943,N_2110,N_3246);
or U9944 (N_9944,N_1741,N_964);
nor U9945 (N_9945,N_102,N_336);
nor U9946 (N_9946,N_2437,N_990);
nand U9947 (N_9947,N_306,N_1911);
and U9948 (N_9948,N_4430,N_1398);
xnor U9949 (N_9949,N_938,N_2892);
nor U9950 (N_9950,N_1582,N_2388);
nor U9951 (N_9951,N_2863,N_1785);
xor U9952 (N_9952,N_470,N_2658);
and U9953 (N_9953,N_3396,N_4203);
nor U9954 (N_9954,N_3658,N_2562);
xnor U9955 (N_9955,N_4805,N_1624);
xnor U9956 (N_9956,N_3435,N_1029);
xor U9957 (N_9957,N_2009,N_4786);
and U9958 (N_9958,N_3740,N_2968);
nor U9959 (N_9959,N_4028,N_1395);
xnor U9960 (N_9960,N_1252,N_2206);
and U9961 (N_9961,N_4263,N_1227);
nand U9962 (N_9962,N_4843,N_4969);
nor U9963 (N_9963,N_3009,N_2214);
and U9964 (N_9964,N_1574,N_4157);
xor U9965 (N_9965,N_2605,N_4760);
nor U9966 (N_9966,N_2256,N_4001);
nor U9967 (N_9967,N_2453,N_2868);
or U9968 (N_9968,N_3309,N_1937);
nand U9969 (N_9969,N_2856,N_4200);
and U9970 (N_9970,N_3948,N_235);
nor U9971 (N_9971,N_1282,N_4314);
xnor U9972 (N_9972,N_737,N_1930);
nand U9973 (N_9973,N_3881,N_1357);
or U9974 (N_9974,N_2929,N_1625);
nor U9975 (N_9975,N_634,N_3116);
xnor U9976 (N_9976,N_4107,N_230);
and U9977 (N_9977,N_121,N_4396);
xnor U9978 (N_9978,N_1924,N_4319);
and U9979 (N_9979,N_400,N_4926);
nor U9980 (N_9980,N_3444,N_3418);
or U9981 (N_9981,N_4647,N_2944);
nand U9982 (N_9982,N_1221,N_1623);
nand U9983 (N_9983,N_4936,N_1224);
xnor U9984 (N_9984,N_1963,N_347);
xor U9985 (N_9985,N_3443,N_1181);
nor U9986 (N_9986,N_762,N_4532);
xnor U9987 (N_9987,N_3425,N_3088);
xnor U9988 (N_9988,N_4995,N_731);
nand U9989 (N_9989,N_1518,N_1184);
nand U9990 (N_9990,N_4527,N_2046);
nor U9991 (N_9991,N_1973,N_2799);
nand U9992 (N_9992,N_1786,N_4203);
and U9993 (N_9993,N_2352,N_4562);
nand U9994 (N_9994,N_3139,N_4232);
xor U9995 (N_9995,N_1129,N_2379);
or U9996 (N_9996,N_3602,N_819);
and U9997 (N_9997,N_4274,N_4220);
nand U9998 (N_9998,N_4196,N_2288);
nor U9999 (N_9999,N_4630,N_1811);
nand U10000 (N_10000,N_5616,N_6364);
xor U10001 (N_10001,N_7823,N_9668);
nand U10002 (N_10002,N_6868,N_9393);
or U10003 (N_10003,N_6897,N_9375);
and U10004 (N_10004,N_7241,N_7066);
and U10005 (N_10005,N_7646,N_8661);
xnor U10006 (N_10006,N_7091,N_8123);
or U10007 (N_10007,N_5738,N_7815);
or U10008 (N_10008,N_5190,N_9550);
or U10009 (N_10009,N_8958,N_7872);
xnor U10010 (N_10010,N_6863,N_8283);
xnor U10011 (N_10011,N_6590,N_5308);
nand U10012 (N_10012,N_6703,N_7858);
and U10013 (N_10013,N_5183,N_8370);
and U10014 (N_10014,N_9605,N_5194);
nor U10015 (N_10015,N_9299,N_5821);
or U10016 (N_10016,N_6041,N_6843);
nor U10017 (N_10017,N_9650,N_9178);
and U10018 (N_10018,N_6690,N_9994);
and U10019 (N_10019,N_5051,N_6930);
xor U10020 (N_10020,N_8048,N_5248);
and U10021 (N_10021,N_5346,N_5794);
nand U10022 (N_10022,N_8392,N_6666);
nand U10023 (N_10023,N_9621,N_7253);
and U10024 (N_10024,N_8256,N_8836);
or U10025 (N_10025,N_8638,N_7111);
nor U10026 (N_10026,N_5586,N_8291);
xnor U10027 (N_10027,N_7520,N_8645);
xor U10028 (N_10028,N_7916,N_7042);
xor U10029 (N_10029,N_9853,N_5438);
nand U10030 (N_10030,N_5154,N_6509);
nand U10031 (N_10031,N_7837,N_9790);
or U10032 (N_10032,N_9579,N_5459);
or U10033 (N_10033,N_8658,N_7511);
nand U10034 (N_10034,N_9279,N_5708);
nor U10035 (N_10035,N_8508,N_9627);
nor U10036 (N_10036,N_9754,N_6893);
nand U10037 (N_10037,N_7279,N_5709);
or U10038 (N_10038,N_9478,N_9339);
xnor U10039 (N_10039,N_7081,N_9047);
and U10040 (N_10040,N_8863,N_7730);
nor U10041 (N_10041,N_6224,N_5788);
or U10042 (N_10042,N_6844,N_6159);
xor U10043 (N_10043,N_8173,N_7099);
or U10044 (N_10044,N_5374,N_5676);
nor U10045 (N_10045,N_8434,N_6322);
or U10046 (N_10046,N_9821,N_5197);
nand U10047 (N_10047,N_6641,N_7806);
xor U10048 (N_10048,N_7501,N_8620);
xnor U10049 (N_10049,N_8980,N_5633);
or U10050 (N_10050,N_5536,N_6846);
nand U10051 (N_10051,N_9083,N_9543);
or U10052 (N_10052,N_6738,N_5960);
nor U10053 (N_10053,N_6866,N_6579);
xnor U10054 (N_10054,N_7365,N_5602);
nor U10055 (N_10055,N_7096,N_5978);
nand U10056 (N_10056,N_6188,N_9611);
nand U10057 (N_10057,N_9155,N_5664);
nand U10058 (N_10058,N_7764,N_9775);
xnor U10059 (N_10059,N_9298,N_5335);
xor U10060 (N_10060,N_8288,N_5947);
and U10061 (N_10061,N_8032,N_9004);
xor U10062 (N_10062,N_7483,N_7670);
and U10063 (N_10063,N_5205,N_9306);
or U10064 (N_10064,N_7804,N_5651);
nor U10065 (N_10065,N_5615,N_8947);
nor U10066 (N_10066,N_8720,N_9364);
or U10067 (N_10067,N_9494,N_7384);
nand U10068 (N_10068,N_5979,N_8169);
and U10069 (N_10069,N_6396,N_6565);
nand U10070 (N_10070,N_9161,N_6127);
nor U10071 (N_10071,N_7084,N_8581);
xor U10072 (N_10072,N_8678,N_8214);
xnor U10073 (N_10073,N_7197,N_5921);
nand U10074 (N_10074,N_9224,N_8106);
or U10075 (N_10075,N_6329,N_8549);
or U10076 (N_10076,N_6153,N_6348);
or U10077 (N_10077,N_9723,N_8145);
xnor U10078 (N_10078,N_8517,N_8026);
xnor U10079 (N_10079,N_6021,N_9071);
and U10080 (N_10080,N_9281,N_8896);
xor U10081 (N_10081,N_8150,N_5007);
and U10082 (N_10082,N_5109,N_9739);
nand U10083 (N_10083,N_6351,N_7246);
nor U10084 (N_10084,N_5299,N_5841);
or U10085 (N_10085,N_7614,N_9832);
and U10086 (N_10086,N_5677,N_6974);
nand U10087 (N_10087,N_7129,N_9244);
or U10088 (N_10088,N_9771,N_6786);
or U10089 (N_10089,N_7296,N_7628);
xnor U10090 (N_10090,N_7065,N_6085);
nor U10091 (N_10091,N_6493,N_8533);
and U10092 (N_10092,N_7106,N_6202);
nor U10093 (N_10093,N_7538,N_6649);
nor U10094 (N_10094,N_5722,N_7925);
nor U10095 (N_10095,N_8138,N_6507);
or U10096 (N_10096,N_8182,N_9219);
xor U10097 (N_10097,N_8418,N_9968);
and U10098 (N_10098,N_7401,N_7469);
nor U10099 (N_10099,N_7947,N_8276);
and U10100 (N_10100,N_7032,N_5010);
and U10101 (N_10101,N_5465,N_7105);
nor U10102 (N_10102,N_5257,N_8779);
nor U10103 (N_10103,N_8860,N_8194);
nor U10104 (N_10104,N_9574,N_8820);
xnor U10105 (N_10105,N_9795,N_5241);
or U10106 (N_10106,N_6244,N_7288);
nor U10107 (N_10107,N_8643,N_5713);
and U10108 (N_10108,N_6007,N_5175);
nand U10109 (N_10109,N_8243,N_6889);
and U10110 (N_10110,N_8640,N_9328);
or U10111 (N_10111,N_9370,N_8302);
nor U10112 (N_10112,N_9991,N_9756);
or U10113 (N_10113,N_8942,N_7229);
nor U10114 (N_10114,N_8295,N_5143);
xor U10115 (N_10115,N_8659,N_7585);
xnor U10116 (N_10116,N_5034,N_6559);
nor U10117 (N_10117,N_8475,N_9648);
nor U10118 (N_10118,N_9144,N_5188);
xnor U10119 (N_10119,N_9384,N_5811);
nor U10120 (N_10120,N_5720,N_6789);
nor U10121 (N_10121,N_8814,N_6157);
nand U10122 (N_10122,N_6773,N_6618);
nor U10123 (N_10123,N_7829,N_6129);
or U10124 (N_10124,N_7661,N_8227);
xor U10125 (N_10125,N_7172,N_9742);
nand U10126 (N_10126,N_5988,N_9410);
or U10127 (N_10127,N_7880,N_5648);
xor U10128 (N_10128,N_6324,N_8154);
nor U10129 (N_10129,N_5073,N_7617);
xnor U10130 (N_10130,N_8927,N_9691);
or U10131 (N_10131,N_6241,N_7681);
or U10132 (N_10132,N_5661,N_7844);
nand U10133 (N_10133,N_9662,N_6549);
nand U10134 (N_10134,N_8285,N_7783);
or U10135 (N_10135,N_9861,N_9072);
and U10136 (N_10136,N_6810,N_8776);
nand U10137 (N_10137,N_6087,N_8058);
or U10138 (N_10138,N_6546,N_6708);
or U10139 (N_10139,N_5642,N_6270);
xor U10140 (N_10140,N_8151,N_5965);
and U10141 (N_10141,N_7315,N_7388);
nor U10142 (N_10142,N_8985,N_5525);
and U10143 (N_10143,N_9931,N_8849);
nand U10144 (N_10144,N_9522,N_8299);
xor U10145 (N_10145,N_6246,N_8641);
and U10146 (N_10146,N_7843,N_9198);
nand U10147 (N_10147,N_6170,N_6382);
nor U10148 (N_10148,N_9115,N_9342);
xnor U10149 (N_10149,N_5009,N_9718);
and U10150 (N_10150,N_8529,N_6257);
nand U10151 (N_10151,N_6659,N_6199);
xnor U10152 (N_10152,N_9194,N_8868);
xor U10153 (N_10153,N_9055,N_8359);
or U10154 (N_10154,N_9112,N_5543);
or U10155 (N_10155,N_5488,N_9639);
nor U10156 (N_10156,N_6760,N_7284);
and U10157 (N_10157,N_8363,N_5740);
nand U10158 (N_10158,N_7849,N_5723);
nand U10159 (N_10159,N_7326,N_8694);
or U10160 (N_10160,N_7477,N_7125);
nor U10161 (N_10161,N_5022,N_7860);
and U10162 (N_10162,N_9831,N_8818);
nor U10163 (N_10163,N_9466,N_8371);
and U10164 (N_10164,N_8767,N_7881);
or U10165 (N_10165,N_9946,N_8937);
xor U10166 (N_10166,N_8401,N_7295);
and U10167 (N_10167,N_7252,N_5231);
nor U10168 (N_10168,N_6342,N_6055);
nand U10169 (N_10169,N_5414,N_6823);
or U10170 (N_10170,N_5354,N_5214);
nand U10171 (N_10171,N_5927,N_8085);
or U10172 (N_10172,N_8551,N_7878);
nand U10173 (N_10173,N_9439,N_7020);
or U10174 (N_10174,N_6784,N_9473);
and U10175 (N_10175,N_5731,N_7183);
nand U10176 (N_10176,N_8804,N_6671);
and U10177 (N_10177,N_9493,N_8773);
nand U10178 (N_10178,N_6992,N_8059);
nand U10179 (N_10179,N_7821,N_8925);
xor U10180 (N_10180,N_8778,N_8889);
nor U10181 (N_10181,N_6265,N_8611);
nor U10182 (N_10182,N_8630,N_5773);
or U10183 (N_10183,N_6636,N_6336);
nand U10184 (N_10184,N_6478,N_6563);
nor U10185 (N_10185,N_6280,N_5764);
xor U10186 (N_10186,N_7165,N_6395);
xnor U10187 (N_10187,N_8156,N_6793);
nor U10188 (N_10188,N_8725,N_6061);
and U10189 (N_10189,N_9955,N_8916);
or U10190 (N_10190,N_6256,N_5429);
nor U10191 (N_10191,N_9412,N_8130);
xnor U10192 (N_10192,N_9699,N_6997);
nand U10193 (N_10193,N_6327,N_5858);
nand U10194 (N_10194,N_6417,N_6587);
and U10195 (N_10195,N_7798,N_7046);
nand U10196 (N_10196,N_9916,N_5765);
or U10197 (N_10197,N_8041,N_5587);
nand U10198 (N_10198,N_8167,N_6027);
nand U10199 (N_10199,N_6093,N_7859);
nor U10200 (N_10200,N_5932,N_5402);
or U10201 (N_10201,N_6956,N_7009);
nand U10202 (N_10202,N_5182,N_9360);
or U10203 (N_10203,N_5513,N_5917);
or U10204 (N_10204,N_6068,N_5741);
nand U10205 (N_10205,N_8310,N_9406);
xnor U10206 (N_10206,N_8437,N_5327);
nand U10207 (N_10207,N_8988,N_5215);
nor U10208 (N_10208,N_8764,N_5044);
or U10209 (N_10209,N_9894,N_5233);
xor U10210 (N_10210,N_5127,N_6536);
nand U10211 (N_10211,N_6436,N_5385);
or U10212 (N_10212,N_8189,N_9285);
xnor U10213 (N_10213,N_9864,N_9401);
or U10214 (N_10214,N_9845,N_6491);
nand U10215 (N_10215,N_7177,N_6977);
nand U10216 (N_10216,N_8811,N_7170);
nand U10217 (N_10217,N_9638,N_7069);
xor U10218 (N_10218,N_7067,N_6980);
and U10219 (N_10219,N_7431,N_5454);
or U10220 (N_10220,N_8729,N_9247);
xnor U10221 (N_10221,N_5470,N_7885);
or U10222 (N_10222,N_6473,N_7529);
and U10223 (N_10223,N_7694,N_9836);
or U10224 (N_10224,N_9202,N_8448);
xnor U10225 (N_10225,N_9517,N_7795);
nand U10226 (N_10226,N_7800,N_7915);
nand U10227 (N_10227,N_8409,N_6313);
xor U10228 (N_10228,N_6943,N_6171);
nand U10229 (N_10229,N_5992,N_6923);
xnor U10230 (N_10230,N_6539,N_8352);
nand U10231 (N_10231,N_6765,N_9231);
and U10232 (N_10232,N_6489,N_8629);
nand U10233 (N_10233,N_6573,N_7419);
nor U10234 (N_10234,N_9180,N_8618);
nand U10235 (N_10235,N_9906,N_8415);
xor U10236 (N_10236,N_8692,N_9663);
or U10237 (N_10237,N_9168,N_7713);
and U10238 (N_10238,N_6919,N_5165);
xnor U10239 (N_10239,N_9600,N_6450);
or U10240 (N_10240,N_7932,N_9307);
xnor U10241 (N_10241,N_7438,N_7963);
and U10242 (N_10242,N_6301,N_8364);
and U10243 (N_10243,N_5972,N_7191);
xor U10244 (N_10244,N_6854,N_7593);
nor U10245 (N_10245,N_5578,N_5173);
xor U10246 (N_10246,N_7664,N_7350);
or U10247 (N_10247,N_6445,N_7826);
and U10248 (N_10248,N_6052,N_8915);
nor U10249 (N_10249,N_7648,N_6469);
or U10250 (N_10250,N_5592,N_7502);
nand U10251 (N_10251,N_8687,N_5029);
and U10252 (N_10252,N_8809,N_8148);
xnor U10253 (N_10253,N_7623,N_8520);
nor U10254 (N_10254,N_6936,N_7410);
and U10255 (N_10255,N_7397,N_9927);
nand U10256 (N_10256,N_5926,N_9564);
nand U10257 (N_10257,N_8003,N_7294);
xor U10258 (N_10258,N_9529,N_6970);
nor U10259 (N_10259,N_8344,N_5036);
or U10260 (N_10260,N_7396,N_8459);
xor U10261 (N_10261,N_5961,N_8757);
xor U10262 (N_10262,N_6277,N_7079);
xor U10263 (N_10263,N_7051,N_6219);
and U10264 (N_10264,N_6033,N_5956);
nand U10265 (N_10265,N_9726,N_6771);
nor U10266 (N_10266,N_5778,N_8708);
and U10267 (N_10267,N_6409,N_7185);
nand U10268 (N_10268,N_5389,N_5507);
or U10269 (N_10269,N_6963,N_8092);
nand U10270 (N_10270,N_7665,N_5087);
or U10271 (N_10271,N_8875,N_5047);
xor U10272 (N_10272,N_7848,N_6135);
or U10273 (N_10273,N_7235,N_7085);
and U10274 (N_10274,N_6133,N_9647);
and U10275 (N_10275,N_7220,N_5069);
xor U10276 (N_10276,N_9447,N_5432);
xnor U10277 (N_10277,N_6837,N_5902);
nand U10278 (N_10278,N_5546,N_9752);
nand U10279 (N_10279,N_5828,N_6415);
nand U10280 (N_10280,N_5099,N_8305);
xor U10281 (N_10281,N_9243,N_6185);
nand U10282 (N_10282,N_8460,N_6353);
xnor U10283 (N_10283,N_5762,N_7811);
and U10284 (N_10284,N_9254,N_7062);
or U10285 (N_10285,N_5217,N_6679);
or U10286 (N_10286,N_5845,N_6914);
and U10287 (N_10287,N_9892,N_6122);
nor U10288 (N_10288,N_8878,N_7583);
and U10289 (N_10289,N_7808,N_7472);
nand U10290 (N_10290,N_5319,N_5487);
xnor U10291 (N_10291,N_9373,N_8225);
nand U10292 (N_10292,N_7465,N_8530);
nand U10293 (N_10293,N_8356,N_6605);
and U10294 (N_10294,N_8810,N_8135);
nor U10295 (N_10295,N_5252,N_9914);
nor U10296 (N_10296,N_9460,N_5137);
and U10297 (N_10297,N_6315,N_7973);
or U10298 (N_10298,N_6676,N_6892);
xor U10299 (N_10299,N_5658,N_8709);
or U10300 (N_10300,N_8616,N_5976);
and U10301 (N_10301,N_5049,N_9264);
nor U10302 (N_10302,N_9278,N_5334);
nor U10303 (N_10303,N_7215,N_9901);
nor U10304 (N_10304,N_9037,N_9159);
or U10305 (N_10305,N_8568,N_7678);
and U10306 (N_10306,N_7600,N_6610);
and U10307 (N_10307,N_8541,N_8478);
nor U10308 (N_10308,N_9897,N_6000);
and U10309 (N_10309,N_5312,N_6288);
xnor U10310 (N_10310,N_9344,N_8715);
nor U10311 (N_10311,N_9998,N_5174);
nor U10312 (N_10312,N_5991,N_8991);
nand U10313 (N_10313,N_5259,N_8768);
and U10314 (N_10314,N_7506,N_7651);
xor U10315 (N_10315,N_8096,N_5830);
and U10316 (N_10316,N_9022,N_7072);
xnor U10317 (N_10317,N_6768,N_9365);
or U10318 (N_10318,N_9077,N_9727);
xor U10319 (N_10319,N_9800,N_8690);
xor U10320 (N_10320,N_8949,N_5311);
nand U10321 (N_10321,N_5056,N_5444);
xor U10322 (N_10322,N_7582,N_7936);
xnor U10323 (N_10323,N_9823,N_6700);
nor U10324 (N_10324,N_6849,N_8490);
nor U10325 (N_10325,N_5847,N_7176);
xnor U10326 (N_10326,N_5508,N_9050);
nor U10327 (N_10327,N_8657,N_5970);
xnor U10328 (N_10328,N_9875,N_7329);
xor U10329 (N_10329,N_8345,N_8296);
or U10330 (N_10330,N_8074,N_7425);
xnor U10331 (N_10331,N_8326,N_5887);
nor U10332 (N_10332,N_7918,N_6542);
nand U10333 (N_10333,N_7551,N_6207);
or U10334 (N_10334,N_6333,N_6780);
nand U10335 (N_10335,N_8236,N_6639);
nand U10336 (N_10336,N_5834,N_5472);
and U10337 (N_10337,N_7702,N_6574);
xnor U10338 (N_10338,N_6148,N_5735);
and U10339 (N_10339,N_5280,N_9965);
nand U10340 (N_10340,N_7910,N_7892);
xnor U10341 (N_10341,N_5761,N_7058);
xnor U10342 (N_10342,N_8978,N_7908);
or U10343 (N_10343,N_5160,N_7662);
and U10344 (N_10344,N_9733,N_6723);
xnor U10345 (N_10345,N_5679,N_5612);
and U10346 (N_10346,N_7059,N_6346);
xnor U10347 (N_10347,N_9415,N_7759);
nand U10348 (N_10348,N_6091,N_7328);
or U10349 (N_10349,N_6198,N_9534);
and U10350 (N_10350,N_5534,N_9936);
and U10351 (N_10351,N_5964,N_6370);
nor U10352 (N_10352,N_6448,N_5668);
and U10353 (N_10353,N_7792,N_9656);
nor U10354 (N_10354,N_5791,N_6883);
nand U10355 (N_10355,N_9961,N_6814);
nor U10356 (N_10356,N_7137,N_9569);
xor U10357 (N_10357,N_7642,N_5207);
xnor U10358 (N_10358,N_9720,N_5085);
nand U10359 (N_10359,N_6677,N_6907);
nand U10360 (N_10360,N_7930,N_9876);
nor U10361 (N_10361,N_6714,N_5732);
xor U10362 (N_10362,N_8405,N_9475);
xnor U10363 (N_10363,N_8484,N_9658);
and U10364 (N_10364,N_9948,N_7391);
nor U10365 (N_10365,N_5206,N_8064);
and U10366 (N_10366,N_6204,N_7337);
and U10367 (N_10367,N_5408,N_5061);
nand U10368 (N_10368,N_7610,N_8115);
and U10369 (N_10369,N_5570,N_9735);
nor U10370 (N_10370,N_8317,N_7174);
nand U10371 (N_10371,N_8321,N_7332);
xor U10372 (N_10372,N_5882,N_8632);
nand U10373 (N_10373,N_8396,N_6707);
nor U10374 (N_10374,N_5656,N_8582);
nor U10375 (N_10375,N_6358,N_9038);
and U10376 (N_10376,N_7960,N_6431);
or U10377 (N_10377,N_8120,N_5617);
nor U10378 (N_10378,N_9666,N_5296);
and U10379 (N_10379,N_6501,N_7970);
nor U10380 (N_10380,N_5219,N_9232);
xor U10381 (N_10381,N_5876,N_9282);
nand U10382 (N_10382,N_7978,N_5718);
nand U10383 (N_10383,N_5613,N_9438);
nor U10384 (N_10384,N_9670,N_7312);
and U10385 (N_10385,N_6177,N_7453);
xnor U10386 (N_10386,N_7727,N_7043);
and U10387 (N_10387,N_9069,N_6060);
or U10388 (N_10388,N_8728,N_6876);
and U10389 (N_10389,N_5637,N_8441);
and U10390 (N_10390,N_8457,N_7500);
xnor U10391 (N_10391,N_7117,N_9193);
xnor U10392 (N_10392,N_5624,N_8410);
nand U10393 (N_10393,N_6350,N_9690);
nand U10394 (N_10394,N_8511,N_5745);
xor U10395 (N_10395,N_5531,N_9111);
nor U10396 (N_10396,N_5383,N_5804);
nand U10397 (N_10397,N_8025,N_5697);
xnor U10398 (N_10398,N_9125,N_5321);
and U10399 (N_10399,N_7011,N_6123);
nand U10400 (N_10400,N_9164,N_7906);
or U10401 (N_10401,N_9429,N_7304);
or U10402 (N_10402,N_8885,N_9041);
nor U10403 (N_10403,N_8908,N_8261);
nor U10404 (N_10404,N_5685,N_6231);
xnor U10405 (N_10405,N_6744,N_8622);
and U10406 (N_10406,N_9082,N_6220);
xnor U10407 (N_10407,N_9986,N_7372);
nor U10408 (N_10408,N_6132,N_8801);
or U10409 (N_10409,N_7080,N_5524);
nand U10410 (N_10410,N_8018,N_7728);
xor U10411 (N_10411,N_9590,N_6235);
and U10412 (N_10412,N_6947,N_5148);
nand U10413 (N_10413,N_8432,N_5066);
or U10414 (N_10414,N_6067,N_6284);
xor U10415 (N_10415,N_5843,N_5393);
and U10416 (N_10416,N_5411,N_5377);
or U10417 (N_10417,N_7797,N_9979);
nand U10418 (N_10418,N_9330,N_9900);
nand U10419 (N_10419,N_5021,N_6236);
nand U10420 (N_10420,N_6142,N_9204);
and U10421 (N_10421,N_9549,N_9217);
xor U10422 (N_10422,N_7673,N_5144);
xor U10423 (N_10423,N_7088,N_9563);
and U10424 (N_10424,N_9815,N_5079);
or U10425 (N_10425,N_6102,N_6195);
and U10426 (N_10426,N_9970,N_5140);
nor U10427 (N_10427,N_7696,N_5116);
or U10428 (N_10428,N_9877,N_9284);
or U10429 (N_10429,N_6016,N_8900);
and U10430 (N_10430,N_9791,N_8703);
nor U10431 (N_10431,N_9486,N_9059);
xor U10432 (N_10432,N_6935,N_9043);
nor U10433 (N_10433,N_7534,N_8961);
xnor U10434 (N_10434,N_5103,N_8117);
and U10435 (N_10435,N_9613,N_7497);
nand U10436 (N_10436,N_9938,N_6733);
nor U10437 (N_10437,N_7112,N_7933);
or U10438 (N_10438,N_9435,N_6113);
xnor U10439 (N_10439,N_7367,N_5490);
nand U10440 (N_10440,N_5417,N_5567);
nor U10441 (N_10441,N_9332,N_5898);
nor U10442 (N_10442,N_7273,N_5118);
or U10443 (N_10443,N_7890,N_8770);
and U10444 (N_10444,N_7341,N_8919);
or U10445 (N_10445,N_7940,N_9758);
and U10446 (N_10446,N_9980,N_5938);
nand U10447 (N_10447,N_9822,N_5042);
nand U10448 (N_10448,N_9976,N_7034);
nand U10449 (N_10449,N_9102,N_8737);
or U10450 (N_10450,N_5657,N_6143);
nor U10451 (N_10451,N_6106,N_8635);
and U10452 (N_10452,N_7269,N_7958);
or U10453 (N_10453,N_7200,N_9380);
or U10454 (N_10454,N_6718,N_6483);
or U10455 (N_10455,N_8741,N_8452);
nand U10456 (N_10456,N_9567,N_9993);
nor U10457 (N_10457,N_5240,N_9424);
nand U10458 (N_10458,N_7285,N_6474);
nand U10459 (N_10459,N_7671,N_9709);
and U10460 (N_10460,N_5552,N_8497);
nor U10461 (N_10461,N_5598,N_9689);
xor U10462 (N_10462,N_6006,N_6108);
xor U10463 (N_10463,N_7943,N_5684);
nand U10464 (N_10464,N_5603,N_6926);
and U10465 (N_10465,N_9989,N_8921);
xor U10466 (N_10466,N_5006,N_7645);
or U10467 (N_10467,N_6971,N_7123);
nor U10468 (N_10468,N_9023,N_7619);
or U10469 (N_10469,N_5807,N_5704);
xnor U10470 (N_10470,N_7725,N_8023);
nor U10471 (N_10471,N_6233,N_7896);
and U10472 (N_10472,N_7173,N_7159);
nor U10473 (N_10473,N_8357,N_8290);
and U10474 (N_10474,N_9325,N_7711);
or U10475 (N_10475,N_8536,N_7983);
and U10476 (N_10476,N_7814,N_5885);
nor U10477 (N_10477,N_7008,N_6203);
nand U10478 (N_10478,N_8255,N_6857);
xor U10479 (N_10479,N_9988,N_9504);
xnor U10480 (N_10480,N_7109,N_5746);
and U10481 (N_10481,N_8580,N_6169);
nor U10482 (N_10482,N_6925,N_9628);
nand U10483 (N_10483,N_8572,N_6865);
nand U10484 (N_10484,N_7460,N_9857);
nor U10485 (N_10485,N_9222,N_5987);
xnor U10486 (N_10486,N_6341,N_5482);
and U10487 (N_10487,N_6609,N_8859);
xor U10488 (N_10488,N_8813,N_9665);
and U10489 (N_10489,N_9996,N_8205);
nand U10490 (N_10490,N_9408,N_9546);
xor U10491 (N_10491,N_8730,N_9766);
and U10492 (N_10492,N_6089,N_9007);
and U10493 (N_10493,N_7620,N_8748);
nor U10494 (N_10494,N_5645,N_9966);
nor U10495 (N_10495,N_5293,N_6529);
xor U10496 (N_10496,N_7423,N_9960);
or U10497 (N_10497,N_5663,N_8465);
xnor U10498 (N_10498,N_6140,N_8648);
nor U10499 (N_10499,N_7498,N_7937);
and U10500 (N_10500,N_9603,N_9964);
or U10501 (N_10501,N_8972,N_7461);
and U10502 (N_10502,N_5986,N_9065);
and U10503 (N_10503,N_5984,N_8506);
xor U10504 (N_10504,N_7692,N_6962);
or U10505 (N_10505,N_7274,N_6267);
or U10506 (N_10506,N_6896,N_7086);
nor U10507 (N_10507,N_6109,N_5258);
nor U10508 (N_10508,N_7602,N_5012);
and U10509 (N_10509,N_6081,N_9602);
or U10510 (N_10510,N_7190,N_9250);
or U10511 (N_10511,N_8537,N_8825);
nand U10512 (N_10512,N_5819,N_7090);
nor U10513 (N_10513,N_6804,N_5925);
xor U10514 (N_10514,N_6011,N_9283);
or U10515 (N_10515,N_8152,N_5519);
nand U10516 (N_10516,N_5413,N_9548);
and U10517 (N_10517,N_8176,N_6022);
nor U10518 (N_10518,N_9388,N_9465);
nand U10519 (N_10519,N_7095,N_6456);
or U10520 (N_10520,N_6015,N_6984);
nor U10521 (N_10521,N_5291,N_9188);
nor U10522 (N_10522,N_6187,N_5264);
or U10523 (N_10523,N_7522,N_8786);
and U10524 (N_10524,N_9308,N_5522);
nor U10525 (N_10525,N_6049,N_9502);
or U10526 (N_10526,N_9463,N_9228);
nand U10527 (N_10527,N_6019,N_6920);
nand U10528 (N_10528,N_9505,N_5798);
or U10529 (N_10529,N_8732,N_6205);
nor U10530 (N_10530,N_5200,N_8063);
and U10531 (N_10531,N_7688,N_6043);
nand U10532 (N_10532,N_6403,N_5147);
xor U10533 (N_10533,N_7243,N_5336);
or U10534 (N_10534,N_6924,N_7809);
nor U10535 (N_10535,N_6595,N_6310);
xor U10536 (N_10536,N_8042,N_7478);
xnor U10537 (N_10537,N_5721,N_8534);
and U10538 (N_10538,N_9664,N_5314);
nand U10539 (N_10539,N_6317,N_6264);
or U10540 (N_10540,N_7734,N_5046);
xnor U10541 (N_10541,N_5496,N_9848);
xnor U10542 (N_10542,N_9302,N_7984);
or U10543 (N_10543,N_5225,N_7537);
nand U10544 (N_10544,N_7803,N_6713);
xor U10545 (N_10545,N_5749,N_6410);
and U10546 (N_10546,N_9941,N_8716);
xor U10547 (N_10547,N_6512,N_7740);
or U10548 (N_10548,N_6615,N_5114);
and U10549 (N_10549,N_5427,N_6429);
nor U10550 (N_10550,N_6175,N_8979);
or U10551 (N_10551,N_9774,N_9196);
nor U10552 (N_10552,N_6819,N_6294);
nand U10553 (N_10553,N_9930,N_9782);
and U10554 (N_10554,N_5246,N_7268);
or U10555 (N_10555,N_9551,N_8734);
nor U10556 (N_10556,N_9451,N_8890);
xnor U10557 (N_10557,N_7709,N_7527);
or U10558 (N_10558,N_7475,N_6519);
nor U10559 (N_10559,N_5260,N_7061);
nand U10560 (N_10560,N_8610,N_5295);
nor U10561 (N_10561,N_6729,N_5348);
or U10562 (N_10562,N_9459,N_9987);
or U10563 (N_10563,N_9803,N_8938);
or U10564 (N_10564,N_5276,N_8793);
and U10565 (N_10565,N_6076,N_8104);
nor U10566 (N_10566,N_7309,N_7652);
xnor U10567 (N_10567,N_6128,N_9044);
xnor U10568 (N_10568,N_6413,N_6378);
xnor U10569 (N_10569,N_9745,N_6518);
or U10570 (N_10570,N_7975,N_5594);
nand U10571 (N_10571,N_9719,N_6162);
nor U10572 (N_10572,N_8078,N_7408);
xor U10573 (N_10573,N_7491,N_8114);
nand U10574 (N_10574,N_9838,N_7541);
xnor U10575 (N_10575,N_8411,N_9274);
xnor U10576 (N_10576,N_5665,N_6423);
xor U10577 (N_10577,N_5196,N_9508);
or U10578 (N_10578,N_8902,N_6062);
nor U10579 (N_10579,N_5908,N_7723);
nor U10580 (N_10580,N_6756,N_5686);
nand U10581 (N_10581,N_5134,N_5055);
nand U10582 (N_10582,N_6726,N_5895);
nor U10583 (N_10583,N_9187,N_9414);
nor U10584 (N_10584,N_7909,N_5981);
xor U10585 (N_10585,N_9345,N_7875);
xor U10586 (N_10586,N_5689,N_5418);
and U10587 (N_10587,N_9507,N_7189);
or U10588 (N_10588,N_7695,N_9552);
nor U10589 (N_10589,N_9352,N_7250);
nor U10590 (N_10590,N_5249,N_9311);
xnor U10591 (N_10591,N_6905,N_6394);
or U10592 (N_10592,N_7038,N_5262);
nand U10593 (N_10593,N_6477,N_5892);
xor U10594 (N_10594,N_7964,N_6800);
xnor U10595 (N_10595,N_9882,N_5511);
nor U10596 (N_10596,N_7802,N_5581);
nor U10597 (N_10597,N_5307,N_9437);
and U10598 (N_10598,N_7373,N_9696);
nand U10599 (N_10599,N_7627,N_7322);
nor U10600 (N_10600,N_5083,N_5434);
or U10601 (N_10601,N_5859,N_8639);
xnor U10602 (N_10602,N_5566,N_6100);
and U10603 (N_10603,N_5191,N_9367);
and U10604 (N_10604,N_9324,N_9619);
xor U10605 (N_10605,N_5093,N_9031);
nor U10606 (N_10606,N_8596,N_5779);
nor U10607 (N_10607,N_8772,N_6721);
xor U10608 (N_10608,N_7649,N_6065);
nand U10609 (N_10609,N_8160,N_9139);
nand U10610 (N_10610,N_5016,N_9954);
and U10611 (N_10611,N_5317,N_7140);
nand U10612 (N_10612,N_5384,N_9121);
or U10613 (N_10613,N_8052,N_7965);
nor U10614 (N_10614,N_9849,N_9098);
or U10615 (N_10615,N_5625,N_6759);
nor U10616 (N_10616,N_6432,N_9515);
nand U10617 (N_10617,N_7004,N_5285);
or U10618 (N_10618,N_7024,N_8808);
or U10619 (N_10619,N_8886,N_5382);
xnor U10620 (N_10620,N_7641,N_7476);
or U10621 (N_10621,N_7594,N_7624);
xor U10622 (N_10622,N_6444,N_8127);
xnor U10623 (N_10623,N_7083,N_5111);
and U10624 (N_10624,N_8547,N_5848);
and U10625 (N_10625,N_5705,N_6577);
nand U10626 (N_10626,N_8828,N_6885);
xnor U10627 (N_10627,N_5867,N_9675);
nand U10628 (N_10628,N_5469,N_7825);
xor U10629 (N_10629,N_9725,N_6331);
xnor U10630 (N_10630,N_5135,N_5652);
nand U10631 (N_10631,N_8469,N_9826);
nor U10632 (N_10632,N_9886,N_6748);
nor U10633 (N_10633,N_9858,N_6172);
or U10634 (N_10634,N_7346,N_5062);
or U10635 (N_10635,N_7644,N_8036);
nand U10636 (N_10636,N_8269,N_8487);
and U10637 (N_10637,N_8994,N_8867);
nand U10638 (N_10638,N_9394,N_5068);
or U10639 (N_10639,N_7758,N_7248);
xor U10640 (N_10640,N_9511,N_7632);
nand U10641 (N_10641,N_9801,N_9851);
nor U10642 (N_10642,N_8724,N_5614);
nand U10643 (N_10643,N_5670,N_5551);
nor U10644 (N_10644,N_8924,N_8525);
nand U10645 (N_10645,N_5201,N_9572);
xor U10646 (N_10646,N_5318,N_9715);
nor U10647 (N_10647,N_9476,N_6945);
nor U10648 (N_10648,N_6894,N_5862);
nand U10649 (N_10649,N_6497,N_9468);
nand U10650 (N_10650,N_9717,N_8824);
nor U10651 (N_10651,N_5700,N_6740);
nor U10652 (N_10652,N_8034,N_9506);
and U10653 (N_10653,N_8304,N_8119);
nand U10654 (N_10654,N_5541,N_8237);
and U10655 (N_10655,N_5903,N_8871);
and U10656 (N_10656,N_6482,N_8791);
and U10657 (N_10657,N_6875,N_7116);
xnor U10658 (N_10658,N_5410,N_6426);
nand U10659 (N_10659,N_7592,N_8598);
or U10660 (N_10660,N_6213,N_6937);
nand U10661 (N_10661,N_7584,N_6741);
xor U10662 (N_10662,N_6105,N_7138);
nor U10663 (N_10663,N_9501,N_6266);
and U10664 (N_10664,N_6226,N_7338);
xor U10665 (N_10665,N_6932,N_7544);
xnor U10666 (N_10666,N_8624,N_6228);
xnor U10667 (N_10667,N_9740,N_8262);
and U10668 (N_10668,N_5937,N_8505);
nor U10669 (N_10669,N_6737,N_5854);
or U10670 (N_10670,N_7251,N_6180);
xnor U10671 (N_10671,N_9266,N_8880);
nand U10672 (N_10672,N_7464,N_9166);
nor U10673 (N_10673,N_5883,N_7546);
nor U10674 (N_10674,N_5582,N_7639);
and U10675 (N_10675,N_5939,N_5888);
nor U10676 (N_10676,N_6416,N_5643);
nor U10677 (N_10677,N_5158,N_7416);
nor U10678 (N_10678,N_9444,N_6553);
or U10679 (N_10679,N_7041,N_9874);
nor U10680 (N_10680,N_5309,N_6138);
and U10681 (N_10681,N_7418,N_6825);
xnor U10682 (N_10682,N_9214,N_6345);
nor U10683 (N_10683,N_5662,N_5271);
nor U10684 (N_10684,N_7002,N_7409);
and U10685 (N_10685,N_5297,N_6107);
xnor U10686 (N_10686,N_9288,N_8858);
nand U10687 (N_10687,N_8492,N_8707);
nand U10688 (N_10688,N_9784,N_7368);
xor U10689 (N_10689,N_6098,N_8765);
or U10690 (N_10690,N_6096,N_9108);
nor U10691 (N_10691,N_9793,N_6428);
nand U10692 (N_10692,N_9070,N_8402);
or U10693 (N_10693,N_7959,N_5835);
nor U10694 (N_10694,N_5038,N_6347);
nand U10695 (N_10695,N_7778,N_6727);
xnor U10696 (N_10696,N_6906,N_5300);
xor U10697 (N_10697,N_8799,N_8670);
xnor U10698 (N_10698,N_7196,N_8368);
nand U10699 (N_10699,N_9385,N_6377);
xnor U10700 (N_10700,N_5366,N_5458);
nand U10701 (N_10701,N_8883,N_5754);
or U10702 (N_10702,N_6330,N_9481);
and U10703 (N_10703,N_5168,N_8588);
xor U10704 (N_10704,N_6717,N_8376);
or U10705 (N_10705,N_6619,N_6375);
xnor U10706 (N_10706,N_7413,N_7850);
nor U10707 (N_10707,N_9489,N_9432);
nor U10708 (N_10708,N_8240,N_8735);
nand U10709 (N_10709,N_6606,N_5405);
and U10710 (N_10710,N_7718,N_5274);
nand U10711 (N_10711,N_7982,N_6167);
or U10712 (N_10712,N_9992,N_6190);
and U10713 (N_10713,N_6523,N_5695);
nor U10714 (N_10714,N_9348,N_5744);
or U10715 (N_10715,N_6766,N_9134);
nand U10716 (N_10716,N_9834,N_6709);
xor U10717 (N_10717,N_7993,N_5237);
or U10718 (N_10718,N_7505,N_6785);
nand U10719 (N_10719,N_8324,N_8408);
nand U10720 (N_10720,N_9737,N_8473);
nor U10721 (N_10721,N_8830,N_6012);
nand U10722 (N_10722,N_6225,N_7863);
xor U10723 (N_10723,N_9918,N_7864);
and U10724 (N_10724,N_7929,N_7554);
xnor U10725 (N_10725,N_9655,N_9181);
and U10726 (N_10726,N_7298,N_8207);
nand U10727 (N_10727,N_5387,N_9702);
nor U10728 (N_10728,N_6869,N_6909);
xor U10729 (N_10729,N_9124,N_5373);
and U10730 (N_10730,N_9568,N_8543);
and U10731 (N_10731,N_7643,N_9387);
nand U10732 (N_10732,N_9555,N_9939);
nand U10733 (N_10733,N_6880,N_6467);
or U10734 (N_10734,N_7580,N_5315);
xor U10735 (N_10735,N_9982,N_6791);
nand U10736 (N_10736,N_8491,N_9674);
and U10737 (N_10737,N_5549,N_5717);
nand U10738 (N_10738,N_6398,N_8564);
nor U10739 (N_10739,N_6982,N_8573);
and U10740 (N_10740,N_7100,N_8854);
nand U10741 (N_10741,N_6693,N_9080);
nand U10742 (N_10742,N_9796,N_7357);
and U10743 (N_10743,N_5812,N_5226);
xor U10744 (N_10744,N_9580,N_5813);
or U10745 (N_10745,N_5039,N_5351);
or U10746 (N_10746,N_8252,N_9607);
nor U10747 (N_10747,N_7299,N_6287);
xor U10748 (N_10748,N_8468,N_9309);
nor U10749 (N_10749,N_8282,N_6155);
nor U10750 (N_10750,N_7640,N_8177);
nand U10751 (N_10751,N_7876,N_9184);
nand U10752 (N_10752,N_8733,N_8004);
and U10753 (N_10753,N_9079,N_6276);
and U10754 (N_10754,N_7221,N_5360);
xor U10755 (N_10755,N_5530,N_5946);
nor U10756 (N_10756,N_7674,N_5035);
xnor U10757 (N_10757,N_6003,N_5953);
or U10758 (N_10758,N_6360,N_7317);
or U10759 (N_10759,N_7587,N_7242);
nor U10760 (N_10760,N_7719,N_7870);
nand U10761 (N_10761,N_6071,N_9208);
nor U10762 (N_10762,N_8222,N_6407);
and U10763 (N_10763,N_6004,N_8646);
xnor U10764 (N_10764,N_8644,N_6210);
xor U10765 (N_10765,N_5714,N_6455);
nor U10766 (N_10766,N_6343,N_9383);
and U10767 (N_10767,N_8249,N_6604);
xnor U10768 (N_10768,N_7601,N_6039);
nor U10769 (N_10769,N_6859,N_8821);
xnor U10770 (N_10770,N_6273,N_8923);
and U10771 (N_10771,N_6758,N_9320);
nand U10772 (N_10772,N_9744,N_7131);
and U10773 (N_10773,N_8178,N_5400);
nand U10774 (N_10774,N_7363,N_7029);
and U10775 (N_10775,N_9837,N_8965);
and U10776 (N_10776,N_7575,N_8954);
xor U10777 (N_10777,N_9827,N_8518);
nand U10778 (N_10778,N_9119,N_5420);
and U10779 (N_10779,N_5537,N_6816);
and U10780 (N_10780,N_7939,N_5292);
or U10781 (N_10781,N_7791,N_6651);
nand U10782 (N_10782,N_6487,N_5577);
nand U10783 (N_10783,N_9855,N_7412);
nor U10784 (N_10784,N_8617,N_9313);
and U10785 (N_10785,N_9684,N_8390);
nand U10786 (N_10786,N_6886,N_5245);
nor U10787 (N_10787,N_5516,N_9780);
nor U10788 (N_10788,N_8327,N_9199);
or U10789 (N_10789,N_6163,N_9683);
nor U10790 (N_10790,N_8726,N_6433);
or U10791 (N_10791,N_5449,N_8973);
and U10792 (N_10792,N_6328,N_8170);
nor U10793 (N_10793,N_5020,N_6682);
nand U10794 (N_10794,N_7204,N_7003);
xor U10795 (N_10795,N_8014,N_7855);
or U10796 (N_10796,N_5120,N_7414);
nand U10797 (N_10797,N_7952,N_6629);
nand U10798 (N_10798,N_6571,N_7181);
xnor U10799 (N_10799,N_9218,N_6811);
nand U10800 (N_10800,N_8855,N_6362);
and U10801 (N_10801,N_7969,N_7167);
nand U10802 (N_10802,N_5952,N_8224);
xor U10803 (N_10803,N_8451,N_6388);
nor U10804 (N_10804,N_9730,N_7547);
nor U10805 (N_10805,N_9593,N_7135);
nor U10806 (N_10806,N_8552,N_8202);
or U10807 (N_10807,N_6083,N_7036);
xor U10808 (N_10808,N_5995,N_8312);
xor U10809 (N_10809,N_7240,N_5910);
and U10810 (N_10810,N_9078,N_9492);
or U10811 (N_10811,N_5263,N_7638);
xor U10812 (N_10812,N_5694,N_9286);
nor U10813 (N_10813,N_7883,N_7914);
xor U10814 (N_10814,N_9879,N_7160);
nand U10815 (N_10815,N_8203,N_7899);
or U10816 (N_10816,N_5730,N_7689);
and U10817 (N_10817,N_6385,N_5502);
nor U10818 (N_10818,N_9523,N_8727);
xnor U10819 (N_10819,N_8272,N_5894);
or U10820 (N_10820,N_8174,N_5907);
or U10821 (N_10821,N_5941,N_6576);
nand U10822 (N_10822,N_9539,N_7463);
nor U10823 (N_10823,N_5451,N_6608);
xor U10824 (N_10824,N_7449,N_8918);
nand U10825 (N_10825,N_6908,N_8917);
and U10826 (N_10826,N_8782,N_9926);
xnor U10827 (N_10827,N_5505,N_5924);
or U10828 (N_10828,N_6249,N_9430);
nor U10829 (N_10829,N_6181,N_6472);
xnor U10830 (N_10830,N_7494,N_7436);
nand U10831 (N_10831,N_9685,N_8936);
nor U10832 (N_10832,N_5660,N_8769);
and U10833 (N_10833,N_9895,N_7218);
nor U10834 (N_10834,N_8619,N_5871);
xor U10835 (N_10835,N_5313,N_6725);
xnor U10836 (N_10836,N_8436,N_9952);
and U10837 (N_10837,N_9708,N_9592);
nor U10838 (N_10838,N_6548,N_7443);
nand U10839 (N_10839,N_7578,N_6769);
and U10840 (N_10840,N_8996,N_7345);
xor U10841 (N_10841,N_5916,N_5906);
and U10842 (N_10842,N_7724,N_7006);
nand U10843 (N_10843,N_8028,N_7133);
nand U10844 (N_10844,N_5209,N_5222);
xnor U10845 (N_10845,N_6630,N_9748);
xor U10846 (N_10846,N_5452,N_7348);
or U10847 (N_10847,N_6505,N_8144);
or U10848 (N_10848,N_7810,N_8147);
and U10849 (N_10849,N_9787,N_8939);
or U10850 (N_10850,N_6533,N_7663);
xnor U10851 (N_10851,N_5901,N_5770);
nand U10852 (N_10852,N_7490,N_6134);
xnor U10853 (N_10853,N_7571,N_6451);
xnor U10854 (N_10854,N_9765,N_8585);
xor U10855 (N_10855,N_5386,N_5833);
nand U10856 (N_10856,N_6299,N_8606);
nand U10857 (N_10857,N_9483,N_5564);
xnor U10858 (N_10858,N_5971,N_5571);
and U10859 (N_10859,N_9958,N_5523);
nand U10860 (N_10860,N_6035,N_7213);
xor U10861 (N_10861,N_6670,N_7776);
nor U10862 (N_10862,N_9423,N_5786);
nor U10863 (N_10863,N_9749,N_9814);
xnor U10864 (N_10864,N_7721,N_8360);
nor U10865 (N_10865,N_8982,N_9346);
xor U10866 (N_10866,N_8131,N_5253);
or U10867 (N_10867,N_8211,N_9084);
and U10868 (N_10868,N_9586,N_7223);
nor U10869 (N_10869,N_9616,N_8971);
xnor U10870 (N_10870,N_9236,N_7745);
xnor U10871 (N_10871,N_7192,N_9226);
xnor U10872 (N_10872,N_6528,N_7087);
or U10873 (N_10873,N_9588,N_9922);
xnor U10874 (N_10874,N_8803,N_6151);
nor U10875 (N_10875,N_6969,N_8655);
nor U10876 (N_10876,N_9978,N_9212);
nor U10877 (N_10877,N_9951,N_7853);
nand U10878 (N_10878,N_9338,N_8171);
nor U10879 (N_10879,N_8608,N_6730);
nor U10880 (N_10880,N_6381,N_9141);
and U10881 (N_10881,N_9792,N_9323);
xnor U10882 (N_10882,N_8609,N_5439);
nor U10883 (N_10883,N_7974,N_7355);
nor U10884 (N_10884,N_8001,N_5478);
nor U10885 (N_10885,N_8446,N_9770);
nand U10886 (N_10886,N_7986,N_9956);
or U10887 (N_10887,N_6805,N_9585);
xor U10888 (N_10888,N_6453,N_8753);
nand U10889 (N_10889,N_5077,N_6904);
nand U10890 (N_10890,N_7166,N_9417);
nor U10891 (N_10891,N_9781,N_9053);
xnor U10892 (N_10892,N_9225,N_8380);
or U10893 (N_10893,N_9227,N_8253);
nor U10894 (N_10894,N_6626,N_5322);
or U10895 (N_10895,N_5088,N_7565);
and U10896 (N_10896,N_5221,N_9104);
and U10897 (N_10897,N_8740,N_9461);
nand U10898 (N_10898,N_6418,N_9025);
nand U10899 (N_10899,N_6544,N_7693);
nor U10900 (N_10900,N_7122,N_8935);
xor U10901 (N_10901,N_9259,N_9477);
or U10902 (N_10902,N_5748,N_8483);
xnor U10903 (N_10903,N_7180,N_5515);
nand U10904 (N_10904,N_9537,N_7270);
or U10905 (N_10905,N_9777,N_5529);
xnor U10906 (N_10906,N_5562,N_9703);
and U10907 (N_10907,N_6018,N_7590);
nand U10908 (N_10908,N_6510,N_9829);
or U10909 (N_10909,N_8081,N_9724);
or U10910 (N_10910,N_7417,N_7726);
nor U10911 (N_10911,N_7679,N_9706);
nand U10912 (N_10912,N_5653,N_6160);
xnor U10913 (N_10913,N_7316,N_7819);
or U10914 (N_10914,N_5878,N_5098);
and U10915 (N_10915,N_5681,N_7115);
xor U10916 (N_10916,N_8493,N_5985);
and U10917 (N_10917,N_9462,N_7566);
or U10918 (N_10918,N_9707,N_7612);
or U10919 (N_10919,N_8197,N_8933);
nor U10920 (N_10920,N_5013,N_6038);
and U10921 (N_10921,N_5498,N_9395);
nor U10922 (N_10922,N_8284,N_7330);
nor U10923 (N_10923,N_7576,N_6545);
nor U10924 (N_10924,N_6818,N_8070);
xor U10925 (N_10925,N_6412,N_9340);
nand U10926 (N_10926,N_6435,N_7247);
or U10927 (N_10927,N_7045,N_6050);
nand U10928 (N_10928,N_9911,N_9381);
nor U10929 (N_10929,N_5509,N_7824);
nor U10930 (N_10930,N_6369,N_9448);
nand U10931 (N_10931,N_5836,N_7754);
and U10932 (N_10932,N_8612,N_6156);
nor U10933 (N_10933,N_5569,N_5994);
xnor U10934 (N_10934,N_7277,N_6080);
and U10935 (N_10935,N_5287,N_5729);
nor U10936 (N_10936,N_9615,N_9148);
xnor U10937 (N_10937,N_7743,N_6503);
nand U10938 (N_10938,N_7622,N_7101);
or U10939 (N_10939,N_5122,N_9403);
nand U10940 (N_10940,N_8467,N_9290);
or U10941 (N_10941,N_9610,N_7056);
or U10942 (N_10942,N_6551,N_7118);
xor U10943 (N_10943,N_7387,N_9769);
nand U10944 (N_10944,N_9880,N_6890);
and U10945 (N_10945,N_8183,N_8652);
xnor U10946 (N_10946,N_6850,N_6036);
and U10947 (N_10947,N_6631,N_7482);
nand U10948 (N_10948,N_6488,N_7075);
xnor U10949 (N_10949,N_6292,N_5289);
or U10950 (N_10950,N_8819,N_5512);
xor U10951 (N_10951,N_5930,N_7254);
nor U10952 (N_10952,N_6521,N_5124);
nand U10953 (N_10953,N_9929,N_9878);
or U10954 (N_10954,N_9713,N_6637);
xnor U10955 (N_10955,N_5796,N_8404);
nand U10956 (N_10956,N_8292,N_9623);
nor U10957 (N_10957,N_7216,N_9625);
or U10958 (N_10958,N_6820,N_8986);
or U10959 (N_10959,N_6365,N_9400);
or U10960 (N_10960,N_9206,N_7716);
nand U10961 (N_10961,N_6598,N_5950);
xor U10962 (N_10962,N_6376,N_6645);
nor U10963 (N_10963,N_8318,N_7238);
nand U10964 (N_10964,N_6653,N_9464);
or U10965 (N_10965,N_8887,N_9779);
nor U10966 (N_10966,N_5627,N_6824);
nor U10967 (N_10967,N_5644,N_8289);
nand U10968 (N_10968,N_7706,N_6583);
xor U10969 (N_10969,N_9519,N_6379);
nand U10970 (N_10970,N_9176,N_9470);
xnor U10971 (N_10971,N_9135,N_9287);
nor U10972 (N_10972,N_5457,N_8009);
or U10973 (N_10973,N_5187,N_6591);
and U10974 (N_10974,N_7690,N_8983);
nor U10975 (N_10975,N_7018,N_5447);
or U10976 (N_10976,N_8242,N_7063);
nand U10977 (N_10977,N_6020,N_5483);
nand U10978 (N_10978,N_7378,N_7746);
and U10979 (N_10979,N_9977,N_5015);
or U10980 (N_10980,N_8097,N_7553);
nor U10981 (N_10981,N_9746,N_5996);
or U10982 (N_10982,N_8223,N_7715);
nand U10983 (N_10983,N_9441,N_9318);
and U10984 (N_10984,N_7919,N_6957);
and U10985 (N_10985,N_6699,N_8850);
or U10986 (N_10986,N_5874,N_5052);
xor U10987 (N_10987,N_8807,N_8743);
xnor U10988 (N_10988,N_9237,N_7898);
and U10989 (N_10989,N_6535,N_5017);
nand U10990 (N_10990,N_9641,N_7891);
xnor U10991 (N_10991,N_5028,N_7941);
nor U10992 (N_10992,N_6704,N_8636);
nand U10993 (N_10993,N_6665,N_9889);
nand U10994 (N_10994,N_6698,N_9015);
nor U10995 (N_10995,N_7184,N_6400);
and U10996 (N_10996,N_6297,N_9201);
and U10997 (N_10997,N_7336,N_9294);
or U10998 (N_10998,N_9912,N_7779);
nand U10999 (N_10999,N_8395,N_9215);
nor U11000 (N_11000,N_6686,N_6763);
and U11001 (N_11001,N_5698,N_7231);
nor U11002 (N_11002,N_8275,N_7325);
or U11003 (N_11003,N_9185,N_9538);
nand U11004 (N_11004,N_5958,N_7005);
nor U11005 (N_11005,N_9671,N_8153);
nand U11006 (N_11006,N_7548,N_8682);
and U11007 (N_11007,N_7540,N_7761);
xor U11008 (N_11008,N_6879,N_5989);
xnor U11009 (N_11009,N_8723,N_7922);
or U11010 (N_11010,N_6309,N_9830);
xor U11011 (N_11011,N_9189,N_8067);
nand U11012 (N_11012,N_6991,N_8334);
or U11013 (N_11013,N_6215,N_8604);
xor U11014 (N_11014,N_8865,N_6044);
and U11015 (N_11015,N_9626,N_6384);
or U11016 (N_11016,N_5203,N_7751);
nand U11017 (N_11017,N_7151,N_5806);
nor U11018 (N_11018,N_7647,N_5824);
nor U11019 (N_11019,N_8649,N_5433);
xor U11020 (N_11020,N_9736,N_5202);
and U11021 (N_11021,N_5846,N_7861);
or U11022 (N_11022,N_5962,N_9935);
nor U11023 (N_11023,N_7000,N_5324);
and U11024 (N_11024,N_5771,N_8847);
and U11025 (N_11025,N_6466,N_8677);
and U11026 (N_11026,N_7558,N_6492);
or U11027 (N_11027,N_6638,N_8674);
nor U11028 (N_11028,N_6513,N_9530);
nor U11029 (N_11029,N_6967,N_9527);
and U11030 (N_11030,N_7630,N_7905);
and U11031 (N_11031,N_6586,N_5279);
xor U11032 (N_11032,N_6298,N_6031);
xor U11033 (N_11033,N_7098,N_6870);
or U11034 (N_11034,N_9907,N_6339);
and U11035 (N_11035,N_9903,N_9583);
nor U11036 (N_11036,N_9272,N_7701);
and U11037 (N_11037,N_9371,N_7769);
xor U11038 (N_11038,N_9075,N_8546);
or U11039 (N_11039,N_6928,N_9404);
and U11040 (N_11040,N_6635,N_8882);
nand U11041 (N_11041,N_7873,N_6537);
or U11042 (N_11042,N_7531,N_5772);
xnor U11043 (N_11043,N_8749,N_8107);
or U11044 (N_11044,N_6147,N_6032);
nor U11045 (N_11045,N_5419,N_6597);
nand U11046 (N_11046,N_9868,N_8869);
nor U11047 (N_11047,N_6575,N_7403);
or U11048 (N_11048,N_6981,N_5707);
xor U11049 (N_11049,N_9110,N_9073);
or U11050 (N_11050,N_6770,N_5110);
xnor U11051 (N_11051,N_7770,N_6502);
nand U11052 (N_11052,N_9036,N_7741);
and U11053 (N_11053,N_8118,N_8191);
xnor U11054 (N_11054,N_7142,N_7481);
nor U11055 (N_11055,N_9866,N_8805);
nand U11056 (N_11056,N_9856,N_6867);
or U11057 (N_11057,N_7389,N_9127);
xnor U11058 (N_11058,N_9681,N_6150);
nand U11059 (N_11059,N_7871,N_8903);
nor U11060 (N_11060,N_6460,N_6821);
nand U11061 (N_11061,N_7426,N_8499);
nand U11062 (N_11062,N_7302,N_5966);
xnor U11063 (N_11063,N_5113,N_7308);
nand U11064 (N_11064,N_7164,N_8566);
xnor U11065 (N_11065,N_5604,N_6757);
nand U11066 (N_11066,N_5371,N_8852);
or U11067 (N_11067,N_5161,N_8424);
or U11068 (N_11068,N_7307,N_8273);
or U11069 (N_11069,N_9734,N_9067);
xor U11070 (N_11070,N_6702,N_9545);
nand U11071 (N_11071,N_9643,N_8998);
nor U11072 (N_11072,N_7816,N_7335);
xor U11073 (N_11073,N_7659,N_9557);
or U11074 (N_11074,N_5302,N_7842);
nor U11075 (N_11075,N_5171,N_7225);
and U11076 (N_11076,N_6827,N_7422);
and U11077 (N_11077,N_7153,N_8705);
and U11078 (N_11078,N_9452,N_7550);
nor U11079 (N_11079,N_6250,N_5065);
or U11080 (N_11080,N_8045,N_5506);
nand U11081 (N_11081,N_7618,N_9885);
nand U11082 (N_11082,N_6166,N_7430);
nand U11083 (N_11083,N_6103,N_8780);
nand U11084 (N_11084,N_5208,N_6623);
xnor U11085 (N_11085,N_9012,N_8400);
nand U11086 (N_11086,N_9617,N_6806);
nor U11087 (N_11087,N_5626,N_7327);
nand U11088 (N_11088,N_8238,N_7840);
or U11089 (N_11089,N_9376,N_8861);
and U11090 (N_11090,N_8679,N_7237);
xor U11091 (N_11091,N_7499,N_5002);
nor U11092 (N_11092,N_8200,N_9773);
nor U11093 (N_11093,N_9389,N_5691);
nand U11094 (N_11094,N_6779,N_7227);
nor U11095 (N_11095,N_9497,N_9509);
nand U11096 (N_11096,N_9357,N_7700);
or U11097 (N_11097,N_8721,N_5370);
and U11098 (N_11098,N_7579,N_9350);
xor U11099 (N_11099,N_9474,N_6034);
or U11100 (N_11100,N_6334,N_8069);
xnor U11101 (N_11101,N_5517,N_8347);
nand U11102 (N_11102,N_5184,N_7306);
xor U11103 (N_11103,N_8835,N_6209);
xor U11104 (N_11104,N_7283,N_9090);
xnor U11105 (N_11105,N_5139,N_9341);
xnor U11106 (N_11106,N_7990,N_7280);
nand U11107 (N_11107,N_5747,N_5595);
nor U11108 (N_11108,N_7893,N_5719);
xnor U11109 (N_11109,N_9928,N_5230);
and U11110 (N_11110,N_9392,N_8193);
and U11111 (N_11111,N_9654,N_9094);
and U11112 (N_11112,N_8035,N_5514);
or U11113 (N_11113,N_5556,N_8691);
nand U11114 (N_11114,N_8239,N_6692);
nor U11115 (N_11115,N_8186,N_7211);
xnor U11116 (N_11116,N_5040,N_5584);
and U11117 (N_11117,N_5967,N_6952);
nor U11118 (N_11118,N_7025,N_6189);
nor U11119 (N_11119,N_6557,N_8134);
nand U11120 (N_11120,N_5933,N_8656);
xor U11121 (N_11121,N_7404,N_9594);
xor U11122 (N_11122,N_6778,N_7733);
and U11123 (N_11123,N_8666,N_5875);
nor U11124 (N_11124,N_5969,N_6663);
or U11125 (N_11125,N_5286,N_9171);
and U11126 (N_11126,N_9056,N_7533);
and U11127 (N_11127,N_7265,N_6746);
and U11128 (N_11128,N_5711,N_9636);
nor U11129 (N_11129,N_7210,N_6295);
or U11130 (N_11130,N_8759,N_6137);
nor U11131 (N_11131,N_8862,N_6602);
xor U11132 (N_11132,N_5473,N_5381);
or U11133 (N_11133,N_7888,N_5618);
nor U11134 (N_11134,N_7782,N_7094);
nand U11135 (N_11135,N_9687,N_9547);
and U11136 (N_11136,N_8952,N_5667);
and U11137 (N_11137,N_5181,N_9416);
or U11138 (N_11138,N_8306,N_8230);
and U11139 (N_11139,N_7300,N_8628);
nor U11140 (N_11140,N_8259,N_6966);
xor U11141 (N_11141,N_8228,N_9409);
nor U11142 (N_11142,N_8823,N_6110);
or U11143 (N_11143,N_6525,N_5575);
xnor U11144 (N_11144,N_9854,N_9216);
nand U11145 (N_11145,N_5075,N_5123);
and U11146 (N_11146,N_5703,N_7015);
and U11147 (N_11147,N_6917,N_9514);
nand U11148 (N_11148,N_7992,N_8569);
or U11149 (N_11149,N_6976,N_6961);
and U11150 (N_11150,N_9152,N_8215);
or U11151 (N_11151,N_9100,N_8141);
or U11152 (N_11152,N_5131,N_7994);
xor U11153 (N_11153,N_5244,N_6938);
nand U11154 (N_11154,N_9757,N_6197);
xor U11155 (N_11155,N_6706,N_6278);
and U11156 (N_11156,N_8163,N_7048);
nor U11157 (N_11157,N_9839,N_6735);
nand U11158 (N_11158,N_7707,N_8962);
or U11159 (N_11159,N_7462,N_8522);
and U11160 (N_11160,N_5934,N_5983);
or U11161 (N_11161,N_5753,N_6005);
nor U11162 (N_11162,N_7515,N_6494);
and U11163 (N_11163,N_7152,N_5622);
nand U11164 (N_11164,N_9265,N_8101);
or U11165 (N_11165,N_9322,N_8165);
and U11166 (N_11166,N_5499,N_6842);
and U11167 (N_11167,N_8043,N_8394);
and U11168 (N_11168,N_8316,N_5095);
and U11169 (N_11169,N_5345,N_6275);
nor U11170 (N_11170,N_7950,N_5683);
nand U11171 (N_11171,N_9300,N_5929);
or U11172 (N_11172,N_9087,N_6126);
xnor U11173 (N_11173,N_8319,N_7657);
xor U11174 (N_11174,N_7496,N_5477);
or U11175 (N_11175,N_7987,N_6125);
nand U11176 (N_11176,N_5119,N_8665);
nor U11177 (N_11177,N_6912,N_5822);
or U11178 (N_11178,N_8265,N_9137);
or U11179 (N_11179,N_7053,N_5816);
or U11180 (N_11180,N_6898,N_5726);
xor U11181 (N_11181,N_8233,N_6515);
nand U11182 (N_11182,N_6534,N_9729);
nand U11183 (N_11183,N_7684,N_9910);
nand U11184 (N_11184,N_8474,N_5097);
or U11185 (N_11185,N_9693,N_7784);
xor U11186 (N_11186,N_9657,N_5769);
or U11187 (N_11187,N_8336,N_8449);
and U11188 (N_11188,N_7560,N_7877);
nand U11189 (N_11189,N_5254,N_6300);
nor U11190 (N_11190,N_5851,N_6078);
nor U11191 (N_11191,N_8963,N_9316);
xnor U11192 (N_11192,N_7712,N_5461);
nor U11193 (N_11193,N_6158,N_5588);
nor U11194 (N_11194,N_7710,N_6307);
and U11195 (N_11195,N_6978,N_9257);
nand U11196 (N_11196,N_7390,N_9997);
nand U11197 (N_11197,N_5437,N_9804);
nand U11198 (N_11198,N_5504,N_7625);
and U11199 (N_11199,N_5343,N_5880);
xor U11200 (N_11200,N_5826,N_8175);
and U11201 (N_11201,N_7073,N_8664);
nand U11202 (N_11202,N_9420,N_5376);
nand U11203 (N_11203,N_5255,N_7698);
nor U11204 (N_11204,N_5674,N_5235);
xor U11205 (N_11205,N_9743,N_9728);
xor U11206 (N_11206,N_9426,N_5805);
and U11207 (N_11207,N_6243,N_5955);
or U11208 (N_11208,N_9981,N_8354);
and U11209 (N_11209,N_9019,N_7291);
nor U11210 (N_11210,N_5421,N_9554);
or U11211 (N_11211,N_8766,N_9315);
or U11212 (N_11212,N_5998,N_6028);
and U11213 (N_11213,N_8597,N_5850);
and U11214 (N_11214,N_5401,N_8565);
and U11215 (N_11215,N_9358,N_6801);
nand U11216 (N_11216,N_7510,N_7862);
xor U11217 (N_11217,N_5579,N_6484);
xor U11218 (N_11218,N_5409,N_7371);
or U11219 (N_11219,N_7369,N_5108);
or U11220 (N_11220,N_8893,N_8633);
xor U11221 (N_11221,N_9118,N_7374);
nor U11222 (N_11222,N_7068,N_6739);
xnor U11223 (N_11223,N_5943,N_6344);
nor U11224 (N_11224,N_7259,N_5863);
or U11225 (N_11225,N_9446,N_9984);
and U11226 (N_11226,N_5787,N_5585);
and U11227 (N_11227,N_9485,N_6355);
nor U11228 (N_11228,N_6131,N_6056);
or U11229 (N_11229,N_5842,N_7492);
and U11230 (N_11230,N_6366,N_6640);
and U11231 (N_11231,N_6047,N_8020);
nor U11232 (N_11232,N_7035,N_7060);
and U11233 (N_11233,N_7382,N_6008);
nor U11234 (N_11234,N_6834,N_8932);
and U11235 (N_11235,N_8920,N_9262);
nand U11236 (N_11236,N_8447,N_6958);
or U11237 (N_11237,N_6987,N_9149);
xnor U11238 (N_11238,N_5340,N_7078);
nand U11239 (N_11239,N_6115,N_8946);
and U11240 (N_11240,N_6675,N_8842);
and U11241 (N_11241,N_6025,N_7320);
nand U11242 (N_11242,N_7411,N_9436);
nor U11243 (N_11243,N_5378,N_6084);
and U11244 (N_11244,N_7989,N_8503);
xnor U11245 (N_11245,N_5538,N_5350);
nand U11246 (N_11246,N_9909,N_8121);
nand U11247 (N_11247,N_5945,N_9454);
xor U11248 (N_11248,N_8831,N_8325);
and U11249 (N_11249,N_7292,N_5646);
nand U11250 (N_11250,N_6374,N_7513);
nor U11251 (N_11251,N_8515,N_6029);
or U11252 (N_11252,N_8526,N_5031);
nor U11253 (N_11253,N_7902,N_8373);
nand U11254 (N_11254,N_5105,N_7186);
nor U11255 (N_11255,N_8399,N_7954);
nor U11256 (N_11256,N_9377,N_7019);
nor U11257 (N_11257,N_9932,N_5860);
nand U11258 (N_11258,N_9536,N_9776);
nand U11259 (N_11259,N_5078,N_5692);
or U11260 (N_11260,N_6775,N_5565);
and U11261 (N_11261,N_5094,N_5316);
nor U11262 (N_11262,N_8075,N_6547);
xnor U11263 (N_11263,N_6251,N_5904);
nor U11264 (N_11264,N_6572,N_6621);
nor U11265 (N_11265,N_8212,N_8198);
nand U11266 (N_11266,N_7976,N_5936);
or U11267 (N_11267,N_6308,N_7206);
nand U11268 (N_11268,N_6490,N_5710);
nor U11269 (N_11269,N_8365,N_9863);
nand U11270 (N_11270,N_7017,N_7442);
or U11271 (N_11271,N_8422,N_8166);
nand U11272 (N_11272,N_7444,N_7033);
and U11273 (N_11273,N_9349,N_9697);
and U11274 (N_11274,N_9695,N_8696);
nor U11275 (N_11275,N_9146,N_7121);
xor U11276 (N_11276,N_7493,N_6554);
and U11277 (N_11277,N_6332,N_6941);
and U11278 (N_11278,N_6681,N_6026);
xnor U11279 (N_11279,N_5817,N_7377);
and U11280 (N_11280,N_6900,N_6731);
nor U11281 (N_11281,N_9934,N_8504);
nor U11282 (N_11282,N_6419,N_9531);
xnor U11283 (N_11283,N_8398,N_8829);
nand U11284 (N_11284,N_6933,N_6486);
xor U11285 (N_11285,N_7996,N_7057);
and U11286 (N_11286,N_9014,N_9632);
xor U11287 (N_11287,N_8355,N_9029);
nand U11288 (N_11288,N_5795,N_5445);
nand U11289 (N_11289,N_5601,N_8464);
nand U11290 (N_11290,N_8684,N_6506);
or U11291 (N_11291,N_8387,N_9013);
or U11292 (N_11292,N_7507,N_7528);
nand U11293 (N_11293,N_6476,N_7828);
and U11294 (N_11294,N_8164,N_8351);
xnor U11295 (N_11295,N_5800,N_8024);
or U11296 (N_11296,N_9597,N_5323);
nand U11297 (N_11297,N_5659,N_5832);
xnor U11298 (N_11298,N_5497,N_9490);
nor U11299 (N_11299,N_6667,N_7010);
nand U11300 (N_11300,N_6411,N_7154);
or U11301 (N_11301,N_6194,N_5533);
xnor U11302 (N_11302,N_8532,N_7903);
and U11303 (N_11303,N_5605,N_7767);
and U11304 (N_11304,N_5492,N_9794);
nand U11305 (N_11305,N_9809,N_9532);
or U11306 (N_11306,N_8683,N_7047);
nor U11307 (N_11307,N_5890,N_9937);
and U11308 (N_11308,N_5948,N_6408);
or U11309 (N_11309,N_7900,N_7729);
xor U11310 (N_11310,N_7607,N_9840);
or U11311 (N_11311,N_7343,N_9872);
nor U11312 (N_11312,N_9609,N_5597);
nor U11313 (N_11313,N_6669,N_5014);
nor U11314 (N_11314,N_9819,N_8625);
or U11315 (N_11315,N_6701,N_8201);
and U11316 (N_11316,N_6877,N_6948);
xnor U11317 (N_11317,N_6634,N_5224);
xnor U11318 (N_11318,N_8480,N_6479);
or U11319 (N_11319,N_5954,N_9612);
or U11320 (N_11320,N_8881,N_8022);
and U11321 (N_11321,N_7703,N_9762);
nand U11322 (N_11322,N_8328,N_6531);
and U11323 (N_11323,N_9898,N_5267);
nor U11324 (N_11324,N_8100,N_6206);
and U11325 (N_11325,N_9716,N_8562);
nor U11326 (N_11326,N_9378,N_9449);
xor U11327 (N_11327,N_9967,N_9560);
xnor U11328 (N_11328,N_7395,N_8462);
or U11329 (N_11329,N_5494,N_6079);
or U11330 (N_11330,N_6835,N_8974);
nor U11331 (N_11331,N_8248,N_7375);
or U11332 (N_11332,N_6051,N_5687);
and U11333 (N_11333,N_8970,N_9985);
and U11334 (N_11334,N_6164,N_8989);
xnor U11335 (N_11335,N_7474,N_6817);
and U11336 (N_11336,N_5220,N_8495);
xnor U11337 (N_11337,N_8669,N_6058);
and U11338 (N_11338,N_7924,N_6985);
nor U11339 (N_11339,N_6628,N_6200);
nand U11340 (N_11340,N_8960,N_8993);
xor U11341 (N_11341,N_8095,N_9785);
nor U11342 (N_11342,N_9329,N_8600);
and U11343 (N_11343,N_5128,N_7889);
xor U11344 (N_11344,N_8812,N_5922);
nor U11345 (N_11345,N_6777,N_7524);
xnor U11346 (N_11346,N_6392,N_7439);
nand U11347 (N_11347,N_8783,N_7485);
nor U11348 (N_11348,N_7832,N_8277);
nand U11349 (N_11349,N_8247,N_7044);
nor U11350 (N_11350,N_5150,N_9445);
or U11351 (N_11351,N_6464,N_9156);
and U11352 (N_11352,N_5060,N_7331);
nand U11353 (N_11353,N_6186,N_8062);
nand U11354 (N_11354,N_9573,N_7406);
or U11355 (N_11355,N_6691,N_5789);
nand U11356 (N_11356,N_6434,N_8758);
nor U11357 (N_11357,N_9778,N_7451);
or U11358 (N_11358,N_6318,N_7901);
nor U11359 (N_11359,N_8554,N_8848);
nand U11360 (N_11360,N_6661,N_7286);
nand U11361 (N_11361,N_9001,N_7911);
or U11362 (N_11362,N_7621,N_8651);
and U11363 (N_11363,N_5096,N_9054);
nor U11364 (N_11364,N_8792,N_7202);
and U11365 (N_11365,N_9113,N_7287);
and U11366 (N_11366,N_7731,N_5159);
xnor U11367 (N_11367,N_7467,N_6973);
nand U11368 (N_11368,N_9116,N_6767);
nand U11369 (N_11369,N_7352,N_5467);
or U11370 (N_11370,N_7786,N_6949);
or U11371 (N_11371,N_6660,N_5169);
xor U11372 (N_11372,N_5560,N_8093);
nand U11373 (N_11373,N_9584,N_9063);
xor U11374 (N_11374,N_5942,N_5380);
or U11375 (N_11375,N_9575,N_9253);
nand U11376 (N_11376,N_9661,N_5369);
nor U11377 (N_11377,N_5780,N_9526);
and U11378 (N_11378,N_6255,N_7126);
and U11379 (N_11379,N_8575,N_8287);
and U11380 (N_11380,N_5357,N_7780);
and U11381 (N_11381,N_5857,N_6192);
nor U11382 (N_11382,N_7456,N_7962);
or U11383 (N_11383,N_8377,N_5232);
and U11384 (N_11384,N_9397,N_7722);
or U11385 (N_11385,N_8550,N_5728);
xnor U11386 (N_11386,N_7680,N_8899);
nor U11387 (N_11387,N_5931,N_6442);
or U11388 (N_11388,N_9209,N_8263);
or U11389 (N_11389,N_9138,N_6001);
nand U11390 (N_11390,N_9319,N_8540);
nor U11391 (N_11391,N_8250,N_8739);
and U11392 (N_11392,N_5392,N_7845);
or U11393 (N_11393,N_5855,N_9917);
nor U11394 (N_11394,N_9343,N_9347);
nand U11395 (N_11395,N_8984,N_7504);
or U11396 (N_11396,N_5797,N_8146);
nand U11397 (N_11397,N_5303,N_6440);
or U11398 (N_11398,N_8775,N_7228);
and U11399 (N_11399,N_7319,N_7926);
and U11400 (N_11400,N_5100,N_5810);
nor U11401 (N_11401,N_5896,N_7434);
nand U11402 (N_11402,N_7907,N_5151);
or U11403 (N_11403,N_7653,N_7561);
xor U11404 (N_11404,N_5001,N_5980);
nor U11405 (N_11405,N_7921,N_7027);
nor U11406 (N_11406,N_6367,N_8542);
nor U11407 (N_11407,N_9871,N_5234);
or U11408 (N_11408,N_8527,N_5185);
and U11409 (N_11409,N_8798,N_6424);
or U11410 (N_11410,N_6500,N_9372);
nor U11411 (N_11411,N_6216,N_9402);
xor U11412 (N_11412,N_6581,N_6566);
or U11413 (N_11413,N_5464,N_8019);
and U11414 (N_11414,N_8901,N_8442);
xor U11415 (N_11415,N_5474,N_9369);
and U11416 (N_11416,N_8578,N_7424);
nor U11417 (N_11417,N_8744,N_8698);
nand U11418 (N_11418,N_6258,N_5540);
nand U11419 (N_11419,N_7574,N_9190);
nand U11420 (N_11420,N_8750,N_7851);
xor U11421 (N_11421,N_8301,N_8603);
xnor U11422 (N_11422,N_9289,N_8082);
xor U11423 (N_11423,N_8660,N_7399);
xnor U11424 (N_11424,N_5344,N_8056);
xnor U11425 (N_11425,N_9427,N_6999);
nand U11426 (N_11426,N_6380,N_7158);
xor U11427 (N_11427,N_5266,N_9652);
and U11428 (N_11428,N_6751,N_6499);
xnor U11429 (N_11429,N_7519,N_7749);
xor U11430 (N_11430,N_8105,N_6650);
and U11431 (N_11431,N_8702,N_6009);
xnor U11432 (N_11432,N_9405,N_7364);
xnor U11433 (N_11433,N_9682,N_9442);
or U11434 (N_11434,N_9088,N_7257);
nor U11435 (N_11435,N_5460,N_8907);
and U11436 (N_11436,N_7697,N_8512);
and U11437 (N_11437,N_6845,N_7049);
nor U11438 (N_11438,N_6279,N_5352);
or U11439 (N_11439,N_9245,N_9544);
nand U11440 (N_11440,N_6030,N_6338);
and U11441 (N_11441,N_7967,N_6217);
xor U11442 (N_11442,N_8593,N_6988);
and U11443 (N_11443,N_8421,N_5911);
xnor U11444 (N_11444,N_6953,N_8476);
xor U11445 (N_11445,N_9630,N_8999);
nand U11446 (N_11446,N_5072,N_7569);
nand U11447 (N_11447,N_8270,N_7516);
or U11448 (N_11448,N_5251,N_6796);
or U11449 (N_11449,N_6613,N_6437);
xnor U11450 (N_11450,N_8268,N_6689);
nand U11451 (N_11451,N_6214,N_5484);
or U11452 (N_11452,N_6734,N_7013);
or U11453 (N_11453,N_8403,N_8461);
nand U11454 (N_11454,N_5416,N_9553);
xor U11455 (N_11455,N_8433,N_7454);
nand U11456 (N_11456,N_7193,N_9487);
nand U11457 (N_11457,N_7774,N_5471);
or U11458 (N_11458,N_7486,N_6141);
nor U11459 (N_11459,N_9558,N_6596);
xnor U11460 (N_11460,N_7222,N_7144);
nand U11461 (N_11461,N_8647,N_5288);
xnor U11462 (N_11462,N_5364,N_9275);
xor U11463 (N_11463,N_5441,N_6480);
and U11464 (N_11464,N_7407,N_5424);
xnor U11465 (N_11465,N_8590,N_6831);
or U11466 (N_11466,N_6524,N_7070);
xor U11467 (N_11467,N_9747,N_6371);
nor U11468 (N_11468,N_5872,N_8426);
nor U11469 (N_11469,N_9221,N_8216);
nor U11470 (N_11470,N_6463,N_5982);
and U11471 (N_11471,N_9645,N_8210);
nor U11472 (N_11472,N_6644,N_6446);
nor U11473 (N_11473,N_6101,N_6323);
nor U11474 (N_11474,N_9714,N_5212);
and U11475 (N_11475,N_8477,N_8558);
and U11476 (N_11476,N_7555,N_6813);
nor U11477 (N_11477,N_5082,N_6260);
or U11478 (N_11478,N_9093,N_5391);
nor U11479 (N_11479,N_5019,N_7102);
nand U11480 (N_11480,N_6002,N_5084);
or U11481 (N_11481,N_6812,N_8232);
nor U11482 (N_11482,N_6320,N_8017);
and U11483 (N_11483,N_7055,N_5839);
and U11484 (N_11484,N_6881,N_6720);
xnor U11485 (N_11485,N_9017,N_9943);
or U11486 (N_11486,N_5256,N_6042);
and U11487 (N_11487,N_9915,N_8340);
nand U11488 (N_11488,N_8472,N_6807);
or U11489 (N_11489,N_9163,N_8440);
nand U11490 (N_11490,N_9355,N_8838);
or U11491 (N_11491,N_8311,N_5742);
xor U11492 (N_11492,N_5975,N_6271);
xor U11493 (N_11493,N_6580,N_7163);
nor U11494 (N_11494,N_9644,N_9825);
nand U11495 (N_11495,N_8417,N_5500);
or U11496 (N_11496,N_6438,N_8992);
nand U11497 (N_11497,N_7082,N_8061);
or U11498 (N_11498,N_7655,N_5186);
or U11499 (N_11499,N_6368,N_7822);
nand U11500 (N_11500,N_8788,N_6569);
nor U11501 (N_11501,N_9233,N_8413);
or U11502 (N_11502,N_6772,N_8877);
xnor U11503 (N_11503,N_5442,N_8898);
or U11504 (N_11504,N_9097,N_6092);
and U11505 (N_11505,N_5905,N_6337);
xor U11506 (N_11506,N_6319,N_5733);
and U11507 (N_11507,N_8374,N_9411);
or U11508 (N_11508,N_9525,N_9556);
or U11509 (N_11509,N_9297,N_9467);
nor U11510 (N_11510,N_5785,N_5064);
xor U11511 (N_11511,N_5693,N_6538);
and U11512 (N_11512,N_7205,N_5715);
xor U11513 (N_11513,N_6139,N_7347);
or U11514 (N_11514,N_9117,N_7275);
and U11515 (N_11515,N_8567,N_8701);
nor U11516 (N_11516,N_9002,N_9162);
nand U11517 (N_11517,N_8241,N_9003);
and U11518 (N_11518,N_9528,N_9920);
xnor U11519 (N_11519,N_8087,N_5870);
and U11520 (N_11520,N_6858,N_6716);
xnor U11521 (N_11521,N_8841,N_8264);
and U11522 (N_11522,N_6146,N_9140);
xor U11523 (N_11523,N_7589,N_7777);
xnor U11524 (N_11524,N_7755,N_8922);
nor U11525 (N_11525,N_8471,N_5453);
or U11526 (N_11526,N_8751,N_5825);
nand U11527 (N_11527,N_8037,N_9211);
nor U11528 (N_11528,N_7935,N_9132);
or U11529 (N_11529,N_7596,N_8361);
and U11530 (N_11530,N_9913,N_6853);
nor U11531 (N_11531,N_5030,N_7968);
and U11532 (N_11532,N_7785,N_8079);
and U11533 (N_11533,N_7934,N_6951);
and U11534 (N_11534,N_8372,N_8080);
xnor U11535 (N_11535,N_5398,N_8884);
and U11536 (N_11536,N_8136,N_9692);
nor U11537 (N_11537,N_8375,N_7256);
nand U11538 (N_11538,N_5757,N_7360);
or U11539 (N_11539,N_8950,N_7928);
nand U11540 (N_11540,N_7658,N_8286);
and U11541 (N_11541,N_7383,N_7834);
xor U11542 (N_11542,N_6354,N_6964);
xor U11543 (N_11543,N_9321,N_7750);
nand U11544 (N_11544,N_8752,N_5059);
and U11545 (N_11545,N_8827,N_9277);
or U11546 (N_11546,N_9258,N_9646);
nor U11547 (N_11547,N_7956,N_8012);
xnor U11548 (N_11548,N_9847,N_8926);
xor U11549 (N_11549,N_6902,N_6934);
xnor U11550 (N_11550,N_7376,N_5403);
and U11551 (N_11551,N_8143,N_8427);
xor U11552 (N_11552,N_5820,N_8254);
and U11553 (N_11553,N_6913,N_5155);
or U11554 (N_11554,N_9120,N_8423);
nand U11555 (N_11555,N_6218,N_6922);
nand U11556 (N_11556,N_9273,N_5759);
nand U11557 (N_11557,N_6862,N_7230);
xor U11558 (N_11558,N_5372,N_8834);
and U11559 (N_11559,N_5269,N_8872);
xor U11560 (N_11560,N_8614,N_7233);
nand U11561 (N_11561,N_5278,N_6261);
nor U11562 (N_11562,N_7114,N_9940);
and U11563 (N_11563,N_9698,N_5548);
or U11564 (N_11564,N_8722,N_8209);
nand U11565 (N_11565,N_9030,N_9434);
nor U11566 (N_11566,N_8840,N_9768);
and U11567 (N_11567,N_6927,N_8876);
and U11568 (N_11568,N_6449,N_9959);
and U11569 (N_11569,N_8839,N_8158);
nor U11570 (N_11570,N_6238,N_7656);
or U11571 (N_11571,N_5840,N_6289);
or U11572 (N_11572,N_7508,N_9192);
nor U11573 (N_11573,N_7568,N_6584);
nand U11574 (N_11574,N_9633,N_6998);
nand U11575 (N_11575,N_5545,N_5365);
nand U11576 (N_11576,N_8260,N_9060);
xnor U11577 (N_11577,N_6305,N_5003);
nor U11578 (N_11578,N_8787,N_9413);
nand U11579 (N_11579,N_8112,N_9705);
and U11580 (N_11580,N_9092,N_7836);
nand U11581 (N_11581,N_9195,N_5527);
and U11582 (N_11582,N_6420,N_6281);
or U11583 (N_11583,N_5132,N_9833);
xnor U11584 (N_11584,N_8667,N_5623);
nor U11585 (N_11585,N_7948,N_5341);
xnor U11586 (N_11586,N_5609,N_9089);
nand U11587 (N_11587,N_9983,N_6282);
or U11588 (N_11588,N_6152,N_7209);
and U11589 (N_11589,N_9230,N_9846);
xnor U11590 (N_11590,N_6747,N_6954);
and U11591 (N_11591,N_8108,N_7669);
and U11592 (N_11592,N_9496,N_6283);
and U11593 (N_11593,N_7854,N_5760);
or U11594 (N_11594,N_6694,N_6552);
or U11595 (N_11595,N_6468,N_5606);
nand U11596 (N_11596,N_8771,N_7799);
nor U11597 (N_11597,N_7040,N_7660);
nor U11598 (N_11598,N_9359,N_8278);
and U11599 (N_11599,N_8332,N_8389);
nand U11600 (N_11600,N_7039,N_5752);
xnor U11601 (N_11601,N_6391,N_6498);
nor U11602 (N_11602,N_9680,N_7763);
xor U11603 (N_11603,N_7768,N_9797);
nand U11604 (N_11604,N_9865,N_8500);
nor U11605 (N_11605,N_5873,N_6683);
nand U11606 (N_11606,N_5353,N_9559);
nor U11607 (N_11607,N_9589,N_6658);
nor U11608 (N_11608,N_9672,N_5758);
nor U11609 (N_11609,N_5923,N_9399);
nand U11610 (N_11610,N_5011,N_8602);
nand U11611 (N_11611,N_5342,N_7362);
xnor U11612 (N_11612,N_9147,N_8414);
or U11613 (N_11613,N_9499,N_6750);
nor U11614 (N_11614,N_8496,N_7260);
xnor U11615 (N_11615,N_8021,N_9040);
or U11616 (N_11616,N_6942,N_7920);
or U11617 (N_11617,N_5918,N_6990);
or U11618 (N_11618,N_8704,N_7668);
or U11619 (N_11619,N_7961,N_5306);
nor U11620 (N_11620,N_6603,N_7503);
nand U11621 (N_11621,N_8626,N_5510);
xnor U11622 (N_11622,N_6104,N_5070);
nor U11623 (N_11623,N_7349,N_8010);
or U11624 (N_11624,N_5672,N_5886);
or U11625 (N_11625,N_9136,N_5521);
nand U11626 (N_11626,N_8443,N_6601);
or U11627 (N_11627,N_9824,N_7356);
or U11628 (N_11628,N_7904,N_8689);
nor U11629 (N_11629,N_7957,N_5889);
nor U11630 (N_11630,N_5736,N_6743);
and U11631 (N_11631,N_7297,N_6086);
nor U11632 (N_11632,N_5261,N_9807);
nor U11633 (N_11633,N_5057,N_8341);
nor U11634 (N_11634,N_7581,N_5792);
nor U11635 (N_11635,N_8125,N_9818);
nand U11636 (N_11636,N_9606,N_9884);
xor U11637 (N_11637,N_6794,N_9925);
or U11638 (N_11638,N_9058,N_8817);
and U11639 (N_11639,N_7214,N_7714);
and U11640 (N_11640,N_8699,N_7219);
and U11641 (N_11641,N_5142,N_9957);
and U11642 (N_11642,N_6182,N_5823);
xor U11643 (N_11643,N_9235,N_5912);
and U11644 (N_11644,N_6485,N_6530);
or U11645 (N_11645,N_6094,N_6234);
nand U11646 (N_11646,N_8895,N_6517);
or U11647 (N_11647,N_5270,N_8397);
nor U11648 (N_11648,N_7635,N_8086);
or U11649 (N_11649,N_8188,N_6873);
nand U11650 (N_11650,N_8124,N_6887);
xor U11651 (N_11651,N_7867,N_7577);
and U11652 (N_11652,N_7266,N_9812);
or U11653 (N_11653,N_7386,N_7473);
xnor U11654 (N_11654,N_5043,N_8761);
or U11655 (N_11655,N_8258,N_9335);
xnor U11656 (N_11656,N_6090,N_5328);
xnor U11657 (N_11657,N_5290,N_6349);
nor U11658 (N_11658,N_5450,N_8055);
nor U11659 (N_11659,N_9353,N_9811);
nor U11660 (N_11660,N_6762,N_7685);
and U11661 (N_11661,N_7379,N_7305);
or U11662 (N_11662,N_7381,N_6040);
xnor U11663 (N_11663,N_8754,N_5803);
xor U11664 (N_11664,N_6860,N_6872);
nor U11665 (N_11665,N_7437,N_8297);
nand U11666 (N_11666,N_7597,N_9686);
nand U11667 (N_11667,N_9182,N_6856);
and U11668 (N_11668,N_8539,N_6511);
xor U11669 (N_11669,N_9893,N_7762);
xor U11670 (N_11670,N_9305,N_9327);
nand U11671 (N_11671,N_9701,N_8425);
and U11672 (N_11672,N_7773,N_7633);
nand U11673 (N_11673,N_5957,N_6674);
nand U11674 (N_11674,N_5763,N_6274);
or U11675 (N_11675,N_8990,N_5634);
nand U11676 (N_11676,N_9006,N_8406);
xor U11677 (N_11677,N_5448,N_7071);
or U11678 (N_11678,N_7563,N_5272);
and U11679 (N_11679,N_9562,N_9620);
or U11680 (N_11680,N_6795,N_7203);
and U11681 (N_11681,N_9576,N_8179);
and U11682 (N_11682,N_7586,N_7030);
nor U11683 (N_11683,N_9174,N_5431);
xnor U11684 (N_11684,N_5138,N_5211);
nand U11685 (N_11685,N_5164,N_6421);
and U11686 (N_11686,N_5641,N_5647);
nor U11687 (N_11687,N_6829,N_9582);
or U11688 (N_11688,N_5325,N_6165);
and U11689 (N_11689,N_5526,N_5133);
or U11690 (N_11690,N_6633,N_9971);
and U11691 (N_11691,N_7487,N_6097);
xor U11692 (N_11692,N_7841,N_6120);
nand U11693 (N_11693,N_8583,N_7261);
nand U11694 (N_11694,N_9337,N_6550);
and U11695 (N_11695,N_9035,N_6520);
xnor U11696 (N_11696,N_5768,N_8481);
or U11697 (N_11697,N_7134,N_5412);
or U11698 (N_11698,N_9249,N_7686);
xor U11699 (N_11699,N_7747,N_6655);
or U11700 (N_11700,N_7380,N_7050);
nand U11701 (N_11701,N_9649,N_6864);
and U11702 (N_11702,N_8444,N_9455);
xnor U11703 (N_11703,N_7139,N_9049);
or U11704 (N_11704,N_6901,N_7591);
xor U11705 (N_11705,N_8463,N_7615);
and U11706 (N_11706,N_8142,N_5145);
or U11707 (N_11707,N_9947,N_5074);
nor U11708 (N_11708,N_6664,N_8016);
xnor U11709 (N_11709,N_9229,N_7521);
or U11710 (N_11710,N_9852,N_7447);
or U11711 (N_11711,N_6193,N_7479);
and U11712 (N_11712,N_8948,N_8746);
xor U11713 (N_11713,N_5590,N_9145);
nand U11714 (N_11714,N_5390,N_5338);
or U11715 (N_11715,N_6179,N_6593);
and U11716 (N_11716,N_5041,N_5395);
nand U11717 (N_11717,N_6099,N_5829);
xnor U11718 (N_11718,N_8535,N_9813);
nand U11719 (N_11719,N_6425,N_9789);
and U11720 (N_11720,N_9034,N_6095);
and U11721 (N_11721,N_6462,N_9191);
or U11722 (N_11722,N_7912,N_9510);
and U11723 (N_11723,N_7314,N_5331);
nor U11724 (N_11724,N_8806,N_5881);
nor U11725 (N_11725,N_6303,N_6815);
xor U11726 (N_11726,N_9520,N_5809);
xnor U11727 (N_11727,N_5476,N_8711);
nor U11728 (N_11728,N_6891,N_8601);
nand U11729 (N_11729,N_7781,N_6589);
xnor U11730 (N_11730,N_8742,N_8385);
xor U11731 (N_11731,N_5172,N_5407);
xor U11732 (N_11732,N_9165,N_9177);
or U11733 (N_11733,N_7110,N_9479);
or U11734 (N_11734,N_5067,N_5216);
xnor U11735 (N_11735,N_9604,N_7595);
or U11736 (N_11736,N_8267,N_6965);
and U11737 (N_11737,N_7420,N_5375);
xnor U11738 (N_11738,N_8346,N_7468);
or U11739 (N_11739,N_6174,N_8015);
nand U11740 (N_11740,N_8894,N_7868);
xnor U11741 (N_11741,N_9456,N_9101);
and U11742 (N_11742,N_8109,N_6208);
or U11743 (N_11743,N_8044,N_6911);
and U11744 (N_11744,N_8339,N_6754);
nor U11745 (N_11745,N_7535,N_8800);
nor U11746 (N_11746,N_9026,N_9081);
nor U11747 (N_11747,N_6059,N_7441);
nor U11748 (N_11748,N_9213,N_7289);
and U11749 (N_11749,N_8846,N_5974);
nand U11750 (N_11750,N_8072,N_7435);
nand U11751 (N_11751,N_8857,N_7525);
and U11752 (N_11752,N_5580,N_6356);
and U11753 (N_11753,N_6836,N_9535);
xnor U11754 (N_11754,N_7212,N_7509);
xor U11755 (N_11755,N_7752,N_9599);
xnor U11756 (N_11756,N_7224,N_6045);
or U11757 (N_11757,N_5629,N_8997);
nor U11758 (N_11758,N_5268,N_9027);
and U11759 (N_11759,N_5026,N_8094);
xnor U11760 (N_11760,N_6111,N_7276);
xnor U11761 (N_11761,N_6470,N_7171);
and U11762 (N_11762,N_6983,N_6222);
or U11763 (N_11763,N_6447,N_7720);
xor U11764 (N_11764,N_7988,N_7869);
and U11765 (N_11765,N_6960,N_5023);
xnor U11766 (N_11766,N_6564,N_9252);
or U11767 (N_11767,N_9518,N_7324);
xnor U11768 (N_11768,N_6242,N_9032);
or U11769 (N_11769,N_7817,N_8246);
xor U11770 (N_11770,N_9843,N_9678);
nand U11771 (N_11771,N_5275,N_7927);
nor U11772 (N_11772,N_8976,N_8393);
nor U11773 (N_11773,N_6643,N_7092);
and U11774 (N_11774,N_9673,N_8910);
and U11775 (N_11775,N_8245,N_5793);
or U11776 (N_11776,N_9020,N_9741);
and U11777 (N_11777,N_5640,N_5666);
nor U11778 (N_11778,N_9704,N_7132);
nor U11779 (N_11779,N_7054,N_6847);
or U11780 (N_11780,N_6048,N_6612);
nor U11781 (N_11781,N_9902,N_9860);
nor U11782 (N_11782,N_7611,N_5204);
xor U11783 (N_11783,N_9009,N_8592);
xnor U11784 (N_11784,N_5050,N_5680);
and U11785 (N_11785,N_6359,N_6495);
nor U11786 (N_11786,N_6268,N_8816);
and U11787 (N_11787,N_5153,N_5935);
or U11788 (N_11788,N_7318,N_8013);
nand U11789 (N_11789,N_9651,N_6642);
xor U11790 (N_11790,N_8544,N_7207);
or U11791 (N_11791,N_8524,N_8968);
nand U11792 (N_11792,N_5739,N_7552);
nand U11793 (N_11793,N_8591,N_8931);
nor U11794 (N_11794,N_6710,N_8333);
nor U11795 (N_11795,N_9450,N_8680);
nor U11796 (N_11796,N_5990,N_6617);
and U11797 (N_11797,N_7609,N_7675);
or U11798 (N_11798,N_6269,N_8892);
nor U11799 (N_11799,N_7169,N_6678);
nand U11800 (N_11800,N_8217,N_8502);
or U11801 (N_11801,N_6514,N_6783);
nor U11802 (N_11802,N_6475,N_6543);
and U11803 (N_11803,N_9363,N_5864);
xnor U11804 (N_11804,N_5808,N_9533);
xnor U11805 (N_11805,N_6316,N_6422);
or U11806 (N_11806,N_6916,N_6724);
xnor U11807 (N_11807,N_6357,N_6684);
and U11808 (N_11808,N_9596,N_7239);
xnor U11809 (N_11809,N_9200,N_9269);
or U11810 (N_11810,N_5080,N_8149);
and U11811 (N_11811,N_7145,N_5193);
nand U11812 (N_11812,N_6871,N_8206);
nor U11813 (N_11813,N_5576,N_8906);
nand U11814 (N_11814,N_9798,N_9457);
or U11815 (N_11815,N_8717,N_8523);
xnor U11816 (N_11816,N_9205,N_7394);
and U11817 (N_11817,N_7429,N_9095);
and U11818 (N_11818,N_7232,N_6237);
or U11819 (N_11819,N_5121,N_8560);
xnor U11820 (N_11820,N_6461,N_9642);
and U11821 (N_11821,N_7788,N_7766);
or U11822 (N_11822,N_8343,N_6168);
and U11823 (N_11823,N_8076,N_8599);
nand U11824 (N_11824,N_6614,N_9304);
xnor U11825 (N_11825,N_9772,N_7631);
nand U11826 (N_11826,N_9712,N_7023);
nand U11827 (N_11827,N_7514,N_6899);
and U11828 (N_11828,N_8486,N_6620);
nand U11829 (N_11829,N_6833,N_9251);
or U11830 (N_11830,N_6687,N_8000);
nor U11831 (N_11831,N_8129,N_7852);
nor U11832 (N_11832,N_8507,N_8762);
nor U11833 (N_11833,N_5639,N_5294);
nand U11834 (N_11834,N_5428,N_9503);
or U11835 (N_11835,N_5696,N_8479);
xnor U11836 (N_11836,N_5363,N_7981);
or U11837 (N_11837,N_7838,N_6454);
nor U11838 (N_11838,N_7831,N_9624);
and U11839 (N_11839,N_8322,N_6993);
nand U11840 (N_11840,N_5115,N_9949);
or U11841 (N_11841,N_5928,N_7361);
nand U11842 (N_11842,N_5126,N_8930);
or U11843 (N_11843,N_9356,N_9908);
nand U11844 (N_11844,N_9870,N_9099);
nor U11845 (N_11845,N_5284,N_5539);
xor U11846 (N_11846,N_9653,N_9351);
or U11847 (N_11847,N_8489,N_8091);
xnor U11848 (N_11848,N_5628,N_8969);
or U11849 (N_11849,N_7650,N_6149);
xnor U11850 (N_11850,N_5004,N_5368);
xnor U11851 (N_11851,N_8196,N_9816);
or U11852 (N_11852,N_8498,N_5048);
nor U11853 (N_11853,N_6959,N_9021);
nand U11854 (N_11854,N_6838,N_5425);
and U11855 (N_11855,N_8168,N_7178);
nand U11856 (N_11856,N_7455,N_8516);
xnor U11857 (N_11857,N_8706,N_6696);
nand U11858 (N_11858,N_5630,N_8300);
nand U11859 (N_11859,N_9755,N_8556);
xnor U11860 (N_11860,N_8007,N_9844);
or U11861 (N_11861,N_8419,N_7398);
xnor U11862 (N_11862,N_6851,N_5818);
nor U11863 (N_11863,N_6262,N_6979);
xor U11864 (N_11864,N_6705,N_7699);
and U11865 (N_11865,N_6457,N_8576);
and U11866 (N_11866,N_9280,N_7980);
xor U11867 (N_11867,N_7208,N_9326);
xor U11868 (N_11868,N_7887,N_6532);
and U11869 (N_11869,N_5844,N_5554);
and U11870 (N_11870,N_9064,N_7542);
xor U11871 (N_11871,N_7977,N_7264);
or U11872 (N_11872,N_5775,N_5058);
xor U11873 (N_11873,N_8445,N_9312);
xnor U11874 (N_11874,N_7789,N_7945);
xnor U11875 (N_11875,N_6657,N_9622);
and U11876 (N_11876,N_9598,N_6290);
or U11877 (N_11877,N_9008,N_9975);
xnor U11878 (N_11878,N_8458,N_7570);
or U11879 (N_11879,N_7857,N_5117);
and U11880 (N_11880,N_5486,N_6918);
or U11881 (N_11881,N_8053,N_8545);
or U11882 (N_11882,N_7677,N_6064);
nand U11883 (N_11883,N_5555,N_5104);
or U11884 (N_11884,N_7488,N_9806);
nand U11885 (N_11885,N_5243,N_6239);
xor U11886 (N_11886,N_8280,N_8088);
nor U11887 (N_11887,N_7446,N_9608);
or U11888 (N_11888,N_7991,N_6625);
and U11889 (N_11889,N_8011,N_5610);
nor U11890 (N_11890,N_5008,N_7894);
nor U11891 (N_11891,N_6372,N_7007);
xnor U11892 (N_11892,N_5891,N_6458);
and U11893 (N_11893,N_7452,N_5238);
nor U11894 (N_11894,N_8229,N_7549);
xnor U11895 (N_11895,N_9905,N_6373);
nand U11896 (N_11896,N_9817,N_9759);
nor U11897 (N_11897,N_8874,N_7148);
xor U11898 (N_11898,N_7953,N_7666);
and U11899 (N_11899,N_5782,N_6540);
nor U11900 (N_11900,N_7001,N_9242);
nor U11901 (N_11901,N_7874,N_9896);
nand U11902 (N_11902,N_7738,N_8266);
and U11903 (N_11903,N_5893,N_6053);
and U11904 (N_11904,N_8235,N_8975);
and U11905 (N_11905,N_8453,N_7471);
nand U11906 (N_11906,N_8455,N_8510);
xor U11907 (N_11907,N_9458,N_8161);
and U11908 (N_11908,N_8219,N_5940);
nor U11909 (N_11909,N_5636,N_6116);
nand U11910 (N_11910,N_6556,N_6161);
or U11911 (N_11911,N_7354,N_5273);
and U11912 (N_11912,N_8358,N_5430);
and U11913 (N_11913,N_7757,N_8668);
xor U11914 (N_11914,N_6719,N_9042);
nor U11915 (N_11915,N_9618,N_8675);
nand U11916 (N_11916,N_7321,N_5170);
or U11917 (N_11917,N_6561,N_5347);
nand U11918 (N_11918,N_6755,N_7199);
nor U11919 (N_11919,N_9131,N_5776);
or U11920 (N_11920,N_5493,N_6600);
or U11921 (N_11921,N_8822,N_5443);
and U11922 (N_11922,N_5362,N_6852);
nor U11923 (N_11923,N_9694,N_8977);
or U11924 (N_11924,N_7428,N_9303);
nand U11925 (N_11925,N_6183,N_8662);
or U11926 (N_11926,N_6075,N_8663);
nand U11927 (N_11927,N_5236,N_7897);
and U11928 (N_11928,N_6401,N_7536);
or U11929 (N_11929,N_6073,N_6839);
xnor U11930 (N_11930,N_7944,N_9962);
nor U11931 (N_11931,N_8595,N_5675);
nand U11932 (N_11932,N_5397,N_6753);
nand U11933 (N_11933,N_7682,N_8833);
nand U11934 (N_11934,N_9086,N_7244);
or U11935 (N_11935,N_9990,N_5701);
nor U11936 (N_11936,N_5997,N_5152);
nor U11937 (N_11937,N_8348,N_6787);
or U11938 (N_11938,N_5129,N_5076);
nand U11939 (N_11939,N_6732,N_8756);
and U11940 (N_11940,N_7637,N_5396);
nand U11941 (N_11941,N_8605,N_8832);
xor U11942 (N_11942,N_8794,N_7805);
and U11943 (N_11943,N_7813,N_9763);
and U11944 (N_11944,N_5339,N_6840);
nor U11945 (N_11945,N_9107,N_5949);
or U11946 (N_11946,N_8320,N_8329);
or U11947 (N_11947,N_9721,N_9354);
xor U11948 (N_11948,N_8362,N_6955);
and U11949 (N_11949,N_7846,N_8218);
and U11950 (N_11950,N_7771,N_8313);
nand U11951 (N_11951,N_9422,N_5333);
nand U11952 (N_11952,N_7093,N_9106);
or U11953 (N_11953,N_9239,N_6752);
nand U11954 (N_11954,N_6745,N_8213);
and U11955 (N_11955,N_9336,N_6402);
or U11956 (N_11956,N_5485,N_6383);
nor U11957 (N_11957,N_9114,N_9142);
xnor U11958 (N_11958,N_6929,N_9210);
or U11959 (N_11959,N_8738,N_6325);
xnor U11960 (N_11960,N_9688,N_5156);
and U11961 (N_11961,N_6680,N_6895);
nor U11962 (N_11962,N_7303,N_5897);
xnor U11963 (N_11963,N_5632,N_8650);
nor U11964 (N_11964,N_7598,N_8342);
nor U11965 (N_11965,N_6616,N_9066);
or U11966 (N_11966,N_7523,N_7466);
nor U11967 (N_11967,N_5125,N_6312);
and U11968 (N_11968,N_8912,N_8928);
or U11969 (N_11969,N_9246,N_6352);
or U11970 (N_11970,N_8132,N_8367);
xnor U11971 (N_11971,N_7796,N_7313);
nor U11972 (N_11972,N_6286,N_7445);
or U11973 (N_11973,N_8429,N_6654);
nor U11974 (N_11974,N_7998,N_7333);
or U11975 (N_11975,N_7097,N_9207);
nand U11976 (N_11976,N_8293,N_6950);
xnor U11977 (N_11977,N_9133,N_7310);
and U11978 (N_11978,N_9731,N_7603);
xor U11979 (N_11979,N_5649,N_7052);
nor U11980 (N_11980,N_8559,N_8049);
nand U11981 (N_11981,N_5162,N_6178);
or U11982 (N_11982,N_8172,N_6761);
xnor U11983 (N_11983,N_8561,N_7194);
nor U11984 (N_11984,N_8494,N_6568);
and U11985 (N_11985,N_7942,N_7127);
nand U11986 (N_11986,N_8563,N_8315);
xor U11987 (N_11987,N_7886,N_9883);
nand U11988 (N_11988,N_5951,N_7281);
or U11989 (N_11989,N_9076,N_8005);
nand U11990 (N_11990,N_7827,N_9919);
nand U11991 (N_11991,N_5491,N_6245);
nor U11992 (N_11992,N_6878,N_9805);
nor U11993 (N_11993,N_8435,N_5756);
nor U11994 (N_11994,N_9333,N_8040);
nand U11995 (N_11995,N_8873,N_5228);
nor U11996 (N_11996,N_7737,N_6173);
nor U11997 (N_11997,N_6023,N_9361);
or U11998 (N_11998,N_8790,N_7931);
nand U11999 (N_11999,N_6285,N_8654);
or U12000 (N_12000,N_9267,N_6541);
or U12001 (N_12001,N_9577,N_8953);
and U12002 (N_12002,N_9255,N_6555);
or U12003 (N_12003,N_9570,N_9167);
or U12004 (N_12004,N_7459,N_6968);
nand U12005 (N_12005,N_7344,N_9640);
and U12006 (N_12006,N_5869,N_5359);
and U12007 (N_12007,N_5489,N_8381);
xor U12008 (N_12008,N_9561,N_8685);
nor U12009 (N_12009,N_9109,N_9301);
nand U12010 (N_12010,N_6311,N_7217);
nand U12011 (N_12011,N_8686,N_6196);
and U12012 (N_12012,N_7448,N_7608);
xnor U12013 (N_12013,N_6405,N_8099);
and U12014 (N_12014,N_5814,N_5356);
nand U12015 (N_12015,N_8891,N_5853);
nand U12016 (N_12016,N_6526,N_9924);
xnor U12017 (N_12017,N_7532,N_8681);
xnor U12018 (N_12018,N_5045,N_7457);
xnor U12019 (N_12019,N_6386,N_8083);
or U12020 (N_12020,N_8431,N_6567);
xor U12021 (N_12021,N_7022,N_7543);
xnor U12022 (N_12022,N_8378,N_5600);
nor U12023 (N_12023,N_9045,N_8844);
xnor U12024 (N_12024,N_8697,N_8030);
or U12025 (N_12025,N_6130,N_9431);
nor U12026 (N_12026,N_9248,N_9179);
or U12027 (N_12027,N_6070,N_8837);
or U12028 (N_12028,N_5024,N_8712);
and U12029 (N_12029,N_5766,N_9172);
nand U12030 (N_12030,N_7108,N_9154);
nor U12031 (N_12031,N_5706,N_8995);
xnor U12032 (N_12032,N_6304,N_6263);
nor U12033 (N_12033,N_7636,N_7530);
nor U12034 (N_12034,N_9471,N_6296);
and U12035 (N_12035,N_9314,N_9151);
nor U12036 (N_12036,N_5856,N_6393);
or U12037 (N_12037,N_8944,N_5394);
and U12038 (N_12038,N_9995,N_5831);
xor U12039 (N_12039,N_8089,N_5227);
nor U12040 (N_12040,N_6247,N_5092);
xnor U12041 (N_12041,N_5166,N_7765);
nand U12042 (N_12042,N_7021,N_8747);
and U12043 (N_12043,N_5239,N_5106);
xnor U12044 (N_12044,N_8870,N_6211);
nor U12045 (N_12045,N_6013,N_8671);
or U12046 (N_12046,N_9122,N_8190);
or U12047 (N_12047,N_7847,N_7120);
and U12048 (N_12048,N_9887,N_9899);
or U12049 (N_12049,N_5849,N_7794);
nand U12050 (N_12050,N_8066,N_7278);
and U12051 (N_12051,N_6888,N_6562);
and U12052 (N_12052,N_6144,N_5558);
and U12053 (N_12053,N_5977,N_9484);
nand U12054 (N_12054,N_7626,N_7732);
xnor U12055 (N_12055,N_7323,N_8571);
or U12056 (N_12056,N_7667,N_8845);
or U12057 (N_12057,N_7128,N_5361);
nand U12058 (N_12058,N_5621,N_9443);
nand U12059 (N_12059,N_7342,N_9760);
nand U12060 (N_12060,N_9331,N_8745);
nand U12061 (N_12061,N_5210,N_5355);
or U12062 (N_12062,N_5446,N_5298);
and U12063 (N_12063,N_6272,N_9521);
or U12064 (N_12064,N_8309,N_8627);
or U12065 (N_12065,N_9061,N_5655);
or U12066 (N_12066,N_9963,N_6254);
and U12067 (N_12067,N_8391,N_7076);
xor U12068 (N_12068,N_9317,N_9587);
and U12069 (N_12069,N_5673,N_9268);
nor U12070 (N_12070,N_9051,N_8350);
and U12071 (N_12071,N_6184,N_6792);
nand U12072 (N_12072,N_7113,N_7866);
and U12073 (N_12073,N_9028,N_8051);
and U12074 (N_12074,N_9368,N_7971);
xor U12075 (N_12075,N_6404,N_9808);
xnor U12076 (N_12076,N_7014,N_5000);
nand U12077 (N_12077,N_5089,N_8528);
nor U12078 (N_12078,N_5503,N_7913);
xnor U12079 (N_12079,N_6939,N_5884);
and U12080 (N_12080,N_8700,N_9068);
or U12081 (N_12081,N_6578,N_5399);
xor U12082 (N_12082,N_7421,N_8157);
xnor U12083 (N_12083,N_9270,N_6306);
or U12084 (N_12084,N_8047,N_8279);
nor U12085 (N_12085,N_8514,N_7282);
xnor U12086 (N_12086,N_5619,N_6841);
nor U12087 (N_12087,N_6232,N_9862);
xnor U12088 (N_12088,N_5468,N_6082);
nor U12089 (N_12089,N_8904,N_8587);
and U12090 (N_12090,N_7234,N_9679);
nand U12091 (N_12091,N_5999,N_8060);
xor U12092 (N_12092,N_8613,N_8688);
xor U12093 (N_12093,N_8068,N_5223);
and U12094 (N_12094,N_6302,N_8607);
or U12095 (N_12095,N_5250,N_5199);
nand U12096 (N_12096,N_9175,N_9105);
and U12097 (N_12097,N_6340,N_8456);
and U12098 (N_12098,N_7064,N_9944);
and U12099 (N_12099,N_7147,N_9296);
nand U12100 (N_12100,N_8470,N_9722);
xor U12101 (N_12101,N_5702,N_5081);
xor U12102 (N_12102,N_8111,N_7556);
or U12103 (N_12103,N_7016,N_5573);
and U12104 (N_12104,N_6828,N_8755);
or U12105 (N_12105,N_5033,N_6230);
or U12106 (N_12106,N_8420,N_9542);
xor U12107 (N_12107,N_6826,N_7351);
xor U12108 (N_12108,N_8959,N_5283);
and U12109 (N_12109,N_6585,N_5535);
and U12110 (N_12110,N_9157,N_5466);
xnor U12111 (N_12111,N_7450,N_9398);
or U12112 (N_12112,N_8226,N_8637);
nor U12113 (N_12113,N_5176,N_9062);
and U12114 (N_12114,N_7150,N_6227);
or U12115 (N_12115,N_6114,N_6361);
nor U12116 (N_12116,N_9016,N_6471);
nor U12117 (N_12117,N_6749,N_7946);
or U12118 (N_12118,N_7353,N_5091);
nand U12119 (N_12119,N_7604,N_6822);
xor U12120 (N_12120,N_5611,N_5163);
or U12121 (N_12121,N_5532,N_7775);
or U12122 (N_12122,N_6648,N_9495);
and U12123 (N_12123,N_8897,N_6465);
or U12124 (N_12124,N_9921,N_7518);
xnor U12125 (N_12125,N_7195,N_8281);
and U12126 (N_12126,N_5620,N_8386);
or U12127 (N_12127,N_5195,N_6240);
and U12128 (N_12128,N_9197,N_9433);
or U12129 (N_12129,N_8133,N_7839);
nor U12130 (N_12130,N_8843,N_9390);
nand U12131 (N_12131,N_6799,N_6024);
or U12132 (N_12132,N_9637,N_6112);
nand U12133 (N_12133,N_6430,N_8653);
nor U12134 (N_12134,N_8071,N_5107);
nand U12135 (N_12135,N_6191,N_7985);
and U12136 (N_12136,N_6406,N_8888);
nand U12137 (N_12137,N_6656,N_5422);
and U12138 (N_12138,N_8785,N_9890);
and U12139 (N_12139,N_6986,N_5404);
xnor U12140 (N_12140,N_5852,N_8574);
or U12141 (N_12141,N_9601,N_5332);
or U12142 (N_12142,N_5149,N_5102);
xor U12143 (N_12143,N_7539,N_8501);
and U12144 (N_12144,N_7787,N_7705);
xnor U12145 (N_12145,N_6248,N_7772);
xnor U12146 (N_12146,N_5329,N_5440);
nand U12147 (N_12147,N_5167,N_6088);
xnor U12148 (N_12148,N_5561,N_8634);
xor U12149 (N_12149,N_9676,N_8251);
xnor U12150 (N_12150,N_7146,N_5837);
nor U12151 (N_12151,N_6994,N_6057);
and U12152 (N_12152,N_8784,N_7179);
and U12153 (N_12153,N_9753,N_6252);
and U12154 (N_12154,N_5572,N_7427);
nand U12155 (N_12155,N_5213,N_8966);
nor U12156 (N_12156,N_5583,N_9869);
or U12157 (N_12157,N_7979,N_6201);
or U12158 (N_12158,N_6861,N_6582);
or U12159 (N_12159,N_5528,N_5456);
and U12160 (N_12160,N_6802,N_6781);
xnor U12161 (N_12161,N_7339,N_5479);
nand U12162 (N_12162,N_5480,N_8488);
or U12163 (N_12163,N_5737,N_7400);
or U12164 (N_12164,N_8879,N_5838);
nor U12165 (N_12165,N_9491,N_8274);
or U12166 (N_12166,N_6560,N_6592);
and U12167 (N_12167,N_9203,N_8538);
or U12168 (N_12168,N_6069,N_7616);
nor U12169 (N_12169,N_8231,N_8159);
nand U12170 (N_12170,N_9710,N_5734);
and U12171 (N_12171,N_9513,N_7103);
nand U12172 (N_12172,N_5018,N_5086);
xor U12173 (N_12173,N_6995,N_5435);
nand U12174 (N_12174,N_8676,N_5063);
nand U12175 (N_12175,N_7567,N_7572);
xnor U12176 (N_12176,N_6588,N_8039);
or U12177 (N_12177,N_6326,N_8098);
nor U12178 (N_12178,N_8008,N_6627);
or U12179 (N_12179,N_9024,N_5277);
or U12180 (N_12180,N_7559,N_7856);
nor U12181 (N_12181,N_9820,N_5247);
nand U12182 (N_12182,N_6830,N_6259);
nand U12183 (N_12183,N_9999,N_7149);
nor U12184 (N_12184,N_5027,N_8519);
nand U12185 (N_12185,N_6975,N_9469);
or U12186 (N_12186,N_8379,N_7717);
and U12187 (N_12187,N_5367,N_9453);
nor U12188 (N_12188,N_8956,N_7917);
nand U12189 (N_12189,N_8416,N_8369);
or U12190 (N_12190,N_6527,N_5157);
nand U12191 (N_12191,N_7290,N_5909);
nor U12192 (N_12192,N_6652,N_9000);
nor U12193 (N_12193,N_8802,N_7938);
xnor U12194 (N_12194,N_9480,N_9516);
nand U12195 (N_12195,N_8774,N_8570);
nor U12196 (N_12196,N_8195,N_5914);
and U12197 (N_12197,N_5455,N_9010);
and U12198 (N_12198,N_7793,N_6624);
nand U12199 (N_12199,N_6808,N_6496);
xnor U12200 (N_12200,N_7161,N_8710);
xor U12201 (N_12201,N_5743,N_9039);
nor U12202 (N_12202,N_9738,N_8271);
nor U12203 (N_12203,N_5090,N_6722);
nand U12204 (N_12204,N_5178,N_5101);
and U12205 (N_12205,N_9153,N_6397);
xor U12206 (N_12206,N_9512,N_7895);
nor U12207 (N_12207,N_5650,N_5305);
xnor U12208 (N_12208,N_9291,N_8162);
and U12209 (N_12209,N_5550,N_7879);
or U12210 (N_12210,N_5229,N_5547);
nand U12211 (N_12211,N_8244,N_6611);
and U12212 (N_12212,N_7818,N_6647);
and U12213 (N_12213,N_9419,N_5865);
nor U12214 (N_12214,N_9126,N_7830);
nor U12215 (N_12215,N_5475,N_5542);
xnor U12216 (N_12216,N_6884,N_7882);
and U12217 (N_12217,N_6441,N_5589);
nand U12218 (N_12218,N_7484,N_7402);
nand U12219 (N_12219,N_7495,N_9972);
xor U12220 (N_12220,N_6321,N_6154);
nor U12221 (N_12221,N_5146,N_6728);
nor U12222 (N_12222,N_6972,N_5179);
xor U12223 (N_12223,N_7599,N_7748);
and U12224 (N_12224,N_8137,N_6074);
or U12225 (N_12225,N_5301,N_8914);
nand U12226 (N_12226,N_8029,N_5520);
xor U12227 (N_12227,N_5727,N_8577);
nor U12228 (N_12228,N_6782,N_7385);
nand U12229 (N_12229,N_6223,N_8466);
or U12230 (N_12230,N_9850,N_9904);
nand U12231 (N_12231,N_8555,N_5599);
or U12232 (N_12232,N_9629,N_9046);
nor U12233 (N_12233,N_7433,N_7301);
xnor U12234 (N_12234,N_8027,N_6788);
nand U12235 (N_12235,N_8795,N_9223);
nor U12236 (N_12236,N_7691,N_6399);
and U12237 (N_12237,N_5462,N_9891);
nor U12238 (N_12238,N_7175,N_7031);
or U12239 (N_12239,N_7742,N_5801);
nor U12240 (N_12240,N_5671,N_7359);
and U12241 (N_12241,N_7470,N_7141);
or U12242 (N_12242,N_7708,N_6253);
and U12243 (N_12243,N_8548,N_8957);
and U12244 (N_12244,N_7995,N_9732);
nand U12245 (N_12245,N_5281,N_7562);
or U12246 (N_12246,N_9123,N_9074);
or U12247 (N_12247,N_9425,N_9379);
nand U12248 (N_12248,N_9482,N_8331);
and U12249 (N_12249,N_8185,N_5973);
nor U12250 (N_12250,N_9974,N_5563);
nand U12251 (N_12251,N_9440,N_7760);
xor U12252 (N_12252,N_9048,N_7634);
nand U12253 (N_12253,N_9143,N_7629);
nand U12254 (N_12254,N_5112,N_5130);
nand U12255 (N_12255,N_9631,N_8731);
nand U12256 (N_12256,N_9396,N_5192);
and U12257 (N_12257,N_8589,N_5242);
nand U12258 (N_12258,N_8383,N_9160);
xnor U12259 (N_12259,N_8221,N_9835);
nand U12260 (N_12260,N_9540,N_6037);
or U12261 (N_12261,N_8439,N_5326);
nor U12262 (N_12262,N_6790,N_9241);
nor U12263 (N_12263,N_8714,N_8713);
nand U12264 (N_12264,N_6594,N_9700);
or U12265 (N_12265,N_8967,N_6711);
or U12266 (N_12266,N_6443,N_7155);
nor U12267 (N_12267,N_8181,N_6121);
nor U12268 (N_12268,N_9595,N_7089);
nand U12269 (N_12269,N_7588,N_9571);
nor U12270 (N_12270,N_6599,N_5568);
or U12271 (N_12271,N_6063,N_5481);
nand U12272 (N_12272,N_8057,N_7258);
nand U12273 (N_12273,N_5415,N_7405);
xor U12274 (N_12274,N_9472,N_6145);
xnor U12275 (N_12275,N_5688,N_9238);
xnor U12276 (N_12276,N_8673,N_7432);
and U12277 (N_12277,N_8257,N_9867);
nor U12278 (N_12278,N_9591,N_7999);
nor U12279 (N_12279,N_6414,N_9945);
and U12280 (N_12280,N_8964,N_8180);
nor U12281 (N_12281,N_9150,N_8826);
and U12282 (N_12282,N_8204,N_5682);
nand U12283 (N_12283,N_9366,N_6046);
xor U12284 (N_12284,N_5774,N_7037);
or U12285 (N_12285,N_8430,N_7271);
nor U12286 (N_12286,N_6459,N_6797);
nor U12287 (N_12287,N_7334,N_9103);
nand U12288 (N_12288,N_5827,N_9240);
nand U12289 (N_12289,N_7255,N_8103);
or U12290 (N_12290,N_9183,N_5993);
nand U12291 (N_12291,N_8781,N_5463);
or U12292 (N_12292,N_8298,N_9362);
xnor U12293 (N_12293,N_5654,N_8695);
and U12294 (N_12294,N_7415,N_6632);
nand U12295 (N_12295,N_8763,N_6882);
xnor U12296 (N_12296,N_6940,N_8777);
or U12297 (N_12297,N_8693,N_9428);
xor U12298 (N_12298,N_5915,N_6697);
nand U12299 (N_12299,N_8719,N_8438);
nor U12300 (N_12300,N_7683,N_5406);
and U12301 (N_12301,N_9186,N_8789);
or U12302 (N_12302,N_5638,N_5678);
xor U12303 (N_12303,N_7676,N_8672);
nand U12304 (N_12304,N_7923,N_7104);
or U12305 (N_12305,N_5815,N_7012);
xnor U12306 (N_12306,N_5349,N_5877);
xnor U12307 (N_12307,N_9386,N_8234);
nand U12308 (N_12308,N_5330,N_8187);
or U12309 (N_12309,N_5716,N_7949);
nand U12310 (N_12310,N_5900,N_7136);
nor U12311 (N_12311,N_9261,N_6736);
and U12312 (N_12312,N_8046,N_6066);
xnor U12313 (N_12313,N_9374,N_6944);
nor U12314 (N_12314,N_8909,N_6742);
nor U12315 (N_12315,N_5690,N_6335);
nor U12316 (N_12316,N_8412,N_6672);
xnor U12317 (N_12317,N_7564,N_7236);
or U12318 (N_12318,N_8531,N_9764);
and U12319 (N_12319,N_8335,N_6176);
nor U12320 (N_12320,N_7835,N_7613);
nand U12321 (N_12321,N_6798,N_8760);
and U12322 (N_12322,N_9881,N_9677);
or U12323 (N_12323,N_8126,N_9751);
or U12324 (N_12324,N_9421,N_9256);
nor U12325 (N_12325,N_5725,N_5755);
nor U12326 (N_12326,N_6522,N_6903);
and U12327 (N_12327,N_8864,N_6776);
and U12328 (N_12328,N_5379,N_9276);
nor U12329 (N_12329,N_8323,N_9234);
nand U12330 (N_12330,N_9888,N_5944);
nand U12331 (N_12331,N_7606,N_8911);
or U12332 (N_12332,N_7654,N_9500);
or U12333 (N_12333,N_6646,N_5054);
and U12334 (N_12334,N_7198,N_6387);
and U12335 (N_12335,N_8615,N_5790);
xnor U12336 (N_12336,N_8943,N_9033);
and U12337 (N_12337,N_8002,N_7272);
nand U12338 (N_12338,N_9799,N_7735);
nand U12339 (N_12339,N_8307,N_6715);
xnor U12340 (N_12340,N_6481,N_8450);
nor U12341 (N_12341,N_6314,N_7739);
xnor U12342 (N_12342,N_5388,N_5053);
or U12343 (N_12343,N_8038,N_7489);
nor U12344 (N_12344,N_9873,N_5699);
and U12345 (N_12345,N_7884,N_8521);
nor U12346 (N_12346,N_5032,N_8220);
xnor U12347 (N_12347,N_8122,N_8553);
and U12348 (N_12348,N_8006,N_7162);
or U12349 (N_12349,N_6212,N_5518);
and U12350 (N_12350,N_7833,N_8102);
or U12351 (N_12351,N_8330,N_8509);
xor U12352 (N_12352,N_7687,N_7557);
or U12353 (N_12353,N_7545,N_8407);
and U12354 (N_12354,N_8054,N_8631);
xnor U12355 (N_12355,N_9271,N_8586);
nand U12356 (N_12356,N_8955,N_8184);
and U12357 (N_12357,N_8337,N_9634);
or U12358 (N_12358,N_9828,N_9407);
nor U12359 (N_12359,N_6390,N_6363);
or U12360 (N_12360,N_5913,N_7440);
and U12361 (N_12361,N_8314,N_8987);
nand U12362 (N_12362,N_9711,N_7807);
nand U12363 (N_12363,N_5802,N_5591);
and U12364 (N_12364,N_7736,N_7801);
nand U12365 (N_12365,N_7188,N_6946);
or U12366 (N_12366,N_9933,N_9841);
or U12367 (N_12367,N_6118,N_9488);
xnor U12368 (N_12368,N_7820,N_6117);
nor U12369 (N_12369,N_8513,N_5919);
and U12370 (N_12370,N_9541,N_6764);
or U12371 (N_12371,N_6622,N_8388);
nor U12372 (N_12372,N_8366,N_5198);
and U12373 (N_12373,N_5751,N_7293);
and U12374 (N_12374,N_6688,N_6439);
nor U12375 (N_12375,N_6389,N_8718);
nand U12376 (N_12376,N_7156,N_7812);
and U12377 (N_12377,N_7187,N_7392);
nor U12378 (N_12378,N_9802,N_8905);
or U12379 (N_12379,N_9667,N_8384);
and U12380 (N_12380,N_6014,N_9310);
and U12381 (N_12381,N_5501,N_7951);
and U12382 (N_12382,N_8941,N_9260);
and U12383 (N_12383,N_7182,N_8033);
and U12384 (N_12384,N_5358,N_6427);
nor U12385 (N_12385,N_8866,N_8308);
xor U12386 (N_12386,N_9660,N_9783);
and U12387 (N_12387,N_9923,N_6712);
or U12388 (N_12388,N_8951,N_8116);
or U12389 (N_12389,N_9659,N_5750);
xnor U12390 (N_12390,N_6124,N_8031);
or U12391 (N_12391,N_5712,N_8856);
xnor U12392 (N_12392,N_8113,N_5559);
nand U12393 (N_12393,N_6010,N_5495);
nand U12394 (N_12394,N_6607,N_5544);
xnor U12395 (N_12395,N_6291,N_8934);
xnor U12396 (N_12396,N_9011,N_6516);
xnor U12397 (N_12397,N_6229,N_5963);
and U12398 (N_12398,N_5783,N_5631);
nand U12399 (N_12399,N_8623,N_7074);
nor U12400 (N_12400,N_6668,N_8155);
nand U12401 (N_12401,N_8594,N_9859);
nand U12402 (N_12402,N_7201,N_8482);
or U12403 (N_12403,N_9169,N_7393);
or U12404 (N_12404,N_8338,N_7744);
nand U12405 (N_12405,N_9578,N_5866);
and U12406 (N_12406,N_5593,N_5608);
nor U12407 (N_12407,N_8084,N_8981);
nand U12408 (N_12408,N_6504,N_7107);
nor U12409 (N_12409,N_5037,N_7753);
xor U12410 (N_12410,N_7366,N_9973);
and U12411 (N_12411,N_8349,N_9091);
nand U12412 (N_12412,N_9292,N_7267);
nand U12413 (N_12413,N_7263,N_9566);
nand U12414 (N_12414,N_9786,N_9810);
or U12415 (N_12415,N_7168,N_5574);
or U12416 (N_12416,N_6874,N_5959);
or U12417 (N_12417,N_9382,N_9614);
and U12418 (N_12418,N_7262,N_6570);
xnor U12419 (N_12419,N_7573,N_8815);
nor U12420 (N_12420,N_8065,N_5304);
xor U12421 (N_12421,N_7966,N_9295);
nand U12422 (N_12422,N_6072,N_9170);
or U12423 (N_12423,N_5799,N_7358);
nor U12424 (N_12424,N_6508,N_5868);
nand U12425 (N_12425,N_9524,N_9418);
xnor U12426 (N_12426,N_7028,N_6774);
xnor U12427 (N_12427,N_7245,N_8736);
xor U12428 (N_12428,N_5218,N_6910);
or U12429 (N_12429,N_9096,N_5426);
xor U12430 (N_12430,N_8642,N_5968);
nand U12431 (N_12431,N_6054,N_7340);
and U12432 (N_12432,N_9005,N_5784);
or U12433 (N_12433,N_8303,N_6848);
or U12434 (N_12434,N_6293,N_6989);
or U12435 (N_12435,N_9220,N_9018);
xnor U12436 (N_12436,N_9391,N_8940);
and U12437 (N_12437,N_7756,N_5282);
or U12438 (N_12438,N_6921,N_7512);
nand U12439 (N_12439,N_7672,N_5635);
or U12440 (N_12440,N_5177,N_7119);
or U12441 (N_12441,N_9565,N_7865);
nor U12442 (N_12442,N_7704,N_5265);
nor U12443 (N_12443,N_8353,N_5423);
nor U12444 (N_12444,N_8199,N_9669);
nand U12445 (N_12445,N_6558,N_6803);
nand U12446 (N_12446,N_9128,N_7311);
xnor U12447 (N_12447,N_6017,N_7226);
nand U12448 (N_12448,N_6832,N_7517);
or U12449 (N_12449,N_6221,N_5669);
nand U12450 (N_12450,N_9750,N_5180);
nand U12451 (N_12451,N_8110,N_5596);
and U12452 (N_12452,N_9842,N_6077);
and U12453 (N_12453,N_5781,N_5899);
nor U12454 (N_12454,N_8557,N_6695);
nand U12455 (N_12455,N_6855,N_9057);
nand U12456 (N_12456,N_8621,N_6452);
nand U12457 (N_12457,N_9635,N_6931);
nor U12458 (N_12458,N_9158,N_6996);
xnor U12459 (N_12459,N_9129,N_9788);
and U12460 (N_12460,N_5777,N_8796);
nor U12461 (N_12461,N_9761,N_8579);
nor U12462 (N_12462,N_9263,N_8853);
nand U12463 (N_12463,N_5724,N_5607);
xnor U12464 (N_12464,N_8382,N_7526);
xnor U12465 (N_12465,N_8050,N_9953);
nor U12466 (N_12466,N_6673,N_8454);
xor U12467 (N_12467,N_5005,N_8851);
or U12468 (N_12468,N_6662,N_9052);
xnor U12469 (N_12469,N_9767,N_9085);
and U12470 (N_12470,N_9130,N_6915);
or U12471 (N_12471,N_7157,N_9581);
nor U12472 (N_12472,N_7955,N_9950);
or U12473 (N_12473,N_7143,N_7480);
or U12474 (N_12474,N_5920,N_8929);
or U12475 (N_12475,N_5767,N_5320);
nor U12476 (N_12476,N_7790,N_5557);
and U12477 (N_12477,N_7458,N_9942);
nand U12478 (N_12478,N_5861,N_7130);
nand U12479 (N_12479,N_5337,N_5136);
xor U12480 (N_12480,N_9498,N_8073);
nor U12481 (N_12481,N_6685,N_8294);
nand U12482 (N_12482,N_5553,N_8192);
or U12483 (N_12483,N_8913,N_9334);
or U12484 (N_12484,N_5189,N_7972);
nor U12485 (N_12485,N_6809,N_7077);
and U12486 (N_12486,N_9173,N_8945);
xor U12487 (N_12487,N_5879,N_8428);
xor U12488 (N_12488,N_8140,N_8584);
nor U12489 (N_12489,N_9969,N_8139);
nor U12490 (N_12490,N_5071,N_5025);
nand U12491 (N_12491,N_7370,N_7249);
or U12492 (N_12492,N_6136,N_5436);
nor U12493 (N_12493,N_8090,N_8797);
and U12494 (N_12494,N_8208,N_7124);
or U12495 (N_12495,N_8077,N_8128);
nor U12496 (N_12496,N_5310,N_5141);
xor U12497 (N_12497,N_7997,N_8485);
xor U12498 (N_12498,N_6119,N_7026);
xor U12499 (N_12499,N_9293,N_7605);
nand U12500 (N_12500,N_7962,N_9552);
nand U12501 (N_12501,N_7648,N_8614);
xnor U12502 (N_12502,N_7668,N_9658);
or U12503 (N_12503,N_9856,N_7462);
nand U12504 (N_12504,N_5449,N_6285);
or U12505 (N_12505,N_5997,N_6679);
nor U12506 (N_12506,N_8946,N_9593);
and U12507 (N_12507,N_5673,N_9573);
nor U12508 (N_12508,N_8622,N_7668);
xor U12509 (N_12509,N_5594,N_6192);
xnor U12510 (N_12510,N_8014,N_7807);
or U12511 (N_12511,N_5459,N_7585);
or U12512 (N_12512,N_6964,N_9919);
xnor U12513 (N_12513,N_9770,N_8293);
or U12514 (N_12514,N_6288,N_6991);
and U12515 (N_12515,N_5829,N_8005);
nand U12516 (N_12516,N_7397,N_9306);
nand U12517 (N_12517,N_9977,N_9630);
nand U12518 (N_12518,N_9939,N_6795);
nand U12519 (N_12519,N_6614,N_5178);
or U12520 (N_12520,N_7353,N_7537);
xor U12521 (N_12521,N_6310,N_6214);
nand U12522 (N_12522,N_7768,N_8843);
xor U12523 (N_12523,N_9601,N_6475);
or U12524 (N_12524,N_5412,N_9258);
and U12525 (N_12525,N_9356,N_5139);
nor U12526 (N_12526,N_9668,N_9474);
xor U12527 (N_12527,N_8126,N_9147);
nor U12528 (N_12528,N_9709,N_9254);
nor U12529 (N_12529,N_8056,N_8841);
and U12530 (N_12530,N_9694,N_8788);
and U12531 (N_12531,N_7135,N_9777);
or U12532 (N_12532,N_6037,N_6341);
xnor U12533 (N_12533,N_6952,N_6303);
xnor U12534 (N_12534,N_6117,N_8144);
and U12535 (N_12535,N_5649,N_7290);
nand U12536 (N_12536,N_9001,N_7235);
and U12537 (N_12537,N_7722,N_5983);
nor U12538 (N_12538,N_7672,N_5771);
or U12539 (N_12539,N_6509,N_9075);
and U12540 (N_12540,N_8368,N_7094);
and U12541 (N_12541,N_5260,N_7681);
xnor U12542 (N_12542,N_5824,N_5159);
and U12543 (N_12543,N_6788,N_7792);
or U12544 (N_12544,N_9786,N_6564);
nor U12545 (N_12545,N_6682,N_5531);
nor U12546 (N_12546,N_7865,N_9764);
or U12547 (N_12547,N_5235,N_8317);
xor U12548 (N_12548,N_6092,N_9557);
nor U12549 (N_12549,N_6031,N_8755);
xor U12550 (N_12550,N_5317,N_9754);
nand U12551 (N_12551,N_9260,N_8735);
xnor U12552 (N_12552,N_6468,N_5075);
or U12553 (N_12553,N_5267,N_8145);
nand U12554 (N_12554,N_7098,N_9436);
and U12555 (N_12555,N_7179,N_9888);
xor U12556 (N_12556,N_6881,N_7816);
or U12557 (N_12557,N_9600,N_8189);
nor U12558 (N_12558,N_9798,N_9566);
nand U12559 (N_12559,N_9316,N_8824);
nand U12560 (N_12560,N_6880,N_6170);
and U12561 (N_12561,N_5445,N_7059);
xnor U12562 (N_12562,N_5329,N_9954);
or U12563 (N_12563,N_6166,N_8126);
and U12564 (N_12564,N_7575,N_6227);
or U12565 (N_12565,N_9947,N_8132);
or U12566 (N_12566,N_7311,N_5901);
nor U12567 (N_12567,N_9408,N_7667);
nand U12568 (N_12568,N_6548,N_7811);
nand U12569 (N_12569,N_6421,N_9498);
and U12570 (N_12570,N_5962,N_7461);
and U12571 (N_12571,N_7603,N_6559);
nand U12572 (N_12572,N_5713,N_9808);
or U12573 (N_12573,N_7498,N_8842);
and U12574 (N_12574,N_8998,N_8501);
or U12575 (N_12575,N_7246,N_7837);
xor U12576 (N_12576,N_9706,N_7960);
nor U12577 (N_12577,N_7060,N_9981);
or U12578 (N_12578,N_9598,N_7752);
or U12579 (N_12579,N_6271,N_5627);
nor U12580 (N_12580,N_7734,N_7566);
nand U12581 (N_12581,N_5056,N_6926);
nand U12582 (N_12582,N_6080,N_7648);
or U12583 (N_12583,N_8373,N_7781);
or U12584 (N_12584,N_9432,N_5970);
or U12585 (N_12585,N_9128,N_5486);
nand U12586 (N_12586,N_6523,N_5653);
xor U12587 (N_12587,N_6192,N_6936);
nor U12588 (N_12588,N_9698,N_7409);
or U12589 (N_12589,N_6681,N_5688);
xnor U12590 (N_12590,N_8066,N_6946);
or U12591 (N_12591,N_7342,N_9059);
and U12592 (N_12592,N_9301,N_7421);
and U12593 (N_12593,N_5567,N_6219);
xor U12594 (N_12594,N_9129,N_9957);
and U12595 (N_12595,N_9956,N_6064);
or U12596 (N_12596,N_8555,N_6497);
nor U12597 (N_12597,N_9971,N_7636);
nand U12598 (N_12598,N_9317,N_8618);
or U12599 (N_12599,N_9596,N_9901);
nor U12600 (N_12600,N_7358,N_8596);
nand U12601 (N_12601,N_8883,N_5829);
nand U12602 (N_12602,N_6601,N_6435);
or U12603 (N_12603,N_6016,N_6303);
nand U12604 (N_12604,N_5904,N_7716);
or U12605 (N_12605,N_7832,N_8689);
nand U12606 (N_12606,N_5356,N_7933);
and U12607 (N_12607,N_7897,N_5595);
xor U12608 (N_12608,N_6528,N_9936);
or U12609 (N_12609,N_5948,N_9574);
or U12610 (N_12610,N_9395,N_9778);
nor U12611 (N_12611,N_8215,N_5365);
or U12612 (N_12612,N_6318,N_6997);
and U12613 (N_12613,N_8117,N_6108);
nor U12614 (N_12614,N_9942,N_9541);
and U12615 (N_12615,N_8079,N_7368);
nor U12616 (N_12616,N_7984,N_6774);
or U12617 (N_12617,N_6981,N_5277);
or U12618 (N_12618,N_8681,N_9479);
nand U12619 (N_12619,N_5267,N_9802);
nor U12620 (N_12620,N_9424,N_7520);
or U12621 (N_12621,N_9282,N_6085);
or U12622 (N_12622,N_8199,N_6938);
nor U12623 (N_12623,N_6197,N_8406);
nand U12624 (N_12624,N_6950,N_9620);
xnor U12625 (N_12625,N_8809,N_7273);
or U12626 (N_12626,N_9025,N_7551);
and U12627 (N_12627,N_7708,N_8467);
and U12628 (N_12628,N_8057,N_9761);
or U12629 (N_12629,N_8739,N_5732);
or U12630 (N_12630,N_5896,N_5683);
or U12631 (N_12631,N_8038,N_6842);
nor U12632 (N_12632,N_6328,N_8065);
xor U12633 (N_12633,N_7268,N_5421);
and U12634 (N_12634,N_8881,N_6476);
nor U12635 (N_12635,N_7298,N_7839);
xor U12636 (N_12636,N_5788,N_9118);
nor U12637 (N_12637,N_9921,N_7880);
xnor U12638 (N_12638,N_7004,N_8731);
xnor U12639 (N_12639,N_8794,N_8877);
nor U12640 (N_12640,N_9051,N_7031);
xnor U12641 (N_12641,N_8859,N_6376);
xnor U12642 (N_12642,N_8369,N_9132);
or U12643 (N_12643,N_8724,N_5963);
or U12644 (N_12644,N_8145,N_7551);
nand U12645 (N_12645,N_7174,N_7050);
nor U12646 (N_12646,N_5862,N_6451);
or U12647 (N_12647,N_6151,N_7468);
or U12648 (N_12648,N_7659,N_5791);
and U12649 (N_12649,N_6503,N_7527);
nand U12650 (N_12650,N_5481,N_8922);
nand U12651 (N_12651,N_8562,N_7817);
and U12652 (N_12652,N_9178,N_6181);
or U12653 (N_12653,N_7627,N_8521);
nor U12654 (N_12654,N_8062,N_7443);
xor U12655 (N_12655,N_5801,N_9669);
or U12656 (N_12656,N_8559,N_5862);
nor U12657 (N_12657,N_5262,N_8340);
nand U12658 (N_12658,N_8440,N_8256);
and U12659 (N_12659,N_9975,N_6488);
nand U12660 (N_12660,N_7294,N_7124);
nand U12661 (N_12661,N_9317,N_6216);
nand U12662 (N_12662,N_7555,N_5339);
xor U12663 (N_12663,N_5424,N_7245);
nand U12664 (N_12664,N_9676,N_7437);
xnor U12665 (N_12665,N_7970,N_5547);
nand U12666 (N_12666,N_9745,N_7878);
nand U12667 (N_12667,N_7055,N_8024);
or U12668 (N_12668,N_8950,N_8606);
nor U12669 (N_12669,N_8625,N_8698);
xnor U12670 (N_12670,N_5650,N_9478);
xnor U12671 (N_12671,N_8754,N_9838);
and U12672 (N_12672,N_9988,N_5227);
nand U12673 (N_12673,N_6114,N_8850);
or U12674 (N_12674,N_8266,N_6127);
and U12675 (N_12675,N_6911,N_5322);
xor U12676 (N_12676,N_8007,N_5283);
and U12677 (N_12677,N_6990,N_8505);
nor U12678 (N_12678,N_8987,N_6462);
or U12679 (N_12679,N_5152,N_5423);
and U12680 (N_12680,N_6547,N_8841);
xor U12681 (N_12681,N_6226,N_5382);
xnor U12682 (N_12682,N_6832,N_7438);
or U12683 (N_12683,N_7092,N_7762);
nor U12684 (N_12684,N_9829,N_5711);
xor U12685 (N_12685,N_6307,N_9926);
nor U12686 (N_12686,N_8572,N_9652);
xnor U12687 (N_12687,N_7569,N_7969);
xor U12688 (N_12688,N_6638,N_7485);
or U12689 (N_12689,N_6532,N_8910);
and U12690 (N_12690,N_7626,N_5669);
xnor U12691 (N_12691,N_6584,N_8448);
nand U12692 (N_12692,N_8921,N_6688);
and U12693 (N_12693,N_8954,N_7538);
or U12694 (N_12694,N_7623,N_9472);
and U12695 (N_12695,N_9257,N_5121);
nor U12696 (N_12696,N_7746,N_6576);
nand U12697 (N_12697,N_7146,N_5891);
or U12698 (N_12698,N_9696,N_9320);
or U12699 (N_12699,N_7360,N_6033);
and U12700 (N_12700,N_6594,N_8345);
or U12701 (N_12701,N_7065,N_8180);
xor U12702 (N_12702,N_5359,N_6934);
nand U12703 (N_12703,N_9007,N_7691);
and U12704 (N_12704,N_6156,N_5702);
or U12705 (N_12705,N_6179,N_7492);
nor U12706 (N_12706,N_5263,N_8732);
xnor U12707 (N_12707,N_5838,N_9033);
xor U12708 (N_12708,N_8902,N_7892);
nand U12709 (N_12709,N_6098,N_6770);
or U12710 (N_12710,N_5575,N_9910);
nor U12711 (N_12711,N_7112,N_9296);
nand U12712 (N_12712,N_8447,N_5691);
xor U12713 (N_12713,N_5058,N_7260);
xor U12714 (N_12714,N_5039,N_8731);
or U12715 (N_12715,N_8922,N_9547);
nand U12716 (N_12716,N_6525,N_7155);
nor U12717 (N_12717,N_9112,N_7575);
and U12718 (N_12718,N_7154,N_5193);
xor U12719 (N_12719,N_6212,N_7032);
or U12720 (N_12720,N_5007,N_6840);
xnor U12721 (N_12721,N_6315,N_5768);
nor U12722 (N_12722,N_6717,N_8442);
nand U12723 (N_12723,N_9899,N_7918);
nor U12724 (N_12724,N_9513,N_5832);
nand U12725 (N_12725,N_8859,N_5419);
or U12726 (N_12726,N_8803,N_8315);
or U12727 (N_12727,N_7338,N_9627);
xnor U12728 (N_12728,N_9415,N_9655);
and U12729 (N_12729,N_8146,N_6074);
nor U12730 (N_12730,N_6342,N_5936);
or U12731 (N_12731,N_5921,N_7569);
and U12732 (N_12732,N_8562,N_5595);
xor U12733 (N_12733,N_6048,N_9257);
nand U12734 (N_12734,N_5273,N_5120);
nor U12735 (N_12735,N_7922,N_6638);
nand U12736 (N_12736,N_7527,N_8493);
xor U12737 (N_12737,N_6238,N_9442);
or U12738 (N_12738,N_8715,N_5797);
and U12739 (N_12739,N_5819,N_6046);
nor U12740 (N_12740,N_6875,N_6487);
or U12741 (N_12741,N_8448,N_5056);
xor U12742 (N_12742,N_8713,N_9607);
and U12743 (N_12743,N_9251,N_8200);
nor U12744 (N_12744,N_7877,N_7359);
or U12745 (N_12745,N_8708,N_8049);
or U12746 (N_12746,N_7163,N_5784);
nand U12747 (N_12747,N_8179,N_7183);
xnor U12748 (N_12748,N_5415,N_9782);
nand U12749 (N_12749,N_9844,N_9472);
and U12750 (N_12750,N_6553,N_5659);
xnor U12751 (N_12751,N_5998,N_7529);
or U12752 (N_12752,N_5057,N_6895);
or U12753 (N_12753,N_8845,N_8972);
nor U12754 (N_12754,N_8015,N_5032);
and U12755 (N_12755,N_5717,N_5035);
and U12756 (N_12756,N_9108,N_8206);
nand U12757 (N_12757,N_8932,N_5229);
or U12758 (N_12758,N_7748,N_9474);
nor U12759 (N_12759,N_6696,N_8089);
nor U12760 (N_12760,N_5338,N_5021);
nor U12761 (N_12761,N_6808,N_6101);
or U12762 (N_12762,N_5664,N_8947);
or U12763 (N_12763,N_9527,N_9241);
and U12764 (N_12764,N_9839,N_5788);
and U12765 (N_12765,N_9324,N_5441);
nand U12766 (N_12766,N_9808,N_5770);
or U12767 (N_12767,N_9637,N_7702);
or U12768 (N_12768,N_7578,N_6496);
or U12769 (N_12769,N_7489,N_9089);
and U12770 (N_12770,N_6573,N_8879);
nand U12771 (N_12771,N_8314,N_7266);
nor U12772 (N_12772,N_8875,N_8294);
or U12773 (N_12773,N_7014,N_7842);
and U12774 (N_12774,N_9778,N_6715);
xor U12775 (N_12775,N_6274,N_7432);
or U12776 (N_12776,N_9596,N_8986);
and U12777 (N_12777,N_7569,N_9313);
and U12778 (N_12778,N_6476,N_6788);
nor U12779 (N_12779,N_9905,N_9822);
and U12780 (N_12780,N_7393,N_9593);
xor U12781 (N_12781,N_9115,N_7442);
nand U12782 (N_12782,N_5409,N_8447);
nor U12783 (N_12783,N_5945,N_6861);
nor U12784 (N_12784,N_5881,N_7890);
xnor U12785 (N_12785,N_5948,N_8599);
xnor U12786 (N_12786,N_6079,N_7449);
nor U12787 (N_12787,N_6574,N_7530);
nor U12788 (N_12788,N_5517,N_9283);
xor U12789 (N_12789,N_9496,N_5384);
and U12790 (N_12790,N_6004,N_5814);
xor U12791 (N_12791,N_6786,N_7014);
and U12792 (N_12792,N_6541,N_9075);
or U12793 (N_12793,N_5652,N_8943);
nor U12794 (N_12794,N_8480,N_8461);
or U12795 (N_12795,N_8422,N_5710);
and U12796 (N_12796,N_6465,N_7394);
nor U12797 (N_12797,N_8843,N_7926);
or U12798 (N_12798,N_5476,N_5158);
or U12799 (N_12799,N_8973,N_6830);
nand U12800 (N_12800,N_8113,N_8039);
or U12801 (N_12801,N_8194,N_7723);
or U12802 (N_12802,N_6420,N_6108);
nor U12803 (N_12803,N_5327,N_6328);
xor U12804 (N_12804,N_5279,N_7520);
and U12805 (N_12805,N_9986,N_5569);
or U12806 (N_12806,N_7281,N_6409);
and U12807 (N_12807,N_7484,N_7043);
and U12808 (N_12808,N_8238,N_8030);
xnor U12809 (N_12809,N_5080,N_5867);
nand U12810 (N_12810,N_8425,N_8306);
nand U12811 (N_12811,N_6871,N_7655);
xnor U12812 (N_12812,N_9349,N_7276);
and U12813 (N_12813,N_6676,N_9613);
xor U12814 (N_12814,N_9444,N_9654);
xnor U12815 (N_12815,N_9982,N_6377);
xnor U12816 (N_12816,N_5687,N_7377);
and U12817 (N_12817,N_5753,N_5762);
and U12818 (N_12818,N_6633,N_9247);
nand U12819 (N_12819,N_9780,N_7213);
nand U12820 (N_12820,N_9388,N_5593);
xor U12821 (N_12821,N_9004,N_5100);
or U12822 (N_12822,N_5191,N_8848);
nor U12823 (N_12823,N_9762,N_8161);
nor U12824 (N_12824,N_6985,N_5774);
nor U12825 (N_12825,N_8504,N_5695);
and U12826 (N_12826,N_7901,N_6447);
or U12827 (N_12827,N_8011,N_7277);
xnor U12828 (N_12828,N_5402,N_9003);
nor U12829 (N_12829,N_7730,N_7434);
nand U12830 (N_12830,N_7455,N_7218);
nand U12831 (N_12831,N_7812,N_5549);
or U12832 (N_12832,N_9491,N_9063);
and U12833 (N_12833,N_6050,N_9342);
and U12834 (N_12834,N_8335,N_7202);
nand U12835 (N_12835,N_6782,N_5695);
nand U12836 (N_12836,N_6967,N_8451);
nor U12837 (N_12837,N_6192,N_9335);
or U12838 (N_12838,N_9448,N_7277);
or U12839 (N_12839,N_6797,N_6912);
nand U12840 (N_12840,N_9246,N_5954);
nand U12841 (N_12841,N_9079,N_8853);
nand U12842 (N_12842,N_5224,N_5221);
nand U12843 (N_12843,N_7683,N_6822);
and U12844 (N_12844,N_5438,N_8572);
xor U12845 (N_12845,N_8404,N_5281);
or U12846 (N_12846,N_6553,N_6787);
xnor U12847 (N_12847,N_8528,N_5201);
or U12848 (N_12848,N_8155,N_8654);
and U12849 (N_12849,N_7625,N_9936);
and U12850 (N_12850,N_6483,N_7233);
or U12851 (N_12851,N_9038,N_9353);
xnor U12852 (N_12852,N_9171,N_8359);
nand U12853 (N_12853,N_7044,N_9801);
and U12854 (N_12854,N_9452,N_8507);
xnor U12855 (N_12855,N_5783,N_6048);
and U12856 (N_12856,N_5099,N_6408);
nor U12857 (N_12857,N_6615,N_8321);
and U12858 (N_12858,N_9153,N_7163);
nand U12859 (N_12859,N_7315,N_7192);
and U12860 (N_12860,N_6554,N_5259);
xor U12861 (N_12861,N_9084,N_7802);
nand U12862 (N_12862,N_5082,N_7005);
or U12863 (N_12863,N_7465,N_7858);
nor U12864 (N_12864,N_8927,N_5240);
xor U12865 (N_12865,N_9940,N_6478);
nand U12866 (N_12866,N_6939,N_6993);
and U12867 (N_12867,N_6956,N_5635);
or U12868 (N_12868,N_6296,N_9834);
xor U12869 (N_12869,N_9704,N_5243);
nand U12870 (N_12870,N_9399,N_5090);
nor U12871 (N_12871,N_7061,N_9432);
and U12872 (N_12872,N_8974,N_8829);
nor U12873 (N_12873,N_9714,N_9255);
xor U12874 (N_12874,N_6520,N_5961);
nor U12875 (N_12875,N_5962,N_6351);
and U12876 (N_12876,N_8764,N_9937);
xor U12877 (N_12877,N_8196,N_7004);
xor U12878 (N_12878,N_9838,N_9165);
xor U12879 (N_12879,N_9280,N_8371);
or U12880 (N_12880,N_7592,N_5402);
nand U12881 (N_12881,N_7756,N_8203);
nand U12882 (N_12882,N_8701,N_5042);
and U12883 (N_12883,N_9194,N_5720);
or U12884 (N_12884,N_6349,N_7535);
nor U12885 (N_12885,N_5328,N_7123);
xor U12886 (N_12886,N_6131,N_9972);
nor U12887 (N_12887,N_6127,N_8023);
nor U12888 (N_12888,N_7924,N_9730);
nor U12889 (N_12889,N_5197,N_8500);
nor U12890 (N_12890,N_6467,N_7701);
nor U12891 (N_12891,N_8171,N_6148);
nor U12892 (N_12892,N_8881,N_6064);
xor U12893 (N_12893,N_7100,N_8488);
nor U12894 (N_12894,N_5671,N_9561);
xor U12895 (N_12895,N_9260,N_9301);
or U12896 (N_12896,N_9403,N_9618);
or U12897 (N_12897,N_6535,N_5862);
nor U12898 (N_12898,N_5022,N_5644);
xor U12899 (N_12899,N_6163,N_7846);
xnor U12900 (N_12900,N_9177,N_5882);
or U12901 (N_12901,N_8164,N_9846);
xnor U12902 (N_12902,N_6098,N_8400);
nand U12903 (N_12903,N_8028,N_8094);
nor U12904 (N_12904,N_5599,N_7394);
xnor U12905 (N_12905,N_7366,N_6898);
nand U12906 (N_12906,N_9821,N_6637);
nor U12907 (N_12907,N_7637,N_7274);
or U12908 (N_12908,N_6632,N_5237);
nor U12909 (N_12909,N_7437,N_9593);
and U12910 (N_12910,N_9312,N_7222);
or U12911 (N_12911,N_9574,N_5420);
and U12912 (N_12912,N_9784,N_8100);
nor U12913 (N_12913,N_6376,N_9457);
nand U12914 (N_12914,N_6629,N_6256);
nor U12915 (N_12915,N_6884,N_7680);
nand U12916 (N_12916,N_7265,N_9926);
and U12917 (N_12917,N_7900,N_7232);
xnor U12918 (N_12918,N_8625,N_9378);
xnor U12919 (N_12919,N_5421,N_7856);
and U12920 (N_12920,N_7426,N_7865);
nor U12921 (N_12921,N_9052,N_9016);
nor U12922 (N_12922,N_5289,N_6069);
nand U12923 (N_12923,N_8853,N_6998);
or U12924 (N_12924,N_7959,N_8125);
nor U12925 (N_12925,N_5483,N_5287);
xor U12926 (N_12926,N_5761,N_5385);
and U12927 (N_12927,N_5488,N_6355);
nand U12928 (N_12928,N_6138,N_9267);
xor U12929 (N_12929,N_7905,N_6057);
nor U12930 (N_12930,N_5510,N_7325);
xnor U12931 (N_12931,N_8121,N_6224);
or U12932 (N_12932,N_6127,N_6410);
or U12933 (N_12933,N_5888,N_6718);
nor U12934 (N_12934,N_9425,N_7938);
nand U12935 (N_12935,N_8157,N_7101);
and U12936 (N_12936,N_8288,N_6317);
nor U12937 (N_12937,N_9684,N_8071);
nand U12938 (N_12938,N_5192,N_7425);
and U12939 (N_12939,N_5457,N_5449);
xor U12940 (N_12940,N_8406,N_7210);
nand U12941 (N_12941,N_9626,N_7065);
nor U12942 (N_12942,N_5488,N_5613);
nor U12943 (N_12943,N_8553,N_7130);
xor U12944 (N_12944,N_6283,N_5164);
nor U12945 (N_12945,N_5872,N_8919);
or U12946 (N_12946,N_9109,N_5244);
or U12947 (N_12947,N_7869,N_5250);
or U12948 (N_12948,N_8106,N_6057);
nand U12949 (N_12949,N_5145,N_8087);
xor U12950 (N_12950,N_6217,N_8589);
nor U12951 (N_12951,N_5826,N_8380);
or U12952 (N_12952,N_9511,N_8177);
or U12953 (N_12953,N_5578,N_6291);
and U12954 (N_12954,N_8687,N_8311);
nor U12955 (N_12955,N_6938,N_8303);
and U12956 (N_12956,N_6389,N_8555);
and U12957 (N_12957,N_8907,N_5564);
and U12958 (N_12958,N_5139,N_5452);
xor U12959 (N_12959,N_7298,N_6109);
and U12960 (N_12960,N_9613,N_8801);
or U12961 (N_12961,N_8412,N_6123);
nand U12962 (N_12962,N_6021,N_6549);
xnor U12963 (N_12963,N_8230,N_9209);
and U12964 (N_12964,N_7706,N_8537);
nand U12965 (N_12965,N_8673,N_8310);
nand U12966 (N_12966,N_9437,N_9086);
and U12967 (N_12967,N_8794,N_6711);
nand U12968 (N_12968,N_6764,N_9497);
nor U12969 (N_12969,N_7464,N_8814);
nand U12970 (N_12970,N_6600,N_8964);
and U12971 (N_12971,N_9103,N_9500);
nor U12972 (N_12972,N_9901,N_6260);
xnor U12973 (N_12973,N_7992,N_6837);
and U12974 (N_12974,N_6116,N_9650);
and U12975 (N_12975,N_5336,N_8184);
nor U12976 (N_12976,N_5885,N_5318);
xor U12977 (N_12977,N_7501,N_7746);
or U12978 (N_12978,N_5648,N_6501);
and U12979 (N_12979,N_8200,N_7548);
nor U12980 (N_12980,N_5419,N_8376);
nand U12981 (N_12981,N_5351,N_5768);
nand U12982 (N_12982,N_6174,N_8574);
or U12983 (N_12983,N_8146,N_9395);
nor U12984 (N_12984,N_8002,N_5113);
nand U12985 (N_12985,N_8328,N_7198);
nor U12986 (N_12986,N_5950,N_7215);
nand U12987 (N_12987,N_6016,N_5423);
and U12988 (N_12988,N_9169,N_9184);
nor U12989 (N_12989,N_7238,N_5548);
or U12990 (N_12990,N_6810,N_9389);
xnor U12991 (N_12991,N_9132,N_7011);
nand U12992 (N_12992,N_6006,N_8937);
nor U12993 (N_12993,N_9063,N_9591);
nor U12994 (N_12994,N_6304,N_5137);
and U12995 (N_12995,N_6536,N_6863);
nor U12996 (N_12996,N_5351,N_8208);
or U12997 (N_12997,N_6999,N_6478);
or U12998 (N_12998,N_9383,N_9603);
xnor U12999 (N_12999,N_7982,N_6467);
and U13000 (N_13000,N_6221,N_9515);
xor U13001 (N_13001,N_9503,N_6964);
or U13002 (N_13002,N_5279,N_9936);
xnor U13003 (N_13003,N_8317,N_7134);
xnor U13004 (N_13004,N_6832,N_5402);
xor U13005 (N_13005,N_8501,N_6538);
or U13006 (N_13006,N_8117,N_6261);
and U13007 (N_13007,N_9482,N_5402);
or U13008 (N_13008,N_7879,N_5899);
or U13009 (N_13009,N_6930,N_5175);
nor U13010 (N_13010,N_8405,N_6577);
nor U13011 (N_13011,N_5264,N_6720);
nand U13012 (N_13012,N_7734,N_7441);
and U13013 (N_13013,N_6569,N_7321);
xor U13014 (N_13014,N_5645,N_5512);
xnor U13015 (N_13015,N_7077,N_9451);
nor U13016 (N_13016,N_6291,N_9852);
nor U13017 (N_13017,N_9700,N_6991);
xor U13018 (N_13018,N_8478,N_5638);
nand U13019 (N_13019,N_9885,N_6683);
nor U13020 (N_13020,N_8170,N_8529);
nor U13021 (N_13021,N_8280,N_8997);
nor U13022 (N_13022,N_6031,N_7919);
nor U13023 (N_13023,N_7659,N_9306);
xnor U13024 (N_13024,N_7033,N_5017);
nand U13025 (N_13025,N_5424,N_6317);
or U13026 (N_13026,N_5909,N_9494);
or U13027 (N_13027,N_8569,N_8632);
nand U13028 (N_13028,N_5113,N_5913);
xor U13029 (N_13029,N_5460,N_8135);
nor U13030 (N_13030,N_5125,N_5526);
nor U13031 (N_13031,N_6809,N_7502);
or U13032 (N_13032,N_6975,N_9124);
nor U13033 (N_13033,N_7849,N_9608);
nor U13034 (N_13034,N_7364,N_9971);
nor U13035 (N_13035,N_5773,N_7897);
xnor U13036 (N_13036,N_8721,N_8095);
nor U13037 (N_13037,N_6099,N_5361);
nand U13038 (N_13038,N_6624,N_8694);
nor U13039 (N_13039,N_9331,N_7794);
or U13040 (N_13040,N_9521,N_9099);
nand U13041 (N_13041,N_6543,N_6603);
and U13042 (N_13042,N_9477,N_8491);
xnor U13043 (N_13043,N_7755,N_8130);
nor U13044 (N_13044,N_8670,N_9669);
and U13045 (N_13045,N_6916,N_9722);
xor U13046 (N_13046,N_6040,N_9170);
and U13047 (N_13047,N_7766,N_5679);
xnor U13048 (N_13048,N_9273,N_6094);
nor U13049 (N_13049,N_7490,N_6621);
nand U13050 (N_13050,N_7012,N_8702);
nand U13051 (N_13051,N_5310,N_8741);
xor U13052 (N_13052,N_9345,N_7140);
nand U13053 (N_13053,N_5373,N_9940);
nor U13054 (N_13054,N_7395,N_9814);
nand U13055 (N_13055,N_5915,N_5803);
nand U13056 (N_13056,N_6852,N_5097);
nor U13057 (N_13057,N_8904,N_5262);
nor U13058 (N_13058,N_8382,N_5644);
nor U13059 (N_13059,N_6323,N_8964);
and U13060 (N_13060,N_6565,N_5128);
xor U13061 (N_13061,N_5001,N_5824);
nor U13062 (N_13062,N_9001,N_7372);
nand U13063 (N_13063,N_9953,N_8066);
nand U13064 (N_13064,N_5782,N_8460);
and U13065 (N_13065,N_6845,N_5290);
and U13066 (N_13066,N_5591,N_5215);
and U13067 (N_13067,N_8948,N_7884);
nand U13068 (N_13068,N_5828,N_5285);
nor U13069 (N_13069,N_9034,N_5575);
nor U13070 (N_13070,N_6315,N_9755);
or U13071 (N_13071,N_5003,N_8386);
xnor U13072 (N_13072,N_9355,N_8282);
or U13073 (N_13073,N_7081,N_5075);
or U13074 (N_13074,N_8382,N_5591);
xor U13075 (N_13075,N_5973,N_9179);
nor U13076 (N_13076,N_7440,N_8740);
xnor U13077 (N_13077,N_7541,N_5300);
nand U13078 (N_13078,N_5051,N_7473);
nor U13079 (N_13079,N_9653,N_7758);
xnor U13080 (N_13080,N_6542,N_7065);
nor U13081 (N_13081,N_9495,N_6662);
or U13082 (N_13082,N_7377,N_7081);
or U13083 (N_13083,N_5308,N_5902);
and U13084 (N_13084,N_5758,N_9327);
nand U13085 (N_13085,N_9386,N_9609);
nor U13086 (N_13086,N_6151,N_6855);
xnor U13087 (N_13087,N_8160,N_7663);
xnor U13088 (N_13088,N_9480,N_9629);
and U13089 (N_13089,N_9862,N_6757);
nand U13090 (N_13090,N_9137,N_6946);
and U13091 (N_13091,N_9578,N_5345);
or U13092 (N_13092,N_6671,N_7236);
nand U13093 (N_13093,N_6810,N_6839);
xnor U13094 (N_13094,N_7665,N_7690);
and U13095 (N_13095,N_5813,N_8653);
nor U13096 (N_13096,N_7494,N_6926);
xor U13097 (N_13097,N_8454,N_8800);
nand U13098 (N_13098,N_8644,N_7736);
or U13099 (N_13099,N_8537,N_7024);
nor U13100 (N_13100,N_9339,N_7715);
or U13101 (N_13101,N_7099,N_6931);
or U13102 (N_13102,N_8762,N_7826);
nand U13103 (N_13103,N_8596,N_8244);
nand U13104 (N_13104,N_6602,N_7403);
xnor U13105 (N_13105,N_7739,N_9255);
xnor U13106 (N_13106,N_9754,N_6685);
and U13107 (N_13107,N_6418,N_5895);
nand U13108 (N_13108,N_7412,N_6295);
nor U13109 (N_13109,N_7440,N_7112);
nor U13110 (N_13110,N_8499,N_7981);
or U13111 (N_13111,N_6977,N_5449);
nor U13112 (N_13112,N_7658,N_9973);
xor U13113 (N_13113,N_8944,N_8416);
nand U13114 (N_13114,N_6664,N_8812);
nor U13115 (N_13115,N_6130,N_6560);
xor U13116 (N_13116,N_5388,N_6724);
nor U13117 (N_13117,N_7253,N_7798);
nor U13118 (N_13118,N_9954,N_7769);
or U13119 (N_13119,N_7174,N_6254);
nor U13120 (N_13120,N_8418,N_6746);
or U13121 (N_13121,N_8702,N_8045);
and U13122 (N_13122,N_6665,N_5612);
xnor U13123 (N_13123,N_7927,N_8272);
xnor U13124 (N_13124,N_6400,N_6845);
and U13125 (N_13125,N_5128,N_7195);
or U13126 (N_13126,N_9133,N_6186);
nand U13127 (N_13127,N_6493,N_9954);
and U13128 (N_13128,N_8212,N_5580);
xnor U13129 (N_13129,N_9927,N_8743);
xnor U13130 (N_13130,N_6242,N_9763);
and U13131 (N_13131,N_8947,N_5255);
xor U13132 (N_13132,N_6919,N_5119);
nand U13133 (N_13133,N_5828,N_8590);
nand U13134 (N_13134,N_5847,N_5322);
nor U13135 (N_13135,N_6552,N_6775);
or U13136 (N_13136,N_5895,N_7108);
and U13137 (N_13137,N_5826,N_5226);
and U13138 (N_13138,N_7236,N_5140);
xor U13139 (N_13139,N_8924,N_9716);
xnor U13140 (N_13140,N_6090,N_5924);
nand U13141 (N_13141,N_5365,N_9561);
and U13142 (N_13142,N_9842,N_9510);
xor U13143 (N_13143,N_5127,N_5345);
or U13144 (N_13144,N_9571,N_6665);
and U13145 (N_13145,N_7236,N_9673);
and U13146 (N_13146,N_9139,N_9353);
nor U13147 (N_13147,N_7408,N_5920);
xor U13148 (N_13148,N_5512,N_7537);
or U13149 (N_13149,N_7468,N_9360);
or U13150 (N_13150,N_6182,N_7939);
nand U13151 (N_13151,N_7646,N_7192);
and U13152 (N_13152,N_6181,N_9234);
or U13153 (N_13153,N_8026,N_7644);
or U13154 (N_13154,N_9539,N_6922);
and U13155 (N_13155,N_7481,N_7101);
nor U13156 (N_13156,N_8550,N_5589);
and U13157 (N_13157,N_7905,N_8965);
and U13158 (N_13158,N_5954,N_8503);
and U13159 (N_13159,N_5320,N_9228);
and U13160 (N_13160,N_5570,N_5385);
or U13161 (N_13161,N_8840,N_9980);
nor U13162 (N_13162,N_9116,N_9445);
or U13163 (N_13163,N_6552,N_8865);
or U13164 (N_13164,N_5283,N_8712);
nor U13165 (N_13165,N_6188,N_6716);
or U13166 (N_13166,N_7626,N_7650);
and U13167 (N_13167,N_7720,N_8539);
or U13168 (N_13168,N_9591,N_8950);
xor U13169 (N_13169,N_9427,N_6737);
nand U13170 (N_13170,N_6499,N_8485);
or U13171 (N_13171,N_8137,N_7927);
xnor U13172 (N_13172,N_7721,N_8029);
or U13173 (N_13173,N_9911,N_9118);
nand U13174 (N_13174,N_6567,N_5034);
xnor U13175 (N_13175,N_5457,N_5453);
and U13176 (N_13176,N_5952,N_9610);
or U13177 (N_13177,N_8390,N_8109);
or U13178 (N_13178,N_8909,N_8045);
nand U13179 (N_13179,N_9460,N_9011);
xor U13180 (N_13180,N_8644,N_7348);
or U13181 (N_13181,N_9055,N_8436);
nand U13182 (N_13182,N_7431,N_5149);
or U13183 (N_13183,N_8098,N_9336);
and U13184 (N_13184,N_8646,N_9490);
xnor U13185 (N_13185,N_7060,N_9092);
nand U13186 (N_13186,N_6446,N_5123);
and U13187 (N_13187,N_9575,N_7399);
nand U13188 (N_13188,N_9930,N_8378);
and U13189 (N_13189,N_7634,N_9379);
and U13190 (N_13190,N_7801,N_5204);
xnor U13191 (N_13191,N_8896,N_5304);
nor U13192 (N_13192,N_6693,N_6960);
or U13193 (N_13193,N_8586,N_9105);
and U13194 (N_13194,N_5159,N_5959);
and U13195 (N_13195,N_7247,N_7697);
nand U13196 (N_13196,N_9068,N_8606);
nor U13197 (N_13197,N_7618,N_6471);
nand U13198 (N_13198,N_7878,N_6631);
or U13199 (N_13199,N_6898,N_5430);
and U13200 (N_13200,N_7479,N_9425);
and U13201 (N_13201,N_8153,N_6282);
and U13202 (N_13202,N_8180,N_7778);
nand U13203 (N_13203,N_6281,N_9704);
nor U13204 (N_13204,N_6154,N_8956);
xnor U13205 (N_13205,N_6429,N_9172);
nor U13206 (N_13206,N_5176,N_8698);
nand U13207 (N_13207,N_7955,N_5079);
nor U13208 (N_13208,N_5316,N_8711);
or U13209 (N_13209,N_9113,N_5789);
or U13210 (N_13210,N_7551,N_8720);
or U13211 (N_13211,N_9821,N_8045);
nand U13212 (N_13212,N_6999,N_7312);
nor U13213 (N_13213,N_6819,N_8611);
xnor U13214 (N_13214,N_8368,N_6680);
and U13215 (N_13215,N_8569,N_5797);
or U13216 (N_13216,N_6592,N_5357);
nand U13217 (N_13217,N_7341,N_5572);
nand U13218 (N_13218,N_5175,N_9927);
and U13219 (N_13219,N_8479,N_5321);
nand U13220 (N_13220,N_5941,N_6634);
nand U13221 (N_13221,N_7821,N_7860);
nand U13222 (N_13222,N_6455,N_6227);
and U13223 (N_13223,N_6307,N_9912);
nand U13224 (N_13224,N_8332,N_7964);
and U13225 (N_13225,N_8523,N_5507);
nand U13226 (N_13226,N_6695,N_5227);
or U13227 (N_13227,N_8190,N_9112);
and U13228 (N_13228,N_7195,N_9946);
xnor U13229 (N_13229,N_6429,N_7826);
nand U13230 (N_13230,N_5292,N_6647);
nand U13231 (N_13231,N_9874,N_6382);
nand U13232 (N_13232,N_9859,N_8214);
or U13233 (N_13233,N_6611,N_6523);
or U13234 (N_13234,N_9140,N_7024);
or U13235 (N_13235,N_9146,N_6152);
and U13236 (N_13236,N_9487,N_7137);
xnor U13237 (N_13237,N_9620,N_8179);
nor U13238 (N_13238,N_7111,N_9624);
nor U13239 (N_13239,N_7849,N_9678);
nand U13240 (N_13240,N_8047,N_6461);
nor U13241 (N_13241,N_5887,N_5579);
xor U13242 (N_13242,N_6325,N_7691);
nand U13243 (N_13243,N_5346,N_5230);
nand U13244 (N_13244,N_5313,N_7361);
or U13245 (N_13245,N_5332,N_6133);
or U13246 (N_13246,N_7691,N_9746);
nand U13247 (N_13247,N_5974,N_5764);
and U13248 (N_13248,N_5461,N_6576);
or U13249 (N_13249,N_7086,N_9306);
or U13250 (N_13250,N_5496,N_8106);
or U13251 (N_13251,N_9819,N_9513);
or U13252 (N_13252,N_6227,N_9876);
or U13253 (N_13253,N_8661,N_8876);
or U13254 (N_13254,N_7104,N_9729);
xor U13255 (N_13255,N_9352,N_9931);
nor U13256 (N_13256,N_5668,N_5648);
xor U13257 (N_13257,N_8880,N_6427);
nor U13258 (N_13258,N_9468,N_9419);
nor U13259 (N_13259,N_8657,N_6791);
or U13260 (N_13260,N_7239,N_8249);
xnor U13261 (N_13261,N_5195,N_9026);
nand U13262 (N_13262,N_8175,N_9487);
or U13263 (N_13263,N_8802,N_5743);
xnor U13264 (N_13264,N_7780,N_5699);
and U13265 (N_13265,N_8726,N_5001);
or U13266 (N_13266,N_9727,N_8168);
nand U13267 (N_13267,N_8360,N_7445);
nor U13268 (N_13268,N_5670,N_6669);
or U13269 (N_13269,N_9210,N_7823);
xnor U13270 (N_13270,N_5092,N_6541);
nand U13271 (N_13271,N_8944,N_6235);
nand U13272 (N_13272,N_5770,N_8313);
and U13273 (N_13273,N_9068,N_9882);
xor U13274 (N_13274,N_8662,N_7000);
nand U13275 (N_13275,N_9558,N_9570);
nand U13276 (N_13276,N_6678,N_6145);
and U13277 (N_13277,N_8711,N_6655);
nor U13278 (N_13278,N_7402,N_7187);
or U13279 (N_13279,N_8269,N_6152);
and U13280 (N_13280,N_9646,N_5679);
and U13281 (N_13281,N_5903,N_9242);
xnor U13282 (N_13282,N_7976,N_6267);
nor U13283 (N_13283,N_9229,N_9640);
xnor U13284 (N_13284,N_7078,N_6780);
or U13285 (N_13285,N_8269,N_5308);
and U13286 (N_13286,N_9934,N_7344);
xnor U13287 (N_13287,N_7291,N_7991);
xor U13288 (N_13288,N_5822,N_7138);
xnor U13289 (N_13289,N_6553,N_8508);
and U13290 (N_13290,N_5421,N_6947);
and U13291 (N_13291,N_7138,N_5828);
and U13292 (N_13292,N_9555,N_6110);
or U13293 (N_13293,N_7571,N_8997);
nor U13294 (N_13294,N_7868,N_6563);
and U13295 (N_13295,N_5410,N_7135);
nor U13296 (N_13296,N_6025,N_8193);
nor U13297 (N_13297,N_9795,N_9488);
and U13298 (N_13298,N_6783,N_9030);
nor U13299 (N_13299,N_8600,N_7899);
and U13300 (N_13300,N_5462,N_8838);
and U13301 (N_13301,N_5767,N_5932);
or U13302 (N_13302,N_7855,N_8782);
xor U13303 (N_13303,N_9864,N_9517);
nor U13304 (N_13304,N_8092,N_5270);
or U13305 (N_13305,N_9740,N_7958);
nor U13306 (N_13306,N_5648,N_5898);
nand U13307 (N_13307,N_7102,N_6376);
nand U13308 (N_13308,N_6433,N_8445);
and U13309 (N_13309,N_7879,N_9639);
nor U13310 (N_13310,N_9264,N_6423);
xnor U13311 (N_13311,N_5125,N_7312);
and U13312 (N_13312,N_7078,N_9119);
or U13313 (N_13313,N_5860,N_5092);
nand U13314 (N_13314,N_9845,N_8477);
or U13315 (N_13315,N_8335,N_6682);
nor U13316 (N_13316,N_8871,N_6704);
nor U13317 (N_13317,N_7080,N_6388);
and U13318 (N_13318,N_5341,N_7887);
nand U13319 (N_13319,N_9460,N_8284);
or U13320 (N_13320,N_9403,N_6637);
xor U13321 (N_13321,N_9792,N_8310);
nor U13322 (N_13322,N_6923,N_7337);
and U13323 (N_13323,N_9727,N_5198);
and U13324 (N_13324,N_6868,N_9521);
xor U13325 (N_13325,N_5537,N_7996);
nand U13326 (N_13326,N_9637,N_5745);
and U13327 (N_13327,N_7327,N_9006);
nand U13328 (N_13328,N_7468,N_7563);
nor U13329 (N_13329,N_6729,N_6364);
nand U13330 (N_13330,N_5222,N_7485);
nand U13331 (N_13331,N_5365,N_5251);
nor U13332 (N_13332,N_7847,N_8227);
nand U13333 (N_13333,N_7948,N_5088);
xnor U13334 (N_13334,N_5890,N_7803);
nor U13335 (N_13335,N_8959,N_5570);
xor U13336 (N_13336,N_6723,N_5506);
nand U13337 (N_13337,N_6733,N_5640);
and U13338 (N_13338,N_8682,N_8606);
xor U13339 (N_13339,N_9685,N_5697);
and U13340 (N_13340,N_7186,N_8187);
and U13341 (N_13341,N_5845,N_6872);
nand U13342 (N_13342,N_5651,N_5215);
nor U13343 (N_13343,N_6071,N_9666);
and U13344 (N_13344,N_9343,N_8154);
xnor U13345 (N_13345,N_7791,N_6067);
and U13346 (N_13346,N_8856,N_7430);
or U13347 (N_13347,N_5705,N_7581);
nand U13348 (N_13348,N_7229,N_7201);
or U13349 (N_13349,N_5135,N_8617);
nor U13350 (N_13350,N_5700,N_5064);
nor U13351 (N_13351,N_7072,N_9721);
nor U13352 (N_13352,N_9329,N_5312);
nor U13353 (N_13353,N_8365,N_5659);
or U13354 (N_13354,N_7703,N_8022);
and U13355 (N_13355,N_6341,N_6026);
nor U13356 (N_13356,N_9540,N_5469);
xor U13357 (N_13357,N_5441,N_9406);
xor U13358 (N_13358,N_6654,N_6316);
nand U13359 (N_13359,N_6281,N_5899);
nand U13360 (N_13360,N_9644,N_6281);
xnor U13361 (N_13361,N_8231,N_6622);
nand U13362 (N_13362,N_5502,N_9638);
and U13363 (N_13363,N_6087,N_9021);
nand U13364 (N_13364,N_6038,N_9017);
and U13365 (N_13365,N_9225,N_5113);
and U13366 (N_13366,N_9109,N_8123);
xor U13367 (N_13367,N_9616,N_8425);
xor U13368 (N_13368,N_9364,N_6439);
xor U13369 (N_13369,N_9001,N_5937);
nand U13370 (N_13370,N_9743,N_6816);
nand U13371 (N_13371,N_5621,N_5980);
and U13372 (N_13372,N_7055,N_8742);
xnor U13373 (N_13373,N_8815,N_5413);
or U13374 (N_13374,N_9116,N_8767);
nand U13375 (N_13375,N_5567,N_9163);
or U13376 (N_13376,N_7146,N_8645);
or U13377 (N_13377,N_5903,N_9862);
and U13378 (N_13378,N_6177,N_5765);
xnor U13379 (N_13379,N_6022,N_6870);
or U13380 (N_13380,N_8113,N_7907);
xnor U13381 (N_13381,N_8336,N_9594);
xor U13382 (N_13382,N_6224,N_9431);
or U13383 (N_13383,N_9789,N_7043);
and U13384 (N_13384,N_6297,N_5622);
or U13385 (N_13385,N_7395,N_8177);
nand U13386 (N_13386,N_5681,N_8320);
xor U13387 (N_13387,N_6658,N_8674);
or U13388 (N_13388,N_6111,N_6886);
or U13389 (N_13389,N_8920,N_6324);
and U13390 (N_13390,N_5415,N_8637);
and U13391 (N_13391,N_8266,N_5323);
nor U13392 (N_13392,N_8266,N_8522);
nand U13393 (N_13393,N_8035,N_8509);
nor U13394 (N_13394,N_8698,N_7203);
xor U13395 (N_13395,N_5697,N_7169);
xor U13396 (N_13396,N_9099,N_9832);
xor U13397 (N_13397,N_5414,N_7295);
or U13398 (N_13398,N_8369,N_5426);
nor U13399 (N_13399,N_6876,N_9438);
nor U13400 (N_13400,N_8563,N_8417);
nor U13401 (N_13401,N_7361,N_6250);
and U13402 (N_13402,N_7976,N_5947);
or U13403 (N_13403,N_6891,N_8093);
or U13404 (N_13404,N_7157,N_9220);
or U13405 (N_13405,N_5181,N_7934);
nor U13406 (N_13406,N_9855,N_8487);
and U13407 (N_13407,N_7505,N_6614);
xnor U13408 (N_13408,N_7346,N_8858);
and U13409 (N_13409,N_7760,N_6342);
nand U13410 (N_13410,N_5517,N_5468);
xor U13411 (N_13411,N_6273,N_5387);
nor U13412 (N_13412,N_9939,N_5904);
and U13413 (N_13413,N_7096,N_5161);
nor U13414 (N_13414,N_8164,N_8296);
xor U13415 (N_13415,N_6618,N_6310);
nor U13416 (N_13416,N_5086,N_5671);
and U13417 (N_13417,N_6096,N_8840);
xor U13418 (N_13418,N_5895,N_9427);
nand U13419 (N_13419,N_5041,N_9712);
xor U13420 (N_13420,N_6665,N_6614);
nor U13421 (N_13421,N_5120,N_8235);
xnor U13422 (N_13422,N_7092,N_6571);
xnor U13423 (N_13423,N_6280,N_7574);
and U13424 (N_13424,N_5634,N_5659);
and U13425 (N_13425,N_5438,N_7387);
and U13426 (N_13426,N_5216,N_8729);
xnor U13427 (N_13427,N_9167,N_8996);
and U13428 (N_13428,N_5742,N_6712);
nand U13429 (N_13429,N_5639,N_6351);
or U13430 (N_13430,N_9771,N_7300);
xnor U13431 (N_13431,N_6664,N_6137);
and U13432 (N_13432,N_8764,N_9203);
and U13433 (N_13433,N_5087,N_5324);
and U13434 (N_13434,N_5465,N_8706);
xor U13435 (N_13435,N_8745,N_9076);
xnor U13436 (N_13436,N_9830,N_8538);
nand U13437 (N_13437,N_9773,N_5227);
and U13438 (N_13438,N_7649,N_5869);
xnor U13439 (N_13439,N_5948,N_8940);
nand U13440 (N_13440,N_7743,N_5129);
and U13441 (N_13441,N_6966,N_7050);
and U13442 (N_13442,N_5711,N_6541);
or U13443 (N_13443,N_8202,N_5381);
and U13444 (N_13444,N_5995,N_5573);
nor U13445 (N_13445,N_8870,N_7776);
xor U13446 (N_13446,N_7313,N_5913);
nand U13447 (N_13447,N_6759,N_7363);
or U13448 (N_13448,N_8438,N_5740);
and U13449 (N_13449,N_8612,N_6412);
nand U13450 (N_13450,N_8948,N_7707);
xor U13451 (N_13451,N_6853,N_6754);
xor U13452 (N_13452,N_8481,N_5358);
nand U13453 (N_13453,N_5144,N_7171);
or U13454 (N_13454,N_6683,N_5588);
nor U13455 (N_13455,N_9965,N_9185);
xor U13456 (N_13456,N_9985,N_9274);
nor U13457 (N_13457,N_7645,N_5939);
nand U13458 (N_13458,N_6975,N_7019);
xor U13459 (N_13459,N_6116,N_7189);
and U13460 (N_13460,N_6589,N_8087);
nand U13461 (N_13461,N_9821,N_7272);
and U13462 (N_13462,N_8281,N_8988);
nor U13463 (N_13463,N_9449,N_6161);
nand U13464 (N_13464,N_8238,N_8085);
nor U13465 (N_13465,N_9528,N_5091);
and U13466 (N_13466,N_8500,N_9082);
or U13467 (N_13467,N_7909,N_5243);
and U13468 (N_13468,N_9044,N_7972);
xnor U13469 (N_13469,N_8226,N_7124);
nand U13470 (N_13470,N_7322,N_5728);
nand U13471 (N_13471,N_6535,N_7934);
xor U13472 (N_13472,N_9766,N_7011);
nand U13473 (N_13473,N_7062,N_8079);
and U13474 (N_13474,N_7442,N_9778);
and U13475 (N_13475,N_7666,N_8014);
and U13476 (N_13476,N_6602,N_9707);
xnor U13477 (N_13477,N_6196,N_6626);
xor U13478 (N_13478,N_6212,N_6779);
nor U13479 (N_13479,N_9911,N_8423);
xor U13480 (N_13480,N_6235,N_6480);
nor U13481 (N_13481,N_8575,N_5899);
or U13482 (N_13482,N_8086,N_6558);
xnor U13483 (N_13483,N_8504,N_7310);
or U13484 (N_13484,N_5084,N_7929);
xnor U13485 (N_13485,N_8750,N_7352);
or U13486 (N_13486,N_7230,N_7382);
or U13487 (N_13487,N_7893,N_7858);
xor U13488 (N_13488,N_6484,N_6345);
or U13489 (N_13489,N_8767,N_9276);
nor U13490 (N_13490,N_9351,N_8719);
or U13491 (N_13491,N_8634,N_9155);
nand U13492 (N_13492,N_8101,N_7435);
and U13493 (N_13493,N_7649,N_6136);
nand U13494 (N_13494,N_8337,N_9073);
nor U13495 (N_13495,N_6951,N_9079);
nand U13496 (N_13496,N_9401,N_8902);
nor U13497 (N_13497,N_6571,N_5988);
xnor U13498 (N_13498,N_8888,N_6842);
or U13499 (N_13499,N_9935,N_8436);
xnor U13500 (N_13500,N_6565,N_5789);
and U13501 (N_13501,N_6824,N_5941);
and U13502 (N_13502,N_7749,N_7598);
xor U13503 (N_13503,N_7157,N_8702);
or U13504 (N_13504,N_5665,N_9059);
or U13505 (N_13505,N_6380,N_5208);
nor U13506 (N_13506,N_8412,N_6312);
nor U13507 (N_13507,N_9458,N_6448);
nor U13508 (N_13508,N_6449,N_9496);
and U13509 (N_13509,N_8857,N_5504);
nor U13510 (N_13510,N_9145,N_9414);
or U13511 (N_13511,N_8487,N_7745);
nand U13512 (N_13512,N_7707,N_6469);
or U13513 (N_13513,N_6857,N_8597);
xor U13514 (N_13514,N_6522,N_5782);
nor U13515 (N_13515,N_8800,N_8584);
nor U13516 (N_13516,N_8183,N_6475);
or U13517 (N_13517,N_6295,N_7402);
xnor U13518 (N_13518,N_7342,N_5734);
and U13519 (N_13519,N_5509,N_5706);
and U13520 (N_13520,N_6990,N_9805);
xnor U13521 (N_13521,N_7262,N_7073);
xnor U13522 (N_13522,N_5979,N_8934);
and U13523 (N_13523,N_6147,N_7344);
nand U13524 (N_13524,N_6297,N_6976);
nand U13525 (N_13525,N_5952,N_8005);
xnor U13526 (N_13526,N_9754,N_6307);
xnor U13527 (N_13527,N_5165,N_7945);
nor U13528 (N_13528,N_5488,N_9269);
nand U13529 (N_13529,N_5751,N_8438);
nor U13530 (N_13530,N_7484,N_6435);
and U13531 (N_13531,N_6231,N_8396);
nand U13532 (N_13532,N_6971,N_5272);
xnor U13533 (N_13533,N_9332,N_6169);
or U13534 (N_13534,N_6024,N_8543);
or U13535 (N_13535,N_7914,N_8844);
xnor U13536 (N_13536,N_7434,N_8176);
xnor U13537 (N_13537,N_8530,N_6272);
xor U13538 (N_13538,N_6425,N_8540);
xor U13539 (N_13539,N_8070,N_5832);
nand U13540 (N_13540,N_8859,N_7800);
nor U13541 (N_13541,N_6812,N_9390);
nor U13542 (N_13542,N_5357,N_9906);
and U13543 (N_13543,N_9977,N_8464);
nor U13544 (N_13544,N_5540,N_5193);
and U13545 (N_13545,N_5742,N_7326);
nor U13546 (N_13546,N_6902,N_5760);
nor U13547 (N_13547,N_6595,N_5134);
xor U13548 (N_13548,N_5265,N_6450);
nand U13549 (N_13549,N_7915,N_7256);
and U13550 (N_13550,N_9584,N_6333);
or U13551 (N_13551,N_6668,N_8644);
nor U13552 (N_13552,N_6624,N_7006);
or U13553 (N_13553,N_6445,N_6993);
xnor U13554 (N_13554,N_6456,N_9565);
and U13555 (N_13555,N_5340,N_9181);
nor U13556 (N_13556,N_9256,N_7754);
nand U13557 (N_13557,N_8248,N_6007);
and U13558 (N_13558,N_6861,N_6647);
nor U13559 (N_13559,N_5963,N_5840);
nor U13560 (N_13560,N_5889,N_9829);
and U13561 (N_13561,N_9402,N_6573);
nand U13562 (N_13562,N_5272,N_6302);
or U13563 (N_13563,N_8579,N_7445);
or U13564 (N_13564,N_7347,N_8293);
and U13565 (N_13565,N_7055,N_7413);
nand U13566 (N_13566,N_8144,N_6629);
xor U13567 (N_13567,N_6009,N_8130);
nand U13568 (N_13568,N_5767,N_8419);
xor U13569 (N_13569,N_6721,N_9949);
nand U13570 (N_13570,N_5183,N_6823);
and U13571 (N_13571,N_8890,N_7299);
and U13572 (N_13572,N_8713,N_5481);
or U13573 (N_13573,N_5055,N_5737);
nand U13574 (N_13574,N_5760,N_5116);
nand U13575 (N_13575,N_5264,N_6933);
nand U13576 (N_13576,N_5100,N_5339);
xor U13577 (N_13577,N_9437,N_7033);
nor U13578 (N_13578,N_8908,N_5317);
nand U13579 (N_13579,N_8622,N_9314);
or U13580 (N_13580,N_8041,N_6079);
and U13581 (N_13581,N_8002,N_7110);
nor U13582 (N_13582,N_8990,N_6662);
and U13583 (N_13583,N_5847,N_7648);
xnor U13584 (N_13584,N_6562,N_5434);
nor U13585 (N_13585,N_9366,N_7528);
xor U13586 (N_13586,N_7070,N_6070);
nand U13587 (N_13587,N_5722,N_6064);
nand U13588 (N_13588,N_8437,N_8248);
nor U13589 (N_13589,N_9238,N_7680);
and U13590 (N_13590,N_6998,N_6477);
nor U13591 (N_13591,N_6251,N_5183);
nand U13592 (N_13592,N_9016,N_8844);
nor U13593 (N_13593,N_5473,N_5196);
or U13594 (N_13594,N_9900,N_9572);
xnor U13595 (N_13595,N_6623,N_9036);
and U13596 (N_13596,N_7711,N_5110);
nand U13597 (N_13597,N_5130,N_8384);
nor U13598 (N_13598,N_6387,N_6617);
xor U13599 (N_13599,N_9943,N_8232);
or U13600 (N_13600,N_6185,N_7521);
nand U13601 (N_13601,N_7700,N_6177);
or U13602 (N_13602,N_6901,N_6432);
nor U13603 (N_13603,N_9628,N_6372);
nand U13604 (N_13604,N_9790,N_5952);
xnor U13605 (N_13605,N_7778,N_9755);
nand U13606 (N_13606,N_8299,N_7244);
xor U13607 (N_13607,N_8858,N_6888);
nor U13608 (N_13608,N_9114,N_7620);
nand U13609 (N_13609,N_9726,N_5322);
or U13610 (N_13610,N_7231,N_9280);
nand U13611 (N_13611,N_9153,N_6642);
or U13612 (N_13612,N_7303,N_5546);
xor U13613 (N_13613,N_5771,N_8629);
and U13614 (N_13614,N_8336,N_6388);
nand U13615 (N_13615,N_7531,N_9556);
and U13616 (N_13616,N_7113,N_7428);
and U13617 (N_13617,N_7762,N_6879);
and U13618 (N_13618,N_9925,N_6072);
or U13619 (N_13619,N_6785,N_9372);
or U13620 (N_13620,N_6337,N_8046);
and U13621 (N_13621,N_9920,N_5738);
xnor U13622 (N_13622,N_5511,N_5298);
and U13623 (N_13623,N_8915,N_6534);
nor U13624 (N_13624,N_9758,N_7139);
nand U13625 (N_13625,N_7230,N_7945);
nand U13626 (N_13626,N_6914,N_7868);
xnor U13627 (N_13627,N_9703,N_6244);
or U13628 (N_13628,N_5347,N_6454);
xnor U13629 (N_13629,N_9064,N_5582);
nand U13630 (N_13630,N_5768,N_6667);
nor U13631 (N_13631,N_6891,N_6836);
nor U13632 (N_13632,N_6354,N_7823);
nor U13633 (N_13633,N_7073,N_8499);
and U13634 (N_13634,N_7331,N_5894);
xnor U13635 (N_13635,N_5794,N_9806);
or U13636 (N_13636,N_5103,N_8967);
and U13637 (N_13637,N_6981,N_5598);
nor U13638 (N_13638,N_8744,N_9116);
xnor U13639 (N_13639,N_7249,N_9373);
xnor U13640 (N_13640,N_5234,N_8148);
xor U13641 (N_13641,N_8956,N_9349);
nand U13642 (N_13642,N_6494,N_5929);
and U13643 (N_13643,N_7277,N_5831);
or U13644 (N_13644,N_6229,N_9468);
xnor U13645 (N_13645,N_6735,N_6186);
or U13646 (N_13646,N_6105,N_6602);
and U13647 (N_13647,N_8488,N_7810);
xnor U13648 (N_13648,N_6198,N_7775);
nand U13649 (N_13649,N_9067,N_9459);
nor U13650 (N_13650,N_5569,N_7373);
nand U13651 (N_13651,N_9388,N_7086);
and U13652 (N_13652,N_6676,N_5660);
xor U13653 (N_13653,N_9811,N_7690);
or U13654 (N_13654,N_7536,N_9955);
and U13655 (N_13655,N_9828,N_5390);
nor U13656 (N_13656,N_6666,N_8128);
nand U13657 (N_13657,N_8496,N_6485);
xor U13658 (N_13658,N_6143,N_5702);
or U13659 (N_13659,N_5989,N_6359);
or U13660 (N_13660,N_9952,N_9637);
and U13661 (N_13661,N_9623,N_7723);
nand U13662 (N_13662,N_8134,N_6622);
nand U13663 (N_13663,N_6825,N_5082);
xnor U13664 (N_13664,N_7888,N_8195);
nand U13665 (N_13665,N_8059,N_9064);
xor U13666 (N_13666,N_5017,N_8419);
nor U13667 (N_13667,N_8580,N_7903);
and U13668 (N_13668,N_9774,N_7717);
nand U13669 (N_13669,N_5888,N_6504);
nand U13670 (N_13670,N_8303,N_7672);
nor U13671 (N_13671,N_9959,N_6979);
nand U13672 (N_13672,N_7218,N_5193);
nand U13673 (N_13673,N_6481,N_9578);
and U13674 (N_13674,N_7266,N_6659);
xnor U13675 (N_13675,N_7928,N_7857);
and U13676 (N_13676,N_7391,N_8695);
and U13677 (N_13677,N_8437,N_8766);
and U13678 (N_13678,N_9327,N_7630);
xor U13679 (N_13679,N_7522,N_5132);
nor U13680 (N_13680,N_7258,N_5598);
xor U13681 (N_13681,N_7467,N_9423);
or U13682 (N_13682,N_8151,N_6741);
and U13683 (N_13683,N_6195,N_9038);
or U13684 (N_13684,N_6217,N_9658);
xnor U13685 (N_13685,N_6553,N_6297);
nand U13686 (N_13686,N_7313,N_8390);
xnor U13687 (N_13687,N_9873,N_9164);
nand U13688 (N_13688,N_6990,N_8109);
and U13689 (N_13689,N_5068,N_5552);
nand U13690 (N_13690,N_5358,N_7228);
nor U13691 (N_13691,N_6355,N_7690);
nand U13692 (N_13692,N_6509,N_9181);
xor U13693 (N_13693,N_5934,N_5623);
nand U13694 (N_13694,N_6773,N_6729);
nand U13695 (N_13695,N_7222,N_7752);
xor U13696 (N_13696,N_5385,N_8639);
and U13697 (N_13697,N_9238,N_5085);
or U13698 (N_13698,N_9707,N_9526);
xor U13699 (N_13699,N_7970,N_6547);
or U13700 (N_13700,N_9204,N_8766);
nor U13701 (N_13701,N_8735,N_5677);
nand U13702 (N_13702,N_9361,N_7600);
xnor U13703 (N_13703,N_9833,N_6925);
xor U13704 (N_13704,N_5952,N_7393);
nand U13705 (N_13705,N_7004,N_6021);
or U13706 (N_13706,N_5881,N_9241);
nor U13707 (N_13707,N_6843,N_8280);
and U13708 (N_13708,N_8997,N_9953);
and U13709 (N_13709,N_5317,N_5535);
nand U13710 (N_13710,N_5068,N_6290);
xnor U13711 (N_13711,N_5674,N_7168);
xor U13712 (N_13712,N_7593,N_9214);
nand U13713 (N_13713,N_6423,N_8311);
and U13714 (N_13714,N_6651,N_9692);
or U13715 (N_13715,N_9908,N_6432);
nor U13716 (N_13716,N_5153,N_7128);
nand U13717 (N_13717,N_5847,N_6682);
xnor U13718 (N_13718,N_5263,N_5876);
nor U13719 (N_13719,N_8920,N_8418);
nand U13720 (N_13720,N_5529,N_7240);
nor U13721 (N_13721,N_8903,N_8164);
and U13722 (N_13722,N_8485,N_6523);
nor U13723 (N_13723,N_5273,N_8044);
nand U13724 (N_13724,N_6364,N_7434);
nor U13725 (N_13725,N_7760,N_9836);
or U13726 (N_13726,N_7630,N_7215);
nor U13727 (N_13727,N_8735,N_5961);
xnor U13728 (N_13728,N_7557,N_9271);
nor U13729 (N_13729,N_6927,N_8472);
nor U13730 (N_13730,N_9260,N_7735);
or U13731 (N_13731,N_6071,N_5450);
or U13732 (N_13732,N_5636,N_8257);
xor U13733 (N_13733,N_8739,N_6525);
xnor U13734 (N_13734,N_9485,N_6725);
nor U13735 (N_13735,N_6411,N_8476);
or U13736 (N_13736,N_5972,N_7491);
nor U13737 (N_13737,N_7093,N_8869);
nor U13738 (N_13738,N_8357,N_9423);
nor U13739 (N_13739,N_7225,N_8008);
and U13740 (N_13740,N_5532,N_8114);
nand U13741 (N_13741,N_9438,N_8557);
nor U13742 (N_13742,N_7025,N_9804);
xnor U13743 (N_13743,N_5684,N_5335);
nor U13744 (N_13744,N_9512,N_8200);
nand U13745 (N_13745,N_8570,N_7728);
nand U13746 (N_13746,N_6465,N_5477);
and U13747 (N_13747,N_5981,N_8838);
and U13748 (N_13748,N_8823,N_6205);
or U13749 (N_13749,N_8021,N_7128);
xnor U13750 (N_13750,N_9383,N_8958);
nand U13751 (N_13751,N_7826,N_9605);
or U13752 (N_13752,N_7036,N_7231);
or U13753 (N_13753,N_8724,N_7841);
xor U13754 (N_13754,N_6804,N_7734);
nor U13755 (N_13755,N_8387,N_7298);
and U13756 (N_13756,N_9815,N_7689);
nor U13757 (N_13757,N_5853,N_9981);
nor U13758 (N_13758,N_9776,N_7502);
nor U13759 (N_13759,N_7349,N_8576);
nor U13760 (N_13760,N_7238,N_8752);
nand U13761 (N_13761,N_6627,N_5132);
xor U13762 (N_13762,N_9505,N_5936);
or U13763 (N_13763,N_7817,N_7927);
or U13764 (N_13764,N_6547,N_9582);
or U13765 (N_13765,N_8564,N_9829);
nand U13766 (N_13766,N_5487,N_7055);
or U13767 (N_13767,N_7558,N_5225);
or U13768 (N_13768,N_8221,N_6493);
nor U13769 (N_13769,N_7402,N_7112);
or U13770 (N_13770,N_7136,N_7839);
nand U13771 (N_13771,N_7781,N_6016);
nand U13772 (N_13772,N_5401,N_8935);
xor U13773 (N_13773,N_6314,N_8102);
and U13774 (N_13774,N_6365,N_5249);
or U13775 (N_13775,N_5737,N_7520);
nor U13776 (N_13776,N_5495,N_8459);
or U13777 (N_13777,N_8564,N_6031);
nand U13778 (N_13778,N_7981,N_6780);
nor U13779 (N_13779,N_9930,N_8154);
xor U13780 (N_13780,N_5135,N_7446);
or U13781 (N_13781,N_8709,N_8590);
xor U13782 (N_13782,N_7580,N_9792);
nand U13783 (N_13783,N_8826,N_5133);
and U13784 (N_13784,N_5355,N_5728);
nand U13785 (N_13785,N_6355,N_8919);
nand U13786 (N_13786,N_6705,N_8111);
or U13787 (N_13787,N_9854,N_8507);
nor U13788 (N_13788,N_6194,N_5425);
xnor U13789 (N_13789,N_6796,N_7149);
nand U13790 (N_13790,N_5496,N_9924);
nor U13791 (N_13791,N_5106,N_8781);
nor U13792 (N_13792,N_7308,N_5266);
or U13793 (N_13793,N_9786,N_6511);
or U13794 (N_13794,N_6850,N_5061);
nand U13795 (N_13795,N_8486,N_5903);
nand U13796 (N_13796,N_5697,N_8955);
and U13797 (N_13797,N_9688,N_8595);
or U13798 (N_13798,N_5665,N_5202);
or U13799 (N_13799,N_9612,N_6487);
nand U13800 (N_13800,N_8653,N_6426);
xnor U13801 (N_13801,N_7198,N_9238);
xnor U13802 (N_13802,N_8119,N_7618);
nand U13803 (N_13803,N_6205,N_8155);
or U13804 (N_13804,N_7282,N_6187);
or U13805 (N_13805,N_8787,N_6109);
nand U13806 (N_13806,N_8453,N_7904);
nand U13807 (N_13807,N_9428,N_7110);
nor U13808 (N_13808,N_8936,N_9092);
or U13809 (N_13809,N_5455,N_5971);
nand U13810 (N_13810,N_6433,N_7324);
nor U13811 (N_13811,N_5710,N_9340);
nand U13812 (N_13812,N_8243,N_9952);
and U13813 (N_13813,N_7667,N_9460);
xor U13814 (N_13814,N_5084,N_7704);
nor U13815 (N_13815,N_9737,N_7366);
xor U13816 (N_13816,N_9458,N_9325);
and U13817 (N_13817,N_6034,N_9541);
or U13818 (N_13818,N_5999,N_9364);
nand U13819 (N_13819,N_9545,N_5715);
nand U13820 (N_13820,N_9283,N_9706);
and U13821 (N_13821,N_7486,N_6217);
nand U13822 (N_13822,N_8288,N_7514);
nor U13823 (N_13823,N_6167,N_7368);
nand U13824 (N_13824,N_9463,N_9955);
xnor U13825 (N_13825,N_6273,N_5139);
nand U13826 (N_13826,N_5771,N_9967);
xnor U13827 (N_13827,N_7314,N_5045);
nand U13828 (N_13828,N_8943,N_5969);
and U13829 (N_13829,N_5528,N_5454);
and U13830 (N_13830,N_8434,N_7808);
or U13831 (N_13831,N_6235,N_8975);
xor U13832 (N_13832,N_6967,N_7434);
and U13833 (N_13833,N_9324,N_9820);
and U13834 (N_13834,N_6187,N_7606);
xor U13835 (N_13835,N_9218,N_9225);
xor U13836 (N_13836,N_5195,N_6762);
or U13837 (N_13837,N_7503,N_8849);
nor U13838 (N_13838,N_8228,N_7869);
and U13839 (N_13839,N_9171,N_5379);
nand U13840 (N_13840,N_8028,N_8770);
xnor U13841 (N_13841,N_5791,N_9040);
nand U13842 (N_13842,N_9686,N_9224);
nand U13843 (N_13843,N_9477,N_9257);
or U13844 (N_13844,N_6267,N_9310);
nand U13845 (N_13845,N_5206,N_6194);
xnor U13846 (N_13846,N_7891,N_9626);
and U13847 (N_13847,N_6785,N_9612);
nand U13848 (N_13848,N_8862,N_9709);
xor U13849 (N_13849,N_8809,N_9655);
nand U13850 (N_13850,N_5823,N_7588);
and U13851 (N_13851,N_6333,N_6472);
nand U13852 (N_13852,N_9361,N_8120);
xor U13853 (N_13853,N_7895,N_7437);
xor U13854 (N_13854,N_9215,N_8900);
or U13855 (N_13855,N_8338,N_6628);
nor U13856 (N_13856,N_7660,N_5210);
or U13857 (N_13857,N_7844,N_8686);
or U13858 (N_13858,N_5862,N_8685);
or U13859 (N_13859,N_5585,N_9779);
nand U13860 (N_13860,N_7454,N_9938);
xor U13861 (N_13861,N_7128,N_6272);
or U13862 (N_13862,N_5453,N_5282);
nand U13863 (N_13863,N_7565,N_9451);
nor U13864 (N_13864,N_8570,N_5823);
xnor U13865 (N_13865,N_9824,N_6477);
nor U13866 (N_13866,N_6406,N_6825);
xor U13867 (N_13867,N_5251,N_9332);
nand U13868 (N_13868,N_6397,N_7341);
nor U13869 (N_13869,N_6144,N_8058);
xnor U13870 (N_13870,N_9414,N_9395);
and U13871 (N_13871,N_8803,N_5827);
and U13872 (N_13872,N_8058,N_7983);
or U13873 (N_13873,N_9531,N_9895);
and U13874 (N_13874,N_6418,N_7428);
xnor U13875 (N_13875,N_7904,N_8731);
and U13876 (N_13876,N_6027,N_7148);
nor U13877 (N_13877,N_9390,N_9952);
nand U13878 (N_13878,N_8791,N_8672);
xnor U13879 (N_13879,N_9016,N_9133);
xnor U13880 (N_13880,N_8621,N_5346);
xnor U13881 (N_13881,N_6417,N_6539);
or U13882 (N_13882,N_6454,N_5186);
or U13883 (N_13883,N_8290,N_6925);
xor U13884 (N_13884,N_9342,N_7013);
and U13885 (N_13885,N_6396,N_9360);
xor U13886 (N_13886,N_9052,N_5643);
nor U13887 (N_13887,N_9486,N_6112);
and U13888 (N_13888,N_7695,N_8630);
or U13889 (N_13889,N_6256,N_5207);
nor U13890 (N_13890,N_6797,N_6842);
xnor U13891 (N_13891,N_6259,N_8909);
and U13892 (N_13892,N_9997,N_6588);
nor U13893 (N_13893,N_8015,N_7392);
or U13894 (N_13894,N_5378,N_7758);
and U13895 (N_13895,N_7476,N_9686);
and U13896 (N_13896,N_7940,N_9419);
or U13897 (N_13897,N_8170,N_6155);
nand U13898 (N_13898,N_6719,N_8724);
nor U13899 (N_13899,N_9254,N_5125);
nor U13900 (N_13900,N_6446,N_6214);
nor U13901 (N_13901,N_7613,N_6914);
nor U13902 (N_13902,N_7174,N_6427);
nand U13903 (N_13903,N_8333,N_5833);
or U13904 (N_13904,N_8098,N_5077);
nand U13905 (N_13905,N_5767,N_6124);
or U13906 (N_13906,N_6005,N_9018);
nand U13907 (N_13907,N_9869,N_5512);
or U13908 (N_13908,N_5844,N_5318);
or U13909 (N_13909,N_6589,N_8127);
and U13910 (N_13910,N_5799,N_8912);
nor U13911 (N_13911,N_5682,N_9085);
xor U13912 (N_13912,N_5375,N_7546);
nor U13913 (N_13913,N_6924,N_9685);
and U13914 (N_13914,N_9517,N_9498);
nand U13915 (N_13915,N_6606,N_9891);
nor U13916 (N_13916,N_9586,N_8830);
or U13917 (N_13917,N_6861,N_7614);
nor U13918 (N_13918,N_7977,N_7486);
nor U13919 (N_13919,N_7107,N_8458);
xnor U13920 (N_13920,N_8008,N_6872);
nor U13921 (N_13921,N_7427,N_8370);
nand U13922 (N_13922,N_8901,N_9467);
and U13923 (N_13923,N_5537,N_9967);
nor U13924 (N_13924,N_9261,N_9697);
or U13925 (N_13925,N_9666,N_6367);
nor U13926 (N_13926,N_6244,N_6981);
xnor U13927 (N_13927,N_6074,N_9312);
nand U13928 (N_13928,N_8900,N_6511);
and U13929 (N_13929,N_9313,N_6465);
nand U13930 (N_13930,N_9435,N_9833);
and U13931 (N_13931,N_5650,N_8302);
nor U13932 (N_13932,N_9228,N_5713);
or U13933 (N_13933,N_5925,N_8786);
nor U13934 (N_13934,N_9359,N_8352);
nor U13935 (N_13935,N_5007,N_5941);
xor U13936 (N_13936,N_5750,N_9333);
nor U13937 (N_13937,N_7643,N_5378);
nor U13938 (N_13938,N_5005,N_7161);
xor U13939 (N_13939,N_9649,N_9333);
and U13940 (N_13940,N_8607,N_7968);
and U13941 (N_13941,N_8984,N_6946);
xor U13942 (N_13942,N_8826,N_5686);
xor U13943 (N_13943,N_7184,N_6534);
xor U13944 (N_13944,N_6028,N_8679);
nor U13945 (N_13945,N_5507,N_6767);
or U13946 (N_13946,N_6110,N_8305);
or U13947 (N_13947,N_8845,N_5036);
nand U13948 (N_13948,N_6298,N_9160);
nor U13949 (N_13949,N_9888,N_8344);
or U13950 (N_13950,N_6124,N_5624);
nor U13951 (N_13951,N_5101,N_6364);
nand U13952 (N_13952,N_5988,N_7509);
xor U13953 (N_13953,N_6054,N_8249);
xnor U13954 (N_13954,N_8859,N_5070);
or U13955 (N_13955,N_8805,N_9285);
nor U13956 (N_13956,N_5740,N_5924);
or U13957 (N_13957,N_5415,N_9561);
or U13958 (N_13958,N_7922,N_5128);
nand U13959 (N_13959,N_8035,N_6195);
nand U13960 (N_13960,N_9907,N_9373);
or U13961 (N_13961,N_8378,N_9352);
xnor U13962 (N_13962,N_5539,N_7882);
nor U13963 (N_13963,N_7807,N_6753);
nand U13964 (N_13964,N_5176,N_5474);
nor U13965 (N_13965,N_5875,N_8144);
or U13966 (N_13966,N_9868,N_7454);
or U13967 (N_13967,N_5931,N_7841);
or U13968 (N_13968,N_8794,N_7178);
xor U13969 (N_13969,N_9030,N_7614);
nor U13970 (N_13970,N_9493,N_8518);
or U13971 (N_13971,N_7003,N_5774);
and U13972 (N_13972,N_5112,N_5927);
xnor U13973 (N_13973,N_6076,N_9434);
and U13974 (N_13974,N_9664,N_8486);
xor U13975 (N_13975,N_5255,N_7429);
nor U13976 (N_13976,N_5620,N_9863);
or U13977 (N_13977,N_6173,N_7717);
nor U13978 (N_13978,N_7450,N_7806);
xor U13979 (N_13979,N_7646,N_9775);
or U13980 (N_13980,N_6966,N_8038);
xnor U13981 (N_13981,N_9523,N_7166);
and U13982 (N_13982,N_6323,N_6056);
and U13983 (N_13983,N_9861,N_8418);
or U13984 (N_13984,N_8112,N_9890);
xor U13985 (N_13985,N_7132,N_9495);
nand U13986 (N_13986,N_9214,N_7344);
or U13987 (N_13987,N_9597,N_8883);
nor U13988 (N_13988,N_5869,N_9502);
nor U13989 (N_13989,N_7383,N_7542);
nand U13990 (N_13990,N_8584,N_7529);
xnor U13991 (N_13991,N_5484,N_6955);
or U13992 (N_13992,N_9758,N_5986);
and U13993 (N_13993,N_6837,N_5894);
and U13994 (N_13994,N_9944,N_7924);
or U13995 (N_13995,N_7732,N_8549);
and U13996 (N_13996,N_9107,N_8011);
or U13997 (N_13997,N_6431,N_5815);
nor U13998 (N_13998,N_8107,N_8336);
nand U13999 (N_13999,N_7515,N_8804);
and U14000 (N_14000,N_8218,N_8219);
or U14001 (N_14001,N_8908,N_5776);
or U14002 (N_14002,N_9261,N_7901);
nand U14003 (N_14003,N_5952,N_9965);
or U14004 (N_14004,N_6730,N_5735);
nor U14005 (N_14005,N_8001,N_9361);
and U14006 (N_14006,N_7381,N_5000);
xnor U14007 (N_14007,N_6086,N_9550);
or U14008 (N_14008,N_5161,N_9334);
xnor U14009 (N_14009,N_9987,N_7112);
and U14010 (N_14010,N_9779,N_5792);
or U14011 (N_14011,N_5339,N_5273);
xnor U14012 (N_14012,N_8628,N_5411);
or U14013 (N_14013,N_5166,N_5636);
nor U14014 (N_14014,N_9556,N_9727);
or U14015 (N_14015,N_9647,N_8229);
nand U14016 (N_14016,N_8292,N_6621);
or U14017 (N_14017,N_6916,N_8968);
nor U14018 (N_14018,N_9221,N_6824);
nor U14019 (N_14019,N_7272,N_5190);
and U14020 (N_14020,N_8590,N_7676);
or U14021 (N_14021,N_5936,N_5388);
nor U14022 (N_14022,N_7823,N_5783);
or U14023 (N_14023,N_9727,N_6739);
nor U14024 (N_14024,N_9381,N_5734);
nand U14025 (N_14025,N_7392,N_5896);
nor U14026 (N_14026,N_8431,N_6502);
xnor U14027 (N_14027,N_8369,N_7248);
nand U14028 (N_14028,N_8932,N_8169);
xnor U14029 (N_14029,N_8564,N_7251);
nor U14030 (N_14030,N_9776,N_8230);
and U14031 (N_14031,N_6001,N_5299);
nand U14032 (N_14032,N_6531,N_5564);
or U14033 (N_14033,N_5482,N_7757);
xor U14034 (N_14034,N_5086,N_5094);
or U14035 (N_14035,N_9812,N_9330);
nand U14036 (N_14036,N_5095,N_5264);
nand U14037 (N_14037,N_5233,N_6902);
nor U14038 (N_14038,N_5763,N_6408);
nor U14039 (N_14039,N_9437,N_9249);
nor U14040 (N_14040,N_6154,N_7550);
nand U14041 (N_14041,N_7665,N_7582);
and U14042 (N_14042,N_9159,N_5348);
and U14043 (N_14043,N_5367,N_5504);
nor U14044 (N_14044,N_6641,N_5945);
xor U14045 (N_14045,N_9369,N_7049);
xor U14046 (N_14046,N_5614,N_9132);
nand U14047 (N_14047,N_6793,N_5312);
nor U14048 (N_14048,N_8726,N_5889);
xnor U14049 (N_14049,N_9663,N_9595);
nor U14050 (N_14050,N_5237,N_7789);
nor U14051 (N_14051,N_7466,N_6372);
nand U14052 (N_14052,N_9275,N_6100);
nand U14053 (N_14053,N_7329,N_5605);
nor U14054 (N_14054,N_5376,N_8799);
and U14055 (N_14055,N_7546,N_7976);
or U14056 (N_14056,N_6607,N_5591);
or U14057 (N_14057,N_6905,N_6397);
nand U14058 (N_14058,N_9916,N_7923);
or U14059 (N_14059,N_7133,N_8106);
xnor U14060 (N_14060,N_8844,N_9616);
nor U14061 (N_14061,N_5593,N_9633);
nor U14062 (N_14062,N_7786,N_8806);
or U14063 (N_14063,N_8948,N_6858);
nand U14064 (N_14064,N_8348,N_6252);
nand U14065 (N_14065,N_5636,N_9196);
and U14066 (N_14066,N_5655,N_7871);
and U14067 (N_14067,N_7217,N_5123);
xnor U14068 (N_14068,N_7024,N_8570);
nor U14069 (N_14069,N_8782,N_5019);
or U14070 (N_14070,N_9877,N_6477);
and U14071 (N_14071,N_9264,N_8039);
nand U14072 (N_14072,N_5271,N_9826);
and U14073 (N_14073,N_5361,N_7930);
xnor U14074 (N_14074,N_5318,N_8462);
and U14075 (N_14075,N_8385,N_5766);
xor U14076 (N_14076,N_7331,N_5957);
nor U14077 (N_14077,N_5413,N_5982);
xor U14078 (N_14078,N_5282,N_6332);
and U14079 (N_14079,N_6235,N_8087);
xnor U14080 (N_14080,N_9649,N_9458);
nor U14081 (N_14081,N_5231,N_7183);
or U14082 (N_14082,N_8573,N_8575);
nor U14083 (N_14083,N_7665,N_9994);
and U14084 (N_14084,N_6616,N_9053);
xnor U14085 (N_14085,N_9175,N_8091);
or U14086 (N_14086,N_8836,N_5587);
nor U14087 (N_14087,N_5049,N_9623);
and U14088 (N_14088,N_9103,N_6943);
nand U14089 (N_14089,N_9338,N_6851);
and U14090 (N_14090,N_7855,N_9255);
and U14091 (N_14091,N_5730,N_7672);
and U14092 (N_14092,N_5463,N_7885);
nand U14093 (N_14093,N_6894,N_6459);
nand U14094 (N_14094,N_8943,N_7880);
or U14095 (N_14095,N_8962,N_5366);
xor U14096 (N_14096,N_7337,N_7003);
xor U14097 (N_14097,N_6290,N_5699);
and U14098 (N_14098,N_7809,N_8009);
or U14099 (N_14099,N_9173,N_8142);
and U14100 (N_14100,N_8879,N_5237);
nand U14101 (N_14101,N_7760,N_6748);
nand U14102 (N_14102,N_6158,N_8566);
xor U14103 (N_14103,N_9334,N_5638);
and U14104 (N_14104,N_5846,N_6350);
nor U14105 (N_14105,N_9776,N_7567);
or U14106 (N_14106,N_9751,N_5621);
or U14107 (N_14107,N_6588,N_8934);
xnor U14108 (N_14108,N_6036,N_9834);
and U14109 (N_14109,N_5044,N_8614);
or U14110 (N_14110,N_8179,N_6019);
or U14111 (N_14111,N_8987,N_8272);
and U14112 (N_14112,N_8654,N_5546);
xnor U14113 (N_14113,N_7130,N_5371);
or U14114 (N_14114,N_9356,N_5131);
nor U14115 (N_14115,N_7007,N_9037);
or U14116 (N_14116,N_7096,N_5424);
or U14117 (N_14117,N_9362,N_5052);
or U14118 (N_14118,N_9050,N_9769);
or U14119 (N_14119,N_9683,N_8829);
nor U14120 (N_14120,N_8033,N_8303);
nor U14121 (N_14121,N_8849,N_6494);
or U14122 (N_14122,N_8407,N_8303);
nand U14123 (N_14123,N_8674,N_8986);
nor U14124 (N_14124,N_6478,N_8357);
nand U14125 (N_14125,N_9420,N_9268);
nor U14126 (N_14126,N_5656,N_8443);
nand U14127 (N_14127,N_9500,N_7358);
xnor U14128 (N_14128,N_9387,N_9345);
nor U14129 (N_14129,N_7532,N_6816);
or U14130 (N_14130,N_5268,N_9420);
and U14131 (N_14131,N_6196,N_9830);
and U14132 (N_14132,N_6742,N_7210);
or U14133 (N_14133,N_6510,N_9885);
and U14134 (N_14134,N_8858,N_7963);
and U14135 (N_14135,N_8209,N_5416);
xor U14136 (N_14136,N_8402,N_8730);
xnor U14137 (N_14137,N_8354,N_8458);
and U14138 (N_14138,N_7539,N_7226);
nor U14139 (N_14139,N_7311,N_8959);
nor U14140 (N_14140,N_5302,N_5702);
nor U14141 (N_14141,N_7483,N_8090);
xnor U14142 (N_14142,N_8262,N_8102);
nor U14143 (N_14143,N_8217,N_9001);
xor U14144 (N_14144,N_6586,N_7319);
nor U14145 (N_14145,N_8037,N_8126);
nor U14146 (N_14146,N_6921,N_5415);
xnor U14147 (N_14147,N_7818,N_5255);
and U14148 (N_14148,N_7143,N_6712);
or U14149 (N_14149,N_5893,N_9504);
nand U14150 (N_14150,N_5978,N_7441);
and U14151 (N_14151,N_7874,N_5399);
nand U14152 (N_14152,N_6375,N_5376);
xor U14153 (N_14153,N_7806,N_6784);
nand U14154 (N_14154,N_8265,N_7226);
xor U14155 (N_14155,N_5586,N_8278);
or U14156 (N_14156,N_5613,N_6405);
nor U14157 (N_14157,N_6996,N_7074);
nand U14158 (N_14158,N_8256,N_5146);
xnor U14159 (N_14159,N_7441,N_8587);
nand U14160 (N_14160,N_6456,N_5459);
or U14161 (N_14161,N_6624,N_8602);
xnor U14162 (N_14162,N_9504,N_5247);
xnor U14163 (N_14163,N_6954,N_7624);
or U14164 (N_14164,N_6372,N_7573);
nor U14165 (N_14165,N_6628,N_6068);
nor U14166 (N_14166,N_5439,N_9071);
and U14167 (N_14167,N_9976,N_5905);
or U14168 (N_14168,N_9178,N_5069);
nand U14169 (N_14169,N_5158,N_8046);
nor U14170 (N_14170,N_6530,N_8016);
nand U14171 (N_14171,N_6152,N_8110);
nand U14172 (N_14172,N_6035,N_7960);
xor U14173 (N_14173,N_6023,N_7448);
or U14174 (N_14174,N_9947,N_6004);
or U14175 (N_14175,N_8323,N_8828);
and U14176 (N_14176,N_5818,N_9281);
and U14177 (N_14177,N_9958,N_8625);
nand U14178 (N_14178,N_9945,N_9440);
and U14179 (N_14179,N_5712,N_8030);
nand U14180 (N_14180,N_9384,N_6558);
or U14181 (N_14181,N_5066,N_8740);
xnor U14182 (N_14182,N_5448,N_6021);
nor U14183 (N_14183,N_7902,N_8823);
xor U14184 (N_14184,N_9432,N_8069);
nor U14185 (N_14185,N_9251,N_8824);
xor U14186 (N_14186,N_8732,N_7647);
nand U14187 (N_14187,N_7968,N_8885);
or U14188 (N_14188,N_8850,N_8043);
or U14189 (N_14189,N_6827,N_9659);
nor U14190 (N_14190,N_6957,N_7384);
xor U14191 (N_14191,N_6440,N_9299);
and U14192 (N_14192,N_5577,N_9423);
nand U14193 (N_14193,N_8497,N_7722);
or U14194 (N_14194,N_9303,N_5852);
and U14195 (N_14195,N_6705,N_7779);
xnor U14196 (N_14196,N_5286,N_6605);
xnor U14197 (N_14197,N_7975,N_9893);
xnor U14198 (N_14198,N_6266,N_5801);
xnor U14199 (N_14199,N_8845,N_5465);
or U14200 (N_14200,N_8911,N_9834);
or U14201 (N_14201,N_8920,N_7092);
nor U14202 (N_14202,N_5874,N_7839);
or U14203 (N_14203,N_8842,N_5366);
nand U14204 (N_14204,N_8266,N_7288);
or U14205 (N_14205,N_9137,N_8786);
and U14206 (N_14206,N_6835,N_6235);
nand U14207 (N_14207,N_9213,N_7892);
nand U14208 (N_14208,N_7404,N_8140);
nand U14209 (N_14209,N_7213,N_6195);
or U14210 (N_14210,N_7704,N_7539);
and U14211 (N_14211,N_6846,N_9067);
or U14212 (N_14212,N_7737,N_5558);
xor U14213 (N_14213,N_8501,N_7138);
xnor U14214 (N_14214,N_9447,N_8161);
nor U14215 (N_14215,N_5812,N_7087);
or U14216 (N_14216,N_9985,N_6092);
nor U14217 (N_14217,N_7592,N_5898);
xor U14218 (N_14218,N_9178,N_6419);
nand U14219 (N_14219,N_9750,N_7843);
and U14220 (N_14220,N_8626,N_5845);
nand U14221 (N_14221,N_6452,N_9994);
and U14222 (N_14222,N_8664,N_7020);
nand U14223 (N_14223,N_8786,N_8288);
xor U14224 (N_14224,N_6215,N_9945);
and U14225 (N_14225,N_5556,N_7599);
xor U14226 (N_14226,N_8471,N_6506);
nor U14227 (N_14227,N_5421,N_5100);
and U14228 (N_14228,N_9836,N_6368);
or U14229 (N_14229,N_7358,N_9810);
nand U14230 (N_14230,N_9720,N_9311);
nor U14231 (N_14231,N_7654,N_9350);
nor U14232 (N_14232,N_8226,N_5866);
and U14233 (N_14233,N_7581,N_9648);
or U14234 (N_14234,N_9933,N_8441);
or U14235 (N_14235,N_5019,N_7961);
nor U14236 (N_14236,N_5446,N_5594);
nand U14237 (N_14237,N_7499,N_5966);
nor U14238 (N_14238,N_6362,N_7037);
and U14239 (N_14239,N_9576,N_9503);
and U14240 (N_14240,N_7038,N_6387);
or U14241 (N_14241,N_6089,N_7316);
nor U14242 (N_14242,N_7604,N_9530);
xnor U14243 (N_14243,N_8834,N_5093);
and U14244 (N_14244,N_8944,N_5858);
and U14245 (N_14245,N_7451,N_7496);
or U14246 (N_14246,N_6553,N_7549);
xnor U14247 (N_14247,N_8652,N_9550);
xnor U14248 (N_14248,N_7468,N_8288);
nor U14249 (N_14249,N_8866,N_8535);
nor U14250 (N_14250,N_7121,N_5085);
nand U14251 (N_14251,N_9056,N_9762);
or U14252 (N_14252,N_7448,N_8200);
or U14253 (N_14253,N_5468,N_5760);
nor U14254 (N_14254,N_8553,N_9705);
xor U14255 (N_14255,N_6642,N_5534);
and U14256 (N_14256,N_5217,N_8395);
xnor U14257 (N_14257,N_6963,N_9460);
and U14258 (N_14258,N_5828,N_9071);
and U14259 (N_14259,N_9894,N_5360);
nand U14260 (N_14260,N_5882,N_9124);
or U14261 (N_14261,N_8626,N_7154);
xnor U14262 (N_14262,N_6714,N_7152);
or U14263 (N_14263,N_7514,N_5420);
or U14264 (N_14264,N_6932,N_7950);
nor U14265 (N_14265,N_8338,N_6970);
xnor U14266 (N_14266,N_5058,N_7751);
nand U14267 (N_14267,N_9459,N_9485);
and U14268 (N_14268,N_7393,N_5826);
or U14269 (N_14269,N_6950,N_7302);
or U14270 (N_14270,N_9720,N_9479);
nor U14271 (N_14271,N_6652,N_5211);
and U14272 (N_14272,N_5385,N_8716);
nor U14273 (N_14273,N_7455,N_5093);
or U14274 (N_14274,N_6554,N_8911);
or U14275 (N_14275,N_9872,N_5559);
nor U14276 (N_14276,N_7230,N_5501);
or U14277 (N_14277,N_9594,N_5877);
nor U14278 (N_14278,N_5494,N_8707);
xnor U14279 (N_14279,N_5796,N_7465);
nor U14280 (N_14280,N_6351,N_6908);
or U14281 (N_14281,N_5177,N_6238);
xnor U14282 (N_14282,N_6373,N_6591);
or U14283 (N_14283,N_6479,N_9727);
nand U14284 (N_14284,N_7046,N_7074);
and U14285 (N_14285,N_5329,N_8485);
and U14286 (N_14286,N_8036,N_8984);
and U14287 (N_14287,N_5533,N_9250);
nor U14288 (N_14288,N_8820,N_7317);
nand U14289 (N_14289,N_8677,N_6921);
xnor U14290 (N_14290,N_7076,N_9188);
xnor U14291 (N_14291,N_8334,N_7078);
xor U14292 (N_14292,N_6615,N_6960);
nor U14293 (N_14293,N_5296,N_7516);
xnor U14294 (N_14294,N_9509,N_5570);
or U14295 (N_14295,N_5361,N_5970);
nand U14296 (N_14296,N_8273,N_9142);
nor U14297 (N_14297,N_6056,N_7693);
nand U14298 (N_14298,N_5442,N_6676);
nand U14299 (N_14299,N_7833,N_9735);
xor U14300 (N_14300,N_5754,N_9618);
xor U14301 (N_14301,N_9731,N_6590);
and U14302 (N_14302,N_8866,N_7243);
and U14303 (N_14303,N_7673,N_7514);
and U14304 (N_14304,N_8655,N_5360);
or U14305 (N_14305,N_5120,N_9119);
or U14306 (N_14306,N_5358,N_6485);
nand U14307 (N_14307,N_5568,N_7642);
nor U14308 (N_14308,N_9292,N_7071);
and U14309 (N_14309,N_7420,N_7063);
nand U14310 (N_14310,N_9903,N_6472);
xor U14311 (N_14311,N_8314,N_6875);
xnor U14312 (N_14312,N_8063,N_8547);
nor U14313 (N_14313,N_9547,N_7398);
nand U14314 (N_14314,N_6391,N_8362);
nand U14315 (N_14315,N_9731,N_7796);
nor U14316 (N_14316,N_9804,N_7640);
or U14317 (N_14317,N_9220,N_9229);
or U14318 (N_14318,N_9606,N_8631);
nand U14319 (N_14319,N_8442,N_6064);
and U14320 (N_14320,N_9985,N_6053);
and U14321 (N_14321,N_6218,N_8184);
xnor U14322 (N_14322,N_9464,N_9788);
nand U14323 (N_14323,N_8082,N_8202);
nor U14324 (N_14324,N_5333,N_6361);
xnor U14325 (N_14325,N_6866,N_9168);
or U14326 (N_14326,N_6551,N_9113);
nand U14327 (N_14327,N_9356,N_7839);
and U14328 (N_14328,N_6814,N_5775);
nor U14329 (N_14329,N_5295,N_5567);
nand U14330 (N_14330,N_6941,N_5276);
nand U14331 (N_14331,N_7407,N_6371);
or U14332 (N_14332,N_7835,N_5737);
xor U14333 (N_14333,N_7233,N_8069);
and U14334 (N_14334,N_8836,N_5912);
nand U14335 (N_14335,N_8947,N_6192);
nand U14336 (N_14336,N_7792,N_6956);
nor U14337 (N_14337,N_7966,N_5400);
xnor U14338 (N_14338,N_6415,N_9934);
nor U14339 (N_14339,N_8840,N_6522);
xnor U14340 (N_14340,N_5254,N_6009);
or U14341 (N_14341,N_6991,N_8603);
nor U14342 (N_14342,N_6502,N_8994);
nand U14343 (N_14343,N_6692,N_6764);
nor U14344 (N_14344,N_6779,N_6522);
nor U14345 (N_14345,N_5893,N_8426);
nand U14346 (N_14346,N_8283,N_6092);
or U14347 (N_14347,N_6048,N_9175);
nand U14348 (N_14348,N_8919,N_6587);
nand U14349 (N_14349,N_9299,N_7894);
nor U14350 (N_14350,N_6249,N_5869);
or U14351 (N_14351,N_6494,N_6138);
and U14352 (N_14352,N_5958,N_7767);
nand U14353 (N_14353,N_7800,N_7355);
nor U14354 (N_14354,N_9259,N_7756);
or U14355 (N_14355,N_8370,N_5651);
xnor U14356 (N_14356,N_6272,N_6632);
nor U14357 (N_14357,N_9791,N_6275);
and U14358 (N_14358,N_6998,N_9956);
or U14359 (N_14359,N_5184,N_8824);
or U14360 (N_14360,N_8768,N_5870);
xor U14361 (N_14361,N_6870,N_8303);
nor U14362 (N_14362,N_5656,N_7406);
nor U14363 (N_14363,N_9357,N_7865);
nand U14364 (N_14364,N_8742,N_9644);
or U14365 (N_14365,N_7405,N_5325);
nand U14366 (N_14366,N_7855,N_7846);
or U14367 (N_14367,N_6584,N_9080);
and U14368 (N_14368,N_6395,N_6267);
nand U14369 (N_14369,N_7165,N_5168);
nor U14370 (N_14370,N_8467,N_6497);
nor U14371 (N_14371,N_7253,N_7833);
or U14372 (N_14372,N_8267,N_5760);
nand U14373 (N_14373,N_6045,N_6971);
and U14374 (N_14374,N_5399,N_5423);
xnor U14375 (N_14375,N_5280,N_6797);
nor U14376 (N_14376,N_8998,N_5425);
and U14377 (N_14377,N_6147,N_5152);
xor U14378 (N_14378,N_9868,N_5466);
or U14379 (N_14379,N_6842,N_9973);
nor U14380 (N_14380,N_9310,N_6268);
nor U14381 (N_14381,N_5774,N_7513);
nor U14382 (N_14382,N_8421,N_6353);
nor U14383 (N_14383,N_8258,N_8166);
xor U14384 (N_14384,N_6232,N_6716);
or U14385 (N_14385,N_8445,N_6585);
or U14386 (N_14386,N_8696,N_9133);
and U14387 (N_14387,N_8148,N_7671);
nand U14388 (N_14388,N_9281,N_7203);
or U14389 (N_14389,N_8695,N_8791);
or U14390 (N_14390,N_6486,N_7117);
nor U14391 (N_14391,N_5573,N_5389);
and U14392 (N_14392,N_6043,N_7659);
xor U14393 (N_14393,N_9318,N_6721);
and U14394 (N_14394,N_7292,N_5279);
xor U14395 (N_14395,N_5703,N_8345);
or U14396 (N_14396,N_6169,N_6002);
xor U14397 (N_14397,N_8465,N_7633);
or U14398 (N_14398,N_5240,N_5912);
nor U14399 (N_14399,N_5158,N_9761);
nor U14400 (N_14400,N_9631,N_6304);
nand U14401 (N_14401,N_8361,N_8944);
xor U14402 (N_14402,N_5841,N_8233);
nor U14403 (N_14403,N_8381,N_8477);
xor U14404 (N_14404,N_8190,N_6310);
or U14405 (N_14405,N_7050,N_5828);
xnor U14406 (N_14406,N_8014,N_6119);
nand U14407 (N_14407,N_9413,N_6925);
xor U14408 (N_14408,N_5558,N_7562);
nor U14409 (N_14409,N_6968,N_9637);
xor U14410 (N_14410,N_8635,N_9110);
nor U14411 (N_14411,N_8223,N_8653);
nor U14412 (N_14412,N_8198,N_8640);
and U14413 (N_14413,N_5148,N_6462);
and U14414 (N_14414,N_7902,N_9418);
xnor U14415 (N_14415,N_7655,N_6993);
or U14416 (N_14416,N_8131,N_8164);
nand U14417 (N_14417,N_8026,N_7007);
and U14418 (N_14418,N_9467,N_6818);
or U14419 (N_14419,N_5900,N_6720);
nand U14420 (N_14420,N_6972,N_9827);
nand U14421 (N_14421,N_7161,N_9242);
xor U14422 (N_14422,N_7277,N_9020);
nand U14423 (N_14423,N_8612,N_5433);
nor U14424 (N_14424,N_8123,N_7630);
nand U14425 (N_14425,N_5118,N_6530);
nor U14426 (N_14426,N_9970,N_6090);
and U14427 (N_14427,N_9710,N_8099);
nor U14428 (N_14428,N_6982,N_9298);
or U14429 (N_14429,N_7934,N_8411);
xnor U14430 (N_14430,N_5330,N_6258);
or U14431 (N_14431,N_6569,N_8796);
nand U14432 (N_14432,N_6521,N_9002);
nor U14433 (N_14433,N_7424,N_8827);
and U14434 (N_14434,N_6698,N_6976);
nand U14435 (N_14435,N_7676,N_6037);
and U14436 (N_14436,N_9234,N_7599);
or U14437 (N_14437,N_5513,N_8666);
nand U14438 (N_14438,N_9497,N_7969);
and U14439 (N_14439,N_7243,N_8125);
xnor U14440 (N_14440,N_9289,N_6096);
and U14441 (N_14441,N_5575,N_7119);
nor U14442 (N_14442,N_9371,N_9613);
nand U14443 (N_14443,N_7891,N_6761);
and U14444 (N_14444,N_8298,N_6014);
xor U14445 (N_14445,N_6118,N_6848);
nor U14446 (N_14446,N_5187,N_8920);
and U14447 (N_14447,N_7773,N_6806);
or U14448 (N_14448,N_7180,N_5409);
xor U14449 (N_14449,N_7152,N_7970);
and U14450 (N_14450,N_6944,N_6351);
or U14451 (N_14451,N_7178,N_7329);
xnor U14452 (N_14452,N_7556,N_9413);
and U14453 (N_14453,N_8344,N_8730);
nor U14454 (N_14454,N_8228,N_7653);
and U14455 (N_14455,N_5989,N_8074);
xnor U14456 (N_14456,N_5639,N_9815);
xnor U14457 (N_14457,N_8977,N_9709);
or U14458 (N_14458,N_9962,N_7620);
nor U14459 (N_14459,N_5284,N_5338);
nand U14460 (N_14460,N_7279,N_7336);
and U14461 (N_14461,N_9505,N_7147);
or U14462 (N_14462,N_6581,N_5658);
or U14463 (N_14463,N_5252,N_8407);
nor U14464 (N_14464,N_7526,N_8781);
xnor U14465 (N_14465,N_5494,N_7658);
nor U14466 (N_14466,N_9357,N_9929);
and U14467 (N_14467,N_5448,N_9286);
nand U14468 (N_14468,N_7673,N_7920);
nand U14469 (N_14469,N_5175,N_6501);
nand U14470 (N_14470,N_5217,N_6580);
xnor U14471 (N_14471,N_6282,N_7254);
nand U14472 (N_14472,N_7512,N_9795);
nor U14473 (N_14473,N_5791,N_5602);
nor U14474 (N_14474,N_9674,N_6769);
xnor U14475 (N_14475,N_5606,N_8975);
nor U14476 (N_14476,N_7057,N_5039);
nand U14477 (N_14477,N_8471,N_5305);
or U14478 (N_14478,N_7558,N_6837);
or U14479 (N_14479,N_8863,N_8374);
nor U14480 (N_14480,N_7480,N_8857);
xnor U14481 (N_14481,N_8618,N_7745);
or U14482 (N_14482,N_8373,N_8932);
xor U14483 (N_14483,N_8297,N_9207);
or U14484 (N_14484,N_5244,N_6046);
or U14485 (N_14485,N_9925,N_9823);
xor U14486 (N_14486,N_7410,N_8578);
nand U14487 (N_14487,N_6158,N_5824);
or U14488 (N_14488,N_6099,N_6064);
and U14489 (N_14489,N_5957,N_9988);
or U14490 (N_14490,N_9863,N_7473);
and U14491 (N_14491,N_5221,N_7135);
or U14492 (N_14492,N_7240,N_6541);
or U14493 (N_14493,N_5105,N_7173);
and U14494 (N_14494,N_6478,N_5428);
xor U14495 (N_14495,N_5311,N_5166);
nand U14496 (N_14496,N_5573,N_5030);
nand U14497 (N_14497,N_5055,N_8433);
or U14498 (N_14498,N_6487,N_5722);
nor U14499 (N_14499,N_6570,N_5098);
or U14500 (N_14500,N_6746,N_8492);
nor U14501 (N_14501,N_6992,N_5462);
and U14502 (N_14502,N_7206,N_9214);
xor U14503 (N_14503,N_9217,N_5826);
nor U14504 (N_14504,N_7273,N_6008);
or U14505 (N_14505,N_5879,N_5082);
nor U14506 (N_14506,N_6277,N_8168);
and U14507 (N_14507,N_8726,N_9335);
xor U14508 (N_14508,N_7702,N_8577);
nand U14509 (N_14509,N_8070,N_7553);
xnor U14510 (N_14510,N_5478,N_9819);
or U14511 (N_14511,N_7308,N_9766);
xnor U14512 (N_14512,N_5628,N_9000);
and U14513 (N_14513,N_6911,N_7286);
or U14514 (N_14514,N_9586,N_7500);
xor U14515 (N_14515,N_9374,N_8163);
and U14516 (N_14516,N_6701,N_8142);
nand U14517 (N_14517,N_8875,N_6978);
and U14518 (N_14518,N_8886,N_7407);
and U14519 (N_14519,N_7788,N_9534);
nand U14520 (N_14520,N_7715,N_8429);
nand U14521 (N_14521,N_7281,N_8206);
xnor U14522 (N_14522,N_8479,N_5435);
nor U14523 (N_14523,N_8984,N_5453);
nand U14524 (N_14524,N_6805,N_8830);
or U14525 (N_14525,N_7100,N_9812);
and U14526 (N_14526,N_8636,N_8993);
or U14527 (N_14527,N_9623,N_5846);
xor U14528 (N_14528,N_8070,N_6651);
or U14529 (N_14529,N_7099,N_8788);
or U14530 (N_14530,N_7718,N_5289);
and U14531 (N_14531,N_8353,N_7305);
nor U14532 (N_14532,N_6423,N_6516);
nand U14533 (N_14533,N_6462,N_6656);
and U14534 (N_14534,N_7875,N_7078);
and U14535 (N_14535,N_5975,N_9165);
nor U14536 (N_14536,N_7006,N_7389);
nor U14537 (N_14537,N_5221,N_7231);
and U14538 (N_14538,N_6700,N_5563);
xnor U14539 (N_14539,N_9507,N_8839);
and U14540 (N_14540,N_5242,N_7622);
nor U14541 (N_14541,N_6767,N_5789);
nor U14542 (N_14542,N_7249,N_8628);
or U14543 (N_14543,N_8527,N_8973);
nand U14544 (N_14544,N_5117,N_6626);
or U14545 (N_14545,N_6853,N_7563);
nand U14546 (N_14546,N_6817,N_8112);
nor U14547 (N_14547,N_6783,N_6809);
xnor U14548 (N_14548,N_9973,N_7142);
or U14549 (N_14549,N_7554,N_5919);
and U14550 (N_14550,N_7782,N_7000);
and U14551 (N_14551,N_8923,N_7143);
or U14552 (N_14552,N_8659,N_9106);
nand U14553 (N_14553,N_5780,N_9226);
and U14554 (N_14554,N_5580,N_5661);
xor U14555 (N_14555,N_5832,N_7150);
and U14556 (N_14556,N_8982,N_7872);
nor U14557 (N_14557,N_9615,N_9477);
and U14558 (N_14558,N_7611,N_6853);
and U14559 (N_14559,N_5253,N_8863);
xnor U14560 (N_14560,N_8505,N_9440);
nand U14561 (N_14561,N_8191,N_5728);
xnor U14562 (N_14562,N_8645,N_5000);
xnor U14563 (N_14563,N_6782,N_7877);
or U14564 (N_14564,N_6080,N_7063);
nor U14565 (N_14565,N_8665,N_6507);
nand U14566 (N_14566,N_8169,N_5671);
nor U14567 (N_14567,N_6682,N_9783);
or U14568 (N_14568,N_7279,N_5407);
or U14569 (N_14569,N_9975,N_9261);
nor U14570 (N_14570,N_6946,N_6815);
xor U14571 (N_14571,N_8095,N_9838);
xnor U14572 (N_14572,N_8097,N_7506);
and U14573 (N_14573,N_7069,N_9826);
nor U14574 (N_14574,N_5698,N_5978);
and U14575 (N_14575,N_9465,N_6336);
nor U14576 (N_14576,N_8449,N_5144);
xnor U14577 (N_14577,N_9854,N_9270);
and U14578 (N_14578,N_8926,N_7652);
or U14579 (N_14579,N_5828,N_6790);
nor U14580 (N_14580,N_9223,N_5199);
nor U14581 (N_14581,N_6772,N_7565);
xor U14582 (N_14582,N_6087,N_5882);
nand U14583 (N_14583,N_9509,N_9049);
and U14584 (N_14584,N_7656,N_9317);
xor U14585 (N_14585,N_5100,N_7987);
xnor U14586 (N_14586,N_6917,N_9059);
nor U14587 (N_14587,N_5955,N_5382);
or U14588 (N_14588,N_5831,N_8467);
or U14589 (N_14589,N_5827,N_5124);
nand U14590 (N_14590,N_9615,N_6836);
or U14591 (N_14591,N_5334,N_6595);
xnor U14592 (N_14592,N_7458,N_8408);
xnor U14593 (N_14593,N_9817,N_8282);
and U14594 (N_14594,N_8164,N_5202);
or U14595 (N_14595,N_5269,N_8054);
or U14596 (N_14596,N_9745,N_8952);
nand U14597 (N_14597,N_7341,N_9791);
nand U14598 (N_14598,N_8725,N_6215);
and U14599 (N_14599,N_9599,N_7095);
xor U14600 (N_14600,N_7992,N_7928);
nand U14601 (N_14601,N_5695,N_7362);
and U14602 (N_14602,N_7071,N_7354);
and U14603 (N_14603,N_9105,N_6247);
and U14604 (N_14604,N_6880,N_7876);
nor U14605 (N_14605,N_8498,N_6124);
or U14606 (N_14606,N_8114,N_6900);
or U14607 (N_14607,N_9837,N_7301);
nand U14608 (N_14608,N_8458,N_6195);
nor U14609 (N_14609,N_7815,N_5681);
and U14610 (N_14610,N_9295,N_5651);
xnor U14611 (N_14611,N_7704,N_6064);
and U14612 (N_14612,N_7713,N_5629);
or U14613 (N_14613,N_7612,N_7528);
xor U14614 (N_14614,N_5226,N_8773);
or U14615 (N_14615,N_5694,N_8222);
xor U14616 (N_14616,N_5459,N_9554);
xor U14617 (N_14617,N_7547,N_6960);
nand U14618 (N_14618,N_6208,N_8049);
and U14619 (N_14619,N_5673,N_5381);
and U14620 (N_14620,N_8196,N_9899);
xor U14621 (N_14621,N_5201,N_8408);
nand U14622 (N_14622,N_7595,N_5862);
nor U14623 (N_14623,N_7573,N_8257);
nand U14624 (N_14624,N_8716,N_5863);
xor U14625 (N_14625,N_8061,N_6395);
nor U14626 (N_14626,N_6891,N_6382);
or U14627 (N_14627,N_8070,N_9796);
and U14628 (N_14628,N_9077,N_8789);
xor U14629 (N_14629,N_7958,N_5766);
nor U14630 (N_14630,N_6511,N_7432);
and U14631 (N_14631,N_5900,N_5791);
and U14632 (N_14632,N_8004,N_9538);
and U14633 (N_14633,N_5015,N_5105);
nor U14634 (N_14634,N_5382,N_9542);
xnor U14635 (N_14635,N_9519,N_7702);
nor U14636 (N_14636,N_7426,N_7749);
xnor U14637 (N_14637,N_9280,N_6841);
or U14638 (N_14638,N_7633,N_9757);
or U14639 (N_14639,N_9963,N_7524);
xnor U14640 (N_14640,N_9521,N_7962);
nor U14641 (N_14641,N_9419,N_5060);
nor U14642 (N_14642,N_8369,N_9877);
nand U14643 (N_14643,N_9290,N_7980);
nor U14644 (N_14644,N_9729,N_8379);
nand U14645 (N_14645,N_6824,N_8414);
or U14646 (N_14646,N_6020,N_6012);
or U14647 (N_14647,N_7842,N_6607);
and U14648 (N_14648,N_6401,N_9324);
and U14649 (N_14649,N_9968,N_9821);
or U14650 (N_14650,N_8999,N_6696);
or U14651 (N_14651,N_9570,N_9298);
and U14652 (N_14652,N_7652,N_5227);
and U14653 (N_14653,N_5319,N_8182);
nor U14654 (N_14654,N_9431,N_9882);
and U14655 (N_14655,N_6193,N_8841);
xnor U14656 (N_14656,N_8849,N_5064);
nor U14657 (N_14657,N_6939,N_5290);
or U14658 (N_14658,N_9041,N_8159);
or U14659 (N_14659,N_7966,N_9431);
nand U14660 (N_14660,N_7302,N_9904);
and U14661 (N_14661,N_5547,N_5027);
nand U14662 (N_14662,N_8554,N_5246);
and U14663 (N_14663,N_8065,N_9699);
nand U14664 (N_14664,N_6209,N_9871);
or U14665 (N_14665,N_5078,N_6272);
nor U14666 (N_14666,N_6992,N_8267);
and U14667 (N_14667,N_7264,N_8145);
nand U14668 (N_14668,N_6136,N_7486);
and U14669 (N_14669,N_7758,N_8538);
or U14670 (N_14670,N_8693,N_5737);
or U14671 (N_14671,N_6766,N_6159);
nand U14672 (N_14672,N_5655,N_6631);
or U14673 (N_14673,N_5829,N_9635);
or U14674 (N_14674,N_8946,N_8009);
xor U14675 (N_14675,N_9355,N_8054);
nand U14676 (N_14676,N_6561,N_5440);
nor U14677 (N_14677,N_5289,N_7122);
or U14678 (N_14678,N_7298,N_5051);
and U14679 (N_14679,N_5375,N_5822);
xnor U14680 (N_14680,N_7129,N_5901);
and U14681 (N_14681,N_9017,N_8400);
nor U14682 (N_14682,N_8495,N_8861);
nor U14683 (N_14683,N_5161,N_6553);
and U14684 (N_14684,N_6446,N_9447);
nand U14685 (N_14685,N_6452,N_8998);
or U14686 (N_14686,N_7183,N_9180);
or U14687 (N_14687,N_8044,N_8264);
or U14688 (N_14688,N_8994,N_9423);
nor U14689 (N_14689,N_6009,N_9853);
nand U14690 (N_14690,N_8784,N_5188);
and U14691 (N_14691,N_9773,N_8273);
xor U14692 (N_14692,N_6672,N_8739);
nor U14693 (N_14693,N_9508,N_6211);
and U14694 (N_14694,N_9414,N_6298);
or U14695 (N_14695,N_7644,N_8739);
xor U14696 (N_14696,N_8527,N_6374);
nand U14697 (N_14697,N_9189,N_6035);
nand U14698 (N_14698,N_6338,N_9040);
nor U14699 (N_14699,N_6664,N_9225);
nor U14700 (N_14700,N_6438,N_5370);
nor U14701 (N_14701,N_7316,N_8208);
nand U14702 (N_14702,N_5468,N_6941);
or U14703 (N_14703,N_6970,N_9948);
and U14704 (N_14704,N_8448,N_8887);
or U14705 (N_14705,N_8682,N_7630);
and U14706 (N_14706,N_9184,N_6608);
nor U14707 (N_14707,N_9749,N_6022);
xor U14708 (N_14708,N_5953,N_7386);
nand U14709 (N_14709,N_8354,N_8049);
nand U14710 (N_14710,N_9411,N_7811);
nor U14711 (N_14711,N_6912,N_7435);
or U14712 (N_14712,N_9669,N_6075);
nand U14713 (N_14713,N_8987,N_5845);
nor U14714 (N_14714,N_6832,N_9618);
or U14715 (N_14715,N_8381,N_9320);
and U14716 (N_14716,N_7591,N_5820);
or U14717 (N_14717,N_8651,N_5589);
or U14718 (N_14718,N_9185,N_9565);
nand U14719 (N_14719,N_9842,N_8511);
nor U14720 (N_14720,N_9955,N_5721);
or U14721 (N_14721,N_7148,N_7785);
or U14722 (N_14722,N_5106,N_8923);
nor U14723 (N_14723,N_5770,N_9228);
nand U14724 (N_14724,N_6966,N_5633);
xor U14725 (N_14725,N_9146,N_7501);
nor U14726 (N_14726,N_7460,N_8767);
or U14727 (N_14727,N_9487,N_9196);
and U14728 (N_14728,N_7287,N_7213);
xor U14729 (N_14729,N_7108,N_9115);
nor U14730 (N_14730,N_7449,N_6416);
nand U14731 (N_14731,N_6103,N_8175);
nor U14732 (N_14732,N_8467,N_8437);
nand U14733 (N_14733,N_7795,N_7567);
and U14734 (N_14734,N_9919,N_5337);
and U14735 (N_14735,N_9396,N_8125);
nand U14736 (N_14736,N_5981,N_9616);
xor U14737 (N_14737,N_9256,N_8338);
and U14738 (N_14738,N_9365,N_8249);
or U14739 (N_14739,N_8367,N_6241);
nand U14740 (N_14740,N_6403,N_9734);
or U14741 (N_14741,N_8991,N_5816);
or U14742 (N_14742,N_7811,N_5355);
nand U14743 (N_14743,N_6050,N_8964);
nand U14744 (N_14744,N_5099,N_5576);
xnor U14745 (N_14745,N_9539,N_8934);
nand U14746 (N_14746,N_9408,N_7137);
nor U14747 (N_14747,N_8512,N_7767);
or U14748 (N_14748,N_5851,N_7013);
and U14749 (N_14749,N_5611,N_9433);
xor U14750 (N_14750,N_7805,N_9862);
nand U14751 (N_14751,N_9095,N_9501);
nor U14752 (N_14752,N_8666,N_7558);
xor U14753 (N_14753,N_8134,N_7204);
nor U14754 (N_14754,N_5670,N_8722);
and U14755 (N_14755,N_5848,N_9436);
xnor U14756 (N_14756,N_8779,N_9092);
nor U14757 (N_14757,N_8238,N_5676);
nand U14758 (N_14758,N_7537,N_5282);
or U14759 (N_14759,N_6775,N_9092);
or U14760 (N_14760,N_6724,N_5591);
nand U14761 (N_14761,N_9123,N_7171);
nor U14762 (N_14762,N_6644,N_6817);
and U14763 (N_14763,N_7295,N_8180);
or U14764 (N_14764,N_7597,N_8799);
and U14765 (N_14765,N_6078,N_9995);
or U14766 (N_14766,N_5390,N_7889);
or U14767 (N_14767,N_9772,N_7727);
or U14768 (N_14768,N_7785,N_9569);
nand U14769 (N_14769,N_9379,N_5735);
xnor U14770 (N_14770,N_7912,N_8605);
nand U14771 (N_14771,N_9399,N_5731);
or U14772 (N_14772,N_6731,N_9408);
or U14773 (N_14773,N_5510,N_6759);
xor U14774 (N_14774,N_5875,N_6969);
or U14775 (N_14775,N_6740,N_7357);
nor U14776 (N_14776,N_8252,N_5823);
xnor U14777 (N_14777,N_9379,N_8753);
xnor U14778 (N_14778,N_8683,N_7745);
nand U14779 (N_14779,N_6568,N_8144);
nor U14780 (N_14780,N_6018,N_9313);
or U14781 (N_14781,N_8380,N_6837);
xor U14782 (N_14782,N_7765,N_6528);
or U14783 (N_14783,N_9641,N_6701);
xnor U14784 (N_14784,N_5482,N_6833);
or U14785 (N_14785,N_6666,N_8313);
nor U14786 (N_14786,N_8678,N_7091);
nor U14787 (N_14787,N_9485,N_9528);
and U14788 (N_14788,N_9143,N_8103);
xnor U14789 (N_14789,N_6529,N_6356);
xor U14790 (N_14790,N_8954,N_5543);
nand U14791 (N_14791,N_8240,N_9712);
xor U14792 (N_14792,N_5230,N_5795);
xnor U14793 (N_14793,N_8489,N_7202);
and U14794 (N_14794,N_6511,N_6876);
and U14795 (N_14795,N_8932,N_6964);
or U14796 (N_14796,N_9618,N_9449);
or U14797 (N_14797,N_5975,N_7077);
nor U14798 (N_14798,N_5725,N_7805);
nor U14799 (N_14799,N_7298,N_9374);
nand U14800 (N_14800,N_5366,N_8438);
nor U14801 (N_14801,N_7146,N_5764);
xnor U14802 (N_14802,N_7867,N_7022);
nor U14803 (N_14803,N_5518,N_6251);
xor U14804 (N_14804,N_7457,N_7154);
xor U14805 (N_14805,N_6568,N_5589);
nor U14806 (N_14806,N_5359,N_8769);
xnor U14807 (N_14807,N_6867,N_5964);
xnor U14808 (N_14808,N_8688,N_8216);
and U14809 (N_14809,N_7325,N_8831);
nand U14810 (N_14810,N_8546,N_5651);
nand U14811 (N_14811,N_7920,N_6009);
xor U14812 (N_14812,N_8232,N_5868);
xnor U14813 (N_14813,N_8656,N_6255);
nand U14814 (N_14814,N_9223,N_9450);
nor U14815 (N_14815,N_6313,N_5027);
nor U14816 (N_14816,N_9408,N_5805);
nand U14817 (N_14817,N_5501,N_6273);
or U14818 (N_14818,N_8916,N_7692);
xor U14819 (N_14819,N_7960,N_7001);
nor U14820 (N_14820,N_8447,N_5871);
or U14821 (N_14821,N_7572,N_7240);
nand U14822 (N_14822,N_9371,N_6887);
or U14823 (N_14823,N_5100,N_7608);
nor U14824 (N_14824,N_9962,N_6942);
or U14825 (N_14825,N_6194,N_8795);
and U14826 (N_14826,N_9308,N_5098);
nor U14827 (N_14827,N_7086,N_7900);
nor U14828 (N_14828,N_8298,N_8979);
xnor U14829 (N_14829,N_8298,N_5217);
xnor U14830 (N_14830,N_5081,N_8899);
or U14831 (N_14831,N_9742,N_5235);
nand U14832 (N_14832,N_8409,N_7784);
nand U14833 (N_14833,N_5711,N_8144);
or U14834 (N_14834,N_5387,N_5444);
nand U14835 (N_14835,N_8020,N_5368);
nor U14836 (N_14836,N_8057,N_9924);
nand U14837 (N_14837,N_5682,N_9392);
nor U14838 (N_14838,N_7718,N_7136);
xnor U14839 (N_14839,N_8838,N_9303);
or U14840 (N_14840,N_8230,N_9986);
nor U14841 (N_14841,N_7087,N_7407);
nand U14842 (N_14842,N_8349,N_5053);
nand U14843 (N_14843,N_8885,N_8720);
and U14844 (N_14844,N_8674,N_5959);
nand U14845 (N_14845,N_9295,N_8668);
and U14846 (N_14846,N_8895,N_6837);
xor U14847 (N_14847,N_6748,N_5781);
nand U14848 (N_14848,N_9902,N_5293);
and U14849 (N_14849,N_7810,N_6135);
and U14850 (N_14850,N_9717,N_9469);
and U14851 (N_14851,N_7452,N_6991);
and U14852 (N_14852,N_7561,N_5139);
xor U14853 (N_14853,N_5296,N_8531);
nand U14854 (N_14854,N_9426,N_8878);
or U14855 (N_14855,N_6237,N_7236);
and U14856 (N_14856,N_9942,N_8065);
nand U14857 (N_14857,N_8866,N_8453);
nor U14858 (N_14858,N_7214,N_9738);
nand U14859 (N_14859,N_8506,N_6536);
nor U14860 (N_14860,N_7021,N_7504);
or U14861 (N_14861,N_5900,N_9126);
and U14862 (N_14862,N_6045,N_9516);
nor U14863 (N_14863,N_6134,N_5914);
nand U14864 (N_14864,N_6895,N_7214);
and U14865 (N_14865,N_7410,N_6796);
xnor U14866 (N_14866,N_9198,N_6727);
xor U14867 (N_14867,N_8063,N_6409);
nand U14868 (N_14868,N_7152,N_9332);
nand U14869 (N_14869,N_7545,N_6086);
xnor U14870 (N_14870,N_9440,N_6914);
nor U14871 (N_14871,N_7857,N_9717);
or U14872 (N_14872,N_5479,N_5032);
nor U14873 (N_14873,N_9612,N_8085);
or U14874 (N_14874,N_5011,N_7502);
and U14875 (N_14875,N_9313,N_5846);
nor U14876 (N_14876,N_9712,N_6903);
xor U14877 (N_14877,N_6189,N_5715);
nand U14878 (N_14878,N_7171,N_9452);
or U14879 (N_14879,N_6765,N_9684);
xnor U14880 (N_14880,N_6223,N_9015);
nand U14881 (N_14881,N_8914,N_6934);
nor U14882 (N_14882,N_9330,N_8469);
nor U14883 (N_14883,N_6918,N_7355);
and U14884 (N_14884,N_9620,N_7856);
and U14885 (N_14885,N_8266,N_8329);
or U14886 (N_14886,N_8787,N_5940);
and U14887 (N_14887,N_8947,N_8989);
or U14888 (N_14888,N_8931,N_7549);
or U14889 (N_14889,N_6443,N_8929);
and U14890 (N_14890,N_5621,N_7037);
nor U14891 (N_14891,N_6453,N_8203);
nor U14892 (N_14892,N_6200,N_7133);
or U14893 (N_14893,N_9583,N_8670);
or U14894 (N_14894,N_8490,N_8425);
nand U14895 (N_14895,N_7527,N_9364);
and U14896 (N_14896,N_7101,N_9886);
nor U14897 (N_14897,N_8221,N_9675);
nand U14898 (N_14898,N_9726,N_5642);
nand U14899 (N_14899,N_5641,N_9779);
xnor U14900 (N_14900,N_7990,N_9824);
and U14901 (N_14901,N_9127,N_6070);
xor U14902 (N_14902,N_7819,N_6729);
nand U14903 (N_14903,N_9932,N_6392);
nand U14904 (N_14904,N_9710,N_6150);
nor U14905 (N_14905,N_8638,N_6902);
or U14906 (N_14906,N_6672,N_6587);
nand U14907 (N_14907,N_5837,N_7692);
or U14908 (N_14908,N_7827,N_8895);
nor U14909 (N_14909,N_5152,N_7005);
xor U14910 (N_14910,N_6312,N_8578);
and U14911 (N_14911,N_6470,N_6360);
or U14912 (N_14912,N_8842,N_9839);
nand U14913 (N_14913,N_6158,N_6026);
xor U14914 (N_14914,N_8878,N_6021);
xnor U14915 (N_14915,N_9389,N_7834);
xnor U14916 (N_14916,N_9030,N_8088);
nand U14917 (N_14917,N_9972,N_9069);
xnor U14918 (N_14918,N_6777,N_5615);
xnor U14919 (N_14919,N_6632,N_7249);
xnor U14920 (N_14920,N_7411,N_9401);
xor U14921 (N_14921,N_5756,N_8387);
nand U14922 (N_14922,N_8541,N_5388);
nor U14923 (N_14923,N_9166,N_6143);
xor U14924 (N_14924,N_7216,N_9979);
nand U14925 (N_14925,N_7629,N_6683);
nand U14926 (N_14926,N_6444,N_8647);
nand U14927 (N_14927,N_6325,N_5808);
nand U14928 (N_14928,N_6203,N_5191);
nor U14929 (N_14929,N_7090,N_5640);
nor U14930 (N_14930,N_5018,N_5699);
nor U14931 (N_14931,N_8766,N_8947);
nand U14932 (N_14932,N_5338,N_8724);
nand U14933 (N_14933,N_8238,N_9863);
nor U14934 (N_14934,N_9394,N_9828);
or U14935 (N_14935,N_8007,N_6737);
and U14936 (N_14936,N_7018,N_5255);
or U14937 (N_14937,N_9119,N_5252);
nand U14938 (N_14938,N_7240,N_9743);
and U14939 (N_14939,N_9659,N_6156);
nor U14940 (N_14940,N_6918,N_5340);
or U14941 (N_14941,N_8137,N_9206);
and U14942 (N_14942,N_7181,N_9431);
or U14943 (N_14943,N_6352,N_7622);
nor U14944 (N_14944,N_9861,N_5503);
nand U14945 (N_14945,N_5249,N_7329);
or U14946 (N_14946,N_5034,N_9791);
or U14947 (N_14947,N_8316,N_8249);
nand U14948 (N_14948,N_8333,N_8463);
or U14949 (N_14949,N_6387,N_5162);
nand U14950 (N_14950,N_9646,N_7421);
xor U14951 (N_14951,N_5053,N_6729);
or U14952 (N_14952,N_5723,N_7124);
and U14953 (N_14953,N_9458,N_5988);
and U14954 (N_14954,N_7453,N_5763);
nor U14955 (N_14955,N_8210,N_7219);
xor U14956 (N_14956,N_8268,N_8245);
nor U14957 (N_14957,N_9165,N_9950);
nand U14958 (N_14958,N_6889,N_6148);
or U14959 (N_14959,N_6015,N_8465);
xor U14960 (N_14960,N_5116,N_7348);
or U14961 (N_14961,N_7015,N_8924);
and U14962 (N_14962,N_6056,N_8915);
nand U14963 (N_14963,N_8500,N_9620);
xnor U14964 (N_14964,N_6462,N_7741);
or U14965 (N_14965,N_8058,N_7488);
nor U14966 (N_14966,N_5330,N_5628);
nand U14967 (N_14967,N_8718,N_6832);
or U14968 (N_14968,N_7846,N_8200);
and U14969 (N_14969,N_6767,N_6511);
xor U14970 (N_14970,N_5566,N_6201);
or U14971 (N_14971,N_7707,N_8302);
nor U14972 (N_14972,N_9754,N_9249);
xnor U14973 (N_14973,N_9052,N_7295);
nand U14974 (N_14974,N_5379,N_9577);
and U14975 (N_14975,N_7324,N_8286);
nor U14976 (N_14976,N_6160,N_7222);
nand U14977 (N_14977,N_6989,N_6745);
or U14978 (N_14978,N_5943,N_8630);
and U14979 (N_14979,N_7136,N_8363);
and U14980 (N_14980,N_5662,N_8927);
nand U14981 (N_14981,N_7093,N_7325);
nor U14982 (N_14982,N_6383,N_6257);
nand U14983 (N_14983,N_7325,N_6204);
nor U14984 (N_14984,N_9684,N_8030);
or U14985 (N_14985,N_5818,N_5562);
nor U14986 (N_14986,N_8051,N_7036);
nand U14987 (N_14987,N_5609,N_5970);
xnor U14988 (N_14988,N_6116,N_7608);
or U14989 (N_14989,N_9631,N_7289);
xnor U14990 (N_14990,N_5455,N_7902);
and U14991 (N_14991,N_8464,N_8758);
nand U14992 (N_14992,N_5524,N_8653);
or U14993 (N_14993,N_8340,N_7667);
nand U14994 (N_14994,N_5477,N_7786);
and U14995 (N_14995,N_8516,N_8964);
nor U14996 (N_14996,N_7226,N_8129);
and U14997 (N_14997,N_6789,N_9394);
or U14998 (N_14998,N_5662,N_8742);
nor U14999 (N_14999,N_7176,N_5736);
and U15000 (N_15000,N_12399,N_10300);
or U15001 (N_15001,N_10749,N_10108);
or U15002 (N_15002,N_13515,N_14456);
nand U15003 (N_15003,N_13660,N_12752);
nor U15004 (N_15004,N_11830,N_11142);
and U15005 (N_15005,N_10505,N_12858);
nand U15006 (N_15006,N_12158,N_14847);
nand U15007 (N_15007,N_10280,N_14152);
or U15008 (N_15008,N_13105,N_11658);
nand U15009 (N_15009,N_12317,N_14066);
nor U15010 (N_15010,N_11898,N_10946);
and U15011 (N_15011,N_12663,N_11162);
nand U15012 (N_15012,N_11764,N_10243);
nor U15013 (N_15013,N_14526,N_12491);
or U15014 (N_15014,N_13494,N_14362);
xnor U15015 (N_15015,N_14041,N_14323);
or U15016 (N_15016,N_12339,N_10561);
and U15017 (N_15017,N_11771,N_12330);
xnor U15018 (N_15018,N_13480,N_10146);
xor U15019 (N_15019,N_12211,N_12885);
nor U15020 (N_15020,N_13240,N_14201);
or U15021 (N_15021,N_13157,N_10544);
and U15022 (N_15022,N_11973,N_10863);
nand U15023 (N_15023,N_14430,N_10499);
nand U15024 (N_15024,N_10275,N_11543);
or U15025 (N_15025,N_12232,N_12954);
and U15026 (N_15026,N_10633,N_13552);
nor U15027 (N_15027,N_14254,N_12168);
xnor U15028 (N_15028,N_14730,N_10770);
xor U15029 (N_15029,N_13910,N_10453);
xnor U15030 (N_15030,N_14422,N_11676);
and U15031 (N_15031,N_13895,N_11605);
and U15032 (N_15032,N_14502,N_14276);
or U15033 (N_15033,N_14772,N_10614);
nor U15034 (N_15034,N_11047,N_11890);
xor U15035 (N_15035,N_11324,N_13947);
nand U15036 (N_15036,N_11222,N_12333);
xnor U15037 (N_15037,N_10820,N_11772);
and U15038 (N_15038,N_12682,N_11647);
nand U15039 (N_15039,N_14272,N_11055);
xor U15040 (N_15040,N_12124,N_12804);
nor U15041 (N_15041,N_10679,N_13846);
nand U15042 (N_15042,N_10455,N_13186);
xnor U15043 (N_15043,N_13449,N_12457);
xor U15044 (N_15044,N_11295,N_13185);
or U15045 (N_15045,N_12262,N_12319);
and U15046 (N_15046,N_12878,N_12697);
or U15047 (N_15047,N_13622,N_11316);
nand U15048 (N_15048,N_13589,N_14259);
and U15049 (N_15049,N_10128,N_12521);
and U15050 (N_15050,N_14590,N_14396);
xnor U15051 (N_15051,N_12868,N_13254);
or U15052 (N_15052,N_10129,N_11422);
nor U15053 (N_15053,N_11573,N_11026);
nor U15054 (N_15054,N_10303,N_11665);
or U15055 (N_15055,N_11419,N_11218);
xor U15056 (N_15056,N_11190,N_12083);
nor U15057 (N_15057,N_11261,N_12283);
nand U15058 (N_15058,N_14770,N_14987);
nand U15059 (N_15059,N_14509,N_11488);
xor U15060 (N_15060,N_12739,N_14186);
and U15061 (N_15061,N_14579,N_13850);
xnor U15062 (N_15062,N_12438,N_14895);
xor U15063 (N_15063,N_14697,N_10061);
nor U15064 (N_15064,N_12583,N_10589);
or U15065 (N_15065,N_13357,N_14615);
nor U15066 (N_15066,N_11394,N_13058);
nand U15067 (N_15067,N_12948,N_13182);
nor U15068 (N_15068,N_11482,N_11352);
nor U15069 (N_15069,N_14985,N_11208);
and U15070 (N_15070,N_10931,N_11972);
nand U15071 (N_15071,N_13626,N_13728);
or U15072 (N_15072,N_11227,N_13315);
nor U15073 (N_15073,N_11072,N_11114);
nand U15074 (N_15074,N_13891,N_11305);
xnor U15075 (N_15075,N_12425,N_14291);
or U15076 (N_15076,N_11291,N_10055);
xnor U15077 (N_15077,N_10639,N_12151);
xnor U15078 (N_15078,N_13423,N_11743);
nor U15079 (N_15079,N_12811,N_11398);
nor U15080 (N_15080,N_11083,N_14085);
or U15081 (N_15081,N_14106,N_13371);
or U15082 (N_15082,N_13924,N_14251);
xor U15083 (N_15083,N_10158,N_12581);
xnor U15084 (N_15084,N_13313,N_14530);
nand U15085 (N_15085,N_11776,N_12516);
nand U15086 (N_15086,N_13279,N_12287);
and U15087 (N_15087,N_14120,N_12869);
or U15088 (N_15088,N_12386,N_13311);
or U15089 (N_15089,N_12767,N_10764);
or U15090 (N_15090,N_13887,N_10439);
or U15091 (N_15091,N_14258,N_14067);
nor U15092 (N_15092,N_10078,N_13642);
nor U15093 (N_15093,N_10757,N_10669);
nand U15094 (N_15094,N_14571,N_10062);
and U15095 (N_15095,N_14607,N_10646);
xnor U15096 (N_15096,N_14787,N_11067);
nand U15097 (N_15097,N_14118,N_12635);
nor U15098 (N_15098,N_10445,N_13390);
xnor U15099 (N_15099,N_11399,N_12022);
and U15100 (N_15100,N_12822,N_10310);
and U15101 (N_15101,N_13573,N_10008);
xor U15102 (N_15102,N_12346,N_12238);
xor U15103 (N_15103,N_11909,N_10379);
nor U15104 (N_15104,N_10793,N_10417);
nor U15105 (N_15105,N_12949,N_14346);
or U15106 (N_15106,N_14551,N_13055);
or U15107 (N_15107,N_12786,N_14942);
or U15108 (N_15108,N_10166,N_12369);
or U15109 (N_15109,N_13419,N_13292);
nor U15110 (N_15110,N_12508,N_13250);
xor U15111 (N_15111,N_11088,N_14282);
nand U15112 (N_15112,N_14388,N_11643);
and U15113 (N_15113,N_11532,N_11683);
xor U15114 (N_15114,N_14614,N_12315);
xnor U15115 (N_15115,N_10352,N_11705);
nand U15116 (N_15116,N_10965,N_12305);
or U15117 (N_15117,N_13147,N_14859);
xor U15118 (N_15118,N_10291,N_12887);
nand U15119 (N_15119,N_12637,N_11477);
or U15120 (N_15120,N_11744,N_14367);
xor U15121 (N_15121,N_12934,N_12031);
or U15122 (N_15122,N_13590,N_13333);
and U15123 (N_15123,N_13676,N_10524);
or U15124 (N_15124,N_11193,N_13782);
nor U15125 (N_15125,N_14052,N_11448);
xor U15126 (N_15126,N_13738,N_12100);
xnor U15127 (N_15127,N_14943,N_12742);
nand U15128 (N_15128,N_10380,N_14515);
xnor U15129 (N_15129,N_13765,N_11124);
and U15130 (N_15130,N_10412,N_10617);
nand U15131 (N_15131,N_14026,N_13392);
xnor U15132 (N_15132,N_12443,N_14944);
or U15133 (N_15133,N_13961,N_10497);
or U15134 (N_15134,N_13032,N_13592);
and U15135 (N_15135,N_12961,N_12833);
nand U15136 (N_15136,N_12906,N_10720);
nor U15137 (N_15137,N_13889,N_13537);
and U15138 (N_15138,N_14431,N_13374);
xor U15139 (N_15139,N_10134,N_14331);
xnor U15140 (N_15140,N_13702,N_14232);
xnor U15141 (N_15141,N_10853,N_11248);
xnor U15142 (N_15142,N_12461,N_12677);
xor U15143 (N_15143,N_12471,N_14593);
nor U15144 (N_15144,N_14602,N_10269);
xnor U15145 (N_15145,N_12827,N_14330);
nand U15146 (N_15146,N_11286,N_14592);
xnor U15147 (N_15147,N_12638,N_11080);
or U15148 (N_15148,N_10001,N_10059);
and U15149 (N_15149,N_12937,N_14700);
nand U15150 (N_15150,N_12033,N_12842);
nand U15151 (N_15151,N_11712,N_10927);
and U15152 (N_15152,N_13249,N_12750);
or U15153 (N_15153,N_10210,N_10758);
and U15154 (N_15154,N_13714,N_13244);
nor U15155 (N_15155,N_13836,N_12215);
xor U15156 (N_15156,N_13065,N_12908);
xor U15157 (N_15157,N_12301,N_14966);
or U15158 (N_15158,N_14872,N_10751);
and U15159 (N_15159,N_10692,N_12228);
xnor U15160 (N_15160,N_14426,N_12907);
or U15161 (N_15161,N_12856,N_12395);
nand U15162 (N_15162,N_11178,N_10294);
nand U15163 (N_15163,N_13927,N_14096);
and U15164 (N_15164,N_10151,N_12819);
or U15165 (N_15165,N_10962,N_11366);
or U15166 (N_15166,N_10356,N_11495);
nor U15167 (N_15167,N_10771,N_14223);
and U15168 (N_15168,N_12536,N_14350);
xnor U15169 (N_15169,N_13863,N_13213);
nand U15170 (N_15170,N_13668,N_13010);
and U15171 (N_15171,N_12094,N_11635);
nor U15172 (N_15172,N_12313,N_10423);
and U15173 (N_15173,N_13726,N_12629);
nand U15174 (N_15174,N_14497,N_14459);
xor U15175 (N_15175,N_12743,N_11803);
nor U15176 (N_15176,N_10986,N_12668);
nor U15177 (N_15177,N_11202,N_14403);
and U15178 (N_15178,N_10244,N_11367);
or U15179 (N_15179,N_14786,N_13657);
xor U15180 (N_15180,N_11622,N_12986);
or U15181 (N_15181,N_13951,N_14364);
nor U15182 (N_15182,N_10349,N_10305);
or U15183 (N_15183,N_13320,N_14691);
or U15184 (N_15184,N_13689,N_10850);
and U15185 (N_15185,N_12029,N_14482);
or U15186 (N_15186,N_13627,N_10107);
or U15187 (N_15187,N_10176,N_13131);
nand U15188 (N_15188,N_12188,N_13168);
and U15189 (N_15189,N_10869,N_11078);
nor U15190 (N_15190,N_10492,N_10807);
or U15191 (N_15191,N_13072,N_14032);
nand U15192 (N_15192,N_11045,N_14470);
or U15193 (N_15193,N_12279,N_12383);
nor U15194 (N_15194,N_14976,N_10823);
nor U15195 (N_15195,N_10640,N_14924);
xor U15196 (N_15196,N_14940,N_14601);
nor U15197 (N_15197,N_12712,N_11581);
nand U15198 (N_15198,N_12701,N_14387);
xnor U15199 (N_15199,N_11356,N_14301);
nand U15200 (N_15200,N_13975,N_11628);
nor U15201 (N_15201,N_13859,N_10095);
or U15202 (N_15202,N_11654,N_12667);
nor U15203 (N_15203,N_13923,N_13766);
nor U15204 (N_15204,N_12327,N_12512);
or U15205 (N_15205,N_11594,N_13183);
nor U15206 (N_15206,N_11907,N_14511);
nor U15207 (N_15207,N_10448,N_14514);
or U15208 (N_15208,N_11309,N_10385);
or U15209 (N_15209,N_14135,N_12639);
or U15210 (N_15210,N_14824,N_13275);
and U15211 (N_15211,N_10367,N_13780);
and U15212 (N_15212,N_13477,N_12787);
or U15213 (N_15213,N_13328,N_10917);
or U15214 (N_15214,N_13653,N_10474);
nand U15215 (N_15215,N_11157,N_12197);
xor U15216 (N_15216,N_10595,N_12883);
or U15217 (N_15217,N_13483,N_11065);
and U15218 (N_15218,N_12746,N_10715);
xor U15219 (N_15219,N_14908,N_12494);
nand U15220 (N_15220,N_14153,N_11423);
or U15221 (N_15221,N_11735,N_14584);
or U15222 (N_15222,N_13302,N_12281);
or U15223 (N_15223,N_12612,N_14823);
or U15224 (N_15224,N_10738,N_10763);
xor U15225 (N_15225,N_14481,N_10112);
nor U15226 (N_15226,N_13406,N_13118);
or U15227 (N_15227,N_14485,N_10289);
nor U15228 (N_15228,N_10317,N_13324);
and U15229 (N_15229,N_11897,N_12765);
xor U15230 (N_15230,N_10264,N_11499);
and U15231 (N_15231,N_14206,N_13683);
and U15232 (N_15232,N_14839,N_13500);
nand U15233 (N_15233,N_13326,N_11273);
xnor U15234 (N_15234,N_13750,N_12651);
or U15235 (N_15235,N_14998,N_12304);
and U15236 (N_15236,N_13002,N_14719);
or U15237 (N_15237,N_11413,N_14705);
nand U15238 (N_15238,N_13097,N_13918);
and U15239 (N_15239,N_13802,N_12077);
nor U15240 (N_15240,N_10558,N_11593);
nand U15241 (N_15241,N_10707,N_12368);
nand U15242 (N_15242,N_10673,N_10579);
nand U15243 (N_15243,N_11652,N_13246);
xor U15244 (N_15244,N_11756,N_11237);
and U15245 (N_15245,N_10875,N_10525);
nor U15246 (N_15246,N_13847,N_12503);
nor U15247 (N_15247,N_11935,N_10753);
and U15248 (N_15248,N_10482,N_12111);
nor U15249 (N_15249,N_10837,N_14308);
nand U15250 (N_15250,N_13277,N_11453);
nor U15251 (N_15251,N_10478,N_10173);
or U15252 (N_15252,N_13337,N_14755);
and U15253 (N_15253,N_14935,N_13070);
or U15254 (N_15254,N_13632,N_12614);
xor U15255 (N_15255,N_12392,N_13022);
nor U15256 (N_15256,N_11904,N_13497);
xor U15257 (N_15257,N_14319,N_14636);
or U15258 (N_15258,N_10967,N_12550);
nor U15259 (N_15259,N_13164,N_10740);
and U15260 (N_15260,N_12467,N_10945);
nor U15261 (N_15261,N_13221,N_10642);
nand U15262 (N_15262,N_14196,N_10442);
nor U15263 (N_15263,N_11836,N_12160);
and U15264 (N_15264,N_14917,N_13753);
and U15265 (N_15265,N_11982,N_12627);
or U15266 (N_15266,N_14270,N_14970);
nand U15267 (N_15267,N_11094,N_14816);
and U15268 (N_15268,N_13485,N_14825);
nor U15269 (N_15269,N_14570,N_14443);
nor U15270 (N_15270,N_12821,N_11504);
or U15271 (N_15271,N_10611,N_13977);
and U15272 (N_15272,N_13742,N_11036);
and U15273 (N_15273,N_14046,N_12388);
xor U15274 (N_15274,N_10301,N_13263);
nand U15275 (N_15275,N_12131,N_14833);
or U15276 (N_15276,N_12174,N_12431);
xnor U15277 (N_15277,N_10159,N_14230);
or U15278 (N_15278,N_14469,N_14296);
nor U15279 (N_15279,N_12788,N_14745);
nor U15280 (N_15280,N_10809,N_10429);
or U15281 (N_15281,N_14284,N_11247);
nand U15282 (N_15282,N_13454,N_13867);
nor U15283 (N_15283,N_10529,N_14465);
and U15284 (N_15284,N_11516,N_13016);
xnor U15285 (N_15285,N_11589,N_12762);
nand U15286 (N_15286,N_10788,N_13893);
nor U15287 (N_15287,N_11782,N_11211);
xor U15288 (N_15288,N_12017,N_13545);
nand U15289 (N_15289,N_10454,N_13703);
xnor U15290 (N_15290,N_11116,N_12873);
xor U15291 (N_15291,N_14081,N_13389);
and U15292 (N_15292,N_13856,N_11707);
nor U15293 (N_15293,N_14265,N_11539);
and U15294 (N_15294,N_12783,N_11929);
nand U15295 (N_15295,N_12432,N_14682);
or U15296 (N_15296,N_12509,N_12236);
and U15297 (N_15297,N_10424,N_11472);
nand U15298 (N_15298,N_10171,N_14894);
and U15299 (N_15299,N_11864,N_11338);
and U15300 (N_15300,N_12926,N_12265);
and U15301 (N_15301,N_12394,N_13038);
and U15302 (N_15302,N_10985,N_12882);
nor U15303 (N_15303,N_14650,N_10415);
or U15304 (N_15304,N_11990,N_13957);
and U15305 (N_15305,N_12705,N_11700);
and U15306 (N_15306,N_13476,N_11892);
and U15307 (N_15307,N_13397,N_11823);
nand U15308 (N_15308,N_10480,N_12059);
nor U15309 (N_15309,N_13945,N_13823);
nor U15310 (N_15310,N_14686,N_13214);
nor U15311 (N_15311,N_11763,N_13430);
xor U15312 (N_15312,N_14712,N_10376);
xor U15313 (N_15313,N_14862,N_12540);
nand U15314 (N_15314,N_12161,N_13414);
or U15315 (N_15315,N_11757,N_14802);
xor U15316 (N_15316,N_10947,N_10189);
xnor U15317 (N_15317,N_11161,N_10290);
nor U15318 (N_15318,N_12271,N_11582);
nor U15319 (N_15319,N_10323,N_11318);
nand U15320 (N_15320,N_11086,N_10401);
or U15321 (N_15321,N_10760,N_12644);
xnor U15322 (N_15322,N_13123,N_11923);
nor U15323 (N_15323,N_11588,N_11385);
or U15324 (N_15324,N_11755,N_14725);
nand U15325 (N_15325,N_14168,N_11052);
nor U15326 (N_15326,N_12881,N_11145);
or U15327 (N_15327,N_12119,N_14058);
xor U15328 (N_15328,N_13739,N_11288);
xor U15329 (N_15329,N_10515,N_11739);
or U15330 (N_15330,N_10369,N_10350);
nand U15331 (N_15331,N_12613,N_14436);
xnor U15332 (N_15332,N_11767,N_12433);
or U15333 (N_15333,N_14905,N_10420);
nor U15334 (N_15334,N_14311,N_13906);
nor U15335 (N_15335,N_10632,N_14218);
nor U15336 (N_15336,N_11528,N_13489);
nand U15337 (N_15337,N_14423,N_11538);
nor U15338 (N_15338,N_14566,N_12844);
or U15339 (N_15339,N_13285,N_12449);
and U15340 (N_15340,N_10657,N_13720);
nor U15341 (N_15341,N_12506,N_14213);
nor U15342 (N_15342,N_12071,N_12547);
and U15343 (N_15343,N_14718,N_10004);
nor U15344 (N_15344,N_12553,N_10926);
nor U15345 (N_15345,N_11691,N_12231);
or U15346 (N_15346,N_11922,N_11396);
or U15347 (N_15347,N_11649,N_10890);
xnor U15348 (N_15348,N_13509,N_11406);
and U15349 (N_15349,N_10325,N_14750);
and U15350 (N_15350,N_12387,N_12798);
xor U15351 (N_15351,N_13564,N_13487);
nand U15352 (N_15352,N_11225,N_14869);
nor U15353 (N_15353,N_13654,N_14377);
nand U15354 (N_15354,N_10954,N_14864);
nor U15355 (N_15355,N_12958,N_11063);
and U15356 (N_15356,N_10086,N_11505);
and U15357 (N_15357,N_11167,N_13042);
and U15358 (N_15358,N_13461,N_12303);
xnor U15359 (N_15359,N_11486,N_10813);
or U15360 (N_15360,N_12711,N_12871);
nand U15361 (N_15361,N_12012,N_14659);
xnor U15362 (N_15362,N_13565,N_14145);
xor U15363 (N_15363,N_14710,N_13257);
nand U15364 (N_15364,N_11426,N_11282);
xnor U15365 (N_15365,N_10025,N_14531);
nand U15366 (N_15366,N_11326,N_13132);
nor U15367 (N_15367,N_13675,N_11489);
nand U15368 (N_15368,N_12441,N_11030);
nor U15369 (N_15369,N_14677,N_13855);
nand U15370 (N_15370,N_10832,N_14844);
and U15371 (N_15371,N_10298,N_11737);
and U15372 (N_15372,N_14982,N_11171);
or U15373 (N_15373,N_12589,N_14332);
xor U15374 (N_15374,N_11098,N_10174);
or U15375 (N_15375,N_14294,N_11424);
or U15376 (N_15376,N_11733,N_13754);
and U15377 (N_15377,N_11337,N_13367);
and U15378 (N_15378,N_14372,N_12987);
nand U15379 (N_15379,N_12836,N_13624);
nand U15380 (N_15380,N_12905,N_12706);
xnor U15381 (N_15381,N_14957,N_14252);
nand U15382 (N_15382,N_12414,N_10012);
or U15383 (N_15383,N_14200,N_14945);
or U15384 (N_15384,N_13190,N_11260);
nor U15385 (N_15385,N_10337,N_11113);
nand U15386 (N_15386,N_12212,N_13471);
nor U15387 (N_15387,N_11913,N_10681);
nor U15388 (N_15388,N_13080,N_13608);
and U15389 (N_15389,N_14398,N_14678);
and U15390 (N_15390,N_14445,N_13712);
nor U15391 (N_15391,N_13770,N_11616);
nor U15392 (N_15392,N_11939,N_11115);
xnor U15393 (N_15393,N_10851,N_11514);
or U15394 (N_15394,N_10929,N_12963);
nand U15395 (N_15395,N_10233,N_14305);
nor U15396 (N_15396,N_10916,N_14407);
xnor U15397 (N_15397,N_12167,N_12631);
nand U15398 (N_15398,N_13448,N_12411);
nand U15399 (N_15399,N_12784,N_11947);
and U15400 (N_15400,N_12585,N_13400);
and U15401 (N_15401,N_11561,N_13351);
or U15402 (N_15402,N_11799,N_12171);
nor U15403 (N_15403,N_13099,N_13540);
xor U15404 (N_15404,N_14438,N_10843);
or U15405 (N_15405,N_12719,N_13974);
or U15406 (N_15406,N_11320,N_10238);
or U15407 (N_15407,N_14297,N_12020);
nor U15408 (N_15408,N_14137,N_11391);
nand U15409 (N_15409,N_13685,N_10214);
xor U15410 (N_15410,N_14635,N_14979);
or U15411 (N_15411,N_12173,N_13452);
or U15412 (N_15412,N_11600,N_14409);
nand U15413 (N_15413,N_12038,N_14932);
and U15414 (N_15414,N_11364,N_10148);
nor U15415 (N_15415,N_13365,N_14897);
xor U15416 (N_15416,N_14871,N_10472);
nand U15417 (N_15417,N_12946,N_11359);
xor U15418 (N_15418,N_13198,N_12766);
nand U15419 (N_15419,N_11794,N_14858);
and U15420 (N_15420,N_12886,N_10773);
nand U15421 (N_15421,N_14010,N_12078);
or U15422 (N_15422,N_12685,N_10718);
nand U15423 (N_15423,N_14586,N_11210);
nand U15424 (N_15424,N_13732,N_10028);
nor U15425 (N_15425,N_10103,N_11149);
nand U15426 (N_15426,N_11006,N_11007);
nor U15427 (N_15427,N_10147,N_10339);
nor U15428 (N_15428,N_13585,N_11376);
nor U15429 (N_15429,N_13443,N_12126);
or U15430 (N_15430,N_12434,N_14554);
nor U15431 (N_15431,N_11666,N_11906);
xor U15432 (N_15432,N_14669,N_11182);
nor U15433 (N_15433,N_13432,N_10992);
nand U15434 (N_15434,N_10712,N_10312);
and U15435 (N_15435,N_10162,N_12807);
nor U15436 (N_15436,N_11977,N_14817);
and U15437 (N_15437,N_11267,N_14204);
and U15438 (N_15438,N_12723,N_10045);
or U15439 (N_15439,N_14778,N_11859);
nor U15440 (N_15440,N_14070,N_14887);
or U15441 (N_15441,N_12349,N_13600);
nand U15442 (N_15442,N_11869,N_11832);
or U15443 (N_15443,N_10844,N_10137);
nand U15444 (N_15444,N_14964,N_14476);
and U15445 (N_15445,N_13299,N_10426);
xnor U15446 (N_15446,N_12282,N_12927);
nor U15447 (N_15447,N_14129,N_10365);
xnor U15448 (N_15448,N_14655,N_12335);
xor U15449 (N_15449,N_10332,N_14140);
xor U15450 (N_15450,N_14537,N_13612);
xnor U15451 (N_15451,N_10039,N_10058);
xor U15452 (N_15452,N_12543,N_13534);
nand U15453 (N_15453,N_12430,N_13857);
and U15454 (N_15454,N_13114,N_14993);
xor U15455 (N_15455,N_11708,N_13015);
or U15456 (N_15456,N_13615,N_12732);
xor U15457 (N_15457,N_11966,N_13422);
or U15458 (N_15458,N_12127,N_13428);
nand U15459 (N_15459,N_12754,N_14611);
xnor U15460 (N_15460,N_13735,N_11546);
xor U15461 (N_15461,N_14587,N_13322);
and U15462 (N_15462,N_11634,N_13794);
and U15463 (N_15463,N_12186,N_14320);
and U15464 (N_15464,N_13405,N_12566);
nand U15465 (N_15465,N_11956,N_11004);
and U15466 (N_15466,N_14811,N_12690);
nor U15467 (N_15467,N_10830,N_13883);
nand U15468 (N_15468,N_12214,N_12735);
nor U15469 (N_15469,N_10647,N_13909);
or U15470 (N_15470,N_13567,N_14048);
or U15471 (N_15471,N_11263,N_12947);
or U15472 (N_15472,N_10622,N_14031);
and U15473 (N_15473,N_13106,N_13352);
or U15474 (N_15474,N_14263,N_12103);
or U15475 (N_15475,N_14182,N_12533);
nor U15476 (N_15476,N_10503,N_13288);
or U15477 (N_15477,N_13259,N_14406);
nor U15478 (N_15478,N_12453,N_14424);
and U15479 (N_15479,N_12177,N_12974);
xor U15480 (N_15480,N_14720,N_14539);
nor U15481 (N_15481,N_10696,N_14925);
or U15482 (N_15482,N_13944,N_13730);
xor U15483 (N_15483,N_13842,N_13764);
nor U15484 (N_15484,N_14955,N_12455);
and U15485 (N_15485,N_12285,N_13629);
xnor U15486 (N_15486,N_14583,N_11428);
xor U15487 (N_15487,N_12004,N_13964);
or U15488 (N_15488,N_13651,N_10315);
or U15489 (N_15489,N_11375,N_11300);
and U15490 (N_15490,N_10723,N_10697);
or U15491 (N_15491,N_10281,N_12359);
nand U15492 (N_15492,N_12251,N_13001);
nand U15493 (N_15493,N_13347,N_13996);
or U15494 (N_15494,N_11595,N_13864);
xor U15495 (N_15495,N_12789,N_14340);
nand U15496 (N_15496,N_14853,N_12603);
xor U15497 (N_15497,N_11431,N_10355);
nand U15498 (N_15498,N_10527,N_14619);
xor U15499 (N_15499,N_10716,N_10441);
xnor U15500 (N_15500,N_14238,N_13937);
and U15501 (N_15501,N_13083,N_11179);
or U15502 (N_15502,N_10610,N_12028);
nand U15503 (N_15503,N_10017,N_11778);
nor U15504 (N_15504,N_11387,N_10919);
or U15505 (N_15505,N_14093,N_14961);
nand U15506 (N_15506,N_11983,N_14017);
or U15507 (N_15507,N_12734,N_11276);
and U15508 (N_15508,N_10040,N_12492);
or U15509 (N_15509,N_10390,N_12615);
xnor U15510 (N_15510,N_10436,N_11801);
or U15511 (N_15511,N_13486,N_13900);
nand U15512 (N_15512,N_14599,N_14901);
nor U15513 (N_15513,N_11382,N_11912);
and U15514 (N_15514,N_11747,N_10063);
or U15515 (N_15515,N_13829,N_12888);
or U15516 (N_15516,N_13303,N_11800);
or U15517 (N_15517,N_12112,N_12135);
or U15518 (N_15518,N_10306,N_12968);
nor U15519 (N_15519,N_14478,N_12420);
and U15520 (N_15520,N_11029,N_11910);
or U15521 (N_15521,N_12448,N_13917);
and U15522 (N_15522,N_12027,N_11810);
nor U15523 (N_15523,N_10272,N_14928);
xnor U15524 (N_15524,N_12475,N_13817);
nor U15525 (N_15525,N_11245,N_12051);
and U15526 (N_15526,N_13911,N_10867);
or U15527 (N_15527,N_10835,N_13308);
and U15528 (N_15528,N_13152,N_13994);
and U15529 (N_15529,N_10921,N_11917);
and U15530 (N_15530,N_10752,N_10204);
nand U15531 (N_15531,N_11637,N_13108);
or U15532 (N_15532,N_12815,N_12445);
xnor U15533 (N_15533,N_12526,N_14488);
nor U15534 (N_15534,N_10286,N_14121);
xor U15535 (N_15535,N_11905,N_12561);
nor U15536 (N_15536,N_10330,N_13920);
and U15537 (N_15537,N_14561,N_10205);
and U15538 (N_15538,N_13044,N_12576);
nor U15539 (N_15539,N_13604,N_12437);
and U15540 (N_15540,N_13075,N_10124);
xnor U15541 (N_15541,N_10794,N_12105);
and U15542 (N_15542,N_10741,N_11963);
and U15543 (N_15543,N_11344,N_13223);
nor U15544 (N_15544,N_14115,N_11854);
nand U15545 (N_15545,N_14100,N_12567);
xor U15546 (N_15546,N_13045,N_12025);
nor U15547 (N_15547,N_13581,N_14075);
nor U15548 (N_15548,N_13151,N_11527);
nand U15549 (N_15549,N_14079,N_13506);
xor U15550 (N_15550,N_12849,N_11024);
xor U15551 (N_15551,N_11661,N_13268);
nor U15552 (N_15552,N_12922,N_14728);
and U15553 (N_15553,N_13695,N_14689);
nand U15554 (N_15554,N_14898,N_11765);
or U15555 (N_15555,N_10140,N_13985);
xnor U15556 (N_15556,N_12917,N_13586);
nand U15557 (N_15557,N_11895,N_13806);
and U15558 (N_15558,N_10701,N_13741);
or U15559 (N_15559,N_13424,N_11241);
or U15560 (N_15560,N_11246,N_12872);
and U15561 (N_15561,N_14312,N_14279);
xnor U15562 (N_15562,N_12249,N_11416);
and U15563 (N_15563,N_11842,N_13662);
or U15564 (N_15564,N_13772,N_11021);
xnor U15565 (N_15565,N_14247,N_11541);
xnor U15566 (N_15566,N_12846,N_12286);
nor U15567 (N_15567,N_14886,N_14373);
nor U15568 (N_15568,N_10842,N_13384);
nand U15569 (N_15569,N_13980,N_10283);
and U15570 (N_15570,N_14298,N_14029);
xor U15571 (N_15571,N_13237,N_12466);
or U15572 (N_15572,N_13174,N_12311);
and U15573 (N_15573,N_10702,N_12674);
xor U15574 (N_15574,N_12074,N_11826);
nand U15575 (N_15575,N_12245,N_12429);
nor U15576 (N_15576,N_10207,N_13402);
xor U15577 (N_15577,N_10666,N_11672);
and U15578 (N_15578,N_11434,N_14777);
nor U15579 (N_15579,N_14920,N_13533);
nor U15580 (N_15580,N_10796,N_11009);
nand U15581 (N_15581,N_13319,N_14535);
and U15582 (N_15582,N_12760,N_13104);
or U15583 (N_15583,N_14314,N_13625);
and U15584 (N_15584,N_13611,N_10398);
and U15585 (N_15585,N_13599,N_12587);
xor U15586 (N_15586,N_13247,N_13159);
nor U15587 (N_15587,N_14333,N_10694);
or U15588 (N_15588,N_14227,N_12224);
nor U15589 (N_15589,N_11223,N_14439);
or U15590 (N_15590,N_13903,N_12267);
and U15591 (N_15591,N_11219,N_13385);
nor U15592 (N_15592,N_13346,N_10498);
nor U15593 (N_15593,N_12847,N_13376);
nor U15594 (N_15594,N_10656,N_14808);
or U15595 (N_15595,N_11148,N_12790);
xor U15596 (N_15596,N_10404,N_12722);
and U15597 (N_15597,N_14739,N_14769);
nand U15598 (N_15598,N_10678,N_10517);
and U15599 (N_15599,N_14848,N_10995);
or U15600 (N_15600,N_13119,N_14670);
nor U15601 (N_15601,N_14374,N_14508);
and U15602 (N_15602,N_11037,N_11452);
or U15603 (N_15603,N_10109,N_12290);
and U15604 (N_15604,N_14713,N_10512);
nor U15605 (N_15605,N_11818,N_11485);
and U15606 (N_15606,N_14338,N_11390);
or U15607 (N_15607,N_13078,N_11031);
nor U15608 (N_15608,N_14412,N_11493);
or U15609 (N_15609,N_12649,N_14214);
nor U15610 (N_15610,N_12733,N_11242);
or U15611 (N_15611,N_14975,N_14130);
xor U15612 (N_15612,N_10858,N_11948);
nor U15613 (N_15613,N_10194,N_12293);
nor U15614 (N_15614,N_12834,N_11138);
or U15615 (N_15615,N_13178,N_10427);
xor U15616 (N_15616,N_14683,N_13301);
and U15617 (N_15617,N_11131,N_14727);
xor U15618 (N_15618,N_11721,N_13136);
nand U15619 (N_15619,N_14237,N_13442);
nor U15620 (N_15620,N_10533,N_12853);
or U15621 (N_15621,N_10138,N_12602);
nor U15622 (N_15622,N_11411,N_11592);
nand U15623 (N_15623,N_13388,N_13807);
nand U15624 (N_15624,N_11348,N_11638);
and U15625 (N_15625,N_11357,N_11839);
or U15626 (N_15626,N_11837,N_13287);
or U15627 (N_15627,N_11613,N_10327);
and U15628 (N_15628,N_13869,N_13678);
or U15629 (N_15629,N_10748,N_12162);
nand U15630 (N_15630,N_10961,N_13434);
and U15631 (N_15631,N_12549,N_13470);
nor U15632 (N_15632,N_13093,N_11609);
and U15633 (N_15633,N_10168,N_12648);
nor U15634 (N_15634,N_11073,N_12799);
xnor U15635 (N_15635,N_12393,N_12715);
nand U15636 (N_15636,N_12852,N_10601);
xnor U15637 (N_15637,N_12796,N_13949);
and U15638 (N_15638,N_10225,N_12951);
or U15639 (N_15639,N_11679,N_12141);
and U15640 (N_15640,N_11953,N_14759);
nor U15641 (N_15641,N_10071,N_10971);
nor U15642 (N_15642,N_10452,N_10990);
or U15643 (N_15643,N_13527,N_14528);
xnor U15644 (N_15644,N_10877,N_11574);
or U15645 (N_15645,N_14241,N_12219);
nor U15646 (N_15646,N_13451,N_14144);
nor U15647 (N_15647,N_12246,N_14468);
nor U15648 (N_15648,N_10022,N_14380);
nor U15649 (N_15649,N_12562,N_11466);
nand U15650 (N_15650,N_10211,N_11621);
or U15651 (N_15651,N_10139,N_11849);
or U15652 (N_15652,N_11979,N_13060);
or U15653 (N_15653,N_10302,N_12073);
xor U15654 (N_15654,N_13597,N_12098);
or U15655 (N_15655,N_12204,N_14874);
nand U15656 (N_15656,N_12725,N_12068);
xor U15657 (N_15657,N_13866,N_10846);
and U15658 (N_15658,N_14513,N_11993);
or U15659 (N_15659,N_11711,N_13825);
nor U15660 (N_15660,N_14801,N_14545);
nand U15661 (N_15661,N_11239,N_12376);
xnor U15662 (N_15662,N_13327,N_10857);
and U15663 (N_15663,N_13046,N_13081);
and U15664 (N_15664,N_10460,N_11667);
xor U15665 (N_15665,N_10469,N_10451);
or U15666 (N_15666,N_11270,N_14889);
nor U15667 (N_15667,N_14868,N_11335);
or U15668 (N_15668,N_11685,N_12984);
nand U15669 (N_15669,N_13746,N_11299);
xor U15670 (N_15670,N_11284,N_13717);
xor U15671 (N_15671,N_11674,N_13531);
or U15672 (N_15672,N_14999,N_13593);
and U15673 (N_15673,N_12539,N_10104);
xnor U15674 (N_15674,N_14836,N_13716);
and U15675 (N_15675,N_10636,N_12478);
nand U15676 (N_15676,N_12679,N_10190);
xor U15677 (N_15677,N_14188,N_10761);
and U15678 (N_15678,N_12298,N_14417);
nor U15679 (N_15679,N_10780,N_12818);
nand U15680 (N_15680,N_14260,N_12625);
nand U15681 (N_15681,N_11623,N_11076);
nor U15682 (N_15682,N_14742,N_14261);
and U15683 (N_15683,N_11134,N_13492);
xnor U15684 (N_15684,N_14235,N_11861);
nand U15685 (N_15685,N_13986,N_12008);
xnor U15686 (N_15686,N_12129,N_13579);
and U15687 (N_15687,N_12751,N_13373);
nand U15688 (N_15688,N_13877,N_13366);
or U15689 (N_15689,N_11975,N_11946);
nand U15690 (N_15690,N_11189,N_12814);
nor U15691 (N_15691,N_11279,N_14968);
or U15692 (N_15692,N_11787,N_12840);
nand U15693 (N_15693,N_12510,N_10331);
or U15694 (N_15694,N_10910,N_12971);
nor U15695 (N_15695,N_10082,N_12314);
and U15696 (N_15696,N_10822,N_10814);
nand U15697 (N_15697,N_10077,N_10607);
nand U15698 (N_15698,N_14919,N_14334);
xor U15699 (N_15699,N_12101,N_14810);
nor U15700 (N_15700,N_12498,N_11327);
and U15701 (N_15701,N_13453,N_10983);
and U15702 (N_15702,N_14208,N_12258);
nor U15703 (N_15703,N_10002,N_12200);
or U15704 (N_15704,N_12604,N_13921);
xnor U15705 (N_15705,N_12756,N_14909);
nand U15706 (N_15706,N_13645,N_14699);
nand U15707 (N_15707,N_13239,N_11534);
xor U15708 (N_15708,N_12120,N_13222);
nor U15709 (N_15709,N_13265,N_11738);
nor U15710 (N_15710,N_12343,N_14444);
nand U15711 (N_15711,N_13172,N_11793);
or U15712 (N_15712,N_10003,N_13577);
nand U15713 (N_15713,N_14781,N_10932);
and U15714 (N_15714,N_12779,N_10542);
nand U15715 (N_15715,N_12709,N_10625);
or U15716 (N_15716,N_14865,N_14049);
xnor U15717 (N_15717,N_12348,N_10840);
and U15718 (N_15718,N_10336,N_11569);
and U15719 (N_15719,N_10049,N_12223);
or U15720 (N_15720,N_14534,N_10627);
nor U15721 (N_15721,N_11846,N_11567);
or U15722 (N_15722,N_14726,N_11215);
and U15723 (N_15723,N_11147,N_13941);
nor U15724 (N_15724,N_12797,N_13267);
and U15725 (N_15725,N_14035,N_13711);
or U15726 (N_15726,N_13833,N_13784);
or U15727 (N_15727,N_11994,N_14741);
or U15728 (N_15728,N_14134,N_14358);
xnor U15729 (N_15729,N_10351,N_11474);
nor U15730 (N_15730,N_14885,N_10963);
and U15731 (N_15731,N_14299,N_14197);
nand U15732 (N_15732,N_13144,N_10587);
nand U15733 (N_15733,N_11777,N_12109);
nand U15734 (N_15734,N_11503,N_10440);
and U15735 (N_15735,N_10043,N_12419);
or U15736 (N_15736,N_13087,N_10488);
nand U15737 (N_15737,N_11120,N_14275);
nand U15738 (N_15738,N_10334,N_13014);
or U15739 (N_15739,N_13000,N_11164);
and U15740 (N_15740,N_11886,N_12745);
and U15741 (N_15741,N_11371,N_10812);
nor U15742 (N_15742,N_12991,N_12334);
nor U15743 (N_15743,N_14797,N_11957);
and U15744 (N_15744,N_14493,N_11749);
xor U15745 (N_15745,N_13583,N_14986);
nor U15746 (N_15746,N_10674,N_11713);
or U15747 (N_15747,N_14819,N_13059);
nor U15748 (N_15748,N_11417,N_12485);
or U15749 (N_15749,N_11958,N_11201);
nor U15750 (N_15750,N_13007,N_12700);
and U15751 (N_15751,N_13227,N_11259);
and U15752 (N_15752,N_11980,N_11028);
nand U15753 (N_15753,N_11401,N_11802);
nand U15754 (N_15754,N_12800,N_12713);
nor U15755 (N_15755,N_14128,N_13258);
nor U15756 (N_15756,N_13523,N_13061);
or U15757 (N_15757,N_11132,N_11696);
nor U15758 (N_15758,N_10018,N_14629);
nor U15759 (N_15759,N_10900,N_10938);
xnor U15760 (N_15760,N_14733,N_11785);
or U15761 (N_15761,N_11105,N_14527);
xor U15762 (N_15762,N_11311,N_13255);
xor U15763 (N_15763,N_10637,N_14496);
and U15764 (N_15764,N_14680,N_10212);
nor U15765 (N_15765,N_14179,N_10768);
xnor U15766 (N_15766,N_14542,N_12698);
or U15767 (N_15767,N_13025,N_11186);
and U15768 (N_15768,N_12046,N_14867);
xnor U15769 (N_15769,N_10406,N_11321);
xnor U15770 (N_15770,N_12143,N_12156);
nor U15771 (N_15771,N_10383,N_14166);
and U15772 (N_15772,N_12076,N_14189);
xnor U15773 (N_15773,N_13541,N_11936);
xnor U15774 (N_15774,N_13340,N_12155);
xnor U15775 (N_15775,N_11862,N_11537);
or U15776 (N_15776,N_12973,N_10106);
xor U15777 (N_15777,N_12525,N_12777);
nor U15778 (N_15778,N_13338,N_14011);
or U15779 (N_15779,N_13012,N_11599);
and U15780 (N_15780,N_11727,N_12897);
nor U15781 (N_15781,N_13993,N_13474);
nand U15782 (N_15782,N_12579,N_14143);
nand U15783 (N_15783,N_14410,N_13875);
xor U15784 (N_15784,N_14002,N_11334);
xor U15785 (N_15785,N_10878,N_10013);
and U15786 (N_15786,N_13068,N_12043);
nand U15787 (N_15787,N_14518,N_10308);
nand U15788 (N_15788,N_12421,N_12225);
xnor U15789 (N_15789,N_13297,N_11780);
nor U15790 (N_15790,N_12716,N_11540);
and U15791 (N_15791,N_12032,N_13049);
xor U15792 (N_15792,N_10603,N_11651);
xor U15793 (N_15793,N_10399,N_14022);
nor U15794 (N_15794,N_13380,N_11885);
xnor U15795 (N_15795,N_11393,N_14714);
nand U15796 (N_15796,N_12375,N_10743);
and U15797 (N_15797,N_13663,N_13630);
nor U15798 (N_15798,N_12356,N_10255);
and U15799 (N_15799,N_11562,N_14946);
and U15800 (N_15800,N_10935,N_10191);
and U15801 (N_15801,N_11217,N_12193);
xor U15802 (N_15802,N_12848,N_10776);
or U15803 (N_15803,N_11629,N_13498);
nand U15804 (N_15804,N_12054,N_13126);
and U15805 (N_15805,N_11119,N_13179);
nor U15806 (N_15806,N_14177,N_12699);
nand U15807 (N_15807,N_12599,N_12026);
xnor U15808 (N_15808,N_10374,N_14501);
xnor U15809 (N_15809,N_13411,N_10872);
xnor U15810 (N_15810,N_11732,N_13673);
nor U15811 (N_15811,N_10127,N_13557);
or U15812 (N_15812,N_12605,N_13816);
nand U15813 (N_15813,N_14666,N_12403);
and U15814 (N_15814,N_12415,N_13011);
nand U15815 (N_15815,N_12276,N_14317);
xor U15816 (N_15816,N_11144,N_12755);
and U15817 (N_15817,N_12190,N_12226);
or U15818 (N_15818,N_11369,N_12391);
nand U15819 (N_15819,N_11444,N_14547);
and U15820 (N_15820,N_12596,N_13379);
xnor U15821 (N_15821,N_12978,N_14101);
nor U15822 (N_15822,N_11571,N_13410);
and U15823 (N_15823,N_11928,N_12941);
nor U15824 (N_15824,N_14731,N_10258);
or U15825 (N_15825,N_12010,N_13804);
nand U15826 (N_15826,N_13518,N_14024);
nor U15827 (N_15827,N_11008,N_10731);
and U15828 (N_15828,N_11308,N_12152);
xor U15829 (N_15829,N_10744,N_12993);
xor U15830 (N_15830,N_10590,N_10239);
xnor U15831 (N_15831,N_10725,N_10056);
or U15832 (N_15832,N_12548,N_14078);
nand U15833 (N_15833,N_10329,N_13047);
xnor U15834 (N_15834,N_11524,N_14827);
nor U15835 (N_15835,N_12955,N_12428);
nor U15836 (N_15836,N_11545,N_12981);
or U15837 (N_15837,N_13215,N_14013);
nor U15838 (N_15838,N_11752,N_13830);
or U15839 (N_15839,N_10364,N_10613);
xor U15840 (N_15840,N_14458,N_13646);
nor U15841 (N_15841,N_14644,N_13345);
xnor U15842 (N_15842,N_12378,N_12239);
and U15843 (N_15843,N_11678,N_11570);
nand U15844 (N_15844,N_10798,N_13938);
and U15845 (N_15845,N_12918,N_14829);
xnor U15846 (N_15846,N_10567,N_13196);
and U15847 (N_15847,N_12364,N_10444);
xor U15848 (N_15848,N_13551,N_13861);
nand U15849 (N_15849,N_11960,N_12592);
or U15850 (N_15850,N_11687,N_10998);
or U15851 (N_15851,N_10729,N_14074);
or U15852 (N_15852,N_12115,N_14280);
or U15853 (N_15853,N_14831,N_14738);
xor U15854 (N_15854,N_12529,N_11896);
and U15855 (N_15855,N_13785,N_13289);
and U15856 (N_15856,N_13293,N_14572);
xnor U15857 (N_15857,N_13238,N_14981);
nor U15858 (N_15858,N_13170,N_13064);
nand U15859 (N_15859,N_13652,N_14375);
and U15860 (N_15860,N_11243,N_11671);
or U15861 (N_15861,N_14640,N_13381);
nand U15862 (N_15862,N_13377,N_13808);
xnor U15863 (N_15863,N_12970,N_13706);
and U15864 (N_15864,N_11441,N_10859);
nand U15865 (N_15865,N_12930,N_13787);
xnor U15866 (N_15866,N_13024,N_12336);
or U15867 (N_15867,N_10093,N_13181);
nand U15868 (N_15868,N_14419,N_13003);
nor U15869 (N_15869,N_11136,N_14693);
xnor U15870 (N_15870,N_13831,N_13074);
nor U15871 (N_15871,N_10130,N_14328);
nand U15872 (N_15872,N_13189,N_12367);
or U15873 (N_15873,N_14161,N_13814);
and U15874 (N_15874,N_12838,N_14385);
nor U15875 (N_15875,N_12048,N_10552);
nor U15876 (N_15876,N_11520,N_13507);
xnor U15877 (N_15877,N_14405,N_10700);
or U15878 (N_15878,N_13135,N_13253);
xor U15879 (N_15879,N_10608,N_10405);
nor U15880 (N_15880,N_13568,N_11058);
and U15881 (N_15881,N_12997,N_12831);
nand U15882 (N_15882,N_12014,N_14064);
nor U15883 (N_15883,N_11329,N_12768);
nand U15884 (N_15884,N_13619,N_14751);
or U15885 (N_15885,N_12707,N_11022);
nor U15886 (N_15886,N_11264,N_14361);
nor U15887 (N_15887,N_14442,N_14606);
nor U15888 (N_15888,N_10953,N_12530);
nand U15889 (N_15889,N_10915,N_10471);
and U15890 (N_15890,N_10661,N_12134);
xor U15891 (N_15891,N_14620,N_10767);
nand U15892 (N_15892,N_13466,N_13006);
nand U15893 (N_15893,N_10321,N_12845);
nand U15894 (N_15894,N_13729,N_13737);
or U15895 (N_15895,N_12154,N_12145);
nor U15896 (N_15896,N_14449,N_12730);
xor U15897 (N_15897,N_12837,N_13363);
nor U15898 (N_15898,N_12240,N_13101);
nor U15899 (N_15899,N_13386,N_10318);
or U15900 (N_15900,N_11544,N_13931);
nor U15901 (N_15901,N_11269,N_11090);
xnor U15902 (N_15902,N_11454,N_11235);
xnor U15903 (N_15903,N_14415,N_13306);
nor U15904 (N_15904,N_14926,N_10247);
and U15905 (N_15905,N_11646,N_13212);
nand U15906 (N_15906,N_13952,N_12950);
nand U15907 (N_15907,N_11551,N_14736);
and U15908 (N_15908,N_12940,N_13062);
nor U15909 (N_15909,N_13946,N_12695);
nand U15910 (N_15910,N_10526,N_10486);
xor U15911 (N_15911,N_10403,N_13691);
nor U15912 (N_15912,N_10123,N_13398);
and U15913 (N_15913,N_10249,N_14402);
and U15914 (N_15914,N_12560,N_12923);
and U15915 (N_15915,N_11563,N_13649);
nor U15916 (N_15916,N_10907,N_13661);
or U15917 (N_15917,N_13089,N_10447);
or U15918 (N_15918,N_11518,N_11192);
nand U15919 (N_15919,N_13446,N_11779);
and U15920 (N_15920,N_10726,N_12969);
nor U15921 (N_15921,N_12338,N_14916);
nor U15922 (N_15922,N_14211,N_11437);
and U15923 (N_15923,N_10540,N_14289);
and U15924 (N_15924,N_14370,N_10048);
or U15925 (N_15925,N_11624,N_14617);
or U15926 (N_15926,N_12601,N_13686);
and U15927 (N_15927,N_13508,N_14596);
nor U15928 (N_15928,N_14117,N_10473);
nor U15929 (N_15929,N_12925,N_12839);
or U15930 (N_15930,N_11568,N_11425);
and U15931 (N_15931,N_11365,N_13153);
and U15932 (N_15932,N_14813,N_14549);
or U15933 (N_15933,N_11769,N_12044);
nor U15934 (N_15934,N_13591,N_14369);
and U15935 (N_15935,N_13030,N_14015);
nand U15936 (N_15936,N_10060,N_13659);
and U15937 (N_15937,N_14336,N_13478);
nor U15938 (N_15938,N_10997,N_12773);
xnor U15939 (N_15939,N_13522,N_10930);
nor U15940 (N_15940,N_11633,N_11469);
and U15941 (N_15941,N_14990,N_11889);
nand U15942 (N_15942,N_12362,N_10889);
and U15943 (N_15943,N_12373,N_14983);
or U15944 (N_15944,N_14321,N_11410);
and U15945 (N_15945,N_11255,N_11536);
nand U15946 (N_15946,N_10711,N_10933);
nand U15947 (N_15947,N_11751,N_13837);
nand U15948 (N_15948,N_11038,N_13110);
and U15949 (N_15949,N_10006,N_12064);
nand U15950 (N_15950,N_11165,N_11554);
nand U15951 (N_15951,N_10409,N_10032);
and U15952 (N_15952,N_10522,N_11498);
nand U15953 (N_15953,N_10596,N_13286);
nand U15954 (N_15954,N_10322,N_10787);
or U15955 (N_15955,N_11996,N_11354);
and U15956 (N_15956,N_12854,N_12332);
xor U15957 (N_15957,N_10880,N_14891);
nand U15958 (N_15958,N_10320,N_10416);
and U15959 (N_15959,N_14181,N_13382);
xnor U15960 (N_15960,N_13283,N_11677);
or U15961 (N_15961,N_10449,N_13133);
and U15962 (N_15962,N_10591,N_13019);
nor U15963 (N_15963,N_10651,N_10792);
and U15964 (N_15964,N_13575,N_13473);
or U15965 (N_15965,N_11035,N_10739);
and U15966 (N_15966,N_13965,N_13270);
or U15967 (N_15967,N_12622,N_10539);
or U15968 (N_15968,N_10005,N_13173);
and U15969 (N_15969,N_11491,N_12021);
nand U15970 (N_15970,N_12914,N_13997);
nand U15971 (N_15971,N_13143,N_13362);
and U15972 (N_15972,N_13566,N_14165);
or U15973 (N_15973,N_14414,N_14348);
nand U15974 (N_15974,N_10852,N_11345);
xor U15975 (N_15975,N_14543,N_14300);
and U15976 (N_15976,N_12148,N_10100);
nand U15977 (N_15977,N_10618,N_10516);
xor U15978 (N_15978,N_13562,N_11251);
or U15979 (N_15979,N_11740,N_11606);
xor U15980 (N_15980,N_14112,N_14382);
nand U15981 (N_15981,N_10357,N_13760);
nor U15982 (N_15982,N_11438,N_10894);
nor U15983 (N_15983,N_10885,N_14012);
or U15984 (N_15984,N_12572,N_12802);
or U15985 (N_15985,N_14339,N_10747);
xnor U15986 (N_15986,N_13169,N_14005);
or U15987 (N_15987,N_10346,N_14344);
and U15988 (N_15988,N_13558,N_14950);
xor U15989 (N_15989,N_14722,N_13282);
and U15990 (N_15990,N_11271,N_10562);
or U15991 (N_15991,N_13820,N_10348);
nand U15992 (N_15992,N_11071,N_14277);
and U15993 (N_15993,N_10149,N_14418);
and U15994 (N_15994,N_13218,N_10262);
nor U15995 (N_15995,N_13331,N_10224);
or U15996 (N_15996,N_11277,N_11230);
xor U15997 (N_15997,N_11585,N_11408);
nor U15998 (N_15998,N_14009,N_13021);
nand U15999 (N_15999,N_11603,N_12903);
or U16000 (N_16000,N_12759,N_12683);
and U16001 (N_16001,N_13339,N_10265);
xnor U16002 (N_16002,N_14567,N_11018);
or U16003 (N_16003,N_13862,N_11377);
nand U16004 (N_16004,N_11742,N_13191);
and U16005 (N_16005,N_14394,N_11126);
and U16006 (N_16006,N_10824,N_10428);
nand U16007 (N_16007,N_14911,N_14517);
xor U16008 (N_16008,N_13694,N_11987);
and U16009 (N_16009,N_11774,N_12781);
nor U16010 (N_16010,N_12618,N_11197);
and U16011 (N_16011,N_11402,N_10037);
or U16012 (N_16012,N_13503,N_12532);
xor U16013 (N_16013,N_13273,N_11092);
nand U16014 (N_16014,N_11648,N_13107);
or U16015 (N_16015,N_14877,N_11507);
nor U16016 (N_16016,N_11169,N_10604);
xnor U16017 (N_16017,N_13519,N_14799);
nor U16018 (N_16018,N_13958,N_12542);
or U16019 (N_16019,N_13640,N_10808);
nand U16020 (N_16020,N_12000,N_13284);
nor U16021 (N_16021,N_14992,N_10196);
or U16022 (N_16022,N_12929,N_12992);
xnor U16023 (N_16023,N_10886,N_13916);
and U16024 (N_16024,N_11060,N_11788);
nand U16025 (N_16025,N_13767,N_12110);
xor U16026 (N_16026,N_13525,N_10970);
nand U16027 (N_16027,N_13821,N_14724);
nor U16028 (N_16028,N_14236,N_14793);
xnor U16029 (N_16029,N_13848,N_12915);
nand U16030 (N_16030,N_13854,N_10242);
nand U16031 (N_16031,N_11280,N_12563);
and U16032 (N_16032,N_11487,N_14735);
xor U16033 (N_16033,N_13360,N_12365);
xor U16034 (N_16034,N_12600,N_12876);
and U16035 (N_16035,N_13844,N_14597);
or U16036 (N_16036,N_11079,N_11597);
xnor U16037 (N_16037,N_12252,N_12647);
nor U16038 (N_16038,N_14524,N_10119);
or U16039 (N_16039,N_12483,N_12088);
nor U16040 (N_16040,N_12544,N_12176);
nor U16041 (N_16041,N_11775,N_14495);
and U16042 (N_16042,N_13563,N_12360);
and U16043 (N_16043,N_13278,N_13845);
nand U16044 (N_16044,N_12666,N_13175);
nand U16045 (N_16045,N_11874,N_10266);
or U16046 (N_16046,N_14631,N_10564);
nand U16047 (N_16047,N_14980,N_14404);
xnor U16048 (N_16048,N_13967,N_11257);
and U16049 (N_16049,N_14873,N_12195);
and U16050 (N_16050,N_12911,N_14267);
or U16051 (N_16051,N_14580,N_11059);
or U16052 (N_16052,N_10382,N_11112);
and U16053 (N_16053,N_11891,N_10578);
and U16054 (N_16054,N_13623,N_10721);
xor U16055 (N_16055,N_14952,N_10023);
nand U16056 (N_16056,N_12608,N_12610);
or U16057 (N_16057,N_11640,N_10710);
xor U16058 (N_16058,N_14127,N_14205);
xor U16059 (N_16059,N_10101,N_14672);
and U16060 (N_16060,N_11578,N_12633);
and U16061 (N_16061,N_10777,N_12326);
or U16062 (N_16062,N_10510,N_14563);
xor U16063 (N_16063,N_10021,N_13018);
and U16064 (N_16064,N_12191,N_11228);
nand U16065 (N_16065,N_10227,N_11806);
or U16066 (N_16066,N_11868,N_14210);
or U16067 (N_16067,N_10905,N_14061);
nor U16068 (N_16068,N_10860,N_10052);
and U16069 (N_16069,N_14965,N_10541);
or U16070 (N_16070,N_13418,N_14668);
nor U16071 (N_16071,N_12199,N_14000);
xnor U16072 (N_16072,N_14600,N_13876);
nand U16073 (N_16073,N_11000,N_11432);
nor U16074 (N_16074,N_12468,N_13325);
nor U16075 (N_16075,N_13165,N_14451);
or U16076 (N_16076,N_10538,N_10016);
or U16077 (N_16077,N_10443,N_10232);
nand U16078 (N_16078,N_12757,N_14390);
or U16079 (N_16079,N_10407,N_12142);
nand U16080 (N_16080,N_11670,N_11011);
or U16081 (N_16081,N_14771,N_13026);
or U16082 (N_16082,N_11343,N_10344);
or U16083 (N_16083,N_13121,N_10027);
xnor U16084 (N_16084,N_12462,N_14622);
or U16085 (N_16085,N_11662,N_13210);
nand U16086 (N_16086,N_12945,N_12890);
and U16087 (N_16087,N_12861,N_13757);
xnor U16088 (N_16088,N_12642,N_13536);
or U16089 (N_16089,N_13233,N_13858);
or U16090 (N_16090,N_13849,N_10116);
nand U16091 (N_16091,N_14162,N_13219);
nor U16092 (N_16092,N_14187,N_10683);
and U16093 (N_16093,N_12006,N_10574);
nor U16094 (N_16094,N_13601,N_12408);
or U16095 (N_16095,N_10906,N_10141);
and U16096 (N_16096,N_13435,N_14960);
xnor U16097 (N_16097,N_12597,N_10942);
or U16098 (N_16098,N_10384,N_11761);
nor U16099 (N_16099,N_13291,N_11322);
nand U16100 (N_16100,N_10387,N_13643);
nand U16101 (N_16101,N_13356,N_11155);
nor U16102 (N_16102,N_13040,N_13130);
and U16103 (N_16103,N_14805,N_11319);
xnor U16104 (N_16104,N_10866,N_13647);
and U16105 (N_16105,N_13404,N_13469);
nor U16106 (N_16106,N_13053,N_12097);
or U16107 (N_16107,N_11641,N_10501);
nand U16108 (N_16108,N_13266,N_10304);
nand U16109 (N_16109,N_12731,N_13948);
nand U16110 (N_16110,N_13439,N_10111);
nand U16111 (N_16111,N_13073,N_13860);
or U16112 (N_16112,N_14562,N_11298);
nand U16113 (N_16113,N_13756,N_11626);
or U16114 (N_16114,N_14335,N_14122);
nand U16115 (N_16115,N_12291,N_11853);
or U16116 (N_16116,N_12764,N_14746);
and U16117 (N_16117,N_14665,N_10616);
xor U16118 (N_16118,N_11128,N_13187);
xnor U16119 (N_16119,N_12708,N_10766);
or U16120 (N_16120,N_11781,N_13835);
nand U16121 (N_16121,N_10221,N_10827);
and U16122 (N_16122,N_10864,N_14073);
xor U16123 (N_16123,N_13809,N_13521);
nand U16124 (N_16124,N_10759,N_13312);
and U16125 (N_16125,N_11753,N_14428);
xor U16126 (N_16126,N_10871,N_12901);
nor U16127 (N_16127,N_11591,N_12341);
or U16128 (N_16128,N_14092,N_11483);
xor U16129 (N_16129,N_14060,N_12864);
or U16130 (N_16130,N_14228,N_12537);
nand U16131 (N_16131,N_14034,N_13744);
or U16132 (N_16132,N_11445,N_11937);
xnor U16133 (N_16133,N_10087,N_10925);
or U16134 (N_16134,N_11106,N_13872);
nor U16135 (N_16135,N_13272,N_13897);
nand U16136 (N_16136,N_14812,N_14480);
xor U16137 (N_16137,N_13798,N_11684);
nand U16138 (N_16138,N_10163,N_12939);
nand U16139 (N_16139,N_13930,N_11418);
xor U16140 (N_16140,N_13749,N_12377);
xnor U16141 (N_16141,N_11463,N_14674);
nor U16142 (N_16142,N_12201,N_13394);
xor U16143 (N_16143,N_14807,N_11682);
xnor U16144 (N_16144,N_14559,N_13020);
nand U16145 (N_16145,N_13868,N_12780);
xnor U16146 (N_16146,N_12385,N_10370);
nor U16147 (N_16147,N_12664,N_12546);
and U16148 (N_16148,N_13224,N_10848);
or U16149 (N_16149,N_10789,N_10605);
nor U16150 (N_16150,N_10342,N_10263);
xor U16151 (N_16151,N_11221,N_14521);
nor U16152 (N_16152,N_13199,N_14837);
xor U16153 (N_16153,N_14499,N_14880);
and U16154 (N_16154,N_13576,N_13618);
nor U16155 (N_16155,N_14190,N_11301);
nand U16156 (N_16156,N_14630,N_14086);
and U16157 (N_16157,N_11368,N_14783);
nor U16158 (N_16158,N_13364,N_10195);
or U16159 (N_16159,N_11433,N_13341);
or U16160 (N_16160,N_10934,N_11360);
or U16161 (N_16161,N_12208,N_12611);
xor U16162 (N_16162,N_14687,N_10620);
and U16163 (N_16163,N_12318,N_12502);
xnor U16164 (N_16164,N_10675,N_14634);
nor U16165 (N_16165,N_14147,N_10670);
and U16166 (N_16166,N_11604,N_11361);
xnor U16167 (N_16167,N_11840,N_13698);
or U16168 (N_16168,N_10650,N_10941);
and U16169 (N_16169,N_13505,N_13617);
xor U16170 (N_16170,N_10582,N_13995);
nor U16171 (N_16171,N_10237,N_11500);
nor U16172 (N_16172,N_14149,N_14984);
nor U16173 (N_16173,N_12328,N_10036);
nand U16174 (N_16174,N_12913,N_10939);
xnor U16175 (N_16175,N_11383,N_14764);
nor U16176 (N_16176,N_11209,N_13109);
nor U16177 (N_16177,N_11576,N_14329);
nand U16178 (N_16178,N_13177,N_12128);
nand U16179 (N_16179,N_10347,N_14794);
or U16180 (N_16180,N_11878,N_11601);
nand U16181 (N_16181,N_12146,N_14884);
nand U16182 (N_16182,N_10928,N_13656);
nand U16183 (N_16183,N_13681,N_10259);
and U16184 (N_16184,N_13350,N_14972);
or U16185 (N_16185,N_14084,N_13580);
nor U16186 (N_16186,N_12659,N_11619);
xnor U16187 (N_16187,N_11475,N_13079);
xor U16188 (N_16188,N_12865,N_10592);
nand U16189 (N_16189,N_12259,N_11893);
nor U16190 (N_16190,N_12480,N_12684);
nand U16191 (N_16191,N_13968,N_13628);
or U16192 (N_16192,N_14822,N_10665);
and U16193 (N_16193,N_12720,N_12686);
or U16194 (N_16194,N_13146,N_11262);
nor U16195 (N_16195,N_11317,N_12275);
or U16196 (N_16196,N_10920,N_12444);
and U16197 (N_16197,N_14685,N_12299);
nor U16198 (N_16198,N_12052,N_12476);
or U16199 (N_16199,N_14021,N_11838);
or U16200 (N_16200,N_10375,N_11468);
and U16201 (N_16201,N_11940,N_13524);
nor U16202 (N_16202,N_11414,N_12710);
and U16203 (N_16203,N_10754,N_11590);
xnor U16204 (N_16204,N_11039,N_12122);
nor U16205 (N_16205,N_10784,N_14220);
nand U16206 (N_16206,N_11884,N_13671);
xor U16207 (N_16207,N_14087,N_14989);
or U16208 (N_16208,N_13048,N_12205);
and U16209 (N_16209,N_10569,N_14949);
and U16210 (N_16210,N_14913,N_12277);
and U16211 (N_16211,N_11988,N_10545);
and U16212 (N_16212,N_13553,N_14063);
nor U16213 (N_16213,N_10668,N_14413);
nand U16214 (N_16214,N_13797,N_14938);
or U16215 (N_16215,N_14702,N_13117);
xnor U16216 (N_16216,N_11281,N_11790);
xnor U16217 (N_16217,N_12966,N_11879);
and U16218 (N_16218,N_12036,N_10185);
or U16219 (N_16219,N_11748,N_11274);
xor U16220 (N_16220,N_14560,N_11351);
nor U16221 (N_16221,N_13548,N_11415);
xor U16222 (N_16222,N_12137,N_13865);
nand U16223 (N_16223,N_10641,N_12851);
nand U16224 (N_16224,N_14224,N_12889);
or U16225 (N_16225,N_14386,N_14749);
xor U16226 (N_16226,N_12456,N_14800);
nor U16227 (N_16227,N_11152,N_10936);
nor U16228 (N_16228,N_10619,N_12322);
xnor U16229 (N_16229,N_13783,N_13762);
or U16230 (N_16230,N_11959,N_14628);
xnor U16231 (N_16231,N_14830,N_13408);
or U16232 (N_16232,N_11798,N_12556);
or U16233 (N_16233,N_10662,N_14638);
nand U16234 (N_16234,N_12352,N_13983);
xnor U16235 (N_16235,N_14732,N_14231);
and U16236 (N_16236,N_10660,N_13606);
or U16237 (N_16237,N_13669,N_11240);
xnor U16238 (N_16238,N_10046,N_11166);
nand U16239 (N_16239,N_14036,N_14595);
and U16240 (N_16240,N_10514,N_14198);
and U16241 (N_16241,N_11584,N_10576);
nor U16242 (N_16242,N_14088,N_11706);
xor U16243 (N_16243,N_12117,N_14605);
nor U16244 (N_16244,N_12626,N_14353);
or U16245 (N_16245,N_14355,N_11660);
nand U16246 (N_16246,N_12087,N_13824);
and U16247 (N_16247,N_10952,N_12912);
xnor U16248 (N_16248,N_13763,N_11949);
or U16249 (N_16249,N_12820,N_12932);
xor U16250 (N_16250,N_13812,N_10724);
or U16251 (N_16251,N_11693,N_13752);
or U16252 (N_16252,N_11234,N_13416);
nand U16253 (N_16253,N_14293,N_13023);
nor U16254 (N_16254,N_11095,N_14657);
and U16255 (N_16255,N_11014,N_10069);
nand U16256 (N_16256,N_10635,N_10693);
and U16257 (N_16257,N_13912,N_13274);
nand U16258 (N_16258,N_10775,N_13493);
nor U16259 (N_16259,N_12234,N_10821);
xnor U16260 (N_16260,N_12196,N_12900);
or U16261 (N_16261,N_10065,N_12013);
and U16262 (N_16262,N_13100,N_13779);
and U16263 (N_16263,N_11888,N_12149);
nor U16264 (N_16264,N_13839,N_12586);
or U16265 (N_16265,N_12093,N_12427);
xnor U16266 (N_16266,N_13425,N_14356);
xnor U16267 (N_16267,N_10340,N_11535);
or U16268 (N_16268,N_10278,N_14467);
nor U16269 (N_16269,N_11697,N_10319);
and U16270 (N_16270,N_11981,N_10508);
or U16271 (N_16271,N_13532,N_12107);
or U16272 (N_16272,N_10493,N_13433);
nand U16273 (N_16273,N_11016,N_11924);
nor U16274 (N_16274,N_13755,N_14875);
nand U16275 (N_16275,N_13991,N_14448);
nand U16276 (N_16276,N_13092,N_11851);
or U16277 (N_16277,N_10819,N_14199);
or U16278 (N_16278,N_14221,N_11724);
xor U16279 (N_16279,N_10598,N_10594);
and U16280 (N_16280,N_14933,N_10270);
nand U16281 (N_16281,N_11968,N_12289);
and U16282 (N_16282,N_13037,N_12121);
xnor U16283 (N_16283,N_10029,N_12640);
xnor U16284 (N_16284,N_11731,N_14327);
or U16285 (N_16285,N_10388,N_14303);
or U16286 (N_16286,N_10957,N_11044);
nand U16287 (N_16287,N_12826,N_12344);
nand U16288 (N_16288,N_13359,N_11522);
nor U16289 (N_16289,N_14643,N_10155);
or U16290 (N_16290,N_11509,N_12965);
or U16291 (N_16291,N_11077,N_12828);
or U16292 (N_16292,N_14878,N_10042);
nor U16293 (N_16293,N_12696,N_14934);
nand U16294 (N_16294,N_13467,N_10612);
and U16295 (N_16295,N_12558,N_13981);
nor U16296 (N_16296,N_11473,N_10908);
or U16297 (N_16297,N_13928,N_13544);
or U16298 (N_16298,N_13602,N_14194);
nand U16299 (N_16299,N_14173,N_11464);
nand U16300 (N_16300,N_12643,N_10914);
xnor U16301 (N_16301,N_11135,N_14785);
or U16302 (N_16302,N_13491,N_10313);
nor U16303 (N_16303,N_11519,N_13090);
and U16304 (N_16304,N_11154,N_12859);
or U16305 (N_16305,N_10170,N_12136);
nor U16306 (N_16306,N_10126,N_11964);
nor U16307 (N_16307,N_13769,N_14948);
nor U16308 (N_16308,N_12809,N_11180);
xnor U16309 (N_16309,N_14429,N_10543);
nand U16310 (N_16310,N_10220,N_10950);
nor U16311 (N_16311,N_11941,N_14658);
nor U16312 (N_16312,N_10252,N_12182);
and U16313 (N_16313,N_10638,N_10431);
and U16314 (N_16314,N_10948,N_10689);
nand U16315 (N_16315,N_13511,N_12687);
and U16316 (N_16316,N_14094,N_14245);
or U16317 (N_16317,N_13307,N_11455);
nand U16318 (N_16318,N_14698,N_12748);
nor U16319 (N_16319,N_14053,N_13736);
nand U16320 (N_16320,N_13088,N_11034);
xor U16321 (N_16321,N_14809,N_13904);
and U16322 (N_16322,N_12055,N_14632);
xnor U16323 (N_16323,N_13256,N_12487);
and U16324 (N_16324,N_10031,N_10671);
xnor U16325 (N_16325,N_10714,N_10341);
and U16326 (N_16326,N_11130,N_11213);
xor U16327 (N_16327,N_12938,N_13502);
or U16328 (N_16328,N_12776,N_12825);
or U16329 (N_16329,N_13276,N_14618);
and U16330 (N_16330,N_14861,N_13125);
nor U16331 (N_16331,N_14054,N_11096);
and U16332 (N_16332,N_10241,N_14707);
nand U16333 (N_16333,N_10389,N_12880);
and U16334 (N_16334,N_10911,N_13017);
xnor U16335 (N_16335,N_14233,N_10236);
and U16336 (N_16336,N_12379,N_11596);
nand U16337 (N_16337,N_12850,N_11350);
nand U16338 (N_16338,N_11049,N_13962);
or U16339 (N_16339,N_14765,N_10437);
nor U16340 (N_16340,N_11292,N_10996);
or U16341 (N_16341,N_14681,N_10188);
nor U16342 (N_16342,N_10581,N_11462);
xnor U16343 (N_16343,N_12307,N_10537);
and U16344 (N_16344,N_12423,N_13664);
nor U16345 (N_16345,N_12841,N_13148);
nor U16346 (N_16346,N_11353,N_12150);
nor U16347 (N_16347,N_10142,N_13790);
and U16348 (N_16348,N_14027,N_13440);
xnor U16349 (N_16349,N_12001,N_10565);
xor U16350 (N_16350,N_13696,N_12769);
and U16351 (N_16351,N_14360,N_13069);
or U16352 (N_16352,N_10799,N_13387);
xor U16353 (N_16353,N_12473,N_13372);
nor U16354 (N_16354,N_11033,N_11081);
or U16355 (N_16355,N_14856,N_14453);
and U16356 (N_16356,N_13932,N_12857);
nor U16357 (N_16357,N_13137,N_10125);
nor U16358 (N_16358,N_13460,N_14098);
and U16359 (N_16359,N_12860,N_11064);
or U16360 (N_16360,N_14729,N_13582);
nor U16361 (N_16361,N_11244,N_13436);
nand U16362 (N_16362,N_11307,N_12069);
nand U16363 (N_16363,N_10088,N_10260);
or U16364 (N_16364,N_12102,N_12738);
xor U16365 (N_16365,N_11550,N_13220);
nand U16366 (N_16366,N_13886,N_10861);
nand U16367 (N_16367,N_10038,N_14274);
or U16368 (N_16368,N_10655,N_11400);
nor U16369 (N_16369,N_10691,N_13468);
xnor U16370 (N_16370,N_12726,N_13043);
nand U16371 (N_16371,N_11627,N_13343);
nand U16372 (N_16372,N_11268,N_14890);
and U16373 (N_16373,N_12075,N_10075);
or U16374 (N_16374,N_13230,N_14363);
nor U16375 (N_16375,N_11548,N_14246);
or U16376 (N_16376,N_11015,N_13834);
xor U16377 (N_16377,N_12108,N_12323);
xor U16378 (N_16378,N_14400,N_14820);
or U16379 (N_16379,N_14490,N_11104);
xor U16380 (N_16380,N_10940,N_13248);
xor U16381 (N_16381,N_12382,N_14503);
nand U16382 (N_16382,N_14633,N_14159);
and U16383 (N_16383,N_14248,N_12928);
or U16384 (N_16384,N_14931,N_13672);
nand U16385 (N_16385,N_12209,N_10999);
and U16386 (N_16386,N_12147,N_13084);
xnor U16387 (N_16387,N_12676,N_11722);
and U16388 (N_16388,N_11863,N_14288);
nor U16389 (N_16389,N_12580,N_11010);
or U16390 (N_16390,N_11358,N_14939);
and U16391 (N_16391,N_14588,N_13631);
nor U16392 (N_16392,N_10296,N_12703);
nand U16393 (N_16393,N_10816,N_13613);
xor U16394 (N_16394,N_10810,N_12458);
xnor U16395 (N_16395,N_11185,N_14715);
nor U16396 (N_16396,N_13251,N_13111);
or U16397 (N_16397,N_10072,N_14007);
and U16398 (N_16398,N_10433,N_10649);
nor U16399 (N_16399,N_11630,N_14664);
nand U16400 (N_16400,N_12380,N_14253);
nand U16401 (N_16401,N_13535,N_13700);
and U16402 (N_16402,N_11330,N_11032);
nand U16403 (N_16403,N_14760,N_13269);
or U16404 (N_16404,N_13290,N_11085);
xor U16405 (N_16405,N_14953,N_13960);
xnor U16406 (N_16406,N_10972,N_13827);
nor U16407 (N_16407,N_14756,N_11962);
nor U16408 (N_16408,N_10234,N_13571);
nand U16409 (N_16409,N_13463,N_11617);
nor U16410 (N_16410,N_10083,N_13141);
or U16411 (N_16411,N_10475,N_14550);
xnor U16412 (N_16412,N_12694,N_12018);
or U16413 (N_16413,N_13225,N_11061);
or U16414 (N_16414,N_11293,N_11025);
xnor U16415 (N_16415,N_13972,N_10969);
and U16416 (N_16416,N_12591,N_13138);
or U16417 (N_16417,N_13342,N_11530);
nand U16418 (N_16418,N_14997,N_14352);
nor U16419 (N_16419,N_10815,N_11355);
and U16420 (N_16420,N_14757,N_14447);
or U16421 (N_16421,N_14016,N_10708);
xor U16422 (N_16422,N_12680,N_14688);
nor U16423 (N_16423,N_10231,N_10630);
and U16424 (N_16424,N_11817,N_11542);
nand U16425 (N_16425,N_12157,N_14761);
nand U16426 (N_16426,N_10899,N_10011);
or U16427 (N_16427,N_12389,N_13873);
and U16428 (N_16428,N_14915,N_11205);
and U16429 (N_16429,N_14018,N_12060);
and U16430 (N_16430,N_11642,N_11883);
nor U16431 (N_16431,N_13731,N_12617);
and U16432 (N_16432,N_10463,N_13096);
xor U16433 (N_16433,N_13605,N_10358);
nor U16434 (N_16434,N_11645,N_11460);
xor U16435 (N_16435,N_12250,N_12524);
xnor U16436 (N_16436,N_12805,N_10621);
and U16437 (N_16437,N_11181,N_11611);
or U16438 (N_16438,N_12358,N_14171);
nor U16439 (N_16439,N_13004,N_13596);
or U16440 (N_16440,N_14870,N_10487);
or U16441 (N_16441,N_12675,N_13777);
xor U16442 (N_16442,N_12396,N_13396);
nor U16443 (N_16443,N_11746,N_11388);
xnor U16444 (N_16444,N_14249,N_10184);
or U16445 (N_16445,N_11212,N_13637);
xnor U16446 (N_16446,N_13353,N_10261);
nor U16447 (N_16447,N_14250,N_14612);
or U16448 (N_16448,N_11143,N_12575);
nor U16449 (N_16449,N_11019,N_11612);
nor U16450 (N_16450,N_11822,N_11556);
xnor U16451 (N_16451,N_13415,N_11156);
nor U16452 (N_16452,N_14876,N_11342);
nand U16453 (N_16453,N_14310,N_10435);
nand U16454 (N_16454,N_14608,N_12130);
or U16455 (N_16455,N_11379,N_12413);
nand U16456 (N_16456,N_11439,N_14072);
and U16457 (N_16457,N_12400,N_12824);
or U16458 (N_16458,N_12541,N_11347);
xor U16459 (N_16459,N_10091,N_13725);
nand U16460 (N_16460,N_12771,N_14457);
nand U16461 (N_16461,N_11188,N_10732);
xor U16462 (N_16462,N_12555,N_10132);
nand U16463 (N_16463,N_14244,N_11786);
nand U16464 (N_16464,N_12569,N_11945);
xor U16465 (N_16465,N_14286,N_11974);
nor U16466 (N_16466,N_12899,N_14838);
xnor U16467 (N_16467,N_11510,N_10098);
xor U16468 (N_16468,N_14089,N_13457);
or U16469 (N_16469,N_14285,N_14850);
and U16470 (N_16470,N_14507,N_11492);
and U16471 (N_16471,N_12653,N_10080);
nor U16472 (N_16472,N_12470,N_14795);
and U16473 (N_16473,N_13899,N_11002);
xnor U16474 (N_16474,N_12843,N_14176);
or U16475 (N_16475,N_11750,N_11087);
nand U16476 (N_16476,N_14494,N_11012);
or U16477 (N_16477,N_11170,N_11146);
xor U16478 (N_16478,N_12056,N_10396);
nor U16479 (N_16479,N_10553,N_11297);
and U16480 (N_16480,N_13271,N_10737);
and U16481 (N_16481,N_11389,N_13234);
or U16482 (N_16482,N_13555,N_10980);
xnor U16483 (N_16483,N_14581,N_12736);
or U16484 (N_16484,N_11392,N_12426);
nand U16485 (N_16485,N_11407,N_14954);
nor U16486 (N_16486,N_12527,N_12998);
xor U16487 (N_16487,N_14239,N_10504);
xor U16488 (N_16488,N_11458,N_12588);
and U16489 (N_16489,N_10699,N_11250);
nor U16490 (N_16490,N_10733,N_14625);
or U16491 (N_16491,N_12657,N_14043);
or U16492 (N_16492,N_13843,N_12390);
nand U16493 (N_16493,N_14826,N_13636);
nand U16494 (N_16494,N_10251,N_12994);
nor U16495 (N_16495,N_12832,N_13727);
and U16496 (N_16496,N_11566,N_10483);
or U16497 (N_16497,N_13517,N_10895);
or U16498 (N_16498,N_13933,N_12003);
nor U16499 (N_16499,N_10834,N_11655);
nand U16500 (N_16500,N_13701,N_12632);
nand U16501 (N_16501,N_12454,N_14671);
nor U16502 (N_16502,N_13479,N_13898);
or U16503 (N_16503,N_12528,N_12654);
and U16504 (N_16504,N_13822,N_10797);
nand U16505 (N_16505,N_14930,N_13679);
nand U16506 (N_16506,N_14896,N_11639);
and U16507 (N_16507,N_12035,N_12517);
or U16508 (N_16508,N_10253,N_10746);
and U16509 (N_16509,N_14226,N_11074);
nor U16510 (N_16510,N_12355,N_13674);
xor U16511 (N_16511,N_14056,N_13245);
and U16512 (N_16512,N_10628,N_14175);
or U16513 (N_16513,N_14734,N_11409);
nand U16514 (N_16514,N_13539,N_12181);
and U16515 (N_16515,N_10411,N_13122);
and U16516 (N_16516,N_14532,N_11698);
nor U16517 (N_16517,N_11632,N_13176);
nand U16518 (N_16518,N_13758,N_10362);
nor U16519 (N_16519,N_12418,N_11908);
xor U16520 (N_16520,N_14240,N_12902);
nand U16521 (N_16521,N_12159,N_13472);
xor U16522 (N_16522,N_10634,N_13036);
xnor U16523 (N_16523,N_13441,N_11723);
xnor U16524 (N_16524,N_10053,N_14163);
nor U16525 (N_16525,N_13094,N_13420);
or U16526 (N_16526,N_13127,N_10913);
and U16527 (N_16527,N_12278,N_11644);
or U16528 (N_16528,N_12179,N_11287);
and U16529 (N_16529,N_12995,N_12628);
nor U16530 (N_16530,N_10378,N_14452);
nand U16531 (N_16531,N_10609,N_11479);
and U16532 (N_16532,N_14434,N_10470);
nor U16533 (N_16533,N_12867,N_12292);
nor U16534 (N_16534,N_14262,N_12086);
and U16535 (N_16535,N_11841,N_13978);
or U16536 (N_16536,N_13456,N_10202);
nor U16537 (N_16537,N_12479,N_14969);
nand U16538 (N_16538,N_10982,N_10988);
nand U16539 (N_16539,N_14821,N_14425);
nand U16540 (N_16540,N_13063,N_13438);
or U16541 (N_16541,N_10688,N_11927);
nand U16542 (N_16542,N_11741,N_12584);
nor U16543 (N_16543,N_13616,N_11843);
and U16544 (N_16544,N_12621,N_13682);
nand U16545 (N_16545,N_13103,N_13751);
and U16546 (N_16546,N_13791,N_14774);
nand U16547 (N_16547,N_11490,N_14568);
or U16548 (N_16548,N_12070,N_12724);
or U16549 (N_16549,N_10070,N_14846);
nor U16550 (N_16550,N_13894,N_13713);
or U16551 (N_16551,N_10811,N_13901);
or U16552 (N_16552,N_11256,N_11512);
or U16553 (N_16553,N_14553,N_13512);
and U16554 (N_16554,N_11100,N_10862);
nor U16555 (N_16555,N_12590,N_10273);
nor U16556 (N_16556,N_11373,N_11374);
xnor U16557 (N_16557,N_11558,N_12057);
nor U16558 (N_16558,N_12194,N_10979);
or U16559 (N_16559,N_12801,N_11494);
nand U16560 (N_16560,N_12091,N_12244);
nor U16561 (N_16561,N_11533,N_11056);
nand U16562 (N_16562,N_14498,N_11620);
or U16563 (N_16563,N_14051,N_12273);
nor U16564 (N_16564,N_11668,N_12505);
or U16565 (N_16565,N_12370,N_12465);
nor U16566 (N_16566,N_11754,N_12870);
xor U16567 (N_16567,N_13056,N_13077);
nor U16568 (N_16568,N_11984,N_10896);
nor U16569 (N_16569,N_13658,N_14684);
nor U16570 (N_16570,N_13113,N_12253);
nand U16571 (N_16571,N_10076,N_10507);
xor U16572 (N_16572,N_10068,N_11159);
and U16573 (N_16573,N_13935,N_14150);
xor U16574 (N_16574,N_14266,N_12545);
nor U16575 (N_16575,N_13989,N_12079);
or U16576 (N_16576,N_11716,N_11625);
and U16577 (N_16577,N_14834,N_10727);
and U16578 (N_16578,N_10150,N_13926);
or U16579 (N_16579,N_12808,N_11795);
nor U16580 (N_16580,N_13793,N_14357);
and U16581 (N_16581,N_13832,N_12577);
nor U16582 (N_16582,N_13431,N_10836);
nor U16583 (N_16583,N_13786,N_13719);
xnor U16584 (N_16584,N_13484,N_11827);
nor U16585 (N_16585,N_12139,N_12325);
nor U16586 (N_16586,N_11306,N_11557);
or U16587 (N_16587,N_11511,N_14174);
or U16588 (N_16588,N_10279,N_13813);
nand U16589 (N_16589,N_13740,N_12823);
or U16590 (N_16590,N_11421,N_12775);
nand U16591 (N_16591,N_12235,N_13620);
or U16592 (N_16592,N_11042,N_12630);
xor U16593 (N_16593,N_12817,N_14849);
nand U16594 (N_16594,N_13609,N_14463);
or U16595 (N_16595,N_13450,N_10135);
nor U16596 (N_16596,N_12893,N_10309);
xor U16597 (N_16597,N_12296,N_11824);
nor U16598 (N_16598,N_13543,N_13264);
nor U16599 (N_16599,N_11703,N_11121);
nand U16600 (N_16600,N_11443,N_14575);
nand U16601 (N_16601,N_12895,N_12125);
xnor U16602 (N_16602,N_11470,N_11195);
nand U16603 (N_16603,N_12910,N_14803);
or U16604 (N_16604,N_14278,N_12357);
and U16605 (N_16605,N_12636,N_12016);
nor U16606 (N_16606,N_10968,N_10377);
nor U16607 (N_16607,N_10229,N_12672);
and U16608 (N_16608,N_11362,N_10769);
and U16609 (N_16609,N_10800,N_14806);
or U16610 (N_16610,N_12407,N_12207);
xor U16611 (N_16611,N_13956,N_10102);
nand U16612 (N_16612,N_13082,N_11476);
nand U16613 (N_16613,N_10547,N_10414);
nor U16614 (N_16614,N_14888,N_12366);
or U16615 (N_16615,N_11046,N_13971);
nor U16616 (N_16616,N_11278,N_14077);
or U16617 (N_16617,N_10571,N_11653);
nand U16618 (N_16618,N_12727,N_13369);
and U16619 (N_16619,N_10187,N_13050);
or U16620 (N_16620,N_14737,N_10786);
nor U16621 (N_16621,N_13488,N_12574);
or U16622 (N_16622,N_12166,N_10736);
and U16623 (N_16623,N_12758,N_13929);
xnor U16624 (N_16624,N_14464,N_11304);
nand U16625 (N_16625,N_13884,N_11820);
nor U16626 (N_16626,N_12652,N_14004);
or U16627 (N_16627,N_10386,N_12409);
nor U16628 (N_16628,N_11107,N_10841);
nor U16629 (N_16629,N_10373,N_10172);
xnor U16630 (N_16630,N_12243,N_14393);
or U16631 (N_16631,N_10402,N_13281);
and U16632 (N_16632,N_12500,N_14391);
and U16633 (N_16633,N_14589,N_12416);
and U16634 (N_16634,N_11919,N_11285);
and U16635 (N_16635,N_11089,N_12744);
nand U16636 (N_16636,N_10430,N_14852);
nand U16637 (N_16637,N_13242,N_14306);
xnor U16638 (N_16638,N_11346,N_14203);
nor U16639 (N_16639,N_14510,N_10254);
nor U16640 (N_16640,N_11991,N_11615);
and U16641 (N_16641,N_14991,N_14354);
and U16642 (N_16642,N_13705,N_13202);
nor U16643 (N_16643,N_12795,N_10778);
nor U16644 (N_16644,N_11961,N_12198);
xnor U16645 (N_16645,N_14860,N_12261);
xor U16646 (N_16646,N_13748,N_10467);
xnor U16647 (N_16647,N_14484,N_11805);
nand U16648 (N_16648,N_10314,N_11252);
or U16649 (N_16649,N_11560,N_13160);
xor U16650 (N_16650,N_10180,N_12670);
nand U16651 (N_16651,N_10511,N_13710);
or U16652 (N_16652,N_12082,N_12952);
xor U16653 (N_16653,N_12439,N_10099);
nand U16654 (N_16654,N_10865,N_13963);
nor U16655 (N_16655,N_13344,N_13039);
and U16656 (N_16656,N_10240,N_14747);
nor U16657 (N_16657,N_12495,N_12497);
nor U16658 (N_16658,N_10393,N_10884);
xor U16659 (N_16659,N_12898,N_11139);
and U16660 (N_16660,N_13095,N_11091);
nand U16661 (N_16661,N_10268,N_13028);
nand U16662 (N_16662,N_10893,N_11610);
nor U16663 (N_16663,N_12140,N_11858);
nand U16664 (N_16664,N_14055,N_13670);
nand U16665 (N_16665,N_11760,N_14910);
or U16666 (N_16666,N_10772,N_13607);
and U16667 (N_16667,N_12988,N_10555);
and U16668 (N_16668,N_12412,N_13621);
nand U16669 (N_16669,N_10575,N_10456);
xor U16670 (N_16670,N_12718,N_12737);
and U16671 (N_16671,N_11172,N_13970);
and U16672 (N_16672,N_13086,N_14552);
or U16673 (N_16673,N_11253,N_13925);
xor U16674 (N_16674,N_14474,N_14798);
nand U16675 (N_16675,N_10870,N_14763);
nand U16676 (N_16676,N_10825,N_14929);
nand U16677 (N_16677,N_11200,N_11232);
or U16678 (N_16678,N_10955,N_12513);
nor U16679 (N_16679,N_14437,N_14744);
nand U16680 (N_16680,N_12920,N_14184);
and U16681 (N_16681,N_10785,N_11339);
nand U16682 (N_16682,N_12650,N_13232);
and U16683 (N_16683,N_11971,N_12866);
nor U16684 (N_16684,N_10178,N_10854);
or U16685 (N_16685,N_13907,N_10418);
and U16686 (N_16686,N_10856,N_13734);
or U16687 (N_16687,N_14268,N_10502);
xor U16688 (N_16688,N_14637,N_13982);
or U16689 (N_16689,N_13697,N_14383);
nor U16690 (N_16690,N_10034,N_11226);
or U16691 (N_16691,N_14408,N_11153);
xor U16692 (N_16692,N_12058,N_13747);
nor U16693 (N_16693,N_11877,N_10532);
nor U16694 (N_16694,N_12656,N_10667);
xor U16695 (N_16695,N_13587,N_11598);
nand U16696 (N_16696,N_10600,N_12309);
and U16697 (N_16697,N_10626,N_14663);
or U16698 (N_16698,N_13677,N_14076);
or U16699 (N_16699,N_10033,N_14609);
and U16700 (N_16700,N_12879,N_10122);
nand U16701 (N_16701,N_13526,N_14971);
and U16702 (N_16702,N_12812,N_14988);
nand U16703 (N_16703,N_11873,N_14216);
nand U16704 (N_16704,N_11497,N_12266);
and U16705 (N_16705,N_12794,N_11506);
or U16706 (N_16706,N_11720,N_14784);
nand U16707 (N_16707,N_13774,N_10989);
nand U16708 (N_16708,N_12402,N_13201);
nor U16709 (N_16709,N_12384,N_14427);
or U16710 (N_16710,N_12085,N_14491);
xnor U16711 (N_16711,N_11954,N_10408);
and U16712 (N_16712,N_11043,N_14169);
nor U16713 (N_16713,N_12464,N_11254);
and U16714 (N_16714,N_14326,N_14900);
nand U16715 (N_16715,N_14906,N_14446);
nor U16716 (N_16716,N_12230,N_12264);
xnor U16717 (N_16717,N_11429,N_11177);
xor U16718 (N_16718,N_12565,N_12302);
and U16719 (N_16719,N_11331,N_11323);
nor U16720 (N_16720,N_13052,N_13704);
or U16721 (N_16721,N_12169,N_10495);
nor U16722 (N_16722,N_10201,N_13329);
xnor U16723 (N_16723,N_14160,N_11266);
xnor U16724 (N_16724,N_10450,N_10144);
nor U16725 (N_16725,N_13349,N_11816);
nand U16726 (N_16726,N_11766,N_11349);
nor U16727 (N_16727,N_10438,N_13973);
nor U16728 (N_16728,N_12089,N_11580);
and U16729 (N_16729,N_10756,N_12728);
and U16730 (N_16730,N_13008,N_10924);
nor U16731 (N_16731,N_14225,N_14273);
and U16732 (N_16732,N_10509,N_14766);
xnor U16733 (N_16733,N_12829,N_12875);
nand U16734 (N_16734,N_11835,N_12417);
or U16735 (N_16735,N_11656,N_14454);
nor U16736 (N_16736,N_14343,N_14315);
xor U16737 (N_16737,N_13578,N_12514);
xor U16738 (N_16738,N_13708,N_14475);
nor U16739 (N_16739,N_10113,N_10169);
or U16740 (N_16740,N_12254,N_14080);
and U16741 (N_16741,N_12624,N_14082);
and U16742 (N_16742,N_13241,N_14042);
and U16743 (N_16743,N_12661,N_13990);
and U16744 (N_16744,N_10425,N_12248);
or U16745 (N_16745,N_11384,N_14136);
or U16746 (N_16746,N_13444,N_10556);
nand U16747 (N_16747,N_11745,N_14538);
xor U16748 (N_16748,N_11521,N_14083);
and U16749 (N_16749,N_12894,N_13163);
and U16750 (N_16750,N_13554,N_12689);
nor U16751 (N_16751,N_13513,N_11183);
xor U16752 (N_16752,N_11013,N_14883);
xor U16753 (N_16753,N_11478,N_14146);
or U16754 (N_16754,N_14899,N_11951);
and U16755 (N_16755,N_14565,N_14706);
nor U16756 (N_16756,N_10909,N_11302);
xor U16757 (N_16757,N_12019,N_13745);
or U16758 (N_16758,N_12740,N_10944);
xor U16759 (N_16759,N_14661,N_14556);
nand U16760 (N_16760,N_14624,N_12507);
nor U16761 (N_16761,N_10073,N_14523);
or U16762 (N_16762,N_14033,N_14753);
xor U16763 (N_16763,N_14395,N_11876);
or U16764 (N_16764,N_10010,N_12175);
and U16765 (N_16765,N_12962,N_11942);
or U16766 (N_16766,N_12288,N_11430);
nor U16767 (N_16767,N_11440,N_12081);
nor U16768 (N_16768,N_12665,N_13112);
nand U16769 (N_16769,N_12065,N_11791);
nand U16770 (N_16770,N_11999,N_10690);
nor U16771 (N_16771,N_11918,N_11380);
xnor U16772 (N_16772,N_14342,N_11659);
nor U16773 (N_16773,N_10728,N_14840);
and U16774 (N_16774,N_10845,N_11758);
or U16775 (N_16775,N_14610,N_12692);
and U16776 (N_16776,N_10226,N_10677);
nand U16777 (N_16777,N_11412,N_14105);
and U16778 (N_16778,N_14978,N_11111);
and U16779 (N_16779,N_12761,N_11734);
xnor U16780 (N_16780,N_13195,N_12072);
or U16781 (N_16781,N_11442,N_10434);
nor U16782 (N_16782,N_14708,N_11174);
or U16783 (N_16783,N_11465,N_14158);
or U16784 (N_16784,N_14365,N_14399);
xor U16785 (N_16785,N_12351,N_10685);
or U16786 (N_16786,N_13722,N_10485);
nand U16787 (N_16787,N_13692,N_11386);
and U16788 (N_16788,N_11513,N_12522);
nand U16789 (N_16789,N_12061,N_10161);
or U16790 (N_16790,N_10833,N_10682);
xor U16791 (N_16791,N_12274,N_13633);
or U16792 (N_16792,N_14178,N_14569);
and U16793 (N_16793,N_12813,N_14519);
xnor U16794 (N_16794,N_10803,N_10276);
nor U16795 (N_16795,N_10496,N_13206);
nor U16796 (N_16796,N_13029,N_12559);
or U16797 (N_16797,N_14466,N_14401);
and U16798 (N_16798,N_10829,N_12573);
and U16799 (N_16799,N_12452,N_11773);
or U16800 (N_16800,N_14345,N_12671);
xor U16801 (N_16801,N_10951,N_10295);
nor U16802 (N_16802,N_13154,N_11099);
and U16803 (N_16803,N_11934,N_14962);
xnor U16804 (N_16804,N_11160,N_13759);
xor U16805 (N_16805,N_11903,N_13150);
nor U16806 (N_16806,N_11041,N_11508);
or U16807 (N_16807,N_12594,N_12956);
nand U16808 (N_16808,N_12778,N_10987);
xnor U16809 (N_16809,N_12960,N_14420);
or U16810 (N_16810,N_11728,N_14768);
or U16811 (N_16811,N_12436,N_12924);
nand U16812 (N_16812,N_12554,N_10117);
nand U16813 (N_16813,N_10354,N_13549);
nor U16814 (N_16814,N_11249,N_11865);
or U16815 (N_16815,N_12582,N_11069);
nor U16816 (N_16816,N_13828,N_11829);
nand U16817 (N_16817,N_13560,N_13304);
nor U16818 (N_16818,N_13569,N_14028);
nand U16819 (N_16819,N_13134,N_12447);
nor U16820 (N_16820,N_13588,N_12308);
or U16821 (N_16821,N_11821,N_14309);
xnor U16822 (N_16822,N_14922,N_11675);
or U16823 (N_16823,N_13709,N_11673);
or U16824 (N_16824,N_13066,N_11730);
xor U16825 (N_16825,N_10554,N_13383);
xnor U16826 (N_16826,N_14557,N_12220);
nand U16827 (N_16827,N_14302,N_13437);
nor U16828 (N_16828,N_13556,N_13690);
or U16829 (N_16829,N_14110,N_14256);
nor U16830 (N_16830,N_10395,N_12964);
and U16831 (N_16831,N_12486,N_11150);
nor U16832 (N_16832,N_11808,N_10847);
xor U16833 (N_16833,N_10762,N_12741);
xor U16834 (N_16834,N_12153,N_10805);
and U16835 (N_16835,N_14855,N_11925);
nand U16836 (N_16836,N_14923,N_10400);
or U16837 (N_16837,N_13655,N_10256);
or U16838 (N_16838,N_11457,N_10114);
or U16839 (N_16839,N_14740,N_10181);
and U16840 (N_16840,N_13209,N_14366);
nor U16841 (N_16841,N_12944,N_14435);
nor U16842 (N_16842,N_13870,N_14656);
xor U16843 (N_16843,N_11997,N_13648);
xor U16844 (N_16844,N_14879,N_14752);
nor U16845 (N_16845,N_14037,N_14325);
nor U16846 (N_16846,N_11529,N_10695);
xor U16847 (N_16847,N_10704,N_14019);
nand U16848 (N_16848,N_13067,N_11718);
nand U16849 (N_16849,N_10782,N_14767);
and U16850 (N_16850,N_12782,N_11435);
nand U16851 (N_16851,N_11614,N_13773);
or U16852 (N_16852,N_13391,N_10044);
or U16853 (N_16853,N_12049,N_12660);
xor U16854 (N_16854,N_13733,N_11911);
nor U16855 (N_16855,N_11807,N_14555);
xnor U16856 (N_16856,N_12217,N_14936);
nor U16857 (N_16857,N_11233,N_13091);
nand U16858 (N_16858,N_10477,N_11176);
xnor U16859 (N_16859,N_12933,N_12874);
and U16860 (N_16860,N_10536,N_12673);
and U16861 (N_16861,N_13801,N_10897);
nand U16862 (N_16862,N_10791,N_14217);
or U16863 (N_16863,N_12662,N_12557);
nand U16864 (N_16864,N_10781,N_14157);
nand U16865 (N_16865,N_10293,N_13413);
nand U16866 (N_16866,N_14647,N_12942);
xor U16867 (N_16867,N_10097,N_12187);
nand U16868 (N_16868,N_14796,N_11333);
xor U16869 (N_16869,N_14099,N_13429);
nand U16870 (N_16870,N_14091,N_13481);
nor U16871 (N_16871,N_14215,N_11783);
and U16872 (N_16872,N_12704,N_12953);
or U16873 (N_16873,N_14780,N_11833);
xnor U16874 (N_16874,N_12578,N_11709);
xnor U16875 (N_16875,N_14307,N_10338);
or U16876 (N_16876,N_13375,N_13323);
and U16877 (N_16877,N_12896,N_12284);
and U16878 (N_16878,N_10465,N_11127);
nor U16879 (N_16879,N_13547,N_11572);
nor U16880 (N_16880,N_12892,N_12269);
nor U16881 (N_16881,N_10156,N_10476);
and U16882 (N_16882,N_14295,N_11992);
and U16883 (N_16883,N_12609,N_10984);
xor U16884 (N_16884,N_13378,N_11191);
or U16885 (N_16885,N_13874,N_13005);
xor U16886 (N_16886,N_12138,N_11914);
xnor U16887 (N_16887,N_10015,N_11848);
xnor U16888 (N_16888,N_10577,N_13908);
xnor U16889 (N_16889,N_12331,N_12669);
or U16890 (N_16890,N_12347,N_11680);
nor U16891 (N_16891,N_11725,N_10307);
and U16892 (N_16892,N_12310,N_10523);
or U16893 (N_16893,N_10120,N_13027);
or U16894 (N_16894,N_13634,N_14776);
or U16895 (N_16895,N_10490,N_14271);
xor U16896 (N_16896,N_12096,N_11602);
xnor U16897 (N_16897,N_11196,N_11265);
xor U16898 (N_16898,N_11275,N_10904);
nor U16899 (N_16899,N_13226,N_14791);
or U16900 (N_16900,N_12009,N_11804);
and U16901 (N_16901,N_13778,N_10245);
nand U16902 (N_16902,N_14782,N_10223);
xor U16903 (N_16903,N_14243,N_10975);
xnor U16904 (N_16904,N_13194,N_14172);
nand U16905 (N_16905,N_14863,N_12272);
nor U16906 (N_16906,N_12090,N_10328);
nand U16907 (N_16907,N_12404,N_10026);
and U16908 (N_16908,N_10222,N_13140);
or U16909 (N_16909,N_11531,N_11001);
and U16910 (N_16910,N_11792,N_10606);
and U16911 (N_16911,N_14138,N_10131);
xor U16912 (N_16912,N_13570,N_10479);
nand U16913 (N_16913,N_11173,N_14500);
nor U16914 (N_16914,N_10672,N_11229);
nor U16915 (N_16915,N_12493,N_14108);
nor U16916 (N_16916,N_11050,N_10432);
nor U16917 (N_16917,N_12484,N_13687);
nor U16918 (N_16918,N_11967,N_14059);
or U16919 (N_16919,N_10966,N_10765);
and U16920 (N_16920,N_10153,N_11815);
and U16921 (N_16921,N_14264,N_14696);
and U16922 (N_16922,N_14675,N_14069);
nand U16923 (N_16923,N_12936,N_10105);
nand U16924 (N_16924,N_12634,N_14604);
or U16925 (N_16925,N_10218,N_10041);
or U16926 (N_16926,N_12222,N_10446);
xnor U16927 (N_16927,N_14141,N_14621);
nand U16928 (N_16928,N_10922,N_11199);
or U16929 (N_16929,N_13203,N_14313);
or U16930 (N_16930,N_13490,N_10874);
xor U16931 (N_16931,N_10468,N_13171);
and U16932 (N_16932,N_11809,N_10466);
or U16933 (N_16933,N_13033,N_14642);
xnor U16934 (N_16934,N_11313,N_11054);
nand U16935 (N_16935,N_12721,N_12534);
xor U16936 (N_16936,N_10826,N_13954);
nand U16937 (N_16937,N_14045,N_14471);
nand U16938 (N_16938,N_13999,N_12324);
nand U16939 (N_16939,N_12463,N_13355);
nand U16940 (N_16940,N_10585,N_14025);
nand U16941 (N_16941,N_11559,N_14116);
xor U16942 (N_16942,N_13688,N_12294);
and U16943 (N_16943,N_13819,N_14341);
and U16944 (N_16944,N_10457,N_10588);
and U16945 (N_16945,N_13841,N_12011);
nand U16946 (N_16946,N_11577,N_10888);
and U16947 (N_16947,N_14578,N_11931);
nor U16948 (N_16948,N_11587,N_14322);
or U16949 (N_16949,N_12982,N_11502);
nand U16950 (N_16950,N_10175,N_11875);
and U16951 (N_16951,N_13644,N_11070);
nor U16952 (N_16952,N_11586,N_13510);
nor U16953 (N_16953,N_11714,N_11312);
xnor U16954 (N_16954,N_10774,N_14164);
or U16955 (N_16955,N_12450,N_12774);
xor U16956 (N_16956,N_12620,N_13776);
nand U16957 (N_16957,N_12496,N_11856);
and U16958 (N_16958,N_13950,N_10217);
and U16959 (N_16959,N_14536,N_13204);
xnor U16960 (N_16960,N_12300,N_13936);
xor U16961 (N_16961,N_10572,N_10654);
nand U16962 (N_16962,N_13162,N_10790);
and U16963 (N_16963,N_11137,N_12990);
and U16964 (N_16964,N_11547,N_10248);
nand U16965 (N_16965,N_13295,N_14522);
nand U16966 (N_16966,N_10143,N_13561);
and U16967 (N_16967,N_13896,N_13158);
nand U16968 (N_16968,N_10883,N_14516);
nand U16969 (N_16969,N_12030,N_11381);
nor U16970 (N_16970,N_13641,N_10177);
and U16971 (N_16971,N_13530,N_10530);
nand U16972 (N_16972,N_12481,N_14290);
and U16973 (N_16973,N_14281,N_14743);
nand U16974 (N_16974,N_11484,N_13913);
or U16975 (N_16975,N_14667,N_12598);
or U16976 (N_16976,N_13496,N_11129);
xor U16977 (N_16977,N_10230,N_13009);
xnor U16978 (N_16978,N_10664,N_14711);
and U16979 (N_16979,N_11496,N_10855);
nor U16980 (N_16980,N_11831,N_11943);
and U16981 (N_16981,N_14479,N_11216);
xnor U16982 (N_16982,N_10519,N_14071);
xor U16983 (N_16983,N_14577,N_14040);
nand U16984 (N_16984,N_13718,N_14156);
xor U16985 (N_16985,N_11989,N_11449);
and U16986 (N_16986,N_11552,N_11020);
and U16987 (N_16987,N_14003,N_11759);
or U16988 (N_16988,N_14142,N_14832);
nor U16989 (N_16989,N_10551,N_10459);
or U16990 (N_16990,N_11926,N_14941);
nand U16991 (N_16991,N_14646,N_13280);
xnor U16992 (N_16992,N_12460,N_13888);
nand U16993 (N_16993,N_13260,N_12446);
nor U16994 (N_16994,N_11944,N_14525);
or U16995 (N_16995,N_13805,N_14411);
or U16996 (N_16996,N_13370,N_11867);
nand U16997 (N_16997,N_12976,N_13955);
or U16998 (N_16998,N_12340,N_10779);
nor U16999 (N_16999,N_12312,N_11397);
xnor U17000 (N_17000,N_12568,N_14185);
xor U17001 (N_17001,N_13666,N_10193);
and U17002 (N_17002,N_13139,N_11976);
nor U17003 (N_17003,N_10287,N_10902);
xor U17004 (N_17004,N_10686,N_12482);
or U17005 (N_17005,N_13217,N_11998);
nor U17006 (N_17006,N_12040,N_10299);
or U17007 (N_17007,N_14455,N_10684);
or U17008 (N_17008,N_13300,N_10292);
nand U17009 (N_17009,N_12931,N_10064);
nand U17010 (N_17010,N_11515,N_14047);
and U17011 (N_17011,N_12165,N_14062);
nor U17012 (N_17012,N_13211,N_11340);
or U17013 (N_17013,N_14209,N_12381);
or U17014 (N_17014,N_12714,N_11461);
nor U17015 (N_17015,N_11870,N_10288);
nor U17016 (N_17016,N_12241,N_11231);
nand U17017 (N_17017,N_14124,N_14023);
xor U17018 (N_17018,N_11880,N_11332);
nor U17019 (N_17019,N_12681,N_12489);
and U17020 (N_17020,N_12050,N_14792);
or U17021 (N_17021,N_11881,N_14921);
nor U17022 (N_17022,N_12499,N_11206);
or U17023 (N_17023,N_11097,N_10200);
and U17024 (N_17024,N_13721,N_14616);
or U17025 (N_17025,N_10285,N_14229);
nor U17026 (N_17026,N_12989,N_14958);
nand U17027 (N_17027,N_11405,N_11336);
nand U17028 (N_17028,N_13458,N_11762);
nand U17029 (N_17029,N_11702,N_13998);
xnor U17030 (N_17030,N_12979,N_10722);
xnor U17031 (N_17031,N_14716,N_13197);
or U17032 (N_17032,N_10597,N_12183);
or U17033 (N_17033,N_11955,N_10359);
and U17034 (N_17034,N_12551,N_10570);
and U17035 (N_17035,N_13723,N_14212);
or U17036 (N_17036,N_11932,N_10978);
xor U17037 (N_17037,N_13156,N_12442);
nor U17038 (N_17038,N_11272,N_13542);
nor U17039 (N_17039,N_12440,N_11108);
and U17040 (N_17040,N_10419,N_12474);
nor U17041 (N_17041,N_13905,N_11436);
xor U17042 (N_17042,N_14773,N_10563);
or U17043 (N_17043,N_12007,N_13368);
nand U17044 (N_17044,N_12354,N_13699);
nor U17045 (N_17045,N_10413,N_12042);
nand U17046 (N_17046,N_10160,N_10007);
or U17047 (N_17047,N_14316,N_14039);
xor U17048 (N_17048,N_10035,N_12297);
or U17049 (N_17049,N_11920,N_11370);
and U17050 (N_17050,N_10372,N_12397);
nor U17051 (N_17051,N_10157,N_14207);
nor U17052 (N_17052,N_11952,N_11549);
nand U17053 (N_17053,N_12717,N_13298);
and U17054 (N_17054,N_14564,N_14558);
nor U17055 (N_17055,N_11950,N_11427);
or U17056 (N_17056,N_13184,N_11900);
or U17057 (N_17057,N_12353,N_11902);
and U17058 (N_17058,N_11102,N_12268);
and U17059 (N_17059,N_13149,N_10277);
or U17060 (N_17060,N_12216,N_10118);
and U17061 (N_17061,N_13761,N_13120);
xnor U17062 (N_17062,N_11310,N_13051);
nand U17063 (N_17063,N_11811,N_13826);
nor U17064 (N_17064,N_14257,N_11467);
and U17065 (N_17065,N_11289,N_12959);
nor U17066 (N_17066,N_13595,N_14102);
xnor U17067 (N_17067,N_13550,N_10531);
or U17068 (N_17068,N_14097,N_11579);
nor U17069 (N_17069,N_10573,N_14520);
or U17070 (N_17070,N_13984,N_12518);
or U17071 (N_17071,N_11103,N_10901);
xnor U17072 (N_17072,N_12985,N_14504);
nand U17073 (N_17073,N_11736,N_14673);
nand U17074 (N_17074,N_13546,N_10520);
xnor U17075 (N_17075,N_14125,N_13902);
or U17076 (N_17076,N_12472,N_14907);
or U17077 (N_17077,N_14546,N_11688);
nand U17078 (N_17078,N_13504,N_13771);
nand U17079 (N_17079,N_10719,N_11328);
nand U17080 (N_17080,N_11341,N_13811);
or U17081 (N_17081,N_10267,N_10518);
nor U17082 (N_17082,N_10876,N_10804);
or U17083 (N_17083,N_14460,N_11978);
or U17084 (N_17084,N_11062,N_11118);
nor U17085 (N_17085,N_11699,N_10923);
xnor U17086 (N_17086,N_10881,N_14654);
nor U17087 (N_17087,N_12227,N_11882);
nor U17088 (N_17088,N_12571,N_10182);
xnor U17089 (N_17089,N_11238,N_14623);
and U17090 (N_17090,N_13316,N_12023);
and U17091 (N_17091,N_11608,N_14104);
nand U17092 (N_17092,N_14030,N_12877);
and U17093 (N_17093,N_13885,N_13128);
nand U17094 (N_17094,N_14512,N_12980);
nor U17095 (N_17095,N_13724,N_10521);
and U17096 (N_17096,N_11296,N_14432);
xnor U17097 (N_17097,N_11938,N_14613);
xnor U17098 (N_17098,N_12024,N_14349);
or U17099 (N_17099,N_11523,N_12435);
nor U17100 (N_17100,N_14912,N_10152);
nand U17101 (N_17101,N_13395,N_10698);
xor U17102 (N_17102,N_10652,N_12321);
nand U17103 (N_17103,N_13976,N_12041);
xnor U17104 (N_17104,N_10311,N_11860);
nand U17105 (N_17105,N_12477,N_14639);
nand U17106 (N_17106,N_14131,N_12270);
or U17107 (N_17107,N_12363,N_13915);
or U17108 (N_17108,N_10887,N_14818);
xor U17109 (N_17109,N_11517,N_14775);
nand U17110 (N_17110,N_11363,N_13528);
nor U17111 (N_17111,N_12144,N_13035);
nand U17112 (N_17112,N_11726,N_11636);
nand U17113 (N_17113,N_13880,N_10734);
or U17114 (N_17114,N_13393,N_11404);
xnor U17115 (N_17115,N_12062,N_10755);
nor U17116 (N_17116,N_12066,N_14598);
nand U17117 (N_17117,N_12229,N_11657);
and U17118 (N_17118,N_12531,N_12039);
or U17119 (N_17119,N_10335,N_12257);
nand U17120 (N_17120,N_12113,N_14892);
xnor U17121 (N_17121,N_10333,N_12793);
and U17122 (N_17122,N_11040,N_12515);
nand U17123 (N_17123,N_12263,N_10014);
xnor U17124 (N_17124,N_14384,N_10392);
nand U17125 (N_17125,N_14754,N_13409);
or U17126 (N_17126,N_12180,N_13076);
nand U17127 (N_17127,N_11717,N_12280);
nand U17128 (N_17128,N_12170,N_14995);
or U17129 (N_17129,N_13922,N_11175);
or U17130 (N_17130,N_14014,N_14378);
or U17131 (N_17131,N_13054,N_14977);
nor U17132 (N_17132,N_11075,N_12350);
and U17133 (N_17133,N_12658,N_11204);
nand U17134 (N_17134,N_14487,N_12691);
nor U17135 (N_17135,N_13638,N_11715);
or U17136 (N_17136,N_14573,N_11395);
or U17137 (N_17137,N_12242,N_11729);
nor U17138 (N_17138,N_11084,N_14114);
nor U17139 (N_17139,N_11825,N_12178);
and U17140 (N_17140,N_11845,N_10838);
nand U17141 (N_17141,N_10535,N_14126);
nor U17142 (N_17142,N_13462,N_12520);
or U17143 (N_17143,N_13361,N_14762);
xnor U17144 (N_17144,N_11631,N_12916);
and U17145 (N_17145,N_10198,N_12256);
nand U17146 (N_17146,N_14154,N_12593);
or U17147 (N_17147,N_11325,N_12306);
and U17148 (N_17148,N_11125,N_13667);
nand U17149 (N_17149,N_12002,N_12255);
and U17150 (N_17150,N_14472,N_13788);
xnor U17151 (N_17151,N_10164,N_14959);
and U17152 (N_17152,N_10030,N_12469);
or U17153 (N_17153,N_13840,N_11378);
or U17154 (N_17154,N_14721,N_13071);
or U17155 (N_17155,N_10019,N_13881);
or U17156 (N_17156,N_13399,N_10381);
and U17157 (N_17157,N_14660,N_12957);
nand U17158 (N_17158,N_13594,N_10994);
xor U17159 (N_17159,N_13775,N_13650);
nand U17160 (N_17160,N_10199,N_14882);
xor U17161 (N_17161,N_11236,N_10096);
nand U17162 (N_17162,N_12063,N_10943);
xnor U17163 (N_17163,N_10964,N_12519);
nor U17164 (N_17164,N_14123,N_14845);
xor U17165 (N_17165,N_10366,N_12999);
nor U17166 (N_17166,N_12005,N_10316);
nor U17167 (N_17167,N_10216,N_10274);
xor U17168 (N_17168,N_11481,N_12164);
nand U17169 (N_17169,N_11093,N_10583);
nor U17170 (N_17170,N_11456,N_11871);
nand U17171 (N_17171,N_14397,N_13796);
or U17172 (N_17172,N_11933,N_14690);
or U17173 (N_17173,N_14857,N_12233);
nor U17174 (N_17174,N_14652,N_14544);
nand U17175 (N_17175,N_12863,N_13216);
or U17176 (N_17176,N_13838,N_11768);
nand U17177 (N_17177,N_14973,N_10500);
nor U17178 (N_17178,N_14337,N_12523);
or U17179 (N_17179,N_14234,N_14283);
and U17180 (N_17180,N_12803,N_10363);
and U17181 (N_17181,N_12806,N_14269);
nand U17182 (N_17182,N_14574,N_12943);
nor U17183 (N_17183,N_14486,N_10183);
xor U17184 (N_17184,N_10993,N_13155);
nand U17185 (N_17185,N_12792,N_11701);
and U17186 (N_17186,N_10528,N_12770);
nand U17187 (N_17187,N_12342,N_14359);
and U17188 (N_17188,N_12114,N_13598);
or U17189 (N_17189,N_14627,N_12037);
and U17190 (N_17190,N_14170,N_10481);
nand U17191 (N_17191,N_10882,N_12345);
and U17192 (N_17192,N_10817,N_13310);
or U17193 (N_17193,N_13421,N_14904);
or U17194 (N_17194,N_12646,N_10458);
or U17195 (N_17195,N_10549,N_11315);
xnor U17196 (N_17196,N_14506,N_13236);
and U17197 (N_17197,N_12749,N_14951);
xor U17198 (N_17198,N_12080,N_12320);
nor U17199 (N_17199,N_12641,N_10179);
xnor U17200 (N_17200,N_10659,N_14963);
nor U17201 (N_17201,N_14505,N_10550);
nor U17202 (N_17202,N_14477,N_10593);
xnor U17203 (N_17203,N_11198,N_11916);
or U17204 (N_17204,N_12034,N_11866);
nand U17205 (N_17205,N_14540,N_14723);
nor U17206 (N_17206,N_13354,N_12118);
nand U17207 (N_17207,N_10513,N_14967);
or U17208 (N_17208,N_13318,N_10215);
and U17209 (N_17209,N_14255,N_12184);
nor U17210 (N_17210,N_11471,N_11372);
nand U17211 (N_17211,N_11027,N_13252);
nor U17212 (N_17212,N_11834,N_10891);
nor U17213 (N_17213,N_12099,N_10324);
and U17214 (N_17214,N_11109,N_12123);
xor U17215 (N_17215,N_12206,N_12511);
or U17216 (N_17216,N_10326,N_14709);
or U17217 (N_17217,N_11480,N_10250);
and U17218 (N_17218,N_13124,N_12623);
and U17219 (N_17219,N_14703,N_12753);
nor U17220 (N_17220,N_12688,N_12401);
and U17221 (N_17221,N_12185,N_10713);
and U17222 (N_17222,N_10839,N_13407);
nor U17223 (N_17223,N_13789,N_10145);
nor U17224 (N_17224,N_10818,N_13358);
xor U17225 (N_17225,N_10206,N_13455);
xnor U17226 (N_17226,N_14119,N_11819);
or U17227 (N_17227,N_13041,N_14008);
xnor U17228 (N_17228,N_14381,N_13336);
and U17229 (N_17229,N_10282,N_11447);
and U17230 (N_17230,N_13584,N_13294);
and U17231 (N_17231,N_11314,N_11526);
and U17232 (N_17232,N_11068,N_10960);
and U17233 (N_17233,N_13853,N_10602);
or U17234 (N_17234,N_10831,N_11694);
nor U17235 (N_17235,N_10973,N_11420);
nor U17236 (N_17236,N_10235,N_10974);
nand U17237 (N_17237,N_14679,N_10956);
xnor U17238 (N_17238,N_11224,N_14351);
nor U17239 (N_17239,N_12459,N_14113);
xor U17240 (N_17240,N_11066,N_10391);
nor U17241 (N_17241,N_14440,N_10795);
nor U17242 (N_17242,N_12095,N_10410);
nor U17243 (N_17243,N_10615,N_12221);
nor U17244 (N_17244,N_11663,N_10566);
xnor U17245 (N_17245,N_14441,N_13321);
and U17246 (N_17246,N_13180,N_14651);
nand U17247 (N_17247,N_11207,N_12329);
nand U17248 (N_17248,N_14779,N_13684);
or U17249 (N_17249,N_12967,N_13330);
or U17250 (N_17250,N_10735,N_14648);
nand U17251 (N_17251,N_14287,N_12260);
nor U17252 (N_17252,N_10009,N_11930);
or U17253 (N_17253,N_13851,N_10653);
nor U17254 (N_17254,N_11303,N_10977);
or U17255 (N_17255,N_10506,N_14167);
or U17256 (N_17256,N_12595,N_10534);
or U17257 (N_17257,N_12116,N_11450);
and U17258 (N_17258,N_11290,N_11692);
nor U17259 (N_17259,N_11828,N_11451);
and U17260 (N_17260,N_12785,N_13348);
nand U17261 (N_17261,N_13538,N_10461);
nand U17262 (N_17262,N_10066,N_14151);
or U17263 (N_17263,N_12791,N_12047);
and U17264 (N_17264,N_14841,N_14851);
nand U17265 (N_17265,N_12371,N_13939);
xnor U17266 (N_17266,N_10879,N_13959);
or U17267 (N_17267,N_10054,N_14814);
nor U17268 (N_17268,N_14815,N_14473);
nor U17269 (N_17269,N_10976,N_11564);
xor U17270 (N_17270,N_13166,N_13969);
nor U17271 (N_17271,N_14902,N_14626);
or U17272 (N_17272,N_10421,N_10154);
nand U17273 (N_17273,N_12816,N_12104);
and U17274 (N_17274,N_14653,N_13200);
and U17275 (N_17275,N_13603,N_13445);
or U17276 (N_17276,N_13979,N_10623);
and U17277 (N_17277,N_11915,N_13482);
or U17278 (N_17278,N_11770,N_13966);
nand U17279 (N_17279,N_14903,N_10959);
nor U17280 (N_17280,N_10020,N_11789);
or U17281 (N_17281,N_14368,N_12501);
nand U17282 (N_17282,N_14937,N_11446);
and U17283 (N_17283,N_12747,N_11690);
nor U17284 (N_17284,N_12337,N_12977);
and U17285 (N_17285,N_13574,N_14842);
nand U17286 (N_17286,N_10750,N_10658);
and U17287 (N_17287,N_10094,N_13495);
or U17288 (N_17288,N_11681,N_10284);
nor U17289 (N_17289,N_14717,N_10208);
or U17290 (N_17290,N_10090,N_12192);
or U17291 (N_17291,N_13261,N_11669);
or U17292 (N_17292,N_14461,N_11575);
xor U17293 (N_17293,N_11168,N_10228);
nand U17294 (N_17294,N_14090,N_10937);
and U17295 (N_17295,N_14389,N_10219);
or U17296 (N_17296,N_12535,N_11151);
or U17297 (N_17297,N_10167,N_10663);
nand U17298 (N_17298,N_11901,N_10898);
and U17299 (N_17299,N_12891,N_11003);
xor U17300 (N_17300,N_14914,N_10648);
nor U17301 (N_17301,N_12538,N_10484);
nor U17302 (N_17302,N_10209,N_12619);
or U17303 (N_17303,N_11553,N_14641);
nand U17304 (N_17304,N_10067,N_10868);
nand U17305 (N_17305,N_10828,N_13781);
xor U17306 (N_17306,N_14001,N_10115);
and U17307 (N_17307,N_14645,N_10643);
or U17308 (N_17308,N_14450,N_10849);
and U17309 (N_17309,N_14068,N_10089);
nor U17310 (N_17310,N_10806,N_10892);
nand U17311 (N_17311,N_11664,N_10092);
xnor U17312 (N_17312,N_12763,N_14585);
or U17313 (N_17313,N_13795,N_13892);
xor U17314 (N_17314,N_13332,N_14649);
or U17315 (N_17315,N_10546,N_13115);
and U17316 (N_17316,N_12830,N_13464);
nor U17317 (N_17317,N_14180,N_11899);
and U17318 (N_17318,N_12424,N_11607);
xnor U17319 (N_17319,N_11141,N_13167);
nand U17320 (N_17320,N_14371,N_13403);
nand U17321 (N_17321,N_14576,N_13085);
or U17322 (N_17322,N_14893,N_13317);
xor U17323 (N_17323,N_13665,N_10717);
nand U17324 (N_17324,N_13309,N_13614);
nor U17325 (N_17325,N_14788,N_14918);
xor U17326 (N_17326,N_10676,N_13878);
xnor U17327 (N_17327,N_13296,N_14065);
nor U17328 (N_17328,N_11023,N_12398);
nand U17329 (N_17329,N_11850,N_10133);
nand U17330 (N_17330,N_14191,N_13768);
nand U17331 (N_17331,N_11459,N_14193);
or U17332 (N_17332,N_14533,N_12855);
nor U17333 (N_17333,N_10110,N_10629);
and U17334 (N_17334,N_13243,N_10121);
nand U17335 (N_17335,N_12189,N_10742);
nand U17336 (N_17336,N_13188,N_14324);
or U17337 (N_17337,N_12045,N_12729);
or U17338 (N_17338,N_12405,N_14662);
and U17339 (N_17339,N_12163,N_14020);
nand U17340 (N_17340,N_14489,N_13335);
nor U17341 (N_17341,N_13914,N_14109);
nor U17342 (N_17342,N_12372,N_10624);
nand U17343 (N_17343,N_11970,N_10051);
nand U17344 (N_17344,N_14492,N_10730);
and U17345 (N_17345,N_13412,N_13852);
nor U17346 (N_17346,N_13229,N_12702);
and U17347 (N_17347,N_13427,N_14582);
and U17348 (N_17348,N_11784,N_14183);
xor U17349 (N_17349,N_14006,N_14927);
xor U17350 (N_17350,N_12451,N_14692);
nor U17351 (N_17351,N_13792,N_10802);
or U17352 (N_17352,N_11565,N_12053);
or U17353 (N_17353,N_10903,N_12316);
nor U17354 (N_17354,N_11894,N_10586);
xnor U17355 (N_17355,N_10360,N_10057);
xor U17356 (N_17356,N_11294,N_13334);
xnor U17357 (N_17357,N_11618,N_11123);
or U17358 (N_17358,N_12106,N_13013);
nor U17359 (N_17359,N_14594,N_14139);
or U17360 (N_17360,N_14038,N_14866);
or U17361 (N_17361,N_14835,N_10706);
xnor U17362 (N_17362,N_14095,N_11887);
nand U17363 (N_17363,N_13305,N_12607);
and U17364 (N_17364,N_10580,N_11813);
and U17365 (N_17365,N_10703,N_13447);
and U17366 (N_17366,N_14195,N_10599);
nor U17367 (N_17367,N_12616,N_12693);
and U17368 (N_17368,N_10491,N_10371);
xor U17369 (N_17369,N_12983,N_13417);
nor U17370 (N_17370,N_12092,N_13871);
and U17371 (N_17371,N_10085,N_13228);
or U17372 (N_17372,N_12210,N_10271);
or U17373 (N_17373,N_10548,N_13145);
and U17374 (N_17374,N_13520,N_11555);
and U17375 (N_17375,N_12422,N_10246);
or U17376 (N_17376,N_13890,N_14994);
nand U17377 (N_17377,N_13988,N_12975);
nor U17378 (N_17378,N_13401,N_13635);
nand U17379 (N_17379,N_11986,N_11650);
xor U17380 (N_17380,N_10801,N_14379);
nor U17381 (N_17381,N_13800,N_14219);
nor U17382 (N_17382,N_12835,N_11855);
or U17383 (N_17383,N_10203,N_12655);
nand U17384 (N_17384,N_11220,N_13879);
and U17385 (N_17385,N_11857,N_13098);
xnor U17386 (N_17386,N_12133,N_14704);
or U17387 (N_17387,N_12921,N_13572);
or U17388 (N_17388,N_13192,N_13529);
nand U17389 (N_17389,N_13940,N_14103);
xor U17390 (N_17390,N_12374,N_12410);
or U17391 (N_17391,N_11852,N_14057);
nor U17392 (N_17392,N_14304,N_11985);
nand U17393 (N_17393,N_13680,N_14843);
nor U17394 (N_17394,N_12132,N_13116);
and U17395 (N_17395,N_14133,N_14155);
nand U17396 (N_17396,N_14676,N_11812);
xor U17397 (N_17397,N_12996,N_13992);
nor U17398 (N_17398,N_11017,N_13235);
or U17399 (N_17399,N_11719,N_14996);
or U17400 (N_17400,N_11163,N_10981);
or U17401 (N_17401,N_10560,N_10912);
xor U17402 (N_17402,N_14694,N_13207);
and U17403 (N_17403,N_14748,N_11048);
or U17404 (N_17404,N_10958,N_13559);
or U17405 (N_17405,N_14044,N_13953);
nor U17406 (N_17406,N_10464,N_13142);
and U17407 (N_17407,N_14421,N_14107);
or U17408 (N_17408,N_10645,N_14416);
and U17409 (N_17409,N_10186,N_13693);
and U17410 (N_17410,N_10192,N_12772);
nand U17411 (N_17411,N_11203,N_10047);
nor U17412 (N_17412,N_13818,N_14789);
nor U17413 (N_17413,N_14376,N_12490);
nand U17414 (N_17414,N_14804,N_12935);
or U17415 (N_17415,N_10949,N_11403);
nor U17416 (N_17416,N_13231,N_11872);
xor U17417 (N_17417,N_13882,N_13514);
nand U17418 (N_17418,N_10687,N_13919);
nand U17419 (N_17419,N_11122,N_10568);
nand U17420 (N_17420,N_13034,N_14828);
nand U17421 (N_17421,N_11158,N_13057);
or U17422 (N_17422,N_12203,N_11583);
nand U17423 (N_17423,N_14483,N_12919);
nand U17424 (N_17424,N_14790,N_10353);
nand U17425 (N_17425,N_13459,N_10081);
xor U17426 (N_17426,N_10024,N_14758);
nand U17427 (N_17427,N_11814,N_13639);
and U17428 (N_17428,N_11695,N_11214);
xnor U17429 (N_17429,N_14192,N_13499);
and U17430 (N_17430,N_10584,N_13799);
or U17431 (N_17431,N_11117,N_12488);
nand U17432 (N_17432,N_11704,N_12172);
xnor U17433 (N_17433,N_11140,N_10297);
xnor U17434 (N_17434,N_14392,N_10000);
xnor U17435 (N_17435,N_11187,N_13161);
nor U17436 (N_17436,N_12202,N_12084);
nand U17437 (N_17437,N_13314,N_11710);
or U17438 (N_17438,N_14433,N_10079);
xor U17439 (N_17439,N_12810,N_10397);
xnor U17440 (N_17440,N_12904,N_12972);
or U17441 (N_17441,N_11847,N_12406);
or U17442 (N_17442,N_12015,N_10165);
nor U17443 (N_17443,N_13987,N_11184);
xnor U17444 (N_17444,N_13815,N_11921);
xor U17445 (N_17445,N_13610,N_14603);
or U17446 (N_17446,N_14202,N_10783);
nor U17447 (N_17447,N_10705,N_14242);
or U17448 (N_17448,N_11005,N_10345);
nor U17449 (N_17449,N_12067,N_14318);
nor U17450 (N_17450,N_11501,N_12564);
nor U17451 (N_17451,N_11053,N_14591);
or U17452 (N_17452,N_11283,N_10197);
or U17453 (N_17453,N_14050,N_13426);
nor U17454 (N_17454,N_14529,N_14974);
nand U17455 (N_17455,N_10557,N_12884);
or U17456 (N_17456,N_14462,N_11796);
nand U17457 (N_17457,N_14695,N_11101);
xor U17458 (N_17458,N_13465,N_11965);
or U17459 (N_17459,N_11995,N_10361);
nand U17460 (N_17460,N_13943,N_13475);
nor U17461 (N_17461,N_14222,N_12504);
nor U17462 (N_17462,N_10462,N_13031);
or U17463 (N_17463,N_11057,N_12218);
nor U17464 (N_17464,N_11133,N_11686);
or U17465 (N_17465,N_14854,N_14347);
xor U17466 (N_17466,N_12606,N_14701);
or U17467 (N_17467,N_14548,N_13205);
and U17468 (N_17468,N_12213,N_10136);
or U17469 (N_17469,N_12361,N_11051);
or U17470 (N_17470,N_11110,N_10394);
nor U17471 (N_17471,N_14541,N_12570);
and U17472 (N_17472,N_13942,N_14111);
or U17473 (N_17473,N_14292,N_10422);
nor U17474 (N_17474,N_14148,N_13707);
xnor U17475 (N_17475,N_12862,N_10644);
or U17476 (N_17476,N_12247,N_13516);
or U17477 (N_17477,N_12678,N_10745);
xnor U17478 (N_17478,N_10494,N_10709);
nor U17479 (N_17479,N_13934,N_10368);
and U17480 (N_17480,N_14881,N_10084);
nor U17481 (N_17481,N_12645,N_11797);
and U17482 (N_17482,N_11194,N_11689);
xor U17483 (N_17483,N_13715,N_13208);
nor U17484 (N_17484,N_10213,N_10074);
xor U17485 (N_17485,N_10559,N_11844);
or U17486 (N_17486,N_13262,N_12552);
and U17487 (N_17487,N_13743,N_13193);
xnor U17488 (N_17488,N_10991,N_10631);
or U17489 (N_17489,N_10489,N_12237);
and U17490 (N_17490,N_10257,N_11525);
or U17491 (N_17491,N_14132,N_10343);
and U17492 (N_17492,N_10050,N_13803);
nand U17493 (N_17493,N_11082,N_10680);
nand U17494 (N_17494,N_14947,N_10918);
nand U17495 (N_17495,N_13501,N_11969);
nor U17496 (N_17496,N_13810,N_14956);
and U17497 (N_17497,N_11258,N_13129);
or U17498 (N_17498,N_12909,N_10873);
nor U17499 (N_17499,N_12295,N_13102);
and U17500 (N_17500,N_12797,N_11862);
or U17501 (N_17501,N_11478,N_12819);
nor U17502 (N_17502,N_10147,N_12220);
or U17503 (N_17503,N_14022,N_14817);
nor U17504 (N_17504,N_11690,N_11909);
nor U17505 (N_17505,N_14717,N_11561);
and U17506 (N_17506,N_10918,N_10949);
nand U17507 (N_17507,N_10737,N_11903);
nor U17508 (N_17508,N_11482,N_14411);
xnor U17509 (N_17509,N_13141,N_10495);
nor U17510 (N_17510,N_13222,N_12165);
xor U17511 (N_17511,N_11929,N_14373);
xor U17512 (N_17512,N_14703,N_13661);
nor U17513 (N_17513,N_14558,N_12740);
xor U17514 (N_17514,N_10367,N_12795);
nor U17515 (N_17515,N_12454,N_13859);
xor U17516 (N_17516,N_13127,N_10713);
nand U17517 (N_17517,N_10531,N_14055);
nor U17518 (N_17518,N_10491,N_12301);
nor U17519 (N_17519,N_10005,N_10647);
nor U17520 (N_17520,N_11291,N_10144);
or U17521 (N_17521,N_13168,N_11395);
xnor U17522 (N_17522,N_11735,N_13815);
nor U17523 (N_17523,N_12839,N_13316);
xor U17524 (N_17524,N_10207,N_11804);
or U17525 (N_17525,N_10863,N_12406);
nor U17526 (N_17526,N_12438,N_14313);
and U17527 (N_17527,N_10979,N_14403);
and U17528 (N_17528,N_13059,N_10379);
and U17529 (N_17529,N_14946,N_13706);
nand U17530 (N_17530,N_12224,N_10028);
or U17531 (N_17531,N_14464,N_11124);
and U17532 (N_17532,N_11554,N_14438);
and U17533 (N_17533,N_11355,N_11341);
or U17534 (N_17534,N_11697,N_13803);
nand U17535 (N_17535,N_10693,N_10639);
and U17536 (N_17536,N_14400,N_14066);
or U17537 (N_17537,N_10217,N_14288);
nand U17538 (N_17538,N_13030,N_14657);
nor U17539 (N_17539,N_14035,N_14130);
xor U17540 (N_17540,N_11740,N_12344);
and U17541 (N_17541,N_10373,N_11198);
nand U17542 (N_17542,N_11209,N_10966);
nand U17543 (N_17543,N_11666,N_14364);
nor U17544 (N_17544,N_14396,N_11012);
xor U17545 (N_17545,N_12843,N_14073);
nand U17546 (N_17546,N_13482,N_13296);
nor U17547 (N_17547,N_13654,N_13204);
xor U17548 (N_17548,N_12584,N_14746);
nand U17549 (N_17549,N_14875,N_11324);
xor U17550 (N_17550,N_13598,N_10722);
nand U17551 (N_17551,N_12864,N_12499);
xnor U17552 (N_17552,N_14791,N_10497);
nor U17553 (N_17553,N_10773,N_14986);
or U17554 (N_17554,N_14029,N_14631);
nor U17555 (N_17555,N_13398,N_13198);
nor U17556 (N_17556,N_13330,N_13569);
and U17557 (N_17557,N_10337,N_12232);
or U17558 (N_17558,N_14769,N_11004);
nand U17559 (N_17559,N_11500,N_11543);
nor U17560 (N_17560,N_10834,N_10263);
nor U17561 (N_17561,N_13195,N_13401);
nand U17562 (N_17562,N_13308,N_11495);
or U17563 (N_17563,N_11888,N_13790);
xor U17564 (N_17564,N_12818,N_13385);
or U17565 (N_17565,N_14318,N_11391);
or U17566 (N_17566,N_13889,N_13478);
nand U17567 (N_17567,N_13390,N_13428);
and U17568 (N_17568,N_10846,N_14208);
xor U17569 (N_17569,N_12989,N_11845);
and U17570 (N_17570,N_10722,N_11669);
nor U17571 (N_17571,N_14313,N_13163);
or U17572 (N_17572,N_11314,N_10985);
xnor U17573 (N_17573,N_13208,N_14800);
nor U17574 (N_17574,N_13145,N_10262);
and U17575 (N_17575,N_12076,N_13504);
or U17576 (N_17576,N_13984,N_14052);
and U17577 (N_17577,N_11106,N_12826);
and U17578 (N_17578,N_14498,N_12814);
and U17579 (N_17579,N_10239,N_14351);
nand U17580 (N_17580,N_10480,N_13058);
xnor U17581 (N_17581,N_13313,N_14048);
xor U17582 (N_17582,N_11716,N_12170);
xnor U17583 (N_17583,N_12208,N_11921);
nor U17584 (N_17584,N_13469,N_10468);
xnor U17585 (N_17585,N_10904,N_13275);
nor U17586 (N_17586,N_11632,N_14520);
nor U17587 (N_17587,N_11673,N_14708);
or U17588 (N_17588,N_11322,N_13901);
and U17589 (N_17589,N_14431,N_11153);
nor U17590 (N_17590,N_12097,N_12551);
or U17591 (N_17591,N_12013,N_13167);
or U17592 (N_17592,N_13247,N_11158);
or U17593 (N_17593,N_13923,N_12182);
or U17594 (N_17594,N_11421,N_11671);
and U17595 (N_17595,N_13950,N_10325);
nor U17596 (N_17596,N_12740,N_11454);
xnor U17597 (N_17597,N_13080,N_11405);
nor U17598 (N_17598,N_13237,N_13136);
and U17599 (N_17599,N_11655,N_10628);
xor U17600 (N_17600,N_13587,N_11078);
and U17601 (N_17601,N_12646,N_11726);
nand U17602 (N_17602,N_11360,N_14760);
nand U17603 (N_17603,N_11696,N_13530);
or U17604 (N_17604,N_14493,N_10796);
nor U17605 (N_17605,N_11949,N_12214);
nor U17606 (N_17606,N_14756,N_10714);
nand U17607 (N_17607,N_10316,N_11329);
nand U17608 (N_17608,N_10564,N_11319);
xor U17609 (N_17609,N_11920,N_10066);
xor U17610 (N_17610,N_12622,N_11699);
and U17611 (N_17611,N_13290,N_12726);
or U17612 (N_17612,N_12994,N_14219);
nand U17613 (N_17613,N_11067,N_12369);
nor U17614 (N_17614,N_10716,N_12564);
or U17615 (N_17615,N_11229,N_11984);
or U17616 (N_17616,N_11918,N_10046);
xor U17617 (N_17617,N_10315,N_12207);
xor U17618 (N_17618,N_11588,N_14681);
and U17619 (N_17619,N_13109,N_10258);
nand U17620 (N_17620,N_12797,N_13051);
and U17621 (N_17621,N_14402,N_13896);
or U17622 (N_17622,N_10295,N_14747);
xor U17623 (N_17623,N_14165,N_10425);
and U17624 (N_17624,N_14509,N_10747);
xnor U17625 (N_17625,N_10654,N_12328);
and U17626 (N_17626,N_13830,N_13832);
nand U17627 (N_17627,N_13882,N_14227);
nor U17628 (N_17628,N_14587,N_13658);
nand U17629 (N_17629,N_10410,N_14054);
xor U17630 (N_17630,N_12861,N_13497);
xor U17631 (N_17631,N_11737,N_11694);
and U17632 (N_17632,N_14081,N_11538);
nor U17633 (N_17633,N_12967,N_12112);
or U17634 (N_17634,N_12773,N_10323);
and U17635 (N_17635,N_12636,N_11649);
xor U17636 (N_17636,N_13604,N_12145);
and U17637 (N_17637,N_13300,N_10583);
nor U17638 (N_17638,N_13725,N_14557);
xor U17639 (N_17639,N_10497,N_12923);
nor U17640 (N_17640,N_10289,N_12725);
nand U17641 (N_17641,N_13747,N_13929);
or U17642 (N_17642,N_11474,N_10862);
or U17643 (N_17643,N_12460,N_10444);
and U17644 (N_17644,N_13090,N_10006);
nand U17645 (N_17645,N_12163,N_13495);
or U17646 (N_17646,N_11055,N_11931);
nand U17647 (N_17647,N_14153,N_10870);
xor U17648 (N_17648,N_13542,N_13932);
and U17649 (N_17649,N_13738,N_14763);
xor U17650 (N_17650,N_12892,N_13448);
and U17651 (N_17651,N_10743,N_12363);
or U17652 (N_17652,N_12998,N_11602);
or U17653 (N_17653,N_10162,N_10616);
nand U17654 (N_17654,N_13813,N_10587);
nor U17655 (N_17655,N_10377,N_12324);
or U17656 (N_17656,N_13020,N_11030);
nand U17657 (N_17657,N_14597,N_11370);
and U17658 (N_17658,N_13943,N_13594);
or U17659 (N_17659,N_11552,N_14101);
nor U17660 (N_17660,N_11358,N_11702);
xnor U17661 (N_17661,N_12974,N_10436);
nor U17662 (N_17662,N_12401,N_11851);
or U17663 (N_17663,N_11750,N_13311);
nand U17664 (N_17664,N_12753,N_11677);
nand U17665 (N_17665,N_12217,N_14087);
xnor U17666 (N_17666,N_11124,N_11486);
nor U17667 (N_17667,N_13831,N_12448);
nand U17668 (N_17668,N_13304,N_10005);
or U17669 (N_17669,N_13590,N_12518);
nor U17670 (N_17670,N_11694,N_12308);
nor U17671 (N_17671,N_10267,N_10854);
nand U17672 (N_17672,N_11327,N_13968);
and U17673 (N_17673,N_14811,N_14038);
nand U17674 (N_17674,N_12281,N_10271);
nor U17675 (N_17675,N_14598,N_13875);
nand U17676 (N_17676,N_13339,N_10133);
and U17677 (N_17677,N_12615,N_12540);
and U17678 (N_17678,N_10677,N_13587);
nand U17679 (N_17679,N_12080,N_11885);
nor U17680 (N_17680,N_10474,N_14846);
nor U17681 (N_17681,N_14586,N_10509);
or U17682 (N_17682,N_10351,N_13763);
or U17683 (N_17683,N_11919,N_13933);
nand U17684 (N_17684,N_13303,N_13821);
nor U17685 (N_17685,N_13863,N_10008);
xnor U17686 (N_17686,N_14119,N_12589);
and U17687 (N_17687,N_10502,N_10607);
nand U17688 (N_17688,N_12450,N_11068);
and U17689 (N_17689,N_14095,N_14398);
nand U17690 (N_17690,N_10203,N_10706);
nor U17691 (N_17691,N_10570,N_14503);
and U17692 (N_17692,N_12277,N_11149);
xor U17693 (N_17693,N_11428,N_13323);
or U17694 (N_17694,N_13493,N_11065);
nor U17695 (N_17695,N_12561,N_10725);
nand U17696 (N_17696,N_11710,N_14069);
xnor U17697 (N_17697,N_13568,N_13668);
and U17698 (N_17698,N_13516,N_10442);
nand U17699 (N_17699,N_12271,N_13888);
and U17700 (N_17700,N_12976,N_12477);
or U17701 (N_17701,N_11514,N_11546);
or U17702 (N_17702,N_11810,N_14714);
nand U17703 (N_17703,N_13814,N_13570);
nand U17704 (N_17704,N_10511,N_14438);
nor U17705 (N_17705,N_11317,N_14660);
xnor U17706 (N_17706,N_13938,N_11591);
xnor U17707 (N_17707,N_10857,N_11818);
and U17708 (N_17708,N_10537,N_10936);
xor U17709 (N_17709,N_11697,N_12520);
or U17710 (N_17710,N_13221,N_13404);
and U17711 (N_17711,N_11876,N_11900);
nand U17712 (N_17712,N_12235,N_12889);
nor U17713 (N_17713,N_13496,N_12805);
xor U17714 (N_17714,N_14999,N_12652);
and U17715 (N_17715,N_10685,N_14272);
or U17716 (N_17716,N_13142,N_14535);
nor U17717 (N_17717,N_12957,N_10382);
and U17718 (N_17718,N_12895,N_12683);
or U17719 (N_17719,N_10089,N_10686);
and U17720 (N_17720,N_11977,N_14438);
or U17721 (N_17721,N_14041,N_14080);
and U17722 (N_17722,N_10216,N_14321);
and U17723 (N_17723,N_11880,N_13157);
and U17724 (N_17724,N_12096,N_10376);
or U17725 (N_17725,N_12347,N_11349);
and U17726 (N_17726,N_13956,N_11922);
or U17727 (N_17727,N_14832,N_13368);
nand U17728 (N_17728,N_10121,N_14645);
or U17729 (N_17729,N_14035,N_11066);
and U17730 (N_17730,N_10449,N_11701);
nor U17731 (N_17731,N_10316,N_10462);
and U17732 (N_17732,N_13035,N_14524);
xnor U17733 (N_17733,N_11503,N_10313);
nor U17734 (N_17734,N_14076,N_10869);
nand U17735 (N_17735,N_10236,N_14887);
or U17736 (N_17736,N_14309,N_14710);
and U17737 (N_17737,N_10040,N_10016);
and U17738 (N_17738,N_13340,N_12937);
and U17739 (N_17739,N_11434,N_10041);
nor U17740 (N_17740,N_13536,N_12647);
xnor U17741 (N_17741,N_12004,N_12601);
or U17742 (N_17742,N_14952,N_11140);
xor U17743 (N_17743,N_14404,N_11205);
or U17744 (N_17744,N_14486,N_11264);
xor U17745 (N_17745,N_14184,N_12910);
nand U17746 (N_17746,N_10815,N_10597);
nand U17747 (N_17747,N_10480,N_14521);
or U17748 (N_17748,N_10834,N_12826);
nand U17749 (N_17749,N_12930,N_12102);
or U17750 (N_17750,N_14193,N_12778);
nor U17751 (N_17751,N_10810,N_14509);
nand U17752 (N_17752,N_11957,N_12671);
or U17753 (N_17753,N_14304,N_11709);
nor U17754 (N_17754,N_13898,N_14842);
nand U17755 (N_17755,N_11181,N_14308);
nand U17756 (N_17756,N_12875,N_13125);
nand U17757 (N_17757,N_14690,N_13786);
or U17758 (N_17758,N_11804,N_13498);
xor U17759 (N_17759,N_10641,N_14033);
or U17760 (N_17760,N_11133,N_13689);
and U17761 (N_17761,N_14155,N_13454);
xor U17762 (N_17762,N_12897,N_10332);
and U17763 (N_17763,N_13513,N_13697);
and U17764 (N_17764,N_14349,N_14954);
or U17765 (N_17765,N_13666,N_14332);
or U17766 (N_17766,N_14207,N_14270);
and U17767 (N_17767,N_10962,N_11456);
and U17768 (N_17768,N_14191,N_13609);
or U17769 (N_17769,N_12540,N_12309);
nor U17770 (N_17770,N_12079,N_14954);
and U17771 (N_17771,N_13422,N_10804);
nand U17772 (N_17772,N_13347,N_14988);
and U17773 (N_17773,N_13559,N_14022);
nand U17774 (N_17774,N_11914,N_12820);
nor U17775 (N_17775,N_10448,N_12819);
nor U17776 (N_17776,N_10307,N_12812);
and U17777 (N_17777,N_12110,N_11676);
or U17778 (N_17778,N_13561,N_14997);
nand U17779 (N_17779,N_13340,N_13003);
and U17780 (N_17780,N_10115,N_14604);
nand U17781 (N_17781,N_13395,N_10457);
nand U17782 (N_17782,N_13080,N_13360);
xnor U17783 (N_17783,N_10581,N_14261);
xor U17784 (N_17784,N_10262,N_14451);
or U17785 (N_17785,N_14813,N_13005);
and U17786 (N_17786,N_11294,N_10796);
nor U17787 (N_17787,N_14598,N_12143);
nor U17788 (N_17788,N_14213,N_14505);
nand U17789 (N_17789,N_10795,N_12894);
or U17790 (N_17790,N_11818,N_12147);
nand U17791 (N_17791,N_10840,N_10265);
or U17792 (N_17792,N_14189,N_14111);
nand U17793 (N_17793,N_11016,N_11573);
or U17794 (N_17794,N_10039,N_12276);
nand U17795 (N_17795,N_11914,N_10015);
nor U17796 (N_17796,N_14337,N_14804);
or U17797 (N_17797,N_11082,N_12544);
nand U17798 (N_17798,N_12076,N_10986);
nand U17799 (N_17799,N_13637,N_14688);
or U17800 (N_17800,N_11368,N_11797);
nor U17801 (N_17801,N_11603,N_12663);
and U17802 (N_17802,N_13039,N_12452);
xnor U17803 (N_17803,N_13078,N_13541);
and U17804 (N_17804,N_14744,N_10179);
and U17805 (N_17805,N_10733,N_10856);
nand U17806 (N_17806,N_14198,N_14034);
or U17807 (N_17807,N_11813,N_10502);
nand U17808 (N_17808,N_12469,N_11132);
xor U17809 (N_17809,N_13291,N_10069);
nor U17810 (N_17810,N_10832,N_12534);
or U17811 (N_17811,N_11821,N_13174);
xor U17812 (N_17812,N_10020,N_11520);
nor U17813 (N_17813,N_13473,N_13153);
and U17814 (N_17814,N_11368,N_13722);
nand U17815 (N_17815,N_11297,N_12261);
xor U17816 (N_17816,N_14706,N_14064);
nor U17817 (N_17817,N_14724,N_11705);
and U17818 (N_17818,N_11371,N_14473);
or U17819 (N_17819,N_12954,N_10101);
xnor U17820 (N_17820,N_13112,N_14604);
xor U17821 (N_17821,N_10950,N_11905);
nand U17822 (N_17822,N_13355,N_10021);
nand U17823 (N_17823,N_12388,N_12802);
xnor U17824 (N_17824,N_11433,N_11843);
or U17825 (N_17825,N_11408,N_13694);
nor U17826 (N_17826,N_10969,N_14887);
nand U17827 (N_17827,N_10489,N_11048);
or U17828 (N_17828,N_13826,N_11206);
nand U17829 (N_17829,N_10478,N_12900);
xnor U17830 (N_17830,N_12346,N_10062);
or U17831 (N_17831,N_12784,N_11604);
nand U17832 (N_17832,N_10876,N_13159);
nor U17833 (N_17833,N_12566,N_10586);
or U17834 (N_17834,N_13412,N_10445);
xor U17835 (N_17835,N_11967,N_14535);
nor U17836 (N_17836,N_14481,N_10639);
xor U17837 (N_17837,N_13106,N_13320);
xnor U17838 (N_17838,N_10512,N_12796);
or U17839 (N_17839,N_12097,N_12508);
and U17840 (N_17840,N_14546,N_12064);
or U17841 (N_17841,N_14213,N_11370);
nor U17842 (N_17842,N_12479,N_10787);
xnor U17843 (N_17843,N_12680,N_12910);
or U17844 (N_17844,N_11127,N_11662);
xor U17845 (N_17845,N_14487,N_14747);
or U17846 (N_17846,N_14793,N_13095);
or U17847 (N_17847,N_12810,N_13526);
nor U17848 (N_17848,N_11876,N_10800);
xor U17849 (N_17849,N_12295,N_11610);
and U17850 (N_17850,N_10610,N_14339);
nor U17851 (N_17851,N_13411,N_11776);
nand U17852 (N_17852,N_10431,N_11512);
nand U17853 (N_17853,N_13082,N_12510);
xor U17854 (N_17854,N_13706,N_10075);
nand U17855 (N_17855,N_13856,N_14966);
nand U17856 (N_17856,N_12881,N_12802);
or U17857 (N_17857,N_14790,N_10611);
nor U17858 (N_17858,N_12176,N_13463);
nor U17859 (N_17859,N_11513,N_12289);
xnor U17860 (N_17860,N_13709,N_14253);
and U17861 (N_17861,N_13859,N_14929);
xnor U17862 (N_17862,N_14999,N_12184);
nor U17863 (N_17863,N_14964,N_11793);
or U17864 (N_17864,N_10661,N_14533);
nand U17865 (N_17865,N_12083,N_13236);
nand U17866 (N_17866,N_12642,N_13346);
xnor U17867 (N_17867,N_10327,N_14780);
or U17868 (N_17868,N_11366,N_14955);
or U17869 (N_17869,N_14897,N_14129);
and U17870 (N_17870,N_12497,N_12964);
xor U17871 (N_17871,N_11148,N_11817);
or U17872 (N_17872,N_11298,N_14177);
nor U17873 (N_17873,N_14001,N_13774);
and U17874 (N_17874,N_14361,N_12025);
xnor U17875 (N_17875,N_13252,N_11693);
or U17876 (N_17876,N_14198,N_11153);
xnor U17877 (N_17877,N_13694,N_11166);
xor U17878 (N_17878,N_13530,N_13468);
xnor U17879 (N_17879,N_11564,N_13591);
and U17880 (N_17880,N_13696,N_12111);
nor U17881 (N_17881,N_10204,N_10552);
or U17882 (N_17882,N_10953,N_13023);
nand U17883 (N_17883,N_14980,N_11691);
or U17884 (N_17884,N_11429,N_13687);
or U17885 (N_17885,N_14381,N_12435);
nand U17886 (N_17886,N_12405,N_11722);
xnor U17887 (N_17887,N_13012,N_11839);
nor U17888 (N_17888,N_11596,N_10044);
nor U17889 (N_17889,N_14072,N_11813);
and U17890 (N_17890,N_12469,N_10328);
nor U17891 (N_17891,N_10538,N_14957);
nand U17892 (N_17892,N_14778,N_12205);
nand U17893 (N_17893,N_14009,N_11786);
xnor U17894 (N_17894,N_11111,N_11794);
nor U17895 (N_17895,N_13244,N_12107);
xnor U17896 (N_17896,N_12408,N_14674);
nor U17897 (N_17897,N_12352,N_13003);
and U17898 (N_17898,N_11439,N_10969);
nor U17899 (N_17899,N_14629,N_14839);
nor U17900 (N_17900,N_10448,N_12688);
nand U17901 (N_17901,N_14935,N_10538);
nand U17902 (N_17902,N_11259,N_12354);
xnor U17903 (N_17903,N_10042,N_10427);
and U17904 (N_17904,N_11623,N_10915);
nand U17905 (N_17905,N_14332,N_10195);
nor U17906 (N_17906,N_11717,N_14259);
nor U17907 (N_17907,N_10874,N_13257);
and U17908 (N_17908,N_14146,N_13158);
nand U17909 (N_17909,N_11026,N_11185);
nor U17910 (N_17910,N_14656,N_14179);
and U17911 (N_17911,N_10992,N_10659);
nand U17912 (N_17912,N_11656,N_10778);
xnor U17913 (N_17913,N_13882,N_10922);
and U17914 (N_17914,N_11828,N_10370);
xor U17915 (N_17915,N_10726,N_12449);
nor U17916 (N_17916,N_11326,N_12178);
and U17917 (N_17917,N_10105,N_11502);
xor U17918 (N_17918,N_11348,N_11641);
or U17919 (N_17919,N_11539,N_13141);
nor U17920 (N_17920,N_12912,N_14488);
nand U17921 (N_17921,N_13391,N_10280);
xnor U17922 (N_17922,N_14472,N_13223);
nor U17923 (N_17923,N_13470,N_13165);
xor U17924 (N_17924,N_13944,N_12889);
nand U17925 (N_17925,N_10823,N_13965);
xnor U17926 (N_17926,N_13272,N_11316);
and U17927 (N_17927,N_12205,N_13247);
xor U17928 (N_17928,N_14559,N_12219);
nand U17929 (N_17929,N_10781,N_12349);
or U17930 (N_17930,N_11082,N_12487);
and U17931 (N_17931,N_14211,N_10712);
or U17932 (N_17932,N_12044,N_14920);
nand U17933 (N_17933,N_12390,N_12527);
xor U17934 (N_17934,N_14311,N_11069);
and U17935 (N_17935,N_10869,N_12874);
nand U17936 (N_17936,N_10124,N_11048);
and U17937 (N_17937,N_14319,N_12214);
and U17938 (N_17938,N_10416,N_13295);
and U17939 (N_17939,N_12282,N_12693);
and U17940 (N_17940,N_13221,N_11683);
nor U17941 (N_17941,N_10864,N_13509);
and U17942 (N_17942,N_11943,N_10133);
nand U17943 (N_17943,N_13550,N_13497);
or U17944 (N_17944,N_11547,N_13351);
or U17945 (N_17945,N_14326,N_11803);
nor U17946 (N_17946,N_14906,N_11887);
xor U17947 (N_17947,N_11718,N_12761);
and U17948 (N_17948,N_10962,N_12038);
or U17949 (N_17949,N_14426,N_11250);
nand U17950 (N_17950,N_13971,N_14835);
nand U17951 (N_17951,N_10489,N_14549);
nand U17952 (N_17952,N_12635,N_13578);
nand U17953 (N_17953,N_12581,N_10060);
nor U17954 (N_17954,N_13841,N_13147);
nand U17955 (N_17955,N_12071,N_14320);
and U17956 (N_17956,N_13725,N_13438);
or U17957 (N_17957,N_12413,N_14614);
xor U17958 (N_17958,N_14817,N_12081);
nand U17959 (N_17959,N_11452,N_10961);
nand U17960 (N_17960,N_13306,N_10118);
nor U17961 (N_17961,N_10949,N_10011);
and U17962 (N_17962,N_13658,N_11430);
and U17963 (N_17963,N_13661,N_10666);
xnor U17964 (N_17964,N_10196,N_12331);
xor U17965 (N_17965,N_14110,N_11802);
xnor U17966 (N_17966,N_13352,N_13063);
xnor U17967 (N_17967,N_12436,N_13386);
xor U17968 (N_17968,N_12211,N_10320);
or U17969 (N_17969,N_14011,N_12360);
nor U17970 (N_17970,N_12272,N_11135);
nor U17971 (N_17971,N_10179,N_12386);
xnor U17972 (N_17972,N_11092,N_14902);
or U17973 (N_17973,N_11625,N_12244);
nor U17974 (N_17974,N_12826,N_11484);
and U17975 (N_17975,N_11493,N_10056);
or U17976 (N_17976,N_12321,N_10839);
and U17977 (N_17977,N_13114,N_10284);
and U17978 (N_17978,N_14392,N_11610);
xnor U17979 (N_17979,N_14121,N_11735);
xnor U17980 (N_17980,N_14234,N_14421);
or U17981 (N_17981,N_10236,N_14538);
nand U17982 (N_17982,N_11319,N_10788);
xor U17983 (N_17983,N_13659,N_11826);
xor U17984 (N_17984,N_14407,N_14919);
and U17985 (N_17985,N_14770,N_10802);
nand U17986 (N_17986,N_13436,N_12584);
or U17987 (N_17987,N_14662,N_12632);
xor U17988 (N_17988,N_14503,N_11668);
or U17989 (N_17989,N_11290,N_12292);
and U17990 (N_17990,N_11639,N_14075);
nor U17991 (N_17991,N_13778,N_14054);
or U17992 (N_17992,N_14777,N_12407);
or U17993 (N_17993,N_13417,N_11281);
xor U17994 (N_17994,N_10922,N_14413);
nor U17995 (N_17995,N_11664,N_13459);
nand U17996 (N_17996,N_10340,N_11321);
and U17997 (N_17997,N_10125,N_11916);
xnor U17998 (N_17998,N_13969,N_13791);
and U17999 (N_17999,N_13067,N_11410);
and U18000 (N_18000,N_12571,N_14646);
xor U18001 (N_18001,N_12233,N_13203);
xor U18002 (N_18002,N_12742,N_11108);
xor U18003 (N_18003,N_13505,N_14210);
nand U18004 (N_18004,N_14455,N_14682);
nor U18005 (N_18005,N_13421,N_14294);
nand U18006 (N_18006,N_13839,N_11418);
nand U18007 (N_18007,N_11821,N_13281);
nor U18008 (N_18008,N_10599,N_12699);
nor U18009 (N_18009,N_10811,N_14422);
and U18010 (N_18010,N_14810,N_11577);
nor U18011 (N_18011,N_14041,N_12820);
xnor U18012 (N_18012,N_10134,N_11027);
xnor U18013 (N_18013,N_14003,N_14536);
nand U18014 (N_18014,N_12251,N_11832);
nor U18015 (N_18015,N_12064,N_12085);
nand U18016 (N_18016,N_11907,N_10332);
and U18017 (N_18017,N_10519,N_10753);
and U18018 (N_18018,N_12506,N_10044);
and U18019 (N_18019,N_13362,N_10342);
xor U18020 (N_18020,N_12458,N_12727);
nand U18021 (N_18021,N_14769,N_14792);
or U18022 (N_18022,N_14768,N_14483);
xor U18023 (N_18023,N_13290,N_11528);
xnor U18024 (N_18024,N_14997,N_13837);
xor U18025 (N_18025,N_14574,N_14638);
xor U18026 (N_18026,N_10591,N_11551);
nand U18027 (N_18027,N_11391,N_13495);
nor U18028 (N_18028,N_10459,N_10085);
or U18029 (N_18029,N_13132,N_14239);
xor U18030 (N_18030,N_12570,N_11791);
or U18031 (N_18031,N_11953,N_13389);
and U18032 (N_18032,N_14187,N_13945);
nor U18033 (N_18033,N_10072,N_14872);
nor U18034 (N_18034,N_11465,N_13572);
xnor U18035 (N_18035,N_10936,N_14335);
nand U18036 (N_18036,N_11282,N_12557);
xor U18037 (N_18037,N_13878,N_13824);
or U18038 (N_18038,N_10801,N_10846);
nor U18039 (N_18039,N_11444,N_14993);
xnor U18040 (N_18040,N_13163,N_12074);
nand U18041 (N_18041,N_12037,N_13380);
and U18042 (N_18042,N_13226,N_11472);
and U18043 (N_18043,N_11744,N_13215);
xor U18044 (N_18044,N_10481,N_12157);
xnor U18045 (N_18045,N_12056,N_13450);
or U18046 (N_18046,N_13784,N_12353);
or U18047 (N_18047,N_10513,N_11950);
or U18048 (N_18048,N_14643,N_13960);
or U18049 (N_18049,N_14808,N_14787);
nand U18050 (N_18050,N_11512,N_12986);
nand U18051 (N_18051,N_10112,N_11946);
or U18052 (N_18052,N_13287,N_10130);
xnor U18053 (N_18053,N_13531,N_12260);
nor U18054 (N_18054,N_13243,N_11449);
xnor U18055 (N_18055,N_14868,N_12020);
or U18056 (N_18056,N_13010,N_14637);
nor U18057 (N_18057,N_11142,N_14971);
and U18058 (N_18058,N_13124,N_11854);
nor U18059 (N_18059,N_12635,N_14215);
and U18060 (N_18060,N_11624,N_11276);
nor U18061 (N_18061,N_14999,N_12561);
and U18062 (N_18062,N_14451,N_13766);
xor U18063 (N_18063,N_13725,N_11423);
nand U18064 (N_18064,N_12653,N_12918);
and U18065 (N_18065,N_11006,N_12456);
nand U18066 (N_18066,N_11771,N_12262);
xnor U18067 (N_18067,N_11726,N_13602);
or U18068 (N_18068,N_14599,N_11802);
nand U18069 (N_18069,N_11137,N_14400);
and U18070 (N_18070,N_10703,N_12184);
and U18071 (N_18071,N_10436,N_11640);
or U18072 (N_18072,N_12513,N_11370);
xor U18073 (N_18073,N_13986,N_11629);
nand U18074 (N_18074,N_13562,N_14361);
nor U18075 (N_18075,N_10643,N_12616);
and U18076 (N_18076,N_11941,N_12884);
and U18077 (N_18077,N_14107,N_11703);
nor U18078 (N_18078,N_12744,N_14257);
or U18079 (N_18079,N_14257,N_10392);
and U18080 (N_18080,N_10634,N_12490);
xnor U18081 (N_18081,N_14072,N_11156);
nor U18082 (N_18082,N_13955,N_12549);
or U18083 (N_18083,N_12740,N_11580);
nand U18084 (N_18084,N_14842,N_10921);
and U18085 (N_18085,N_13959,N_10705);
nand U18086 (N_18086,N_12894,N_13938);
xor U18087 (N_18087,N_13833,N_12916);
or U18088 (N_18088,N_11019,N_14467);
and U18089 (N_18089,N_12155,N_13942);
nor U18090 (N_18090,N_10610,N_11993);
nor U18091 (N_18091,N_11904,N_10056);
nor U18092 (N_18092,N_12419,N_10079);
nand U18093 (N_18093,N_13371,N_10223);
xor U18094 (N_18094,N_12466,N_14274);
and U18095 (N_18095,N_10985,N_14615);
nand U18096 (N_18096,N_14259,N_12399);
nand U18097 (N_18097,N_12169,N_10833);
or U18098 (N_18098,N_10765,N_14949);
xor U18099 (N_18099,N_14859,N_14768);
nor U18100 (N_18100,N_10819,N_10343);
or U18101 (N_18101,N_14564,N_14750);
nor U18102 (N_18102,N_12943,N_14012);
nor U18103 (N_18103,N_14803,N_14931);
and U18104 (N_18104,N_14970,N_13555);
and U18105 (N_18105,N_13302,N_14666);
or U18106 (N_18106,N_13913,N_12345);
nand U18107 (N_18107,N_12645,N_10681);
nor U18108 (N_18108,N_10679,N_10473);
nor U18109 (N_18109,N_11112,N_11978);
nand U18110 (N_18110,N_13483,N_13669);
xor U18111 (N_18111,N_10877,N_12166);
nand U18112 (N_18112,N_12391,N_13598);
nand U18113 (N_18113,N_11151,N_13813);
and U18114 (N_18114,N_11532,N_10252);
and U18115 (N_18115,N_13790,N_14412);
nor U18116 (N_18116,N_11411,N_12999);
xor U18117 (N_18117,N_13821,N_14761);
nor U18118 (N_18118,N_11263,N_14699);
and U18119 (N_18119,N_10402,N_11688);
xor U18120 (N_18120,N_12353,N_11407);
or U18121 (N_18121,N_10958,N_11462);
xor U18122 (N_18122,N_12777,N_13140);
xor U18123 (N_18123,N_11975,N_13552);
nand U18124 (N_18124,N_10818,N_14460);
nand U18125 (N_18125,N_12851,N_10895);
nand U18126 (N_18126,N_14475,N_10523);
nor U18127 (N_18127,N_12406,N_14355);
nand U18128 (N_18128,N_11456,N_14818);
nor U18129 (N_18129,N_13037,N_14177);
nor U18130 (N_18130,N_10603,N_10509);
nor U18131 (N_18131,N_11506,N_11083);
nor U18132 (N_18132,N_11883,N_14928);
nand U18133 (N_18133,N_11760,N_12910);
xnor U18134 (N_18134,N_13827,N_14430);
nand U18135 (N_18135,N_14267,N_13262);
xnor U18136 (N_18136,N_12169,N_12381);
nor U18137 (N_18137,N_10746,N_11489);
and U18138 (N_18138,N_12520,N_14387);
or U18139 (N_18139,N_14934,N_13674);
xnor U18140 (N_18140,N_13776,N_10956);
and U18141 (N_18141,N_14460,N_10693);
xor U18142 (N_18142,N_12334,N_14522);
or U18143 (N_18143,N_10700,N_12363);
nor U18144 (N_18144,N_14619,N_10571);
nor U18145 (N_18145,N_14605,N_13175);
or U18146 (N_18146,N_12226,N_14429);
and U18147 (N_18147,N_14270,N_13075);
nand U18148 (N_18148,N_12284,N_10189);
nand U18149 (N_18149,N_13385,N_11390);
or U18150 (N_18150,N_10149,N_11739);
nand U18151 (N_18151,N_14500,N_10621);
or U18152 (N_18152,N_12513,N_12399);
and U18153 (N_18153,N_13621,N_10231);
nor U18154 (N_18154,N_14050,N_11952);
nor U18155 (N_18155,N_10809,N_13249);
or U18156 (N_18156,N_14986,N_10759);
nor U18157 (N_18157,N_10988,N_11567);
and U18158 (N_18158,N_13511,N_10317);
xor U18159 (N_18159,N_10942,N_10041);
xor U18160 (N_18160,N_14157,N_12037);
xor U18161 (N_18161,N_12803,N_14464);
xor U18162 (N_18162,N_14606,N_14246);
nand U18163 (N_18163,N_13403,N_11850);
nand U18164 (N_18164,N_12807,N_12745);
nor U18165 (N_18165,N_14616,N_13420);
and U18166 (N_18166,N_14075,N_10114);
nor U18167 (N_18167,N_12544,N_12768);
or U18168 (N_18168,N_10412,N_10335);
nor U18169 (N_18169,N_10591,N_10952);
nand U18170 (N_18170,N_14060,N_13404);
nand U18171 (N_18171,N_13012,N_13268);
xnor U18172 (N_18172,N_14231,N_14348);
or U18173 (N_18173,N_12780,N_13296);
or U18174 (N_18174,N_12635,N_13872);
or U18175 (N_18175,N_13432,N_13569);
and U18176 (N_18176,N_10945,N_10553);
xor U18177 (N_18177,N_10020,N_11996);
nand U18178 (N_18178,N_12763,N_13710);
nor U18179 (N_18179,N_10792,N_13581);
nand U18180 (N_18180,N_13457,N_14719);
nand U18181 (N_18181,N_11032,N_14155);
nor U18182 (N_18182,N_12814,N_12779);
and U18183 (N_18183,N_13376,N_14313);
xnor U18184 (N_18184,N_11602,N_10971);
and U18185 (N_18185,N_14457,N_10448);
nor U18186 (N_18186,N_14888,N_12604);
xor U18187 (N_18187,N_11160,N_14196);
nor U18188 (N_18188,N_10518,N_14117);
xnor U18189 (N_18189,N_13267,N_14309);
xor U18190 (N_18190,N_14428,N_11933);
and U18191 (N_18191,N_12701,N_11727);
nor U18192 (N_18192,N_11303,N_14366);
and U18193 (N_18193,N_13698,N_14712);
and U18194 (N_18194,N_10716,N_10215);
xnor U18195 (N_18195,N_14810,N_13335);
nor U18196 (N_18196,N_13593,N_12360);
xnor U18197 (N_18197,N_12927,N_11744);
and U18198 (N_18198,N_12504,N_11118);
or U18199 (N_18199,N_11250,N_10384);
and U18200 (N_18200,N_10908,N_11047);
nand U18201 (N_18201,N_13456,N_10625);
or U18202 (N_18202,N_10836,N_12135);
nand U18203 (N_18203,N_12314,N_12755);
nand U18204 (N_18204,N_14797,N_12658);
or U18205 (N_18205,N_13104,N_12567);
or U18206 (N_18206,N_13948,N_12246);
nand U18207 (N_18207,N_12661,N_14817);
or U18208 (N_18208,N_13817,N_12994);
nand U18209 (N_18209,N_11888,N_12587);
or U18210 (N_18210,N_14646,N_13560);
xor U18211 (N_18211,N_13815,N_14127);
nand U18212 (N_18212,N_12232,N_12539);
xnor U18213 (N_18213,N_13744,N_14269);
or U18214 (N_18214,N_14175,N_10115);
or U18215 (N_18215,N_11221,N_12759);
nand U18216 (N_18216,N_12737,N_13530);
and U18217 (N_18217,N_10680,N_10979);
or U18218 (N_18218,N_13603,N_13852);
nor U18219 (N_18219,N_10598,N_14609);
or U18220 (N_18220,N_13035,N_14487);
and U18221 (N_18221,N_14554,N_13534);
nand U18222 (N_18222,N_13602,N_12764);
and U18223 (N_18223,N_11511,N_14843);
nor U18224 (N_18224,N_14189,N_12742);
xor U18225 (N_18225,N_12864,N_12013);
nor U18226 (N_18226,N_14613,N_10857);
and U18227 (N_18227,N_13372,N_11808);
and U18228 (N_18228,N_13407,N_14578);
and U18229 (N_18229,N_13586,N_12602);
nand U18230 (N_18230,N_13105,N_14382);
or U18231 (N_18231,N_12761,N_13591);
nor U18232 (N_18232,N_11047,N_12775);
nor U18233 (N_18233,N_14970,N_14944);
xnor U18234 (N_18234,N_12429,N_14383);
or U18235 (N_18235,N_13088,N_12983);
xnor U18236 (N_18236,N_10157,N_14617);
and U18237 (N_18237,N_10679,N_12723);
or U18238 (N_18238,N_12761,N_12312);
and U18239 (N_18239,N_14630,N_11314);
or U18240 (N_18240,N_14660,N_13740);
nor U18241 (N_18241,N_14957,N_13138);
nand U18242 (N_18242,N_13639,N_12233);
nor U18243 (N_18243,N_14326,N_12083);
xor U18244 (N_18244,N_10750,N_12116);
and U18245 (N_18245,N_11988,N_12102);
nor U18246 (N_18246,N_11765,N_13584);
nand U18247 (N_18247,N_14940,N_12003);
and U18248 (N_18248,N_11491,N_14428);
nand U18249 (N_18249,N_11809,N_10157);
nand U18250 (N_18250,N_10842,N_14459);
and U18251 (N_18251,N_11949,N_13967);
or U18252 (N_18252,N_14155,N_14089);
xor U18253 (N_18253,N_10442,N_13664);
and U18254 (N_18254,N_10069,N_10827);
nand U18255 (N_18255,N_12170,N_10546);
or U18256 (N_18256,N_11755,N_13531);
or U18257 (N_18257,N_13847,N_10609);
xor U18258 (N_18258,N_13596,N_12444);
or U18259 (N_18259,N_13936,N_14833);
xnor U18260 (N_18260,N_14634,N_10955);
xor U18261 (N_18261,N_10413,N_10997);
and U18262 (N_18262,N_12656,N_12873);
xnor U18263 (N_18263,N_11465,N_13110);
or U18264 (N_18264,N_14595,N_10876);
xor U18265 (N_18265,N_13152,N_13779);
and U18266 (N_18266,N_11536,N_14464);
nand U18267 (N_18267,N_14272,N_14051);
and U18268 (N_18268,N_10169,N_11672);
and U18269 (N_18269,N_10466,N_12804);
nand U18270 (N_18270,N_14354,N_14673);
nand U18271 (N_18271,N_13490,N_12574);
or U18272 (N_18272,N_12218,N_10416);
or U18273 (N_18273,N_12323,N_13953);
xnor U18274 (N_18274,N_11943,N_10388);
nor U18275 (N_18275,N_12581,N_11751);
and U18276 (N_18276,N_11057,N_11284);
or U18277 (N_18277,N_13274,N_14461);
and U18278 (N_18278,N_10287,N_10441);
xnor U18279 (N_18279,N_11805,N_12495);
or U18280 (N_18280,N_14006,N_11810);
or U18281 (N_18281,N_14016,N_12686);
nor U18282 (N_18282,N_11341,N_13409);
or U18283 (N_18283,N_11541,N_10482);
and U18284 (N_18284,N_13595,N_11638);
and U18285 (N_18285,N_11631,N_12917);
xor U18286 (N_18286,N_13551,N_11973);
xor U18287 (N_18287,N_12488,N_14048);
and U18288 (N_18288,N_12635,N_13412);
nand U18289 (N_18289,N_14145,N_14002);
and U18290 (N_18290,N_13483,N_12966);
xnor U18291 (N_18291,N_11278,N_11399);
and U18292 (N_18292,N_11844,N_14926);
or U18293 (N_18293,N_13538,N_12329);
nor U18294 (N_18294,N_11598,N_11826);
nand U18295 (N_18295,N_14560,N_14096);
nor U18296 (N_18296,N_10543,N_13833);
xor U18297 (N_18297,N_10038,N_14651);
nor U18298 (N_18298,N_13876,N_11633);
or U18299 (N_18299,N_12215,N_11805);
nand U18300 (N_18300,N_11179,N_10030);
xnor U18301 (N_18301,N_13565,N_11538);
nand U18302 (N_18302,N_12831,N_13388);
xnor U18303 (N_18303,N_13110,N_11475);
xor U18304 (N_18304,N_11781,N_13718);
and U18305 (N_18305,N_13553,N_12362);
nand U18306 (N_18306,N_14042,N_12318);
or U18307 (N_18307,N_11151,N_13583);
nor U18308 (N_18308,N_10484,N_13080);
and U18309 (N_18309,N_10873,N_14828);
or U18310 (N_18310,N_10216,N_13670);
nor U18311 (N_18311,N_11495,N_10932);
xor U18312 (N_18312,N_12961,N_10966);
nand U18313 (N_18313,N_12759,N_13499);
or U18314 (N_18314,N_13908,N_12214);
or U18315 (N_18315,N_14049,N_10238);
nand U18316 (N_18316,N_12294,N_10360);
and U18317 (N_18317,N_10017,N_14720);
nor U18318 (N_18318,N_10648,N_12657);
nor U18319 (N_18319,N_12227,N_13081);
nand U18320 (N_18320,N_12609,N_11377);
and U18321 (N_18321,N_13893,N_13622);
nor U18322 (N_18322,N_13777,N_13392);
nand U18323 (N_18323,N_14222,N_11729);
nor U18324 (N_18324,N_13667,N_12904);
and U18325 (N_18325,N_11705,N_12566);
or U18326 (N_18326,N_14787,N_14609);
or U18327 (N_18327,N_14716,N_11063);
xor U18328 (N_18328,N_10630,N_13931);
or U18329 (N_18329,N_14025,N_13738);
xnor U18330 (N_18330,N_11312,N_12679);
or U18331 (N_18331,N_13124,N_10311);
nor U18332 (N_18332,N_12584,N_12037);
nand U18333 (N_18333,N_10868,N_14659);
nand U18334 (N_18334,N_10678,N_14901);
or U18335 (N_18335,N_13696,N_11317);
nand U18336 (N_18336,N_14764,N_14340);
nand U18337 (N_18337,N_10794,N_13307);
xnor U18338 (N_18338,N_12471,N_13031);
nand U18339 (N_18339,N_10142,N_14123);
nand U18340 (N_18340,N_14777,N_14119);
nand U18341 (N_18341,N_12404,N_12622);
nor U18342 (N_18342,N_11378,N_13268);
xnor U18343 (N_18343,N_13584,N_12428);
xnor U18344 (N_18344,N_14094,N_11349);
or U18345 (N_18345,N_11259,N_13118);
and U18346 (N_18346,N_11772,N_14333);
or U18347 (N_18347,N_10469,N_12601);
and U18348 (N_18348,N_12789,N_14874);
xnor U18349 (N_18349,N_12047,N_13985);
nor U18350 (N_18350,N_12980,N_10218);
nand U18351 (N_18351,N_11256,N_10018);
xor U18352 (N_18352,N_13888,N_10790);
or U18353 (N_18353,N_13865,N_10103);
nand U18354 (N_18354,N_13696,N_11740);
nand U18355 (N_18355,N_14948,N_13574);
or U18356 (N_18356,N_14400,N_14812);
xnor U18357 (N_18357,N_14659,N_11259);
or U18358 (N_18358,N_11696,N_11814);
nor U18359 (N_18359,N_14228,N_12619);
nand U18360 (N_18360,N_11909,N_11185);
nand U18361 (N_18361,N_13014,N_11112);
xnor U18362 (N_18362,N_11854,N_13854);
xnor U18363 (N_18363,N_14148,N_14383);
or U18364 (N_18364,N_13912,N_12106);
xor U18365 (N_18365,N_13018,N_13224);
nand U18366 (N_18366,N_14838,N_14351);
nand U18367 (N_18367,N_10943,N_10773);
nor U18368 (N_18368,N_14740,N_11731);
nand U18369 (N_18369,N_11630,N_14729);
and U18370 (N_18370,N_12553,N_13287);
or U18371 (N_18371,N_13071,N_11817);
or U18372 (N_18372,N_11998,N_13735);
nand U18373 (N_18373,N_10058,N_10893);
or U18374 (N_18374,N_14180,N_10744);
xor U18375 (N_18375,N_10888,N_12265);
xnor U18376 (N_18376,N_13053,N_11547);
nor U18377 (N_18377,N_12923,N_13428);
xor U18378 (N_18378,N_12434,N_14502);
or U18379 (N_18379,N_14899,N_12367);
nand U18380 (N_18380,N_12892,N_12897);
nor U18381 (N_18381,N_10505,N_11111);
and U18382 (N_18382,N_11427,N_14608);
nor U18383 (N_18383,N_10907,N_14181);
and U18384 (N_18384,N_14637,N_10215);
nand U18385 (N_18385,N_12771,N_14214);
nor U18386 (N_18386,N_13159,N_12576);
and U18387 (N_18387,N_11263,N_13091);
xor U18388 (N_18388,N_12357,N_12944);
and U18389 (N_18389,N_13177,N_12484);
and U18390 (N_18390,N_11555,N_11890);
or U18391 (N_18391,N_14989,N_12813);
nor U18392 (N_18392,N_12069,N_11677);
nor U18393 (N_18393,N_12047,N_10773);
nand U18394 (N_18394,N_11582,N_14122);
nor U18395 (N_18395,N_14605,N_10798);
xor U18396 (N_18396,N_14761,N_13184);
or U18397 (N_18397,N_10894,N_13230);
and U18398 (N_18398,N_11799,N_12920);
nor U18399 (N_18399,N_12650,N_13929);
nor U18400 (N_18400,N_14814,N_13746);
xor U18401 (N_18401,N_11276,N_12150);
nand U18402 (N_18402,N_11785,N_10783);
xor U18403 (N_18403,N_11724,N_12976);
or U18404 (N_18404,N_14308,N_14884);
xnor U18405 (N_18405,N_10375,N_10546);
or U18406 (N_18406,N_12017,N_13329);
or U18407 (N_18407,N_12508,N_10665);
xor U18408 (N_18408,N_11597,N_12487);
nor U18409 (N_18409,N_12785,N_10138);
xnor U18410 (N_18410,N_12385,N_11232);
nor U18411 (N_18411,N_14015,N_10231);
and U18412 (N_18412,N_14136,N_13895);
and U18413 (N_18413,N_11034,N_11792);
xor U18414 (N_18414,N_12398,N_13632);
nand U18415 (N_18415,N_11754,N_10622);
and U18416 (N_18416,N_13608,N_14383);
xor U18417 (N_18417,N_13368,N_10576);
or U18418 (N_18418,N_14965,N_12307);
or U18419 (N_18419,N_12049,N_12025);
nor U18420 (N_18420,N_13872,N_10440);
and U18421 (N_18421,N_14967,N_10494);
or U18422 (N_18422,N_14243,N_12708);
nor U18423 (N_18423,N_11714,N_14176);
or U18424 (N_18424,N_11744,N_11743);
xnor U18425 (N_18425,N_12109,N_10387);
xnor U18426 (N_18426,N_11821,N_12648);
xor U18427 (N_18427,N_13164,N_11497);
nor U18428 (N_18428,N_14841,N_10607);
nor U18429 (N_18429,N_13209,N_10525);
or U18430 (N_18430,N_12462,N_13428);
xor U18431 (N_18431,N_10290,N_10306);
and U18432 (N_18432,N_10241,N_12939);
nor U18433 (N_18433,N_14536,N_13458);
xor U18434 (N_18434,N_12005,N_12900);
xnor U18435 (N_18435,N_11199,N_14158);
and U18436 (N_18436,N_12700,N_11951);
and U18437 (N_18437,N_11968,N_12818);
nand U18438 (N_18438,N_11623,N_13192);
or U18439 (N_18439,N_12529,N_10519);
nand U18440 (N_18440,N_12351,N_14009);
nor U18441 (N_18441,N_13459,N_13274);
nand U18442 (N_18442,N_13419,N_12815);
or U18443 (N_18443,N_13383,N_10279);
xor U18444 (N_18444,N_14344,N_11224);
or U18445 (N_18445,N_10918,N_12364);
xnor U18446 (N_18446,N_10077,N_13809);
and U18447 (N_18447,N_11043,N_10610);
xnor U18448 (N_18448,N_13575,N_12215);
nor U18449 (N_18449,N_10896,N_12558);
and U18450 (N_18450,N_13008,N_10476);
nand U18451 (N_18451,N_11756,N_14349);
or U18452 (N_18452,N_14541,N_11448);
nor U18453 (N_18453,N_11608,N_11315);
nand U18454 (N_18454,N_13658,N_11457);
or U18455 (N_18455,N_14350,N_12532);
nand U18456 (N_18456,N_12511,N_13134);
xnor U18457 (N_18457,N_12369,N_10232);
nand U18458 (N_18458,N_11207,N_13787);
nand U18459 (N_18459,N_13674,N_13482);
and U18460 (N_18460,N_14174,N_10642);
and U18461 (N_18461,N_10471,N_10718);
nor U18462 (N_18462,N_11349,N_12776);
xor U18463 (N_18463,N_14668,N_13045);
or U18464 (N_18464,N_14575,N_12719);
or U18465 (N_18465,N_14231,N_14217);
and U18466 (N_18466,N_11881,N_14728);
and U18467 (N_18467,N_13658,N_13535);
nor U18468 (N_18468,N_10036,N_10574);
and U18469 (N_18469,N_11837,N_10668);
and U18470 (N_18470,N_11328,N_10357);
and U18471 (N_18471,N_12880,N_13527);
xnor U18472 (N_18472,N_10202,N_12682);
or U18473 (N_18473,N_13691,N_10227);
or U18474 (N_18474,N_10129,N_14740);
and U18475 (N_18475,N_13892,N_14286);
nor U18476 (N_18476,N_12199,N_11120);
xor U18477 (N_18477,N_14189,N_14676);
nor U18478 (N_18478,N_12081,N_10181);
xor U18479 (N_18479,N_13222,N_11632);
and U18480 (N_18480,N_10510,N_10952);
or U18481 (N_18481,N_11255,N_14875);
and U18482 (N_18482,N_12837,N_14472);
nor U18483 (N_18483,N_14043,N_12607);
nor U18484 (N_18484,N_14897,N_13361);
nand U18485 (N_18485,N_11700,N_10478);
nand U18486 (N_18486,N_12854,N_10881);
xor U18487 (N_18487,N_11049,N_11213);
xor U18488 (N_18488,N_12287,N_12060);
nor U18489 (N_18489,N_10602,N_10991);
or U18490 (N_18490,N_14363,N_13240);
nor U18491 (N_18491,N_12164,N_12293);
and U18492 (N_18492,N_11950,N_13306);
or U18493 (N_18493,N_12772,N_12349);
nand U18494 (N_18494,N_13033,N_13732);
xnor U18495 (N_18495,N_13409,N_13182);
and U18496 (N_18496,N_13216,N_13219);
or U18497 (N_18497,N_13500,N_13196);
and U18498 (N_18498,N_11671,N_11289);
or U18499 (N_18499,N_12130,N_12320);
xor U18500 (N_18500,N_13002,N_14401);
nor U18501 (N_18501,N_11231,N_11959);
nand U18502 (N_18502,N_11672,N_13708);
nand U18503 (N_18503,N_10342,N_12710);
or U18504 (N_18504,N_11594,N_10207);
nor U18505 (N_18505,N_13429,N_10152);
and U18506 (N_18506,N_11680,N_10195);
nand U18507 (N_18507,N_13172,N_14936);
nor U18508 (N_18508,N_12121,N_13836);
nand U18509 (N_18509,N_13659,N_12871);
nand U18510 (N_18510,N_14022,N_12225);
or U18511 (N_18511,N_10445,N_12892);
xor U18512 (N_18512,N_10097,N_13487);
nand U18513 (N_18513,N_13723,N_11771);
xor U18514 (N_18514,N_11087,N_11090);
and U18515 (N_18515,N_10615,N_12363);
xnor U18516 (N_18516,N_11871,N_14012);
xnor U18517 (N_18517,N_14866,N_14562);
and U18518 (N_18518,N_11526,N_10839);
or U18519 (N_18519,N_14045,N_13901);
and U18520 (N_18520,N_11006,N_11183);
and U18521 (N_18521,N_14697,N_10749);
nand U18522 (N_18522,N_10958,N_12284);
or U18523 (N_18523,N_12686,N_12445);
and U18524 (N_18524,N_10752,N_10653);
xnor U18525 (N_18525,N_14214,N_14996);
or U18526 (N_18526,N_14278,N_10495);
and U18527 (N_18527,N_13367,N_10434);
xnor U18528 (N_18528,N_11068,N_14689);
or U18529 (N_18529,N_13122,N_11997);
and U18530 (N_18530,N_13705,N_14552);
or U18531 (N_18531,N_13342,N_10335);
and U18532 (N_18532,N_13566,N_11733);
nor U18533 (N_18533,N_13140,N_11862);
nand U18534 (N_18534,N_12123,N_10492);
nor U18535 (N_18535,N_12054,N_10930);
or U18536 (N_18536,N_11548,N_10475);
nor U18537 (N_18537,N_10457,N_14875);
or U18538 (N_18538,N_13703,N_13845);
or U18539 (N_18539,N_13864,N_10593);
xor U18540 (N_18540,N_12370,N_11841);
nor U18541 (N_18541,N_12386,N_11058);
xnor U18542 (N_18542,N_12974,N_13743);
nor U18543 (N_18543,N_13705,N_11623);
nand U18544 (N_18544,N_13990,N_13350);
nor U18545 (N_18545,N_11565,N_10568);
or U18546 (N_18546,N_12966,N_13374);
nand U18547 (N_18547,N_11496,N_14351);
nor U18548 (N_18548,N_13091,N_14514);
or U18549 (N_18549,N_13939,N_11165);
nand U18550 (N_18550,N_11143,N_10732);
and U18551 (N_18551,N_12490,N_13608);
xor U18552 (N_18552,N_11122,N_13023);
and U18553 (N_18553,N_14079,N_11639);
or U18554 (N_18554,N_12625,N_11223);
and U18555 (N_18555,N_11917,N_10289);
or U18556 (N_18556,N_10655,N_14914);
or U18557 (N_18557,N_13947,N_14155);
xnor U18558 (N_18558,N_13323,N_11869);
and U18559 (N_18559,N_12880,N_11428);
and U18560 (N_18560,N_14600,N_10048);
nor U18561 (N_18561,N_11592,N_10962);
or U18562 (N_18562,N_13205,N_13819);
or U18563 (N_18563,N_13893,N_14597);
or U18564 (N_18564,N_11193,N_12993);
and U18565 (N_18565,N_12874,N_13410);
xor U18566 (N_18566,N_11084,N_14984);
nand U18567 (N_18567,N_10480,N_11349);
xor U18568 (N_18568,N_11658,N_10638);
or U18569 (N_18569,N_10897,N_14756);
nor U18570 (N_18570,N_14935,N_12165);
nor U18571 (N_18571,N_10366,N_14030);
nor U18572 (N_18572,N_13100,N_10460);
and U18573 (N_18573,N_14587,N_10926);
nor U18574 (N_18574,N_13228,N_10290);
or U18575 (N_18575,N_13392,N_14987);
or U18576 (N_18576,N_10236,N_11207);
nor U18577 (N_18577,N_10691,N_10301);
or U18578 (N_18578,N_13352,N_12863);
and U18579 (N_18579,N_13219,N_10978);
xor U18580 (N_18580,N_11172,N_13822);
and U18581 (N_18581,N_12229,N_14421);
or U18582 (N_18582,N_10388,N_10608);
nand U18583 (N_18583,N_10622,N_13648);
nand U18584 (N_18584,N_13559,N_13719);
nor U18585 (N_18585,N_11796,N_13178);
xnor U18586 (N_18586,N_14049,N_11484);
and U18587 (N_18587,N_13653,N_12602);
or U18588 (N_18588,N_10865,N_13551);
xnor U18589 (N_18589,N_10626,N_11573);
and U18590 (N_18590,N_12501,N_10673);
nand U18591 (N_18591,N_10124,N_11102);
nor U18592 (N_18592,N_14744,N_11679);
nor U18593 (N_18593,N_14437,N_12936);
nand U18594 (N_18594,N_12829,N_11953);
and U18595 (N_18595,N_14979,N_10748);
nand U18596 (N_18596,N_12373,N_10687);
nand U18597 (N_18597,N_12785,N_10705);
xnor U18598 (N_18598,N_11944,N_11662);
or U18599 (N_18599,N_10062,N_13744);
nand U18600 (N_18600,N_14573,N_11484);
or U18601 (N_18601,N_13382,N_11064);
nor U18602 (N_18602,N_14000,N_11045);
nor U18603 (N_18603,N_10514,N_10808);
and U18604 (N_18604,N_10412,N_12986);
nor U18605 (N_18605,N_12168,N_10094);
or U18606 (N_18606,N_13316,N_11563);
xor U18607 (N_18607,N_11821,N_14566);
xnor U18608 (N_18608,N_14109,N_10781);
nor U18609 (N_18609,N_11569,N_10641);
nand U18610 (N_18610,N_12766,N_11102);
or U18611 (N_18611,N_14586,N_11454);
and U18612 (N_18612,N_12778,N_14626);
nor U18613 (N_18613,N_13523,N_13794);
nor U18614 (N_18614,N_14371,N_11638);
or U18615 (N_18615,N_14050,N_12727);
xnor U18616 (N_18616,N_11038,N_10094);
xnor U18617 (N_18617,N_13071,N_12884);
or U18618 (N_18618,N_11234,N_10392);
and U18619 (N_18619,N_13919,N_14777);
or U18620 (N_18620,N_11226,N_14624);
nor U18621 (N_18621,N_14183,N_10632);
or U18622 (N_18622,N_12230,N_10834);
or U18623 (N_18623,N_14363,N_14727);
nor U18624 (N_18624,N_12849,N_13075);
xor U18625 (N_18625,N_12130,N_11944);
and U18626 (N_18626,N_14447,N_13532);
or U18627 (N_18627,N_11311,N_11087);
xor U18628 (N_18628,N_11415,N_11989);
nor U18629 (N_18629,N_12892,N_13355);
nor U18630 (N_18630,N_14944,N_10597);
nor U18631 (N_18631,N_11299,N_13684);
and U18632 (N_18632,N_10415,N_14403);
xnor U18633 (N_18633,N_13105,N_13058);
xnor U18634 (N_18634,N_10360,N_13021);
or U18635 (N_18635,N_14693,N_11141);
or U18636 (N_18636,N_12562,N_11295);
nand U18637 (N_18637,N_10061,N_13367);
and U18638 (N_18638,N_13661,N_10741);
and U18639 (N_18639,N_11219,N_11460);
nand U18640 (N_18640,N_14671,N_11273);
or U18641 (N_18641,N_14289,N_13255);
nor U18642 (N_18642,N_14678,N_10796);
or U18643 (N_18643,N_14654,N_10885);
xnor U18644 (N_18644,N_10195,N_14641);
xnor U18645 (N_18645,N_13091,N_14577);
nand U18646 (N_18646,N_11882,N_13251);
nand U18647 (N_18647,N_10952,N_14726);
and U18648 (N_18648,N_12103,N_12975);
nor U18649 (N_18649,N_12837,N_11437);
xor U18650 (N_18650,N_12699,N_14371);
nand U18651 (N_18651,N_12471,N_12574);
nor U18652 (N_18652,N_12280,N_13026);
xnor U18653 (N_18653,N_13622,N_14399);
or U18654 (N_18654,N_12534,N_14630);
xnor U18655 (N_18655,N_12740,N_13471);
and U18656 (N_18656,N_11605,N_13309);
or U18657 (N_18657,N_12028,N_13473);
nand U18658 (N_18658,N_11426,N_11297);
or U18659 (N_18659,N_12840,N_13060);
and U18660 (N_18660,N_11178,N_13155);
or U18661 (N_18661,N_14391,N_13110);
and U18662 (N_18662,N_12792,N_11664);
nand U18663 (N_18663,N_12600,N_14382);
and U18664 (N_18664,N_14986,N_14727);
and U18665 (N_18665,N_10019,N_14391);
or U18666 (N_18666,N_11715,N_13777);
nor U18667 (N_18667,N_14909,N_10404);
nor U18668 (N_18668,N_14079,N_11988);
xor U18669 (N_18669,N_12801,N_13471);
nand U18670 (N_18670,N_14777,N_13671);
and U18671 (N_18671,N_14401,N_14078);
nand U18672 (N_18672,N_14551,N_11720);
nand U18673 (N_18673,N_13165,N_11301);
and U18674 (N_18674,N_11295,N_12097);
and U18675 (N_18675,N_11443,N_12830);
xnor U18676 (N_18676,N_13709,N_11719);
xor U18677 (N_18677,N_10292,N_13813);
or U18678 (N_18678,N_14698,N_14459);
nor U18679 (N_18679,N_11515,N_13906);
nor U18680 (N_18680,N_13267,N_14349);
or U18681 (N_18681,N_10226,N_11338);
nor U18682 (N_18682,N_12903,N_13744);
or U18683 (N_18683,N_11429,N_11736);
nand U18684 (N_18684,N_12064,N_10163);
and U18685 (N_18685,N_14570,N_13991);
and U18686 (N_18686,N_13098,N_10955);
nand U18687 (N_18687,N_14349,N_13363);
nor U18688 (N_18688,N_11179,N_10599);
nand U18689 (N_18689,N_13101,N_11367);
or U18690 (N_18690,N_11104,N_13832);
nand U18691 (N_18691,N_13747,N_10776);
nor U18692 (N_18692,N_10506,N_11793);
and U18693 (N_18693,N_10081,N_12220);
and U18694 (N_18694,N_14279,N_13983);
and U18695 (N_18695,N_14905,N_12730);
nand U18696 (N_18696,N_12826,N_10368);
or U18697 (N_18697,N_14425,N_11295);
nand U18698 (N_18698,N_11382,N_10675);
nor U18699 (N_18699,N_11259,N_10373);
nor U18700 (N_18700,N_11492,N_10398);
xnor U18701 (N_18701,N_13667,N_11334);
and U18702 (N_18702,N_14075,N_13558);
or U18703 (N_18703,N_10522,N_10539);
nand U18704 (N_18704,N_14157,N_13474);
nor U18705 (N_18705,N_13367,N_11063);
xnor U18706 (N_18706,N_14282,N_12087);
and U18707 (N_18707,N_11377,N_12345);
xnor U18708 (N_18708,N_14141,N_14022);
or U18709 (N_18709,N_10330,N_10466);
nor U18710 (N_18710,N_14806,N_10805);
nor U18711 (N_18711,N_14113,N_12603);
xnor U18712 (N_18712,N_10457,N_11010);
nand U18713 (N_18713,N_11751,N_11065);
xnor U18714 (N_18714,N_14827,N_13707);
and U18715 (N_18715,N_10546,N_14066);
or U18716 (N_18716,N_12206,N_14747);
nand U18717 (N_18717,N_13839,N_14657);
and U18718 (N_18718,N_14885,N_12156);
and U18719 (N_18719,N_11948,N_14567);
nand U18720 (N_18720,N_12226,N_11248);
and U18721 (N_18721,N_13303,N_13352);
nor U18722 (N_18722,N_13366,N_12831);
nand U18723 (N_18723,N_10594,N_14164);
or U18724 (N_18724,N_14652,N_10738);
and U18725 (N_18725,N_14538,N_10577);
or U18726 (N_18726,N_12037,N_10987);
xnor U18727 (N_18727,N_12925,N_13830);
nor U18728 (N_18728,N_12105,N_12035);
xnor U18729 (N_18729,N_14544,N_11099);
nor U18730 (N_18730,N_13664,N_14600);
and U18731 (N_18731,N_14074,N_10570);
and U18732 (N_18732,N_13323,N_11522);
or U18733 (N_18733,N_10449,N_14139);
nand U18734 (N_18734,N_14863,N_11077);
or U18735 (N_18735,N_10110,N_13213);
nor U18736 (N_18736,N_14342,N_14686);
nand U18737 (N_18737,N_13671,N_12505);
nor U18738 (N_18738,N_10664,N_13022);
xor U18739 (N_18739,N_10041,N_11768);
nor U18740 (N_18740,N_14675,N_11546);
nor U18741 (N_18741,N_13324,N_12017);
or U18742 (N_18742,N_14979,N_14476);
xor U18743 (N_18743,N_14784,N_13139);
or U18744 (N_18744,N_10745,N_14450);
nor U18745 (N_18745,N_12581,N_10653);
and U18746 (N_18746,N_12114,N_14320);
or U18747 (N_18747,N_12321,N_13018);
nor U18748 (N_18748,N_14271,N_10213);
and U18749 (N_18749,N_13101,N_11536);
and U18750 (N_18750,N_10108,N_11402);
xnor U18751 (N_18751,N_13997,N_14354);
nor U18752 (N_18752,N_13769,N_13299);
nand U18753 (N_18753,N_12413,N_12119);
xnor U18754 (N_18754,N_10810,N_12465);
nor U18755 (N_18755,N_14326,N_10302);
and U18756 (N_18756,N_10875,N_14706);
and U18757 (N_18757,N_14270,N_10417);
xnor U18758 (N_18758,N_12951,N_14547);
nor U18759 (N_18759,N_11837,N_11359);
xnor U18760 (N_18760,N_14419,N_13481);
xnor U18761 (N_18761,N_10075,N_13957);
nor U18762 (N_18762,N_10329,N_14008);
xnor U18763 (N_18763,N_13605,N_10176);
xor U18764 (N_18764,N_10628,N_12798);
nand U18765 (N_18765,N_14518,N_11581);
or U18766 (N_18766,N_13184,N_10440);
nand U18767 (N_18767,N_10289,N_13007);
nand U18768 (N_18768,N_12405,N_14586);
nor U18769 (N_18769,N_11007,N_11551);
xor U18770 (N_18770,N_13334,N_10723);
xor U18771 (N_18771,N_11663,N_10884);
nor U18772 (N_18772,N_14398,N_13905);
nor U18773 (N_18773,N_10719,N_12680);
or U18774 (N_18774,N_11844,N_13501);
or U18775 (N_18775,N_10303,N_10586);
or U18776 (N_18776,N_13679,N_14935);
nor U18777 (N_18777,N_11531,N_14169);
nor U18778 (N_18778,N_10473,N_14735);
and U18779 (N_18779,N_14863,N_12934);
xor U18780 (N_18780,N_12128,N_12133);
and U18781 (N_18781,N_14494,N_10812);
xor U18782 (N_18782,N_13011,N_14008);
and U18783 (N_18783,N_11580,N_13411);
nor U18784 (N_18784,N_13414,N_14519);
nand U18785 (N_18785,N_14593,N_13788);
xnor U18786 (N_18786,N_11868,N_14054);
and U18787 (N_18787,N_12659,N_10063);
nor U18788 (N_18788,N_10939,N_14678);
xor U18789 (N_18789,N_13669,N_10711);
nand U18790 (N_18790,N_13418,N_12565);
nor U18791 (N_18791,N_12202,N_11000);
nand U18792 (N_18792,N_10440,N_12895);
or U18793 (N_18793,N_10925,N_13339);
xor U18794 (N_18794,N_11642,N_12372);
nand U18795 (N_18795,N_13293,N_14675);
or U18796 (N_18796,N_14295,N_14852);
or U18797 (N_18797,N_11640,N_13288);
nor U18798 (N_18798,N_12575,N_10036);
nor U18799 (N_18799,N_12876,N_10306);
nand U18800 (N_18800,N_13706,N_14365);
nor U18801 (N_18801,N_11921,N_10060);
xnor U18802 (N_18802,N_14851,N_13034);
or U18803 (N_18803,N_11220,N_10180);
xnor U18804 (N_18804,N_10047,N_13494);
nor U18805 (N_18805,N_12957,N_10947);
or U18806 (N_18806,N_10423,N_10947);
nor U18807 (N_18807,N_11815,N_13117);
nor U18808 (N_18808,N_13488,N_11685);
xor U18809 (N_18809,N_13882,N_14123);
and U18810 (N_18810,N_13456,N_13186);
xnor U18811 (N_18811,N_13508,N_14579);
or U18812 (N_18812,N_10970,N_11357);
and U18813 (N_18813,N_10459,N_14157);
nand U18814 (N_18814,N_13382,N_10385);
nand U18815 (N_18815,N_13674,N_11855);
nor U18816 (N_18816,N_12135,N_13642);
and U18817 (N_18817,N_11500,N_13320);
nor U18818 (N_18818,N_12055,N_14303);
nor U18819 (N_18819,N_10202,N_13182);
nand U18820 (N_18820,N_14975,N_11474);
nand U18821 (N_18821,N_14700,N_11886);
or U18822 (N_18822,N_13037,N_10624);
xor U18823 (N_18823,N_10518,N_12862);
xor U18824 (N_18824,N_11962,N_14310);
nor U18825 (N_18825,N_12174,N_10164);
xor U18826 (N_18826,N_14488,N_12310);
and U18827 (N_18827,N_10662,N_10292);
xor U18828 (N_18828,N_11572,N_14023);
nor U18829 (N_18829,N_12738,N_14744);
nand U18830 (N_18830,N_10394,N_12480);
nand U18831 (N_18831,N_12941,N_13923);
and U18832 (N_18832,N_14579,N_10493);
xor U18833 (N_18833,N_12448,N_10372);
nor U18834 (N_18834,N_13774,N_13198);
or U18835 (N_18835,N_13945,N_12370);
xnor U18836 (N_18836,N_11683,N_13319);
and U18837 (N_18837,N_10560,N_13279);
nor U18838 (N_18838,N_11915,N_12183);
nand U18839 (N_18839,N_10273,N_13733);
or U18840 (N_18840,N_13076,N_12888);
nand U18841 (N_18841,N_12965,N_10709);
xor U18842 (N_18842,N_13478,N_11938);
nor U18843 (N_18843,N_11057,N_10852);
xnor U18844 (N_18844,N_10033,N_14722);
or U18845 (N_18845,N_13749,N_11318);
or U18846 (N_18846,N_13042,N_14917);
and U18847 (N_18847,N_13404,N_13038);
or U18848 (N_18848,N_10040,N_12987);
nand U18849 (N_18849,N_10988,N_12230);
and U18850 (N_18850,N_14313,N_11319);
nand U18851 (N_18851,N_11153,N_13761);
nand U18852 (N_18852,N_14296,N_13757);
or U18853 (N_18853,N_12424,N_11463);
or U18854 (N_18854,N_11348,N_13873);
and U18855 (N_18855,N_13416,N_13013);
xnor U18856 (N_18856,N_12199,N_12931);
nand U18857 (N_18857,N_13379,N_13171);
xnor U18858 (N_18858,N_12678,N_12200);
nor U18859 (N_18859,N_14553,N_11916);
xnor U18860 (N_18860,N_10023,N_11973);
or U18861 (N_18861,N_10302,N_11452);
nand U18862 (N_18862,N_10864,N_11528);
or U18863 (N_18863,N_14500,N_12161);
nand U18864 (N_18864,N_11105,N_12109);
xnor U18865 (N_18865,N_14947,N_14801);
nor U18866 (N_18866,N_13158,N_10888);
and U18867 (N_18867,N_12994,N_13292);
nor U18868 (N_18868,N_10255,N_11543);
xor U18869 (N_18869,N_12163,N_13497);
or U18870 (N_18870,N_13150,N_11851);
xnor U18871 (N_18871,N_11881,N_10571);
nor U18872 (N_18872,N_13388,N_11060);
nand U18873 (N_18873,N_13187,N_14523);
nand U18874 (N_18874,N_11876,N_14481);
or U18875 (N_18875,N_10498,N_14590);
or U18876 (N_18876,N_11263,N_11052);
and U18877 (N_18877,N_11089,N_13805);
nor U18878 (N_18878,N_11062,N_14333);
and U18879 (N_18879,N_10017,N_11537);
xnor U18880 (N_18880,N_11214,N_13733);
xnor U18881 (N_18881,N_10372,N_10057);
nor U18882 (N_18882,N_10174,N_11630);
nor U18883 (N_18883,N_11592,N_10139);
xnor U18884 (N_18884,N_13787,N_10843);
or U18885 (N_18885,N_14911,N_11799);
or U18886 (N_18886,N_12603,N_11842);
nor U18887 (N_18887,N_14310,N_12533);
nand U18888 (N_18888,N_13874,N_14163);
xnor U18889 (N_18889,N_13076,N_10046);
nand U18890 (N_18890,N_12502,N_14010);
nor U18891 (N_18891,N_12680,N_12982);
and U18892 (N_18892,N_13730,N_11448);
nor U18893 (N_18893,N_10027,N_12285);
or U18894 (N_18894,N_12883,N_10967);
nor U18895 (N_18895,N_10857,N_12960);
xor U18896 (N_18896,N_11925,N_11011);
and U18897 (N_18897,N_14288,N_11136);
xor U18898 (N_18898,N_14463,N_13874);
nand U18899 (N_18899,N_12031,N_14674);
or U18900 (N_18900,N_13670,N_13533);
nand U18901 (N_18901,N_11214,N_14344);
and U18902 (N_18902,N_11212,N_11926);
nand U18903 (N_18903,N_13776,N_14887);
xor U18904 (N_18904,N_12085,N_12199);
or U18905 (N_18905,N_14648,N_14182);
nand U18906 (N_18906,N_12332,N_13010);
or U18907 (N_18907,N_14183,N_13939);
or U18908 (N_18908,N_14132,N_11215);
or U18909 (N_18909,N_13671,N_14438);
nand U18910 (N_18910,N_12765,N_14379);
nor U18911 (N_18911,N_12253,N_14419);
xnor U18912 (N_18912,N_12614,N_14452);
and U18913 (N_18913,N_10002,N_11564);
and U18914 (N_18914,N_12833,N_14511);
or U18915 (N_18915,N_10560,N_11617);
and U18916 (N_18916,N_13874,N_10409);
nor U18917 (N_18917,N_11796,N_13682);
and U18918 (N_18918,N_14836,N_13343);
nor U18919 (N_18919,N_13772,N_12605);
or U18920 (N_18920,N_10819,N_12231);
nor U18921 (N_18921,N_10018,N_13715);
nor U18922 (N_18922,N_11862,N_13111);
xor U18923 (N_18923,N_10538,N_10178);
or U18924 (N_18924,N_12972,N_11676);
or U18925 (N_18925,N_13946,N_11011);
xnor U18926 (N_18926,N_10553,N_11803);
nand U18927 (N_18927,N_10793,N_10742);
or U18928 (N_18928,N_10082,N_14870);
nand U18929 (N_18929,N_14101,N_13973);
nor U18930 (N_18930,N_11825,N_12162);
or U18931 (N_18931,N_13952,N_10415);
or U18932 (N_18932,N_13908,N_14049);
or U18933 (N_18933,N_14749,N_11249);
nor U18934 (N_18934,N_11636,N_10010);
nor U18935 (N_18935,N_13523,N_12495);
nand U18936 (N_18936,N_14099,N_12503);
nand U18937 (N_18937,N_13608,N_12792);
and U18938 (N_18938,N_13839,N_13092);
and U18939 (N_18939,N_12701,N_13708);
and U18940 (N_18940,N_13089,N_14802);
or U18941 (N_18941,N_10333,N_13124);
and U18942 (N_18942,N_11773,N_11761);
and U18943 (N_18943,N_12845,N_13433);
and U18944 (N_18944,N_11712,N_13629);
or U18945 (N_18945,N_10314,N_13360);
nor U18946 (N_18946,N_11601,N_10445);
or U18947 (N_18947,N_11451,N_12163);
nor U18948 (N_18948,N_11024,N_11678);
and U18949 (N_18949,N_14859,N_11765);
and U18950 (N_18950,N_13724,N_12786);
nand U18951 (N_18951,N_10630,N_13215);
xnor U18952 (N_18952,N_13938,N_12383);
xor U18953 (N_18953,N_11379,N_14434);
xor U18954 (N_18954,N_10569,N_14387);
and U18955 (N_18955,N_11995,N_14036);
nand U18956 (N_18956,N_10053,N_10346);
xor U18957 (N_18957,N_11813,N_13331);
and U18958 (N_18958,N_13677,N_13069);
or U18959 (N_18959,N_14600,N_12672);
nand U18960 (N_18960,N_10743,N_13855);
nand U18961 (N_18961,N_12683,N_12138);
nor U18962 (N_18962,N_13060,N_13422);
xnor U18963 (N_18963,N_10019,N_11446);
xnor U18964 (N_18964,N_12593,N_14420);
xor U18965 (N_18965,N_12867,N_10055);
or U18966 (N_18966,N_13016,N_13743);
and U18967 (N_18967,N_11739,N_12856);
nand U18968 (N_18968,N_12876,N_14383);
nand U18969 (N_18969,N_13464,N_13872);
nor U18970 (N_18970,N_13723,N_10109);
and U18971 (N_18971,N_12905,N_12025);
and U18972 (N_18972,N_13155,N_12992);
and U18973 (N_18973,N_11916,N_14873);
or U18974 (N_18974,N_10942,N_11144);
nor U18975 (N_18975,N_10044,N_10557);
and U18976 (N_18976,N_10414,N_10909);
or U18977 (N_18977,N_10062,N_13792);
nor U18978 (N_18978,N_14002,N_12224);
or U18979 (N_18979,N_11766,N_13606);
or U18980 (N_18980,N_12015,N_10682);
xor U18981 (N_18981,N_13979,N_13931);
xnor U18982 (N_18982,N_13808,N_10809);
and U18983 (N_18983,N_11954,N_13554);
nand U18984 (N_18984,N_10801,N_12113);
nor U18985 (N_18985,N_10203,N_11275);
nand U18986 (N_18986,N_14353,N_11595);
or U18987 (N_18987,N_12993,N_13378);
xor U18988 (N_18988,N_12333,N_14619);
and U18989 (N_18989,N_12204,N_12419);
and U18990 (N_18990,N_13366,N_13341);
and U18991 (N_18991,N_14810,N_11389);
or U18992 (N_18992,N_13815,N_13413);
or U18993 (N_18993,N_12629,N_11015);
nand U18994 (N_18994,N_13670,N_11248);
and U18995 (N_18995,N_11469,N_10179);
nand U18996 (N_18996,N_11010,N_10709);
xnor U18997 (N_18997,N_13104,N_11006);
or U18998 (N_18998,N_13686,N_11350);
nand U18999 (N_18999,N_12240,N_12385);
nand U19000 (N_19000,N_11127,N_12468);
nor U19001 (N_19001,N_12093,N_12734);
and U19002 (N_19002,N_11331,N_11761);
nand U19003 (N_19003,N_11371,N_10676);
and U19004 (N_19004,N_10837,N_10172);
nor U19005 (N_19005,N_13583,N_14743);
or U19006 (N_19006,N_10089,N_14255);
nor U19007 (N_19007,N_13947,N_12123);
xor U19008 (N_19008,N_12738,N_11633);
xor U19009 (N_19009,N_11553,N_13704);
nor U19010 (N_19010,N_14753,N_13156);
and U19011 (N_19011,N_12632,N_11471);
nor U19012 (N_19012,N_11323,N_13762);
and U19013 (N_19013,N_10054,N_10155);
and U19014 (N_19014,N_14420,N_12644);
nand U19015 (N_19015,N_14794,N_12807);
or U19016 (N_19016,N_13830,N_12561);
nor U19017 (N_19017,N_13105,N_11086);
nor U19018 (N_19018,N_12745,N_12609);
nor U19019 (N_19019,N_14863,N_12331);
and U19020 (N_19020,N_12346,N_12558);
xnor U19021 (N_19021,N_14042,N_12224);
and U19022 (N_19022,N_14482,N_12258);
xor U19023 (N_19023,N_12878,N_11236);
or U19024 (N_19024,N_10609,N_14093);
or U19025 (N_19025,N_10168,N_14512);
nor U19026 (N_19026,N_13602,N_11316);
xnor U19027 (N_19027,N_14435,N_10737);
nand U19028 (N_19028,N_12977,N_11609);
xnor U19029 (N_19029,N_12531,N_13121);
nand U19030 (N_19030,N_11084,N_11228);
or U19031 (N_19031,N_14848,N_13101);
nor U19032 (N_19032,N_14910,N_13401);
nand U19033 (N_19033,N_13010,N_12139);
nor U19034 (N_19034,N_13437,N_13702);
nand U19035 (N_19035,N_13385,N_12071);
nor U19036 (N_19036,N_14608,N_10330);
and U19037 (N_19037,N_12099,N_12942);
nor U19038 (N_19038,N_10097,N_11048);
nand U19039 (N_19039,N_14556,N_10494);
or U19040 (N_19040,N_13030,N_14948);
nand U19041 (N_19041,N_13040,N_12852);
or U19042 (N_19042,N_12723,N_10761);
and U19043 (N_19043,N_12587,N_12683);
xnor U19044 (N_19044,N_13085,N_11493);
nand U19045 (N_19045,N_11753,N_10260);
and U19046 (N_19046,N_10663,N_12203);
nor U19047 (N_19047,N_14226,N_13947);
xnor U19048 (N_19048,N_13757,N_13608);
xor U19049 (N_19049,N_13565,N_12356);
nor U19050 (N_19050,N_10507,N_13968);
and U19051 (N_19051,N_10245,N_12135);
nor U19052 (N_19052,N_11592,N_13795);
or U19053 (N_19053,N_13926,N_11426);
xor U19054 (N_19054,N_10985,N_14606);
and U19055 (N_19055,N_11216,N_11207);
nand U19056 (N_19056,N_12683,N_14559);
xnor U19057 (N_19057,N_11068,N_14043);
nor U19058 (N_19058,N_12271,N_11517);
and U19059 (N_19059,N_10971,N_13599);
nand U19060 (N_19060,N_13575,N_11609);
xor U19061 (N_19061,N_12305,N_10673);
nor U19062 (N_19062,N_12012,N_13782);
xnor U19063 (N_19063,N_11595,N_14693);
nand U19064 (N_19064,N_11513,N_13623);
nor U19065 (N_19065,N_10933,N_12295);
nor U19066 (N_19066,N_14791,N_10926);
nor U19067 (N_19067,N_10335,N_12266);
and U19068 (N_19068,N_10933,N_14714);
and U19069 (N_19069,N_14944,N_10155);
and U19070 (N_19070,N_13327,N_10066);
or U19071 (N_19071,N_10839,N_14975);
or U19072 (N_19072,N_10633,N_11596);
nand U19073 (N_19073,N_14509,N_14335);
and U19074 (N_19074,N_14825,N_12467);
nand U19075 (N_19075,N_12475,N_13217);
xnor U19076 (N_19076,N_10479,N_10183);
and U19077 (N_19077,N_11441,N_12478);
or U19078 (N_19078,N_14378,N_12180);
nor U19079 (N_19079,N_13839,N_12529);
or U19080 (N_19080,N_12593,N_11373);
xor U19081 (N_19081,N_13288,N_13507);
nor U19082 (N_19082,N_12769,N_12435);
nand U19083 (N_19083,N_10449,N_11028);
and U19084 (N_19084,N_13278,N_14200);
and U19085 (N_19085,N_12560,N_13266);
nand U19086 (N_19086,N_10557,N_13736);
nand U19087 (N_19087,N_11855,N_13133);
nand U19088 (N_19088,N_14929,N_10757);
or U19089 (N_19089,N_12154,N_14147);
or U19090 (N_19090,N_13851,N_13854);
and U19091 (N_19091,N_10827,N_10390);
xor U19092 (N_19092,N_13907,N_10225);
nor U19093 (N_19093,N_11600,N_13077);
or U19094 (N_19094,N_10589,N_14826);
xor U19095 (N_19095,N_13474,N_13087);
xnor U19096 (N_19096,N_12868,N_10221);
xor U19097 (N_19097,N_11939,N_14818);
xor U19098 (N_19098,N_14729,N_14531);
nor U19099 (N_19099,N_12059,N_13208);
and U19100 (N_19100,N_12839,N_10170);
xnor U19101 (N_19101,N_14159,N_14967);
nand U19102 (N_19102,N_11872,N_11565);
nor U19103 (N_19103,N_13537,N_13541);
nand U19104 (N_19104,N_13661,N_10297);
xor U19105 (N_19105,N_14778,N_14663);
and U19106 (N_19106,N_12782,N_14792);
and U19107 (N_19107,N_10892,N_12507);
nand U19108 (N_19108,N_10463,N_10792);
nand U19109 (N_19109,N_11463,N_14718);
and U19110 (N_19110,N_10363,N_11794);
nor U19111 (N_19111,N_10725,N_13561);
nand U19112 (N_19112,N_12834,N_10819);
or U19113 (N_19113,N_10723,N_10997);
xor U19114 (N_19114,N_13903,N_13090);
nand U19115 (N_19115,N_10676,N_13612);
or U19116 (N_19116,N_13404,N_12742);
nand U19117 (N_19117,N_10291,N_12067);
or U19118 (N_19118,N_14243,N_12829);
xnor U19119 (N_19119,N_14546,N_14814);
or U19120 (N_19120,N_12213,N_14023);
or U19121 (N_19121,N_11621,N_13596);
or U19122 (N_19122,N_10178,N_10957);
nand U19123 (N_19123,N_11340,N_12937);
nor U19124 (N_19124,N_11382,N_14850);
or U19125 (N_19125,N_11214,N_12622);
nand U19126 (N_19126,N_14814,N_10911);
nor U19127 (N_19127,N_13945,N_12211);
xnor U19128 (N_19128,N_13564,N_12972);
xor U19129 (N_19129,N_10086,N_14729);
nand U19130 (N_19130,N_12122,N_11281);
nor U19131 (N_19131,N_14481,N_14258);
xor U19132 (N_19132,N_14508,N_12464);
and U19133 (N_19133,N_10649,N_10874);
or U19134 (N_19134,N_13679,N_14308);
xor U19135 (N_19135,N_10035,N_13203);
xor U19136 (N_19136,N_10662,N_12175);
nor U19137 (N_19137,N_14886,N_12737);
nor U19138 (N_19138,N_11481,N_12834);
xor U19139 (N_19139,N_10630,N_11660);
nor U19140 (N_19140,N_10984,N_10681);
xor U19141 (N_19141,N_10576,N_11026);
and U19142 (N_19142,N_12070,N_12804);
nor U19143 (N_19143,N_10910,N_11543);
and U19144 (N_19144,N_14069,N_11270);
nor U19145 (N_19145,N_14183,N_10746);
xnor U19146 (N_19146,N_10241,N_11418);
nor U19147 (N_19147,N_10488,N_11530);
and U19148 (N_19148,N_11765,N_10167);
nand U19149 (N_19149,N_10609,N_14128);
or U19150 (N_19150,N_12907,N_14764);
or U19151 (N_19151,N_10891,N_10440);
nand U19152 (N_19152,N_10105,N_11639);
or U19153 (N_19153,N_13877,N_13278);
xor U19154 (N_19154,N_10956,N_10967);
nand U19155 (N_19155,N_11408,N_11847);
and U19156 (N_19156,N_12504,N_10049);
or U19157 (N_19157,N_13726,N_12155);
nor U19158 (N_19158,N_10828,N_13140);
or U19159 (N_19159,N_14576,N_12498);
nor U19160 (N_19160,N_13776,N_14923);
nor U19161 (N_19161,N_14585,N_14318);
nor U19162 (N_19162,N_10360,N_13162);
and U19163 (N_19163,N_14263,N_11591);
nor U19164 (N_19164,N_11394,N_10973);
and U19165 (N_19165,N_14672,N_11619);
nand U19166 (N_19166,N_11865,N_11597);
nor U19167 (N_19167,N_14341,N_11303);
nor U19168 (N_19168,N_12357,N_14019);
or U19169 (N_19169,N_12044,N_12218);
and U19170 (N_19170,N_13304,N_12037);
or U19171 (N_19171,N_11488,N_12149);
nor U19172 (N_19172,N_12742,N_14697);
xor U19173 (N_19173,N_12957,N_14063);
nand U19174 (N_19174,N_13520,N_10274);
xor U19175 (N_19175,N_13447,N_11288);
nand U19176 (N_19176,N_10749,N_14965);
and U19177 (N_19177,N_10681,N_13911);
xor U19178 (N_19178,N_11837,N_13023);
or U19179 (N_19179,N_11989,N_12859);
nor U19180 (N_19180,N_14517,N_10748);
or U19181 (N_19181,N_10596,N_13765);
nand U19182 (N_19182,N_14712,N_10887);
and U19183 (N_19183,N_11583,N_12843);
xnor U19184 (N_19184,N_11540,N_11032);
nor U19185 (N_19185,N_10268,N_10503);
nand U19186 (N_19186,N_14177,N_13629);
and U19187 (N_19187,N_11345,N_13641);
xor U19188 (N_19188,N_14772,N_12885);
xor U19189 (N_19189,N_14086,N_13105);
and U19190 (N_19190,N_13586,N_13961);
nor U19191 (N_19191,N_13059,N_14306);
and U19192 (N_19192,N_10360,N_13560);
nand U19193 (N_19193,N_11242,N_12519);
xor U19194 (N_19194,N_12501,N_13615);
or U19195 (N_19195,N_12124,N_14642);
xnor U19196 (N_19196,N_10074,N_12222);
xnor U19197 (N_19197,N_13557,N_13299);
or U19198 (N_19198,N_13099,N_13736);
nand U19199 (N_19199,N_13465,N_12795);
nand U19200 (N_19200,N_13541,N_13554);
and U19201 (N_19201,N_11789,N_12577);
xnor U19202 (N_19202,N_10843,N_10524);
nor U19203 (N_19203,N_11108,N_12787);
and U19204 (N_19204,N_14186,N_14072);
or U19205 (N_19205,N_11472,N_12953);
or U19206 (N_19206,N_14730,N_12543);
or U19207 (N_19207,N_13794,N_12996);
and U19208 (N_19208,N_12217,N_10320);
nand U19209 (N_19209,N_12239,N_14138);
or U19210 (N_19210,N_13572,N_12860);
xnor U19211 (N_19211,N_10507,N_12375);
and U19212 (N_19212,N_11789,N_10975);
and U19213 (N_19213,N_10139,N_14506);
or U19214 (N_19214,N_13051,N_10090);
and U19215 (N_19215,N_12056,N_12620);
nor U19216 (N_19216,N_12843,N_14022);
nor U19217 (N_19217,N_13563,N_14411);
nand U19218 (N_19218,N_12775,N_13547);
xnor U19219 (N_19219,N_11912,N_14838);
nand U19220 (N_19220,N_13019,N_12996);
nand U19221 (N_19221,N_12473,N_13833);
nand U19222 (N_19222,N_10903,N_13154);
and U19223 (N_19223,N_14621,N_14504);
and U19224 (N_19224,N_11506,N_11761);
or U19225 (N_19225,N_10985,N_14155);
or U19226 (N_19226,N_14511,N_10885);
or U19227 (N_19227,N_13320,N_11298);
nand U19228 (N_19228,N_14322,N_13227);
nand U19229 (N_19229,N_14068,N_13971);
nand U19230 (N_19230,N_10206,N_12803);
and U19231 (N_19231,N_14028,N_11148);
and U19232 (N_19232,N_11377,N_14781);
xnor U19233 (N_19233,N_10537,N_12415);
and U19234 (N_19234,N_10979,N_14010);
xnor U19235 (N_19235,N_12993,N_11499);
and U19236 (N_19236,N_10643,N_11252);
nand U19237 (N_19237,N_12282,N_10280);
xor U19238 (N_19238,N_13617,N_14865);
nor U19239 (N_19239,N_11787,N_13489);
and U19240 (N_19240,N_13713,N_13190);
xnor U19241 (N_19241,N_11048,N_13039);
nand U19242 (N_19242,N_10405,N_11313);
and U19243 (N_19243,N_13260,N_14149);
xnor U19244 (N_19244,N_11140,N_11327);
nor U19245 (N_19245,N_12758,N_10503);
or U19246 (N_19246,N_13255,N_14219);
nand U19247 (N_19247,N_14794,N_13306);
or U19248 (N_19248,N_13579,N_11310);
nand U19249 (N_19249,N_14271,N_10837);
xor U19250 (N_19250,N_11398,N_11284);
and U19251 (N_19251,N_13715,N_12501);
nor U19252 (N_19252,N_14029,N_13395);
and U19253 (N_19253,N_12927,N_13033);
and U19254 (N_19254,N_10479,N_11443);
or U19255 (N_19255,N_12940,N_11276);
nand U19256 (N_19256,N_12116,N_12971);
xnor U19257 (N_19257,N_10688,N_10634);
nor U19258 (N_19258,N_10424,N_12144);
nor U19259 (N_19259,N_10977,N_13494);
or U19260 (N_19260,N_13259,N_13030);
xnor U19261 (N_19261,N_13762,N_11171);
nor U19262 (N_19262,N_10466,N_13376);
nand U19263 (N_19263,N_11678,N_13990);
nor U19264 (N_19264,N_11498,N_12080);
nand U19265 (N_19265,N_11068,N_14504);
and U19266 (N_19266,N_12115,N_12668);
nand U19267 (N_19267,N_10466,N_11834);
and U19268 (N_19268,N_10059,N_11969);
nand U19269 (N_19269,N_10717,N_14938);
and U19270 (N_19270,N_11100,N_12193);
or U19271 (N_19271,N_10772,N_12220);
nand U19272 (N_19272,N_12295,N_11980);
or U19273 (N_19273,N_10671,N_14622);
or U19274 (N_19274,N_11876,N_14169);
nand U19275 (N_19275,N_10064,N_13805);
nand U19276 (N_19276,N_10491,N_10523);
nand U19277 (N_19277,N_14109,N_12692);
and U19278 (N_19278,N_10117,N_14382);
nor U19279 (N_19279,N_14759,N_10439);
or U19280 (N_19280,N_12100,N_10063);
and U19281 (N_19281,N_10012,N_12004);
or U19282 (N_19282,N_10359,N_13604);
xnor U19283 (N_19283,N_13725,N_13454);
or U19284 (N_19284,N_14299,N_11974);
nor U19285 (N_19285,N_13065,N_14195);
nand U19286 (N_19286,N_14095,N_11800);
xor U19287 (N_19287,N_12362,N_12248);
xor U19288 (N_19288,N_12307,N_12071);
nor U19289 (N_19289,N_11313,N_13433);
nor U19290 (N_19290,N_13023,N_13222);
and U19291 (N_19291,N_11456,N_12528);
nor U19292 (N_19292,N_14582,N_13628);
and U19293 (N_19293,N_11170,N_10864);
xnor U19294 (N_19294,N_10115,N_12554);
xor U19295 (N_19295,N_11906,N_14103);
xor U19296 (N_19296,N_11959,N_12189);
xor U19297 (N_19297,N_14381,N_12000);
xor U19298 (N_19298,N_10346,N_11981);
and U19299 (N_19299,N_13338,N_14792);
and U19300 (N_19300,N_11959,N_10173);
xor U19301 (N_19301,N_11263,N_10555);
nand U19302 (N_19302,N_11217,N_13897);
or U19303 (N_19303,N_14496,N_10967);
nor U19304 (N_19304,N_11346,N_10146);
nor U19305 (N_19305,N_14437,N_10327);
or U19306 (N_19306,N_14402,N_13046);
nand U19307 (N_19307,N_13855,N_11857);
and U19308 (N_19308,N_13793,N_10417);
or U19309 (N_19309,N_12050,N_11810);
xor U19310 (N_19310,N_13112,N_12223);
or U19311 (N_19311,N_10769,N_13124);
nand U19312 (N_19312,N_13737,N_12990);
xnor U19313 (N_19313,N_10279,N_12907);
or U19314 (N_19314,N_11762,N_10963);
xor U19315 (N_19315,N_14936,N_13848);
nor U19316 (N_19316,N_11592,N_13930);
nand U19317 (N_19317,N_11741,N_10053);
or U19318 (N_19318,N_12106,N_13231);
and U19319 (N_19319,N_11210,N_10285);
nor U19320 (N_19320,N_11140,N_13127);
nor U19321 (N_19321,N_10200,N_13797);
or U19322 (N_19322,N_12781,N_10612);
nand U19323 (N_19323,N_14458,N_12047);
or U19324 (N_19324,N_13556,N_12553);
nor U19325 (N_19325,N_10101,N_10692);
or U19326 (N_19326,N_12213,N_14478);
and U19327 (N_19327,N_12939,N_14367);
xnor U19328 (N_19328,N_10862,N_10849);
and U19329 (N_19329,N_11995,N_11099);
nand U19330 (N_19330,N_10658,N_13722);
and U19331 (N_19331,N_12980,N_14922);
and U19332 (N_19332,N_14325,N_14137);
and U19333 (N_19333,N_13426,N_10466);
xnor U19334 (N_19334,N_13144,N_12176);
nor U19335 (N_19335,N_13335,N_13694);
nand U19336 (N_19336,N_11623,N_13395);
xor U19337 (N_19337,N_12785,N_11365);
or U19338 (N_19338,N_10313,N_12202);
nor U19339 (N_19339,N_14534,N_13367);
and U19340 (N_19340,N_10927,N_12134);
xnor U19341 (N_19341,N_10978,N_12056);
nor U19342 (N_19342,N_12182,N_12082);
nor U19343 (N_19343,N_11114,N_10913);
and U19344 (N_19344,N_12496,N_13322);
or U19345 (N_19345,N_14430,N_12742);
or U19346 (N_19346,N_14325,N_14441);
xor U19347 (N_19347,N_12118,N_12427);
nand U19348 (N_19348,N_13368,N_11368);
nand U19349 (N_19349,N_13372,N_13929);
nand U19350 (N_19350,N_14349,N_10245);
or U19351 (N_19351,N_13028,N_11347);
or U19352 (N_19352,N_12125,N_11744);
nand U19353 (N_19353,N_12266,N_10410);
xnor U19354 (N_19354,N_11697,N_11378);
and U19355 (N_19355,N_12143,N_11040);
and U19356 (N_19356,N_10903,N_12263);
nor U19357 (N_19357,N_13682,N_12849);
or U19358 (N_19358,N_10480,N_11122);
or U19359 (N_19359,N_14965,N_11963);
xnor U19360 (N_19360,N_13752,N_11463);
nor U19361 (N_19361,N_10366,N_14143);
or U19362 (N_19362,N_11337,N_11474);
xnor U19363 (N_19363,N_13682,N_10638);
xor U19364 (N_19364,N_14610,N_14256);
nand U19365 (N_19365,N_12593,N_10120);
or U19366 (N_19366,N_10460,N_13684);
nor U19367 (N_19367,N_12497,N_14218);
xor U19368 (N_19368,N_12315,N_13912);
or U19369 (N_19369,N_10811,N_10100);
and U19370 (N_19370,N_10587,N_10473);
xor U19371 (N_19371,N_11906,N_13331);
or U19372 (N_19372,N_14861,N_14740);
xnor U19373 (N_19373,N_11970,N_11148);
nor U19374 (N_19374,N_11121,N_14020);
xor U19375 (N_19375,N_10572,N_11394);
nor U19376 (N_19376,N_13691,N_14644);
or U19377 (N_19377,N_12450,N_14050);
and U19378 (N_19378,N_13183,N_13871);
nand U19379 (N_19379,N_14768,N_10534);
nor U19380 (N_19380,N_12428,N_10402);
and U19381 (N_19381,N_13049,N_10385);
xor U19382 (N_19382,N_14275,N_13378);
and U19383 (N_19383,N_14253,N_14541);
xor U19384 (N_19384,N_14429,N_10928);
nor U19385 (N_19385,N_11924,N_13729);
and U19386 (N_19386,N_11541,N_14575);
xnor U19387 (N_19387,N_10157,N_10513);
nor U19388 (N_19388,N_13236,N_13569);
nor U19389 (N_19389,N_12423,N_10459);
nand U19390 (N_19390,N_12961,N_13749);
and U19391 (N_19391,N_12181,N_12711);
nor U19392 (N_19392,N_14753,N_10631);
nor U19393 (N_19393,N_14771,N_11398);
nand U19394 (N_19394,N_12749,N_12864);
nand U19395 (N_19395,N_11905,N_13973);
nor U19396 (N_19396,N_12246,N_10272);
nor U19397 (N_19397,N_11829,N_14743);
nor U19398 (N_19398,N_13477,N_11103);
nor U19399 (N_19399,N_13798,N_12418);
and U19400 (N_19400,N_10200,N_13413);
nand U19401 (N_19401,N_10076,N_13983);
nor U19402 (N_19402,N_10482,N_12939);
nand U19403 (N_19403,N_13054,N_14006);
and U19404 (N_19404,N_12965,N_12709);
nor U19405 (N_19405,N_12899,N_11048);
and U19406 (N_19406,N_14814,N_10394);
nand U19407 (N_19407,N_10788,N_11848);
or U19408 (N_19408,N_12672,N_12019);
and U19409 (N_19409,N_12187,N_14532);
nor U19410 (N_19410,N_10735,N_11547);
or U19411 (N_19411,N_12180,N_12747);
and U19412 (N_19412,N_11826,N_10312);
xor U19413 (N_19413,N_10500,N_10987);
and U19414 (N_19414,N_14576,N_14035);
or U19415 (N_19415,N_13748,N_13938);
or U19416 (N_19416,N_14184,N_10113);
and U19417 (N_19417,N_14338,N_12342);
or U19418 (N_19418,N_12009,N_10691);
xor U19419 (N_19419,N_13809,N_11328);
and U19420 (N_19420,N_13943,N_10103);
nand U19421 (N_19421,N_10927,N_14066);
nor U19422 (N_19422,N_10271,N_10355);
nor U19423 (N_19423,N_14892,N_13853);
nand U19424 (N_19424,N_14538,N_10131);
xnor U19425 (N_19425,N_12466,N_12992);
and U19426 (N_19426,N_12205,N_13654);
nand U19427 (N_19427,N_11732,N_11120);
nor U19428 (N_19428,N_10360,N_10396);
nor U19429 (N_19429,N_11222,N_10907);
xor U19430 (N_19430,N_11098,N_11186);
nand U19431 (N_19431,N_12477,N_14736);
xnor U19432 (N_19432,N_11172,N_14688);
xor U19433 (N_19433,N_12263,N_12909);
xnor U19434 (N_19434,N_11724,N_14024);
nand U19435 (N_19435,N_11218,N_12729);
nand U19436 (N_19436,N_13549,N_14073);
or U19437 (N_19437,N_13479,N_11715);
nor U19438 (N_19438,N_11833,N_12464);
nand U19439 (N_19439,N_13058,N_13018);
or U19440 (N_19440,N_14181,N_13591);
or U19441 (N_19441,N_10391,N_11901);
and U19442 (N_19442,N_11061,N_13809);
and U19443 (N_19443,N_12050,N_13051);
nor U19444 (N_19444,N_10456,N_10901);
or U19445 (N_19445,N_13907,N_10835);
nand U19446 (N_19446,N_11530,N_13519);
xor U19447 (N_19447,N_12886,N_11962);
nand U19448 (N_19448,N_13875,N_10485);
and U19449 (N_19449,N_14137,N_10952);
or U19450 (N_19450,N_11874,N_11296);
or U19451 (N_19451,N_14837,N_13332);
and U19452 (N_19452,N_14688,N_10675);
xor U19453 (N_19453,N_12680,N_11234);
or U19454 (N_19454,N_12001,N_10750);
nand U19455 (N_19455,N_11701,N_10833);
xor U19456 (N_19456,N_12588,N_14993);
xor U19457 (N_19457,N_12685,N_14872);
and U19458 (N_19458,N_13176,N_14324);
or U19459 (N_19459,N_14703,N_14303);
xor U19460 (N_19460,N_12595,N_14456);
nand U19461 (N_19461,N_10631,N_12467);
and U19462 (N_19462,N_12454,N_13715);
and U19463 (N_19463,N_13790,N_14386);
and U19464 (N_19464,N_10197,N_11452);
and U19465 (N_19465,N_11472,N_14961);
xor U19466 (N_19466,N_14171,N_13843);
or U19467 (N_19467,N_10025,N_11595);
nor U19468 (N_19468,N_10681,N_12266);
nand U19469 (N_19469,N_10850,N_10381);
nand U19470 (N_19470,N_10424,N_12313);
nor U19471 (N_19471,N_14338,N_11445);
or U19472 (N_19472,N_12427,N_10295);
nor U19473 (N_19473,N_12022,N_13794);
and U19474 (N_19474,N_11688,N_12248);
and U19475 (N_19475,N_12527,N_11266);
or U19476 (N_19476,N_14373,N_14195);
xor U19477 (N_19477,N_10207,N_12376);
or U19478 (N_19478,N_10123,N_13026);
or U19479 (N_19479,N_10398,N_13317);
nor U19480 (N_19480,N_11806,N_12494);
or U19481 (N_19481,N_14945,N_10780);
nand U19482 (N_19482,N_10889,N_12425);
xor U19483 (N_19483,N_13985,N_14927);
nand U19484 (N_19484,N_11302,N_11922);
xor U19485 (N_19485,N_10706,N_12421);
xnor U19486 (N_19486,N_13723,N_11581);
nand U19487 (N_19487,N_14662,N_14077);
nand U19488 (N_19488,N_13110,N_11042);
xor U19489 (N_19489,N_12119,N_11086);
xnor U19490 (N_19490,N_12643,N_13636);
nand U19491 (N_19491,N_13771,N_12119);
nand U19492 (N_19492,N_13297,N_13271);
nor U19493 (N_19493,N_12775,N_14571);
nor U19494 (N_19494,N_13963,N_13151);
nand U19495 (N_19495,N_11099,N_14188);
nand U19496 (N_19496,N_14191,N_12090);
nor U19497 (N_19497,N_14494,N_10382);
or U19498 (N_19498,N_13824,N_12563);
xnor U19499 (N_19499,N_13920,N_10624);
xnor U19500 (N_19500,N_14236,N_14787);
nor U19501 (N_19501,N_13177,N_13558);
or U19502 (N_19502,N_10648,N_12726);
nor U19503 (N_19503,N_13487,N_10345);
or U19504 (N_19504,N_13347,N_13521);
or U19505 (N_19505,N_10604,N_10743);
or U19506 (N_19506,N_12667,N_10923);
xor U19507 (N_19507,N_14315,N_11758);
xor U19508 (N_19508,N_13173,N_10441);
xor U19509 (N_19509,N_10487,N_13792);
nand U19510 (N_19510,N_11025,N_14300);
nand U19511 (N_19511,N_14210,N_14162);
xor U19512 (N_19512,N_13612,N_10068);
xnor U19513 (N_19513,N_14603,N_11300);
nor U19514 (N_19514,N_13411,N_12080);
or U19515 (N_19515,N_13624,N_10735);
and U19516 (N_19516,N_10335,N_12185);
or U19517 (N_19517,N_12491,N_12266);
xnor U19518 (N_19518,N_11946,N_11903);
nor U19519 (N_19519,N_11670,N_14804);
and U19520 (N_19520,N_14638,N_12147);
nand U19521 (N_19521,N_14337,N_13369);
or U19522 (N_19522,N_12802,N_11270);
xnor U19523 (N_19523,N_13151,N_12322);
nand U19524 (N_19524,N_14617,N_13189);
or U19525 (N_19525,N_14119,N_11792);
xor U19526 (N_19526,N_12213,N_13061);
nor U19527 (N_19527,N_11591,N_14287);
nor U19528 (N_19528,N_12433,N_10461);
or U19529 (N_19529,N_13523,N_11403);
nor U19530 (N_19530,N_13985,N_14874);
nand U19531 (N_19531,N_11472,N_11643);
and U19532 (N_19532,N_10262,N_10768);
nand U19533 (N_19533,N_10679,N_12477);
xnor U19534 (N_19534,N_11960,N_11948);
and U19535 (N_19535,N_13610,N_13886);
nand U19536 (N_19536,N_12696,N_13981);
or U19537 (N_19537,N_10555,N_12968);
nand U19538 (N_19538,N_12600,N_10829);
nor U19539 (N_19539,N_14608,N_13833);
and U19540 (N_19540,N_10906,N_11794);
xnor U19541 (N_19541,N_14364,N_11400);
nor U19542 (N_19542,N_14773,N_14640);
xnor U19543 (N_19543,N_13512,N_13523);
nor U19544 (N_19544,N_11743,N_14596);
nand U19545 (N_19545,N_10661,N_13322);
and U19546 (N_19546,N_12923,N_14490);
xnor U19547 (N_19547,N_14159,N_10807);
xnor U19548 (N_19548,N_10387,N_11178);
xnor U19549 (N_19549,N_13040,N_12445);
xor U19550 (N_19550,N_11249,N_11140);
or U19551 (N_19551,N_12206,N_10332);
or U19552 (N_19552,N_14598,N_11540);
nand U19553 (N_19553,N_13414,N_14008);
or U19554 (N_19554,N_11474,N_14329);
and U19555 (N_19555,N_10206,N_11212);
nor U19556 (N_19556,N_11660,N_13117);
and U19557 (N_19557,N_12421,N_10962);
and U19558 (N_19558,N_10683,N_13802);
xor U19559 (N_19559,N_13221,N_13255);
nor U19560 (N_19560,N_11268,N_12011);
nand U19561 (N_19561,N_13142,N_14935);
nand U19562 (N_19562,N_14143,N_12205);
xnor U19563 (N_19563,N_12421,N_10132);
and U19564 (N_19564,N_10101,N_10639);
nand U19565 (N_19565,N_13731,N_10766);
nand U19566 (N_19566,N_14048,N_13523);
nand U19567 (N_19567,N_12591,N_12084);
nor U19568 (N_19568,N_11774,N_13735);
nand U19569 (N_19569,N_12649,N_10410);
nand U19570 (N_19570,N_10760,N_12616);
nor U19571 (N_19571,N_12972,N_14295);
or U19572 (N_19572,N_12358,N_11364);
nand U19573 (N_19573,N_10615,N_11158);
nor U19574 (N_19574,N_11361,N_11528);
xor U19575 (N_19575,N_13462,N_13023);
xor U19576 (N_19576,N_10615,N_14339);
nor U19577 (N_19577,N_12190,N_14794);
and U19578 (N_19578,N_14446,N_10724);
nor U19579 (N_19579,N_14745,N_12132);
and U19580 (N_19580,N_14919,N_13439);
nor U19581 (N_19581,N_10259,N_14634);
or U19582 (N_19582,N_10443,N_12364);
or U19583 (N_19583,N_13663,N_11905);
nand U19584 (N_19584,N_14192,N_10441);
nand U19585 (N_19585,N_12292,N_13675);
and U19586 (N_19586,N_14707,N_13218);
nor U19587 (N_19587,N_11914,N_14392);
xor U19588 (N_19588,N_10112,N_11365);
or U19589 (N_19589,N_12067,N_13643);
xor U19590 (N_19590,N_10801,N_14709);
nor U19591 (N_19591,N_14342,N_12824);
nor U19592 (N_19592,N_13508,N_11532);
xor U19593 (N_19593,N_13845,N_11191);
nor U19594 (N_19594,N_14608,N_14200);
nor U19595 (N_19595,N_10777,N_12053);
nand U19596 (N_19596,N_12077,N_14090);
xor U19597 (N_19597,N_10444,N_14987);
or U19598 (N_19598,N_14158,N_12931);
or U19599 (N_19599,N_11540,N_10200);
or U19600 (N_19600,N_11631,N_10157);
or U19601 (N_19601,N_12537,N_10106);
and U19602 (N_19602,N_10084,N_11067);
and U19603 (N_19603,N_13444,N_13792);
nor U19604 (N_19604,N_14824,N_14330);
nand U19605 (N_19605,N_10790,N_13010);
or U19606 (N_19606,N_10527,N_12902);
nor U19607 (N_19607,N_10653,N_11765);
nor U19608 (N_19608,N_13979,N_11108);
xor U19609 (N_19609,N_11180,N_10938);
or U19610 (N_19610,N_12547,N_11353);
nor U19611 (N_19611,N_11957,N_12151);
nand U19612 (N_19612,N_14240,N_14705);
or U19613 (N_19613,N_11778,N_11575);
or U19614 (N_19614,N_10406,N_12414);
xnor U19615 (N_19615,N_13864,N_12700);
nor U19616 (N_19616,N_12532,N_13905);
nor U19617 (N_19617,N_12709,N_11641);
nand U19618 (N_19618,N_13037,N_12920);
and U19619 (N_19619,N_12832,N_10406);
nor U19620 (N_19620,N_14189,N_10266);
nor U19621 (N_19621,N_12192,N_11256);
nand U19622 (N_19622,N_10363,N_14018);
xnor U19623 (N_19623,N_10173,N_13492);
and U19624 (N_19624,N_10233,N_12263);
xor U19625 (N_19625,N_12131,N_13279);
xnor U19626 (N_19626,N_10994,N_10734);
and U19627 (N_19627,N_10835,N_14788);
nand U19628 (N_19628,N_10789,N_11018);
nor U19629 (N_19629,N_10582,N_13712);
or U19630 (N_19630,N_10759,N_13419);
or U19631 (N_19631,N_14449,N_13854);
nor U19632 (N_19632,N_10657,N_12899);
nand U19633 (N_19633,N_14050,N_12603);
xor U19634 (N_19634,N_12356,N_12006);
xnor U19635 (N_19635,N_11064,N_10501);
nand U19636 (N_19636,N_13049,N_11078);
nand U19637 (N_19637,N_10646,N_11471);
or U19638 (N_19638,N_13398,N_13356);
and U19639 (N_19639,N_10835,N_14353);
or U19640 (N_19640,N_14751,N_11050);
nor U19641 (N_19641,N_11491,N_13630);
nand U19642 (N_19642,N_10983,N_14187);
or U19643 (N_19643,N_12480,N_13433);
nor U19644 (N_19644,N_11946,N_12782);
and U19645 (N_19645,N_14286,N_11967);
or U19646 (N_19646,N_13553,N_12918);
xnor U19647 (N_19647,N_10973,N_14566);
and U19648 (N_19648,N_13355,N_12396);
or U19649 (N_19649,N_12803,N_12786);
and U19650 (N_19650,N_13456,N_10121);
nor U19651 (N_19651,N_11476,N_13069);
nor U19652 (N_19652,N_10569,N_11893);
nor U19653 (N_19653,N_13291,N_14768);
and U19654 (N_19654,N_12926,N_13355);
or U19655 (N_19655,N_13907,N_14120);
and U19656 (N_19656,N_14779,N_10861);
nor U19657 (N_19657,N_14821,N_11308);
nand U19658 (N_19658,N_13275,N_12678);
and U19659 (N_19659,N_14551,N_11032);
nor U19660 (N_19660,N_12980,N_13784);
or U19661 (N_19661,N_10440,N_14314);
nor U19662 (N_19662,N_11662,N_13553);
nand U19663 (N_19663,N_12239,N_14341);
nor U19664 (N_19664,N_10885,N_13678);
or U19665 (N_19665,N_13049,N_14792);
nor U19666 (N_19666,N_13370,N_10200);
and U19667 (N_19667,N_10839,N_12554);
and U19668 (N_19668,N_14269,N_10680);
and U19669 (N_19669,N_12883,N_14567);
nand U19670 (N_19670,N_14010,N_14270);
nor U19671 (N_19671,N_12565,N_10400);
xnor U19672 (N_19672,N_14491,N_13265);
and U19673 (N_19673,N_10464,N_10903);
and U19674 (N_19674,N_10226,N_12198);
and U19675 (N_19675,N_14019,N_11290);
and U19676 (N_19676,N_13877,N_10652);
or U19677 (N_19677,N_12314,N_12839);
xor U19678 (N_19678,N_10436,N_11904);
nor U19679 (N_19679,N_11986,N_13553);
nor U19680 (N_19680,N_14234,N_10979);
nor U19681 (N_19681,N_10272,N_10378);
or U19682 (N_19682,N_11110,N_13178);
xor U19683 (N_19683,N_12557,N_12188);
nor U19684 (N_19684,N_11540,N_14684);
nor U19685 (N_19685,N_10708,N_12040);
and U19686 (N_19686,N_14408,N_11850);
and U19687 (N_19687,N_13540,N_14324);
and U19688 (N_19688,N_14582,N_10651);
nor U19689 (N_19689,N_13812,N_12242);
or U19690 (N_19690,N_14253,N_14044);
xnor U19691 (N_19691,N_11436,N_13237);
and U19692 (N_19692,N_11070,N_12346);
nand U19693 (N_19693,N_12677,N_11098);
xnor U19694 (N_19694,N_10726,N_12626);
nand U19695 (N_19695,N_14044,N_10624);
or U19696 (N_19696,N_13379,N_10999);
or U19697 (N_19697,N_14607,N_13993);
or U19698 (N_19698,N_12543,N_10906);
and U19699 (N_19699,N_10455,N_10903);
nor U19700 (N_19700,N_11010,N_10581);
nand U19701 (N_19701,N_10364,N_11095);
or U19702 (N_19702,N_14831,N_12365);
nand U19703 (N_19703,N_13202,N_12103);
and U19704 (N_19704,N_12503,N_10916);
nand U19705 (N_19705,N_14256,N_13877);
nand U19706 (N_19706,N_12155,N_14087);
nor U19707 (N_19707,N_13039,N_13372);
nand U19708 (N_19708,N_14354,N_10609);
or U19709 (N_19709,N_10677,N_10978);
and U19710 (N_19710,N_12002,N_10020);
and U19711 (N_19711,N_12971,N_14269);
and U19712 (N_19712,N_11778,N_11395);
nand U19713 (N_19713,N_12886,N_11893);
nand U19714 (N_19714,N_14601,N_12531);
xor U19715 (N_19715,N_13975,N_14405);
nand U19716 (N_19716,N_13481,N_10469);
nor U19717 (N_19717,N_13896,N_13878);
and U19718 (N_19718,N_11721,N_10469);
nand U19719 (N_19719,N_12089,N_10627);
nand U19720 (N_19720,N_10790,N_11533);
and U19721 (N_19721,N_14286,N_11386);
nand U19722 (N_19722,N_14197,N_11838);
xor U19723 (N_19723,N_10345,N_11139);
xnor U19724 (N_19724,N_11046,N_10997);
xor U19725 (N_19725,N_14116,N_14440);
xnor U19726 (N_19726,N_14402,N_13658);
nand U19727 (N_19727,N_13017,N_11707);
or U19728 (N_19728,N_14117,N_13670);
nand U19729 (N_19729,N_13223,N_11824);
or U19730 (N_19730,N_12140,N_10396);
xnor U19731 (N_19731,N_14024,N_10758);
nor U19732 (N_19732,N_12897,N_10220);
nor U19733 (N_19733,N_12024,N_13426);
and U19734 (N_19734,N_12650,N_11306);
or U19735 (N_19735,N_13619,N_14887);
and U19736 (N_19736,N_10512,N_13643);
xnor U19737 (N_19737,N_11495,N_11024);
nand U19738 (N_19738,N_11279,N_14605);
and U19739 (N_19739,N_14006,N_14193);
nand U19740 (N_19740,N_14649,N_13450);
and U19741 (N_19741,N_10056,N_12098);
or U19742 (N_19742,N_13793,N_14483);
xor U19743 (N_19743,N_12419,N_13660);
nand U19744 (N_19744,N_11213,N_10810);
and U19745 (N_19745,N_12354,N_14554);
and U19746 (N_19746,N_11076,N_12251);
xnor U19747 (N_19747,N_14609,N_14807);
or U19748 (N_19748,N_10099,N_11664);
and U19749 (N_19749,N_14521,N_13555);
and U19750 (N_19750,N_14967,N_12230);
or U19751 (N_19751,N_14982,N_12211);
xnor U19752 (N_19752,N_12953,N_12092);
and U19753 (N_19753,N_12876,N_13151);
nor U19754 (N_19754,N_10800,N_11243);
nand U19755 (N_19755,N_10827,N_10084);
and U19756 (N_19756,N_12870,N_14132);
or U19757 (N_19757,N_10605,N_11032);
nand U19758 (N_19758,N_12911,N_14234);
nor U19759 (N_19759,N_11520,N_14394);
and U19760 (N_19760,N_14819,N_14706);
nand U19761 (N_19761,N_14827,N_11191);
xnor U19762 (N_19762,N_12184,N_10430);
xor U19763 (N_19763,N_14042,N_13271);
xor U19764 (N_19764,N_14729,N_12022);
or U19765 (N_19765,N_13399,N_14899);
nand U19766 (N_19766,N_12644,N_13856);
nand U19767 (N_19767,N_10517,N_13069);
or U19768 (N_19768,N_12788,N_13949);
or U19769 (N_19769,N_11163,N_10478);
nor U19770 (N_19770,N_13385,N_10070);
nor U19771 (N_19771,N_11981,N_14905);
nor U19772 (N_19772,N_11903,N_14537);
nand U19773 (N_19773,N_14945,N_13764);
and U19774 (N_19774,N_10473,N_14822);
nand U19775 (N_19775,N_13688,N_12845);
and U19776 (N_19776,N_11091,N_13939);
nor U19777 (N_19777,N_11590,N_10713);
xor U19778 (N_19778,N_10401,N_11604);
or U19779 (N_19779,N_11444,N_14751);
xnor U19780 (N_19780,N_10822,N_13657);
xor U19781 (N_19781,N_12149,N_12268);
nand U19782 (N_19782,N_11606,N_12825);
xnor U19783 (N_19783,N_14989,N_10394);
xnor U19784 (N_19784,N_13896,N_10538);
xnor U19785 (N_19785,N_13076,N_10808);
nand U19786 (N_19786,N_13030,N_10829);
or U19787 (N_19787,N_14863,N_11517);
or U19788 (N_19788,N_12953,N_14117);
and U19789 (N_19789,N_13845,N_10609);
and U19790 (N_19790,N_11811,N_10260);
nor U19791 (N_19791,N_13977,N_11334);
nand U19792 (N_19792,N_11293,N_11121);
nand U19793 (N_19793,N_14151,N_13718);
xnor U19794 (N_19794,N_10436,N_13607);
and U19795 (N_19795,N_12405,N_13770);
and U19796 (N_19796,N_12145,N_13181);
or U19797 (N_19797,N_10606,N_14825);
xnor U19798 (N_19798,N_14441,N_10728);
nand U19799 (N_19799,N_14564,N_10578);
nand U19800 (N_19800,N_10624,N_12767);
nand U19801 (N_19801,N_14243,N_14170);
and U19802 (N_19802,N_11968,N_14186);
or U19803 (N_19803,N_11753,N_12765);
nand U19804 (N_19804,N_14056,N_14437);
xnor U19805 (N_19805,N_10504,N_13864);
and U19806 (N_19806,N_14028,N_12342);
and U19807 (N_19807,N_11334,N_12852);
nor U19808 (N_19808,N_12748,N_14798);
nor U19809 (N_19809,N_11914,N_13096);
and U19810 (N_19810,N_13903,N_13618);
nor U19811 (N_19811,N_13515,N_14643);
nor U19812 (N_19812,N_11948,N_14883);
xor U19813 (N_19813,N_11529,N_12520);
or U19814 (N_19814,N_13633,N_11910);
nor U19815 (N_19815,N_13511,N_12303);
nand U19816 (N_19816,N_10864,N_12447);
or U19817 (N_19817,N_12659,N_11019);
xnor U19818 (N_19818,N_10931,N_10508);
xnor U19819 (N_19819,N_13152,N_14365);
nand U19820 (N_19820,N_12452,N_13544);
or U19821 (N_19821,N_12615,N_12428);
nand U19822 (N_19822,N_12293,N_13297);
or U19823 (N_19823,N_14689,N_11179);
xor U19824 (N_19824,N_12882,N_10345);
or U19825 (N_19825,N_12627,N_11419);
nor U19826 (N_19826,N_14321,N_13393);
and U19827 (N_19827,N_12596,N_11707);
nand U19828 (N_19828,N_13776,N_12512);
or U19829 (N_19829,N_13809,N_13353);
and U19830 (N_19830,N_12169,N_11273);
and U19831 (N_19831,N_13164,N_11746);
or U19832 (N_19832,N_10898,N_10732);
nor U19833 (N_19833,N_12885,N_13196);
nor U19834 (N_19834,N_13283,N_14243);
nand U19835 (N_19835,N_12561,N_14466);
nor U19836 (N_19836,N_14434,N_14617);
nand U19837 (N_19837,N_13309,N_13672);
or U19838 (N_19838,N_13387,N_10342);
nand U19839 (N_19839,N_10190,N_12253);
and U19840 (N_19840,N_13831,N_13822);
nand U19841 (N_19841,N_14286,N_14453);
and U19842 (N_19842,N_11270,N_11272);
or U19843 (N_19843,N_10038,N_13371);
xnor U19844 (N_19844,N_11406,N_11044);
and U19845 (N_19845,N_14431,N_11817);
nor U19846 (N_19846,N_14352,N_12545);
or U19847 (N_19847,N_14673,N_12380);
and U19848 (N_19848,N_12850,N_10324);
nor U19849 (N_19849,N_10634,N_12003);
nand U19850 (N_19850,N_11271,N_13635);
or U19851 (N_19851,N_11278,N_13311);
and U19852 (N_19852,N_11412,N_12031);
and U19853 (N_19853,N_11557,N_10905);
xnor U19854 (N_19854,N_12272,N_10481);
nand U19855 (N_19855,N_11063,N_13488);
and U19856 (N_19856,N_11331,N_10496);
or U19857 (N_19857,N_14904,N_13222);
xnor U19858 (N_19858,N_13031,N_11131);
nand U19859 (N_19859,N_10859,N_14061);
or U19860 (N_19860,N_14271,N_10793);
nor U19861 (N_19861,N_10608,N_11382);
and U19862 (N_19862,N_13562,N_10050);
nand U19863 (N_19863,N_13676,N_14326);
and U19864 (N_19864,N_11259,N_11170);
and U19865 (N_19865,N_10307,N_14826);
and U19866 (N_19866,N_10035,N_10282);
nor U19867 (N_19867,N_13858,N_13121);
and U19868 (N_19868,N_12122,N_12386);
and U19869 (N_19869,N_12820,N_10312);
or U19870 (N_19870,N_12520,N_14864);
nand U19871 (N_19871,N_11463,N_10030);
and U19872 (N_19872,N_10310,N_10198);
xnor U19873 (N_19873,N_11390,N_14545);
or U19874 (N_19874,N_13188,N_14501);
and U19875 (N_19875,N_12967,N_10272);
nand U19876 (N_19876,N_12740,N_13120);
nand U19877 (N_19877,N_10465,N_11139);
or U19878 (N_19878,N_10441,N_12507);
nand U19879 (N_19879,N_10761,N_10199);
nand U19880 (N_19880,N_10612,N_11754);
xnor U19881 (N_19881,N_13258,N_14096);
xnor U19882 (N_19882,N_13940,N_10888);
xnor U19883 (N_19883,N_14106,N_14564);
and U19884 (N_19884,N_10789,N_13834);
or U19885 (N_19885,N_14964,N_12298);
xor U19886 (N_19886,N_12052,N_11300);
nor U19887 (N_19887,N_12653,N_12134);
or U19888 (N_19888,N_11889,N_11247);
and U19889 (N_19889,N_12072,N_13830);
and U19890 (N_19890,N_14305,N_14093);
nand U19891 (N_19891,N_12626,N_11475);
xnor U19892 (N_19892,N_12570,N_11842);
and U19893 (N_19893,N_11346,N_14086);
xor U19894 (N_19894,N_14807,N_12732);
and U19895 (N_19895,N_11451,N_11154);
or U19896 (N_19896,N_13575,N_11982);
xor U19897 (N_19897,N_10026,N_11260);
or U19898 (N_19898,N_12017,N_12862);
xor U19899 (N_19899,N_11573,N_12960);
nor U19900 (N_19900,N_11914,N_12372);
and U19901 (N_19901,N_13330,N_12845);
xnor U19902 (N_19902,N_12315,N_14002);
and U19903 (N_19903,N_10308,N_10729);
or U19904 (N_19904,N_13666,N_10404);
xor U19905 (N_19905,N_13369,N_12815);
or U19906 (N_19906,N_11572,N_14586);
nor U19907 (N_19907,N_10184,N_14345);
nor U19908 (N_19908,N_14662,N_14528);
xnor U19909 (N_19909,N_12483,N_14163);
nand U19910 (N_19910,N_10097,N_10963);
or U19911 (N_19911,N_13268,N_11722);
and U19912 (N_19912,N_12830,N_14269);
nor U19913 (N_19913,N_10319,N_10905);
or U19914 (N_19914,N_14205,N_10339);
and U19915 (N_19915,N_13453,N_14550);
nand U19916 (N_19916,N_13880,N_12355);
and U19917 (N_19917,N_12760,N_12482);
or U19918 (N_19918,N_10318,N_11337);
nor U19919 (N_19919,N_14828,N_12871);
or U19920 (N_19920,N_13426,N_11362);
nor U19921 (N_19921,N_13181,N_14304);
nor U19922 (N_19922,N_14701,N_11855);
nor U19923 (N_19923,N_10715,N_13496);
nor U19924 (N_19924,N_10769,N_13142);
nand U19925 (N_19925,N_14518,N_13368);
or U19926 (N_19926,N_13648,N_13741);
xnor U19927 (N_19927,N_10662,N_11935);
nand U19928 (N_19928,N_10763,N_10420);
nor U19929 (N_19929,N_10258,N_12400);
xnor U19930 (N_19930,N_10206,N_13103);
nand U19931 (N_19931,N_10956,N_11413);
nand U19932 (N_19932,N_12758,N_12085);
xor U19933 (N_19933,N_12488,N_10374);
and U19934 (N_19934,N_10500,N_10122);
nor U19935 (N_19935,N_10786,N_13944);
nor U19936 (N_19936,N_11344,N_13262);
nor U19937 (N_19937,N_14111,N_11478);
and U19938 (N_19938,N_14849,N_14809);
nor U19939 (N_19939,N_10974,N_11073);
nand U19940 (N_19940,N_11333,N_10961);
xor U19941 (N_19941,N_10062,N_12427);
nor U19942 (N_19942,N_10392,N_14666);
xor U19943 (N_19943,N_13853,N_14521);
and U19944 (N_19944,N_12032,N_13228);
xnor U19945 (N_19945,N_11739,N_14122);
nand U19946 (N_19946,N_13491,N_10074);
nor U19947 (N_19947,N_12615,N_12207);
and U19948 (N_19948,N_12895,N_12167);
or U19949 (N_19949,N_13020,N_11318);
nor U19950 (N_19950,N_10482,N_13074);
nor U19951 (N_19951,N_10013,N_10168);
xor U19952 (N_19952,N_13035,N_10321);
and U19953 (N_19953,N_12007,N_11909);
nand U19954 (N_19954,N_10086,N_12856);
nand U19955 (N_19955,N_10845,N_11965);
nor U19956 (N_19956,N_14034,N_14718);
nand U19957 (N_19957,N_14050,N_14630);
nor U19958 (N_19958,N_10106,N_14181);
and U19959 (N_19959,N_14392,N_12715);
or U19960 (N_19960,N_13595,N_14544);
and U19961 (N_19961,N_14011,N_13078);
and U19962 (N_19962,N_11431,N_13864);
nand U19963 (N_19963,N_12868,N_14919);
or U19964 (N_19964,N_13305,N_13630);
xnor U19965 (N_19965,N_14136,N_10128);
and U19966 (N_19966,N_10475,N_14269);
or U19967 (N_19967,N_11611,N_10548);
or U19968 (N_19968,N_10765,N_12182);
and U19969 (N_19969,N_10552,N_10629);
and U19970 (N_19970,N_13994,N_12700);
nand U19971 (N_19971,N_12178,N_10617);
or U19972 (N_19972,N_10741,N_13384);
nor U19973 (N_19973,N_10742,N_12671);
and U19974 (N_19974,N_13285,N_11695);
nor U19975 (N_19975,N_14257,N_13318);
nor U19976 (N_19976,N_11879,N_11473);
nor U19977 (N_19977,N_12612,N_11609);
nor U19978 (N_19978,N_10117,N_10048);
or U19979 (N_19979,N_14893,N_13517);
and U19980 (N_19980,N_12887,N_11149);
nor U19981 (N_19981,N_12523,N_11133);
nor U19982 (N_19982,N_12491,N_13235);
nand U19983 (N_19983,N_13899,N_14697);
nor U19984 (N_19984,N_10396,N_12306);
and U19985 (N_19985,N_12977,N_10552);
or U19986 (N_19986,N_10910,N_10636);
nand U19987 (N_19987,N_11824,N_12763);
and U19988 (N_19988,N_13114,N_13557);
or U19989 (N_19989,N_14866,N_14250);
nor U19990 (N_19990,N_13368,N_14975);
nand U19991 (N_19991,N_14493,N_13490);
nand U19992 (N_19992,N_12247,N_13628);
and U19993 (N_19993,N_12475,N_14861);
xor U19994 (N_19994,N_11840,N_12971);
nor U19995 (N_19995,N_14521,N_12123);
nand U19996 (N_19996,N_10237,N_10739);
and U19997 (N_19997,N_14874,N_11684);
or U19998 (N_19998,N_11049,N_11065);
nor U19999 (N_19999,N_11110,N_12749);
or UO_0 (O_0,N_15710,N_19617);
and UO_1 (O_1,N_18081,N_19751);
nand UO_2 (O_2,N_16684,N_19685);
nand UO_3 (O_3,N_17027,N_15010);
and UO_4 (O_4,N_16113,N_15014);
nand UO_5 (O_5,N_15229,N_16369);
and UO_6 (O_6,N_19802,N_18139);
xor UO_7 (O_7,N_18187,N_16501);
nor UO_8 (O_8,N_16022,N_16583);
and UO_9 (O_9,N_15082,N_15916);
nor UO_10 (O_10,N_19240,N_17508);
and UO_11 (O_11,N_19303,N_17936);
or UO_12 (O_12,N_18802,N_19811);
or UO_13 (O_13,N_19420,N_19052);
xnor UO_14 (O_14,N_15070,N_18817);
and UO_15 (O_15,N_17011,N_16476);
and UO_16 (O_16,N_16582,N_17776);
xnor UO_17 (O_17,N_16338,N_17827);
and UO_18 (O_18,N_18264,N_16855);
nand UO_19 (O_19,N_15434,N_15911);
nand UO_20 (O_20,N_15749,N_17933);
xor UO_21 (O_21,N_17147,N_19600);
or UO_22 (O_22,N_17145,N_17480);
xnor UO_23 (O_23,N_19196,N_16693);
or UO_24 (O_24,N_18011,N_16445);
xor UO_25 (O_25,N_19020,N_15816);
and UO_26 (O_26,N_16879,N_18166);
xnor UO_27 (O_27,N_15269,N_16614);
xor UO_28 (O_28,N_15473,N_16701);
or UO_29 (O_29,N_16480,N_18303);
and UO_30 (O_30,N_19011,N_15400);
xnor UO_31 (O_31,N_17451,N_16366);
or UO_32 (O_32,N_19306,N_16176);
and UO_33 (O_33,N_18189,N_17959);
or UO_34 (O_34,N_19923,N_16413);
nor UO_35 (O_35,N_17173,N_19559);
nor UO_36 (O_36,N_18798,N_17984);
nor UO_37 (O_37,N_16279,N_15969);
nor UO_38 (O_38,N_19079,N_18651);
xor UO_39 (O_39,N_18128,N_16987);
nand UO_40 (O_40,N_16499,N_15041);
nor UO_41 (O_41,N_15696,N_17526);
or UO_42 (O_42,N_18067,N_17511);
xnor UO_43 (O_43,N_19129,N_16695);
nand UO_44 (O_44,N_18119,N_17719);
xor UO_45 (O_45,N_19267,N_17676);
and UO_46 (O_46,N_17646,N_18679);
and UO_47 (O_47,N_18814,N_18546);
nand UO_48 (O_48,N_15510,N_17167);
xor UO_49 (O_49,N_16159,N_18034);
and UO_50 (O_50,N_17236,N_16929);
nor UO_51 (O_51,N_18244,N_17649);
nand UO_52 (O_52,N_15884,N_17643);
or UO_53 (O_53,N_17603,N_15075);
or UO_54 (O_54,N_18813,N_19987);
and UO_55 (O_55,N_19193,N_17450);
or UO_56 (O_56,N_17928,N_15745);
and UO_57 (O_57,N_18626,N_19487);
and UO_58 (O_58,N_19167,N_18270);
and UO_59 (O_59,N_18513,N_16985);
nor UO_60 (O_60,N_17999,N_18292);
nor UO_61 (O_61,N_16149,N_17578);
nand UO_62 (O_62,N_15479,N_15942);
nor UO_63 (O_63,N_18967,N_15828);
nor UO_64 (O_64,N_15809,N_16566);
xor UO_65 (O_65,N_19309,N_17822);
nor UO_66 (O_66,N_19631,N_18394);
xnor UO_67 (O_67,N_17447,N_17121);
and UO_68 (O_68,N_19755,N_19288);
or UO_69 (O_69,N_16624,N_15088);
nand UO_70 (O_70,N_15414,N_16542);
xor UO_71 (O_71,N_16729,N_16672);
nand UO_72 (O_72,N_16337,N_16331);
nand UO_73 (O_73,N_17668,N_19615);
or UO_74 (O_74,N_17044,N_16291);
or UO_75 (O_75,N_17046,N_17925);
and UO_76 (O_76,N_16535,N_15464);
xor UO_77 (O_77,N_15830,N_16112);
or UO_78 (O_78,N_15917,N_17478);
nand UO_79 (O_79,N_16759,N_16452);
and UO_80 (O_80,N_15735,N_17003);
nand UO_81 (O_81,N_19355,N_15602);
xor UO_82 (O_82,N_19155,N_18017);
or UO_83 (O_83,N_15819,N_18257);
or UO_84 (O_84,N_15701,N_19806);
and UO_85 (O_85,N_15871,N_16037);
nand UO_86 (O_86,N_16004,N_17358);
or UO_87 (O_87,N_16286,N_17782);
nand UO_88 (O_88,N_17886,N_19455);
or UO_89 (O_89,N_16343,N_17378);
nand UO_90 (O_90,N_15035,N_15033);
xnor UO_91 (O_91,N_17878,N_16241);
and UO_92 (O_92,N_17891,N_19710);
nand UO_93 (O_93,N_15939,N_18425);
xnor UO_94 (O_94,N_16088,N_18082);
or UO_95 (O_95,N_17919,N_19488);
or UO_96 (O_96,N_16812,N_17519);
or UO_97 (O_97,N_17188,N_18560);
and UO_98 (O_98,N_15507,N_17852);
and UO_99 (O_99,N_17013,N_19745);
nor UO_100 (O_100,N_17118,N_16714);
nor UO_101 (O_101,N_18952,N_18921);
or UO_102 (O_102,N_19440,N_16899);
or UO_103 (O_103,N_17471,N_15240);
nor UO_104 (O_104,N_18735,N_17061);
nand UO_105 (O_105,N_19367,N_18621);
nor UO_106 (O_106,N_18485,N_16754);
and UO_107 (O_107,N_16458,N_19604);
and UO_108 (O_108,N_15896,N_16340);
or UO_109 (O_109,N_15202,N_17197);
or UO_110 (O_110,N_17665,N_15586);
and UO_111 (O_111,N_17140,N_19870);
nor UO_112 (O_112,N_15505,N_19407);
or UO_113 (O_113,N_19023,N_17353);
or UO_114 (O_114,N_15151,N_19042);
nor UO_115 (O_115,N_16206,N_16243);
and UO_116 (O_116,N_19852,N_16650);
nand UO_117 (O_117,N_19966,N_19032);
and UO_118 (O_118,N_16951,N_17718);
or UO_119 (O_119,N_17360,N_17997);
or UO_120 (O_120,N_17179,N_19706);
nand UO_121 (O_121,N_15419,N_18252);
and UO_122 (O_122,N_19606,N_15245);
nor UO_123 (O_123,N_19709,N_17018);
xnor UO_124 (O_124,N_18795,N_15213);
nand UO_125 (O_125,N_15885,N_18910);
nor UO_126 (O_126,N_17650,N_18765);
xor UO_127 (O_127,N_15108,N_15738);
or UO_128 (O_128,N_18509,N_17418);
nor UO_129 (O_129,N_16454,N_18037);
nand UO_130 (O_130,N_15937,N_17555);
or UO_131 (O_131,N_17338,N_16664);
or UO_132 (O_132,N_18995,N_17271);
nor UO_133 (O_133,N_17726,N_17024);
and UO_134 (O_134,N_17692,N_15962);
nor UO_135 (O_135,N_16975,N_19383);
or UO_136 (O_136,N_19738,N_19195);
xnor UO_137 (O_137,N_19978,N_15998);
xnor UO_138 (O_138,N_17998,N_16101);
nor UO_139 (O_139,N_15160,N_18065);
and UO_140 (O_140,N_18584,N_17007);
nor UO_141 (O_141,N_19117,N_15221);
xor UO_142 (O_142,N_18341,N_15277);
or UO_143 (O_143,N_16405,N_18980);
nor UO_144 (O_144,N_15592,N_15704);
or UO_145 (O_145,N_19910,N_19329);
nor UO_146 (O_146,N_18785,N_16376);
nor UO_147 (O_147,N_15433,N_18520);
and UO_148 (O_148,N_19858,N_19874);
or UO_149 (O_149,N_15188,N_16526);
nor UO_150 (O_150,N_19499,N_15069);
and UO_151 (O_151,N_19323,N_17505);
nand UO_152 (O_152,N_15226,N_17309);
and UO_153 (O_153,N_16442,N_16511);
and UO_154 (O_154,N_16947,N_18276);
nand UO_155 (O_155,N_17085,N_15036);
xnor UO_156 (O_156,N_18871,N_17843);
or UO_157 (O_157,N_17564,N_17513);
nand UO_158 (O_158,N_19156,N_15282);
and UO_159 (O_159,N_19918,N_18984);
xnor UO_160 (O_160,N_18863,N_16562);
xnor UO_161 (O_161,N_15583,N_16744);
and UO_162 (O_162,N_16649,N_16383);
or UO_163 (O_163,N_17272,N_17452);
and UO_164 (O_164,N_16140,N_16568);
or UO_165 (O_165,N_16743,N_17386);
nor UO_166 (O_166,N_19444,N_16519);
xor UO_167 (O_167,N_17401,N_18340);
xor UO_168 (O_168,N_17324,N_19299);
or UO_169 (O_169,N_18183,N_15945);
xor UO_170 (O_170,N_19562,N_16199);
and UO_171 (O_171,N_18171,N_18841);
nor UO_172 (O_172,N_18527,N_17135);
and UO_173 (O_173,N_16127,N_16916);
xor UO_174 (O_174,N_16411,N_19467);
or UO_175 (O_175,N_19392,N_19097);
nand UO_176 (O_176,N_16406,N_18196);
nand UO_177 (O_177,N_16006,N_19312);
nor UO_178 (O_178,N_16441,N_16725);
nand UO_179 (O_179,N_18456,N_15827);
or UO_180 (O_180,N_15593,N_16756);
nor UO_181 (O_181,N_15632,N_17050);
or UO_182 (O_182,N_16742,N_19231);
nand UO_183 (O_183,N_15255,N_19399);
xor UO_184 (O_184,N_17940,N_18610);
nor UO_185 (O_185,N_17503,N_18205);
nand UO_186 (O_186,N_15997,N_15214);
nand UO_187 (O_187,N_19753,N_16021);
and UO_188 (O_188,N_16749,N_17512);
nand UO_189 (O_189,N_16457,N_16153);
nand UO_190 (O_190,N_18322,N_16886);
and UO_191 (O_191,N_16934,N_18231);
nand UO_192 (O_192,N_16385,N_15365);
nand UO_193 (O_193,N_16887,N_15117);
or UO_194 (O_194,N_15989,N_16196);
nand UO_195 (O_195,N_18224,N_15242);
nor UO_196 (O_196,N_17181,N_16118);
or UO_197 (O_197,N_16137,N_18290);
nor UO_198 (O_198,N_15778,N_16048);
nor UO_199 (O_199,N_15781,N_16086);
xor UO_200 (O_200,N_17254,N_15006);
and UO_201 (O_201,N_17711,N_18049);
nand UO_202 (O_202,N_19175,N_18991);
xor UO_203 (O_203,N_15483,N_17784);
xnor UO_204 (O_204,N_17339,N_15284);
and UO_205 (O_205,N_17906,N_17681);
and UO_206 (O_206,N_17337,N_16601);
and UO_207 (O_207,N_19841,N_19327);
nand UO_208 (O_208,N_15297,N_17120);
nor UO_209 (O_209,N_18478,N_17746);
and UO_210 (O_210,N_17388,N_19892);
or UO_211 (O_211,N_19985,N_16166);
xor UO_212 (O_212,N_17908,N_19668);
and UO_213 (O_213,N_19743,N_18226);
nand UO_214 (O_214,N_16261,N_17515);
and UO_215 (O_215,N_18346,N_16786);
or UO_216 (O_216,N_17602,N_15115);
xor UO_217 (O_217,N_16090,N_19242);
and UO_218 (O_218,N_17652,N_18764);
nor UO_219 (O_219,N_15785,N_17045);
nand UO_220 (O_220,N_16438,N_15791);
nand UO_221 (O_221,N_18745,N_19948);
and UO_222 (O_222,N_18315,N_17960);
nand UO_223 (O_223,N_19408,N_17020);
nand UO_224 (O_224,N_19979,N_18946);
and UO_225 (O_225,N_18014,N_18959);
or UO_226 (O_226,N_18783,N_15216);
xor UO_227 (O_227,N_16348,N_19236);
xor UO_228 (O_228,N_15110,N_17365);
xor UO_229 (O_229,N_15148,N_18801);
nor UO_230 (O_230,N_16505,N_18089);
xnor UO_231 (O_231,N_16641,N_15042);
nand UO_232 (O_232,N_15085,N_17675);
and UO_233 (O_233,N_16180,N_19610);
or UO_234 (O_234,N_19908,N_19211);
nor UO_235 (O_235,N_17481,N_18644);
or UO_236 (O_236,N_18739,N_19378);
xnor UO_237 (O_237,N_17553,N_18353);
xnor UO_238 (O_238,N_19699,N_16707);
xor UO_239 (O_239,N_17009,N_15840);
nor UO_240 (O_240,N_19532,N_17761);
nand UO_241 (O_241,N_19316,N_15319);
xnor UO_242 (O_242,N_18488,N_15420);
xor UO_243 (O_243,N_15577,N_19273);
nor UO_244 (O_244,N_18040,N_18678);
nand UO_245 (O_245,N_19104,N_18650);
and UO_246 (O_246,N_15888,N_16081);
nor UO_247 (O_247,N_19254,N_15988);
or UO_248 (O_248,N_16859,N_19914);
xor UO_249 (O_249,N_16470,N_19977);
or UO_250 (O_250,N_17751,N_18668);
and UO_251 (O_251,N_17422,N_17196);
nand UO_252 (O_252,N_15984,N_18230);
xor UO_253 (O_253,N_17441,N_19125);
and UO_254 (O_254,N_17204,N_19655);
nor UO_255 (O_255,N_19425,N_15671);
or UO_256 (O_256,N_15002,N_16804);
nor UO_257 (O_257,N_16528,N_15258);
and UO_258 (O_258,N_19111,N_19774);
and UO_259 (O_259,N_19581,N_15973);
and UO_260 (O_260,N_19109,N_19641);
and UO_261 (O_261,N_18579,N_15086);
nand UO_262 (O_262,N_18329,N_17707);
nor UO_263 (O_263,N_17224,N_18361);
nor UO_264 (O_264,N_18084,N_15266);
or UO_265 (O_265,N_19522,N_15619);
xnor UO_266 (O_266,N_18707,N_18595);
nand UO_267 (O_267,N_17619,N_17715);
nor UO_268 (O_268,N_17752,N_16163);
or UO_269 (O_269,N_19274,N_15542);
nand UO_270 (O_270,N_15679,N_15303);
nand UO_271 (O_271,N_18135,N_16254);
nor UO_272 (O_272,N_15625,N_16753);
and UO_273 (O_273,N_18298,N_16388);
or UO_274 (O_274,N_18255,N_18807);
or UO_275 (O_275,N_17632,N_19215);
and UO_276 (O_276,N_16828,N_19661);
xnor UO_277 (O_277,N_16606,N_18815);
or UO_278 (O_278,N_19570,N_19415);
nor UO_279 (O_279,N_18146,N_18725);
nand UO_280 (O_280,N_19761,N_15180);
nand UO_281 (O_281,N_19374,N_16970);
or UO_282 (O_282,N_16238,N_15311);
nor UO_283 (O_283,N_17357,N_18327);
nor UO_284 (O_284,N_17396,N_18381);
and UO_285 (O_285,N_15415,N_17053);
xnor UO_286 (O_286,N_16067,N_17202);
or UO_287 (O_287,N_15579,N_19915);
nand UO_288 (O_288,N_17740,N_15407);
and UO_289 (O_289,N_18313,N_18943);
nand UO_290 (O_290,N_19742,N_19447);
xnor UO_291 (O_291,N_17443,N_19543);
or UO_292 (O_292,N_17833,N_15802);
and UO_293 (O_293,N_18345,N_15392);
or UO_294 (O_294,N_15126,N_15775);
xor UO_295 (O_295,N_18287,N_15015);
nor UO_296 (O_296,N_15178,N_18080);
nand UO_297 (O_297,N_17763,N_17333);
and UO_298 (O_298,N_18306,N_19103);
xnor UO_299 (O_299,N_19807,N_18951);
xnor UO_300 (O_300,N_15253,N_15243);
xnor UO_301 (O_301,N_17221,N_15683);
xor UO_302 (O_302,N_16773,N_16586);
xnor UO_303 (O_303,N_17484,N_15922);
nor UO_304 (O_304,N_16322,N_16824);
or UO_305 (O_305,N_19095,N_18372);
nor UO_306 (O_306,N_18699,N_18486);
nor UO_307 (O_307,N_16801,N_19851);
xor UO_308 (O_308,N_17657,N_19503);
or UO_309 (O_309,N_15804,N_17395);
or UO_310 (O_310,N_19347,N_18583);
xnor UO_311 (O_311,N_15474,N_17530);
nor UO_312 (O_312,N_17245,N_16817);
xor UO_313 (O_313,N_15780,N_17030);
nor UO_314 (O_314,N_17177,N_19839);
nor UO_315 (O_315,N_17504,N_18142);
nand UO_316 (O_316,N_16724,N_17762);
nor UO_317 (O_317,N_17473,N_15629);
or UO_318 (O_318,N_19217,N_17971);
or UO_319 (O_319,N_17647,N_15661);
xor UO_320 (O_320,N_19625,N_19334);
xor UO_321 (O_321,N_16897,N_17436);
or UO_322 (O_322,N_18923,N_18338);
nor UO_323 (O_323,N_16246,N_17622);
or UO_324 (O_324,N_18222,N_18413);
xnor UO_325 (O_325,N_19465,N_16121);
or UO_326 (O_326,N_17713,N_17556);
and UO_327 (O_327,N_17359,N_18335);
and UO_328 (O_328,N_18444,N_15893);
xor UO_329 (O_329,N_19331,N_18240);
nor UO_330 (O_330,N_15454,N_15448);
xor UO_331 (O_331,N_19076,N_15210);
and UO_332 (O_332,N_19278,N_16215);
xor UO_333 (O_333,N_15318,N_16307);
or UO_334 (O_334,N_15891,N_18009);
and UO_335 (O_335,N_16507,N_16330);
nor UO_336 (O_336,N_19438,N_17062);
nor UO_337 (O_337,N_18866,N_16533);
xor UO_338 (O_338,N_15784,N_18518);
nor UO_339 (O_339,N_17258,N_18574);
nand UO_340 (O_340,N_16293,N_19897);
nand UO_341 (O_341,N_19946,N_16625);
nand UO_342 (O_342,N_17788,N_16155);
nor UO_343 (O_343,N_15990,N_19726);
or UO_344 (O_344,N_17539,N_15307);
or UO_345 (O_345,N_16545,N_19065);
or UO_346 (O_346,N_19439,N_17280);
nor UO_347 (O_347,N_18956,N_18855);
nor UO_348 (O_348,N_18818,N_17616);
xor UO_349 (O_349,N_15825,N_15799);
and UO_350 (O_350,N_17077,N_15516);
nor UO_351 (O_351,N_18682,N_19257);
or UO_352 (O_352,N_19000,N_18124);
xnor UO_353 (O_353,N_16135,N_16613);
nor UO_354 (O_354,N_16755,N_16425);
nor UO_355 (O_355,N_19994,N_16837);
xnor UO_356 (O_356,N_19101,N_17694);
nand UO_357 (O_357,N_16058,N_19171);
and UO_358 (O_358,N_19575,N_18487);
or UO_359 (O_359,N_18368,N_19492);
nor UO_360 (O_360,N_15107,N_17461);
nand UO_361 (O_361,N_16997,N_18021);
xnor UO_362 (O_362,N_17310,N_16680);
or UO_363 (O_363,N_17318,N_15196);
and UO_364 (O_364,N_15543,N_18777);
nand UO_365 (O_365,N_16678,N_18157);
and UO_366 (O_366,N_19703,N_17305);
or UO_367 (O_367,N_15821,N_15480);
xnor UO_368 (O_368,N_15983,N_19805);
xor UO_369 (O_369,N_15912,N_19293);
and UO_370 (O_370,N_16265,N_17114);
and UO_371 (O_371,N_15718,N_18551);
xnor UO_372 (O_372,N_18378,N_16979);
xor UO_373 (O_373,N_16077,N_18191);
and UO_374 (O_374,N_16621,N_19632);
and UO_375 (O_375,N_18968,N_18778);
xor UO_376 (O_376,N_18896,N_19188);
nor UO_377 (O_377,N_15100,N_15466);
and UO_378 (O_378,N_18402,N_15947);
nor UO_379 (O_379,N_18672,N_18105);
and UO_380 (O_380,N_16633,N_15789);
and UO_381 (O_381,N_15571,N_17232);
xnor UO_382 (O_382,N_19014,N_17312);
nor UO_383 (O_383,N_17157,N_18359);
xnor UO_384 (O_384,N_19018,N_18319);
nor UO_385 (O_385,N_17950,N_18704);
nand UO_386 (O_386,N_15032,N_15688);
and UO_387 (O_387,N_18248,N_19132);
nor UO_388 (O_388,N_17986,N_18688);
nor UO_389 (O_389,N_17001,N_17308);
nor UO_390 (O_390,N_16219,N_17262);
nor UO_391 (O_391,N_17385,N_16675);
xnor UO_392 (O_392,N_16658,N_19370);
or UO_393 (O_393,N_18627,N_17685);
or UO_394 (O_394,N_17845,N_18429);
xor UO_395 (O_395,N_19635,N_15299);
xor UO_396 (O_396,N_16025,N_18380);
nor UO_397 (O_397,N_19343,N_17509);
or UO_398 (O_398,N_19265,N_16648);
xnor UO_399 (O_399,N_18806,N_18772);
nor UO_400 (O_400,N_17489,N_17809);
and UO_401 (O_401,N_15605,N_19158);
nand UO_402 (O_402,N_17335,N_17522);
and UO_403 (O_403,N_16467,N_15451);
or UO_404 (O_404,N_16436,N_15295);
or UO_405 (O_405,N_17220,N_18902);
and UO_406 (O_406,N_18919,N_15664);
nor UO_407 (O_407,N_16989,N_16604);
xor UO_408 (O_408,N_17412,N_15271);
nor UO_409 (O_409,N_15757,N_18751);
nand UO_410 (O_410,N_18177,N_16292);
xnor UO_411 (O_411,N_15022,N_15192);
or UO_412 (O_412,N_15157,N_18388);
nor UO_413 (O_413,N_19813,N_16204);
or UO_414 (O_414,N_19473,N_16775);
xor UO_415 (O_415,N_15410,N_16356);
nor UO_416 (O_416,N_18883,N_17356);
nor UO_417 (O_417,N_17648,N_19785);
or UO_418 (O_418,N_18730,N_19022);
and UO_419 (O_419,N_18092,N_16561);
and UO_420 (O_420,N_15967,N_17783);
or UO_421 (O_421,N_19759,N_16637);
or UO_422 (O_422,N_16083,N_17945);
nand UO_423 (O_423,N_17417,N_17824);
nor UO_424 (O_424,N_15074,N_16799);
and UO_425 (O_425,N_19024,N_16095);
and UO_426 (O_426,N_17880,N_15000);
nand UO_427 (O_427,N_18630,N_15076);
and UO_428 (O_428,N_19768,N_19667);
and UO_429 (O_429,N_16638,N_17642);
nand UO_430 (O_430,N_18199,N_16008);
xnor UO_431 (O_431,N_19563,N_16785);
and UO_432 (O_432,N_16209,N_19163);
xnor UO_433 (O_433,N_18983,N_16080);
or UO_434 (O_434,N_19074,N_16765);
nand UO_435 (O_435,N_15404,N_19174);
or UO_436 (O_436,N_19388,N_16418);
nand UO_437 (O_437,N_15970,N_18022);
nand UO_438 (O_438,N_17801,N_18097);
and UO_439 (O_439,N_17311,N_16298);
xor UO_440 (O_440,N_19162,N_16666);
nand UO_441 (O_441,N_19249,N_15156);
nand UO_442 (O_442,N_19234,N_16409);
nor UO_443 (O_443,N_16214,N_19494);
nand UO_444 (O_444,N_18590,N_18998);
and UO_445 (O_445,N_19855,N_19300);
and UO_446 (O_446,N_16757,N_16966);
xor UO_447 (O_447,N_19422,N_16056);
or UO_448 (O_448,N_18779,N_16160);
nand UO_449 (O_449,N_17319,N_15720);
nand UO_450 (O_450,N_16361,N_19790);
or UO_451 (O_451,N_15397,N_17545);
and UO_452 (O_452,N_16740,N_18834);
xnor UO_453 (O_453,N_18517,N_17689);
or UO_454 (O_454,N_15247,N_16818);
xnor UO_455 (O_455,N_18305,N_18564);
xnor UO_456 (O_456,N_15875,N_18571);
and UO_457 (O_457,N_17372,N_18843);
nor UO_458 (O_458,N_16456,N_15061);
nand UO_459 (O_459,N_15955,N_15128);
nand UO_460 (O_460,N_17592,N_16651);
nor UO_461 (O_461,N_16731,N_19148);
nor UO_462 (O_462,N_16096,N_17837);
and UO_463 (O_463,N_15012,N_19044);
nor UO_464 (O_464,N_16807,N_19474);
xor UO_465 (O_465,N_18819,N_19723);
and UO_466 (O_466,N_19212,N_18709);
nor UO_467 (O_467,N_19143,N_19634);
nor UO_468 (O_468,N_18749,N_16882);
nor UO_469 (O_469,N_16866,N_16794);
nand UO_470 (O_470,N_18864,N_19800);
or UO_471 (O_471,N_18603,N_15325);
or UO_472 (O_472,N_16884,N_15315);
or UO_473 (O_473,N_19630,N_17819);
or UO_474 (O_474,N_17369,N_16247);
xnor UO_475 (O_475,N_15452,N_16244);
or UO_476 (O_476,N_16381,N_16446);
or UO_477 (O_477,N_15626,N_18304);
xor UO_478 (O_478,N_15852,N_16889);
xnor UO_479 (O_479,N_19033,N_15232);
or UO_480 (O_480,N_15470,N_17091);
nand UO_481 (O_481,N_15693,N_17695);
or UO_482 (O_482,N_18179,N_18963);
and UO_483 (O_483,N_18193,N_18930);
nand UO_484 (O_484,N_18442,N_16796);
xnor UO_485 (O_485,N_15486,N_19502);
nor UO_486 (O_486,N_16784,N_18985);
xnor UO_487 (O_487,N_18198,N_16850);
nand UO_488 (O_488,N_15901,N_19861);
xor UO_489 (O_489,N_15235,N_18903);
nor UO_490 (O_490,N_15152,N_19721);
nor UO_491 (O_491,N_16888,N_16375);
and UO_492 (O_492,N_18625,N_17735);
nor UO_493 (O_493,N_15844,N_16401);
and UO_494 (O_494,N_15238,N_15961);
nor UO_495 (O_495,N_16833,N_15575);
nand UO_496 (O_496,N_16974,N_19192);
and UO_497 (O_497,N_16208,N_16061);
xnor UO_498 (O_498,N_19886,N_17777);
nor UO_499 (O_499,N_18750,N_19172);
xnor UO_500 (O_500,N_17332,N_18992);
nand UO_501 (O_501,N_19798,N_19989);
xnor UO_502 (O_502,N_19823,N_15034);
nand UO_503 (O_503,N_15659,N_17292);
and UO_504 (O_504,N_15106,N_17209);
and UO_505 (O_505,N_16657,N_15905);
and UO_506 (O_506,N_16876,N_16468);
nor UO_507 (O_507,N_17610,N_19657);
or UO_508 (O_508,N_17206,N_19816);
and UO_509 (O_509,N_18636,N_16602);
nor UO_510 (O_510,N_16363,N_18892);
nor UO_511 (O_511,N_15143,N_15546);
xor UO_512 (O_512,N_17573,N_16721);
nor UO_513 (O_513,N_17529,N_18858);
nand UO_514 (O_514,N_17798,N_17769);
xnor UO_515 (O_515,N_15662,N_17191);
nand UO_516 (O_516,N_16977,N_18835);
or UO_517 (O_517,N_17421,N_19070);
or UO_518 (O_518,N_17387,N_17823);
nand UO_519 (O_519,N_16047,N_15021);
nand UO_520 (O_520,N_18587,N_16632);
or UO_521 (O_521,N_19339,N_17818);
nor UO_522 (O_522,N_18182,N_17458);
nor UO_523 (O_523,N_19366,N_18743);
nor UO_524 (O_524,N_17551,N_19958);
or UO_525 (O_525,N_15494,N_15599);
nand UO_526 (O_526,N_15829,N_18950);
xor UO_527 (O_527,N_15264,N_16120);
xor UO_528 (O_528,N_15123,N_19894);
nand UO_529 (O_529,N_18033,N_16301);
nand UO_530 (O_530,N_18717,N_18647);
nand UO_531 (O_531,N_16747,N_17313);
xnor UO_532 (O_532,N_15324,N_19119);
xnor UO_533 (O_533,N_18877,N_16549);
nor UO_534 (O_534,N_17037,N_15567);
nand UO_535 (O_535,N_19490,N_19963);
nor UO_536 (O_536,N_19666,N_15281);
xnor UO_537 (O_537,N_18804,N_19950);
xor UO_538 (O_538,N_17170,N_16892);
xor UO_539 (O_539,N_15949,N_18406);
or UO_540 (O_540,N_15093,N_16865);
or UO_541 (O_541,N_16350,N_16252);
and UO_542 (O_542,N_18047,N_19066);
nand UO_543 (O_543,N_16688,N_18170);
nor UO_544 (O_544,N_16847,N_15341);
nand UO_545 (O_545,N_15564,N_15615);
or UO_546 (O_546,N_16642,N_16465);
nand UO_547 (O_547,N_16768,N_17717);
and UO_548 (O_548,N_16921,N_17344);
or UO_549 (O_549,N_19670,N_15956);
nand UO_550 (O_550,N_18716,N_19324);
nand UO_551 (O_551,N_19636,N_15294);
or UO_552 (O_552,N_19810,N_19648);
and UO_553 (O_553,N_17724,N_18667);
nand UO_554 (O_554,N_16548,N_16198);
xor UO_555 (O_555,N_19788,N_19660);
xor UO_556 (O_556,N_16779,N_19508);
nor UO_557 (O_557,N_18161,N_19483);
nor UO_558 (O_558,N_19954,N_16798);
and UO_559 (O_559,N_19009,N_19133);
nand UO_560 (O_560,N_18853,N_15897);
or UO_561 (O_561,N_17065,N_18206);
and UO_562 (O_562,N_19593,N_18087);
nand UO_563 (O_563,N_19762,N_16100);
nand UO_564 (O_564,N_16555,N_17446);
nor UO_565 (O_565,N_19973,N_18781);
nand UO_566 (O_566,N_17099,N_19206);
or UO_567 (O_567,N_19582,N_17576);
xnor UO_568 (O_568,N_18070,N_17340);
or UO_569 (O_569,N_15389,N_19523);
or UO_570 (O_570,N_18803,N_15976);
nand UO_571 (O_571,N_19498,N_17423);
xor UO_572 (O_572,N_19772,N_15886);
nor UO_573 (O_573,N_15184,N_17587);
nand UO_574 (O_574,N_19822,N_18615);
nor UO_575 (O_575,N_17314,N_15608);
nand UO_576 (O_576,N_17403,N_17918);
or UO_577 (O_577,N_17976,N_17259);
nand UO_578 (O_578,N_16332,N_19199);
nand UO_579 (O_579,N_16060,N_17031);
nor UO_580 (O_580,N_19345,N_15487);
nand UO_581 (O_581,N_19750,N_16028);
or UO_582 (O_582,N_17049,N_17122);
or UO_583 (O_583,N_18862,N_18144);
nor UO_584 (O_584,N_15136,N_19385);
or UO_585 (O_585,N_17470,N_15648);
and UO_586 (O_586,N_18234,N_19041);
nand UO_587 (O_587,N_16339,N_17190);
or UO_588 (O_588,N_17688,N_18575);
and UO_589 (O_589,N_15119,N_19019);
or UO_590 (O_590,N_19786,N_15761);
and UO_591 (O_591,N_16864,N_16584);
or UO_592 (O_592,N_16314,N_16302);
or UO_593 (O_593,N_18484,N_17912);
and UO_594 (O_594,N_19400,N_19244);
nor UO_595 (O_595,N_16032,N_17656);
nand UO_596 (O_596,N_19725,N_18763);
xnor UO_597 (O_597,N_16427,N_18282);
nand UO_598 (O_598,N_17770,N_16591);
xnor UO_599 (O_599,N_16769,N_16861);
and UO_600 (O_600,N_17267,N_19882);
xnor UO_601 (O_601,N_16952,N_17463);
or UO_602 (O_602,N_17345,N_19951);
nand UO_603 (O_603,N_19746,N_15934);
nor UO_604 (O_604,N_19854,N_17698);
and UO_605 (O_605,N_16956,N_17705);
or UO_606 (O_606,N_17596,N_16092);
xor UO_607 (O_607,N_16187,N_16079);
or UO_608 (O_608,N_19732,N_15124);
nor UO_609 (O_609,N_15173,N_19221);
and UO_610 (O_610,N_17017,N_16231);
or UO_611 (O_611,N_17864,N_17542);
nor UO_612 (O_612,N_15142,N_16108);
nand UO_613 (O_613,N_15368,N_15455);
nor UO_614 (O_614,N_18140,N_19459);
nand UO_615 (O_615,N_17832,N_16829);
or UO_616 (O_616,N_15737,N_16644);
or UO_617 (O_617,N_18917,N_16116);
nand UO_618 (O_618,N_19237,N_17103);
or UO_619 (O_619,N_17620,N_18354);
xnor UO_620 (O_620,N_18324,N_19921);
and UO_621 (O_621,N_16394,N_16421);
and UO_622 (O_622,N_18759,N_15438);
and UO_623 (O_623,N_17281,N_18606);
and UO_624 (O_624,N_15861,N_16821);
nand UO_625 (O_625,N_18570,N_15332);
nor UO_626 (O_626,N_17948,N_17393);
nor UO_627 (O_627,N_19929,N_18639);
and UO_628 (O_628,N_15944,N_17426);
xor UO_629 (O_629,N_18540,N_17606);
nor UO_630 (O_630,N_18929,N_16111);
nor UO_631 (O_631,N_19749,N_18366);
or UO_632 (O_632,N_18659,N_17854);
nand UO_633 (O_633,N_15587,N_17400);
nand UO_634 (O_634,N_15375,N_15753);
nor UO_635 (O_635,N_19296,N_16854);
or UO_636 (O_636,N_15026,N_16210);
nand UO_637 (O_637,N_18993,N_19509);
nor UO_638 (O_638,N_18350,N_15766);
nand UO_639 (O_639,N_18620,N_15306);
nor UO_640 (O_640,N_16697,N_15639);
and UO_641 (O_641,N_17149,N_19353);
nor UO_642 (O_642,N_19281,N_16251);
nand UO_643 (O_643,N_19614,N_16572);
nor UO_644 (O_644,N_18357,N_15752);
nand UO_645 (O_645,N_18057,N_19341);
and UO_646 (O_646,N_17138,N_15146);
xor UO_647 (O_647,N_17856,N_18130);
xnor UO_648 (O_648,N_15550,N_18094);
or UO_649 (O_649,N_18673,N_17466);
nand UO_650 (O_650,N_17584,N_15951);
xnor UO_651 (O_651,N_17494,N_18100);
nand UO_652 (O_652,N_16915,N_17525);
nand UO_653 (O_653,N_17828,N_17315);
or UO_654 (O_654,N_15687,N_16577);
xnor UO_655 (O_655,N_18348,N_16391);
or UO_656 (O_656,N_17535,N_18577);
nor UO_657 (O_657,N_18794,N_16239);
and UO_658 (O_658,N_17733,N_17076);
nand UO_659 (O_659,N_16663,N_16700);
nor UO_660 (O_660,N_18782,N_15660);
nor UO_661 (O_661,N_18856,N_19818);
nand UO_662 (O_662,N_17263,N_19866);
or UO_663 (O_663,N_18960,N_18294);
or UO_664 (O_664,N_19491,N_19332);
or UO_665 (O_665,N_17364,N_19776);
and UO_666 (O_666,N_16453,N_18529);
xor UO_667 (O_667,N_15529,N_18916);
or UO_668 (O_668,N_17483,N_19702);
xnor UO_669 (O_669,N_15628,N_15925);
xnor UO_670 (O_670,N_19071,N_19814);
and UO_671 (O_671,N_17902,N_19917);
nor UO_672 (O_672,N_15528,N_19016);
xor UO_673 (O_673,N_17618,N_18432);
nand UO_674 (O_674,N_15812,N_17589);
or UO_675 (O_675,N_15059,N_16287);
xnor UO_676 (O_676,N_16727,N_15851);
nor UO_677 (O_677,N_16217,N_19737);
nand UO_678 (O_678,N_17704,N_18336);
or UO_679 (O_679,N_18133,N_18965);
nor UO_680 (O_680,N_16455,N_17303);
nor UO_681 (O_681,N_19149,N_17496);
nor UO_682 (O_682,N_17904,N_15726);
or UO_683 (O_683,N_16509,N_15762);
xor UO_684 (O_684,N_15337,N_18543);
xor UO_685 (O_685,N_18440,N_17939);
xnor UO_686 (O_686,N_15918,N_18131);
nor UO_687 (O_687,N_18349,N_18530);
nand UO_688 (O_688,N_19120,N_16440);
or UO_689 (O_689,N_15674,N_16321);
nand UO_690 (O_690,N_19927,N_19185);
nand UO_691 (O_691,N_15904,N_15388);
or UO_692 (O_692,N_16546,N_15794);
nor UO_693 (O_693,N_17992,N_15963);
nand UO_694 (O_694,N_16563,N_19243);
and UO_695 (O_695,N_18347,N_15073);
nand UO_696 (O_696,N_19466,N_19724);
nand UO_697 (O_697,N_15159,N_17322);
nand UO_698 (O_698,N_17175,N_19679);
nor UO_699 (O_699,N_15333,N_15199);
or UO_700 (O_700,N_17270,N_17568);
and UO_701 (O_701,N_19787,N_17932);
nor UO_702 (O_702,N_16203,N_16573);
nand UO_703 (O_703,N_16143,N_18729);
and UO_704 (O_704,N_18611,N_17035);
nand UO_705 (O_705,N_17946,N_15728);
nor UO_706 (O_706,N_17217,N_17241);
or UO_707 (O_707,N_18568,N_19624);
nand UO_708 (O_708,N_17516,N_16610);
nor UO_709 (O_709,N_15083,N_15902);
and UO_710 (O_710,N_19521,N_18150);
or UO_711 (O_711,N_19134,N_19205);
xor UO_712 (O_712,N_19409,N_17575);
nor UO_713 (O_713,N_15072,N_16868);
or UO_714 (O_714,N_16525,N_15362);
nor UO_715 (O_715,N_17638,N_18296);
nor UO_716 (O_716,N_16983,N_16129);
nand UO_717 (O_717,N_16462,N_18439);
nor UO_718 (O_718,N_15097,N_19611);
xnor UO_719 (O_719,N_19107,N_19552);
and UO_720 (O_720,N_17462,N_15598);
nor UO_721 (O_721,N_15658,N_17178);
or UO_722 (O_722,N_18427,N_19294);
xnor UO_723 (O_723,N_19775,N_19556);
or UO_724 (O_724,N_16071,N_16170);
and UO_725 (O_725,N_16726,N_17894);
and UO_726 (O_726,N_18412,N_15363);
nor UO_727 (O_727,N_17370,N_18711);
nand UO_728 (O_728,N_15624,N_16598);
nand UO_729 (O_729,N_15894,N_18790);
xor UO_730 (O_730,N_16539,N_15430);
nor UO_731 (O_731,N_15800,N_19609);
or UO_732 (O_732,N_15244,N_17794);
nand UO_733 (O_733,N_18403,N_17449);
or UO_734 (O_734,N_19393,N_19313);
and UO_735 (O_735,N_19933,N_17821);
or UO_736 (O_736,N_15037,N_17243);
nor UO_737 (O_737,N_15876,N_15469);
or UO_738 (O_738,N_15447,N_19390);
nand UO_739 (O_739,N_19857,N_18163);
and UO_740 (O_740,N_18538,N_18370);
nor UO_741 (O_741,N_17947,N_19803);
nor UO_742 (O_742,N_16805,N_15964);
nand UO_743 (O_743,N_16288,N_15864);
nor UO_744 (O_744,N_15919,N_15521);
xnor UO_745 (O_745,N_17022,N_19029);
or UO_746 (O_746,N_16554,N_16216);
nor UO_747 (O_747,N_18332,N_19371);
and UO_748 (O_748,N_15843,N_18986);
and UO_749 (O_749,N_16191,N_18724);
xnor UO_750 (O_750,N_16969,N_16420);
nand UO_751 (O_751,N_17870,N_15038);
nand UO_752 (O_752,N_19949,N_16627);
xor UO_753 (O_753,N_17234,N_19184);
and UO_754 (O_754,N_18333,N_18300);
nor UO_755 (O_755,N_18326,N_19869);
nand UO_756 (O_756,N_16578,N_19991);
xnor UO_757 (O_757,N_16668,N_15217);
nand UO_758 (O_758,N_19122,N_18512);
xnor UO_759 (O_759,N_15280,N_19154);
and UO_760 (O_760,N_16762,N_19115);
nor UO_761 (O_761,N_18955,N_17993);
xor UO_762 (O_762,N_19769,N_16075);
xor UO_763 (O_763,N_19691,N_15060);
xor UO_764 (O_764,N_15842,N_15446);
nand UO_765 (O_765,N_16848,N_16609);
and UO_766 (O_766,N_19030,N_17490);
nand UO_767 (O_767,N_15096,N_18238);
nor UO_768 (O_768,N_19649,N_17414);
nand UO_769 (O_769,N_18153,N_17246);
nor UO_770 (O_770,N_16910,N_18670);
nand UO_771 (O_771,N_17488,N_17104);
nand UO_772 (O_772,N_16270,N_19178);
or UO_773 (O_773,N_16103,N_18462);
or UO_774 (O_774,N_19250,N_18516);
or UO_775 (O_775,N_18715,N_17774);
xor UO_776 (O_776,N_16115,N_17789);
nand UO_777 (O_777,N_15534,N_18526);
and UO_778 (O_778,N_17922,N_15838);
or UO_779 (O_779,N_15690,N_17198);
xor UO_780 (O_780,N_16820,N_19027);
or UO_781 (O_781,N_15686,N_19144);
nor UO_782 (O_782,N_18797,N_19336);
and UO_783 (O_783,N_16995,N_18645);
nand UO_784 (O_784,N_16349,N_16702);
or UO_785 (O_785,N_16410,N_16367);
or UO_786 (O_786,N_19573,N_16679);
or UO_787 (O_787,N_16109,N_16493);
nand UO_788 (O_788,N_17745,N_17295);
or UO_789 (O_789,N_18355,N_17226);
xor UO_790 (O_790,N_18592,N_15672);
xor UO_791 (O_791,N_19186,N_16093);
xnor UO_792 (O_792,N_19358,N_17969);
and UO_793 (O_793,N_18812,N_17212);
xnor UO_794 (O_794,N_16106,N_16323);
and UO_795 (O_795,N_15548,N_19626);
or UO_796 (O_796,N_17874,N_19865);
nand UO_797 (O_797,N_18113,N_15262);
or UO_798 (O_798,N_16014,N_17631);
xnor UO_799 (O_799,N_17980,N_19714);
or UO_800 (O_800,N_15461,N_16389);
xnor UO_801 (O_801,N_19675,N_18865);
xnor UO_802 (O_802,N_16268,N_15504);
and UO_803 (O_803,N_16932,N_16502);
nand UO_804 (O_804,N_19911,N_17128);
and UO_805 (O_805,N_15808,N_18820);
nor UO_806 (O_806,N_16515,N_18573);
nor UO_807 (O_807,N_17144,N_16057);
and UO_808 (O_808,N_19191,N_19940);
or UO_809 (O_809,N_17693,N_15774);
and UO_810 (O_810,N_17566,N_19613);
or UO_811 (O_811,N_15999,N_18691);
nand UO_812 (O_812,N_19261,N_16169);
xnor UO_813 (O_813,N_19005,N_16173);
and UO_814 (O_814,N_16863,N_19239);
or UO_815 (O_815,N_17732,N_16819);
and UO_816 (O_816,N_15760,N_17189);
and UO_817 (O_817,N_15767,N_15064);
xnor UO_818 (O_818,N_19646,N_18767);
xor UO_819 (O_819,N_16962,N_15936);
and UO_820 (O_820,N_15870,N_18385);
or UO_821 (O_821,N_18503,N_16575);
nor UO_822 (O_822,N_19245,N_16541);
or UO_823 (O_823,N_16296,N_17349);
or UO_824 (O_824,N_18054,N_19380);
and UO_825 (O_825,N_17662,N_16760);
nor UO_826 (O_826,N_18331,N_16556);
nor UO_827 (O_827,N_19357,N_15031);
xor UO_828 (O_828,N_15348,N_16950);
or UO_829 (O_829,N_19403,N_19896);
nor UO_830 (O_830,N_15177,N_15820);
or UO_831 (O_831,N_16414,N_17432);
or UO_832 (O_832,N_18101,N_19411);
nor UO_833 (O_833,N_18619,N_18665);
xor UO_834 (O_834,N_16233,N_18000);
nor UO_835 (O_835,N_15650,N_17601);
nor UO_836 (O_836,N_17230,N_15371);
xnor UO_837 (O_837,N_19549,N_19280);
nor UO_838 (O_838,N_16655,N_17962);
or UO_839 (O_839,N_16961,N_19123);
xnor UO_840 (O_840,N_17607,N_17302);
nor UO_841 (O_841,N_17038,N_18379);
or UO_842 (O_842,N_16774,N_16630);
and UO_843 (O_843,N_18774,N_18410);
nand UO_844 (O_844,N_19596,N_19526);
or UO_845 (O_845,N_15783,N_19326);
xnor UO_846 (O_846,N_17909,N_16124);
and UO_847 (O_847,N_17014,N_15111);
nand UO_848 (O_848,N_19633,N_15302);
and UO_849 (O_849,N_16844,N_16567);
nand UO_850 (O_850,N_17916,N_16384);
nand UO_851 (O_851,N_16326,N_17899);
nand UO_852 (O_852,N_17559,N_17126);
and UO_853 (O_853,N_16920,N_17588);
or UO_854 (O_854,N_15130,N_18249);
xnor UO_855 (O_855,N_15519,N_16905);
and UO_856 (O_856,N_18056,N_15621);
and UO_857 (O_857,N_17176,N_17944);
nand UO_858 (O_858,N_18243,N_18239);
nand UO_859 (O_859,N_18038,N_15358);
or UO_860 (O_860,N_16737,N_19879);
xnor UO_861 (O_861,N_15200,N_19418);
xor UO_862 (O_862,N_16840,N_18849);
nand UO_863 (O_863,N_18036,N_16599);
and UO_864 (O_864,N_19228,N_16551);
xor UO_865 (O_865,N_15646,N_16091);
nand UO_866 (O_866,N_18154,N_18758);
or UO_867 (O_867,N_19840,N_17621);
nor UO_868 (O_868,N_19317,N_19092);
nor UO_869 (O_869,N_16249,N_17090);
and UO_870 (O_870,N_15638,N_16119);
and UO_871 (O_871,N_15403,N_18316);
nor UO_872 (O_872,N_15715,N_16946);
and UO_873 (O_873,N_18184,N_17273);
or UO_874 (O_874,N_18301,N_18589);
nor UO_875 (O_875,N_19398,N_18784);
xor UO_876 (O_876,N_16144,N_18118);
nand UO_877 (O_877,N_19015,N_15330);
nand UO_878 (O_878,N_18068,N_18576);
or UO_879 (O_879,N_17219,N_19693);
nor UO_880 (O_880,N_15406,N_19102);
nand UO_881 (O_881,N_17965,N_17070);
xnor UO_882 (O_882,N_18111,N_16938);
or UO_883 (O_883,N_15614,N_18974);
nand UO_884 (O_884,N_19121,N_16053);
nor UO_885 (O_885,N_17785,N_18824);
xor UO_886 (O_886,N_16716,N_19099);
nand UO_887 (O_887,N_19934,N_19684);
xor UO_888 (O_888,N_16589,N_15530);
nand UO_889 (O_889,N_17889,N_15429);
and UO_890 (O_890,N_17686,N_19671);
xnor UO_891 (O_891,N_15369,N_16033);
and UO_892 (O_892,N_19381,N_17497);
or UO_893 (O_893,N_19077,N_19352);
nand UO_894 (O_894,N_19583,N_18713);
nand UO_895 (O_895,N_18024,N_15865);
or UO_896 (O_896,N_18596,N_19295);
nand UO_897 (O_897,N_19860,N_16912);
or UO_898 (O_898,N_19848,N_18999);
and UO_899 (O_899,N_18528,N_16971);
xnor UO_900 (O_900,N_18554,N_18497);
nor UO_901 (O_901,N_16174,N_17722);
xor UO_902 (O_902,N_19782,N_15048);
nor UO_903 (O_903,N_15313,N_18531);
xnor UO_904 (O_904,N_19876,N_16276);
nand UO_905 (O_905,N_18174,N_16178);
nand UO_906 (O_906,N_17355,N_18095);
or UO_907 (O_907,N_17139,N_19087);
and UO_908 (O_908,N_15959,N_18123);
nor UO_909 (O_909,N_15730,N_16162);
and UO_910 (O_910,N_17987,N_16131);
and UO_911 (O_911,N_17875,N_16372);
or UO_912 (O_912,N_18307,N_19862);
and UO_913 (O_913,N_18941,N_15334);
and UO_914 (O_914,N_17039,N_15977);
nor UO_915 (O_915,N_19203,N_19391);
or UO_916 (O_916,N_18547,N_19975);
xnor UO_917 (O_917,N_17392,N_15225);
and UO_918 (O_918,N_19678,N_16054);
nand UO_919 (O_919,N_15351,N_17475);
nand UO_920 (O_920,N_19727,N_18190);
nor UO_921 (O_921,N_15727,N_18703);
nand UO_922 (O_922,N_16133,N_15338);
or UO_923 (O_923,N_17042,N_19766);
and UO_924 (O_924,N_18280,N_15622);
nor UO_925 (O_925,N_19255,N_15004);
xor UO_926 (O_926,N_15382,N_19821);
xnor UO_927 (O_927,N_18483,N_16225);
nor UO_928 (O_928,N_16134,N_16473);
nor UO_929 (O_929,N_17768,N_19595);
nand UO_930 (O_930,N_17760,N_18386);
or UO_931 (O_931,N_15355,N_16087);
and UO_932 (O_932,N_18117,N_16933);
and UO_933 (O_933,N_19961,N_15276);
and UO_934 (O_934,N_18842,N_18544);
and UO_935 (O_935,N_16487,N_18475);
nand UO_936 (O_936,N_19981,N_17536);
nor UO_937 (O_937,N_16514,N_18210);
nand UO_938 (O_938,N_17457,N_16992);
nand UO_939 (O_939,N_16795,N_17269);
xor UO_940 (O_940,N_15555,N_19713);
nand UO_941 (O_941,N_15257,N_18376);
nor UO_942 (O_942,N_19112,N_18897);
nand UO_943 (O_943,N_18233,N_15765);
and UO_944 (O_944,N_16229,N_18756);
and UO_945 (O_945,N_15943,N_18689);
and UO_946 (O_946,N_17216,N_18811);
xnor UO_947 (O_947,N_16289,N_19001);
nand UO_948 (O_948,N_16588,N_16895);
nor UO_949 (O_949,N_15668,N_16097);
xnor UO_950 (O_950,N_19262,N_15782);
nand UO_951 (O_951,N_16618,N_18532);
and UO_952 (O_952,N_19401,N_15699);
nand UO_953 (O_953,N_18887,N_17795);
nor UO_954 (O_954,N_19771,N_18474);
and UO_955 (O_955,N_19431,N_15537);
nor UO_956 (O_956,N_17203,N_15310);
nor UO_957 (O_957,N_17859,N_15920);
nand UO_958 (O_958,N_16732,N_19815);
nor UO_959 (O_959,N_16558,N_16161);
xor UO_960 (O_960,N_17866,N_18660);
or UO_961 (O_961,N_18975,N_15163);
xnor UO_962 (O_962,N_16141,N_19365);
nand UO_963 (O_963,N_15853,N_16510);
xnor UO_964 (O_964,N_16362,N_19568);
nor UO_965 (O_965,N_18035,N_16942);
nand UO_966 (O_966,N_15071,N_17005);
xnor UO_967 (O_967,N_17171,N_16965);
and UO_968 (O_968,N_18077,N_19157);
nor UO_969 (O_969,N_17143,N_18468);
xor UO_970 (O_970,N_19485,N_18695);
or UO_971 (O_971,N_19489,N_19168);
and UO_972 (O_972,N_16463,N_18364);
xnor UO_973 (O_973,N_18136,N_16565);
nand UO_974 (O_974,N_18681,N_19656);
xor UO_975 (O_975,N_19047,N_18289);
or UO_976 (O_976,N_16464,N_16433);
and UO_977 (O_977,N_17691,N_19264);
nand UO_978 (O_978,N_17667,N_15049);
and UO_979 (O_979,N_17187,N_17670);
nand UO_980 (O_980,N_15869,N_16851);
or UO_981 (O_981,N_15203,N_15491);
or UO_982 (O_982,N_16240,N_16479);
xor UO_983 (O_983,N_17199,N_16940);
nor UO_984 (O_984,N_17594,N_15669);
nor UO_985 (O_985,N_16781,N_15527);
or UO_986 (O_986,N_19867,N_17164);
and UO_987 (O_987,N_19531,N_18700);
xnor UO_988 (O_988,N_19376,N_17796);
nand UO_989 (O_989,N_19793,N_18362);
and UO_990 (O_990,N_15175,N_16399);
or UO_991 (O_991,N_19328,N_19972);
nor UO_992 (O_992,N_15952,N_17533);
and UO_993 (O_993,N_19687,N_18601);
nand UO_994 (O_994,N_18521,N_16357);
xnor UO_995 (O_995,N_16272,N_15931);
xor UO_996 (O_996,N_18821,N_16474);
xnor UO_997 (O_997,N_15533,N_15515);
or UO_998 (O_998,N_18492,N_16671);
and UO_999 (O_999,N_17054,N_17560);
nand UO_1000 (O_1000,N_18330,N_15899);
nand UO_1001 (O_1001,N_18055,N_18640);
and UO_1002 (O_1002,N_17808,N_16038);
xnor UO_1003 (O_1003,N_16311,N_18078);
and UO_1004 (O_1004,N_17229,N_17056);
or UO_1005 (O_1005,N_18563,N_17931);
and UO_1006 (O_1006,N_18216,N_16936);
or UO_1007 (O_1007,N_19748,N_18708);
xor UO_1008 (O_1008,N_19850,N_18433);
nor UO_1009 (O_1009,N_15771,N_19246);
nand UO_1010 (O_1010,N_16228,N_18500);
xnor UO_1011 (O_1011,N_19898,N_18796);
or UO_1012 (O_1012,N_17865,N_17160);
and UO_1013 (O_1013,N_18297,N_18467);
nor UO_1014 (O_1014,N_18940,N_18876);
and UO_1015 (O_1015,N_19757,N_19833);
nor UO_1016 (O_1016,N_17844,N_17781);
and UO_1017 (O_1017,N_15431,N_16506);
or UO_1018 (O_1018,N_17362,N_15971);
nand UO_1019 (O_1019,N_18605,N_17098);
nor UO_1020 (O_1020,N_15239,N_15364);
nor UO_1021 (O_1021,N_19453,N_17399);
or UO_1022 (O_1022,N_19202,N_19789);
nand UO_1023 (O_1023,N_15320,N_16559);
xor UO_1024 (O_1024,N_16984,N_18480);
xor UO_1025 (O_1025,N_19662,N_17180);
nand UO_1026 (O_1026,N_17208,N_16705);
nand UO_1027 (O_1027,N_19616,N_15713);
or UO_1028 (O_1028,N_15681,N_18489);
or UO_1029 (O_1029,N_17384,N_19063);
or UO_1030 (O_1030,N_17394,N_15653);
and UO_1031 (O_1031,N_17923,N_16631);
and UO_1032 (O_1032,N_15395,N_18453);
nand UO_1033 (O_1033,N_17373,N_18868);
or UO_1034 (O_1034,N_18541,N_16919);
nor UO_1035 (O_1035,N_17244,N_19939);
nand UO_1036 (O_1036,N_19218,N_19553);
and UO_1037 (O_1037,N_16557,N_17977);
xnor UO_1038 (O_1038,N_15929,N_15181);
nor UO_1039 (O_1039,N_17137,N_18395);
nand UO_1040 (O_1040,N_18145,N_19462);
and UO_1041 (O_1041,N_17755,N_15572);
and UO_1042 (O_1042,N_19216,N_19213);
xnor UO_1043 (O_1043,N_18504,N_19627);
nand UO_1044 (O_1044,N_15205,N_18706);
or UO_1045 (O_1045,N_15803,N_16593);
or UO_1046 (O_1046,N_19470,N_19253);
or UO_1047 (O_1047,N_17994,N_19895);
nand UO_1048 (O_1048,N_16128,N_18323);
nand UO_1049 (O_1049,N_17968,N_17849);
and UO_1050 (O_1050,N_17156,N_15974);
and UO_1051 (O_1051,N_17445,N_18069);
xnor UO_1052 (O_1052,N_18775,N_16619);
nand UO_1053 (O_1053,N_15994,N_17093);
xnor UO_1054 (O_1054,N_15168,N_15995);
and UO_1055 (O_1055,N_17352,N_16981);
xor UO_1056 (O_1056,N_15025,N_17900);
nand UO_1057 (O_1057,N_15722,N_15468);
nand UO_1058 (O_1058,N_17379,N_16012);
or UO_1059 (O_1059,N_15568,N_19534);
nor UO_1060 (O_1060,N_16574,N_15409);
and UO_1061 (O_1061,N_18649,N_17141);
nand UO_1062 (O_1062,N_18229,N_17807);
and UO_1063 (O_1063,N_18490,N_18981);
nand UO_1064 (O_1064,N_18156,N_15539);
and UO_1065 (O_1065,N_16481,N_15517);
or UO_1066 (O_1066,N_18494,N_19209);
nor UO_1067 (O_1067,N_18692,N_15790);
nand UO_1068 (O_1068,N_15029,N_16669);
or UO_1069 (O_1069,N_16154,N_18642);
xor UO_1070 (O_1070,N_15134,N_15304);
and UO_1071 (O_1071,N_19402,N_18854);
nand UO_1072 (O_1072,N_18760,N_17115);
xnor UO_1073 (O_1073,N_15377,N_18221);
nor UO_1074 (O_1074,N_18769,N_17211);
xnor UO_1075 (O_1075,N_18552,N_15485);
xnor UO_1076 (O_1076,N_19128,N_15347);
xnor UO_1077 (O_1077,N_16715,N_17233);
nand UO_1078 (O_1078,N_16665,N_17964);
nand UO_1079 (O_1079,N_15366,N_18891);
nor UO_1080 (O_1080,N_15845,N_16530);
nand UO_1081 (O_1081,N_18629,N_17609);
nand UO_1082 (O_1082,N_18032,N_18558);
xor UO_1083 (O_1083,N_18398,N_16224);
nand UO_1084 (O_1084,N_16242,N_16423);
xnor UO_1085 (O_1085,N_16027,N_16745);
xor UO_1086 (O_1086,N_18328,N_16232);
and UO_1087 (O_1087,N_15023,N_18934);
or UO_1088 (O_1088,N_18823,N_17151);
xor UO_1089 (O_1089,N_18408,N_17872);
nor UO_1090 (O_1090,N_19599,N_15471);
nor UO_1091 (O_1091,N_17835,N_17636);
xnor UO_1092 (O_1092,N_19145,N_16064);
nand UO_1093 (O_1093,N_19962,N_16041);
or UO_1094 (O_1094,N_15185,N_19728);
or UO_1095 (O_1095,N_16415,N_16310);
nor UO_1096 (O_1096,N_19504,N_17102);
or UO_1097 (O_1097,N_18091,N_17679);
nand UO_1098 (O_1098,N_17772,N_17957);
or UO_1099 (O_1099,N_19008,N_15408);
or UO_1100 (O_1100,N_19586,N_17625);
or UO_1101 (O_1101,N_17534,N_15256);
nor UO_1102 (O_1102,N_17334,N_19820);
nand UO_1103 (O_1103,N_17354,N_18250);
and UO_1104 (O_1104,N_17557,N_15401);
nor UO_1105 (O_1105,N_19082,N_17701);
nor UO_1106 (O_1106,N_18599,N_17249);
or UO_1107 (O_1107,N_16597,N_17064);
nor UO_1108 (O_1108,N_17336,N_15573);
nand UO_1109 (O_1109,N_17738,N_17391);
xor UO_1110 (O_1110,N_15231,N_19437);
xor UO_1111 (O_1111,N_18634,N_18367);
and UO_1112 (O_1112,N_18508,N_16342);
nor UO_1113 (O_1113,N_16635,N_16211);
nor UO_1114 (O_1114,N_15705,N_18083);
nor UO_1115 (O_1115,N_18878,N_18565);
and UO_1116 (O_1116,N_18585,N_19471);
or UO_1117 (O_1117,N_16494,N_16175);
xor UO_1118 (O_1118,N_18405,N_17599);
or UO_1119 (O_1119,N_15387,N_19151);
or UO_1120 (O_1120,N_16250,N_17291);
xnor UO_1121 (O_1121,N_19628,N_16834);
nor UO_1122 (O_1122,N_18218,N_16891);
xor UO_1123 (O_1123,N_18225,N_18793);
nor UO_1124 (O_1124,N_16063,N_15416);
xnor UO_1125 (O_1125,N_17851,N_15317);
nand UO_1126 (O_1126,N_15801,N_16581);
or UO_1127 (O_1127,N_18616,N_19007);
xor UO_1128 (O_1128,N_19464,N_17266);
xor UO_1129 (O_1129,N_17377,N_15798);
nand UO_1130 (O_1130,N_15709,N_19905);
nor UO_1131 (O_1131,N_18125,N_19735);
nand UO_1132 (O_1132,N_18694,N_17025);
and UO_1133 (O_1133,N_18013,N_19574);
nor UO_1134 (O_1134,N_18519,N_17708);
xor UO_1135 (O_1135,N_19935,N_19389);
and UO_1136 (O_1136,N_19956,N_19873);
nor UO_1137 (O_1137,N_17831,N_16878);
or UO_1138 (O_1138,N_18122,N_15103);
xnor UO_1139 (O_1139,N_18160,N_19477);
or UO_1140 (O_1140,N_15526,N_19204);
or UO_1141 (O_1141,N_16084,N_16517);
and UO_1142 (O_1142,N_19550,N_17210);
nand UO_1143 (O_1143,N_16909,N_18373);
or UO_1144 (O_1144,N_15992,N_18602);
and UO_1145 (O_1145,N_18771,N_15698);
or UO_1146 (O_1146,N_15930,N_19536);
xor UO_1147 (O_1147,N_16303,N_16498);
nand UO_1148 (O_1148,N_19118,N_15417);
xnor UO_1149 (O_1149,N_17780,N_16652);
and UO_1150 (O_1150,N_15068,N_15009);
nand UO_1151 (O_1151,N_15565,N_16189);
xor UO_1152 (O_1152,N_16235,N_17847);
or UO_1153 (O_1153,N_17067,N_19368);
or UO_1154 (O_1154,N_19754,N_15744);
or UO_1155 (O_1155,N_19792,N_15102);
nand UO_1156 (O_1156,N_15211,N_17404);
nor UO_1157 (O_1157,N_19524,N_15763);
xor UO_1158 (O_1158,N_18352,N_19139);
or UO_1159 (O_1159,N_19758,N_17888);
xnor UO_1160 (O_1160,N_19463,N_15147);
or UO_1161 (O_1161,N_15091,N_18074);
xnor UO_1162 (O_1162,N_18426,N_19971);
or UO_1163 (O_1163,N_18015,N_15261);
and UO_1164 (O_1164,N_18211,N_16939);
nand UO_1165 (O_1165,N_17806,N_18586);
or UO_1166 (O_1166,N_18663,N_18465);
or UO_1167 (O_1167,N_15524,N_19277);
or UO_1168 (O_1168,N_15370,N_16082);
and UO_1169 (O_1169,N_15691,N_16294);
or UO_1170 (O_1170,N_19912,N_19048);
nor UO_1171 (O_1171,N_18988,N_19608);
xor UO_1172 (O_1172,N_16869,N_19672);
xor UO_1173 (O_1173,N_16312,N_15176);
or UO_1174 (O_1174,N_15795,N_18905);
and UO_1175 (O_1175,N_18050,N_19592);
nor UO_1176 (O_1176,N_17283,N_17626);
nand UO_1177 (O_1177,N_17558,N_16908);
nand UO_1178 (O_1178,N_17136,N_18176);
nor UO_1179 (O_1179,N_15354,N_15326);
or UO_1180 (O_1180,N_18957,N_17346);
nand UO_1181 (O_1181,N_18253,N_15815);
nand UO_1182 (O_1182,N_19469,N_16392);
or UO_1183 (O_1183,N_16924,N_19302);
nor UO_1184 (O_1184,N_19747,N_19137);
xnor UO_1185 (O_1185,N_16422,N_17570);
xor UO_1186 (O_1186,N_19441,N_15652);
nand UO_1187 (O_1187,N_18132,N_16158);
and UO_1188 (O_1188,N_15328,N_15016);
nor UO_1189 (O_1189,N_16386,N_15522);
xnor UO_1190 (O_1190,N_15857,N_18237);
or UO_1191 (O_1191,N_18646,N_17048);
nor UO_1192 (O_1192,N_15298,N_17240);
xnor UO_1193 (O_1193,N_19645,N_17696);
nor UO_1194 (O_1194,N_16746,N_17506);
and UO_1195 (O_1195,N_18653,N_17836);
or UO_1196 (O_1196,N_15495,N_17456);
nand UO_1197 (O_1197,N_16777,N_19055);
or UO_1198 (O_1198,N_17967,N_15978);
nand UO_1199 (O_1199,N_17867,N_15296);
nor UO_1200 (O_1200,N_18151,N_16945);
nand UO_1201 (O_1201,N_16266,N_15055);
or UO_1202 (O_1202,N_18514,N_17682);
nor UO_1203 (O_1203,N_15725,N_18027);
nor UO_1204 (O_1204,N_17300,N_18360);
nor UO_1205 (O_1205,N_15270,N_17406);
nand UO_1206 (O_1206,N_19603,N_15305);
nand UO_1207 (O_1207,N_19752,N_17075);
nand UO_1208 (O_1208,N_15046,N_15352);
xor UO_1209 (O_1209,N_15116,N_17304);
or UO_1210 (O_1210,N_19406,N_15024);
nand UO_1211 (O_1211,N_16333,N_19756);
xnor UO_1212 (O_1212,N_19472,N_18661);
and UO_1213 (O_1213,N_19936,N_17361);
and UO_1214 (O_1214,N_19276,N_18914);
nand UO_1215 (O_1215,N_19829,N_16157);
xor UO_1216 (O_1216,N_18321,N_15858);
nor UO_1217 (O_1217,N_19878,N_15260);
nand UO_1218 (O_1218,N_19773,N_19607);
xor UO_1219 (O_1219,N_15972,N_19944);
xor UO_1220 (O_1220,N_18375,N_17868);
nor UO_1221 (O_1221,N_18654,N_16190);
nand UO_1222 (O_1222,N_19967,N_16104);
xor UO_1223 (O_1223,N_18384,N_15848);
nand UO_1224 (O_1224,N_18420,N_15098);
and UO_1225 (O_1225,N_19964,N_18273);
and UO_1226 (O_1226,N_16281,N_16790);
or UO_1227 (O_1227,N_17942,N_15538);
and UO_1228 (O_1228,N_15856,N_16720);
and UO_1229 (O_1229,N_18137,N_18578);
nor UO_1230 (O_1230,N_19241,N_19555);
or UO_1231 (O_1231,N_17008,N_18662);
or UO_1232 (O_1232,N_17963,N_15212);
and UO_1233 (O_1233,N_17581,N_18926);
xnor UO_1234 (O_1234,N_17063,N_15289);
xor UO_1235 (O_1235,N_18874,N_17678);
xnor UO_1236 (O_1236,N_16316,N_15913);
and UO_1237 (O_1237,N_16089,N_18044);
or UO_1238 (O_1238,N_18268,N_15450);
and UO_1239 (O_1239,N_15062,N_15950);
xor UO_1240 (O_1240,N_18641,N_17207);
xnor UO_1241 (O_1241,N_17464,N_15595);
or UO_1242 (O_1242,N_19643,N_15862);
or UO_1243 (O_1243,N_17611,N_16674);
or UO_1244 (O_1244,N_17877,N_17424);
xnor UO_1245 (O_1245,N_19397,N_19224);
or UO_1246 (O_1246,N_19259,N_19834);
and UO_1247 (O_1247,N_19292,N_16380);
nor UO_1248 (O_1248,N_17804,N_18311);
or UO_1249 (O_1249,N_18344,N_15224);
or UO_1250 (O_1250,N_17973,N_18597);
nor UO_1251 (O_1251,N_19301,N_15553);
nor UO_1252 (O_1252,N_19075,N_16313);
nand UO_1253 (O_1253,N_15489,N_17124);
and UO_1254 (O_1254,N_16875,N_19516);
nand UO_1255 (O_1255,N_18173,N_19637);
and UO_1256 (O_1256,N_16264,N_19955);
xnor UO_1257 (O_1257,N_15356,N_18752);
nor UO_1258 (O_1258,N_15367,N_18265);
xnor UO_1259 (O_1259,N_16317,N_18003);
xor UO_1260 (O_1260,N_15141,N_18904);
or UO_1261 (O_1261,N_17812,N_19493);
xor UO_1262 (O_1262,N_18299,N_17651);
xor UO_1263 (O_1263,N_18826,N_17083);
nor UO_1264 (O_1264,N_15149,N_15569);
nor UO_1265 (O_1265,N_19387,N_16085);
and UO_1266 (O_1266,N_15908,N_16615);
nand UO_1267 (O_1267,N_18058,N_18523);
xnor UO_1268 (O_1268,N_16491,N_17930);
nor UO_1269 (O_1269,N_17758,N_15499);
nor UO_1270 (O_1270,N_15906,N_18569);
nand UO_1271 (O_1271,N_16262,N_19779);
nand UO_1272 (O_1272,N_17803,N_17907);
and UO_1273 (O_1273,N_19893,N_19297);
xnor UO_1274 (O_1274,N_16478,N_19435);
xnor UO_1275 (O_1275,N_17978,N_18899);
xnor UO_1276 (O_1276,N_19995,N_16398);
xnor UO_1277 (O_1277,N_19739,N_16955);
or UO_1278 (O_1278,N_18073,N_15607);
nor UO_1279 (O_1279,N_16653,N_18466);
or UO_1280 (O_1280,N_17084,N_18409);
or UO_1281 (O_1281,N_17433,N_18086);
or UO_1282 (O_1282,N_19808,N_15850);
xor UO_1283 (O_1283,N_15359,N_15169);
xnor UO_1284 (O_1284,N_17627,N_19653);
and UO_1285 (O_1285,N_18099,N_15559);
and UO_1286 (O_1286,N_15393,N_17153);
and UO_1287 (O_1287,N_19223,N_17477);
xor UO_1288 (O_1288,N_18622,N_19664);
nand UO_1289 (O_1289,N_18746,N_18913);
or UO_1290 (O_1290,N_17152,N_15574);
nor UO_1291 (O_1291,N_16894,N_17943);
or UO_1292 (O_1292,N_16990,N_17500);
nand UO_1293 (O_1293,N_16201,N_19229);
xor UO_1294 (O_1294,N_19394,N_17368);
xnor UO_1295 (O_1295,N_18567,N_16448);
or UO_1296 (O_1296,N_19043,N_17524);
and UO_1297 (O_1297,N_17850,N_18604);
and UO_1298 (O_1298,N_18016,N_19744);
nand UO_1299 (O_1299,N_18258,N_19530);
and UO_1300 (O_1300,N_17917,N_16736);
nand UO_1301 (O_1301,N_17855,N_15343);
nand UO_1302 (O_1302,N_17472,N_15007);
nor UO_1303 (O_1303,N_18045,N_16177);
nand UO_1304 (O_1304,N_17869,N_16661);
nand UO_1305 (O_1305,N_16107,N_17052);
xnor UO_1306 (O_1306,N_18079,N_15837);
nor UO_1307 (O_1307,N_19410,N_17802);
nand UO_1308 (O_1308,N_16982,N_19529);
and UO_1309 (O_1309,N_16328,N_15703);
nand UO_1310 (O_1310,N_17348,N_18898);
and UO_1311 (O_1311,N_18591,N_18127);
nor UO_1312 (O_1312,N_16278,N_19554);
nor UO_1313 (O_1313,N_16527,N_16944);
or UO_1314 (O_1314,N_15716,N_16327);
nand UO_1315 (O_1315,N_18428,N_19452);
xor UO_1316 (O_1316,N_17430,N_15719);
or UO_1317 (O_1317,N_15566,N_17753);
xnor UO_1318 (O_1318,N_16171,N_16988);
or UO_1319 (O_1319,N_19567,N_17021);
or UO_1320 (O_1320,N_16184,N_19590);
nor UO_1321 (O_1321,N_19062,N_17970);
nor UO_1322 (O_1322,N_19619,N_19767);
nand UO_1323 (O_1323,N_18915,N_15314);
and UO_1324 (O_1324,N_15481,N_17161);
nand UO_1325 (O_1325,N_17951,N_16904);
nor UO_1326 (O_1326,N_15020,N_16145);
or UO_1327 (O_1327,N_17666,N_19252);
or UO_1328 (O_1328,N_17507,N_17431);
and UO_1329 (O_1329,N_17754,N_15924);
nor UO_1330 (O_1330,N_17501,N_15019);
or UO_1331 (O_1331,N_19513,N_19618);
or UO_1332 (O_1332,N_19701,N_18928);
or UO_1333 (O_1333,N_17903,N_16741);
nor UO_1334 (O_1334,N_16403,N_16748);
nand UO_1335 (O_1335,N_19338,N_16670);
or UO_1336 (O_1336,N_18635,N_18515);
and UO_1337 (O_1337,N_18220,N_16906);
and UO_1338 (O_1338,N_16284,N_16205);
nor UO_1339 (O_1339,N_19373,N_19528);
or UO_1340 (O_1340,N_18369,N_19997);
xor UO_1341 (O_1341,N_18121,N_15807);
nand UO_1342 (O_1342,N_16416,N_18680);
nand UO_1343 (O_1343,N_16044,N_16019);
nor UO_1344 (O_1344,N_15127,N_18768);
nor UO_1345 (O_1345,N_17285,N_15768);
nor UO_1346 (O_1346,N_19160,N_16183);
nor UO_1347 (O_1347,N_16791,N_16656);
or UO_1348 (O_1348,N_16055,N_17108);
or UO_1349 (O_1349,N_18582,N_16329);
xnor UO_1350 (O_1350,N_15230,N_16858);
nor UO_1351 (O_1351,N_16489,N_15309);
nor UO_1352 (O_1352,N_18805,N_19369);
nor UO_1353 (O_1353,N_17786,N_17731);
nand UO_1354 (O_1354,N_19650,N_18736);
xnor UO_1355 (O_1355,N_17468,N_15635);
and UO_1356 (O_1356,N_19430,N_17119);
and UO_1357 (O_1357,N_18857,N_17004);
nand UO_1358 (O_1358,N_17323,N_16136);
or UO_1359 (O_1359,N_16787,N_16274);
nor UO_1360 (O_1360,N_16553,N_16838);
nor UO_1361 (O_1361,N_19478,N_16396);
and UO_1362 (O_1362,N_15228,N_15590);
and UO_1363 (O_1363,N_16550,N_18830);
nand UO_1364 (O_1364,N_17653,N_18972);
nand UO_1365 (O_1365,N_17684,N_17146);
and UO_1366 (O_1366,N_19809,N_19537);
nand UO_1367 (O_1367,N_19990,N_17749);
xor UO_1368 (O_1368,N_19461,N_19928);
or UO_1369 (O_1369,N_19176,N_15927);
nand UO_1370 (O_1370,N_16750,N_15932);
nand UO_1371 (O_1371,N_18652,N_17383);
xor UO_1372 (O_1372,N_15576,N_19564);
nor UO_1373 (O_1373,N_18482,N_16911);
nor UO_1374 (O_1374,N_17097,N_18446);
or UO_1375 (O_1375,N_19396,N_15208);
or UO_1376 (O_1376,N_18188,N_19770);
nor UO_1377 (O_1377,N_19640,N_16043);
and UO_1378 (O_1378,N_19225,N_16980);
and UO_1379 (O_1379,N_16622,N_18836);
nor UO_1380 (O_1380,N_16437,N_16778);
and UO_1381 (O_1381,N_16841,N_17474);
or UO_1382 (O_1382,N_18062,N_19141);
nor UO_1383 (O_1383,N_17562,N_17407);
xor UO_1384 (O_1384,N_19417,N_19012);
and UO_1385 (O_1385,N_18391,N_18371);
and UO_1386 (O_1386,N_18051,N_15993);
nand UO_1387 (O_1387,N_16797,N_17523);
and UO_1388 (O_1388,N_19922,N_19169);
and UO_1389 (O_1389,N_15237,N_16523);
nor UO_1390 (O_1390,N_15741,N_19853);
and UO_1391 (O_1391,N_18770,N_17897);
nor UO_1392 (O_1392,N_15056,N_19342);
xor UO_1393 (O_1393,N_17597,N_15165);
or UO_1394 (O_1394,N_17615,N_15077);
xnor UO_1395 (O_1395,N_15960,N_19717);
nor UO_1396 (O_1396,N_17012,N_18977);
nand UO_1397 (O_1397,N_16857,N_17257);
nor UO_1398 (O_1398,N_15779,N_19899);
and UO_1399 (O_1399,N_18533,N_15087);
nor UO_1400 (O_1400,N_18126,N_18256);
and UO_1401 (O_1401,N_17476,N_16370);
nand UO_1402 (O_1402,N_18675,N_19197);
nand UO_1403 (O_1403,N_18741,N_15603);
nor UO_1404 (O_1404,N_18840,N_15946);
nor UO_1405 (O_1405,N_16913,N_18906);
nand UO_1406 (O_1406,N_17510,N_15439);
nor UO_1407 (O_1407,N_16130,N_19318);
xnor UO_1408 (O_1408,N_16831,N_18447);
nor UO_1409 (O_1409,N_15874,N_15613);
xnor UO_1410 (O_1410,N_15585,N_19812);
nand UO_1411 (O_1411,N_19348,N_17107);
nand UO_1412 (O_1412,N_19527,N_16529);
nand UO_1413 (O_1413,N_19587,N_17890);
nand UO_1414 (O_1414,N_15105,N_19644);
nand UO_1415 (O_1415,N_15385,N_16698);
and UO_1416 (O_1416,N_18870,N_15435);
nor UO_1417 (O_1417,N_19965,N_17736);
nor UO_1418 (O_1418,N_15011,N_17325);
nor UO_1419 (O_1419,N_15051,N_16881);
or UO_1420 (O_1420,N_18194,N_15425);
nor UO_1421 (O_1421,N_17853,N_19970);
or UO_1422 (O_1422,N_17183,N_15349);
xor UO_1423 (O_1423,N_19938,N_16883);
and UO_1424 (O_1424,N_15125,N_15506);
and UO_1425 (O_1425,N_17116,N_16290);
and UO_1426 (O_1426,N_15708,N_15496);
and UO_1427 (O_1427,N_15787,N_18738);
nor UO_1428 (O_1428,N_16722,N_19654);
nor UO_1429 (O_1429,N_17434,N_17057);
xnor UO_1430 (O_1430,N_18120,N_15810);
nor UO_1431 (O_1431,N_17814,N_15694);
xor UO_1432 (O_1432,N_18685,N_16607);
xor UO_1433 (O_1433,N_17982,N_15290);
xor UO_1434 (O_1434,N_15316,N_16072);
and UO_1435 (O_1435,N_15723,N_16538);
and UO_1436 (O_1436,N_17934,N_19232);
or UO_1437 (O_1437,N_16049,N_18020);
and UO_1438 (O_1438,N_18023,N_17296);
nor UO_1439 (O_1439,N_17341,N_17282);
nor UO_1440 (O_1440,N_17567,N_16400);
nand UO_1441 (O_1441,N_19924,N_15402);
nand UO_1442 (O_1442,N_17593,N_16826);
nor UO_1443 (O_1443,N_15003,N_17663);
or UO_1444 (O_1444,N_16234,N_16763);
nor UO_1445 (O_1445,N_15047,N_16371);
nor UO_1446 (O_1446,N_19916,N_19871);
nor UO_1447 (O_1447,N_16504,N_19360);
xnor UO_1448 (O_1448,N_16540,N_16334);
and UO_1449 (O_1449,N_16186,N_18042);
and UO_1450 (O_1450,N_18076,N_16412);
and UO_1451 (O_1451,N_16587,N_17420);
and UO_1452 (O_1452,N_17425,N_18096);
nor UO_1453 (O_1453,N_18501,N_15702);
nand UO_1454 (O_1454,N_18666,N_18026);
xor UO_1455 (O_1455,N_19765,N_15441);
or UO_1456 (O_1456,N_19919,N_16230);
nor UO_1457 (O_1457,N_19993,N_18912);
nand UO_1458 (O_1458,N_19872,N_18971);
nand UO_1459 (O_1459,N_17816,N_16717);
nand UO_1460 (O_1460,N_15655,N_19450);
nand UO_1461 (O_1461,N_16193,N_16378);
and UO_1462 (O_1462,N_15114,N_15540);
nand UO_1463 (O_1463,N_16706,N_18809);
nand UO_1464 (O_1464,N_18557,N_18404);
or UO_1465 (O_1465,N_16534,N_16431);
nand UO_1466 (O_1466,N_18334,N_15288);
or UO_1467 (O_1467,N_18112,N_17123);
or UO_1468 (O_1468,N_17953,N_17201);
xor UO_1469 (O_1469,N_16220,N_16432);
nand UO_1470 (O_1470,N_18227,N_16918);
or UO_1471 (O_1471,N_15322,N_19310);
nor UO_1472 (O_1472,N_19142,N_18476);
nor UO_1473 (O_1473,N_19605,N_19856);
nand UO_1474 (O_1474,N_15769,N_15039);
nand UO_1475 (O_1475,N_18850,N_19495);
nor UO_1476 (O_1476,N_17287,N_15544);
xor UO_1477 (O_1477,N_19548,N_17000);
or UO_1478 (O_1478,N_18712,N_17910);
and UO_1479 (O_1479,N_15684,N_16023);
and UO_1480 (O_1480,N_15651,N_19969);
nor UO_1481 (O_1481,N_15005,N_17629);
xor UO_1482 (O_1482,N_15113,N_18178);
or UO_1483 (O_1483,N_18267,N_16634);
xnor UO_1484 (O_1484,N_16018,N_17690);
or UO_1485 (O_1485,N_16694,N_18236);
and UO_1486 (O_1486,N_15424,N_19036);
nor UO_1487 (O_1487,N_19058,N_17680);
or UO_1488 (O_1488,N_18399,N_17306);
and UO_1489 (O_1489,N_15751,N_18423);
nand UO_1490 (O_1490,N_15511,N_18285);
or UO_1491 (O_1491,N_17142,N_18085);
nor UO_1492 (O_1492,N_19138,N_18436);
or UO_1493 (O_1493,N_18202,N_19926);
or UO_1494 (O_1494,N_19432,N_16877);
nand UO_1495 (O_1495,N_15518,N_19538);
xnor UO_1496 (O_1496,N_15109,N_15584);
or UO_1497 (O_1497,N_17612,N_17235);
and UO_1498 (O_1498,N_19510,N_17380);
xor UO_1499 (O_1499,N_18158,N_18260);
and UO_1500 (O_1500,N_17773,N_18192);
or UO_1501 (O_1501,N_16245,N_15881);
nor UO_1502 (O_1502,N_19694,N_18293);
and UO_1503 (O_1503,N_19337,N_18839);
xnor UO_1504 (O_1504,N_15909,N_19943);
nor UO_1505 (O_1505,N_18935,N_16776);
xor UO_1506 (O_1506,N_17829,N_16138);
xor UO_1507 (O_1507,N_19824,N_17195);
or UO_1508 (O_1508,N_18002,N_17860);
and UO_1509 (O_1509,N_17927,N_18838);
nand UO_1510 (O_1510,N_17743,N_15278);
nand UO_1511 (O_1511,N_18175,N_16029);
nand UO_1512 (O_1512,N_15182,N_15101);
and UO_1513 (O_1513,N_17096,N_19364);
and UO_1514 (O_1514,N_19113,N_17182);
and UO_1515 (O_1515,N_19194,N_17073);
or UO_1516 (O_1516,N_17429,N_15456);
nand UO_1517 (O_1517,N_15773,N_16690);
xor UO_1518 (O_1518,N_16495,N_19159);
and UO_1519 (O_1519,N_16257,N_16972);
or UO_1520 (O_1520,N_17527,N_16842);
nor UO_1521 (O_1521,N_18918,N_15161);
or UO_1522 (O_1522,N_18816,N_16815);
xnor UO_1523 (O_1523,N_18908,N_15953);
or UO_1524 (O_1524,N_15339,N_19269);
or UO_1525 (O_1525,N_19105,N_18669);
or UO_1526 (O_1526,N_15251,N_15879);
and UO_1527 (O_1527,N_17074,N_18200);
or UO_1528 (O_1528,N_15140,N_18832);
xor UO_1529 (O_1529,N_16450,N_17614);
and UO_1530 (O_1530,N_17482,N_19711);
nand UO_1531 (O_1531,N_16353,N_18223);
or UO_1532 (O_1532,N_15818,N_16074);
and UO_1533 (O_1533,N_18938,N_15656);
nand UO_1534 (O_1534,N_15965,N_17712);
nor UO_1535 (O_1535,N_19424,N_18947);
nor UO_1536 (O_1536,N_18415,N_17112);
xnor UO_1537 (O_1537,N_16005,N_16922);
nor UO_1538 (O_1538,N_15193,N_15411);
nand UO_1539 (O_1539,N_18534,N_15440);
and UO_1540 (O_1540,N_18687,N_15903);
xnor UO_1541 (O_1541,N_17734,N_19697);
xor UO_1542 (O_1542,N_18499,N_19804);
and UO_1543 (O_1543,N_17747,N_18786);
and UO_1544 (O_1544,N_15501,N_19585);
or UO_1545 (O_1545,N_19136,N_19346);
and UO_1546 (O_1546,N_19497,N_15154);
xor UO_1547 (O_1547,N_18228,N_15636);
or UO_1548 (O_1548,N_15855,N_15236);
nor UO_1549 (O_1549,N_16236,N_16148);
and UO_1550 (O_1550,N_19947,N_15721);
nor UO_1551 (O_1551,N_19976,N_19073);
or UO_1552 (O_1552,N_16600,N_18656);
xnor UO_1553 (O_1553,N_15259,N_15080);
or UO_1554 (O_1554,N_16358,N_19986);
nor UO_1555 (O_1555,N_18624,N_18944);
or UO_1556 (O_1556,N_18808,N_17032);
nor UO_1557 (O_1557,N_16802,N_15954);
xor UO_1558 (O_1558,N_19308,N_19566);
and UO_1559 (O_1559,N_17671,N_17081);
nor UO_1560 (O_1560,N_16890,N_19201);
or UO_1561 (O_1561,N_16062,N_17106);
xnor UO_1562 (O_1562,N_19046,N_15189);
xnor UO_1563 (O_1563,N_17059,N_18147);
or UO_1564 (O_1564,N_15907,N_17218);
nand UO_1565 (O_1565,N_18880,N_18374);
xnor UO_1566 (O_1566,N_18631,N_16299);
xor UO_1567 (O_1567,N_16346,N_17591);
xor UO_1568 (O_1568,N_16318,N_19428);
nand UO_1569 (O_1569,N_19026,N_18648);
or UO_1570 (O_1570,N_18421,N_15167);
and UO_1571 (O_1571,N_18072,N_16213);
nor UO_1572 (O_1572,N_17730,N_16803);
and UO_1573 (O_1573,N_18978,N_16991);
nor UO_1574 (O_1574,N_15283,N_15545);
nor UO_1575 (O_1575,N_15935,N_18901);
and UO_1576 (O_1576,N_17518,N_17748);
and UO_1577 (O_1577,N_18046,N_19340);
nor UO_1578 (O_1578,N_16728,N_15153);
nand UO_1579 (O_1579,N_18525,N_16711);
or UO_1580 (O_1580,N_18325,N_16424);
nor UO_1581 (O_1581,N_19542,N_15895);
nor UO_1582 (O_1582,N_17491,N_17101);
nand UO_1583 (O_1583,N_19795,N_17834);
xnor UO_1584 (O_1584,N_17168,N_19064);
nor UO_1585 (O_1585,N_15292,N_15991);
or UO_1586 (O_1586,N_16304,N_15413);
or UO_1587 (O_1587,N_15308,N_15476);
xor UO_1588 (O_1588,N_18443,N_17028);
nand UO_1589 (O_1589,N_15531,N_16002);
xnor UO_1590 (O_1590,N_17645,N_16628);
or UO_1591 (O_1591,N_16319,N_16179);
nor UO_1592 (O_1592,N_16165,N_17498);
or UO_1593 (O_1593,N_15321,N_15792);
or UO_1594 (O_1594,N_16957,N_17659);
nor UO_1595 (O_1595,N_15596,N_17550);
or UO_1596 (O_1596,N_15860,N_17725);
and UO_1597 (O_1597,N_19189,N_16194);
and UO_1598 (O_1598,N_16521,N_19059);
xnor UO_1599 (O_1599,N_19091,N_17985);
nand UO_1600 (O_1600,N_19688,N_17604);
nand UO_1601 (O_1601,N_15265,N_16341);
nor UO_1602 (O_1602,N_16069,N_19889);
xor UO_1603 (O_1603,N_17879,N_16123);
nand UO_1604 (O_1604,N_18457,N_17131);
nor UO_1605 (O_1605,N_15171,N_16218);
or UO_1606 (O_1606,N_18608,N_19330);
nand UO_1607 (O_1607,N_15557,N_19106);
nand UO_1608 (O_1608,N_16114,N_19844);
and UO_1609 (O_1609,N_16896,N_15287);
or UO_1610 (O_1610,N_16237,N_15645);
and UO_1611 (O_1611,N_15509,N_17739);
or UO_1612 (O_1612,N_18431,N_16893);
or UO_1613 (O_1613,N_18039,N_15044);
nand UO_1614 (O_1614,N_18028,N_17658);
xor UO_1615 (O_1615,N_16735,N_19025);
and UO_1616 (O_1616,N_18737,N_15018);
nor UO_1617 (O_1617,N_19220,N_15824);
or UO_1618 (O_1618,N_16719,N_17639);
nand UO_1619 (O_1619,N_16395,N_16862);
xnor UO_1620 (O_1620,N_18748,N_17723);
and UO_1621 (O_1621,N_15868,N_17487);
or UO_1622 (O_1622,N_18469,N_19621);
xnor UO_1623 (O_1623,N_15467,N_15523);
and UO_1624 (O_1624,N_17237,N_15987);
nand UO_1625 (O_1625,N_16042,N_15386);
nor UO_1626 (O_1626,N_17842,N_19796);
nand UO_1627 (O_1627,N_17268,N_17531);
and UO_1628 (O_1628,N_19561,N_19454);
xor UO_1629 (O_1629,N_17826,N_19124);
and UO_1630 (O_1630,N_19476,N_15285);
nor UO_1631 (O_1631,N_18464,N_17405);
nor UO_1632 (O_1632,N_19569,N_18885);
xor UO_1633 (O_1633,N_19442,N_18396);
xor UO_1634 (O_1634,N_19427,N_17882);
nor UO_1635 (O_1635,N_16325,N_17742);
nand UO_1636 (O_1636,N_16564,N_16710);
nor UO_1637 (O_1637,N_17617,N_18511);
or UO_1638 (O_1638,N_18152,N_18686);
nor UO_1639 (O_1639,N_15541,N_19511);
and UO_1640 (O_1640,N_19279,N_17342);
nor UO_1641 (O_1641,N_19864,N_19010);
or UO_1642 (O_1642,N_16917,N_19891);
and UO_1643 (O_1643,N_16126,N_16345);
and UO_1644 (O_1644,N_16552,N_16485);
nand UO_1645 (O_1645,N_18788,N_15707);
or UO_1646 (O_1646,N_19960,N_15381);
nor UO_1647 (O_1647,N_18262,N_19520);
or UO_1648 (O_1648,N_19588,N_18064);
nand UO_1649 (O_1649,N_15345,N_17460);
nand UO_1650 (O_1650,N_16305,N_15252);
nor UO_1651 (O_1651,N_16667,N_18454);
nor UO_1652 (O_1652,N_16512,N_17382);
xor UO_1653 (O_1653,N_16611,N_19291);
xor UO_1654 (O_1654,N_15197,N_15329);
or UO_1655 (O_1655,N_18419,N_15610);
nand UO_1656 (O_1656,N_16034,N_19089);
xnor UO_1657 (O_1657,N_15137,N_18614);
nand UO_1658 (O_1658,N_19620,N_15547);
or UO_1659 (O_1659,N_18041,N_18861);
nand UO_1660 (O_1660,N_16659,N_15027);
xor UO_1661 (O_1661,N_19825,N_18109);
and UO_1662 (O_1662,N_17439,N_16682);
and UO_1663 (O_1663,N_16031,N_19446);
xor UO_1664 (O_1664,N_18933,N_19760);
or UO_1665 (O_1665,N_19069,N_17169);
nor UO_1666 (O_1666,N_18937,N_19045);
nand UO_1667 (O_1667,N_17375,N_18789);
or UO_1668 (O_1668,N_15618,N_17415);
xnor UO_1669 (O_1669,N_17637,N_19130);
and UO_1670 (O_1670,N_16612,N_16752);
xnor UO_1671 (O_1671,N_18235,N_19888);
nor UO_1672 (O_1672,N_15268,N_15788);
xor UO_1673 (O_1673,N_18397,N_19161);
xor UO_1674 (O_1674,N_18472,N_19913);
nand UO_1675 (O_1675,N_15186,N_16212);
xor UO_1676 (O_1676,N_18149,N_18791);
xor UO_1677 (O_1677,N_16703,N_17321);
nand UO_1678 (O_1678,N_16685,N_19349);
nor UO_1679 (O_1679,N_15642,N_16000);
nand UO_1680 (O_1680,N_16923,N_18010);
xor UO_1681 (O_1681,N_15673,N_18674);
nor UO_1682 (O_1682,N_16767,N_19037);
xor UO_1683 (O_1683,N_16522,N_16579);
nand UO_1684 (O_1684,N_15667,N_17577);
nor UO_1685 (O_1685,N_15198,N_16146);
nor UO_1686 (O_1686,N_17440,N_18498);
and UO_1687 (O_1687,N_16402,N_18232);
or UO_1688 (O_1688,N_19004,N_17565);
nand UO_1689 (O_1689,N_18848,N_19325);
and UO_1690 (O_1690,N_16903,N_16182);
nor UO_1691 (O_1691,N_15449,N_17502);
or UO_1692 (O_1692,N_16207,N_16935);
nor UO_1693 (O_1693,N_15084,N_15336);
xnor UO_1694 (O_1694,N_16636,N_18623);
nor UO_1695 (O_1695,N_19481,N_19716);
and UO_1696 (O_1696,N_17087,N_18677);
nand UO_1697 (O_1697,N_18291,N_19843);
or UO_1698 (O_1698,N_19594,N_19571);
nand UO_1699 (O_1699,N_19356,N_17154);
nand UO_1700 (O_1700,N_17493,N_19404);
nor UO_1701 (O_1701,N_15836,N_17929);
xor UO_1702 (O_1702,N_19890,N_16846);
nor UO_1703 (O_1703,N_18780,N_15459);
and UO_1704 (O_1704,N_16925,N_19475);
nand UO_1705 (O_1705,N_15301,N_18728);
nand UO_1706 (O_1706,N_18363,N_18958);
nor UO_1707 (O_1707,N_17117,N_19885);
nand UO_1708 (O_1708,N_16931,N_16595);
nor UO_1709 (O_1709,N_18104,N_15215);
nand UO_1710 (O_1710,N_19434,N_19248);
xnor UO_1711 (O_1711,N_17225,N_17709);
and UO_1712 (O_1712,N_19539,N_17413);
or UO_1713 (O_1713,N_18437,N_15172);
nor UO_1714 (O_1714,N_16483,N_19395);
xor UO_1715 (O_1715,N_18005,N_16065);
nand UO_1716 (O_1716,N_15986,N_18754);
nand UO_1717 (O_1717,N_17060,N_18833);
nor UO_1718 (O_1718,N_19230,N_18477);
nand UO_1719 (O_1719,N_18496,N_17437);
nand UO_1720 (O_1720,N_18657,N_15928);
or UO_1721 (O_1721,N_17111,N_19942);
and UO_1722 (O_1722,N_19419,N_15145);
or UO_1723 (O_1723,N_19484,N_17885);
or UO_1724 (O_1724,N_18102,N_15560);
or UO_1725 (O_1725,N_17015,N_17279);
nor UO_1726 (O_1726,N_19482,N_19781);
nand UO_1727 (O_1727,N_15512,N_16051);
or UO_1728 (O_1728,N_19405,N_17194);
xor UO_1729 (O_1729,N_18618,N_15353);
nand UO_1730 (O_1730,N_18723,N_17793);
nand UO_1731 (O_1731,N_17608,N_19429);
nand UO_1732 (O_1732,N_18561,N_17130);
or UO_1733 (O_1733,N_17041,N_19287);
and UO_1734 (O_1734,N_16789,N_19135);
nand UO_1735 (O_1735,N_18452,N_17654);
xnor UO_1736 (O_1736,N_15873,N_16508);
and UO_1737 (O_1737,N_15248,N_19622);
xnor UO_1738 (O_1738,N_17248,N_19021);
and UO_1739 (O_1739,N_17664,N_17148);
and UO_1740 (O_1740,N_18390,N_17402);
and UO_1741 (O_1741,N_15996,N_18970);
nor UO_1742 (O_1742,N_15095,N_15556);
or UO_1743 (O_1743,N_19705,N_18658);
nand UO_1744 (O_1744,N_15457,N_15859);
or UO_1745 (O_1745,N_17016,N_16772);
and UO_1746 (O_1746,N_18277,N_19651);
xor UO_1747 (O_1747,N_15422,N_19031);
or UO_1748 (O_1748,N_17544,N_19284);
xor UO_1749 (O_1749,N_17876,N_15558);
xor UO_1750 (O_1750,N_18925,N_16937);
nor UO_1751 (O_1751,N_18450,N_16978);
xor UO_1752 (O_1752,N_18761,N_18684);
nand UO_1753 (O_1753,N_18945,N_19642);
xor UO_1754 (O_1754,N_18911,N_16428);
or UO_1755 (O_1755,N_16164,N_16699);
nor UO_1756 (O_1756,N_15090,N_17630);
xor UO_1757 (O_1757,N_18263,N_18266);
nor UO_1758 (O_1758,N_17316,N_15764);
nor UO_1759 (O_1759,N_18559,N_18459);
nand UO_1760 (O_1760,N_16050,N_16094);
xor UO_1761 (O_1761,N_19183,N_16605);
xor UO_1762 (O_1762,N_18302,N_17883);
nor UO_1763 (O_1763,N_16419,N_15081);
and UO_1764 (O_1764,N_18894,N_19584);
or UO_1765 (O_1765,N_16282,N_17605);
and UO_1766 (O_1766,N_17155,N_15350);
or UO_1767 (O_1767,N_15398,N_16335);
xor UO_1768 (O_1768,N_19256,N_16686);
xor UO_1769 (O_1769,N_16998,N_17033);
nand UO_1770 (O_1770,N_16393,N_17242);
nand UO_1771 (O_1771,N_15490,N_17389);
nor UO_1772 (O_1772,N_15759,N_15166);
xor UO_1773 (O_1773,N_16016,N_15331);
and UO_1774 (O_1774,N_15312,N_17956);
xor UO_1775 (O_1775,N_17264,N_16076);
xor UO_1776 (O_1776,N_19902,N_18907);
nand UO_1777 (O_1777,N_18438,N_17981);
nor UO_1778 (O_1778,N_17901,N_18734);
and UO_1779 (O_1779,N_19681,N_17983);
xnor UO_1780 (O_1780,N_17775,N_17486);
and UO_1781 (O_1781,N_15663,N_17521);
and UO_1782 (O_1782,N_19777,N_15832);
and UO_1783 (O_1783,N_16430,N_17683);
or UO_1784 (O_1784,N_16202,N_19333);
nand UO_1785 (O_1785,N_19505,N_16900);
or UO_1786 (O_1786,N_15617,N_17920);
nand UO_1787 (O_1787,N_16813,N_18030);
or UO_1788 (O_1788,N_18043,N_16839);
xor UO_1789 (O_1789,N_16885,N_17172);
nand UO_1790 (O_1790,N_17376,N_18288);
xor UO_1791 (O_1791,N_19315,N_16640);
nor UO_1792 (O_1792,N_16964,N_19819);
nand UO_1793 (O_1793,N_16200,N_19413);
xnor UO_1794 (O_1794,N_17790,N_18683);
nor UO_1795 (O_1795,N_18822,N_16352);
or UO_1796 (O_1796,N_17129,N_16078);
and UO_1797 (O_1797,N_15670,N_19695);
xnor UO_1798 (O_1798,N_16277,N_16660);
and UO_1799 (O_1799,N_18792,N_19006);
xnor UO_1800 (O_1800,N_15640,N_16608);
or UO_1801 (O_1801,N_15588,N_18365);
nor UO_1802 (O_1802,N_16039,N_15396);
nor UO_1803 (O_1803,N_18875,N_15497);
and UO_1804 (O_1804,N_15187,N_15478);
or UO_1805 (O_1805,N_17623,N_19577);
xnor UO_1806 (O_1806,N_17125,N_18869);
xor UO_1807 (O_1807,N_19845,N_15740);
or UO_1808 (O_1808,N_18505,N_17517);
nand UO_1809 (O_1809,N_18542,N_16426);
and UO_1810 (O_1810,N_18283,N_15833);
nor UO_1811 (O_1811,N_18481,N_15882);
nor UO_1812 (O_1812,N_16168,N_15361);
nor UO_1813 (O_1813,N_19002,N_18110);
nor UO_1814 (O_1814,N_17213,N_17937);
xnor UO_1815 (O_1815,N_19268,N_17540);
and UO_1816 (O_1816,N_16696,N_18164);
nand UO_1817 (O_1817,N_16195,N_17086);
or UO_1818 (O_1818,N_15045,N_18545);
or UO_1819 (O_1819,N_15915,N_16676);
nand UO_1820 (O_1820,N_16275,N_19733);
and UO_1821 (O_1821,N_17861,N_18275);
or UO_1822 (O_1822,N_19535,N_18637);
and UO_1823 (O_1823,N_18048,N_16324);
and UO_1824 (O_1824,N_16860,N_16692);
xnor UO_1825 (O_1825,N_19039,N_15346);
xor UO_1826 (O_1826,N_18159,N_17294);
nand UO_1827 (O_1827,N_19351,N_15094);
nor UO_1828 (O_1828,N_18867,N_18416);
nand UO_1829 (O_1829,N_16308,N_17455);
or UO_1830 (O_1830,N_19061,N_15129);
nand UO_1831 (O_1831,N_15463,N_16172);
nor UO_1832 (O_1832,N_18722,N_16960);
xor UO_1833 (O_1833,N_16260,N_17792);
nor UO_1834 (O_1834,N_15549,N_19591);
or UO_1835 (O_1835,N_15724,N_16516);
nand UO_1836 (O_1836,N_16927,N_15883);
or UO_1837 (O_1837,N_15164,N_15484);
nor UO_1838 (O_1838,N_18195,N_16560);
xnor UO_1839 (O_1839,N_19883,N_19496);
or UO_1840 (O_1840,N_18018,N_15551);
and UO_1841 (O_1841,N_16782,N_17674);
nand UO_1842 (O_1842,N_18180,N_16449);
and UO_1843 (O_1843,N_18090,N_17779);
and UO_1844 (O_1844,N_17741,N_19335);
nand UO_1845 (O_1845,N_16073,N_19093);
or UO_1846 (O_1846,N_15150,N_19468);
and UO_1847 (O_1847,N_15122,N_19959);
or UO_1848 (O_1848,N_15135,N_17989);
nand UO_1849 (O_1849,N_16117,N_19219);
xor UO_1850 (O_1850,N_18308,N_16843);
nor UO_1851 (O_1851,N_16132,N_18927);
nor UO_1852 (O_1852,N_15604,N_16930);
nor UO_1853 (O_1853,N_16949,N_16806);
or UO_1854 (O_1854,N_15985,N_18628);
nor UO_1855 (O_1855,N_19837,N_16783);
or UO_1856 (O_1856,N_17633,N_15249);
xnor UO_1857 (O_1857,N_18463,N_15979);
nand UO_1858 (O_1858,N_19344,N_17817);
and UO_1859 (O_1859,N_16309,N_18417);
nor UO_1860 (O_1860,N_19589,N_18810);
and UO_1861 (O_1861,N_17469,N_17080);
nand UO_1862 (O_1862,N_17766,N_19057);
xor UO_1863 (O_1863,N_17600,N_18172);
and UO_1864 (O_1864,N_18031,N_15914);
or UO_1865 (O_1865,N_15594,N_18007);
xnor UO_1866 (O_1866,N_18594,N_17347);
nor UO_1867 (O_1867,N_17825,N_16513);
nor UO_1868 (O_1868,N_17979,N_17109);
nor UO_1869 (O_1869,N_15758,N_15194);
nor UO_1870 (O_1870,N_18358,N_16867);
and UO_1871 (O_1871,N_17192,N_15383);
or UO_1872 (O_1872,N_15532,N_17499);
nor UO_1873 (O_1873,N_15427,N_19233);
xnor UO_1874 (O_1874,N_17438,N_18994);
and UO_1875 (O_1875,N_18148,N_15170);
and UO_1876 (O_1876,N_15814,N_19941);
xnor UO_1877 (O_1877,N_18441,N_15938);
or UO_1878 (O_1878,N_15412,N_15878);
xor UO_1879 (O_1879,N_19096,N_15063);
xnor UO_1880 (O_1880,N_19601,N_15372);
or UO_1881 (O_1881,N_17250,N_17810);
nand UO_1882 (O_1882,N_18053,N_19980);
and UO_1883 (O_1883,N_17677,N_15391);
or UO_1884 (O_1884,N_16359,N_17585);
nor UO_1885 (O_1885,N_16730,N_16497);
xnor UO_1886 (O_1886,N_19384,N_16066);
nor UO_1887 (O_1887,N_16592,N_15887);
xnor UO_1888 (O_1888,N_18106,N_19547);
and UO_1889 (O_1889,N_16662,N_18664);
xor UO_1890 (O_1890,N_16382,N_16654);
nand UO_1891 (O_1891,N_19996,N_18400);
nand UO_1892 (O_1892,N_19013,N_16377);
nor UO_1893 (O_1893,N_16738,N_16536);
nor UO_1894 (O_1894,N_16928,N_18310);
and UO_1895 (O_1895,N_16110,N_17905);
nor UO_1896 (O_1896,N_19179,N_19017);
or UO_1897 (O_1897,N_15849,N_15877);
or UO_1898 (O_1898,N_15054,N_18882);
and UO_1899 (O_1899,N_15104,N_15697);
or UO_1900 (O_1900,N_18458,N_19127);
xor UO_1901 (O_1901,N_16181,N_19669);
nor UO_1902 (O_1902,N_15898,N_16941);
xnor UO_1903 (O_1903,N_17442,N_17113);
and UO_1904 (O_1904,N_19708,N_17791);
or UO_1905 (O_1905,N_17628,N_18964);
nand UO_1906 (O_1906,N_19377,N_19999);
or UO_1907 (O_1907,N_15811,N_16417);
nor UO_1908 (O_1908,N_16492,N_16761);
nor UO_1909 (O_1909,N_19658,N_19147);
xor UO_1910 (O_1910,N_15195,N_18342);
nor UO_1911 (O_1911,N_17514,N_15606);
nand UO_1912 (O_1912,N_16827,N_16068);
nand UO_1913 (O_1913,N_18726,N_18580);
nand UO_1914 (O_1914,N_16629,N_19412);
nor UO_1915 (O_1915,N_19925,N_17846);
and UO_1916 (O_1916,N_19457,N_15711);
nand UO_1917 (O_1917,N_15133,N_16870);
nor UO_1918 (O_1918,N_18138,N_17887);
or UO_1919 (O_1919,N_15772,N_15535);
nand UO_1920 (O_1920,N_18553,N_19827);
nand UO_1921 (O_1921,N_16780,N_18422);
or UO_1922 (O_1922,N_18939,N_15207);
or UO_1923 (O_1923,N_16967,N_16253);
or UO_1924 (O_1924,N_18259,N_18214);
and UO_1925 (O_1925,N_19260,N_15250);
nand UO_1926 (O_1926,N_18633,N_18212);
nor UO_1927 (O_1927,N_19909,N_19763);
nand UO_1928 (O_1928,N_18757,N_19131);
nor UO_1929 (O_1929,N_15654,N_17757);
nand UO_1930 (O_1930,N_19778,N_16477);
nand UO_1931 (O_1931,N_16347,N_16766);
or UO_1932 (O_1932,N_19696,N_19187);
nor UO_1933 (O_1933,N_17286,N_17289);
or UO_1934 (O_1934,N_15712,N_18019);
nand UO_1935 (O_1935,N_17941,N_15139);
nand UO_1936 (O_1936,N_17841,N_17896);
xor UO_1937 (O_1937,N_18506,N_15597);
or UO_1938 (O_1938,N_18979,N_17991);
xor UO_1939 (O_1939,N_15390,N_19953);
nor UO_1940 (O_1940,N_19580,N_15513);
nand UO_1941 (O_1941,N_18219,N_17071);
and UO_1942 (O_1942,N_17105,N_19579);
xnor UO_1943 (O_1943,N_18286,N_19797);
xor UO_1944 (O_1944,N_19718,N_16354);
nor UO_1945 (O_1945,N_19266,N_15616);
nor UO_1946 (O_1946,N_16373,N_18655);
xor UO_1947 (O_1947,N_15222,N_18389);
nand UO_1948 (O_1948,N_18461,N_19181);
xnor UO_1949 (O_1949,N_18181,N_17094);
xnor UO_1950 (O_1950,N_17938,N_15847);
xnor UO_1951 (O_1951,N_18613,N_17127);
xor UO_1952 (O_1952,N_15957,N_17913);
xor UO_1953 (O_1953,N_19226,N_18888);
xor UO_1954 (O_1954,N_19088,N_16712);
and UO_1955 (O_1955,N_19114,N_19551);
xnor UO_1956 (O_1956,N_16035,N_17002);
xnor UO_1957 (O_1957,N_18800,N_15327);
nand UO_1958 (O_1958,N_16267,N_15846);
or UO_1959 (O_1959,N_15966,N_17238);
nand UO_1960 (O_1960,N_17703,N_15428);
nand UO_1961 (O_1961,N_18281,N_18245);
xnor UO_1962 (O_1962,N_18382,N_19835);
nor UO_1963 (O_1963,N_18448,N_19182);
and UO_1964 (O_1964,N_15743,N_16524);
nand UO_1965 (O_1965,N_15831,N_18884);
and UO_1966 (O_1966,N_19612,N_15910);
nor UO_1967 (O_1967,N_18107,N_15234);
nand UO_1968 (O_1968,N_15866,N_16677);
xnor UO_1969 (O_1969,N_19448,N_18522);
or UO_1970 (O_1970,N_16125,N_17298);
or UO_1971 (O_1971,N_18799,N_19707);
or UO_1972 (O_1972,N_18860,N_18383);
nand UO_1973 (O_1973,N_19307,N_16973);
or UO_1974 (O_1974,N_16010,N_19519);
nor UO_1975 (O_1975,N_15817,N_17554);
and UO_1976 (O_1976,N_16704,N_18976);
and UO_1977 (O_1977,N_15736,N_18418);
nor UO_1978 (O_1978,N_15941,N_16902);
nand UO_1979 (O_1979,N_18588,N_17019);
nor UO_1980 (O_1980,N_19321,N_15079);
nor UO_1981 (O_1981,N_19140,N_18909);
xnor UO_1982 (O_1982,N_18312,N_15677);
xor UO_1983 (O_1983,N_19690,N_17448);
nor UO_1984 (O_1984,N_17223,N_16444);
xor UO_1985 (O_1985,N_15092,N_17996);
or UO_1986 (O_1986,N_18451,N_17546);
xor UO_1987 (O_1987,N_16739,N_17068);
nand UO_1988 (O_1988,N_18114,N_15756);
xnor UO_1989 (O_1989,N_15692,N_19049);
nand UO_1990 (O_1990,N_18581,N_18676);
xnor UO_1991 (O_1991,N_15067,N_19623);
xor UO_1992 (O_1992,N_16800,N_15357);
nand UO_1993 (O_1993,N_19081,N_16872);
or UO_1994 (O_1994,N_17036,N_15968);
or UO_1995 (O_1995,N_19517,N_17408);
nor UO_1996 (O_1996,N_17961,N_16823);
and UO_1997 (O_1997,N_17366,N_18008);
and UO_1998 (O_1998,N_17528,N_17390);
and UO_1999 (O_1999,N_19285,N_18859);
xor UO_2000 (O_2000,N_17228,N_16976);
and UO_2001 (O_2001,N_15340,N_19152);
nor UO_2002 (O_2002,N_19945,N_16404);
or UO_2003 (O_2003,N_15373,N_18279);
xor UO_2004 (O_2004,N_16429,N_17288);
and UO_2005 (O_2005,N_16271,N_15254);
nand UO_2006 (O_2006,N_17256,N_18982);
or UO_2007 (O_2007,N_17026,N_17572);
nor UO_2008 (O_2008,N_17326,N_19416);
or UO_2009 (O_2009,N_18025,N_18550);
and UO_2010 (O_2010,N_19984,N_15323);
xor UO_2011 (O_2011,N_19998,N_18787);
nand UO_2012 (O_2012,N_17893,N_19900);
or UO_2013 (O_2013,N_18873,N_15233);
nand UO_2014 (O_2014,N_19177,N_19875);
xnor UO_2015 (O_2015,N_15443,N_15678);
nand UO_2016 (O_2016,N_15514,N_19734);
or UO_2017 (O_2017,N_17330,N_16596);
xnor UO_2018 (O_2018,N_15601,N_15676);
or UO_2019 (O_2019,N_19674,N_18537);
and UO_2020 (O_2020,N_19683,N_15631);
xor UO_2021 (O_2021,N_18762,N_17317);
and UO_2022 (O_2022,N_19164,N_19198);
xnor UO_2023 (O_2023,N_18829,N_17293);
xor UO_2024 (O_2024,N_17397,N_19040);
nand UO_2025 (O_2025,N_15796,N_16531);
xnor UO_2026 (O_2026,N_15948,N_19283);
or UO_2027 (O_2027,N_15426,N_19165);
nand UO_2028 (O_2028,N_19932,N_16003);
and UO_2029 (O_2029,N_15138,N_15612);
nand UO_2030 (O_2030,N_18562,N_18948);
xor UO_2031 (O_2031,N_19314,N_15839);
nand UO_2032 (O_2032,N_16543,N_15477);
xor UO_2033 (O_2033,N_18337,N_15458);
xor UO_2034 (O_2034,N_16407,N_16256);
xnor UO_2035 (O_2035,N_17580,N_18638);
or UO_2036 (O_2036,N_19507,N_17275);
or UO_2037 (O_2037,N_19060,N_15854);
nand UO_2038 (O_2038,N_15641,N_19034);
or UO_2039 (O_2039,N_15380,N_19423);
xnor UO_2040 (O_2040,N_19525,N_18401);
nand UO_2041 (O_2041,N_18742,N_18987);
and UO_2042 (O_2042,N_16447,N_15344);
nand UO_2043 (O_2043,N_15561,N_19173);
xor UO_2044 (O_2044,N_18430,N_16365);
xnor UO_2045 (O_2045,N_19863,N_15300);
nand UO_2046 (O_2046,N_19712,N_16300);
nor UO_2047 (O_2047,N_15981,N_18209);
or UO_2048 (O_2048,N_18954,N_16188);
and UO_2049 (O_2049,N_19372,N_15777);
nand UO_2050 (O_2050,N_18851,N_16223);
nand UO_2051 (O_2051,N_19207,N_19982);
and UO_2052 (O_2052,N_15685,N_16792);
nor UO_2053 (O_2053,N_16469,N_17428);
xnor UO_2054 (O_2054,N_16098,N_17231);
nand UO_2055 (O_2055,N_16151,N_18535);
nor UO_2056 (O_2056,N_16963,N_17066);
and UO_2057 (O_2057,N_17830,N_17673);
xnor UO_2058 (O_2058,N_15498,N_15630);
nor UO_2059 (O_2059,N_16059,N_17069);
and UO_2060 (O_2060,N_18942,N_16360);
nor UO_2061 (O_2061,N_15643,N_18612);
or UO_2062 (O_2062,N_15342,N_15890);
nor UO_2063 (O_2063,N_15378,N_18714);
or UO_2064 (O_2064,N_19363,N_17914);
nor UO_2065 (O_2065,N_15374,N_19359);
nand UO_2066 (O_2066,N_17552,N_15432);
nor UO_2067 (O_2067,N_15562,N_15376);
or UO_2068 (O_2068,N_19028,N_16954);
and UO_2069 (O_2069,N_15384,N_16248);
or UO_2070 (O_2070,N_17586,N_16689);
or UO_2071 (O_2071,N_15017,N_19783);
nor UO_2072 (O_2072,N_18377,N_19799);
nand UO_2073 (O_2073,N_16387,N_17737);
nand UO_2074 (O_2074,N_16811,N_16484);
xnor UO_2075 (O_2075,N_15360,N_16280);
xor UO_2076 (O_2076,N_15013,N_16460);
nand UO_2077 (O_2077,N_19304,N_17079);
nor UO_2078 (O_2078,N_16482,N_16733);
nand UO_2079 (O_2079,N_15099,N_18339);
xor UO_2080 (O_2080,N_15637,N_19722);
or UO_2081 (O_2081,N_17100,N_16379);
and UO_2082 (O_2082,N_16490,N_19479);
and UO_2083 (O_2083,N_16355,N_19686);
nor UO_2084 (O_2084,N_17158,N_18524);
and UO_2085 (O_2085,N_18710,N_18776);
nor UO_2086 (O_2086,N_19859,N_18207);
and UO_2087 (O_2087,N_18698,N_19638);
nor UO_2088 (O_2088,N_17023,N_18598);
nand UO_2089 (O_2089,N_17343,N_16152);
nor UO_2090 (O_2090,N_19068,N_18996);
and UO_2091 (O_2091,N_18702,N_16646);
nand UO_2092 (O_2092,N_18837,N_15001);
and UO_2093 (O_2093,N_17174,N_16681);
and UO_2094 (O_2094,N_19486,N_16691);
and UO_2095 (O_2095,N_17547,N_18261);
or UO_2096 (O_2096,N_19680,N_19729);
nand UO_2097 (O_2097,N_18314,N_17260);
and UO_2098 (O_2098,N_16320,N_16898);
nand UO_2099 (O_2099,N_15008,N_19038);
nand UO_2100 (O_2100,N_16570,N_19298);
and UO_2101 (O_2101,N_17419,N_18893);
and UO_2102 (O_2102,N_17040,N_16295);
nand UO_2103 (O_2103,N_16156,N_18507);
xor UO_2104 (O_2104,N_17699,N_17955);
and UO_2105 (O_2105,N_16569,N_16708);
nor UO_2106 (O_2106,N_17571,N_17541);
xor UO_2107 (O_2107,N_15620,N_18572);
nor UO_2108 (O_2108,N_17029,N_18169);
or UO_2109 (O_2109,N_16273,N_16576);
xnor UO_2110 (O_2110,N_15241,N_18251);
and UO_2111 (O_2111,N_17857,N_18766);
xnor UO_2112 (O_2112,N_18061,N_15813);
xor UO_2113 (O_2113,N_18052,N_15206);
nor UO_2114 (O_2114,N_17398,N_19354);
and UO_2115 (O_2115,N_18932,N_18881);
nand UO_2116 (O_2116,N_15131,N_17058);
nor UO_2117 (O_2117,N_18747,N_19846);
xor UO_2118 (O_2118,N_17492,N_19515);
nor UO_2119 (O_2119,N_18071,N_16434);
and UO_2120 (O_2120,N_19272,N_19700);
xnor UO_2121 (O_2121,N_16283,N_18847);
or UO_2122 (O_2122,N_15279,N_19050);
and UO_2123 (O_2123,N_19362,N_15900);
or UO_2124 (O_2124,N_19200,N_16751);
nor UO_2125 (O_2125,N_15179,N_15209);
and UO_2126 (O_2126,N_16771,N_15052);
or UO_2127 (O_2127,N_18536,N_19035);
nand UO_2128 (O_2128,N_16687,N_18115);
nand UO_2129 (O_2129,N_18318,N_19663);
nor UO_2130 (O_2130,N_16788,N_16999);
nand UO_2131 (O_2131,N_19235,N_15570);
nand UO_2132 (O_2132,N_15926,N_18949);
nand UO_2133 (O_2133,N_16390,N_16901);
nor UO_2134 (O_2134,N_17839,N_19051);
and UO_2135 (O_2135,N_18479,N_16880);
xnor UO_2136 (O_2136,N_16197,N_17644);
nor UO_2137 (O_2137,N_19263,N_15589);
and UO_2138 (O_2138,N_19078,N_19836);
or UO_2139 (O_2139,N_17583,N_18886);
nor UO_2140 (O_2140,N_18098,N_15742);
and UO_2141 (O_2141,N_19375,N_17276);
or UO_2142 (O_2142,N_17714,N_16263);
or UO_2143 (O_2143,N_17767,N_15118);
xor UO_2144 (O_2144,N_15582,N_18548);
and UO_2145 (O_2145,N_17367,N_15158);
nand UO_2146 (O_2146,N_15421,N_16825);
or UO_2147 (O_2147,N_15591,N_18697);
or UO_2148 (O_2148,N_17915,N_18414);
and UO_2149 (O_2149,N_17687,N_16011);
and UO_2150 (O_2150,N_19558,N_18727);
nor UO_2151 (O_2151,N_15120,N_17277);
or UO_2152 (O_2152,N_15246,N_15460);
xnor UO_2153 (O_2153,N_16808,N_18732);
nor UO_2154 (O_2154,N_15940,N_15508);
and UO_2155 (O_2155,N_15445,N_18201);
nor UO_2156 (O_2156,N_19436,N_16645);
and UO_2157 (O_2157,N_17952,N_18493);
xnor UO_2158 (O_2158,N_18831,N_16585);
nor UO_2159 (O_2159,N_15482,N_17184);
nand UO_2160 (O_2160,N_19698,N_19868);
nor UO_2161 (O_2161,N_16643,N_18773);
and UO_2162 (O_2162,N_15112,N_19153);
nor UO_2163 (O_2163,N_19881,N_15706);
nand UO_2164 (O_2164,N_19560,N_16227);
xnor UO_2165 (O_2165,N_19180,N_17805);
xnor UO_2166 (O_2166,N_16832,N_16167);
xor UO_2167 (O_2167,N_17706,N_16142);
nand UO_2168 (O_2168,N_17222,N_19514);
nor UO_2169 (O_2169,N_16472,N_17655);
nand UO_2170 (O_2170,N_18351,N_17350);
xnor UO_2171 (O_2171,N_17239,N_16459);
or UO_2172 (O_2172,N_19930,N_18141);
or UO_2173 (O_2173,N_17034,N_18671);
or UO_2174 (O_2174,N_18167,N_18495);
nand UO_2175 (O_2175,N_15634,N_17253);
nand UO_2176 (O_2176,N_15649,N_15050);
nor UO_2177 (O_2177,N_19832,N_15666);
or UO_2178 (O_2178,N_16683,N_15272);
nor UO_2179 (O_2179,N_17165,N_17975);
or UO_2180 (O_2180,N_16718,N_19289);
xor UO_2181 (O_2181,N_15700,N_16046);
or UO_2182 (O_2182,N_16351,N_18060);
nor UO_2183 (O_2183,N_18063,N_17520);
nand UO_2184 (O_2184,N_19817,N_19665);
or UO_2185 (O_2185,N_19828,N_19842);
xnor UO_2186 (O_2186,N_16364,N_18066);
nor UO_2187 (O_2187,N_19449,N_18936);
nor UO_2188 (O_2188,N_15739,N_15223);
nor UO_2189 (O_2189,N_15057,N_15058);
and UO_2190 (O_2190,N_16958,N_15066);
nand UO_2191 (O_2191,N_18460,N_17435);
or UO_2192 (O_2192,N_17214,N_17327);
nand UO_2193 (O_2193,N_16793,N_15174);
nor UO_2194 (O_2194,N_17274,N_15492);
nand UO_2195 (O_2195,N_17661,N_18203);
or UO_2196 (O_2196,N_17727,N_17459);
nor UO_2197 (O_2197,N_17720,N_16518);
and UO_2198 (O_2198,N_18733,N_15732);
nor UO_2199 (O_2199,N_16221,N_17205);
xor UO_2200 (O_2200,N_18844,N_19083);
nor UO_2201 (O_2201,N_16040,N_16856);
or UO_2202 (O_2202,N_16723,N_18555);
xor UO_2203 (O_2203,N_17261,N_15227);
or UO_2204 (O_2204,N_18320,N_17089);
or UO_2205 (O_2205,N_19275,N_16734);
or UO_2206 (O_2206,N_16537,N_18556);
or UO_2207 (O_2207,N_17815,N_19305);
or UO_2208 (O_2208,N_15554,N_19053);
nor UO_2209 (O_2209,N_19794,N_19565);
xnor UO_2210 (O_2210,N_18116,N_17787);
xnor UO_2211 (O_2211,N_15680,N_18278);
xnor UO_2212 (O_2212,N_16026,N_17881);
or UO_2213 (O_2213,N_15053,N_15797);
nand UO_2214 (O_2214,N_18134,N_17186);
or UO_2215 (O_2215,N_17166,N_17863);
xor UO_2216 (O_2216,N_16547,N_18889);
and UO_2217 (O_2217,N_16852,N_18720);
or UO_2218 (O_2218,N_17549,N_17132);
and UO_2219 (O_2219,N_18924,N_17574);
xnor UO_2220 (O_2220,N_19545,N_16500);
xor UO_2221 (O_2221,N_18966,N_17563);
and UO_2222 (O_2222,N_18445,N_17756);
xor UO_2223 (O_2223,N_17595,N_16443);
or UO_2224 (O_2224,N_19546,N_18029);
xor UO_2225 (O_2225,N_16344,N_19166);
and UO_2226 (O_2226,N_18424,N_17873);
nor UO_2227 (O_2227,N_19270,N_16147);
nor UO_2228 (O_2228,N_15695,N_19451);
nor UO_2229 (O_2229,N_16397,N_17444);
and UO_2230 (O_2230,N_16874,N_18449);
and UO_2231 (O_2231,N_19659,N_16907);
nand UO_2232 (O_2232,N_15089,N_16914);
xor UO_2233 (O_2233,N_17092,N_19831);
xnor UO_2234 (O_2234,N_18284,N_17995);
xor UO_2235 (O_2235,N_19784,N_16709);
and UO_2236 (O_2236,N_19386,N_16647);
xnor UO_2237 (O_2237,N_16639,N_15379);
nand UO_2238 (O_2238,N_16269,N_15750);
and UO_2239 (O_2239,N_19421,N_15488);
or UO_2240 (O_2240,N_19901,N_15657);
and UO_2241 (O_2241,N_18247,N_17800);
nand UO_2242 (O_2242,N_17660,N_19080);
and UO_2243 (O_2243,N_18744,N_18434);
nand UO_2244 (O_2244,N_18317,N_19639);
xnor UO_2245 (O_2245,N_15030,N_15921);
or UO_2246 (O_2246,N_17110,N_18731);
nor UO_2247 (O_2247,N_15980,N_18004);
nand UO_2248 (O_2248,N_15748,N_15436);
or UO_2249 (O_2249,N_18103,N_15776);
nand UO_2250 (O_2250,N_16030,N_15754);
and UO_2251 (O_2251,N_15144,N_15647);
nand UO_2252 (O_2252,N_16408,N_15275);
and UO_2253 (O_2253,N_16036,N_16617);
and UO_2254 (O_2254,N_17532,N_18241);
or UO_2255 (O_2255,N_19920,N_18246);
nor UO_2256 (O_2256,N_18471,N_18162);
and UO_2257 (O_2257,N_17778,N_19271);
nor UO_2258 (O_2258,N_19880,N_15623);
nor UO_2259 (O_2259,N_19673,N_19715);
xor UO_2260 (O_2260,N_17764,N_17410);
or UO_2261 (O_2261,N_19458,N_17797);
nor UO_2262 (O_2262,N_17467,N_15525);
nand UO_2263 (O_2263,N_15453,N_16673);
and UO_2264 (O_2264,N_18890,N_17838);
xnor UO_2265 (O_2265,N_16020,N_19952);
xnor UO_2266 (O_2266,N_16770,N_19190);
nor UO_2267 (O_2267,N_18186,N_17926);
nor UO_2268 (O_2268,N_18108,N_18006);
and UO_2269 (O_2269,N_17884,N_18197);
and UO_2270 (O_2270,N_15923,N_17265);
and UO_2271 (O_2271,N_17078,N_15078);
and UO_2272 (O_2272,N_19286,N_19719);
xnor UO_2273 (O_2273,N_17454,N_18088);
xnor UO_2274 (O_2274,N_18705,N_16475);
nor UO_2275 (O_2275,N_15633,N_19572);
nand UO_2276 (O_2276,N_16185,N_15933);
xnor UO_2277 (O_2277,N_17958,N_18411);
nand UO_2278 (O_2278,N_17374,N_18828);
nor UO_2279 (O_2279,N_15204,N_18549);
nand UO_2280 (O_2280,N_17954,N_18740);
nand UO_2281 (O_2281,N_16102,N_17465);
nand UO_2282 (O_2282,N_16451,N_19282);
xnor UO_2283 (O_2283,N_17537,N_18502);
nand UO_2284 (O_2284,N_15274,N_19576);
and UO_2285 (O_2285,N_19108,N_16024);
xnor UO_2286 (O_2286,N_17892,N_15293);
and UO_2287 (O_2287,N_19056,N_17159);
or UO_2288 (O_2288,N_19720,N_16544);
nor UO_2289 (O_2289,N_17227,N_19445);
or UO_2290 (O_2290,N_19319,N_17862);
nor UO_2291 (O_2291,N_15823,N_19741);
nand UO_2292 (O_2292,N_19238,N_15581);
or UO_2293 (O_2293,N_19094,N_15155);
xnor UO_2294 (O_2294,N_15675,N_17453);
nor UO_2295 (O_2295,N_16070,N_19838);
and UO_2296 (O_2296,N_16603,N_17935);
nand UO_2297 (O_2297,N_19877,N_17744);
nand UO_2298 (O_2298,N_18920,N_16520);
and UO_2299 (O_2299,N_16873,N_15806);
and UO_2300 (O_2300,N_19597,N_15734);
or UO_2301 (O_2301,N_15834,N_19460);
xnor UO_2302 (O_2302,N_15219,N_19100);
or UO_2303 (O_2303,N_17972,N_15578);
and UO_2304 (O_2304,N_16368,N_18393);
and UO_2305 (O_2305,N_15399,N_19533);
nor UO_2306 (O_2306,N_18962,N_16486);
nand UO_2307 (O_2307,N_16015,N_19247);
or UO_2308 (O_2308,N_15132,N_16968);
xor UO_2309 (O_2309,N_17974,N_19085);
nor UO_2310 (O_2310,N_15465,N_17051);
xor UO_2311 (O_2311,N_15880,N_16285);
nor UO_2312 (O_2312,N_18309,N_15291);
xor UO_2313 (O_2313,N_17728,N_19906);
nor UO_2314 (O_2314,N_16986,N_18185);
and UO_2315 (O_2315,N_19443,N_18204);
and UO_2316 (O_2316,N_18846,N_18491);
and UO_2317 (O_2317,N_16713,N_15755);
and UO_2318 (O_2318,N_19433,N_15394);
nand UO_2319 (O_2319,N_16835,N_18953);
nor UO_2320 (O_2320,N_15273,N_19647);
nor UO_2321 (O_2321,N_16471,N_19957);
xor UO_2322 (O_2322,N_18215,N_17043);
or UO_2323 (O_2323,N_17331,N_17301);
xor UO_2324 (O_2324,N_16496,N_18690);
or UO_2325 (O_2325,N_16503,N_19830);
nor UO_2326 (O_2326,N_19506,N_18997);
or UO_2327 (O_2327,N_19764,N_18845);
and UO_2328 (O_2328,N_19937,N_17134);
nor UO_2329 (O_2329,N_19054,N_19736);
and UO_2330 (O_2330,N_19426,N_17427);
and UO_2331 (O_2331,N_19320,N_16816);
or UO_2332 (O_2332,N_18217,N_19801);
or UO_2333 (O_2333,N_19557,N_18969);
xnor UO_2334 (O_2334,N_15043,N_18879);
nand UO_2335 (O_2335,N_16017,N_18129);
or UO_2336 (O_2336,N_18470,N_16435);
nor UO_2337 (O_2337,N_18473,N_16045);
nor UO_2338 (O_2338,N_15503,N_17409);
nand UO_2339 (O_2339,N_19414,N_19731);
nand UO_2340 (O_2340,N_18387,N_16139);
or UO_2341 (O_2341,N_18852,N_15335);
nor UO_2342 (O_2342,N_15475,N_17133);
or UO_2343 (O_2343,N_18961,N_15982);
nand UO_2344 (O_2344,N_15423,N_19578);
nand UO_2345 (O_2345,N_18271,N_15442);
and UO_2346 (O_2346,N_17624,N_16150);
xnor UO_2347 (O_2347,N_19849,N_16809);
xnor UO_2348 (O_2348,N_18989,N_17949);
nor UO_2349 (O_2349,N_15552,N_17924);
nor UO_2350 (O_2350,N_15201,N_17895);
or UO_2351 (O_2351,N_17672,N_15267);
and UO_2352 (O_2352,N_16439,N_17479);
xnor UO_2353 (O_2353,N_18274,N_17613);
xor UO_2354 (O_2354,N_15867,N_17858);
nor UO_2355 (O_2355,N_19150,N_17088);
nor UO_2356 (O_2356,N_16052,N_17590);
nor UO_2357 (O_2357,N_18718,N_17729);
nor UO_2358 (O_2358,N_17721,N_15121);
and UO_2359 (O_2359,N_19086,N_18755);
xor UO_2360 (O_2360,N_16336,N_18343);
xnor UO_2361 (O_2361,N_15563,N_19931);
and UO_2362 (O_2362,N_18165,N_17716);
or UO_2363 (O_2363,N_19677,N_16461);
and UO_2364 (O_2364,N_15472,N_17848);
nand UO_2365 (O_2365,N_15580,N_18242);
xor UO_2366 (O_2366,N_19907,N_16315);
and UO_2367 (O_2367,N_19251,N_17840);
and UO_2368 (O_2368,N_17416,N_19780);
or UO_2369 (O_2369,N_17299,N_17640);
or UO_2370 (O_2370,N_19098,N_18900);
or UO_2371 (O_2371,N_15958,N_17307);
nor UO_2372 (O_2372,N_18566,N_18012);
nor UO_2373 (O_2373,N_17820,N_18600);
and UO_2374 (O_2374,N_19689,N_15220);
nand UO_2375 (O_2375,N_18696,N_15493);
and UO_2376 (O_2376,N_17871,N_15731);
nand UO_2377 (O_2377,N_18753,N_18208);
and UO_2378 (O_2378,N_15040,N_15191);
and UO_2379 (O_2379,N_16488,N_16845);
xnor UO_2380 (O_2380,N_18269,N_17095);
or UO_2381 (O_2381,N_17215,N_15872);
nor UO_2382 (O_2382,N_18455,N_15611);
xnor UO_2383 (O_2383,N_15826,N_16959);
xnor UO_2384 (O_2384,N_19730,N_18701);
xor UO_2385 (O_2385,N_17641,N_19512);
xor UO_2386 (O_2386,N_19208,N_17538);
nor UO_2387 (O_2387,N_16192,N_17700);
nor UO_2388 (O_2388,N_16297,N_18539);
nand UO_2389 (O_2389,N_15502,N_17278);
nor UO_2390 (O_2390,N_18632,N_15536);
nand UO_2391 (O_2391,N_16830,N_18593);
or UO_2392 (O_2392,N_15747,N_16001);
nand UO_2393 (O_2393,N_17082,N_19682);
or UO_2394 (O_2394,N_15500,N_19544);
nand UO_2395 (O_2395,N_16620,N_15822);
and UO_2396 (O_2396,N_16996,N_17710);
or UO_2397 (O_2397,N_19847,N_16764);
nor UO_2398 (O_2398,N_15729,N_19214);
and UO_2399 (O_2399,N_17799,N_17561);
xnor UO_2400 (O_2400,N_18643,N_18922);
nand UO_2401 (O_2401,N_15714,N_17911);
and UO_2402 (O_2402,N_19116,N_15263);
xnor UO_2403 (O_2403,N_18392,N_19210);
and UO_2404 (O_2404,N_15444,N_15835);
xnor UO_2405 (O_2405,N_19992,N_17329);
nor UO_2406 (O_2406,N_19290,N_17251);
or UO_2407 (O_2407,N_19361,N_17055);
or UO_2408 (O_2408,N_16994,N_17495);
nor UO_2409 (O_2409,N_18155,N_18827);
xnor UO_2410 (O_2410,N_17150,N_19311);
or UO_2411 (O_2411,N_17702,N_19126);
or UO_2412 (O_2412,N_19541,N_18435);
xnor UO_2413 (O_2413,N_15520,N_17988);
nand UO_2414 (O_2414,N_16623,N_18059);
xor UO_2415 (O_2415,N_17252,N_17921);
xnor UO_2416 (O_2416,N_19903,N_16571);
nand UO_2417 (O_2417,N_16926,N_18075);
nor UO_2418 (O_2418,N_17200,N_17163);
nor UO_2419 (O_2419,N_19692,N_19350);
nor UO_2420 (O_2420,N_19740,N_18973);
or UO_2421 (O_2421,N_17750,N_18721);
nor UO_2422 (O_2422,N_16849,N_18609);
or UO_2423 (O_2423,N_19676,N_19540);
nor UO_2424 (O_2424,N_15190,N_15975);
or UO_2425 (O_2425,N_16222,N_17255);
nand UO_2426 (O_2426,N_16258,N_15627);
or UO_2427 (O_2427,N_17543,N_18001);
nor UO_2428 (O_2428,N_17328,N_19322);
xnor UO_2429 (O_2429,N_15863,N_17363);
nor UO_2430 (O_2430,N_19791,N_18872);
nor UO_2431 (O_2431,N_15405,N_15609);
and UO_2432 (O_2432,N_15183,N_19518);
nand UO_2433 (O_2433,N_17297,N_15418);
nand UO_2434 (O_2434,N_19072,N_18510);
xnor UO_2435 (O_2435,N_17898,N_16594);
nand UO_2436 (O_2436,N_16626,N_16099);
xor UO_2437 (O_2437,N_17813,N_16993);
nand UO_2438 (O_2438,N_15746,N_17990);
nor UO_2439 (O_2439,N_15770,N_16814);
nor UO_2440 (O_2440,N_18607,N_17185);
nor UO_2441 (O_2441,N_19170,N_18719);
nor UO_2442 (O_2442,N_19222,N_19988);
or UO_2443 (O_2443,N_19500,N_16532);
and UO_2444 (O_2444,N_16616,N_17193);
and UO_2445 (O_2445,N_17569,N_19826);
xor UO_2446 (O_2446,N_19629,N_17598);
or UO_2447 (O_2447,N_15286,N_16374);
or UO_2448 (O_2448,N_16822,N_17635);
nand UO_2449 (O_2449,N_18825,N_19084);
nor UO_2450 (O_2450,N_15689,N_18143);
xor UO_2451 (O_2451,N_17320,N_15841);
nor UO_2452 (O_2452,N_17811,N_15717);
or UO_2453 (O_2453,N_15162,N_15065);
nor UO_2454 (O_2454,N_19456,N_19704);
and UO_2455 (O_2455,N_15892,N_17485);
xnor UO_2456 (O_2456,N_16466,N_19090);
and UO_2457 (O_2457,N_17290,N_16836);
and UO_2458 (O_2458,N_17351,N_15218);
nand UO_2459 (O_2459,N_16948,N_17006);
nor UO_2460 (O_2460,N_19379,N_18093);
nand UO_2461 (O_2461,N_16009,N_15665);
and UO_2462 (O_2462,N_16259,N_18213);
or UO_2463 (O_2463,N_17548,N_16226);
or UO_2464 (O_2464,N_18254,N_19983);
or UO_2465 (O_2465,N_15644,N_19258);
xnor UO_2466 (O_2466,N_19598,N_18168);
nand UO_2467 (O_2467,N_17582,N_15028);
xor UO_2468 (O_2468,N_16871,N_15437);
or UO_2469 (O_2469,N_16306,N_19887);
or UO_2470 (O_2470,N_17765,N_16758);
xnor UO_2471 (O_2471,N_19974,N_19884);
nand UO_2472 (O_2472,N_17634,N_19146);
and UO_2473 (O_2473,N_15733,N_17047);
nand UO_2474 (O_2474,N_16122,N_16580);
xor UO_2475 (O_2475,N_19067,N_16105);
and UO_2476 (O_2476,N_16943,N_18407);
and UO_2477 (O_2477,N_17284,N_18356);
nand UO_2478 (O_2478,N_16590,N_19652);
nand UO_2479 (O_2479,N_19968,N_15682);
nand UO_2480 (O_2480,N_18693,N_16810);
or UO_2481 (O_2481,N_18931,N_17411);
nor UO_2482 (O_2482,N_15600,N_16853);
nand UO_2483 (O_2483,N_18295,N_15889);
and UO_2484 (O_2484,N_19904,N_15805);
nor UO_2485 (O_2485,N_17381,N_18990);
nand UO_2486 (O_2486,N_17247,N_19382);
nand UO_2487 (O_2487,N_17771,N_17697);
nand UO_2488 (O_2488,N_17371,N_18895);
or UO_2489 (O_2489,N_16953,N_15786);
and UO_2490 (O_2490,N_17579,N_15793);
nand UO_2491 (O_2491,N_16013,N_15462);
and UO_2492 (O_2492,N_17162,N_19227);
and UO_2493 (O_2493,N_17010,N_16255);
nor UO_2494 (O_2494,N_17669,N_16007);
nor UO_2495 (O_2495,N_17759,N_17072);
and UO_2496 (O_2496,N_19480,N_19110);
nor UO_2497 (O_2497,N_18617,N_19003);
and UO_2498 (O_2498,N_19501,N_19602);
nor UO_2499 (O_2499,N_18272,N_17966);
endmodule