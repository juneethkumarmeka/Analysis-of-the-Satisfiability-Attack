module basic_1500_15000_2000_30_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xnor U0 (N_0,In_418,In_1495);
nor U1 (N_1,In_1387,In_605);
or U2 (N_2,In_987,In_1084);
nand U3 (N_3,In_566,In_1176);
xnor U4 (N_4,In_792,In_247);
xnor U5 (N_5,In_230,In_635);
xor U6 (N_6,In_306,In_30);
xor U7 (N_7,In_406,In_1494);
or U8 (N_8,In_165,In_1185);
xnor U9 (N_9,In_217,In_1386);
or U10 (N_10,In_1160,In_424);
and U11 (N_11,In_385,In_1313);
or U12 (N_12,In_696,In_262);
nor U13 (N_13,In_117,In_768);
and U14 (N_14,In_494,In_1461);
or U15 (N_15,In_1279,In_1326);
xnor U16 (N_16,In_4,In_807);
xnor U17 (N_17,In_1329,In_958);
xnor U18 (N_18,In_878,In_622);
or U19 (N_19,In_1257,In_1009);
nor U20 (N_20,In_1147,In_389);
or U21 (N_21,In_382,In_826);
and U22 (N_22,In_911,In_121);
and U23 (N_23,In_1366,In_320);
nand U24 (N_24,In_1002,In_741);
or U25 (N_25,In_1209,In_81);
and U26 (N_26,In_1324,In_1454);
or U27 (N_27,In_1229,In_162);
nor U28 (N_28,In_840,In_334);
and U29 (N_29,In_1096,In_575);
and U30 (N_30,In_538,In_1402);
xnor U31 (N_31,In_962,In_920);
and U32 (N_32,In_875,In_1303);
or U33 (N_33,In_539,In_1050);
xor U34 (N_34,In_409,In_1021);
nor U35 (N_35,In_1417,In_1424);
nand U36 (N_36,In_791,In_435);
xnor U37 (N_37,In_747,In_816);
or U38 (N_38,In_1478,In_1413);
and U39 (N_39,In_1211,In_1379);
and U40 (N_40,In_500,In_1374);
or U41 (N_41,In_924,In_432);
nor U42 (N_42,In_3,In_785);
nor U43 (N_43,In_896,In_993);
or U44 (N_44,In_1441,In_227);
and U45 (N_45,In_940,In_1108);
nand U46 (N_46,In_110,In_443);
nor U47 (N_47,In_1213,In_813);
nor U48 (N_48,In_1104,In_65);
and U49 (N_49,In_136,In_748);
nand U50 (N_50,In_482,In_877);
nand U51 (N_51,In_1281,In_1252);
nor U52 (N_52,In_34,In_862);
nand U53 (N_53,In_1051,In_508);
nand U54 (N_54,In_995,In_914);
or U55 (N_55,In_98,In_808);
xnor U56 (N_56,In_810,In_1450);
nor U57 (N_57,In_362,In_664);
xnor U58 (N_58,In_327,In_207);
or U59 (N_59,In_451,In_304);
and U60 (N_60,In_1451,In_905);
nand U61 (N_61,In_388,In_1492);
xnor U62 (N_62,In_1129,In_1218);
xnor U63 (N_63,In_574,In_111);
nand U64 (N_64,In_44,In_1354);
or U65 (N_65,In_883,In_867);
and U66 (N_66,In_767,In_1106);
nand U67 (N_67,In_673,In_314);
nand U68 (N_68,In_1091,In_787);
nand U69 (N_69,In_533,In_233);
nor U70 (N_70,In_75,In_1190);
xnor U71 (N_71,In_1238,In_194);
and U72 (N_72,In_977,In_51);
xnor U73 (N_73,In_1166,In_448);
nand U74 (N_74,In_980,In_1119);
xor U75 (N_75,In_1315,In_704);
and U76 (N_76,In_1156,In_1223);
nor U77 (N_77,In_737,In_1275);
or U78 (N_78,In_1282,In_1003);
or U79 (N_79,In_967,In_5);
nand U80 (N_80,In_1477,In_359);
or U81 (N_81,In_373,In_293);
and U82 (N_82,In_880,In_687);
xnor U83 (N_83,In_559,In_232);
nor U84 (N_84,In_1433,In_377);
and U85 (N_85,In_665,In_1423);
xor U86 (N_86,In_918,In_1369);
and U87 (N_87,In_209,In_534);
or U88 (N_88,In_28,In_1428);
or U89 (N_89,In_1042,In_1037);
nand U90 (N_90,In_1469,In_490);
or U91 (N_91,In_70,In_1388);
xnor U92 (N_92,In_321,In_229);
xor U93 (N_93,In_954,In_512);
nor U94 (N_94,In_922,In_1353);
nand U95 (N_95,In_436,In_268);
and U96 (N_96,In_1311,In_547);
xnor U97 (N_97,In_108,In_1270);
and U98 (N_98,In_771,In_1491);
nand U99 (N_99,In_403,In_295);
and U100 (N_100,In_433,In_1352);
nor U101 (N_101,In_367,In_1340);
and U102 (N_102,In_356,In_1309);
nor U103 (N_103,In_583,In_953);
xnor U104 (N_104,In_1331,In_35);
and U105 (N_105,In_908,In_511);
nor U106 (N_106,In_568,In_560);
nor U107 (N_107,In_1253,In_438);
or U108 (N_108,In_659,In_838);
nor U109 (N_109,In_931,In_1343);
nand U110 (N_110,In_1112,In_1310);
nand U111 (N_111,In_1152,In_1400);
or U112 (N_112,In_469,In_1090);
xnor U113 (N_113,In_1382,In_796);
xor U114 (N_114,In_1248,In_671);
xor U115 (N_115,In_1196,In_1116);
nand U116 (N_116,In_139,In_899);
xnor U117 (N_117,In_928,In_604);
xnor U118 (N_118,In_729,In_856);
xnor U119 (N_119,In_1154,In_1010);
or U120 (N_120,In_509,In_1406);
or U121 (N_121,In_1101,In_173);
xor U122 (N_122,In_542,In_532);
or U123 (N_123,In_1027,In_910);
and U124 (N_124,In_1055,In_739);
or U125 (N_125,In_750,In_20);
or U126 (N_126,In_379,In_755);
nor U127 (N_127,In_1225,In_1466);
nand U128 (N_128,In_290,In_156);
and U129 (N_129,In_322,In_1484);
nand U130 (N_130,In_812,In_161);
nand U131 (N_131,In_530,In_917);
nor U132 (N_132,In_1173,In_1134);
nor U133 (N_133,In_1345,In_346);
and U134 (N_134,In_1066,In_834);
or U135 (N_135,In_240,In_393);
or U136 (N_136,In_541,In_1078);
and U137 (N_137,In_1180,In_468);
nand U138 (N_138,In_986,In_292);
or U139 (N_139,In_841,In_853);
or U140 (N_140,In_636,In_1498);
xor U141 (N_141,In_1452,In_109);
xnor U142 (N_142,In_1422,In_397);
and U143 (N_143,In_1170,In_46);
nor U144 (N_144,In_624,In_378);
and U145 (N_145,In_545,In_666);
nand U146 (N_146,In_1483,In_42);
nand U147 (N_147,In_573,In_514);
nor U148 (N_148,In_186,In_572);
nor U149 (N_149,In_90,In_855);
nor U150 (N_150,In_582,In_383);
nand U151 (N_151,In_353,In_1140);
nor U152 (N_152,In_129,In_844);
and U153 (N_153,In_594,In_523);
nand U154 (N_154,In_1219,In_657);
or U155 (N_155,In_1305,In_72);
nand U156 (N_156,In_447,In_1363);
nor U157 (N_157,In_502,In_239);
xor U158 (N_158,In_1316,In_1202);
xor U159 (N_159,In_1060,In_1321);
nand U160 (N_160,In_1032,In_1086);
and U161 (N_161,In_47,In_159);
xnor U162 (N_162,In_219,In_1039);
or U163 (N_163,In_31,In_215);
or U164 (N_164,In_256,In_1377);
nand U165 (N_165,In_115,In_53);
nand U166 (N_166,In_332,In_688);
nor U167 (N_167,In_872,In_1485);
xor U168 (N_168,In_1040,In_658);
nand U169 (N_169,In_1464,In_780);
nor U170 (N_170,In_835,In_350);
or U171 (N_171,In_93,In_1144);
or U172 (N_172,In_39,In_630);
and U173 (N_173,In_43,In_416);
nand U174 (N_174,In_1214,In_1);
nor U175 (N_175,In_1193,In_479);
xor U176 (N_176,In_1067,In_309);
nand U177 (N_177,In_176,In_1189);
nor U178 (N_178,In_1221,In_260);
nor U179 (N_179,In_1399,In_1022);
nor U180 (N_180,In_374,In_1472);
or U181 (N_181,In_596,In_331);
or U182 (N_182,In_354,In_312);
nor U183 (N_183,In_1023,In_1094);
xor U184 (N_184,In_943,In_372);
xnor U185 (N_185,In_158,In_59);
and U186 (N_186,In_1325,In_626);
xor U187 (N_187,In_287,In_86);
nand U188 (N_188,In_1224,In_777);
xnor U189 (N_189,In_618,In_839);
and U190 (N_190,In_628,In_632);
and U191 (N_191,In_722,In_776);
and U192 (N_192,In_22,In_930);
nor U193 (N_193,In_452,In_1162);
xnor U194 (N_194,In_932,In_307);
nand U195 (N_195,In_1421,In_1163);
and U196 (N_196,In_1474,In_646);
and U197 (N_197,In_1332,In_198);
nand U198 (N_198,In_781,In_773);
nor U199 (N_199,In_836,In_1085);
or U200 (N_200,In_728,In_1007);
xor U201 (N_201,In_806,In_1459);
xnor U202 (N_202,In_553,In_1103);
or U203 (N_203,In_692,In_1360);
and U204 (N_204,In_540,In_990);
or U205 (N_205,In_315,In_302);
nand U206 (N_206,In_764,In_1470);
xnor U207 (N_207,In_801,In_455);
nand U208 (N_208,In_2,In_1264);
or U209 (N_209,In_351,In_1235);
or U210 (N_210,In_927,In_818);
or U211 (N_211,In_689,In_339);
nand U212 (N_212,In_276,In_1008);
xor U213 (N_213,In_711,In_137);
nor U214 (N_214,In_1114,In_1174);
nand U215 (N_215,In_874,In_184);
or U216 (N_216,In_425,In_846);
nand U217 (N_217,In_654,In_49);
xnor U218 (N_218,In_495,In_994);
xnor U219 (N_219,In_484,In_513);
nand U220 (N_220,In_685,In_141);
and U221 (N_221,In_651,In_1398);
or U222 (N_222,In_555,In_399);
nor U223 (N_223,In_1337,In_525);
nor U224 (N_224,In_1390,In_1043);
xor U225 (N_225,In_1208,In_99);
xnor U226 (N_226,In_1287,In_992);
nand U227 (N_227,In_1053,In_1294);
xor U228 (N_228,In_714,In_167);
or U229 (N_229,In_890,In_1304);
nor U230 (N_230,In_316,In_69);
xnor U231 (N_231,In_820,In_178);
or U232 (N_232,In_1151,In_1299);
nand U233 (N_233,In_611,In_253);
or U234 (N_234,In_1327,In_480);
xor U235 (N_235,In_355,In_644);
and U236 (N_236,In_613,In_193);
or U237 (N_237,In_1188,In_580);
nor U238 (N_238,In_1099,In_675);
nand U239 (N_239,In_516,In_446);
nand U240 (N_240,In_570,In_1442);
and U241 (N_241,In_631,In_1240);
or U242 (N_242,In_1014,In_213);
and U243 (N_243,In_1026,In_978);
nor U244 (N_244,In_832,In_1284);
and U245 (N_245,In_338,In_1195);
nand U246 (N_246,In_1271,In_882);
nor U247 (N_247,In_865,In_1395);
xor U248 (N_248,In_984,In_133);
and U249 (N_249,In_981,In_454);
nand U250 (N_250,In_1100,In_1490);
or U251 (N_251,In_745,In_705);
and U252 (N_252,In_847,In_1226);
nand U253 (N_253,In_422,In_629);
nand U254 (N_254,In_721,In_788);
or U255 (N_255,In_916,In_888);
nand U256 (N_256,In_677,In_674);
or U257 (N_257,In_172,In_437);
xnor U258 (N_258,In_868,In_243);
and U259 (N_259,In_182,In_32);
nor U260 (N_260,In_261,In_458);
or U261 (N_261,In_1447,In_933);
nor U262 (N_262,In_171,In_1348);
nor U263 (N_263,In_1231,In_1045);
xnor U264 (N_264,In_1404,In_1462);
nand U265 (N_265,In_1121,In_1164);
nand U266 (N_266,In_1093,In_274);
and U267 (N_267,In_58,In_491);
nand U268 (N_268,In_799,In_515);
and U269 (N_269,In_174,In_1089);
nor U270 (N_270,In_348,In_1247);
xnor U271 (N_271,In_778,In_441);
nor U272 (N_272,In_627,In_301);
nand U273 (N_273,In_380,In_770);
xnor U274 (N_274,In_474,In_1035);
or U275 (N_275,In_1475,In_1342);
nand U276 (N_276,In_1250,In_623);
or U277 (N_277,In_333,In_848);
or U278 (N_278,In_858,In_752);
or U279 (N_279,In_1128,In_1307);
or U280 (N_280,In_1471,In_1254);
xnor U281 (N_281,In_54,In_1286);
nor U282 (N_282,In_585,In_38);
xor U283 (N_283,In_279,In_597);
nand U284 (N_284,In_1361,In_466);
xnor U285 (N_285,In_57,In_886);
and U286 (N_286,In_1298,In_1088);
or U287 (N_287,In_794,In_36);
nor U288 (N_288,In_1041,In_386);
xor U289 (N_289,In_563,In_1130);
or U290 (N_290,In_1083,In_548);
and U291 (N_291,In_531,In_1308);
nand U292 (N_292,In_1277,In_617);
and U293 (N_293,In_445,In_1206);
nor U294 (N_294,In_470,In_1172);
nand U295 (N_295,In_1062,In_1312);
xor U296 (N_296,In_1443,In_970);
xor U297 (N_297,In_13,In_395);
nand U298 (N_298,In_979,In_985);
nor U299 (N_299,In_588,In_1239);
or U300 (N_300,In_518,In_119);
nand U301 (N_301,In_400,In_77);
or U302 (N_302,In_1059,In_786);
and U303 (N_303,In_947,In_569);
and U304 (N_304,In_1110,In_1444);
xnor U305 (N_305,In_1124,In_1065);
xnor U306 (N_306,In_1434,In_486);
and U307 (N_307,In_100,In_889);
nand U308 (N_308,In_1052,In_1063);
nand U309 (N_309,In_189,In_138);
nor U310 (N_310,In_343,In_414);
or U311 (N_311,In_740,In_676);
xnor U312 (N_312,In_1259,In_122);
xnor U313 (N_313,In_699,In_619);
nand U314 (N_314,In_701,In_1155);
and U315 (N_315,In_1350,In_1159);
or U316 (N_316,In_906,In_505);
nand U317 (N_317,In_11,In_64);
nand U318 (N_318,In_344,In_29);
or U319 (N_319,In_96,In_1457);
xnor U320 (N_320,In_811,In_706);
xnor U321 (N_321,In_303,In_358);
nor U322 (N_322,In_1030,In_702);
and U323 (N_323,In_814,In_423);
or U324 (N_324,In_1412,In_1430);
and U325 (N_325,In_74,In_1216);
xor U326 (N_326,In_1427,In_1126);
nor U327 (N_327,In_12,In_146);
xor U328 (N_328,In_459,In_370);
and U329 (N_329,In_413,In_1161);
nand U330 (N_330,In_761,In_1105);
nand U331 (N_331,In_703,In_1047);
nand U332 (N_332,In_203,In_444);
or U333 (N_333,In_1455,In_1048);
and U334 (N_334,In_528,In_1426);
xnor U335 (N_335,In_1463,In_427);
or U336 (N_336,In_913,In_123);
and U337 (N_337,In_997,In_625);
nand U338 (N_338,In_960,In_242);
xnor U339 (N_339,In_881,In_1033);
xor U340 (N_340,In_1397,In_113);
nor U341 (N_341,In_550,In_1482);
xor U342 (N_342,In_145,In_396);
and U343 (N_343,In_250,In_1258);
or U344 (N_344,In_1265,In_163);
nor U345 (N_345,In_349,In_1031);
or U346 (N_346,In_285,In_1356);
nand U347 (N_347,In_1073,In_61);
nor U348 (N_348,In_1346,In_255);
and U349 (N_349,In_45,In_536);
and U350 (N_350,In_510,In_328);
nor U351 (N_351,In_475,In_1192);
or U352 (N_352,In_252,In_1168);
nor U353 (N_353,In_895,In_340);
or U354 (N_354,In_1291,In_1292);
xnor U355 (N_355,In_1107,In_754);
xor U356 (N_356,In_1013,In_1232);
nand U357 (N_357,In_601,In_1347);
nor U358 (N_358,In_1237,In_465);
nor U359 (N_359,In_873,In_843);
nand U360 (N_360,In_1302,In_254);
nor U361 (N_361,In_376,In_937);
nor U362 (N_362,In_185,In_234);
nand U363 (N_363,In_1488,In_949);
nand U364 (N_364,In_1001,In_713);
and U365 (N_365,In_1285,In_1446);
nand U366 (N_366,In_420,In_214);
xor U367 (N_367,In_892,In_825);
nor U368 (N_368,In_1288,In_1210);
xor U369 (N_369,In_743,In_1025);
nor U370 (N_370,In_154,In_957);
and U371 (N_371,In_744,In_151);
and U372 (N_372,In_576,In_1380);
xnor U373 (N_373,In_1336,In_206);
or U374 (N_374,In_488,In_827);
nand U375 (N_375,In_700,In_1268);
nor U376 (N_376,In_1137,In_1038);
or U377 (N_377,In_246,In_37);
xor U378 (N_378,In_948,In_817);
nand U379 (N_379,In_524,In_612);
nor U380 (N_380,In_211,In_639);
xnor U381 (N_381,In_736,In_589);
xor U382 (N_382,In_996,In_181);
xnor U383 (N_383,In_1165,In_1297);
xnor U384 (N_384,In_270,In_439);
or U385 (N_385,In_945,In_128);
nand U386 (N_386,In_1368,In_1143);
and U387 (N_387,In_1314,In_1330);
and U388 (N_388,In_595,In_352);
nand U389 (N_389,In_134,In_652);
xnor U390 (N_390,In_118,In_879);
nor U391 (N_391,In_600,In_105);
nor U392 (N_392,In_415,In_294);
or U393 (N_393,In_1317,In_772);
nor U394 (N_394,In_650,In_160);
and U395 (N_395,In_802,In_222);
nor U396 (N_396,In_1068,In_989);
xor U397 (N_397,In_80,In_1389);
or U398 (N_398,In_1373,In_1006);
xor U399 (N_399,In_564,In_691);
xor U400 (N_400,In_670,In_935);
nand U401 (N_401,In_1004,In_106);
nand U402 (N_402,In_140,In_1328);
and U403 (N_403,In_763,In_1000);
and U404 (N_404,In_697,In_1236);
nand U405 (N_405,In_976,In_830);
and U406 (N_406,In_815,In_602);
xnor U407 (N_407,In_912,In_790);
nor U408 (N_408,In_24,In_387);
nor U409 (N_409,In_730,In_1344);
and U410 (N_410,In_599,In_135);
or U411 (N_411,In_503,In_567);
and U412 (N_412,In_1245,In_1425);
nand U413 (N_413,In_963,In_237);
nand U414 (N_414,In_1132,In_1102);
nand U415 (N_415,In_384,In_633);
xor U416 (N_416,In_296,In_166);
xor U417 (N_417,In_708,In_1355);
nor U418 (N_418,In_831,In_1179);
or U419 (N_419,In_537,In_1175);
nor U420 (N_420,In_342,In_824);
nor U421 (N_421,In_760,In_1109);
and U422 (N_422,In_690,In_769);
or U423 (N_423,In_766,In_1320);
and U424 (N_424,In_265,In_891);
or U425 (N_425,In_212,In_190);
and U426 (N_426,In_324,In_381);
and U427 (N_427,In_762,In_197);
nand U428 (N_428,In_800,In_21);
nor U429 (N_429,In_1489,In_734);
nor U430 (N_430,In_1295,In_919);
xnor U431 (N_431,In_551,In_62);
nand U432 (N_432,In_1234,In_968);
and U433 (N_433,In_955,In_1016);
or U434 (N_434,In_1394,In_1028);
or U435 (N_435,In_1197,In_249);
nand U436 (N_436,In_392,In_1158);
xnor U437 (N_437,In_477,In_749);
xor U438 (N_438,In_609,In_608);
nor U439 (N_439,In_73,In_1269);
or U440 (N_440,In_394,In_757);
and U441 (N_441,In_1411,In_404);
nand U442 (N_442,In_1449,In_586);
or U443 (N_443,In_854,In_1097);
nor U444 (N_444,In_1177,In_91);
xnor U445 (N_445,In_823,In_876);
or U446 (N_446,In_89,In_526);
and U447 (N_447,In_1203,In_1181);
or U448 (N_448,In_1212,In_1015);
nand U449 (N_449,In_485,In_1333);
nor U450 (N_450,In_1157,In_578);
nor U451 (N_451,In_988,In_1359);
nor U452 (N_452,In_1499,In_467);
or U453 (N_453,In_201,In_756);
or U454 (N_454,In_1262,In_695);
nand U455 (N_455,In_647,In_263);
nand U456 (N_456,In_923,In_1391);
nor U457 (N_457,In_1241,In_10);
or U458 (N_458,In_504,In_668);
xor U459 (N_459,In_637,In_126);
nand U460 (N_460,In_308,In_92);
or U461 (N_461,In_869,In_456);
nand U462 (N_462,In_860,In_614);
or U463 (N_463,In_300,In_842);
and U464 (N_464,In_733,In_1044);
or U465 (N_465,In_6,In_731);
xor U466 (N_466,In_1358,In_1448);
nor U467 (N_467,In_152,In_598);
nand U468 (N_468,In_535,In_1420);
and U469 (N_469,In_492,In_1123);
xor U470 (N_470,In_1473,In_481);
and U471 (N_471,In_732,In_1242);
nand U472 (N_472,In_476,In_1408);
or U473 (N_473,In_707,In_1133);
nor U474 (N_474,In_549,In_775);
nor U475 (N_475,In_1149,In_774);
xor U476 (N_476,In_1187,In_643);
xnor U477 (N_477,In_1334,In_1362);
nor U478 (N_478,In_669,In_1456);
xnor U479 (N_479,In_148,In_983);
nand U480 (N_480,In_257,In_871);
or U481 (N_481,In_421,In_1255);
or U482 (N_482,In_956,In_884);
or U483 (N_483,In_297,In_921);
nand U484 (N_484,In_1020,In_837);
xor U485 (N_485,In_1077,In_408);
nor U486 (N_486,In_584,In_236);
nor U487 (N_487,In_765,In_710);
and U488 (N_488,In_323,In_116);
and U489 (N_489,In_593,In_942);
xor U490 (N_490,In_1263,In_1364);
nor U491 (N_491,In_1409,In_202);
nor U492 (N_492,In_972,In_1115);
xor U493 (N_493,In_907,In_144);
nor U494 (N_494,In_1375,In_1465);
xor U495 (N_495,In_1293,In_241);
or U496 (N_496,In_822,In_1246);
nand U497 (N_497,In_1372,In_506);
or U498 (N_498,In_759,In_78);
or U499 (N_499,In_195,In_661);
and U500 (N_500,N_423,In_1403);
and U501 (N_501,N_481,N_74);
nand U502 (N_502,In_187,N_63);
or U503 (N_503,In_391,In_71);
or U504 (N_504,N_110,N_102);
nand U505 (N_505,In_944,N_419);
nand U506 (N_506,In_264,N_27);
nor U507 (N_507,In_196,N_60);
and U508 (N_508,N_208,N_100);
xor U509 (N_509,In_753,In_280);
nand U510 (N_510,In_1069,N_255);
or U511 (N_511,In_68,In_901);
nor U512 (N_512,In_1205,N_471);
nor U513 (N_513,In_587,In_335);
nor U514 (N_514,In_147,In_1410);
nand U515 (N_515,In_517,In_1487);
nor U516 (N_516,N_300,N_249);
xor U517 (N_517,In_1228,In_590);
xor U518 (N_518,In_366,N_80);
nand U519 (N_519,N_253,In_55);
and U520 (N_520,In_544,In_1251);
xnor U521 (N_521,N_496,In_63);
and U522 (N_522,In_678,In_1319);
nand U523 (N_523,In_371,In_804);
and U524 (N_524,N_393,N_85);
nor U525 (N_525,N_164,In_1061);
nor U526 (N_526,In_1445,In_803);
nand U527 (N_527,In_1335,In_951);
or U528 (N_528,N_205,N_143);
xor U529 (N_529,In_667,N_166);
and U530 (N_530,N_141,N_17);
nand U531 (N_531,In_417,N_95);
and U532 (N_532,In_859,N_397);
nor U533 (N_533,N_324,N_349);
or U534 (N_534,N_189,N_363);
and U535 (N_535,In_1056,N_429);
nand U536 (N_536,In_1057,N_308);
and U537 (N_537,In_709,N_207);
nand U538 (N_538,In_223,N_172);
and U539 (N_539,In_473,In_1049);
nand U540 (N_540,N_284,N_46);
and U541 (N_541,In_1092,N_402);
or U542 (N_542,N_92,In_337);
and U543 (N_543,N_335,In_7);
and U544 (N_544,In_607,In_1118);
nand U545 (N_545,N_354,N_332);
nand U546 (N_546,In_430,In_120);
xor U547 (N_547,In_199,In_15);
or U548 (N_548,In_925,N_64);
or U549 (N_549,In_798,In_1167);
xnor U550 (N_550,N_137,In_56);
and U551 (N_551,N_269,In_738);
and U552 (N_552,N_304,In_735);
nand U553 (N_553,In_1376,N_420);
or U554 (N_554,In_1436,In_961);
or U555 (N_555,N_438,N_279);
and U556 (N_556,In_489,N_190);
nand U557 (N_557,N_406,N_10);
nor U558 (N_558,In_1098,In_1186);
and U559 (N_559,In_718,N_366);
or U560 (N_560,N_453,N_61);
or U561 (N_561,In_902,N_182);
nor U562 (N_562,In_683,In_1249);
nand U563 (N_563,In_851,In_1468);
nand U564 (N_564,N_358,In_1435);
nor U565 (N_565,N_160,In_1381);
xor U566 (N_566,N_67,N_474);
nor U567 (N_567,In_149,In_499);
and U568 (N_568,In_929,N_458);
and U569 (N_569,N_243,In_210);
xor U570 (N_570,N_168,In_936);
nand U571 (N_571,In_1146,N_186);
xnor U572 (N_572,In_1183,In_224);
nor U573 (N_573,In_1351,In_1318);
xnor U574 (N_574,In_1029,N_370);
nor U575 (N_575,N_202,In_231);
or U576 (N_576,In_282,N_181);
and U577 (N_577,In_1017,In_169);
and U578 (N_578,In_175,In_833);
and U579 (N_579,N_56,In_464);
nand U580 (N_580,N_199,N_16);
nor U581 (N_581,N_380,In_431);
nand U582 (N_582,N_396,N_162);
and U583 (N_583,N_177,N_153);
and U584 (N_584,In_900,N_219);
or U585 (N_585,N_57,In_496);
or U586 (N_586,N_360,In_561);
and U587 (N_587,N_84,In_797);
nand U588 (N_588,In_1385,N_326);
or U589 (N_589,In_1138,N_30);
xnor U590 (N_590,N_22,In_375);
and U591 (N_591,In_426,N_359);
nor U592 (N_592,N_197,In_1497);
nor U593 (N_593,In_969,N_337);
and U594 (N_594,N_444,In_157);
xnor U595 (N_595,In_1079,In_1024);
nor U596 (N_596,N_464,In_226);
xnor U597 (N_597,In_318,N_422);
and U598 (N_598,In_410,N_55);
and U599 (N_599,N_302,N_105);
or U600 (N_600,In_894,N_131);
or U601 (N_601,N_480,N_367);
and U602 (N_602,In_76,N_231);
xnor U603 (N_603,In_789,In_758);
xor U604 (N_604,N_263,In_104);
nor U605 (N_605,N_355,N_62);
nor U606 (N_606,N_362,In_522);
and U607 (N_607,In_1034,N_407);
nand U608 (N_608,In_95,In_1125);
nand U609 (N_609,In_390,N_94);
nand U610 (N_610,In_1046,In_926);
xor U611 (N_611,N_493,In_1111);
nor U612 (N_612,In_663,In_861);
and U613 (N_613,N_456,In_245);
nand U614 (N_614,N_11,N_118);
and U615 (N_615,In_1439,In_67);
xnor U616 (N_616,In_982,N_233);
or U617 (N_617,N_436,In_1200);
or U618 (N_618,N_216,N_51);
xor U619 (N_619,N_434,In_720);
xnor U620 (N_620,N_313,In_606);
and U621 (N_621,N_303,In_850);
xor U622 (N_622,N_20,In_952);
nand U623 (N_623,In_974,N_482);
and U624 (N_624,N_491,In_1198);
and U625 (N_625,In_112,In_405);
xnor U626 (N_626,N_221,N_340);
xor U627 (N_627,N_203,In_571);
and U628 (N_628,In_716,In_401);
and U629 (N_629,N_364,In_472);
and U630 (N_630,In_153,N_490);
and U631 (N_631,In_497,N_239);
xnor U632 (N_632,N_375,N_169);
or U633 (N_633,In_897,N_476);
and U634 (N_634,In_1058,N_472);
and U635 (N_635,N_274,In_724);
nor U636 (N_636,In_793,In_603);
nand U637 (N_637,N_191,In_17);
xnor U638 (N_638,In_521,N_214);
xor U639 (N_639,In_281,N_33);
or U640 (N_640,In_784,In_529);
or U641 (N_641,In_562,N_385);
and U642 (N_642,In_218,In_1267);
and U643 (N_643,In_1012,N_247);
nand U644 (N_644,N_350,In_336);
nand U645 (N_645,N_250,N_45);
or U646 (N_646,In_552,In_1178);
or U647 (N_647,In_84,N_0);
xnor U648 (N_648,N_187,In_102);
or U649 (N_649,N_123,In_275);
or U650 (N_650,In_1323,N_399);
and U651 (N_651,In_1429,In_1064);
nand U652 (N_652,In_272,N_180);
nand U653 (N_653,In_471,In_330);
xnor U654 (N_654,In_107,N_310);
or U655 (N_655,N_37,N_414);
nor U656 (N_656,In_325,N_201);
nand U657 (N_657,In_1150,In_1215);
xnor U658 (N_658,N_365,N_449);
and U659 (N_659,N_14,N_122);
or U660 (N_660,In_681,N_416);
xnor U661 (N_661,N_451,In_640);
nand U662 (N_662,In_1171,N_212);
nor U663 (N_663,N_356,N_381);
nand U664 (N_664,In_819,In_319);
nand U665 (N_665,In_546,In_1306);
or U666 (N_666,In_1054,In_964);
xnor U667 (N_667,N_192,N_383);
and U668 (N_668,In_1357,In_188);
and U669 (N_669,N_28,In_428);
nand U670 (N_670,N_38,In_999);
and U671 (N_671,In_1407,N_394);
or U672 (N_672,N_138,In_1071);
xnor U673 (N_673,In_1438,In_579);
nand U674 (N_674,In_939,In_938);
and U675 (N_675,N_401,N_165);
xor U676 (N_676,N_489,N_116);
or U677 (N_677,In_8,N_264);
or U678 (N_678,N_13,N_254);
nor U679 (N_679,N_409,N_79);
nor U680 (N_680,N_1,N_232);
nand U681 (N_681,N_430,N_391);
xor U682 (N_682,In_25,In_1371);
or U683 (N_683,N_140,In_1437);
nand U684 (N_684,In_893,In_1182);
and U685 (N_685,N_159,N_178);
nor U686 (N_686,In_60,In_180);
xor U687 (N_687,N_48,N_344);
nor U688 (N_688,In_79,In_440);
xor U689 (N_689,N_150,In_1036);
xnor U690 (N_690,N_29,In_723);
nand U691 (N_691,In_909,N_148);
or U692 (N_692,In_341,N_227);
nor U693 (N_693,In_192,N_352);
or U694 (N_694,In_1070,In_291);
and U695 (N_695,N_196,N_188);
nor U696 (N_696,In_0,In_1396);
and U697 (N_697,In_183,N_135);
xor U698 (N_698,In_965,In_1383);
or U699 (N_699,In_719,In_1432);
or U700 (N_700,N_19,N_68);
nor U701 (N_701,N_157,N_54);
nand U702 (N_702,N_301,N_467);
or U703 (N_703,In_1074,N_432);
xor U704 (N_704,N_259,In_1220);
nand U705 (N_705,N_114,N_257);
and U706 (N_706,In_903,N_7);
nand U707 (N_707,N_70,N_147);
and U708 (N_708,N_377,N_320);
or U709 (N_709,N_44,N_183);
and U710 (N_710,N_328,N_107);
nand U711 (N_711,In_273,In_288);
nand U712 (N_712,In_1479,N_98);
nand U713 (N_713,N_75,In_672);
xor U714 (N_714,N_316,In_1272);
and U715 (N_715,N_455,In_179);
xnor U716 (N_716,N_58,N_198);
or U717 (N_717,N_241,N_31);
and U718 (N_718,N_53,N_106);
nand U719 (N_719,In_591,N_59);
nor U720 (N_720,N_446,N_440);
nor U721 (N_721,N_325,N_109);
and U722 (N_722,In_238,N_305);
nor U723 (N_723,N_111,N_224);
nor U724 (N_724,N_479,In_1266);
nor U725 (N_725,N_124,In_1486);
and U726 (N_726,In_648,N_431);
or U727 (N_727,N_357,N_194);
nor U728 (N_728,In_204,In_170);
and U729 (N_729,N_104,In_1260);
and U730 (N_730,N_39,N_195);
nor U731 (N_731,N_171,N_8);
and U732 (N_732,In_205,In_1191);
xnor U733 (N_733,In_368,N_336);
or U734 (N_734,N_353,In_1136);
or U735 (N_735,In_662,In_33);
nand U736 (N_736,In_1230,In_103);
nor U737 (N_737,N_272,In_1153);
nor U738 (N_738,N_285,In_26);
and U739 (N_739,In_277,In_40);
nand U740 (N_740,N_175,In_18);
nor U741 (N_741,N_3,N_132);
nand U742 (N_742,In_751,In_1290);
nand U743 (N_743,N_488,N_435);
nor U744 (N_744,N_266,N_345);
xnor U745 (N_745,In_1300,N_441);
nand U746 (N_746,N_234,N_379);
nor U747 (N_747,N_91,N_428);
nand U748 (N_748,In_870,In_660);
nor U749 (N_749,N_77,In_130);
and U750 (N_750,N_478,N_297);
xnor U751 (N_751,N_462,N_348);
xor U752 (N_752,In_1278,N_12);
nand U753 (N_753,In_150,In_1467);
nor U754 (N_754,In_363,N_41);
xor U755 (N_755,In_649,In_821);
xnor U756 (N_756,N_466,N_258);
and U757 (N_757,In_345,In_244);
or U758 (N_758,In_326,N_323);
xor U759 (N_759,N_475,In_934);
nor U760 (N_760,N_448,In_1139);
and U761 (N_761,In_317,N_477);
and U762 (N_762,In_1072,N_331);
nor U763 (N_763,N_69,In_1122);
xor U764 (N_764,N_442,In_191);
and U765 (N_765,N_82,In_398);
nor U766 (N_766,In_1405,N_412);
xor U767 (N_767,N_373,In_863);
and U768 (N_768,In_887,In_1243);
nor U769 (N_769,In_271,N_389);
or U770 (N_770,N_152,In_682);
nor U771 (N_771,N_204,N_282);
nor U772 (N_772,In_615,N_42);
and U773 (N_773,N_411,In_971);
xor U774 (N_774,In_1204,N_267);
nand U775 (N_775,In_305,In_463);
nor U776 (N_776,In_828,In_442);
nor U777 (N_777,In_1095,In_365);
and U778 (N_778,N_215,In_1365);
or U779 (N_779,N_170,N_314);
nand U780 (N_780,N_403,N_156);
and U781 (N_781,In_941,N_312);
nand U782 (N_782,N_400,N_83);
and U783 (N_783,In_1131,In_82);
or U784 (N_784,N_32,N_268);
and U785 (N_785,In_200,In_259);
and U786 (N_786,N_343,N_230);
or U787 (N_787,N_71,In_727);
xor U788 (N_788,N_483,N_463);
nor U789 (N_789,N_176,In_852);
and U790 (N_790,In_1082,In_1120);
nor U791 (N_791,N_261,In_1075);
and U792 (N_792,In_487,In_298);
xor U793 (N_793,N_387,N_73);
xnor U794 (N_794,In_898,N_315);
or U795 (N_795,N_418,N_103);
and U796 (N_796,In_1087,N_174);
or U797 (N_797,N_398,In_1256);
nor U798 (N_798,In_114,N_236);
and U799 (N_799,In_131,In_483);
or U800 (N_800,N_445,N_386);
nor U801 (N_801,In_97,In_1117);
nand U802 (N_802,N_142,N_473);
or U803 (N_803,In_23,In_1018);
and U804 (N_804,In_998,In_726);
nand U805 (N_805,N_220,N_86);
nand U806 (N_806,In_1416,In_866);
or U807 (N_807,In_124,N_498);
and U808 (N_808,N_361,In_556);
nand U809 (N_809,N_43,N_163);
or U810 (N_810,In_991,N_151);
xor U811 (N_811,In_680,N_161);
nand U812 (N_812,In_1019,In_1207);
and U813 (N_813,In_283,N_346);
and U814 (N_814,N_417,In_641);
nand U815 (N_815,In_1496,N_256);
and U816 (N_816,N_211,N_40);
nor U817 (N_817,N_283,N_72);
nand U818 (N_818,In_1480,N_287);
nand U819 (N_819,N_78,N_321);
and U820 (N_820,N_288,N_395);
nand U821 (N_821,N_134,In_1481);
nor U822 (N_822,In_783,In_27);
or U823 (N_823,N_213,N_155);
nand U824 (N_824,In_1460,In_1201);
nor U825 (N_825,In_1378,In_507);
xor U826 (N_826,In_1142,In_610);
and U827 (N_827,N_112,In_717);
nand U828 (N_828,N_465,In_216);
nand U829 (N_829,In_829,N_145);
nor U830 (N_830,N_497,N_52);
and U831 (N_831,In_310,N_468);
nor U832 (N_832,In_1113,In_357);
nor U833 (N_833,N_470,N_265);
xor U834 (N_834,In_16,In_1261);
nand U835 (N_835,In_554,N_88);
nor U836 (N_836,In_1274,N_244);
xor U837 (N_837,In_87,N_329);
or U838 (N_838,In_712,N_371);
or U839 (N_839,N_173,N_278);
and U840 (N_840,N_139,N_421);
xor U841 (N_841,N_65,In_1453);
or U842 (N_842,In_177,In_656);
nand U843 (N_843,In_1169,In_1401);
and U844 (N_844,N_494,In_299);
and U845 (N_845,In_845,In_693);
nand U846 (N_846,N_99,N_291);
xnor U847 (N_847,In_746,In_616);
nand U848 (N_848,N_119,N_499);
xnor U849 (N_849,In_1194,N_36);
nor U850 (N_850,N_390,N_115);
nor U851 (N_851,In_809,In_1141);
or U852 (N_852,N_5,N_90);
or U853 (N_853,N_81,N_484);
or U854 (N_854,N_18,N_382);
and U855 (N_855,In_402,N_342);
and U856 (N_856,N_469,In_450);
or U857 (N_857,N_130,In_1367);
or U858 (N_858,In_1392,N_225);
and U859 (N_859,In_1418,N_235);
nand U860 (N_860,N_295,In_411);
nand U861 (N_861,N_289,N_210);
xnor U862 (N_862,In_1415,N_281);
nor U863 (N_863,In_267,N_228);
nor U864 (N_864,In_85,N_218);
xor U865 (N_865,In_407,N_487);
nor U866 (N_866,In_565,N_76);
or U867 (N_867,N_369,In_1370);
nor U868 (N_868,In_125,N_6);
or U869 (N_869,In_501,In_251);
or U870 (N_870,N_9,In_684);
and U871 (N_871,In_142,N_306);
nand U872 (N_872,N_251,In_313);
or U873 (N_873,N_368,N_437);
nand U874 (N_874,In_258,N_299);
and U875 (N_875,In_1273,In_155);
or U876 (N_876,N_426,N_184);
nand U877 (N_877,N_273,N_454);
xor U878 (N_878,In_14,N_129);
or U879 (N_879,N_23,N_439);
or U880 (N_880,In_266,In_225);
and U881 (N_881,N_117,N_330);
nor U882 (N_882,In_1233,In_715);
nand U883 (N_883,In_1414,In_694);
or U884 (N_884,In_621,N_179);
xnor U885 (N_885,N_223,In_973);
xor U886 (N_886,N_410,N_35);
and U887 (N_887,In_950,In_1148);
nand U888 (N_888,In_94,N_378);
or U889 (N_889,In_143,N_424);
or U890 (N_890,N_319,In_1005);
xor U891 (N_891,N_185,N_87);
xnor U892 (N_892,N_93,N_322);
and U893 (N_893,In_1322,N_144);
nand U894 (N_894,N_270,N_425);
nand U895 (N_895,In_462,N_347);
and U896 (N_896,In_1440,In_1244);
or U897 (N_897,In_453,N_433);
and U898 (N_898,N_461,In_1081);
and U899 (N_899,In_101,In_1135);
or U900 (N_900,N_133,N_149);
xor U901 (N_901,N_460,N_376);
and U902 (N_902,N_125,In_904);
xnor U903 (N_903,N_49,N_338);
xnor U904 (N_904,In_634,In_329);
xor U905 (N_905,In_1289,N_495);
xnor U906 (N_906,In_1080,N_24);
or U907 (N_907,N_66,In_429);
xor U908 (N_908,N_318,N_108);
nand U909 (N_909,In_1011,In_1349);
or U910 (N_910,N_146,In_360);
xnor U911 (N_911,In_1341,In_478);
or U912 (N_912,N_262,In_966);
nand U913 (N_913,In_132,N_327);
xor U914 (N_914,N_276,N_4);
xor U915 (N_915,N_293,In_946);
or U916 (N_916,In_686,N_206);
nand U917 (N_917,In_1476,N_277);
xnor U918 (N_918,N_209,In_364);
nand U919 (N_919,In_1393,N_271);
nor U920 (N_920,In_164,N_238);
nor U921 (N_921,N_374,In_557);
nand U922 (N_922,N_334,In_864);
nand U923 (N_923,In_642,In_48);
and U924 (N_924,In_289,In_221);
and U925 (N_925,N_492,In_461);
or U926 (N_926,In_88,In_269);
nand U927 (N_927,In_1493,In_127);
and U928 (N_928,N_275,In_725);
nand U929 (N_929,In_208,In_9);
xnor U930 (N_930,N_245,N_237);
nand U931 (N_931,In_168,In_369);
and U932 (N_932,N_120,N_47);
nand U933 (N_933,In_558,In_449);
xnor U934 (N_934,In_1296,In_975);
nor U935 (N_935,In_278,In_857);
or U936 (N_936,N_286,N_372);
and U937 (N_937,N_298,In_1458);
nor U938 (N_938,N_447,In_1280);
or U939 (N_939,In_527,N_296);
nand U940 (N_940,In_1199,N_127);
nor U941 (N_941,In_653,N_309);
and U942 (N_942,In_543,In_460);
xnor U943 (N_943,In_361,N_404);
and U944 (N_944,In_1217,In_248);
nand U945 (N_945,In_220,N_217);
nand U946 (N_946,In_1339,In_779);
or U947 (N_947,In_655,N_89);
or U948 (N_948,In_83,N_240);
or U949 (N_949,N_260,In_805);
xor U950 (N_950,In_782,N_311);
nand U951 (N_951,In_519,In_1145);
nor U952 (N_952,N_450,In_742);
and U953 (N_953,N_34,N_113);
xor U954 (N_954,N_246,In_19);
and U955 (N_955,N_459,N_317);
nand U956 (N_956,In_577,N_252);
nand U957 (N_957,In_885,N_339);
nand U958 (N_958,In_645,In_638);
or U959 (N_959,N_413,In_498);
nand U960 (N_960,N_158,In_419);
nand U961 (N_961,N_486,In_235);
and U962 (N_962,In_1227,N_351);
nand U963 (N_963,In_284,In_1222);
nor U964 (N_964,N_193,In_620);
xor U965 (N_965,N_292,N_25);
or U966 (N_966,N_392,In_698);
and U967 (N_967,In_286,N_408);
xor U968 (N_968,In_1431,N_294);
nor U969 (N_969,In_1076,N_229);
nand U970 (N_970,In_679,In_52);
or U971 (N_971,N_388,N_384);
nand U972 (N_972,In_1419,N_341);
nor U973 (N_973,In_592,N_307);
and U974 (N_974,N_457,N_154);
xnor U975 (N_975,N_290,In_412);
xor U976 (N_976,In_228,In_1276);
or U977 (N_977,In_581,N_333);
or U978 (N_978,N_21,In_849);
nand U979 (N_979,In_457,In_311);
or U980 (N_980,N_50,In_1301);
xor U981 (N_981,N_200,N_405);
nand U982 (N_982,N_126,N_427);
nand U983 (N_983,In_520,In_959);
nand U984 (N_984,N_167,In_41);
xnor U985 (N_985,N_226,N_128);
nand U986 (N_986,N_121,N_242);
or U987 (N_987,N_485,In_915);
nand U988 (N_988,In_66,N_415);
and U989 (N_989,N_222,N_443);
xor U990 (N_990,N_136,N_280);
and U991 (N_991,N_15,In_795);
nor U992 (N_992,N_2,In_1184);
nand U993 (N_993,In_434,In_1283);
and U994 (N_994,N_96,In_1127);
and U995 (N_995,In_493,N_452);
nand U996 (N_996,In_1384,In_50);
xnor U997 (N_997,In_347,N_26);
nand U998 (N_998,N_101,N_97);
xor U999 (N_999,N_248,In_1338);
nor U1000 (N_1000,N_833,N_701);
nor U1001 (N_1001,N_773,N_920);
and U1002 (N_1002,N_868,N_763);
or U1003 (N_1003,N_932,N_681);
and U1004 (N_1004,N_623,N_887);
and U1005 (N_1005,N_737,N_893);
nor U1006 (N_1006,N_759,N_640);
nor U1007 (N_1007,N_591,N_855);
xor U1008 (N_1008,N_999,N_775);
and U1009 (N_1009,N_930,N_965);
nor U1010 (N_1010,N_794,N_718);
and U1011 (N_1011,N_538,N_940);
nand U1012 (N_1012,N_552,N_814);
and U1013 (N_1013,N_757,N_629);
xnor U1014 (N_1014,N_533,N_957);
xnor U1015 (N_1015,N_805,N_791);
xnor U1016 (N_1016,N_960,N_822);
or U1017 (N_1017,N_558,N_783);
or U1018 (N_1018,N_747,N_691);
and U1019 (N_1019,N_816,N_735);
and U1020 (N_1020,N_955,N_636);
nor U1021 (N_1021,N_653,N_981);
and U1022 (N_1022,N_795,N_508);
nand U1023 (N_1023,N_535,N_670);
xor U1024 (N_1024,N_871,N_689);
and U1025 (N_1025,N_943,N_549);
nand U1026 (N_1026,N_996,N_669);
nor U1027 (N_1027,N_824,N_534);
nand U1028 (N_1028,N_873,N_577);
nand U1029 (N_1029,N_821,N_774);
nor U1030 (N_1030,N_739,N_634);
or U1031 (N_1031,N_726,N_556);
xnor U1032 (N_1032,N_786,N_892);
and U1033 (N_1033,N_844,N_576);
nand U1034 (N_1034,N_611,N_647);
nand U1035 (N_1035,N_537,N_870);
or U1036 (N_1036,N_764,N_730);
and U1037 (N_1037,N_727,N_622);
xor U1038 (N_1038,N_595,N_638);
nand U1039 (N_1039,N_696,N_505);
or U1040 (N_1040,N_582,N_706);
nand U1041 (N_1041,N_586,N_863);
and U1042 (N_1042,N_842,N_800);
nor U1043 (N_1043,N_978,N_846);
nand U1044 (N_1044,N_583,N_880);
nor U1045 (N_1045,N_801,N_555);
or U1046 (N_1046,N_803,N_649);
and U1047 (N_1047,N_515,N_808);
and U1048 (N_1048,N_919,N_547);
and U1049 (N_1049,N_904,N_948);
nor U1050 (N_1050,N_756,N_839);
or U1051 (N_1051,N_849,N_657);
nor U1052 (N_1052,N_915,N_709);
xnor U1053 (N_1053,N_598,N_780);
xor U1054 (N_1054,N_970,N_881);
and U1055 (N_1055,N_778,N_787);
nand U1056 (N_1056,N_541,N_543);
xnor U1057 (N_1057,N_722,N_946);
xor U1058 (N_1058,N_924,N_605);
nand U1059 (N_1059,N_607,N_788);
or U1060 (N_1060,N_864,N_560);
nand U1061 (N_1061,N_620,N_914);
and U1062 (N_1062,N_652,N_516);
nor U1063 (N_1063,N_518,N_765);
nand U1064 (N_1064,N_719,N_677);
and U1065 (N_1065,N_832,N_967);
xor U1066 (N_1066,N_521,N_989);
xor U1067 (N_1067,N_771,N_974);
nor U1068 (N_1068,N_553,N_702);
nor U1069 (N_1069,N_950,N_897);
and U1070 (N_1070,N_713,N_966);
nand U1071 (N_1071,N_606,N_721);
xor U1072 (N_1072,N_826,N_860);
and U1073 (N_1073,N_831,N_712);
xor U1074 (N_1074,N_650,N_777);
or U1075 (N_1075,N_819,N_520);
nand U1076 (N_1076,N_615,N_990);
nor U1077 (N_1077,N_517,N_768);
nor U1078 (N_1078,N_628,N_933);
or U1079 (N_1079,N_898,N_852);
nor U1080 (N_1080,N_512,N_663);
nor U1081 (N_1081,N_841,N_890);
nor U1082 (N_1082,N_857,N_593);
xnor U1083 (N_1083,N_834,N_891);
nor U1084 (N_1084,N_529,N_858);
and U1085 (N_1085,N_971,N_980);
and U1086 (N_1086,N_559,N_761);
nand U1087 (N_1087,N_690,N_813);
nor U1088 (N_1088,N_804,N_720);
and U1089 (N_1089,N_776,N_542);
and U1090 (N_1090,N_987,N_716);
or U1091 (N_1091,N_679,N_878);
or U1092 (N_1092,N_995,N_729);
and U1093 (N_1093,N_790,N_641);
xnor U1094 (N_1094,N_835,N_988);
or U1095 (N_1095,N_725,N_711);
and U1096 (N_1096,N_997,N_953);
xnor U1097 (N_1097,N_902,N_926);
xnor U1098 (N_1098,N_564,N_745);
xnor U1099 (N_1099,N_956,N_962);
and U1100 (N_1100,N_917,N_665);
and U1101 (N_1101,N_947,N_928);
xor U1102 (N_1102,N_500,N_862);
nor U1103 (N_1103,N_646,N_799);
or U1104 (N_1104,N_883,N_810);
or U1105 (N_1105,N_596,N_548);
and U1106 (N_1106,N_982,N_993);
nand U1107 (N_1107,N_662,N_510);
nor U1108 (N_1108,N_744,N_900);
nor U1109 (N_1109,N_554,N_884);
and U1110 (N_1110,N_886,N_624);
or U1111 (N_1111,N_557,N_680);
and U1112 (N_1112,N_700,N_659);
nor U1113 (N_1113,N_861,N_837);
and U1114 (N_1114,N_600,N_710);
nor U1115 (N_1115,N_545,N_695);
or U1116 (N_1116,N_676,N_723);
and U1117 (N_1117,N_941,N_699);
or U1118 (N_1118,N_825,N_736);
and U1119 (N_1119,N_575,N_642);
xor U1120 (N_1120,N_977,N_707);
nor U1121 (N_1121,N_877,N_895);
and U1122 (N_1122,N_668,N_530);
or U1123 (N_1123,N_644,N_683);
nor U1124 (N_1124,N_592,N_762);
and U1125 (N_1125,N_798,N_551);
or U1126 (N_1126,N_621,N_632);
xor U1127 (N_1127,N_903,N_760);
nand U1128 (N_1128,N_686,N_567);
or U1129 (N_1129,N_626,N_572);
or U1130 (N_1130,N_708,N_931);
xor U1131 (N_1131,N_963,N_589);
xor U1132 (N_1132,N_751,N_525);
nor U1133 (N_1133,N_934,N_918);
nand U1134 (N_1134,N_938,N_513);
or U1135 (N_1135,N_850,N_655);
or U1136 (N_1136,N_975,N_630);
and U1137 (N_1137,N_879,N_692);
and U1138 (N_1138,N_563,N_748);
nor U1139 (N_1139,N_531,N_532);
nor U1140 (N_1140,N_927,N_882);
nand U1141 (N_1141,N_627,N_829);
and U1142 (N_1142,N_767,N_945);
and U1143 (N_1143,N_579,N_769);
nor U1144 (N_1144,N_840,N_675);
xor U1145 (N_1145,N_867,N_610);
nand U1146 (N_1146,N_984,N_565);
and U1147 (N_1147,N_848,N_820);
and U1148 (N_1148,N_958,N_601);
nor U1149 (N_1149,N_754,N_590);
and U1150 (N_1150,N_694,N_571);
or U1151 (N_1151,N_509,N_703);
nand U1152 (N_1152,N_588,N_865);
and U1153 (N_1153,N_986,N_845);
and U1154 (N_1154,N_522,N_648);
and U1155 (N_1155,N_929,N_942);
and U1156 (N_1156,N_847,N_830);
xor U1157 (N_1157,N_959,N_750);
xnor U1158 (N_1158,N_749,N_580);
and U1159 (N_1159,N_753,N_985);
nand U1160 (N_1160,N_734,N_746);
nor U1161 (N_1161,N_869,N_639);
nor U1162 (N_1162,N_672,N_550);
xor U1163 (N_1163,N_608,N_523);
nor U1164 (N_1164,N_823,N_570);
and U1165 (N_1165,N_802,N_766);
or U1166 (N_1166,N_501,N_876);
nor U1167 (N_1167,N_910,N_674);
xnor U1168 (N_1168,N_514,N_740);
nand U1169 (N_1169,N_643,N_617);
nor U1170 (N_1170,N_685,N_658);
and U1171 (N_1171,N_717,N_952);
nor U1172 (N_1172,N_896,N_954);
nand U1173 (N_1173,N_507,N_998);
xnor U1174 (N_1174,N_797,N_859);
xnor U1175 (N_1175,N_687,N_939);
xnor U1176 (N_1176,N_752,N_673);
and U1177 (N_1177,N_526,N_809);
nand U1178 (N_1178,N_854,N_528);
or U1179 (N_1179,N_781,N_504);
nand U1180 (N_1180,N_866,N_656);
xor U1181 (N_1181,N_594,N_603);
nor U1182 (N_1182,N_964,N_540);
xor U1183 (N_1183,N_705,N_782);
or U1184 (N_1184,N_875,N_568);
nor U1185 (N_1185,N_697,N_561);
xor U1186 (N_1186,N_732,N_524);
xnor U1187 (N_1187,N_874,N_923);
and U1188 (N_1188,N_581,N_664);
xor U1189 (N_1189,N_693,N_992);
and U1190 (N_1190,N_812,N_502);
xor U1191 (N_1191,N_573,N_838);
xor U1192 (N_1192,N_843,N_618);
or U1193 (N_1193,N_885,N_704);
and U1194 (N_1194,N_968,N_613);
or U1195 (N_1195,N_894,N_602);
nor U1196 (N_1196,N_836,N_536);
nand U1197 (N_1197,N_973,N_574);
nor U1198 (N_1198,N_637,N_546);
nor U1199 (N_1199,N_544,N_682);
and U1200 (N_1200,N_566,N_738);
nor U1201 (N_1201,N_935,N_527);
xor U1202 (N_1202,N_944,N_913);
nand U1203 (N_1203,N_585,N_949);
xnor U1204 (N_1204,N_625,N_916);
xnor U1205 (N_1205,N_772,N_667);
xnor U1206 (N_1206,N_912,N_951);
nand U1207 (N_1207,N_569,N_827);
or U1208 (N_1208,N_660,N_969);
xnor U1209 (N_1209,N_724,N_806);
and U1210 (N_1210,N_907,N_856);
nor U1211 (N_1211,N_743,N_784);
or U1212 (N_1212,N_792,N_818);
or U1213 (N_1213,N_714,N_811);
or U1214 (N_1214,N_853,N_922);
or U1215 (N_1215,N_645,N_909);
nor U1216 (N_1216,N_631,N_688);
and U1217 (N_1217,N_506,N_651);
or U1218 (N_1218,N_728,N_936);
and U1219 (N_1219,N_901,N_991);
xnor U1220 (N_1220,N_614,N_539);
and U1221 (N_1221,N_889,N_511);
and U1222 (N_1222,N_961,N_587);
nand U1223 (N_1223,N_684,N_976);
nand U1224 (N_1224,N_872,N_562);
or U1225 (N_1225,N_619,N_789);
or U1226 (N_1226,N_888,N_817);
nand U1227 (N_1227,N_599,N_731);
nand U1228 (N_1228,N_578,N_633);
nand U1229 (N_1229,N_742,N_815);
and U1230 (N_1230,N_807,N_906);
nor U1231 (N_1231,N_678,N_983);
and U1232 (N_1232,N_925,N_793);
nor U1233 (N_1233,N_796,N_828);
nor U1234 (N_1234,N_921,N_899);
nand U1235 (N_1235,N_911,N_612);
and U1236 (N_1236,N_661,N_654);
nor U1237 (N_1237,N_604,N_908);
and U1238 (N_1238,N_715,N_851);
or U1239 (N_1239,N_698,N_972);
or U1240 (N_1240,N_741,N_503);
or U1241 (N_1241,N_666,N_785);
and U1242 (N_1242,N_905,N_979);
nor U1243 (N_1243,N_733,N_584);
and U1244 (N_1244,N_770,N_519);
nand U1245 (N_1245,N_758,N_609);
nand U1246 (N_1246,N_755,N_597);
nand U1247 (N_1247,N_937,N_779);
xnor U1248 (N_1248,N_994,N_616);
and U1249 (N_1249,N_635,N_671);
nand U1250 (N_1250,N_644,N_816);
nand U1251 (N_1251,N_549,N_988);
and U1252 (N_1252,N_824,N_983);
xnor U1253 (N_1253,N_972,N_567);
or U1254 (N_1254,N_842,N_817);
or U1255 (N_1255,N_705,N_621);
or U1256 (N_1256,N_684,N_913);
or U1257 (N_1257,N_730,N_773);
nand U1258 (N_1258,N_884,N_997);
nand U1259 (N_1259,N_734,N_573);
or U1260 (N_1260,N_810,N_605);
nand U1261 (N_1261,N_945,N_771);
and U1262 (N_1262,N_967,N_689);
and U1263 (N_1263,N_683,N_858);
nand U1264 (N_1264,N_749,N_841);
or U1265 (N_1265,N_892,N_896);
nand U1266 (N_1266,N_543,N_862);
xor U1267 (N_1267,N_570,N_921);
nand U1268 (N_1268,N_563,N_506);
xnor U1269 (N_1269,N_594,N_940);
and U1270 (N_1270,N_580,N_947);
or U1271 (N_1271,N_915,N_950);
nor U1272 (N_1272,N_814,N_933);
nor U1273 (N_1273,N_804,N_677);
or U1274 (N_1274,N_851,N_889);
or U1275 (N_1275,N_615,N_933);
nand U1276 (N_1276,N_945,N_732);
nand U1277 (N_1277,N_541,N_713);
nand U1278 (N_1278,N_598,N_732);
or U1279 (N_1279,N_653,N_990);
and U1280 (N_1280,N_818,N_649);
nor U1281 (N_1281,N_603,N_926);
xnor U1282 (N_1282,N_800,N_651);
and U1283 (N_1283,N_743,N_725);
nand U1284 (N_1284,N_764,N_715);
nor U1285 (N_1285,N_528,N_901);
nand U1286 (N_1286,N_615,N_504);
nor U1287 (N_1287,N_929,N_884);
or U1288 (N_1288,N_844,N_928);
nor U1289 (N_1289,N_801,N_918);
nor U1290 (N_1290,N_727,N_787);
nand U1291 (N_1291,N_924,N_825);
or U1292 (N_1292,N_972,N_766);
and U1293 (N_1293,N_930,N_731);
xor U1294 (N_1294,N_786,N_585);
and U1295 (N_1295,N_533,N_677);
nand U1296 (N_1296,N_833,N_552);
or U1297 (N_1297,N_757,N_724);
xor U1298 (N_1298,N_854,N_860);
or U1299 (N_1299,N_794,N_959);
or U1300 (N_1300,N_899,N_645);
or U1301 (N_1301,N_614,N_717);
and U1302 (N_1302,N_743,N_785);
and U1303 (N_1303,N_871,N_903);
xnor U1304 (N_1304,N_866,N_804);
nor U1305 (N_1305,N_911,N_556);
nor U1306 (N_1306,N_729,N_862);
nor U1307 (N_1307,N_778,N_766);
xnor U1308 (N_1308,N_593,N_817);
xor U1309 (N_1309,N_723,N_788);
or U1310 (N_1310,N_940,N_519);
nand U1311 (N_1311,N_836,N_971);
xor U1312 (N_1312,N_525,N_845);
or U1313 (N_1313,N_929,N_606);
xor U1314 (N_1314,N_965,N_851);
or U1315 (N_1315,N_875,N_852);
and U1316 (N_1316,N_900,N_925);
and U1317 (N_1317,N_970,N_637);
nor U1318 (N_1318,N_655,N_968);
or U1319 (N_1319,N_802,N_809);
or U1320 (N_1320,N_962,N_649);
nor U1321 (N_1321,N_739,N_672);
xor U1322 (N_1322,N_904,N_507);
nand U1323 (N_1323,N_678,N_592);
xnor U1324 (N_1324,N_780,N_910);
and U1325 (N_1325,N_691,N_997);
or U1326 (N_1326,N_680,N_675);
nor U1327 (N_1327,N_886,N_533);
nand U1328 (N_1328,N_816,N_791);
xor U1329 (N_1329,N_601,N_910);
and U1330 (N_1330,N_582,N_945);
nor U1331 (N_1331,N_612,N_689);
xor U1332 (N_1332,N_862,N_672);
xor U1333 (N_1333,N_725,N_814);
nor U1334 (N_1334,N_889,N_613);
nor U1335 (N_1335,N_732,N_805);
nand U1336 (N_1336,N_879,N_935);
nand U1337 (N_1337,N_826,N_768);
or U1338 (N_1338,N_722,N_562);
or U1339 (N_1339,N_678,N_714);
nand U1340 (N_1340,N_879,N_992);
xor U1341 (N_1341,N_960,N_808);
or U1342 (N_1342,N_627,N_622);
nand U1343 (N_1343,N_762,N_677);
nor U1344 (N_1344,N_815,N_940);
xnor U1345 (N_1345,N_858,N_633);
nand U1346 (N_1346,N_927,N_600);
nor U1347 (N_1347,N_710,N_922);
nor U1348 (N_1348,N_684,N_564);
nand U1349 (N_1349,N_876,N_915);
nand U1350 (N_1350,N_988,N_594);
or U1351 (N_1351,N_720,N_539);
nor U1352 (N_1352,N_898,N_825);
or U1353 (N_1353,N_627,N_697);
nor U1354 (N_1354,N_669,N_814);
nand U1355 (N_1355,N_883,N_947);
nand U1356 (N_1356,N_549,N_955);
nand U1357 (N_1357,N_831,N_564);
xnor U1358 (N_1358,N_663,N_866);
xnor U1359 (N_1359,N_538,N_546);
xnor U1360 (N_1360,N_713,N_501);
xnor U1361 (N_1361,N_987,N_732);
and U1362 (N_1362,N_868,N_803);
nor U1363 (N_1363,N_560,N_708);
nor U1364 (N_1364,N_888,N_862);
nand U1365 (N_1365,N_712,N_570);
or U1366 (N_1366,N_715,N_924);
nor U1367 (N_1367,N_816,N_518);
xor U1368 (N_1368,N_963,N_517);
xor U1369 (N_1369,N_751,N_843);
nand U1370 (N_1370,N_544,N_580);
or U1371 (N_1371,N_647,N_898);
or U1372 (N_1372,N_900,N_725);
or U1373 (N_1373,N_843,N_987);
and U1374 (N_1374,N_852,N_794);
xnor U1375 (N_1375,N_641,N_737);
xnor U1376 (N_1376,N_870,N_914);
nor U1377 (N_1377,N_661,N_990);
xnor U1378 (N_1378,N_966,N_587);
xor U1379 (N_1379,N_715,N_775);
or U1380 (N_1380,N_580,N_672);
nor U1381 (N_1381,N_809,N_789);
and U1382 (N_1382,N_526,N_874);
or U1383 (N_1383,N_596,N_902);
nor U1384 (N_1384,N_964,N_999);
nor U1385 (N_1385,N_796,N_692);
or U1386 (N_1386,N_998,N_938);
nand U1387 (N_1387,N_981,N_889);
nor U1388 (N_1388,N_513,N_559);
or U1389 (N_1389,N_627,N_761);
nand U1390 (N_1390,N_660,N_922);
and U1391 (N_1391,N_990,N_579);
or U1392 (N_1392,N_915,N_596);
nor U1393 (N_1393,N_806,N_712);
xor U1394 (N_1394,N_943,N_606);
xor U1395 (N_1395,N_774,N_753);
or U1396 (N_1396,N_851,N_663);
xor U1397 (N_1397,N_682,N_767);
or U1398 (N_1398,N_600,N_632);
and U1399 (N_1399,N_570,N_824);
and U1400 (N_1400,N_795,N_634);
nand U1401 (N_1401,N_956,N_885);
and U1402 (N_1402,N_526,N_673);
or U1403 (N_1403,N_948,N_911);
nand U1404 (N_1404,N_786,N_634);
xor U1405 (N_1405,N_907,N_745);
xnor U1406 (N_1406,N_981,N_843);
nand U1407 (N_1407,N_656,N_540);
nor U1408 (N_1408,N_827,N_978);
and U1409 (N_1409,N_847,N_559);
and U1410 (N_1410,N_698,N_740);
nor U1411 (N_1411,N_575,N_551);
nand U1412 (N_1412,N_501,N_764);
nor U1413 (N_1413,N_546,N_829);
nand U1414 (N_1414,N_911,N_838);
nand U1415 (N_1415,N_507,N_840);
nor U1416 (N_1416,N_806,N_841);
nand U1417 (N_1417,N_510,N_663);
and U1418 (N_1418,N_509,N_765);
xnor U1419 (N_1419,N_812,N_586);
or U1420 (N_1420,N_511,N_515);
nand U1421 (N_1421,N_940,N_832);
nand U1422 (N_1422,N_817,N_558);
nand U1423 (N_1423,N_570,N_659);
or U1424 (N_1424,N_729,N_581);
or U1425 (N_1425,N_971,N_555);
or U1426 (N_1426,N_779,N_879);
nor U1427 (N_1427,N_703,N_719);
and U1428 (N_1428,N_820,N_833);
or U1429 (N_1429,N_869,N_664);
and U1430 (N_1430,N_785,N_528);
nand U1431 (N_1431,N_779,N_717);
nor U1432 (N_1432,N_876,N_973);
xor U1433 (N_1433,N_792,N_819);
nand U1434 (N_1434,N_937,N_983);
and U1435 (N_1435,N_816,N_752);
and U1436 (N_1436,N_873,N_736);
nand U1437 (N_1437,N_814,N_903);
and U1438 (N_1438,N_577,N_661);
xor U1439 (N_1439,N_747,N_845);
or U1440 (N_1440,N_652,N_597);
nand U1441 (N_1441,N_578,N_980);
nand U1442 (N_1442,N_522,N_667);
nor U1443 (N_1443,N_996,N_723);
and U1444 (N_1444,N_908,N_687);
xor U1445 (N_1445,N_734,N_917);
nor U1446 (N_1446,N_786,N_903);
xor U1447 (N_1447,N_965,N_885);
nor U1448 (N_1448,N_654,N_613);
and U1449 (N_1449,N_557,N_624);
or U1450 (N_1450,N_507,N_962);
nand U1451 (N_1451,N_597,N_647);
xnor U1452 (N_1452,N_767,N_836);
and U1453 (N_1453,N_811,N_812);
and U1454 (N_1454,N_823,N_897);
or U1455 (N_1455,N_861,N_949);
nor U1456 (N_1456,N_780,N_885);
or U1457 (N_1457,N_731,N_660);
nand U1458 (N_1458,N_860,N_613);
or U1459 (N_1459,N_807,N_655);
nor U1460 (N_1460,N_500,N_738);
or U1461 (N_1461,N_619,N_598);
xor U1462 (N_1462,N_640,N_833);
and U1463 (N_1463,N_824,N_575);
nand U1464 (N_1464,N_720,N_964);
or U1465 (N_1465,N_534,N_677);
nor U1466 (N_1466,N_896,N_877);
or U1467 (N_1467,N_602,N_860);
nand U1468 (N_1468,N_736,N_546);
or U1469 (N_1469,N_636,N_819);
or U1470 (N_1470,N_944,N_501);
nor U1471 (N_1471,N_887,N_874);
or U1472 (N_1472,N_711,N_889);
nand U1473 (N_1473,N_590,N_728);
nand U1474 (N_1474,N_876,N_563);
or U1475 (N_1475,N_794,N_643);
nand U1476 (N_1476,N_580,N_716);
or U1477 (N_1477,N_538,N_787);
nand U1478 (N_1478,N_752,N_505);
nand U1479 (N_1479,N_768,N_861);
or U1480 (N_1480,N_543,N_670);
and U1481 (N_1481,N_513,N_789);
nor U1482 (N_1482,N_783,N_571);
nor U1483 (N_1483,N_694,N_632);
xor U1484 (N_1484,N_507,N_841);
nand U1485 (N_1485,N_648,N_917);
and U1486 (N_1486,N_951,N_500);
xnor U1487 (N_1487,N_745,N_768);
nand U1488 (N_1488,N_955,N_517);
and U1489 (N_1489,N_591,N_959);
nor U1490 (N_1490,N_957,N_558);
and U1491 (N_1491,N_609,N_960);
and U1492 (N_1492,N_803,N_853);
nor U1493 (N_1493,N_952,N_672);
nand U1494 (N_1494,N_945,N_621);
or U1495 (N_1495,N_514,N_627);
nor U1496 (N_1496,N_946,N_790);
xnor U1497 (N_1497,N_664,N_953);
nor U1498 (N_1498,N_628,N_673);
or U1499 (N_1499,N_547,N_670);
xor U1500 (N_1500,N_1372,N_1055);
or U1501 (N_1501,N_1194,N_1152);
xnor U1502 (N_1502,N_1149,N_1123);
nand U1503 (N_1503,N_1090,N_1038);
and U1504 (N_1504,N_1078,N_1366);
and U1505 (N_1505,N_1488,N_1013);
or U1506 (N_1506,N_1105,N_1432);
xor U1507 (N_1507,N_1018,N_1180);
and U1508 (N_1508,N_1251,N_1408);
xor U1509 (N_1509,N_1178,N_1283);
nor U1510 (N_1510,N_1080,N_1276);
and U1511 (N_1511,N_1231,N_1493);
xor U1512 (N_1512,N_1325,N_1181);
xor U1513 (N_1513,N_1222,N_1484);
xnor U1514 (N_1514,N_1371,N_1050);
and U1515 (N_1515,N_1249,N_1328);
and U1516 (N_1516,N_1310,N_1485);
and U1517 (N_1517,N_1095,N_1256);
nor U1518 (N_1518,N_1011,N_1244);
nand U1519 (N_1519,N_1499,N_1397);
or U1520 (N_1520,N_1386,N_1461);
or U1521 (N_1521,N_1111,N_1028);
nand U1522 (N_1522,N_1466,N_1370);
nor U1523 (N_1523,N_1179,N_1447);
or U1524 (N_1524,N_1395,N_1435);
or U1525 (N_1525,N_1393,N_1046);
xor U1526 (N_1526,N_1066,N_1341);
nor U1527 (N_1527,N_1198,N_1073);
and U1528 (N_1528,N_1155,N_1462);
or U1529 (N_1529,N_1245,N_1048);
and U1530 (N_1530,N_1496,N_1443);
xnor U1531 (N_1531,N_1188,N_1166);
nor U1532 (N_1532,N_1103,N_1426);
and U1533 (N_1533,N_1262,N_1373);
nand U1534 (N_1534,N_1148,N_1479);
xor U1535 (N_1535,N_1380,N_1071);
nor U1536 (N_1536,N_1475,N_1312);
nor U1537 (N_1537,N_1032,N_1278);
and U1538 (N_1538,N_1202,N_1431);
and U1539 (N_1539,N_1324,N_1137);
nand U1540 (N_1540,N_1117,N_1357);
nor U1541 (N_1541,N_1215,N_1346);
xor U1542 (N_1542,N_1454,N_1124);
or U1543 (N_1543,N_1107,N_1358);
xor U1544 (N_1544,N_1410,N_1045);
nand U1545 (N_1545,N_1472,N_1131);
nand U1546 (N_1546,N_1322,N_1250);
or U1547 (N_1547,N_1405,N_1189);
xor U1548 (N_1548,N_1171,N_1470);
or U1549 (N_1549,N_1333,N_1340);
or U1550 (N_1550,N_1182,N_1449);
or U1551 (N_1551,N_1337,N_1116);
xor U1552 (N_1552,N_1343,N_1265);
and U1553 (N_1553,N_1368,N_1299);
nor U1554 (N_1554,N_1017,N_1186);
xor U1555 (N_1555,N_1026,N_1455);
xnor U1556 (N_1556,N_1204,N_1412);
xor U1557 (N_1557,N_1275,N_1438);
xnor U1558 (N_1558,N_1062,N_1396);
or U1559 (N_1559,N_1375,N_1390);
or U1560 (N_1560,N_1169,N_1154);
nand U1561 (N_1561,N_1218,N_1453);
and U1562 (N_1562,N_1318,N_1075);
nor U1563 (N_1563,N_1331,N_1269);
nor U1564 (N_1564,N_1361,N_1112);
or U1565 (N_1565,N_1162,N_1190);
nand U1566 (N_1566,N_1126,N_1404);
nand U1567 (N_1567,N_1019,N_1293);
nand U1568 (N_1568,N_1016,N_1012);
and U1569 (N_1569,N_1321,N_1000);
xor U1570 (N_1570,N_1238,N_1350);
nor U1571 (N_1571,N_1139,N_1138);
nand U1572 (N_1572,N_1351,N_1211);
and U1573 (N_1573,N_1237,N_1482);
xor U1574 (N_1574,N_1196,N_1216);
or U1575 (N_1575,N_1077,N_1260);
nor U1576 (N_1576,N_1206,N_1439);
nand U1577 (N_1577,N_1392,N_1086);
or U1578 (N_1578,N_1052,N_1021);
nand U1579 (N_1579,N_1460,N_1213);
or U1580 (N_1580,N_1008,N_1414);
nor U1581 (N_1581,N_1301,N_1199);
or U1582 (N_1582,N_1286,N_1415);
nand U1583 (N_1583,N_1130,N_1458);
or U1584 (N_1584,N_1221,N_1184);
nand U1585 (N_1585,N_1474,N_1441);
and U1586 (N_1586,N_1161,N_1029);
nor U1587 (N_1587,N_1489,N_1072);
xor U1588 (N_1588,N_1342,N_1445);
xor U1589 (N_1589,N_1413,N_1291);
nor U1590 (N_1590,N_1156,N_1088);
xor U1591 (N_1591,N_1335,N_1409);
nor U1592 (N_1592,N_1151,N_1022);
and U1593 (N_1593,N_1259,N_1074);
nor U1594 (N_1594,N_1121,N_1239);
nand U1595 (N_1595,N_1175,N_1243);
and U1596 (N_1596,N_1360,N_1434);
xor U1597 (N_1597,N_1314,N_1159);
nor U1598 (N_1598,N_1058,N_1132);
xor U1599 (N_1599,N_1354,N_1091);
nor U1600 (N_1600,N_1287,N_1427);
nor U1601 (N_1601,N_1320,N_1036);
nor U1602 (N_1602,N_1102,N_1030);
and U1603 (N_1603,N_1068,N_1400);
and U1604 (N_1604,N_1307,N_1120);
and U1605 (N_1605,N_1254,N_1134);
or U1606 (N_1606,N_1067,N_1349);
xor U1607 (N_1607,N_1290,N_1469);
and U1608 (N_1608,N_1228,N_1150);
nand U1609 (N_1609,N_1060,N_1119);
nor U1610 (N_1610,N_1407,N_1429);
nor U1611 (N_1611,N_1428,N_1172);
and U1612 (N_1612,N_1140,N_1356);
nor U1613 (N_1613,N_1035,N_1145);
and U1614 (N_1614,N_1200,N_1096);
xnor U1615 (N_1615,N_1279,N_1133);
and U1616 (N_1616,N_1402,N_1344);
nand U1617 (N_1617,N_1258,N_1118);
nand U1618 (N_1618,N_1348,N_1195);
and U1619 (N_1619,N_1197,N_1127);
nor U1620 (N_1620,N_1025,N_1101);
and U1621 (N_1621,N_1252,N_1329);
xor U1622 (N_1622,N_1212,N_1332);
and U1623 (N_1623,N_1316,N_1083);
nand U1624 (N_1624,N_1064,N_1241);
xor U1625 (N_1625,N_1033,N_1242);
xnor U1626 (N_1626,N_1113,N_1494);
and U1627 (N_1627,N_1217,N_1006);
nor U1628 (N_1628,N_1277,N_1153);
nor U1629 (N_1629,N_1085,N_1492);
nor U1630 (N_1630,N_1367,N_1053);
or U1631 (N_1631,N_1388,N_1313);
xnor U1632 (N_1632,N_1135,N_1236);
or U1633 (N_1633,N_1302,N_1323);
and U1634 (N_1634,N_1024,N_1311);
and U1635 (N_1635,N_1420,N_1487);
xor U1636 (N_1636,N_1285,N_1230);
nand U1637 (N_1637,N_1143,N_1417);
or U1638 (N_1638,N_1480,N_1292);
or U1639 (N_1639,N_1020,N_1491);
nor U1640 (N_1640,N_1391,N_1057);
xor U1641 (N_1641,N_1339,N_1266);
or U1642 (N_1642,N_1082,N_1300);
or U1643 (N_1643,N_1468,N_1257);
or U1644 (N_1644,N_1289,N_1023);
xnor U1645 (N_1645,N_1129,N_1224);
nand U1646 (N_1646,N_1295,N_1003);
or U1647 (N_1647,N_1015,N_1108);
nand U1648 (N_1648,N_1205,N_1010);
xnor U1649 (N_1649,N_1097,N_1219);
nor U1650 (N_1650,N_1208,N_1442);
and U1651 (N_1651,N_1183,N_1079);
nand U1652 (N_1652,N_1170,N_1115);
nand U1653 (N_1653,N_1065,N_1042);
nand U1654 (N_1654,N_1220,N_1041);
and U1655 (N_1655,N_1362,N_1471);
and U1656 (N_1656,N_1355,N_1389);
xor U1657 (N_1657,N_1384,N_1319);
or U1658 (N_1658,N_1326,N_1037);
xor U1659 (N_1659,N_1309,N_1353);
nor U1660 (N_1660,N_1187,N_1398);
xor U1661 (N_1661,N_1114,N_1306);
nor U1662 (N_1662,N_1363,N_1305);
nor U1663 (N_1663,N_1210,N_1359);
and U1664 (N_1664,N_1247,N_1061);
nor U1665 (N_1665,N_1270,N_1002);
xnor U1666 (N_1666,N_1044,N_1059);
and U1667 (N_1667,N_1416,N_1467);
nor U1668 (N_1668,N_1490,N_1007);
and U1669 (N_1669,N_1418,N_1076);
xor U1670 (N_1670,N_1282,N_1478);
or U1671 (N_1671,N_1040,N_1089);
nor U1672 (N_1672,N_1125,N_1165);
xor U1673 (N_1673,N_1261,N_1092);
or U1674 (N_1674,N_1225,N_1255);
xor U1675 (N_1675,N_1448,N_1164);
nand U1676 (N_1676,N_1268,N_1174);
or U1677 (N_1677,N_1436,N_1147);
or U1678 (N_1678,N_1288,N_1450);
xnor U1679 (N_1679,N_1476,N_1419);
nor U1680 (N_1680,N_1226,N_1176);
and U1681 (N_1681,N_1377,N_1433);
xor U1682 (N_1682,N_1203,N_1142);
and U1683 (N_1683,N_1483,N_1034);
nand U1684 (N_1684,N_1387,N_1157);
nand U1685 (N_1685,N_1146,N_1223);
and U1686 (N_1686,N_1136,N_1235);
and U1687 (N_1687,N_1336,N_1451);
nand U1688 (N_1688,N_1168,N_1347);
or U1689 (N_1689,N_1069,N_1274);
nor U1690 (N_1690,N_1338,N_1369);
or U1691 (N_1691,N_1303,N_1411);
or U1692 (N_1692,N_1498,N_1296);
nor U1693 (N_1693,N_1284,N_1141);
nor U1694 (N_1694,N_1234,N_1081);
nor U1695 (N_1695,N_1158,N_1444);
nand U1696 (N_1696,N_1177,N_1173);
nand U1697 (N_1697,N_1214,N_1106);
or U1698 (N_1698,N_1457,N_1122);
nand U1699 (N_1699,N_1049,N_1423);
and U1700 (N_1700,N_1163,N_1009);
and U1701 (N_1701,N_1110,N_1463);
or U1702 (N_1702,N_1263,N_1233);
nand U1703 (N_1703,N_1464,N_1031);
or U1704 (N_1704,N_1063,N_1334);
or U1705 (N_1705,N_1465,N_1253);
xnor U1706 (N_1706,N_1481,N_1424);
nor U1707 (N_1707,N_1425,N_1001);
xnor U1708 (N_1708,N_1298,N_1452);
nand U1709 (N_1709,N_1193,N_1403);
or U1710 (N_1710,N_1229,N_1185);
nor U1711 (N_1711,N_1376,N_1308);
xor U1712 (N_1712,N_1128,N_1051);
nand U1713 (N_1713,N_1273,N_1232);
and U1714 (N_1714,N_1459,N_1495);
and U1715 (N_1715,N_1039,N_1437);
nand U1716 (N_1716,N_1246,N_1227);
and U1717 (N_1717,N_1486,N_1027);
nand U1718 (N_1718,N_1381,N_1473);
xor U1719 (N_1719,N_1379,N_1192);
nand U1720 (N_1720,N_1297,N_1281);
or U1721 (N_1721,N_1374,N_1382);
nand U1722 (N_1722,N_1345,N_1385);
nand U1723 (N_1723,N_1248,N_1327);
xor U1724 (N_1724,N_1271,N_1047);
nor U1725 (N_1725,N_1005,N_1167);
or U1726 (N_1726,N_1207,N_1209);
and U1727 (N_1727,N_1456,N_1421);
xnor U1728 (N_1728,N_1430,N_1098);
nor U1729 (N_1729,N_1440,N_1056);
and U1730 (N_1730,N_1330,N_1004);
nor U1731 (N_1731,N_1422,N_1264);
or U1732 (N_1732,N_1267,N_1054);
and U1733 (N_1733,N_1087,N_1014);
nor U1734 (N_1734,N_1104,N_1317);
xor U1735 (N_1735,N_1070,N_1084);
xnor U1736 (N_1736,N_1272,N_1378);
nand U1737 (N_1737,N_1144,N_1094);
or U1738 (N_1738,N_1352,N_1191);
and U1739 (N_1739,N_1401,N_1399);
nand U1740 (N_1740,N_1294,N_1477);
and U1741 (N_1741,N_1109,N_1160);
or U1742 (N_1742,N_1497,N_1365);
and U1743 (N_1743,N_1315,N_1406);
and U1744 (N_1744,N_1364,N_1304);
or U1745 (N_1745,N_1383,N_1446);
nand U1746 (N_1746,N_1043,N_1280);
nand U1747 (N_1747,N_1099,N_1093);
xnor U1748 (N_1748,N_1100,N_1240);
nor U1749 (N_1749,N_1394,N_1201);
xnor U1750 (N_1750,N_1097,N_1469);
and U1751 (N_1751,N_1222,N_1200);
nand U1752 (N_1752,N_1367,N_1189);
xor U1753 (N_1753,N_1045,N_1018);
nor U1754 (N_1754,N_1493,N_1139);
nand U1755 (N_1755,N_1224,N_1427);
and U1756 (N_1756,N_1445,N_1088);
nand U1757 (N_1757,N_1013,N_1010);
nand U1758 (N_1758,N_1030,N_1392);
nand U1759 (N_1759,N_1220,N_1127);
or U1760 (N_1760,N_1101,N_1185);
nand U1761 (N_1761,N_1135,N_1273);
nor U1762 (N_1762,N_1361,N_1454);
nor U1763 (N_1763,N_1325,N_1380);
or U1764 (N_1764,N_1047,N_1388);
nand U1765 (N_1765,N_1126,N_1280);
or U1766 (N_1766,N_1037,N_1468);
or U1767 (N_1767,N_1358,N_1325);
or U1768 (N_1768,N_1169,N_1192);
xnor U1769 (N_1769,N_1185,N_1212);
or U1770 (N_1770,N_1195,N_1112);
and U1771 (N_1771,N_1081,N_1025);
nand U1772 (N_1772,N_1360,N_1400);
nor U1773 (N_1773,N_1299,N_1098);
xnor U1774 (N_1774,N_1038,N_1282);
and U1775 (N_1775,N_1155,N_1445);
xor U1776 (N_1776,N_1072,N_1375);
nand U1777 (N_1777,N_1233,N_1130);
nand U1778 (N_1778,N_1158,N_1449);
and U1779 (N_1779,N_1490,N_1010);
nor U1780 (N_1780,N_1332,N_1017);
and U1781 (N_1781,N_1311,N_1285);
nand U1782 (N_1782,N_1292,N_1087);
nand U1783 (N_1783,N_1287,N_1077);
and U1784 (N_1784,N_1158,N_1397);
nand U1785 (N_1785,N_1036,N_1195);
and U1786 (N_1786,N_1056,N_1357);
and U1787 (N_1787,N_1149,N_1377);
and U1788 (N_1788,N_1432,N_1387);
or U1789 (N_1789,N_1494,N_1224);
nor U1790 (N_1790,N_1420,N_1154);
nand U1791 (N_1791,N_1106,N_1265);
and U1792 (N_1792,N_1048,N_1054);
nor U1793 (N_1793,N_1227,N_1016);
nand U1794 (N_1794,N_1110,N_1050);
or U1795 (N_1795,N_1232,N_1362);
xnor U1796 (N_1796,N_1483,N_1057);
or U1797 (N_1797,N_1094,N_1194);
nor U1798 (N_1798,N_1014,N_1156);
xnor U1799 (N_1799,N_1019,N_1204);
and U1800 (N_1800,N_1455,N_1119);
nand U1801 (N_1801,N_1426,N_1252);
nor U1802 (N_1802,N_1060,N_1460);
and U1803 (N_1803,N_1009,N_1070);
nand U1804 (N_1804,N_1034,N_1248);
xnor U1805 (N_1805,N_1314,N_1388);
nand U1806 (N_1806,N_1249,N_1421);
nor U1807 (N_1807,N_1461,N_1499);
or U1808 (N_1808,N_1324,N_1171);
and U1809 (N_1809,N_1259,N_1140);
nand U1810 (N_1810,N_1257,N_1286);
xor U1811 (N_1811,N_1416,N_1237);
xnor U1812 (N_1812,N_1494,N_1106);
nand U1813 (N_1813,N_1163,N_1329);
xnor U1814 (N_1814,N_1434,N_1305);
nand U1815 (N_1815,N_1128,N_1331);
or U1816 (N_1816,N_1236,N_1041);
or U1817 (N_1817,N_1045,N_1469);
nand U1818 (N_1818,N_1039,N_1349);
or U1819 (N_1819,N_1413,N_1313);
or U1820 (N_1820,N_1080,N_1295);
nor U1821 (N_1821,N_1019,N_1394);
nor U1822 (N_1822,N_1164,N_1136);
nor U1823 (N_1823,N_1250,N_1167);
or U1824 (N_1824,N_1364,N_1136);
xnor U1825 (N_1825,N_1358,N_1030);
nor U1826 (N_1826,N_1436,N_1249);
nor U1827 (N_1827,N_1437,N_1221);
nand U1828 (N_1828,N_1038,N_1221);
xnor U1829 (N_1829,N_1375,N_1489);
xnor U1830 (N_1830,N_1296,N_1404);
nand U1831 (N_1831,N_1181,N_1069);
nor U1832 (N_1832,N_1126,N_1159);
nor U1833 (N_1833,N_1410,N_1481);
and U1834 (N_1834,N_1411,N_1394);
nor U1835 (N_1835,N_1229,N_1245);
nor U1836 (N_1836,N_1038,N_1020);
and U1837 (N_1837,N_1031,N_1454);
or U1838 (N_1838,N_1417,N_1132);
xor U1839 (N_1839,N_1410,N_1110);
and U1840 (N_1840,N_1117,N_1135);
and U1841 (N_1841,N_1466,N_1457);
nor U1842 (N_1842,N_1438,N_1056);
and U1843 (N_1843,N_1269,N_1495);
xnor U1844 (N_1844,N_1484,N_1189);
xnor U1845 (N_1845,N_1146,N_1438);
nand U1846 (N_1846,N_1352,N_1160);
xnor U1847 (N_1847,N_1431,N_1361);
xor U1848 (N_1848,N_1476,N_1156);
xor U1849 (N_1849,N_1015,N_1044);
nor U1850 (N_1850,N_1035,N_1330);
xor U1851 (N_1851,N_1057,N_1161);
nand U1852 (N_1852,N_1443,N_1287);
or U1853 (N_1853,N_1416,N_1034);
xor U1854 (N_1854,N_1279,N_1129);
nand U1855 (N_1855,N_1169,N_1239);
nand U1856 (N_1856,N_1258,N_1291);
nor U1857 (N_1857,N_1205,N_1039);
or U1858 (N_1858,N_1112,N_1160);
nand U1859 (N_1859,N_1123,N_1026);
nand U1860 (N_1860,N_1158,N_1495);
xnor U1861 (N_1861,N_1059,N_1154);
nor U1862 (N_1862,N_1362,N_1057);
and U1863 (N_1863,N_1093,N_1019);
nor U1864 (N_1864,N_1310,N_1134);
and U1865 (N_1865,N_1219,N_1020);
nand U1866 (N_1866,N_1385,N_1190);
nor U1867 (N_1867,N_1199,N_1359);
nor U1868 (N_1868,N_1003,N_1103);
or U1869 (N_1869,N_1257,N_1143);
nand U1870 (N_1870,N_1331,N_1291);
nor U1871 (N_1871,N_1295,N_1358);
nor U1872 (N_1872,N_1425,N_1061);
xnor U1873 (N_1873,N_1088,N_1238);
or U1874 (N_1874,N_1040,N_1108);
xnor U1875 (N_1875,N_1040,N_1121);
or U1876 (N_1876,N_1014,N_1045);
or U1877 (N_1877,N_1159,N_1285);
xnor U1878 (N_1878,N_1413,N_1279);
or U1879 (N_1879,N_1106,N_1228);
nand U1880 (N_1880,N_1310,N_1354);
nor U1881 (N_1881,N_1269,N_1123);
xnor U1882 (N_1882,N_1024,N_1016);
and U1883 (N_1883,N_1215,N_1352);
xnor U1884 (N_1884,N_1265,N_1111);
or U1885 (N_1885,N_1267,N_1155);
and U1886 (N_1886,N_1479,N_1402);
or U1887 (N_1887,N_1331,N_1320);
and U1888 (N_1888,N_1442,N_1419);
xnor U1889 (N_1889,N_1248,N_1487);
nand U1890 (N_1890,N_1072,N_1162);
nand U1891 (N_1891,N_1018,N_1407);
xnor U1892 (N_1892,N_1091,N_1165);
nand U1893 (N_1893,N_1008,N_1177);
xor U1894 (N_1894,N_1088,N_1389);
and U1895 (N_1895,N_1173,N_1038);
nor U1896 (N_1896,N_1383,N_1201);
nor U1897 (N_1897,N_1473,N_1230);
or U1898 (N_1898,N_1232,N_1343);
nand U1899 (N_1899,N_1029,N_1124);
nor U1900 (N_1900,N_1001,N_1117);
or U1901 (N_1901,N_1158,N_1235);
and U1902 (N_1902,N_1032,N_1440);
nor U1903 (N_1903,N_1039,N_1390);
or U1904 (N_1904,N_1277,N_1021);
xor U1905 (N_1905,N_1248,N_1277);
and U1906 (N_1906,N_1496,N_1457);
xnor U1907 (N_1907,N_1040,N_1134);
and U1908 (N_1908,N_1072,N_1105);
nor U1909 (N_1909,N_1185,N_1264);
or U1910 (N_1910,N_1067,N_1061);
nand U1911 (N_1911,N_1157,N_1174);
xor U1912 (N_1912,N_1123,N_1230);
and U1913 (N_1913,N_1452,N_1012);
xor U1914 (N_1914,N_1282,N_1143);
xnor U1915 (N_1915,N_1348,N_1286);
and U1916 (N_1916,N_1413,N_1305);
xor U1917 (N_1917,N_1038,N_1051);
xor U1918 (N_1918,N_1221,N_1208);
nand U1919 (N_1919,N_1322,N_1249);
or U1920 (N_1920,N_1257,N_1431);
and U1921 (N_1921,N_1339,N_1323);
nand U1922 (N_1922,N_1056,N_1388);
nor U1923 (N_1923,N_1226,N_1072);
or U1924 (N_1924,N_1336,N_1256);
nor U1925 (N_1925,N_1246,N_1200);
xnor U1926 (N_1926,N_1253,N_1282);
nor U1927 (N_1927,N_1277,N_1255);
or U1928 (N_1928,N_1296,N_1410);
or U1929 (N_1929,N_1188,N_1181);
or U1930 (N_1930,N_1388,N_1026);
nor U1931 (N_1931,N_1001,N_1371);
nand U1932 (N_1932,N_1373,N_1222);
or U1933 (N_1933,N_1013,N_1024);
or U1934 (N_1934,N_1391,N_1176);
and U1935 (N_1935,N_1418,N_1388);
xor U1936 (N_1936,N_1488,N_1334);
nor U1937 (N_1937,N_1261,N_1380);
xnor U1938 (N_1938,N_1369,N_1485);
xor U1939 (N_1939,N_1464,N_1037);
xnor U1940 (N_1940,N_1162,N_1033);
or U1941 (N_1941,N_1214,N_1293);
or U1942 (N_1942,N_1450,N_1277);
nor U1943 (N_1943,N_1115,N_1089);
xor U1944 (N_1944,N_1150,N_1230);
xor U1945 (N_1945,N_1024,N_1125);
nor U1946 (N_1946,N_1432,N_1161);
and U1947 (N_1947,N_1176,N_1394);
nor U1948 (N_1948,N_1374,N_1254);
nand U1949 (N_1949,N_1455,N_1152);
or U1950 (N_1950,N_1335,N_1426);
nand U1951 (N_1951,N_1185,N_1432);
or U1952 (N_1952,N_1006,N_1397);
nand U1953 (N_1953,N_1078,N_1198);
nor U1954 (N_1954,N_1345,N_1466);
and U1955 (N_1955,N_1224,N_1042);
nor U1956 (N_1956,N_1227,N_1226);
nor U1957 (N_1957,N_1283,N_1168);
nor U1958 (N_1958,N_1110,N_1078);
nand U1959 (N_1959,N_1027,N_1454);
and U1960 (N_1960,N_1210,N_1113);
nor U1961 (N_1961,N_1180,N_1005);
and U1962 (N_1962,N_1007,N_1179);
xnor U1963 (N_1963,N_1439,N_1013);
nand U1964 (N_1964,N_1003,N_1140);
xnor U1965 (N_1965,N_1258,N_1035);
nor U1966 (N_1966,N_1492,N_1341);
xor U1967 (N_1967,N_1434,N_1455);
nand U1968 (N_1968,N_1492,N_1143);
xor U1969 (N_1969,N_1122,N_1367);
and U1970 (N_1970,N_1316,N_1368);
xor U1971 (N_1971,N_1182,N_1289);
or U1972 (N_1972,N_1494,N_1152);
nand U1973 (N_1973,N_1025,N_1122);
nand U1974 (N_1974,N_1059,N_1321);
nand U1975 (N_1975,N_1217,N_1028);
or U1976 (N_1976,N_1242,N_1177);
nand U1977 (N_1977,N_1161,N_1383);
nor U1978 (N_1978,N_1360,N_1117);
nor U1979 (N_1979,N_1093,N_1213);
and U1980 (N_1980,N_1034,N_1436);
and U1981 (N_1981,N_1146,N_1131);
or U1982 (N_1982,N_1359,N_1238);
or U1983 (N_1983,N_1025,N_1398);
xnor U1984 (N_1984,N_1420,N_1448);
nand U1985 (N_1985,N_1077,N_1024);
nor U1986 (N_1986,N_1451,N_1335);
or U1987 (N_1987,N_1481,N_1178);
and U1988 (N_1988,N_1182,N_1417);
or U1989 (N_1989,N_1031,N_1123);
nand U1990 (N_1990,N_1091,N_1318);
or U1991 (N_1991,N_1260,N_1467);
or U1992 (N_1992,N_1351,N_1475);
xor U1993 (N_1993,N_1204,N_1497);
nand U1994 (N_1994,N_1057,N_1354);
nand U1995 (N_1995,N_1245,N_1318);
nand U1996 (N_1996,N_1427,N_1494);
nand U1997 (N_1997,N_1344,N_1086);
nand U1998 (N_1998,N_1458,N_1480);
xor U1999 (N_1999,N_1254,N_1497);
nand U2000 (N_2000,N_1974,N_1944);
nand U2001 (N_2001,N_1768,N_1928);
and U2002 (N_2002,N_1758,N_1842);
and U2003 (N_2003,N_1604,N_1714);
or U2004 (N_2004,N_1733,N_1794);
or U2005 (N_2005,N_1547,N_1700);
nand U2006 (N_2006,N_1906,N_1596);
xnor U2007 (N_2007,N_1601,N_1507);
or U2008 (N_2008,N_1579,N_1615);
and U2009 (N_2009,N_1975,N_1514);
or U2010 (N_2010,N_1911,N_1875);
and U2011 (N_2011,N_1500,N_1959);
and U2012 (N_2012,N_1755,N_1605);
xnor U2013 (N_2013,N_1722,N_1947);
nor U2014 (N_2014,N_1843,N_1982);
and U2015 (N_2015,N_1719,N_1993);
or U2016 (N_2016,N_1820,N_1930);
nor U2017 (N_2017,N_1724,N_1955);
and U2018 (N_2018,N_1771,N_1608);
xor U2019 (N_2019,N_1616,N_1828);
and U2020 (N_2020,N_1582,N_1581);
xnor U2021 (N_2021,N_1584,N_1528);
xor U2022 (N_2022,N_1574,N_1738);
nor U2023 (N_2023,N_1643,N_1648);
and U2024 (N_2024,N_1872,N_1578);
or U2025 (N_2025,N_1512,N_1832);
nand U2026 (N_2026,N_1566,N_1718);
or U2027 (N_2027,N_1545,N_1894);
nor U2028 (N_2028,N_1675,N_1992);
and U2029 (N_2029,N_1709,N_1732);
nor U2030 (N_2030,N_1798,N_1671);
or U2031 (N_2031,N_1573,N_1884);
or U2032 (N_2032,N_1904,N_1531);
xor U2033 (N_2033,N_1867,N_1551);
and U2034 (N_2034,N_1897,N_1589);
xnor U2035 (N_2035,N_1987,N_1864);
and U2036 (N_2036,N_1692,N_1971);
xnor U2037 (N_2037,N_1723,N_1515);
and U2038 (N_2038,N_1857,N_1602);
or U2039 (N_2039,N_1599,N_1854);
xor U2040 (N_2040,N_1552,N_1740);
or U2041 (N_2041,N_1782,N_1815);
xnor U2042 (N_2042,N_1795,N_1681);
and U2043 (N_2043,N_1802,N_1583);
nand U2044 (N_2044,N_1696,N_1543);
xnor U2045 (N_2045,N_1655,N_1684);
nand U2046 (N_2046,N_1770,N_1878);
nor U2047 (N_2047,N_1754,N_1918);
or U2048 (N_2048,N_1970,N_1535);
nand U2049 (N_2049,N_1988,N_1610);
nand U2050 (N_2050,N_1935,N_1707);
or U2051 (N_2051,N_1873,N_1606);
or U2052 (N_2052,N_1699,N_1855);
xnor U2053 (N_2053,N_1949,N_1806);
and U2054 (N_2054,N_1862,N_1640);
xor U2055 (N_2055,N_1533,N_1627);
xor U2056 (N_2056,N_1680,N_1886);
or U2057 (N_2057,N_1939,N_1952);
or U2058 (N_2058,N_1649,N_1711);
or U2059 (N_2059,N_1568,N_1662);
or U2060 (N_2060,N_1563,N_1560);
nand U2061 (N_2061,N_1816,N_1876);
nand U2062 (N_2062,N_1990,N_1863);
xnor U2063 (N_2063,N_1851,N_1837);
or U2064 (N_2064,N_1965,N_1659);
or U2065 (N_2065,N_1529,N_1505);
and U2066 (N_2066,N_1978,N_1669);
and U2067 (N_2067,N_1634,N_1870);
nor U2068 (N_2068,N_1629,N_1916);
and U2069 (N_2069,N_1750,N_1540);
xor U2070 (N_2070,N_1951,N_1565);
nand U2071 (N_2071,N_1549,N_1539);
nand U2072 (N_2072,N_1548,N_1747);
xnor U2073 (N_2073,N_1799,N_1660);
xnor U2074 (N_2074,N_1597,N_1869);
xnor U2075 (N_2075,N_1912,N_1979);
nor U2076 (N_2076,N_1695,N_1541);
or U2077 (N_2077,N_1801,N_1800);
nand U2078 (N_2078,N_1907,N_1923);
or U2079 (N_2079,N_1763,N_1858);
xor U2080 (N_2080,N_1623,N_1729);
nand U2081 (N_2081,N_1698,N_1668);
nor U2082 (N_2082,N_1968,N_1509);
and U2083 (N_2083,N_1829,N_1690);
xor U2084 (N_2084,N_1960,N_1956);
nand U2085 (N_2085,N_1645,N_1778);
xor U2086 (N_2086,N_1663,N_1734);
nor U2087 (N_2087,N_1989,N_1622);
xor U2088 (N_2088,N_1845,N_1553);
nand U2089 (N_2089,N_1950,N_1586);
nor U2090 (N_2090,N_1892,N_1787);
and U2091 (N_2091,N_1694,N_1761);
nand U2092 (N_2092,N_1591,N_1577);
nand U2093 (N_2093,N_1941,N_1967);
or U2094 (N_2094,N_1880,N_1969);
nand U2095 (N_2095,N_1670,N_1929);
xor U2096 (N_2096,N_1716,N_1953);
nor U2097 (N_2097,N_1635,N_1721);
or U2098 (N_2098,N_1691,N_1883);
nor U2099 (N_2099,N_1748,N_1945);
nor U2100 (N_2100,N_1779,N_1926);
nor U2101 (N_2101,N_1677,N_1644);
and U2102 (N_2102,N_1920,N_1785);
xnor U2103 (N_2103,N_1558,N_1784);
xor U2104 (N_2104,N_1847,N_1961);
nor U2105 (N_2105,N_1537,N_1637);
or U2106 (N_2106,N_1585,N_1809);
or U2107 (N_2107,N_1532,N_1713);
nor U2108 (N_2108,N_1885,N_1625);
or U2109 (N_2109,N_1592,N_1527);
or U2110 (N_2110,N_1773,N_1756);
or U2111 (N_2111,N_1933,N_1852);
or U2112 (N_2112,N_1510,N_1877);
or U2113 (N_2113,N_1708,N_1913);
nor U2114 (N_2114,N_1751,N_1501);
nand U2115 (N_2115,N_1924,N_1991);
and U2116 (N_2116,N_1664,N_1697);
nor U2117 (N_2117,N_1818,N_1575);
nand U2118 (N_2118,N_1672,N_1946);
or U2119 (N_2119,N_1521,N_1679);
nor U2120 (N_2120,N_1861,N_1780);
nor U2121 (N_2121,N_1834,N_1922);
xor U2122 (N_2122,N_1827,N_1631);
xor U2123 (N_2123,N_1618,N_1673);
nor U2124 (N_2124,N_1859,N_1735);
or U2125 (N_2125,N_1890,N_1641);
nor U2126 (N_2126,N_1686,N_1749);
nand U2127 (N_2127,N_1972,N_1817);
and U2128 (N_2128,N_1525,N_1665);
and U2129 (N_2129,N_1942,N_1797);
nor U2130 (N_2130,N_1905,N_1737);
and U2131 (N_2131,N_1676,N_1710);
and U2132 (N_2132,N_1588,N_1746);
and U2133 (N_2133,N_1772,N_1628);
or U2134 (N_2134,N_1931,N_1919);
or U2135 (N_2135,N_1638,N_1661);
and U2136 (N_2136,N_1893,N_1726);
nor U2137 (N_2137,N_1976,N_1587);
and U2138 (N_2138,N_1590,N_1594);
nor U2139 (N_2139,N_1874,N_1813);
and U2140 (N_2140,N_1986,N_1717);
nand U2141 (N_2141,N_1511,N_1614);
xnor U2142 (N_2142,N_1682,N_1776);
and U2143 (N_2143,N_1999,N_1788);
or U2144 (N_2144,N_1725,N_1774);
nor U2145 (N_2145,N_1712,N_1745);
or U2146 (N_2146,N_1538,N_1572);
xnor U2147 (N_2147,N_1506,N_1765);
xor U2148 (N_2148,N_1781,N_1825);
nand U2149 (N_2149,N_1998,N_1812);
and U2150 (N_2150,N_1938,N_1838);
and U2151 (N_2151,N_1936,N_1766);
or U2152 (N_2152,N_1612,N_1642);
and U2153 (N_2153,N_1789,N_1569);
nor U2154 (N_2154,N_1567,N_1613);
and U2155 (N_2155,N_1636,N_1657);
nor U2156 (N_2156,N_1977,N_1503);
nand U2157 (N_2157,N_1757,N_1759);
xor U2158 (N_2158,N_1819,N_1792);
xor U2159 (N_2159,N_1621,N_1666);
nand U2160 (N_2160,N_1524,N_1674);
or U2161 (N_2161,N_1775,N_1846);
or U2162 (N_2162,N_1513,N_1542);
xor U2163 (N_2163,N_1849,N_1727);
or U2164 (N_2164,N_1685,N_1767);
or U2165 (N_2165,N_1954,N_1518);
nand U2166 (N_2166,N_1948,N_1925);
nor U2167 (N_2167,N_1814,N_1915);
nor U2168 (N_2168,N_1517,N_1632);
and U2169 (N_2169,N_1791,N_1653);
or U2170 (N_2170,N_1624,N_1887);
and U2171 (N_2171,N_1576,N_1881);
nor U2172 (N_2172,N_1957,N_1804);
nand U2173 (N_2173,N_1561,N_1688);
nand U2174 (N_2174,N_1902,N_1871);
nand U2175 (N_2175,N_1620,N_1562);
and U2176 (N_2176,N_1995,N_1731);
and U2177 (N_2177,N_1609,N_1571);
nand U2178 (N_2178,N_1830,N_1764);
nand U2179 (N_2179,N_1536,N_1652);
and U2180 (N_2180,N_1996,N_1777);
xor U2181 (N_2181,N_1706,N_1811);
xnor U2182 (N_2182,N_1753,N_1654);
nor U2183 (N_2183,N_1580,N_1502);
nor U2184 (N_2184,N_1983,N_1639);
nand U2185 (N_2185,N_1909,N_1557);
xor U2186 (N_2186,N_1667,N_1600);
or U2187 (N_2187,N_1914,N_1937);
nand U2188 (N_2188,N_1530,N_1656);
or U2189 (N_2189,N_1964,N_1522);
xnor U2190 (N_2190,N_1687,N_1651);
and U2191 (N_2191,N_1626,N_1848);
nor U2192 (N_2192,N_1963,N_1921);
nor U2193 (N_2193,N_1683,N_1808);
or U2194 (N_2194,N_1720,N_1833);
or U2195 (N_2195,N_1559,N_1888);
nand U2196 (N_2196,N_1526,N_1554);
xor U2197 (N_2197,N_1895,N_1630);
xor U2198 (N_2198,N_1901,N_1899);
or U2199 (N_2199,N_1927,N_1516);
nor U2200 (N_2200,N_1932,N_1633);
xnor U2201 (N_2201,N_1891,N_1519);
nor U2202 (N_2202,N_1822,N_1715);
or U2203 (N_2203,N_1984,N_1689);
xor U2204 (N_2204,N_1856,N_1985);
and U2205 (N_2205,N_1934,N_1910);
and U2206 (N_2206,N_1744,N_1783);
or U2207 (N_2207,N_1900,N_1742);
or U2208 (N_2208,N_1598,N_1958);
xor U2209 (N_2209,N_1841,N_1940);
nor U2210 (N_2210,N_1619,N_1850);
or U2211 (N_2211,N_1693,N_1807);
xor U2212 (N_2212,N_1823,N_1603);
xor U2213 (N_2213,N_1917,N_1844);
and U2214 (N_2214,N_1981,N_1769);
nor U2215 (N_2215,N_1617,N_1546);
and U2216 (N_2216,N_1550,N_1879);
nor U2217 (N_2217,N_1810,N_1839);
nor U2218 (N_2218,N_1647,N_1865);
nand U2219 (N_2219,N_1728,N_1882);
xor U2220 (N_2220,N_1966,N_1534);
nor U2221 (N_2221,N_1831,N_1860);
and U2222 (N_2222,N_1611,N_1903);
or U2223 (N_2223,N_1824,N_1980);
xnor U2224 (N_2224,N_1973,N_1730);
or U2225 (N_2225,N_1650,N_1835);
and U2226 (N_2226,N_1853,N_1821);
nand U2227 (N_2227,N_1760,N_1703);
xnor U2228 (N_2228,N_1658,N_1504);
xnor U2229 (N_2229,N_1866,N_1908);
or U2230 (N_2230,N_1762,N_1508);
or U2231 (N_2231,N_1646,N_1741);
nor U2232 (N_2232,N_1898,N_1994);
xor U2233 (N_2233,N_1868,N_1826);
nand U2234 (N_2234,N_1796,N_1962);
nand U2235 (N_2235,N_1840,N_1593);
xnor U2236 (N_2236,N_1544,N_1555);
or U2237 (N_2237,N_1889,N_1556);
nor U2238 (N_2238,N_1595,N_1678);
or U2239 (N_2239,N_1607,N_1896);
or U2240 (N_2240,N_1786,N_1997);
and U2241 (N_2241,N_1805,N_1701);
xnor U2242 (N_2242,N_1705,N_1704);
nand U2243 (N_2243,N_1570,N_1790);
and U2244 (N_2244,N_1943,N_1743);
and U2245 (N_2245,N_1836,N_1752);
nand U2246 (N_2246,N_1564,N_1793);
and U2247 (N_2247,N_1523,N_1739);
nand U2248 (N_2248,N_1520,N_1736);
nor U2249 (N_2249,N_1702,N_1803);
or U2250 (N_2250,N_1753,N_1968);
or U2251 (N_2251,N_1770,N_1937);
xnor U2252 (N_2252,N_1857,N_1874);
or U2253 (N_2253,N_1625,N_1584);
xnor U2254 (N_2254,N_1509,N_1738);
xnor U2255 (N_2255,N_1512,N_1989);
nand U2256 (N_2256,N_1543,N_1668);
and U2257 (N_2257,N_1843,N_1730);
xor U2258 (N_2258,N_1513,N_1790);
xor U2259 (N_2259,N_1901,N_1524);
nand U2260 (N_2260,N_1960,N_1579);
nand U2261 (N_2261,N_1884,N_1603);
nand U2262 (N_2262,N_1531,N_1597);
and U2263 (N_2263,N_1698,N_1851);
xor U2264 (N_2264,N_1884,N_1781);
and U2265 (N_2265,N_1579,N_1770);
or U2266 (N_2266,N_1862,N_1722);
or U2267 (N_2267,N_1861,N_1996);
nand U2268 (N_2268,N_1610,N_1690);
and U2269 (N_2269,N_1586,N_1547);
xnor U2270 (N_2270,N_1717,N_1545);
or U2271 (N_2271,N_1563,N_1741);
xor U2272 (N_2272,N_1769,N_1797);
or U2273 (N_2273,N_1521,N_1524);
and U2274 (N_2274,N_1529,N_1614);
nor U2275 (N_2275,N_1867,N_1896);
nand U2276 (N_2276,N_1723,N_1629);
or U2277 (N_2277,N_1608,N_1607);
or U2278 (N_2278,N_1827,N_1898);
xor U2279 (N_2279,N_1810,N_1851);
and U2280 (N_2280,N_1782,N_1786);
xor U2281 (N_2281,N_1591,N_1629);
xnor U2282 (N_2282,N_1607,N_1690);
nor U2283 (N_2283,N_1943,N_1800);
or U2284 (N_2284,N_1767,N_1662);
nand U2285 (N_2285,N_1852,N_1795);
xnor U2286 (N_2286,N_1701,N_1540);
nor U2287 (N_2287,N_1652,N_1834);
and U2288 (N_2288,N_1853,N_1671);
or U2289 (N_2289,N_1503,N_1608);
xnor U2290 (N_2290,N_1616,N_1818);
and U2291 (N_2291,N_1876,N_1693);
nand U2292 (N_2292,N_1713,N_1682);
or U2293 (N_2293,N_1609,N_1520);
xnor U2294 (N_2294,N_1572,N_1819);
nor U2295 (N_2295,N_1708,N_1594);
nor U2296 (N_2296,N_1694,N_1601);
or U2297 (N_2297,N_1786,N_1573);
and U2298 (N_2298,N_1993,N_1877);
nand U2299 (N_2299,N_1611,N_1745);
nand U2300 (N_2300,N_1998,N_1944);
and U2301 (N_2301,N_1655,N_1895);
or U2302 (N_2302,N_1549,N_1869);
nor U2303 (N_2303,N_1549,N_1799);
xor U2304 (N_2304,N_1788,N_1654);
or U2305 (N_2305,N_1929,N_1824);
and U2306 (N_2306,N_1759,N_1780);
nor U2307 (N_2307,N_1550,N_1555);
xnor U2308 (N_2308,N_1995,N_1508);
xnor U2309 (N_2309,N_1812,N_1623);
xnor U2310 (N_2310,N_1804,N_1781);
nor U2311 (N_2311,N_1748,N_1734);
nor U2312 (N_2312,N_1918,N_1766);
nor U2313 (N_2313,N_1986,N_1958);
nor U2314 (N_2314,N_1773,N_1870);
nand U2315 (N_2315,N_1980,N_1806);
nand U2316 (N_2316,N_1777,N_1893);
and U2317 (N_2317,N_1820,N_1846);
and U2318 (N_2318,N_1854,N_1774);
nor U2319 (N_2319,N_1500,N_1798);
and U2320 (N_2320,N_1600,N_1609);
and U2321 (N_2321,N_1888,N_1718);
nor U2322 (N_2322,N_1742,N_1925);
and U2323 (N_2323,N_1654,N_1527);
nor U2324 (N_2324,N_1875,N_1855);
and U2325 (N_2325,N_1607,N_1732);
or U2326 (N_2326,N_1597,N_1522);
nand U2327 (N_2327,N_1857,N_1876);
xnor U2328 (N_2328,N_1891,N_1919);
or U2329 (N_2329,N_1650,N_1812);
nor U2330 (N_2330,N_1574,N_1946);
nand U2331 (N_2331,N_1821,N_1543);
nor U2332 (N_2332,N_1863,N_1882);
xor U2333 (N_2333,N_1705,N_1917);
or U2334 (N_2334,N_1750,N_1820);
nor U2335 (N_2335,N_1722,N_1769);
xor U2336 (N_2336,N_1658,N_1970);
nor U2337 (N_2337,N_1664,N_1626);
or U2338 (N_2338,N_1871,N_1866);
and U2339 (N_2339,N_1945,N_1534);
xnor U2340 (N_2340,N_1535,N_1548);
or U2341 (N_2341,N_1532,N_1756);
and U2342 (N_2342,N_1965,N_1535);
nor U2343 (N_2343,N_1591,N_1936);
nor U2344 (N_2344,N_1779,N_1716);
xor U2345 (N_2345,N_1659,N_1784);
and U2346 (N_2346,N_1791,N_1762);
nor U2347 (N_2347,N_1866,N_1957);
or U2348 (N_2348,N_1502,N_1747);
nand U2349 (N_2349,N_1745,N_1987);
xnor U2350 (N_2350,N_1509,N_1690);
nor U2351 (N_2351,N_1561,N_1880);
or U2352 (N_2352,N_1829,N_1889);
or U2353 (N_2353,N_1955,N_1878);
and U2354 (N_2354,N_1871,N_1933);
and U2355 (N_2355,N_1852,N_1579);
and U2356 (N_2356,N_1635,N_1997);
xor U2357 (N_2357,N_1962,N_1770);
or U2358 (N_2358,N_1601,N_1653);
or U2359 (N_2359,N_1870,N_1735);
nor U2360 (N_2360,N_1607,N_1908);
and U2361 (N_2361,N_1934,N_1889);
nand U2362 (N_2362,N_1842,N_1651);
nand U2363 (N_2363,N_1570,N_1520);
xnor U2364 (N_2364,N_1952,N_1812);
nor U2365 (N_2365,N_1653,N_1647);
nand U2366 (N_2366,N_1551,N_1652);
nor U2367 (N_2367,N_1931,N_1656);
nor U2368 (N_2368,N_1575,N_1988);
nand U2369 (N_2369,N_1658,N_1761);
xnor U2370 (N_2370,N_1996,N_1779);
or U2371 (N_2371,N_1505,N_1510);
xor U2372 (N_2372,N_1676,N_1818);
and U2373 (N_2373,N_1563,N_1957);
nor U2374 (N_2374,N_1641,N_1638);
or U2375 (N_2375,N_1526,N_1650);
nand U2376 (N_2376,N_1778,N_1913);
and U2377 (N_2377,N_1757,N_1534);
and U2378 (N_2378,N_1622,N_1781);
or U2379 (N_2379,N_1578,N_1771);
nor U2380 (N_2380,N_1525,N_1983);
or U2381 (N_2381,N_1715,N_1783);
xnor U2382 (N_2382,N_1955,N_1995);
and U2383 (N_2383,N_1531,N_1952);
and U2384 (N_2384,N_1974,N_1953);
or U2385 (N_2385,N_1818,N_1990);
or U2386 (N_2386,N_1680,N_1810);
nor U2387 (N_2387,N_1921,N_1717);
and U2388 (N_2388,N_1944,N_1513);
nor U2389 (N_2389,N_1859,N_1633);
nand U2390 (N_2390,N_1694,N_1581);
and U2391 (N_2391,N_1634,N_1525);
nor U2392 (N_2392,N_1789,N_1972);
xnor U2393 (N_2393,N_1842,N_1686);
nor U2394 (N_2394,N_1524,N_1615);
nor U2395 (N_2395,N_1658,N_1732);
or U2396 (N_2396,N_1569,N_1594);
nor U2397 (N_2397,N_1510,N_1850);
and U2398 (N_2398,N_1709,N_1692);
and U2399 (N_2399,N_1706,N_1976);
or U2400 (N_2400,N_1966,N_1911);
nor U2401 (N_2401,N_1884,N_1893);
and U2402 (N_2402,N_1774,N_1557);
and U2403 (N_2403,N_1667,N_1889);
nand U2404 (N_2404,N_1903,N_1853);
nand U2405 (N_2405,N_1544,N_1923);
nand U2406 (N_2406,N_1514,N_1919);
or U2407 (N_2407,N_1692,N_1768);
xnor U2408 (N_2408,N_1845,N_1523);
nand U2409 (N_2409,N_1801,N_1700);
or U2410 (N_2410,N_1863,N_1870);
and U2411 (N_2411,N_1859,N_1522);
or U2412 (N_2412,N_1721,N_1886);
or U2413 (N_2413,N_1947,N_1672);
xnor U2414 (N_2414,N_1547,N_1944);
nor U2415 (N_2415,N_1884,N_1840);
nor U2416 (N_2416,N_1591,N_1599);
or U2417 (N_2417,N_1526,N_1904);
or U2418 (N_2418,N_1705,N_1646);
nand U2419 (N_2419,N_1943,N_1787);
and U2420 (N_2420,N_1883,N_1748);
and U2421 (N_2421,N_1964,N_1754);
xnor U2422 (N_2422,N_1905,N_1694);
xor U2423 (N_2423,N_1776,N_1794);
or U2424 (N_2424,N_1826,N_1836);
and U2425 (N_2425,N_1600,N_1970);
xnor U2426 (N_2426,N_1573,N_1844);
and U2427 (N_2427,N_1592,N_1735);
and U2428 (N_2428,N_1972,N_1941);
nor U2429 (N_2429,N_1897,N_1776);
nor U2430 (N_2430,N_1918,N_1844);
xnor U2431 (N_2431,N_1899,N_1514);
nor U2432 (N_2432,N_1585,N_1656);
or U2433 (N_2433,N_1689,N_1566);
xnor U2434 (N_2434,N_1971,N_1710);
or U2435 (N_2435,N_1581,N_1781);
nor U2436 (N_2436,N_1717,N_1605);
or U2437 (N_2437,N_1556,N_1758);
nor U2438 (N_2438,N_1960,N_1742);
and U2439 (N_2439,N_1935,N_1516);
xnor U2440 (N_2440,N_1980,N_1804);
nand U2441 (N_2441,N_1557,N_1824);
xor U2442 (N_2442,N_1557,N_1706);
nor U2443 (N_2443,N_1717,N_1681);
nand U2444 (N_2444,N_1640,N_1879);
or U2445 (N_2445,N_1528,N_1738);
xnor U2446 (N_2446,N_1741,N_1880);
xor U2447 (N_2447,N_1986,N_1881);
nand U2448 (N_2448,N_1852,N_1934);
xor U2449 (N_2449,N_1614,N_1863);
nand U2450 (N_2450,N_1904,N_1903);
and U2451 (N_2451,N_1989,N_1927);
nor U2452 (N_2452,N_1784,N_1941);
xnor U2453 (N_2453,N_1640,N_1641);
nand U2454 (N_2454,N_1818,N_1908);
and U2455 (N_2455,N_1981,N_1714);
and U2456 (N_2456,N_1858,N_1535);
nand U2457 (N_2457,N_1795,N_1776);
nor U2458 (N_2458,N_1546,N_1649);
and U2459 (N_2459,N_1951,N_1959);
xnor U2460 (N_2460,N_1531,N_1828);
and U2461 (N_2461,N_1928,N_1807);
xnor U2462 (N_2462,N_1744,N_1580);
nand U2463 (N_2463,N_1977,N_1972);
or U2464 (N_2464,N_1949,N_1698);
or U2465 (N_2465,N_1541,N_1954);
or U2466 (N_2466,N_1810,N_1620);
or U2467 (N_2467,N_1828,N_1835);
nor U2468 (N_2468,N_1660,N_1676);
and U2469 (N_2469,N_1529,N_1849);
nor U2470 (N_2470,N_1665,N_1567);
nor U2471 (N_2471,N_1789,N_1905);
and U2472 (N_2472,N_1511,N_1549);
xor U2473 (N_2473,N_1863,N_1891);
nand U2474 (N_2474,N_1930,N_1830);
and U2475 (N_2475,N_1785,N_1571);
nor U2476 (N_2476,N_1816,N_1964);
or U2477 (N_2477,N_1696,N_1787);
xnor U2478 (N_2478,N_1963,N_1741);
or U2479 (N_2479,N_1859,N_1585);
xnor U2480 (N_2480,N_1547,N_1953);
and U2481 (N_2481,N_1544,N_1530);
xor U2482 (N_2482,N_1832,N_1967);
nor U2483 (N_2483,N_1929,N_1844);
xor U2484 (N_2484,N_1880,N_1709);
or U2485 (N_2485,N_1584,N_1596);
nor U2486 (N_2486,N_1633,N_1896);
xor U2487 (N_2487,N_1884,N_1887);
or U2488 (N_2488,N_1842,N_1601);
and U2489 (N_2489,N_1534,N_1575);
nor U2490 (N_2490,N_1616,N_1640);
nand U2491 (N_2491,N_1720,N_1526);
xor U2492 (N_2492,N_1917,N_1873);
xor U2493 (N_2493,N_1543,N_1990);
nand U2494 (N_2494,N_1999,N_1820);
nor U2495 (N_2495,N_1633,N_1892);
or U2496 (N_2496,N_1597,N_1549);
xnor U2497 (N_2497,N_1871,N_1982);
nor U2498 (N_2498,N_1951,N_1646);
and U2499 (N_2499,N_1727,N_1819);
or U2500 (N_2500,N_2420,N_2382);
nand U2501 (N_2501,N_2256,N_2439);
nor U2502 (N_2502,N_2099,N_2298);
xnor U2503 (N_2503,N_2111,N_2491);
or U2504 (N_2504,N_2026,N_2338);
nor U2505 (N_2505,N_2047,N_2407);
xor U2506 (N_2506,N_2335,N_2159);
xnor U2507 (N_2507,N_2147,N_2363);
xor U2508 (N_2508,N_2336,N_2202);
nor U2509 (N_2509,N_2135,N_2480);
xor U2510 (N_2510,N_2218,N_2304);
and U2511 (N_2511,N_2217,N_2090);
and U2512 (N_2512,N_2376,N_2467);
or U2513 (N_2513,N_2284,N_2232);
xor U2514 (N_2514,N_2416,N_2456);
and U2515 (N_2515,N_2316,N_2007);
and U2516 (N_2516,N_2216,N_2380);
nand U2517 (N_2517,N_2487,N_2044);
and U2518 (N_2518,N_2103,N_2091);
nor U2519 (N_2519,N_2200,N_2072);
or U2520 (N_2520,N_2328,N_2124);
or U2521 (N_2521,N_2411,N_2194);
or U2522 (N_2522,N_2449,N_2378);
nand U2523 (N_2523,N_2285,N_2349);
xor U2524 (N_2524,N_2353,N_2027);
or U2525 (N_2525,N_2471,N_2119);
and U2526 (N_2526,N_2485,N_2224);
nand U2527 (N_2527,N_2451,N_2190);
and U2528 (N_2528,N_2136,N_2122);
and U2529 (N_2529,N_2412,N_2023);
nand U2530 (N_2530,N_2199,N_2259);
and U2531 (N_2531,N_2235,N_2362);
or U2532 (N_2532,N_2141,N_2022);
and U2533 (N_2533,N_2277,N_2418);
nor U2534 (N_2534,N_2292,N_2038);
xnor U2535 (N_2535,N_2080,N_2071);
xnor U2536 (N_2536,N_2058,N_2461);
nor U2537 (N_2537,N_2050,N_2036);
or U2538 (N_2538,N_2230,N_2064);
and U2539 (N_2539,N_2466,N_2358);
nand U2540 (N_2540,N_2400,N_2186);
and U2541 (N_2541,N_2178,N_2000);
nor U2542 (N_2542,N_2372,N_2245);
and U2543 (N_2543,N_2315,N_2016);
nor U2544 (N_2544,N_2265,N_2401);
and U2545 (N_2545,N_2383,N_2484);
xnor U2546 (N_2546,N_2116,N_2436);
nand U2547 (N_2547,N_2289,N_2323);
or U2548 (N_2548,N_2348,N_2029);
xnor U2549 (N_2549,N_2221,N_2121);
nand U2550 (N_2550,N_2215,N_2396);
and U2551 (N_2551,N_2322,N_2021);
and U2552 (N_2552,N_2425,N_2214);
or U2553 (N_2553,N_2492,N_2053);
or U2554 (N_2554,N_2048,N_2426);
nor U2555 (N_2555,N_2321,N_2477);
xor U2556 (N_2556,N_2301,N_2033);
xnor U2557 (N_2557,N_2414,N_2249);
xnor U2558 (N_2558,N_2431,N_2138);
xor U2559 (N_2559,N_2435,N_2389);
or U2560 (N_2560,N_2294,N_2248);
nor U2561 (N_2561,N_2433,N_2197);
xnor U2562 (N_2562,N_2409,N_2052);
or U2563 (N_2563,N_2127,N_2102);
and U2564 (N_2564,N_2094,N_2476);
xor U2565 (N_2565,N_2278,N_2276);
xnor U2566 (N_2566,N_2137,N_2337);
or U2567 (N_2567,N_2191,N_2165);
nand U2568 (N_2568,N_2281,N_2454);
and U2569 (N_2569,N_2092,N_2062);
nand U2570 (N_2570,N_2231,N_2371);
and U2571 (N_2571,N_2143,N_2089);
or U2572 (N_2572,N_2262,N_2464);
nor U2573 (N_2573,N_2452,N_2209);
xnor U2574 (N_2574,N_2307,N_2297);
or U2575 (N_2575,N_2341,N_2188);
xor U2576 (N_2576,N_2360,N_2157);
xnor U2577 (N_2577,N_2192,N_2057);
nor U2578 (N_2578,N_2446,N_2145);
xnor U2579 (N_2579,N_2126,N_2160);
xnor U2580 (N_2580,N_2210,N_2242);
and U2581 (N_2581,N_2074,N_2282);
nand U2582 (N_2582,N_2110,N_2101);
and U2583 (N_2583,N_2437,N_2238);
xnor U2584 (N_2584,N_2302,N_2333);
nand U2585 (N_2585,N_2253,N_2104);
nor U2586 (N_2586,N_2331,N_2151);
nand U2587 (N_2587,N_2076,N_2049);
xor U2588 (N_2588,N_2004,N_2061);
nor U2589 (N_2589,N_2489,N_2447);
xnor U2590 (N_2590,N_2299,N_2334);
and U2591 (N_2591,N_2014,N_2370);
nor U2592 (N_2592,N_2406,N_2403);
nand U2593 (N_2593,N_2324,N_2228);
nor U2594 (N_2594,N_2320,N_2252);
nor U2595 (N_2595,N_2070,N_2394);
xor U2596 (N_2596,N_2329,N_2438);
or U2597 (N_2597,N_2390,N_2077);
nor U2598 (N_2598,N_2035,N_2402);
and U2599 (N_2599,N_2114,N_2379);
xor U2600 (N_2600,N_2440,N_2313);
or U2601 (N_2601,N_2069,N_2280);
nand U2602 (N_2602,N_2481,N_2240);
nand U2603 (N_2603,N_2486,N_2196);
nand U2604 (N_2604,N_2012,N_2290);
xor U2605 (N_2605,N_2266,N_2010);
and U2606 (N_2606,N_2375,N_2120);
xnor U2607 (N_2607,N_2352,N_2171);
xnor U2608 (N_2608,N_2041,N_2312);
nand U2609 (N_2609,N_2350,N_2330);
nor U2610 (N_2610,N_2434,N_2208);
nand U2611 (N_2611,N_2155,N_2493);
nor U2612 (N_2612,N_2028,N_2172);
nor U2613 (N_2613,N_2270,N_2150);
nor U2614 (N_2614,N_2325,N_2180);
and U2615 (N_2615,N_2462,N_2239);
and U2616 (N_2616,N_2459,N_2195);
or U2617 (N_2617,N_2243,N_2156);
and U2618 (N_2618,N_2413,N_2347);
and U2619 (N_2619,N_2332,N_2293);
xnor U2620 (N_2620,N_2123,N_2204);
and U2621 (N_2621,N_2494,N_2129);
nor U2622 (N_2622,N_2223,N_2274);
nand U2623 (N_2623,N_2286,N_2109);
xnor U2624 (N_2624,N_2475,N_2001);
nor U2625 (N_2625,N_2220,N_2490);
nand U2626 (N_2626,N_2246,N_2343);
nor U2627 (N_2627,N_2306,N_2113);
and U2628 (N_2628,N_2055,N_2042);
nor U2629 (N_2629,N_2257,N_2258);
nand U2630 (N_2630,N_2283,N_2139);
nor U2631 (N_2631,N_2065,N_2279);
and U2632 (N_2632,N_2152,N_2233);
or U2633 (N_2633,N_2189,N_2067);
and U2634 (N_2634,N_2496,N_2162);
and U2635 (N_2635,N_2020,N_2305);
or U2636 (N_2636,N_2309,N_2207);
and U2637 (N_2637,N_2032,N_2193);
xor U2638 (N_2638,N_2128,N_2002);
and U2639 (N_2639,N_2013,N_2039);
and U2640 (N_2640,N_2388,N_2166);
and U2641 (N_2641,N_2268,N_2263);
nor U2642 (N_2642,N_2345,N_2030);
nand U2643 (N_2643,N_2460,N_2131);
xnor U2644 (N_2644,N_2125,N_2455);
or U2645 (N_2645,N_2408,N_2497);
xnor U2646 (N_2646,N_2018,N_2108);
xnor U2647 (N_2647,N_2140,N_2154);
nand U2648 (N_2648,N_2198,N_2112);
nor U2649 (N_2649,N_2359,N_2219);
or U2650 (N_2650,N_2398,N_2317);
xnor U2651 (N_2651,N_2469,N_2222);
and U2652 (N_2652,N_2167,N_2149);
and U2653 (N_2653,N_2450,N_2342);
xnor U2654 (N_2654,N_2424,N_2303);
nand U2655 (N_2655,N_2133,N_2097);
or U2656 (N_2656,N_2176,N_2213);
nor U2657 (N_2657,N_2373,N_2339);
or U2658 (N_2658,N_2311,N_2254);
nand U2659 (N_2659,N_2374,N_2478);
nor U2660 (N_2660,N_2326,N_2273);
and U2661 (N_2661,N_2444,N_2272);
xnor U2662 (N_2662,N_2314,N_2310);
and U2663 (N_2663,N_2095,N_2499);
nand U2664 (N_2664,N_2453,N_2443);
or U2665 (N_2665,N_2083,N_2264);
nor U2666 (N_2666,N_2073,N_2115);
nor U2667 (N_2667,N_2244,N_2473);
and U2668 (N_2668,N_2153,N_2184);
xnor U2669 (N_2669,N_2146,N_2463);
nand U2670 (N_2670,N_2054,N_2130);
and U2671 (N_2671,N_2170,N_2386);
nor U2672 (N_2672,N_2185,N_2479);
nor U2673 (N_2673,N_2361,N_2287);
or U2674 (N_2674,N_2187,N_2367);
nor U2675 (N_2675,N_2488,N_2066);
or U2676 (N_2676,N_2393,N_2237);
nor U2677 (N_2677,N_2148,N_2368);
xnor U2678 (N_2678,N_2106,N_2031);
nor U2679 (N_2679,N_2037,N_2465);
nand U2680 (N_2680,N_2483,N_2419);
xnor U2681 (N_2681,N_2201,N_2441);
xor U2682 (N_2682,N_2005,N_2346);
nor U2683 (N_2683,N_2043,N_2107);
and U2684 (N_2684,N_2340,N_2397);
and U2685 (N_2685,N_2024,N_2075);
nor U2686 (N_2686,N_2288,N_2079);
and U2687 (N_2687,N_2399,N_2429);
nor U2688 (N_2688,N_2236,N_2448);
nand U2689 (N_2689,N_2025,N_2247);
xor U2690 (N_2690,N_2051,N_2096);
xnor U2691 (N_2691,N_2468,N_2100);
nand U2692 (N_2692,N_2181,N_2445);
nor U2693 (N_2693,N_2161,N_2269);
or U2694 (N_2694,N_2430,N_2060);
nand U2695 (N_2695,N_2068,N_2255);
nor U2696 (N_2696,N_2175,N_2087);
or U2697 (N_2697,N_2319,N_2251);
nand U2698 (N_2698,N_2117,N_2495);
and U2699 (N_2699,N_2387,N_2144);
xnor U2700 (N_2700,N_2212,N_2019);
nor U2701 (N_2701,N_2011,N_2085);
nand U2702 (N_2702,N_2470,N_2300);
and U2703 (N_2703,N_2275,N_2142);
xor U2704 (N_2704,N_2006,N_2369);
or U2705 (N_2705,N_2169,N_2182);
or U2706 (N_2706,N_2250,N_2098);
nand U2707 (N_2707,N_2017,N_2134);
and U2708 (N_2708,N_2009,N_2457);
or U2709 (N_2709,N_2183,N_2498);
or U2710 (N_2710,N_2211,N_2405);
nor U2711 (N_2711,N_2410,N_2357);
and U2712 (N_2712,N_2327,N_2179);
nand U2713 (N_2713,N_2442,N_2234);
nand U2714 (N_2714,N_2040,N_2415);
nand U2715 (N_2715,N_2428,N_2088);
or U2716 (N_2716,N_2295,N_2105);
nor U2717 (N_2717,N_2391,N_2356);
nand U2718 (N_2718,N_2260,N_2422);
and U2719 (N_2719,N_2404,N_2377);
nand U2720 (N_2720,N_2417,N_2432);
or U2721 (N_2721,N_2177,N_2059);
nand U2722 (N_2722,N_2308,N_2366);
xnor U2723 (N_2723,N_2226,N_2427);
or U2724 (N_2724,N_2034,N_2365);
and U2725 (N_2725,N_2385,N_2351);
nand U2726 (N_2726,N_2164,N_2227);
nand U2727 (N_2727,N_2173,N_2163);
nand U2728 (N_2728,N_2271,N_2364);
nand U2729 (N_2729,N_2384,N_2081);
nand U2730 (N_2730,N_2086,N_2132);
and U2731 (N_2731,N_2206,N_2296);
and U2732 (N_2732,N_2056,N_2158);
and U2733 (N_2733,N_2003,N_2118);
nand U2734 (N_2734,N_2472,N_2291);
nor U2735 (N_2735,N_2241,N_2225);
xnor U2736 (N_2736,N_2395,N_2093);
or U2737 (N_2737,N_2015,N_2168);
nor U2738 (N_2738,N_2423,N_2229);
xor U2739 (N_2739,N_2355,N_2392);
or U2740 (N_2740,N_2174,N_2205);
nor U2741 (N_2741,N_2046,N_2318);
nand U2742 (N_2742,N_2261,N_2008);
xor U2743 (N_2743,N_2421,N_2084);
nand U2744 (N_2744,N_2482,N_2063);
xor U2745 (N_2745,N_2458,N_2474);
nand U2746 (N_2746,N_2203,N_2344);
xor U2747 (N_2747,N_2082,N_2354);
nor U2748 (N_2748,N_2045,N_2381);
or U2749 (N_2749,N_2267,N_2078);
nand U2750 (N_2750,N_2178,N_2391);
xor U2751 (N_2751,N_2263,N_2434);
or U2752 (N_2752,N_2033,N_2351);
and U2753 (N_2753,N_2024,N_2334);
nor U2754 (N_2754,N_2234,N_2406);
nor U2755 (N_2755,N_2323,N_2163);
xor U2756 (N_2756,N_2021,N_2295);
or U2757 (N_2757,N_2262,N_2156);
or U2758 (N_2758,N_2117,N_2366);
and U2759 (N_2759,N_2197,N_2066);
nor U2760 (N_2760,N_2026,N_2325);
or U2761 (N_2761,N_2122,N_2499);
or U2762 (N_2762,N_2460,N_2165);
xor U2763 (N_2763,N_2210,N_2159);
and U2764 (N_2764,N_2499,N_2129);
nand U2765 (N_2765,N_2473,N_2030);
nand U2766 (N_2766,N_2137,N_2261);
nand U2767 (N_2767,N_2116,N_2322);
nor U2768 (N_2768,N_2421,N_2311);
xnor U2769 (N_2769,N_2086,N_2346);
nand U2770 (N_2770,N_2150,N_2235);
or U2771 (N_2771,N_2220,N_2181);
nor U2772 (N_2772,N_2423,N_2166);
or U2773 (N_2773,N_2184,N_2302);
xor U2774 (N_2774,N_2106,N_2128);
nor U2775 (N_2775,N_2097,N_2241);
xor U2776 (N_2776,N_2076,N_2066);
and U2777 (N_2777,N_2311,N_2164);
xor U2778 (N_2778,N_2096,N_2252);
nor U2779 (N_2779,N_2236,N_2461);
or U2780 (N_2780,N_2140,N_2278);
and U2781 (N_2781,N_2140,N_2064);
and U2782 (N_2782,N_2386,N_2069);
or U2783 (N_2783,N_2136,N_2263);
nor U2784 (N_2784,N_2337,N_2202);
nand U2785 (N_2785,N_2016,N_2266);
or U2786 (N_2786,N_2144,N_2147);
nor U2787 (N_2787,N_2097,N_2319);
xnor U2788 (N_2788,N_2215,N_2430);
xnor U2789 (N_2789,N_2253,N_2147);
and U2790 (N_2790,N_2435,N_2023);
and U2791 (N_2791,N_2321,N_2156);
and U2792 (N_2792,N_2298,N_2414);
xnor U2793 (N_2793,N_2256,N_2436);
nand U2794 (N_2794,N_2157,N_2213);
xnor U2795 (N_2795,N_2436,N_2327);
nand U2796 (N_2796,N_2388,N_2037);
or U2797 (N_2797,N_2228,N_2497);
nand U2798 (N_2798,N_2199,N_2446);
xor U2799 (N_2799,N_2152,N_2497);
or U2800 (N_2800,N_2203,N_2184);
xnor U2801 (N_2801,N_2372,N_2142);
nand U2802 (N_2802,N_2498,N_2210);
xor U2803 (N_2803,N_2252,N_2219);
xor U2804 (N_2804,N_2102,N_2115);
nor U2805 (N_2805,N_2077,N_2071);
nor U2806 (N_2806,N_2384,N_2412);
xor U2807 (N_2807,N_2283,N_2069);
or U2808 (N_2808,N_2219,N_2212);
nor U2809 (N_2809,N_2446,N_2172);
and U2810 (N_2810,N_2483,N_2339);
and U2811 (N_2811,N_2044,N_2238);
and U2812 (N_2812,N_2048,N_2265);
nor U2813 (N_2813,N_2166,N_2259);
xor U2814 (N_2814,N_2159,N_2144);
and U2815 (N_2815,N_2266,N_2111);
or U2816 (N_2816,N_2423,N_2227);
and U2817 (N_2817,N_2285,N_2037);
and U2818 (N_2818,N_2445,N_2015);
or U2819 (N_2819,N_2492,N_2340);
or U2820 (N_2820,N_2336,N_2411);
nor U2821 (N_2821,N_2048,N_2299);
xnor U2822 (N_2822,N_2234,N_2451);
xor U2823 (N_2823,N_2036,N_2340);
nand U2824 (N_2824,N_2386,N_2262);
xnor U2825 (N_2825,N_2007,N_2169);
or U2826 (N_2826,N_2217,N_2283);
and U2827 (N_2827,N_2285,N_2154);
nor U2828 (N_2828,N_2476,N_2331);
or U2829 (N_2829,N_2018,N_2138);
nor U2830 (N_2830,N_2395,N_2074);
or U2831 (N_2831,N_2414,N_2120);
nor U2832 (N_2832,N_2067,N_2287);
xor U2833 (N_2833,N_2275,N_2199);
xor U2834 (N_2834,N_2480,N_2171);
nand U2835 (N_2835,N_2045,N_2430);
nand U2836 (N_2836,N_2499,N_2353);
xnor U2837 (N_2837,N_2009,N_2212);
or U2838 (N_2838,N_2318,N_2282);
xnor U2839 (N_2839,N_2248,N_2180);
or U2840 (N_2840,N_2389,N_2029);
and U2841 (N_2841,N_2403,N_2221);
and U2842 (N_2842,N_2221,N_2198);
xnor U2843 (N_2843,N_2154,N_2249);
xor U2844 (N_2844,N_2065,N_2357);
xor U2845 (N_2845,N_2311,N_2093);
and U2846 (N_2846,N_2326,N_2434);
and U2847 (N_2847,N_2111,N_2367);
nor U2848 (N_2848,N_2201,N_2071);
xor U2849 (N_2849,N_2451,N_2345);
nand U2850 (N_2850,N_2499,N_2264);
xor U2851 (N_2851,N_2345,N_2224);
nand U2852 (N_2852,N_2044,N_2351);
nor U2853 (N_2853,N_2275,N_2229);
nor U2854 (N_2854,N_2110,N_2220);
nand U2855 (N_2855,N_2291,N_2461);
and U2856 (N_2856,N_2393,N_2432);
nand U2857 (N_2857,N_2039,N_2238);
nand U2858 (N_2858,N_2311,N_2430);
or U2859 (N_2859,N_2328,N_2337);
nor U2860 (N_2860,N_2035,N_2328);
nand U2861 (N_2861,N_2409,N_2160);
nand U2862 (N_2862,N_2258,N_2025);
and U2863 (N_2863,N_2287,N_2248);
xor U2864 (N_2864,N_2247,N_2411);
xor U2865 (N_2865,N_2041,N_2286);
xnor U2866 (N_2866,N_2091,N_2139);
and U2867 (N_2867,N_2383,N_2397);
nor U2868 (N_2868,N_2096,N_2300);
nand U2869 (N_2869,N_2222,N_2288);
and U2870 (N_2870,N_2096,N_2254);
or U2871 (N_2871,N_2491,N_2479);
and U2872 (N_2872,N_2094,N_2149);
xnor U2873 (N_2873,N_2129,N_2029);
or U2874 (N_2874,N_2105,N_2141);
nand U2875 (N_2875,N_2350,N_2041);
xor U2876 (N_2876,N_2105,N_2171);
and U2877 (N_2877,N_2432,N_2130);
and U2878 (N_2878,N_2144,N_2253);
and U2879 (N_2879,N_2281,N_2245);
nor U2880 (N_2880,N_2334,N_2336);
nor U2881 (N_2881,N_2494,N_2092);
nor U2882 (N_2882,N_2155,N_2093);
nor U2883 (N_2883,N_2012,N_2417);
or U2884 (N_2884,N_2361,N_2436);
nor U2885 (N_2885,N_2291,N_2139);
and U2886 (N_2886,N_2378,N_2154);
and U2887 (N_2887,N_2018,N_2374);
nand U2888 (N_2888,N_2306,N_2470);
or U2889 (N_2889,N_2138,N_2042);
and U2890 (N_2890,N_2195,N_2441);
or U2891 (N_2891,N_2143,N_2153);
nand U2892 (N_2892,N_2236,N_2490);
or U2893 (N_2893,N_2492,N_2360);
xnor U2894 (N_2894,N_2491,N_2431);
nand U2895 (N_2895,N_2326,N_2130);
and U2896 (N_2896,N_2243,N_2047);
or U2897 (N_2897,N_2045,N_2297);
and U2898 (N_2898,N_2184,N_2011);
and U2899 (N_2899,N_2097,N_2277);
nor U2900 (N_2900,N_2418,N_2414);
nand U2901 (N_2901,N_2363,N_2197);
and U2902 (N_2902,N_2490,N_2347);
nor U2903 (N_2903,N_2224,N_2292);
xnor U2904 (N_2904,N_2244,N_2145);
nand U2905 (N_2905,N_2293,N_2394);
nand U2906 (N_2906,N_2393,N_2363);
and U2907 (N_2907,N_2164,N_2369);
and U2908 (N_2908,N_2480,N_2369);
or U2909 (N_2909,N_2244,N_2222);
xnor U2910 (N_2910,N_2145,N_2197);
and U2911 (N_2911,N_2354,N_2249);
or U2912 (N_2912,N_2185,N_2044);
nor U2913 (N_2913,N_2455,N_2204);
xnor U2914 (N_2914,N_2290,N_2423);
xor U2915 (N_2915,N_2453,N_2498);
nor U2916 (N_2916,N_2044,N_2107);
and U2917 (N_2917,N_2446,N_2432);
nor U2918 (N_2918,N_2062,N_2014);
or U2919 (N_2919,N_2468,N_2094);
or U2920 (N_2920,N_2487,N_2080);
nor U2921 (N_2921,N_2183,N_2198);
and U2922 (N_2922,N_2200,N_2457);
and U2923 (N_2923,N_2313,N_2284);
xnor U2924 (N_2924,N_2147,N_2074);
nand U2925 (N_2925,N_2309,N_2493);
nand U2926 (N_2926,N_2441,N_2025);
nand U2927 (N_2927,N_2293,N_2083);
and U2928 (N_2928,N_2112,N_2255);
nand U2929 (N_2929,N_2496,N_2385);
and U2930 (N_2930,N_2000,N_2318);
xnor U2931 (N_2931,N_2135,N_2476);
nand U2932 (N_2932,N_2051,N_2069);
and U2933 (N_2933,N_2215,N_2271);
nand U2934 (N_2934,N_2120,N_2103);
xor U2935 (N_2935,N_2360,N_2261);
nor U2936 (N_2936,N_2240,N_2492);
nand U2937 (N_2937,N_2261,N_2102);
and U2938 (N_2938,N_2285,N_2299);
or U2939 (N_2939,N_2257,N_2169);
xor U2940 (N_2940,N_2422,N_2134);
nand U2941 (N_2941,N_2224,N_2246);
nand U2942 (N_2942,N_2231,N_2276);
and U2943 (N_2943,N_2357,N_2247);
and U2944 (N_2944,N_2406,N_2419);
and U2945 (N_2945,N_2082,N_2098);
nor U2946 (N_2946,N_2025,N_2026);
nor U2947 (N_2947,N_2323,N_2340);
and U2948 (N_2948,N_2256,N_2135);
nand U2949 (N_2949,N_2198,N_2485);
or U2950 (N_2950,N_2311,N_2428);
nand U2951 (N_2951,N_2294,N_2274);
xor U2952 (N_2952,N_2277,N_2376);
and U2953 (N_2953,N_2467,N_2413);
nor U2954 (N_2954,N_2324,N_2349);
and U2955 (N_2955,N_2398,N_2235);
xor U2956 (N_2956,N_2131,N_2321);
nor U2957 (N_2957,N_2177,N_2363);
xor U2958 (N_2958,N_2017,N_2144);
nor U2959 (N_2959,N_2000,N_2132);
nor U2960 (N_2960,N_2022,N_2404);
nor U2961 (N_2961,N_2206,N_2311);
and U2962 (N_2962,N_2450,N_2475);
nor U2963 (N_2963,N_2173,N_2236);
xor U2964 (N_2964,N_2446,N_2490);
nand U2965 (N_2965,N_2484,N_2174);
nor U2966 (N_2966,N_2474,N_2001);
and U2967 (N_2967,N_2356,N_2069);
nand U2968 (N_2968,N_2158,N_2438);
nand U2969 (N_2969,N_2393,N_2448);
nand U2970 (N_2970,N_2288,N_2403);
or U2971 (N_2971,N_2494,N_2270);
nor U2972 (N_2972,N_2194,N_2031);
nand U2973 (N_2973,N_2063,N_2168);
nand U2974 (N_2974,N_2254,N_2028);
xor U2975 (N_2975,N_2347,N_2452);
nor U2976 (N_2976,N_2117,N_2059);
and U2977 (N_2977,N_2156,N_2091);
or U2978 (N_2978,N_2181,N_2039);
nand U2979 (N_2979,N_2480,N_2132);
and U2980 (N_2980,N_2446,N_2011);
and U2981 (N_2981,N_2427,N_2160);
and U2982 (N_2982,N_2127,N_2470);
and U2983 (N_2983,N_2164,N_2018);
nor U2984 (N_2984,N_2203,N_2373);
nor U2985 (N_2985,N_2033,N_2053);
nand U2986 (N_2986,N_2152,N_2207);
or U2987 (N_2987,N_2411,N_2095);
nand U2988 (N_2988,N_2356,N_2060);
xnor U2989 (N_2989,N_2211,N_2237);
xor U2990 (N_2990,N_2325,N_2215);
and U2991 (N_2991,N_2265,N_2298);
nor U2992 (N_2992,N_2397,N_2245);
nor U2993 (N_2993,N_2070,N_2415);
nand U2994 (N_2994,N_2183,N_2458);
nand U2995 (N_2995,N_2276,N_2272);
nand U2996 (N_2996,N_2027,N_2259);
nor U2997 (N_2997,N_2424,N_2204);
nand U2998 (N_2998,N_2417,N_2200);
nand U2999 (N_2999,N_2043,N_2208);
or U3000 (N_3000,N_2713,N_2641);
and U3001 (N_3001,N_2507,N_2828);
xor U3002 (N_3002,N_2801,N_2673);
nor U3003 (N_3003,N_2881,N_2595);
and U3004 (N_3004,N_2958,N_2675);
nor U3005 (N_3005,N_2726,N_2626);
nor U3006 (N_3006,N_2657,N_2703);
nand U3007 (N_3007,N_2830,N_2516);
nor U3008 (N_3008,N_2520,N_2632);
xnor U3009 (N_3009,N_2667,N_2878);
xnor U3010 (N_3010,N_2658,N_2571);
nand U3011 (N_3011,N_2739,N_2977);
or U3012 (N_3012,N_2802,N_2775);
or U3013 (N_3013,N_2690,N_2748);
xnor U3014 (N_3014,N_2751,N_2765);
nor U3015 (N_3015,N_2888,N_2646);
xor U3016 (N_3016,N_2897,N_2973);
nand U3017 (N_3017,N_2866,N_2609);
nor U3018 (N_3018,N_2962,N_2928);
or U3019 (N_3019,N_2665,N_2678);
nor U3020 (N_3020,N_2944,N_2939);
or U3021 (N_3021,N_2959,N_2603);
or U3022 (N_3022,N_2808,N_2887);
nor U3023 (N_3023,N_2594,N_2687);
or U3024 (N_3024,N_2870,N_2600);
nand U3025 (N_3025,N_2532,N_2738);
nand U3026 (N_3026,N_2554,N_2776);
nor U3027 (N_3027,N_2869,N_2994);
xor U3028 (N_3028,N_2503,N_2653);
or U3029 (N_3029,N_2895,N_2607);
nor U3030 (N_3030,N_2548,N_2976);
nor U3031 (N_3031,N_2831,N_2664);
xnor U3032 (N_3032,N_2833,N_2654);
nor U3033 (N_3033,N_2922,N_2649);
nand U3034 (N_3034,N_2982,N_2832);
and U3035 (N_3035,N_2631,N_2968);
xnor U3036 (N_3036,N_2911,N_2645);
nand U3037 (N_3037,N_2935,N_2834);
and U3038 (N_3038,N_2555,N_2744);
or U3039 (N_3039,N_2597,N_2666);
or U3040 (N_3040,N_2588,N_2708);
nand U3041 (N_3041,N_2860,N_2582);
nand U3042 (N_3042,N_2947,N_2937);
and U3043 (N_3043,N_2795,N_2576);
xor U3044 (N_3044,N_2586,N_2515);
nand U3045 (N_3045,N_2877,N_2952);
nor U3046 (N_3046,N_2818,N_2696);
and U3047 (N_3047,N_2538,N_2731);
nor U3048 (N_3048,N_2622,N_2508);
nand U3049 (N_3049,N_2916,N_2855);
and U3050 (N_3050,N_2505,N_2661);
nor U3051 (N_3051,N_2745,N_2787);
xor U3052 (N_3052,N_2593,N_2559);
or U3053 (N_3053,N_2697,N_2788);
nor U3054 (N_3054,N_2543,N_2931);
nand U3055 (N_3055,N_2913,N_2615);
xor U3056 (N_3056,N_2614,N_2761);
xnor U3057 (N_3057,N_2647,N_2894);
nand U3058 (N_3058,N_2898,N_2572);
nand U3059 (N_3059,N_2602,N_2964);
and U3060 (N_3060,N_2517,N_2813);
and U3061 (N_3061,N_2610,N_2840);
and U3062 (N_3062,N_2906,N_2784);
nor U3063 (N_3063,N_2825,N_2810);
nor U3064 (N_3064,N_2735,N_2552);
nor U3065 (N_3065,N_2768,N_2770);
xor U3066 (N_3066,N_2752,N_2565);
or U3067 (N_3067,N_2868,N_2859);
or U3068 (N_3068,N_2587,N_2606);
nor U3069 (N_3069,N_2778,N_2749);
nand U3070 (N_3070,N_2852,N_2652);
xnor U3071 (N_3071,N_2642,N_2670);
xor U3072 (N_3072,N_2978,N_2758);
or U3073 (N_3073,N_2635,N_2953);
or U3074 (N_3074,N_2680,N_2707);
or U3075 (N_3075,N_2643,N_2996);
nand U3076 (N_3076,N_2955,N_2500);
xnor U3077 (N_3077,N_2817,N_2943);
xnor U3078 (N_3078,N_2717,N_2779);
and U3079 (N_3079,N_2890,N_2527);
nor U3080 (N_3080,N_2736,N_2743);
xor U3081 (N_3081,N_2692,N_2562);
nor U3082 (N_3082,N_2721,N_2545);
nor U3083 (N_3083,N_2710,N_2793);
nor U3084 (N_3084,N_2669,N_2984);
xnor U3085 (N_3085,N_2725,N_2811);
nor U3086 (N_3086,N_2522,N_2742);
or U3087 (N_3087,N_2704,N_2974);
and U3088 (N_3088,N_2618,N_2836);
or U3089 (N_3089,N_2957,N_2938);
xnor U3090 (N_3090,N_2750,N_2566);
nand U3091 (N_3091,N_2530,N_2858);
xor U3092 (N_3092,N_2722,N_2961);
or U3093 (N_3093,N_2907,N_2542);
or U3094 (N_3094,N_2567,N_2676);
nor U3095 (N_3095,N_2910,N_2519);
or U3096 (N_3096,N_2843,N_2620);
nor U3097 (N_3097,N_2526,N_2728);
and U3098 (N_3098,N_2668,N_2790);
nor U3099 (N_3099,N_2573,N_2874);
xnor U3100 (N_3100,N_2989,N_2783);
nand U3101 (N_3101,N_2891,N_2908);
nand U3102 (N_3102,N_2863,N_2899);
xor U3103 (N_3103,N_2629,N_2556);
and U3104 (N_3104,N_2915,N_2763);
or U3105 (N_3105,N_2700,N_2585);
nand U3106 (N_3106,N_2772,N_2826);
nor U3107 (N_3107,N_2659,N_2900);
or U3108 (N_3108,N_2862,N_2988);
xor U3109 (N_3109,N_2674,N_2809);
xnor U3110 (N_3110,N_2794,N_2592);
and U3111 (N_3111,N_2934,N_2577);
or U3112 (N_3112,N_2814,N_2997);
nor U3113 (N_3113,N_2510,N_2789);
nor U3114 (N_3114,N_2621,N_2812);
and U3115 (N_3115,N_2716,N_2861);
nor U3116 (N_3116,N_2589,N_2917);
and U3117 (N_3117,N_2979,N_2693);
nand U3118 (N_3118,N_2655,N_2564);
and U3119 (N_3119,N_2901,N_2511);
and U3120 (N_3120,N_2966,N_2998);
nor U3121 (N_3121,N_2702,N_2912);
xnor U3122 (N_3122,N_2651,N_2625);
nor U3123 (N_3123,N_2771,N_2921);
nor U3124 (N_3124,N_2804,N_2925);
or U3125 (N_3125,N_2537,N_2681);
nor U3126 (N_3126,N_2981,N_2648);
nor U3127 (N_3127,N_2807,N_2549);
nor U3128 (N_3128,N_2838,N_2924);
nand U3129 (N_3129,N_2756,N_2963);
or U3130 (N_3130,N_2927,N_2942);
nand U3131 (N_3131,N_2506,N_2767);
and U3132 (N_3132,N_2521,N_2960);
and U3133 (N_3133,N_2580,N_2584);
nor U3134 (N_3134,N_2839,N_2701);
nand U3135 (N_3135,N_2617,N_2920);
or U3136 (N_3136,N_2724,N_2769);
or U3137 (N_3137,N_2513,N_2883);
and U3138 (N_3138,N_2746,N_2672);
or U3139 (N_3139,N_2841,N_2579);
xor U3140 (N_3140,N_2885,N_2914);
and U3141 (N_3141,N_2623,N_2558);
nand U3142 (N_3142,N_2705,N_2876);
and U3143 (N_3143,N_2821,N_2853);
xnor U3144 (N_3144,N_2764,N_2777);
and U3145 (N_3145,N_2820,N_2611);
nor U3146 (N_3146,N_2598,N_2972);
xor U3147 (N_3147,N_2636,N_2849);
or U3148 (N_3148,N_2850,N_2509);
nand U3149 (N_3149,N_2941,N_2754);
xnor U3150 (N_3150,N_2946,N_2682);
nor U3151 (N_3151,N_2786,N_2936);
nor U3152 (N_3152,N_2695,N_2759);
nor U3153 (N_3153,N_2683,N_2686);
or U3154 (N_3154,N_2546,N_2842);
or U3155 (N_3155,N_2684,N_2685);
and U3156 (N_3156,N_2835,N_2797);
and U3157 (N_3157,N_2837,N_2715);
nand U3158 (N_3158,N_2956,N_2590);
nor U3159 (N_3159,N_2766,N_2711);
or U3160 (N_3160,N_2905,N_2528);
or U3161 (N_3161,N_2949,N_2827);
nor U3162 (N_3162,N_2604,N_2923);
nand U3163 (N_3163,N_2741,N_2985);
xor U3164 (N_3164,N_2718,N_2514);
or U3165 (N_3165,N_2940,N_2755);
nor U3166 (N_3166,N_2930,N_2965);
nand U3167 (N_3167,N_2918,N_2539);
or U3168 (N_3168,N_2829,N_2563);
and U3169 (N_3169,N_2689,N_2677);
nor U3170 (N_3170,N_2541,N_2523);
and U3171 (N_3171,N_2706,N_2720);
nor U3172 (N_3172,N_2879,N_2656);
nand U3173 (N_3173,N_2889,N_2524);
and U3174 (N_3174,N_2823,N_2760);
or U3175 (N_3175,N_2815,N_2660);
nor U3176 (N_3176,N_2525,N_2926);
xor U3177 (N_3177,N_2583,N_2799);
or U3178 (N_3178,N_2990,N_2805);
or U3179 (N_3179,N_2662,N_2730);
or U3180 (N_3180,N_2747,N_2872);
and U3181 (N_3181,N_2613,N_2803);
nand U3182 (N_3182,N_2574,N_2856);
nand U3183 (N_3183,N_2847,N_2599);
nand U3184 (N_3184,N_2688,N_2634);
nand U3185 (N_3185,N_2624,N_2719);
and U3186 (N_3186,N_2550,N_2848);
or U3187 (N_3187,N_2800,N_2581);
nor U3188 (N_3188,N_2774,N_2630);
and U3189 (N_3189,N_2529,N_2954);
xor U3190 (N_3190,N_2986,N_2864);
xor U3191 (N_3191,N_2798,N_2865);
or U3192 (N_3192,N_2640,N_2857);
nor U3193 (N_3193,N_2873,N_2904);
nor U3194 (N_3194,N_2551,N_2951);
nand U3195 (N_3195,N_2845,N_2557);
xnor U3196 (N_3196,N_2547,N_2533);
and U3197 (N_3197,N_2570,N_2737);
nand U3198 (N_3198,N_2792,N_2502);
or U3199 (N_3199,N_2727,N_2919);
nand U3200 (N_3200,N_2971,N_2663);
and U3201 (N_3201,N_2619,N_2757);
nand U3202 (N_3202,N_2992,N_2773);
xnor U3203 (N_3203,N_2560,N_2782);
nor U3204 (N_3204,N_2644,N_2886);
or U3205 (N_3205,N_2882,N_2867);
xor U3206 (N_3206,N_2540,N_2819);
and U3207 (N_3207,N_2995,N_2780);
nor U3208 (N_3208,N_2753,N_2679);
and U3209 (N_3209,N_2762,N_2723);
nand U3210 (N_3210,N_2531,N_2544);
nand U3211 (N_3211,N_2699,N_2638);
xnor U3212 (N_3212,N_2608,N_2933);
or U3213 (N_3213,N_2884,N_2796);
and U3214 (N_3214,N_2824,N_2822);
and U3215 (N_3215,N_2712,N_2875);
or U3216 (N_3216,N_2909,N_2851);
and U3217 (N_3217,N_2639,N_2880);
nor U3218 (N_3218,N_2578,N_2892);
or U3219 (N_3219,N_2732,N_2650);
and U3220 (N_3220,N_2627,N_2781);
or U3221 (N_3221,N_2991,N_2893);
nor U3222 (N_3222,N_2993,N_2628);
or U3223 (N_3223,N_2637,N_2987);
xnor U3224 (N_3224,N_2999,N_2512);
and U3225 (N_3225,N_2535,N_2569);
nor U3226 (N_3226,N_2871,N_2501);
nand U3227 (N_3227,N_2948,N_2575);
nor U3228 (N_3228,N_2734,N_2816);
xor U3229 (N_3229,N_2945,N_2691);
and U3230 (N_3230,N_2967,N_2729);
nor U3231 (N_3231,N_2929,N_2561);
nor U3232 (N_3232,N_2785,N_2932);
xor U3233 (N_3233,N_2504,N_2846);
and U3234 (N_3234,N_2553,N_2903);
nor U3235 (N_3235,N_2975,N_2591);
and U3236 (N_3236,N_2950,N_2709);
xor U3237 (N_3237,N_2854,N_2740);
xor U3238 (N_3238,N_2536,N_2534);
and U3239 (N_3239,N_2733,N_2844);
nand U3240 (N_3240,N_2671,N_2791);
or U3241 (N_3241,N_2605,N_2896);
nor U3242 (N_3242,N_2806,N_2969);
nand U3243 (N_3243,N_2601,N_2596);
and U3244 (N_3244,N_2980,N_2633);
and U3245 (N_3245,N_2970,N_2616);
nand U3246 (N_3246,N_2983,N_2568);
or U3247 (N_3247,N_2902,N_2694);
xnor U3248 (N_3248,N_2714,N_2698);
and U3249 (N_3249,N_2612,N_2518);
and U3250 (N_3250,N_2855,N_2630);
nor U3251 (N_3251,N_2636,N_2798);
nand U3252 (N_3252,N_2964,N_2917);
or U3253 (N_3253,N_2538,N_2858);
xnor U3254 (N_3254,N_2748,N_2815);
or U3255 (N_3255,N_2774,N_2970);
xnor U3256 (N_3256,N_2526,N_2977);
nand U3257 (N_3257,N_2606,N_2729);
or U3258 (N_3258,N_2674,N_2966);
and U3259 (N_3259,N_2809,N_2938);
or U3260 (N_3260,N_2698,N_2861);
nor U3261 (N_3261,N_2781,N_2552);
nand U3262 (N_3262,N_2789,N_2587);
nor U3263 (N_3263,N_2524,N_2636);
nor U3264 (N_3264,N_2512,N_2678);
or U3265 (N_3265,N_2919,N_2715);
xnor U3266 (N_3266,N_2783,N_2834);
nand U3267 (N_3267,N_2679,N_2923);
or U3268 (N_3268,N_2977,N_2519);
and U3269 (N_3269,N_2747,N_2536);
and U3270 (N_3270,N_2833,N_2622);
or U3271 (N_3271,N_2824,N_2937);
nor U3272 (N_3272,N_2667,N_2809);
or U3273 (N_3273,N_2513,N_2934);
nor U3274 (N_3274,N_2858,N_2503);
or U3275 (N_3275,N_2617,N_2668);
and U3276 (N_3276,N_2667,N_2916);
xor U3277 (N_3277,N_2610,N_2974);
or U3278 (N_3278,N_2871,N_2758);
nand U3279 (N_3279,N_2646,N_2704);
xnor U3280 (N_3280,N_2831,N_2573);
and U3281 (N_3281,N_2755,N_2764);
nand U3282 (N_3282,N_2794,N_2957);
xor U3283 (N_3283,N_2541,N_2731);
or U3284 (N_3284,N_2926,N_2642);
nand U3285 (N_3285,N_2628,N_2626);
nand U3286 (N_3286,N_2887,N_2673);
nor U3287 (N_3287,N_2542,N_2951);
xor U3288 (N_3288,N_2575,N_2660);
or U3289 (N_3289,N_2710,N_2559);
nand U3290 (N_3290,N_2502,N_2645);
or U3291 (N_3291,N_2840,N_2508);
or U3292 (N_3292,N_2959,N_2682);
nor U3293 (N_3293,N_2861,N_2741);
nor U3294 (N_3294,N_2660,N_2933);
xor U3295 (N_3295,N_2983,N_2888);
nor U3296 (N_3296,N_2570,N_2664);
or U3297 (N_3297,N_2879,N_2692);
or U3298 (N_3298,N_2626,N_2795);
and U3299 (N_3299,N_2630,N_2767);
nand U3300 (N_3300,N_2635,N_2592);
xnor U3301 (N_3301,N_2847,N_2608);
nand U3302 (N_3302,N_2540,N_2877);
xor U3303 (N_3303,N_2628,N_2924);
or U3304 (N_3304,N_2785,N_2832);
and U3305 (N_3305,N_2502,N_2757);
nor U3306 (N_3306,N_2700,N_2509);
xor U3307 (N_3307,N_2657,N_2533);
nand U3308 (N_3308,N_2957,N_2924);
nand U3309 (N_3309,N_2737,N_2726);
xnor U3310 (N_3310,N_2961,N_2787);
nor U3311 (N_3311,N_2509,N_2735);
nor U3312 (N_3312,N_2843,N_2876);
nand U3313 (N_3313,N_2549,N_2600);
nor U3314 (N_3314,N_2696,N_2546);
nor U3315 (N_3315,N_2630,N_2652);
and U3316 (N_3316,N_2605,N_2812);
or U3317 (N_3317,N_2933,N_2611);
nor U3318 (N_3318,N_2795,N_2751);
or U3319 (N_3319,N_2768,N_2821);
nor U3320 (N_3320,N_2661,N_2557);
xnor U3321 (N_3321,N_2998,N_2879);
nor U3322 (N_3322,N_2526,N_2966);
nor U3323 (N_3323,N_2549,N_2585);
or U3324 (N_3324,N_2989,N_2509);
nor U3325 (N_3325,N_2807,N_2595);
xor U3326 (N_3326,N_2911,N_2656);
and U3327 (N_3327,N_2857,N_2801);
nor U3328 (N_3328,N_2556,N_2681);
and U3329 (N_3329,N_2548,N_2509);
and U3330 (N_3330,N_2744,N_2551);
or U3331 (N_3331,N_2961,N_2898);
nor U3332 (N_3332,N_2917,N_2984);
xor U3333 (N_3333,N_2771,N_2694);
and U3334 (N_3334,N_2792,N_2809);
or U3335 (N_3335,N_2841,N_2557);
or U3336 (N_3336,N_2986,N_2729);
and U3337 (N_3337,N_2831,N_2593);
and U3338 (N_3338,N_2938,N_2647);
or U3339 (N_3339,N_2821,N_2532);
and U3340 (N_3340,N_2719,N_2603);
xor U3341 (N_3341,N_2658,N_2999);
or U3342 (N_3342,N_2936,N_2592);
or U3343 (N_3343,N_2998,N_2546);
and U3344 (N_3344,N_2523,N_2823);
nand U3345 (N_3345,N_2772,N_2916);
and U3346 (N_3346,N_2958,N_2788);
or U3347 (N_3347,N_2924,N_2925);
nand U3348 (N_3348,N_2639,N_2773);
nor U3349 (N_3349,N_2605,N_2984);
nor U3350 (N_3350,N_2942,N_2728);
nor U3351 (N_3351,N_2513,N_2926);
nand U3352 (N_3352,N_2535,N_2783);
or U3353 (N_3353,N_2835,N_2897);
nand U3354 (N_3354,N_2760,N_2681);
and U3355 (N_3355,N_2973,N_2591);
or U3356 (N_3356,N_2545,N_2734);
nand U3357 (N_3357,N_2621,N_2959);
xnor U3358 (N_3358,N_2779,N_2723);
nor U3359 (N_3359,N_2843,N_2604);
or U3360 (N_3360,N_2592,N_2504);
and U3361 (N_3361,N_2896,N_2812);
or U3362 (N_3362,N_2837,N_2981);
or U3363 (N_3363,N_2787,N_2907);
nand U3364 (N_3364,N_2926,N_2734);
nand U3365 (N_3365,N_2559,N_2619);
xor U3366 (N_3366,N_2768,N_2869);
xnor U3367 (N_3367,N_2946,N_2520);
and U3368 (N_3368,N_2554,N_2627);
and U3369 (N_3369,N_2947,N_2938);
xor U3370 (N_3370,N_2527,N_2724);
or U3371 (N_3371,N_2808,N_2668);
or U3372 (N_3372,N_2869,N_2598);
and U3373 (N_3373,N_2543,N_2785);
or U3374 (N_3374,N_2695,N_2501);
nand U3375 (N_3375,N_2626,N_2931);
xnor U3376 (N_3376,N_2981,N_2714);
and U3377 (N_3377,N_2535,N_2666);
and U3378 (N_3378,N_2553,N_2584);
and U3379 (N_3379,N_2516,N_2835);
or U3380 (N_3380,N_2630,N_2584);
nor U3381 (N_3381,N_2778,N_2880);
xor U3382 (N_3382,N_2665,N_2640);
or U3383 (N_3383,N_2732,N_2964);
and U3384 (N_3384,N_2625,N_2844);
and U3385 (N_3385,N_2958,N_2552);
or U3386 (N_3386,N_2527,N_2561);
nor U3387 (N_3387,N_2594,N_2966);
nor U3388 (N_3388,N_2831,N_2742);
and U3389 (N_3389,N_2875,N_2828);
nor U3390 (N_3390,N_2741,N_2651);
xor U3391 (N_3391,N_2996,N_2648);
xor U3392 (N_3392,N_2758,N_2646);
nand U3393 (N_3393,N_2639,N_2573);
xor U3394 (N_3394,N_2711,N_2923);
nor U3395 (N_3395,N_2992,N_2841);
nor U3396 (N_3396,N_2910,N_2980);
xor U3397 (N_3397,N_2836,N_2682);
nor U3398 (N_3398,N_2784,N_2501);
nor U3399 (N_3399,N_2848,N_2973);
or U3400 (N_3400,N_2809,N_2525);
or U3401 (N_3401,N_2619,N_2693);
nor U3402 (N_3402,N_2820,N_2869);
or U3403 (N_3403,N_2966,N_2893);
nor U3404 (N_3404,N_2923,N_2950);
nor U3405 (N_3405,N_2616,N_2639);
nor U3406 (N_3406,N_2866,N_2622);
xnor U3407 (N_3407,N_2962,N_2711);
nor U3408 (N_3408,N_2844,N_2843);
and U3409 (N_3409,N_2579,N_2978);
nand U3410 (N_3410,N_2969,N_2824);
or U3411 (N_3411,N_2618,N_2596);
nor U3412 (N_3412,N_2611,N_2718);
nand U3413 (N_3413,N_2810,N_2799);
or U3414 (N_3414,N_2976,N_2990);
or U3415 (N_3415,N_2622,N_2694);
nor U3416 (N_3416,N_2827,N_2921);
or U3417 (N_3417,N_2999,N_2812);
or U3418 (N_3418,N_2561,N_2574);
nor U3419 (N_3419,N_2743,N_2767);
xor U3420 (N_3420,N_2634,N_2783);
nand U3421 (N_3421,N_2711,N_2774);
xor U3422 (N_3422,N_2692,N_2805);
nand U3423 (N_3423,N_2896,N_2952);
nand U3424 (N_3424,N_2577,N_2769);
or U3425 (N_3425,N_2688,N_2908);
nor U3426 (N_3426,N_2550,N_2799);
xor U3427 (N_3427,N_2902,N_2926);
nor U3428 (N_3428,N_2746,N_2748);
nor U3429 (N_3429,N_2604,N_2893);
nand U3430 (N_3430,N_2807,N_2774);
or U3431 (N_3431,N_2800,N_2552);
nor U3432 (N_3432,N_2911,N_2688);
xnor U3433 (N_3433,N_2621,N_2706);
nor U3434 (N_3434,N_2833,N_2930);
xor U3435 (N_3435,N_2501,N_2697);
nor U3436 (N_3436,N_2983,N_2828);
nor U3437 (N_3437,N_2599,N_2724);
or U3438 (N_3438,N_2820,N_2874);
nor U3439 (N_3439,N_2656,N_2598);
and U3440 (N_3440,N_2675,N_2756);
and U3441 (N_3441,N_2977,N_2797);
and U3442 (N_3442,N_2859,N_2945);
xor U3443 (N_3443,N_2803,N_2835);
or U3444 (N_3444,N_2834,N_2866);
and U3445 (N_3445,N_2827,N_2600);
and U3446 (N_3446,N_2695,N_2633);
nor U3447 (N_3447,N_2588,N_2785);
and U3448 (N_3448,N_2649,N_2969);
or U3449 (N_3449,N_2856,N_2739);
nor U3450 (N_3450,N_2589,N_2660);
and U3451 (N_3451,N_2805,N_2959);
xnor U3452 (N_3452,N_2797,N_2923);
nand U3453 (N_3453,N_2692,N_2720);
nor U3454 (N_3454,N_2782,N_2963);
and U3455 (N_3455,N_2762,N_2691);
or U3456 (N_3456,N_2539,N_2695);
nand U3457 (N_3457,N_2968,N_2863);
nor U3458 (N_3458,N_2973,N_2541);
xnor U3459 (N_3459,N_2692,N_2864);
nand U3460 (N_3460,N_2937,N_2674);
nor U3461 (N_3461,N_2932,N_2896);
or U3462 (N_3462,N_2570,N_2938);
and U3463 (N_3463,N_2792,N_2785);
nand U3464 (N_3464,N_2889,N_2660);
nand U3465 (N_3465,N_2569,N_2614);
and U3466 (N_3466,N_2805,N_2640);
and U3467 (N_3467,N_2984,N_2665);
xor U3468 (N_3468,N_2788,N_2922);
xor U3469 (N_3469,N_2835,N_2892);
nor U3470 (N_3470,N_2921,N_2933);
or U3471 (N_3471,N_2689,N_2930);
nand U3472 (N_3472,N_2671,N_2584);
and U3473 (N_3473,N_2938,N_2813);
and U3474 (N_3474,N_2756,N_2591);
xor U3475 (N_3475,N_2680,N_2760);
or U3476 (N_3476,N_2627,N_2574);
xnor U3477 (N_3477,N_2522,N_2531);
nor U3478 (N_3478,N_2811,N_2642);
nand U3479 (N_3479,N_2721,N_2535);
and U3480 (N_3480,N_2977,N_2585);
xnor U3481 (N_3481,N_2700,N_2672);
or U3482 (N_3482,N_2646,N_2572);
or U3483 (N_3483,N_2876,N_2666);
and U3484 (N_3484,N_2800,N_2503);
and U3485 (N_3485,N_2959,N_2881);
or U3486 (N_3486,N_2796,N_2588);
xor U3487 (N_3487,N_2901,N_2548);
or U3488 (N_3488,N_2984,N_2835);
and U3489 (N_3489,N_2529,N_2571);
nand U3490 (N_3490,N_2505,N_2566);
nor U3491 (N_3491,N_2595,N_2682);
nand U3492 (N_3492,N_2967,N_2904);
and U3493 (N_3493,N_2656,N_2571);
or U3494 (N_3494,N_2742,N_2526);
nand U3495 (N_3495,N_2940,N_2555);
or U3496 (N_3496,N_2776,N_2725);
and U3497 (N_3497,N_2718,N_2767);
or U3498 (N_3498,N_2945,N_2557);
xor U3499 (N_3499,N_2919,N_2883);
xnor U3500 (N_3500,N_3130,N_3304);
xor U3501 (N_3501,N_3102,N_3122);
and U3502 (N_3502,N_3178,N_3242);
nor U3503 (N_3503,N_3456,N_3053);
nor U3504 (N_3504,N_3087,N_3054);
nand U3505 (N_3505,N_3416,N_3103);
and U3506 (N_3506,N_3414,N_3355);
nor U3507 (N_3507,N_3124,N_3104);
or U3508 (N_3508,N_3361,N_3489);
or U3509 (N_3509,N_3186,N_3234);
nor U3510 (N_3510,N_3192,N_3310);
nand U3511 (N_3511,N_3026,N_3040);
or U3512 (N_3512,N_3145,N_3386);
and U3513 (N_3513,N_3332,N_3455);
xnor U3514 (N_3514,N_3008,N_3101);
nand U3515 (N_3515,N_3035,N_3482);
or U3516 (N_3516,N_3410,N_3084);
xnor U3517 (N_3517,N_3289,N_3014);
nand U3518 (N_3518,N_3062,N_3225);
nor U3519 (N_3519,N_3315,N_3346);
nor U3520 (N_3520,N_3058,N_3016);
xnor U3521 (N_3521,N_3193,N_3251);
nand U3522 (N_3522,N_3350,N_3415);
xnor U3523 (N_3523,N_3172,N_3345);
and U3524 (N_3524,N_3190,N_3140);
nor U3525 (N_3525,N_3268,N_3454);
nand U3526 (N_3526,N_3316,N_3002);
and U3527 (N_3527,N_3433,N_3137);
nor U3528 (N_3528,N_3215,N_3487);
nor U3529 (N_3529,N_3167,N_3152);
and U3530 (N_3530,N_3179,N_3387);
nand U3531 (N_3531,N_3371,N_3453);
xor U3532 (N_3532,N_3119,N_3282);
nor U3533 (N_3533,N_3088,N_3470);
nand U3534 (N_3534,N_3363,N_3318);
nor U3535 (N_3535,N_3370,N_3066);
or U3536 (N_3536,N_3442,N_3078);
nand U3537 (N_3537,N_3471,N_3430);
or U3538 (N_3538,N_3202,N_3207);
xor U3539 (N_3539,N_3177,N_3074);
nor U3540 (N_3540,N_3422,N_3080);
nor U3541 (N_3541,N_3176,N_3025);
xor U3542 (N_3542,N_3254,N_3075);
and U3543 (N_3543,N_3280,N_3153);
xor U3544 (N_3544,N_3438,N_3314);
xor U3545 (N_3545,N_3391,N_3162);
nand U3546 (N_3546,N_3312,N_3020);
nor U3547 (N_3547,N_3379,N_3108);
and U3548 (N_3548,N_3443,N_3231);
xor U3549 (N_3549,N_3417,N_3060);
nand U3550 (N_3550,N_3271,N_3405);
or U3551 (N_3551,N_3352,N_3419);
or U3552 (N_3552,N_3056,N_3079);
or U3553 (N_3553,N_3073,N_3490);
or U3554 (N_3554,N_3129,N_3019);
nor U3555 (N_3555,N_3121,N_3156);
xnor U3556 (N_3556,N_3126,N_3406);
nand U3557 (N_3557,N_3384,N_3321);
xor U3558 (N_3558,N_3399,N_3045);
xor U3559 (N_3559,N_3389,N_3021);
or U3560 (N_3560,N_3360,N_3206);
nor U3561 (N_3561,N_3498,N_3340);
nand U3562 (N_3562,N_3181,N_3032);
or U3563 (N_3563,N_3277,N_3009);
nor U3564 (N_3564,N_3013,N_3089);
xor U3565 (N_3565,N_3267,N_3434);
and U3566 (N_3566,N_3022,N_3180);
or U3567 (N_3567,N_3086,N_3402);
nor U3568 (N_3568,N_3157,N_3241);
nand U3569 (N_3569,N_3467,N_3291);
nand U3570 (N_3570,N_3418,N_3359);
xor U3571 (N_3571,N_3049,N_3283);
nand U3572 (N_3572,N_3237,N_3376);
nand U3573 (N_3573,N_3123,N_3472);
or U3574 (N_3574,N_3023,N_3462);
nor U3575 (N_3575,N_3059,N_3091);
or U3576 (N_3576,N_3041,N_3496);
or U3577 (N_3577,N_3311,N_3128);
nor U3578 (N_3578,N_3497,N_3463);
and U3579 (N_3579,N_3229,N_3136);
xnor U3580 (N_3580,N_3293,N_3432);
nand U3581 (N_3581,N_3252,N_3249);
nand U3582 (N_3582,N_3302,N_3184);
xnor U3583 (N_3583,N_3048,N_3199);
xor U3584 (N_3584,N_3243,N_3174);
nand U3585 (N_3585,N_3272,N_3003);
and U3586 (N_3586,N_3147,N_3439);
nand U3587 (N_3587,N_3480,N_3459);
nand U3588 (N_3588,N_3495,N_3475);
nor U3589 (N_3589,N_3211,N_3191);
or U3590 (N_3590,N_3110,N_3135);
nand U3591 (N_3591,N_3149,N_3465);
and U3592 (N_3592,N_3208,N_3077);
xnor U3593 (N_3593,N_3245,N_3292);
or U3594 (N_3594,N_3468,N_3423);
nand U3595 (N_3595,N_3161,N_3481);
or U3596 (N_3596,N_3165,N_3256);
and U3597 (N_3597,N_3188,N_3004);
or U3598 (N_3598,N_3330,N_3483);
xor U3599 (N_3599,N_3300,N_3365);
or U3600 (N_3600,N_3261,N_3341);
xor U3601 (N_3601,N_3431,N_3220);
nand U3602 (N_3602,N_3440,N_3201);
nor U3603 (N_3603,N_3445,N_3285);
nor U3604 (N_3604,N_3063,N_3114);
nand U3605 (N_3605,N_3115,N_3297);
nand U3606 (N_3606,N_3353,N_3466);
or U3607 (N_3607,N_3164,N_3037);
or U3608 (N_3608,N_3150,N_3185);
nor U3609 (N_3609,N_3117,N_3239);
nor U3610 (N_3610,N_3067,N_3082);
or U3611 (N_3611,N_3120,N_3322);
xor U3612 (N_3612,N_3112,N_3055);
or U3613 (N_3613,N_3027,N_3069);
nand U3614 (N_3614,N_3036,N_3044);
nor U3615 (N_3615,N_3362,N_3017);
nor U3616 (N_3616,N_3326,N_3295);
and U3617 (N_3617,N_3388,N_3336);
xor U3618 (N_3618,N_3170,N_3342);
or U3619 (N_3619,N_3486,N_3448);
nor U3620 (N_3620,N_3046,N_3427);
or U3621 (N_3621,N_3477,N_3307);
nand U3622 (N_3622,N_3327,N_3141);
nand U3623 (N_3623,N_3118,N_3401);
or U3624 (N_3624,N_3096,N_3323);
nand U3625 (N_3625,N_3047,N_3380);
nor U3626 (N_3626,N_3093,N_3085);
xnor U3627 (N_3627,N_3383,N_3375);
nand U3628 (N_3628,N_3024,N_3007);
or U3629 (N_3629,N_3042,N_3368);
xnor U3630 (N_3630,N_3499,N_3043);
nand U3631 (N_3631,N_3488,N_3226);
xor U3632 (N_3632,N_3457,N_3424);
or U3633 (N_3633,N_3100,N_3484);
and U3634 (N_3634,N_3052,N_3446);
xnor U3635 (N_3635,N_3298,N_3214);
nand U3636 (N_3636,N_3250,N_3319);
nor U3637 (N_3637,N_3038,N_3366);
xnor U3638 (N_3638,N_3491,N_3494);
and U3639 (N_3639,N_3294,N_3284);
nor U3640 (N_3640,N_3068,N_3255);
and U3641 (N_3641,N_3274,N_3286);
and U3642 (N_3642,N_3348,N_3182);
xnor U3643 (N_3643,N_3447,N_3394);
xnor U3644 (N_3644,N_3218,N_3273);
or U3645 (N_3645,N_3473,N_3325);
xnor U3646 (N_3646,N_3479,N_3263);
and U3647 (N_3647,N_3364,N_3260);
xnor U3648 (N_3648,N_3236,N_3476);
nor U3649 (N_3649,N_3143,N_3175);
xnor U3650 (N_3650,N_3264,N_3339);
nand U3651 (N_3651,N_3328,N_3381);
or U3652 (N_3652,N_3219,N_3372);
nor U3653 (N_3653,N_3374,N_3265);
and U3654 (N_3654,N_3144,N_3299);
or U3655 (N_3655,N_3051,N_3148);
or U3656 (N_3656,N_3400,N_3278);
nor U3657 (N_3657,N_3397,N_3194);
nor U3658 (N_3658,N_3006,N_3411);
or U3659 (N_3659,N_3138,N_3099);
and U3660 (N_3660,N_3478,N_3493);
nor U3661 (N_3661,N_3171,N_3428);
or U3662 (N_3662,N_3158,N_3132);
nor U3663 (N_3663,N_3213,N_3195);
nor U3664 (N_3664,N_3398,N_3395);
and U3665 (N_3665,N_3151,N_3449);
nand U3666 (N_3666,N_3262,N_3358);
nand U3667 (N_3667,N_3458,N_3308);
nor U3668 (N_3668,N_3306,N_3098);
nor U3669 (N_3669,N_3238,N_3270);
and U3670 (N_3670,N_3197,N_3113);
nor U3671 (N_3671,N_3131,N_3061);
nand U3672 (N_3672,N_3216,N_3065);
nand U3673 (N_3673,N_3469,N_3246);
nor U3674 (N_3674,N_3109,N_3451);
and U3675 (N_3675,N_3076,N_3441);
nor U3676 (N_3676,N_3240,N_3000);
nand U3677 (N_3677,N_3257,N_3039);
and U3678 (N_3678,N_3413,N_3015);
nor U3679 (N_3679,N_3189,N_3373);
nand U3680 (N_3680,N_3247,N_3222);
and U3681 (N_3681,N_3357,N_3233);
or U3682 (N_3682,N_3309,N_3349);
xnor U3683 (N_3683,N_3166,N_3116);
nand U3684 (N_3684,N_3337,N_3356);
xnor U3685 (N_3685,N_3452,N_3369);
or U3686 (N_3686,N_3403,N_3196);
nand U3687 (N_3687,N_3198,N_3317);
xor U3688 (N_3688,N_3155,N_3212);
and U3689 (N_3689,N_3425,N_3460);
or U3690 (N_3690,N_3146,N_3377);
nor U3691 (N_3691,N_3324,N_3169);
nor U3692 (N_3692,N_3031,N_3094);
xor U3693 (N_3693,N_3407,N_3029);
or U3694 (N_3694,N_3354,N_3097);
xnor U3695 (N_3695,N_3072,N_3335);
or U3696 (N_3696,N_3071,N_3276);
nor U3697 (N_3697,N_3392,N_3107);
or U3698 (N_3698,N_3227,N_3351);
nand U3699 (N_3699,N_3203,N_3296);
xor U3700 (N_3700,N_3092,N_3288);
nor U3701 (N_3701,N_3139,N_3244);
or U3702 (N_3702,N_3183,N_3279);
xnor U3703 (N_3703,N_3010,N_3232);
nand U3704 (N_3704,N_3313,N_3168);
nor U3705 (N_3705,N_3485,N_3050);
or U3706 (N_3706,N_3421,N_3070);
nand U3707 (N_3707,N_3134,N_3492);
or U3708 (N_3708,N_3287,N_3329);
and U3709 (N_3709,N_3106,N_3303);
xor U3710 (N_3710,N_3334,N_3200);
nor U3711 (N_3711,N_3159,N_3253);
nand U3712 (N_3712,N_3223,N_3301);
xnor U3713 (N_3713,N_3436,N_3393);
nor U3714 (N_3714,N_3001,N_3011);
or U3715 (N_3715,N_3111,N_3133);
nand U3716 (N_3716,N_3224,N_3018);
nand U3717 (N_3717,N_3034,N_3281);
or U3718 (N_3718,N_3464,N_3005);
nor U3719 (N_3719,N_3333,N_3331);
nand U3720 (N_3720,N_3305,N_3230);
and U3721 (N_3721,N_3028,N_3344);
xor U3722 (N_3722,N_3266,N_3338);
xor U3723 (N_3723,N_3221,N_3064);
and U3724 (N_3724,N_3474,N_3127);
xnor U3725 (N_3725,N_3426,N_3275);
and U3726 (N_3726,N_3033,N_3409);
or U3727 (N_3727,N_3095,N_3081);
nor U3728 (N_3728,N_3320,N_3429);
and U3729 (N_3729,N_3347,N_3187);
and U3730 (N_3730,N_3396,N_3125);
and U3731 (N_3731,N_3412,N_3378);
nor U3732 (N_3732,N_3205,N_3173);
nand U3733 (N_3733,N_3259,N_3444);
or U3734 (N_3734,N_3209,N_3258);
nor U3735 (N_3735,N_3160,N_3090);
or U3736 (N_3736,N_3404,N_3235);
xor U3737 (N_3737,N_3269,N_3154);
xor U3738 (N_3738,N_3385,N_3408);
and U3739 (N_3739,N_3105,N_3343);
nor U3740 (N_3740,N_3057,N_3435);
nor U3741 (N_3741,N_3290,N_3437);
nand U3742 (N_3742,N_3204,N_3217);
nand U3743 (N_3743,N_3382,N_3450);
and U3744 (N_3744,N_3248,N_3163);
nor U3745 (N_3745,N_3210,N_3367);
or U3746 (N_3746,N_3142,N_3228);
xor U3747 (N_3747,N_3030,N_3390);
or U3748 (N_3748,N_3083,N_3420);
xor U3749 (N_3749,N_3461,N_3012);
nor U3750 (N_3750,N_3354,N_3310);
and U3751 (N_3751,N_3469,N_3021);
nand U3752 (N_3752,N_3000,N_3360);
or U3753 (N_3753,N_3316,N_3084);
nor U3754 (N_3754,N_3109,N_3025);
nand U3755 (N_3755,N_3348,N_3490);
nor U3756 (N_3756,N_3440,N_3224);
or U3757 (N_3757,N_3448,N_3105);
nand U3758 (N_3758,N_3329,N_3378);
xor U3759 (N_3759,N_3334,N_3183);
or U3760 (N_3760,N_3401,N_3333);
nand U3761 (N_3761,N_3150,N_3266);
or U3762 (N_3762,N_3219,N_3187);
nor U3763 (N_3763,N_3364,N_3142);
nand U3764 (N_3764,N_3348,N_3419);
xnor U3765 (N_3765,N_3141,N_3329);
xnor U3766 (N_3766,N_3067,N_3246);
or U3767 (N_3767,N_3056,N_3304);
xnor U3768 (N_3768,N_3494,N_3171);
nand U3769 (N_3769,N_3253,N_3206);
and U3770 (N_3770,N_3244,N_3238);
and U3771 (N_3771,N_3388,N_3375);
nor U3772 (N_3772,N_3296,N_3488);
xor U3773 (N_3773,N_3335,N_3461);
xor U3774 (N_3774,N_3188,N_3291);
nand U3775 (N_3775,N_3309,N_3124);
xor U3776 (N_3776,N_3244,N_3440);
nor U3777 (N_3777,N_3347,N_3192);
or U3778 (N_3778,N_3211,N_3158);
nand U3779 (N_3779,N_3199,N_3209);
and U3780 (N_3780,N_3173,N_3026);
and U3781 (N_3781,N_3356,N_3227);
xnor U3782 (N_3782,N_3064,N_3345);
xnor U3783 (N_3783,N_3403,N_3133);
nor U3784 (N_3784,N_3094,N_3408);
nor U3785 (N_3785,N_3491,N_3442);
nor U3786 (N_3786,N_3194,N_3448);
nand U3787 (N_3787,N_3456,N_3066);
nand U3788 (N_3788,N_3122,N_3036);
nor U3789 (N_3789,N_3085,N_3070);
or U3790 (N_3790,N_3444,N_3382);
nor U3791 (N_3791,N_3031,N_3027);
and U3792 (N_3792,N_3251,N_3083);
xor U3793 (N_3793,N_3481,N_3446);
and U3794 (N_3794,N_3145,N_3055);
nor U3795 (N_3795,N_3485,N_3349);
xor U3796 (N_3796,N_3333,N_3147);
or U3797 (N_3797,N_3061,N_3326);
nor U3798 (N_3798,N_3159,N_3464);
and U3799 (N_3799,N_3188,N_3161);
and U3800 (N_3800,N_3290,N_3402);
nor U3801 (N_3801,N_3101,N_3361);
xor U3802 (N_3802,N_3391,N_3204);
and U3803 (N_3803,N_3403,N_3269);
or U3804 (N_3804,N_3344,N_3449);
xnor U3805 (N_3805,N_3153,N_3416);
or U3806 (N_3806,N_3427,N_3482);
and U3807 (N_3807,N_3369,N_3000);
nand U3808 (N_3808,N_3128,N_3196);
or U3809 (N_3809,N_3212,N_3219);
nor U3810 (N_3810,N_3080,N_3491);
and U3811 (N_3811,N_3358,N_3078);
nor U3812 (N_3812,N_3293,N_3374);
nand U3813 (N_3813,N_3267,N_3175);
nand U3814 (N_3814,N_3102,N_3467);
or U3815 (N_3815,N_3338,N_3172);
nor U3816 (N_3816,N_3127,N_3409);
xnor U3817 (N_3817,N_3059,N_3019);
or U3818 (N_3818,N_3191,N_3199);
nand U3819 (N_3819,N_3047,N_3234);
or U3820 (N_3820,N_3429,N_3227);
and U3821 (N_3821,N_3037,N_3497);
or U3822 (N_3822,N_3221,N_3104);
nand U3823 (N_3823,N_3371,N_3473);
nor U3824 (N_3824,N_3145,N_3426);
and U3825 (N_3825,N_3203,N_3346);
nor U3826 (N_3826,N_3381,N_3269);
and U3827 (N_3827,N_3309,N_3299);
nand U3828 (N_3828,N_3136,N_3148);
and U3829 (N_3829,N_3244,N_3310);
nand U3830 (N_3830,N_3147,N_3324);
and U3831 (N_3831,N_3134,N_3199);
xnor U3832 (N_3832,N_3387,N_3215);
or U3833 (N_3833,N_3464,N_3239);
or U3834 (N_3834,N_3258,N_3277);
nor U3835 (N_3835,N_3368,N_3094);
xnor U3836 (N_3836,N_3321,N_3005);
nand U3837 (N_3837,N_3191,N_3162);
xnor U3838 (N_3838,N_3376,N_3339);
xnor U3839 (N_3839,N_3342,N_3437);
or U3840 (N_3840,N_3173,N_3062);
nand U3841 (N_3841,N_3466,N_3025);
or U3842 (N_3842,N_3263,N_3218);
nor U3843 (N_3843,N_3367,N_3093);
and U3844 (N_3844,N_3475,N_3451);
or U3845 (N_3845,N_3017,N_3078);
and U3846 (N_3846,N_3202,N_3191);
nor U3847 (N_3847,N_3493,N_3356);
and U3848 (N_3848,N_3013,N_3497);
nor U3849 (N_3849,N_3018,N_3414);
xnor U3850 (N_3850,N_3431,N_3404);
and U3851 (N_3851,N_3411,N_3084);
nor U3852 (N_3852,N_3488,N_3447);
and U3853 (N_3853,N_3288,N_3113);
xor U3854 (N_3854,N_3282,N_3448);
nand U3855 (N_3855,N_3378,N_3011);
and U3856 (N_3856,N_3226,N_3396);
nor U3857 (N_3857,N_3310,N_3482);
nand U3858 (N_3858,N_3243,N_3471);
or U3859 (N_3859,N_3366,N_3417);
and U3860 (N_3860,N_3334,N_3401);
nand U3861 (N_3861,N_3358,N_3291);
or U3862 (N_3862,N_3189,N_3375);
xnor U3863 (N_3863,N_3429,N_3479);
and U3864 (N_3864,N_3157,N_3482);
and U3865 (N_3865,N_3341,N_3246);
xnor U3866 (N_3866,N_3333,N_3257);
nor U3867 (N_3867,N_3341,N_3406);
xor U3868 (N_3868,N_3327,N_3212);
xor U3869 (N_3869,N_3029,N_3164);
xnor U3870 (N_3870,N_3224,N_3095);
and U3871 (N_3871,N_3180,N_3021);
or U3872 (N_3872,N_3430,N_3483);
nand U3873 (N_3873,N_3077,N_3378);
nand U3874 (N_3874,N_3355,N_3202);
nor U3875 (N_3875,N_3168,N_3224);
xor U3876 (N_3876,N_3053,N_3398);
or U3877 (N_3877,N_3331,N_3202);
nand U3878 (N_3878,N_3481,N_3268);
nor U3879 (N_3879,N_3163,N_3231);
and U3880 (N_3880,N_3140,N_3036);
xor U3881 (N_3881,N_3327,N_3439);
or U3882 (N_3882,N_3023,N_3402);
nand U3883 (N_3883,N_3265,N_3419);
nor U3884 (N_3884,N_3393,N_3361);
and U3885 (N_3885,N_3232,N_3391);
xor U3886 (N_3886,N_3489,N_3271);
nand U3887 (N_3887,N_3047,N_3001);
and U3888 (N_3888,N_3185,N_3127);
xnor U3889 (N_3889,N_3247,N_3290);
xnor U3890 (N_3890,N_3139,N_3152);
xor U3891 (N_3891,N_3436,N_3493);
or U3892 (N_3892,N_3015,N_3395);
xnor U3893 (N_3893,N_3244,N_3138);
nand U3894 (N_3894,N_3242,N_3082);
or U3895 (N_3895,N_3160,N_3118);
and U3896 (N_3896,N_3037,N_3383);
or U3897 (N_3897,N_3459,N_3150);
nand U3898 (N_3898,N_3074,N_3463);
xor U3899 (N_3899,N_3142,N_3373);
and U3900 (N_3900,N_3323,N_3292);
xor U3901 (N_3901,N_3226,N_3054);
nor U3902 (N_3902,N_3000,N_3263);
or U3903 (N_3903,N_3124,N_3147);
nand U3904 (N_3904,N_3357,N_3026);
xor U3905 (N_3905,N_3169,N_3312);
and U3906 (N_3906,N_3463,N_3380);
and U3907 (N_3907,N_3354,N_3431);
xor U3908 (N_3908,N_3262,N_3385);
nand U3909 (N_3909,N_3405,N_3440);
nand U3910 (N_3910,N_3120,N_3250);
xnor U3911 (N_3911,N_3289,N_3041);
nor U3912 (N_3912,N_3142,N_3297);
or U3913 (N_3913,N_3452,N_3160);
or U3914 (N_3914,N_3369,N_3074);
nor U3915 (N_3915,N_3391,N_3327);
nor U3916 (N_3916,N_3419,N_3095);
nor U3917 (N_3917,N_3306,N_3007);
and U3918 (N_3918,N_3192,N_3087);
and U3919 (N_3919,N_3061,N_3053);
and U3920 (N_3920,N_3028,N_3286);
xnor U3921 (N_3921,N_3259,N_3008);
or U3922 (N_3922,N_3045,N_3055);
nand U3923 (N_3923,N_3201,N_3004);
nand U3924 (N_3924,N_3117,N_3022);
nor U3925 (N_3925,N_3175,N_3296);
or U3926 (N_3926,N_3401,N_3203);
nor U3927 (N_3927,N_3304,N_3168);
and U3928 (N_3928,N_3112,N_3283);
and U3929 (N_3929,N_3000,N_3059);
or U3930 (N_3930,N_3262,N_3329);
and U3931 (N_3931,N_3363,N_3018);
nand U3932 (N_3932,N_3392,N_3371);
nor U3933 (N_3933,N_3411,N_3232);
nand U3934 (N_3934,N_3406,N_3157);
nor U3935 (N_3935,N_3362,N_3331);
nor U3936 (N_3936,N_3010,N_3245);
nor U3937 (N_3937,N_3286,N_3347);
or U3938 (N_3938,N_3196,N_3425);
or U3939 (N_3939,N_3041,N_3024);
or U3940 (N_3940,N_3195,N_3489);
and U3941 (N_3941,N_3001,N_3177);
nand U3942 (N_3942,N_3349,N_3263);
nand U3943 (N_3943,N_3228,N_3490);
and U3944 (N_3944,N_3162,N_3188);
and U3945 (N_3945,N_3170,N_3438);
and U3946 (N_3946,N_3333,N_3498);
nand U3947 (N_3947,N_3489,N_3487);
or U3948 (N_3948,N_3365,N_3061);
xnor U3949 (N_3949,N_3383,N_3377);
nor U3950 (N_3950,N_3192,N_3176);
and U3951 (N_3951,N_3452,N_3049);
nor U3952 (N_3952,N_3297,N_3434);
xnor U3953 (N_3953,N_3005,N_3214);
and U3954 (N_3954,N_3199,N_3127);
nand U3955 (N_3955,N_3116,N_3001);
and U3956 (N_3956,N_3110,N_3227);
and U3957 (N_3957,N_3025,N_3150);
nand U3958 (N_3958,N_3432,N_3224);
or U3959 (N_3959,N_3398,N_3303);
xnor U3960 (N_3960,N_3287,N_3331);
and U3961 (N_3961,N_3236,N_3104);
and U3962 (N_3962,N_3000,N_3362);
nand U3963 (N_3963,N_3254,N_3123);
and U3964 (N_3964,N_3078,N_3213);
nor U3965 (N_3965,N_3449,N_3475);
or U3966 (N_3966,N_3249,N_3232);
xor U3967 (N_3967,N_3010,N_3026);
and U3968 (N_3968,N_3342,N_3401);
xor U3969 (N_3969,N_3494,N_3353);
nor U3970 (N_3970,N_3179,N_3100);
or U3971 (N_3971,N_3321,N_3304);
nand U3972 (N_3972,N_3308,N_3150);
or U3973 (N_3973,N_3381,N_3022);
nand U3974 (N_3974,N_3372,N_3383);
or U3975 (N_3975,N_3444,N_3007);
nor U3976 (N_3976,N_3137,N_3325);
or U3977 (N_3977,N_3339,N_3360);
xnor U3978 (N_3978,N_3399,N_3156);
and U3979 (N_3979,N_3227,N_3133);
xnor U3980 (N_3980,N_3389,N_3237);
xor U3981 (N_3981,N_3163,N_3372);
and U3982 (N_3982,N_3340,N_3348);
nand U3983 (N_3983,N_3178,N_3369);
or U3984 (N_3984,N_3106,N_3019);
and U3985 (N_3985,N_3158,N_3194);
nand U3986 (N_3986,N_3464,N_3026);
or U3987 (N_3987,N_3304,N_3080);
and U3988 (N_3988,N_3457,N_3303);
and U3989 (N_3989,N_3038,N_3121);
xor U3990 (N_3990,N_3157,N_3132);
and U3991 (N_3991,N_3456,N_3474);
or U3992 (N_3992,N_3421,N_3231);
and U3993 (N_3993,N_3189,N_3044);
xnor U3994 (N_3994,N_3108,N_3146);
xnor U3995 (N_3995,N_3114,N_3034);
xnor U3996 (N_3996,N_3376,N_3299);
nand U3997 (N_3997,N_3490,N_3444);
nor U3998 (N_3998,N_3123,N_3067);
nor U3999 (N_3999,N_3039,N_3327);
nand U4000 (N_4000,N_3742,N_3777);
nor U4001 (N_4001,N_3881,N_3971);
nor U4002 (N_4002,N_3940,N_3835);
or U4003 (N_4003,N_3723,N_3868);
xnor U4004 (N_4004,N_3876,N_3690);
nand U4005 (N_4005,N_3936,N_3529);
and U4006 (N_4006,N_3902,N_3925);
nand U4007 (N_4007,N_3806,N_3755);
or U4008 (N_4008,N_3786,N_3536);
nand U4009 (N_4009,N_3981,N_3888);
nor U4010 (N_4010,N_3696,N_3964);
or U4011 (N_4011,N_3886,N_3804);
xor U4012 (N_4012,N_3930,N_3542);
nand U4013 (N_4013,N_3519,N_3524);
nor U4014 (N_4014,N_3707,N_3657);
nor U4015 (N_4015,N_3992,N_3669);
and U4016 (N_4016,N_3679,N_3824);
nor U4017 (N_4017,N_3948,N_3665);
and U4018 (N_4018,N_3721,N_3820);
xnor U4019 (N_4019,N_3602,N_3763);
nor U4020 (N_4020,N_3705,N_3676);
nand U4021 (N_4021,N_3849,N_3965);
and U4022 (N_4022,N_3697,N_3648);
and U4023 (N_4023,N_3923,N_3924);
nor U4024 (N_4024,N_3810,N_3644);
nor U4025 (N_4025,N_3984,N_3689);
nor U4026 (N_4026,N_3627,N_3630);
nand U4027 (N_4027,N_3727,N_3905);
xnor U4028 (N_4028,N_3512,N_3551);
nor U4029 (N_4029,N_3634,N_3548);
or U4030 (N_4030,N_3867,N_3584);
nor U4031 (N_4031,N_3739,N_3861);
or U4032 (N_4032,N_3507,N_3539);
xor U4033 (N_4033,N_3660,N_3842);
nand U4034 (N_4034,N_3891,N_3526);
or U4035 (N_4035,N_3558,N_3675);
xor U4036 (N_4036,N_3744,N_3972);
nor U4037 (N_4037,N_3811,N_3621);
xnor U4038 (N_4038,N_3698,N_3614);
nand U4039 (N_4039,N_3986,N_3822);
or U4040 (N_4040,N_3979,N_3784);
nand U4041 (N_4041,N_3569,N_3762);
and U4042 (N_4042,N_3625,N_3737);
or U4043 (N_4043,N_3833,N_3677);
or U4044 (N_4044,N_3795,N_3870);
nand U4045 (N_4045,N_3903,N_3642);
nand U4046 (N_4046,N_3785,N_3720);
xnor U4047 (N_4047,N_3606,N_3758);
nor U4048 (N_4048,N_3793,N_3543);
and U4049 (N_4049,N_3946,N_3504);
or U4050 (N_4050,N_3559,N_3699);
or U4051 (N_4051,N_3717,N_3538);
and U4052 (N_4052,N_3848,N_3666);
nand U4053 (N_4053,N_3686,N_3568);
nor U4054 (N_4054,N_3550,N_3920);
and U4055 (N_4055,N_3658,N_3729);
xnor U4056 (N_4056,N_3780,N_3670);
nand U4057 (N_4057,N_3791,N_3710);
nor U4058 (N_4058,N_3748,N_3577);
nor U4059 (N_4059,N_3818,N_3672);
and U4060 (N_4060,N_3706,N_3546);
and U4061 (N_4061,N_3598,N_3893);
and U4062 (N_4062,N_3638,N_3917);
xnor U4063 (N_4063,N_3600,N_3812);
xnor U4064 (N_4064,N_3772,N_3899);
nor U4065 (N_4065,N_3643,N_3572);
nand U4066 (N_4066,N_3574,N_3622);
and U4067 (N_4067,N_3927,N_3667);
or U4068 (N_4068,N_3735,N_3975);
and U4069 (N_4069,N_3910,N_3592);
nor U4070 (N_4070,N_3631,N_3637);
xor U4071 (N_4071,N_3553,N_3745);
nor U4072 (N_4072,N_3957,N_3581);
and U4073 (N_4073,N_3513,N_3534);
nor U4074 (N_4074,N_3884,N_3852);
nand U4075 (N_4075,N_3915,N_3912);
or U4076 (N_4076,N_3753,N_3839);
or U4077 (N_4077,N_3950,N_3716);
or U4078 (N_4078,N_3759,N_3809);
and U4079 (N_4079,N_3654,N_3864);
nand U4080 (N_4080,N_3547,N_3599);
xor U4081 (N_4081,N_3858,N_3766);
or U4082 (N_4082,N_3929,N_3846);
or U4083 (N_4083,N_3647,N_3503);
nor U4084 (N_4084,N_3952,N_3828);
or U4085 (N_4085,N_3892,N_3770);
xnor U4086 (N_4086,N_3983,N_3540);
or U4087 (N_4087,N_3958,N_3961);
and U4088 (N_4088,N_3973,N_3595);
nor U4089 (N_4089,N_3969,N_3904);
and U4090 (N_4090,N_3555,N_3500);
nand U4091 (N_4091,N_3573,N_3712);
xnor U4092 (N_4092,N_3931,N_3640);
xnor U4093 (N_4093,N_3943,N_3635);
or U4094 (N_4094,N_3545,N_3794);
nand U4095 (N_4095,N_3875,N_3510);
xnor U4096 (N_4096,N_3750,N_3781);
or U4097 (N_4097,N_3819,N_3956);
or U4098 (N_4098,N_3731,N_3934);
xnor U4099 (N_4099,N_3531,N_3516);
and U4100 (N_4100,N_3563,N_3857);
nor U4101 (N_4101,N_3985,N_3798);
xor U4102 (N_4102,N_3808,N_3757);
nand U4103 (N_4103,N_3799,N_3709);
nor U4104 (N_4104,N_3556,N_3746);
and U4105 (N_4105,N_3837,N_3995);
and U4106 (N_4106,N_3562,N_3702);
nor U4107 (N_4107,N_3575,N_3724);
and U4108 (N_4108,N_3501,N_3692);
nor U4109 (N_4109,N_3897,N_3653);
xor U4110 (N_4110,N_3756,N_3880);
or U4111 (N_4111,N_3775,N_3589);
or U4112 (N_4112,N_3741,N_3652);
nand U4113 (N_4113,N_3518,N_3747);
and U4114 (N_4114,N_3845,N_3722);
or U4115 (N_4115,N_3728,N_3982);
nand U4116 (N_4116,N_3841,N_3951);
xor U4117 (N_4117,N_3738,N_3919);
nor U4118 (N_4118,N_3769,N_3678);
nor U4119 (N_4119,N_3871,N_3847);
or U4120 (N_4120,N_3998,N_3913);
and U4121 (N_4121,N_3792,N_3655);
nand U4122 (N_4122,N_3552,N_3645);
nand U4123 (N_4123,N_3898,N_3856);
or U4124 (N_4124,N_3715,N_3609);
nor U4125 (N_4125,N_3520,N_3901);
and U4126 (N_4126,N_3937,N_3761);
nand U4127 (N_4127,N_3854,N_3869);
or U4128 (N_4128,N_3713,N_3585);
nand U4129 (N_4129,N_3887,N_3734);
xor U4130 (N_4130,N_3586,N_3607);
or U4131 (N_4131,N_3821,N_3541);
xor U4132 (N_4132,N_3743,N_3908);
and U4133 (N_4133,N_3576,N_3850);
xnor U4134 (N_4134,N_3521,N_3608);
nand U4135 (N_4135,N_3671,N_3900);
nand U4136 (N_4136,N_3649,N_3774);
or U4137 (N_4137,N_3523,N_3840);
nor U4138 (N_4138,N_3974,N_3588);
xor U4139 (N_4139,N_3883,N_3947);
and U4140 (N_4140,N_3853,N_3954);
nor U4141 (N_4141,N_3613,N_3687);
and U4142 (N_4142,N_3966,N_3612);
or U4143 (N_4143,N_3796,N_3719);
xor U4144 (N_4144,N_3656,N_3522);
nor U4145 (N_4145,N_3767,N_3661);
or U4146 (N_4146,N_3610,N_3790);
and U4147 (N_4147,N_3980,N_3659);
and U4148 (N_4148,N_3859,N_3771);
and U4149 (N_4149,N_3663,N_3506);
and U4150 (N_4150,N_3571,N_3977);
and U4151 (N_4151,N_3616,N_3967);
xor U4152 (N_4152,N_3801,N_3527);
nor U4153 (N_4153,N_3560,N_3693);
and U4154 (N_4154,N_3619,N_3752);
nand U4155 (N_4155,N_3681,N_3914);
nor U4156 (N_4156,N_3736,N_3844);
nand U4157 (N_4157,N_3528,N_3933);
and U4158 (N_4158,N_3578,N_3830);
nand U4159 (N_4159,N_3911,N_3593);
or U4160 (N_4160,N_3673,N_3829);
or U4161 (N_4161,N_3511,N_3641);
nor U4162 (N_4162,N_3976,N_3565);
xor U4163 (N_4163,N_3909,N_3749);
or U4164 (N_4164,N_3800,N_3895);
xor U4165 (N_4165,N_3962,N_3873);
or U4166 (N_4166,N_3508,N_3872);
nor U4167 (N_4167,N_3685,N_3751);
nand U4168 (N_4168,N_3580,N_3623);
nand U4169 (N_4169,N_3944,N_3726);
or U4170 (N_4170,N_3683,N_3968);
and U4171 (N_4171,N_3587,N_3926);
nor U4172 (N_4172,N_3618,N_3544);
and U4173 (N_4173,N_3561,N_3814);
and U4174 (N_4174,N_3803,N_3664);
or U4175 (N_4175,N_3651,N_3788);
nand U4176 (N_4176,N_3994,N_3918);
nand U4177 (N_4177,N_3955,N_3807);
nand U4178 (N_4178,N_3636,N_3805);
or U4179 (N_4179,N_3557,N_3832);
and U4180 (N_4180,N_3570,N_3953);
or U4181 (N_4181,N_3760,N_3620);
xor U4182 (N_4182,N_3894,N_3714);
xor U4183 (N_4183,N_3650,N_3999);
nand U4184 (N_4184,N_3684,N_3502);
nor U4185 (N_4185,N_3896,N_3783);
nand U4186 (N_4186,N_3533,N_3970);
nand U4187 (N_4187,N_3789,N_3567);
and U4188 (N_4188,N_3802,N_3855);
xnor U4189 (N_4189,N_3626,N_3554);
or U4190 (N_4190,N_3776,N_3691);
xnor U4191 (N_4191,N_3990,N_3989);
nand U4192 (N_4192,N_3996,N_3532);
and U4193 (N_4193,N_3997,N_3773);
and U4194 (N_4194,N_3674,N_3711);
nand U4195 (N_4195,N_3597,N_3725);
or U4196 (N_4196,N_3765,N_3708);
nor U4197 (N_4197,N_3514,N_3718);
and U4198 (N_4198,N_3525,N_3566);
xnor U4199 (N_4199,N_3831,N_3703);
xnor U4200 (N_4200,N_3787,N_3991);
and U4201 (N_4201,N_3701,N_3617);
or U4202 (N_4202,N_3704,N_3843);
and U4203 (N_4203,N_3993,N_3695);
nor U4204 (N_4204,N_3764,N_3509);
and U4205 (N_4205,N_3963,N_3959);
nor U4206 (N_4206,N_3945,N_3604);
or U4207 (N_4207,N_3863,N_3987);
or U4208 (N_4208,N_3564,N_3879);
xnor U4209 (N_4209,N_3916,N_3505);
nand U4210 (N_4210,N_3732,N_3932);
xnor U4211 (N_4211,N_3632,N_3688);
nor U4212 (N_4212,N_3834,N_3633);
or U4213 (N_4213,N_3938,N_3583);
and U4214 (N_4214,N_3815,N_3885);
xnor U4215 (N_4215,N_3823,N_3537);
or U4216 (N_4216,N_3860,N_3935);
and U4217 (N_4217,N_3579,N_3827);
nand U4218 (N_4218,N_3939,N_3549);
or U4219 (N_4219,N_3639,N_3889);
xor U4220 (N_4220,N_3668,N_3906);
nor U4221 (N_4221,N_3836,N_3694);
and U4222 (N_4222,N_3624,N_3817);
nand U4223 (N_4223,N_3662,N_3682);
and U4224 (N_4224,N_3605,N_3768);
nand U4225 (N_4225,N_3535,N_3596);
nand U4226 (N_4226,N_3960,N_3582);
nor U4227 (N_4227,N_3878,N_3730);
or U4228 (N_4228,N_3590,N_3611);
or U4229 (N_4229,N_3825,N_3646);
and U4230 (N_4230,N_3942,N_3591);
or U4231 (N_4231,N_3700,N_3921);
nor U4232 (N_4232,N_3740,N_3754);
nand U4233 (N_4233,N_3779,N_3922);
nor U4234 (N_4234,N_3866,N_3778);
or U4235 (N_4235,N_3928,N_3949);
nor U4236 (N_4236,N_3877,N_3882);
nand U4237 (N_4237,N_3594,N_3629);
nand U4238 (N_4238,N_3615,N_3515);
or U4239 (N_4239,N_3890,N_3601);
and U4240 (N_4240,N_3816,N_3517);
xor U4241 (N_4241,N_3941,N_3628);
nand U4242 (N_4242,N_3603,N_3988);
and U4243 (N_4243,N_3851,N_3874);
and U4244 (N_4244,N_3797,N_3865);
nand U4245 (N_4245,N_3862,N_3838);
or U4246 (N_4246,N_3530,N_3978);
nand U4247 (N_4247,N_3680,N_3782);
or U4248 (N_4248,N_3826,N_3733);
and U4249 (N_4249,N_3907,N_3813);
xnor U4250 (N_4250,N_3724,N_3948);
nand U4251 (N_4251,N_3680,N_3821);
and U4252 (N_4252,N_3622,N_3605);
nor U4253 (N_4253,N_3630,N_3905);
nor U4254 (N_4254,N_3584,N_3546);
nor U4255 (N_4255,N_3548,N_3547);
xnor U4256 (N_4256,N_3726,N_3667);
nand U4257 (N_4257,N_3542,N_3595);
and U4258 (N_4258,N_3793,N_3901);
nand U4259 (N_4259,N_3781,N_3563);
or U4260 (N_4260,N_3555,N_3766);
nand U4261 (N_4261,N_3705,N_3742);
nor U4262 (N_4262,N_3675,N_3524);
and U4263 (N_4263,N_3678,N_3554);
or U4264 (N_4264,N_3614,N_3670);
or U4265 (N_4265,N_3547,N_3698);
or U4266 (N_4266,N_3839,N_3745);
nand U4267 (N_4267,N_3748,N_3663);
nor U4268 (N_4268,N_3871,N_3766);
nor U4269 (N_4269,N_3943,N_3667);
xnor U4270 (N_4270,N_3640,N_3661);
nor U4271 (N_4271,N_3833,N_3531);
xnor U4272 (N_4272,N_3608,N_3656);
and U4273 (N_4273,N_3516,N_3873);
nor U4274 (N_4274,N_3562,N_3737);
nor U4275 (N_4275,N_3545,N_3795);
nor U4276 (N_4276,N_3862,N_3641);
nand U4277 (N_4277,N_3947,N_3831);
nor U4278 (N_4278,N_3568,N_3888);
nand U4279 (N_4279,N_3563,N_3560);
xnor U4280 (N_4280,N_3674,N_3598);
and U4281 (N_4281,N_3574,N_3778);
nor U4282 (N_4282,N_3740,N_3757);
nor U4283 (N_4283,N_3806,N_3856);
nand U4284 (N_4284,N_3700,N_3948);
or U4285 (N_4285,N_3783,N_3631);
xor U4286 (N_4286,N_3863,N_3551);
nand U4287 (N_4287,N_3861,N_3879);
nand U4288 (N_4288,N_3921,N_3626);
nand U4289 (N_4289,N_3653,N_3537);
and U4290 (N_4290,N_3740,N_3636);
nor U4291 (N_4291,N_3517,N_3965);
or U4292 (N_4292,N_3598,N_3755);
or U4293 (N_4293,N_3921,N_3721);
nand U4294 (N_4294,N_3546,N_3857);
or U4295 (N_4295,N_3842,N_3716);
nor U4296 (N_4296,N_3592,N_3673);
or U4297 (N_4297,N_3788,N_3572);
and U4298 (N_4298,N_3958,N_3630);
and U4299 (N_4299,N_3648,N_3862);
nand U4300 (N_4300,N_3576,N_3947);
xnor U4301 (N_4301,N_3937,N_3668);
and U4302 (N_4302,N_3888,N_3920);
or U4303 (N_4303,N_3511,N_3822);
or U4304 (N_4304,N_3655,N_3791);
nand U4305 (N_4305,N_3828,N_3861);
nor U4306 (N_4306,N_3644,N_3760);
and U4307 (N_4307,N_3891,N_3839);
or U4308 (N_4308,N_3814,N_3880);
xnor U4309 (N_4309,N_3833,N_3947);
or U4310 (N_4310,N_3988,N_3661);
nand U4311 (N_4311,N_3888,N_3606);
xnor U4312 (N_4312,N_3520,N_3664);
or U4313 (N_4313,N_3759,N_3616);
xor U4314 (N_4314,N_3767,N_3624);
nor U4315 (N_4315,N_3531,N_3602);
xor U4316 (N_4316,N_3592,N_3684);
and U4317 (N_4317,N_3552,N_3942);
or U4318 (N_4318,N_3826,N_3858);
xnor U4319 (N_4319,N_3935,N_3869);
nand U4320 (N_4320,N_3844,N_3723);
nor U4321 (N_4321,N_3761,N_3931);
and U4322 (N_4322,N_3893,N_3618);
nand U4323 (N_4323,N_3723,N_3668);
nand U4324 (N_4324,N_3711,N_3976);
nor U4325 (N_4325,N_3541,N_3787);
xnor U4326 (N_4326,N_3794,N_3581);
nand U4327 (N_4327,N_3627,N_3575);
or U4328 (N_4328,N_3622,N_3581);
nand U4329 (N_4329,N_3655,N_3595);
or U4330 (N_4330,N_3601,N_3602);
nand U4331 (N_4331,N_3644,N_3737);
and U4332 (N_4332,N_3791,N_3938);
nand U4333 (N_4333,N_3863,N_3916);
nand U4334 (N_4334,N_3743,N_3850);
nor U4335 (N_4335,N_3849,N_3578);
and U4336 (N_4336,N_3843,N_3942);
nand U4337 (N_4337,N_3581,N_3986);
nor U4338 (N_4338,N_3859,N_3929);
xor U4339 (N_4339,N_3819,N_3984);
nor U4340 (N_4340,N_3631,N_3727);
or U4341 (N_4341,N_3966,N_3809);
nand U4342 (N_4342,N_3546,N_3799);
xnor U4343 (N_4343,N_3953,N_3626);
nand U4344 (N_4344,N_3860,N_3817);
nand U4345 (N_4345,N_3943,N_3652);
nor U4346 (N_4346,N_3994,N_3752);
or U4347 (N_4347,N_3596,N_3608);
nor U4348 (N_4348,N_3805,N_3789);
or U4349 (N_4349,N_3940,N_3545);
and U4350 (N_4350,N_3789,N_3982);
nand U4351 (N_4351,N_3897,N_3817);
xor U4352 (N_4352,N_3718,N_3899);
or U4353 (N_4353,N_3994,N_3778);
nand U4354 (N_4354,N_3718,N_3666);
and U4355 (N_4355,N_3707,N_3966);
and U4356 (N_4356,N_3963,N_3933);
nand U4357 (N_4357,N_3529,N_3798);
xor U4358 (N_4358,N_3707,N_3558);
and U4359 (N_4359,N_3628,N_3638);
nand U4360 (N_4360,N_3558,N_3829);
or U4361 (N_4361,N_3890,N_3540);
xor U4362 (N_4362,N_3614,N_3542);
xnor U4363 (N_4363,N_3685,N_3683);
nor U4364 (N_4364,N_3542,N_3837);
nand U4365 (N_4365,N_3620,N_3792);
and U4366 (N_4366,N_3619,N_3962);
nand U4367 (N_4367,N_3805,N_3782);
and U4368 (N_4368,N_3939,N_3783);
xnor U4369 (N_4369,N_3904,N_3975);
or U4370 (N_4370,N_3943,N_3614);
xor U4371 (N_4371,N_3602,N_3994);
or U4372 (N_4372,N_3713,N_3885);
xnor U4373 (N_4373,N_3785,N_3834);
nand U4374 (N_4374,N_3648,N_3554);
nor U4375 (N_4375,N_3781,N_3692);
and U4376 (N_4376,N_3908,N_3945);
nor U4377 (N_4377,N_3948,N_3989);
nor U4378 (N_4378,N_3513,N_3599);
or U4379 (N_4379,N_3997,N_3510);
and U4380 (N_4380,N_3505,N_3864);
xnor U4381 (N_4381,N_3816,N_3659);
or U4382 (N_4382,N_3818,N_3522);
xnor U4383 (N_4383,N_3607,N_3977);
nand U4384 (N_4384,N_3728,N_3833);
xnor U4385 (N_4385,N_3514,N_3666);
nor U4386 (N_4386,N_3941,N_3826);
and U4387 (N_4387,N_3890,N_3801);
or U4388 (N_4388,N_3855,N_3946);
and U4389 (N_4389,N_3526,N_3577);
xor U4390 (N_4390,N_3886,N_3717);
and U4391 (N_4391,N_3813,N_3680);
nor U4392 (N_4392,N_3954,N_3938);
nor U4393 (N_4393,N_3585,N_3644);
xnor U4394 (N_4394,N_3732,N_3664);
and U4395 (N_4395,N_3563,N_3612);
xnor U4396 (N_4396,N_3724,N_3528);
xor U4397 (N_4397,N_3972,N_3913);
nor U4398 (N_4398,N_3647,N_3563);
nand U4399 (N_4399,N_3512,N_3796);
nand U4400 (N_4400,N_3988,N_3523);
nand U4401 (N_4401,N_3826,N_3516);
nand U4402 (N_4402,N_3828,N_3758);
and U4403 (N_4403,N_3924,N_3583);
nand U4404 (N_4404,N_3543,N_3937);
or U4405 (N_4405,N_3826,N_3847);
nor U4406 (N_4406,N_3580,N_3634);
nand U4407 (N_4407,N_3964,N_3851);
and U4408 (N_4408,N_3543,N_3963);
and U4409 (N_4409,N_3534,N_3963);
and U4410 (N_4410,N_3969,N_3711);
or U4411 (N_4411,N_3868,N_3968);
and U4412 (N_4412,N_3980,N_3866);
xnor U4413 (N_4413,N_3973,N_3752);
xor U4414 (N_4414,N_3789,N_3987);
xnor U4415 (N_4415,N_3733,N_3869);
or U4416 (N_4416,N_3729,N_3841);
and U4417 (N_4417,N_3853,N_3606);
xnor U4418 (N_4418,N_3793,N_3728);
or U4419 (N_4419,N_3610,N_3652);
nor U4420 (N_4420,N_3772,N_3760);
nand U4421 (N_4421,N_3661,N_3555);
and U4422 (N_4422,N_3975,N_3621);
xnor U4423 (N_4423,N_3571,N_3588);
nand U4424 (N_4424,N_3673,N_3579);
xnor U4425 (N_4425,N_3598,N_3725);
nand U4426 (N_4426,N_3659,N_3695);
or U4427 (N_4427,N_3620,N_3606);
nand U4428 (N_4428,N_3705,N_3504);
xor U4429 (N_4429,N_3579,N_3986);
and U4430 (N_4430,N_3992,N_3855);
xnor U4431 (N_4431,N_3682,N_3676);
and U4432 (N_4432,N_3721,N_3513);
nor U4433 (N_4433,N_3927,N_3505);
or U4434 (N_4434,N_3553,N_3769);
nor U4435 (N_4435,N_3575,N_3985);
and U4436 (N_4436,N_3585,N_3500);
xnor U4437 (N_4437,N_3636,N_3787);
nand U4438 (N_4438,N_3861,N_3974);
and U4439 (N_4439,N_3989,N_3703);
or U4440 (N_4440,N_3886,N_3589);
nand U4441 (N_4441,N_3510,N_3702);
nand U4442 (N_4442,N_3884,N_3930);
nor U4443 (N_4443,N_3911,N_3586);
nor U4444 (N_4444,N_3575,N_3957);
and U4445 (N_4445,N_3588,N_3660);
nand U4446 (N_4446,N_3689,N_3786);
and U4447 (N_4447,N_3803,N_3863);
nor U4448 (N_4448,N_3599,N_3729);
nor U4449 (N_4449,N_3674,N_3546);
or U4450 (N_4450,N_3604,N_3552);
and U4451 (N_4451,N_3619,N_3745);
nor U4452 (N_4452,N_3974,N_3939);
or U4453 (N_4453,N_3814,N_3665);
nor U4454 (N_4454,N_3662,N_3860);
nor U4455 (N_4455,N_3999,N_3975);
nand U4456 (N_4456,N_3752,N_3708);
nor U4457 (N_4457,N_3670,N_3630);
and U4458 (N_4458,N_3818,N_3745);
nor U4459 (N_4459,N_3738,N_3642);
nor U4460 (N_4460,N_3746,N_3513);
or U4461 (N_4461,N_3687,N_3511);
nor U4462 (N_4462,N_3675,N_3637);
or U4463 (N_4463,N_3731,N_3523);
or U4464 (N_4464,N_3945,N_3587);
nor U4465 (N_4465,N_3839,N_3951);
and U4466 (N_4466,N_3924,N_3575);
or U4467 (N_4467,N_3720,N_3522);
and U4468 (N_4468,N_3610,N_3961);
nand U4469 (N_4469,N_3906,N_3531);
and U4470 (N_4470,N_3985,N_3776);
and U4471 (N_4471,N_3666,N_3685);
nand U4472 (N_4472,N_3550,N_3588);
and U4473 (N_4473,N_3621,N_3698);
and U4474 (N_4474,N_3922,N_3708);
nor U4475 (N_4475,N_3719,N_3906);
nand U4476 (N_4476,N_3949,N_3650);
nand U4477 (N_4477,N_3532,N_3615);
nor U4478 (N_4478,N_3731,N_3770);
nor U4479 (N_4479,N_3785,N_3775);
or U4480 (N_4480,N_3802,N_3633);
xnor U4481 (N_4481,N_3903,N_3806);
or U4482 (N_4482,N_3537,N_3528);
or U4483 (N_4483,N_3795,N_3657);
or U4484 (N_4484,N_3846,N_3738);
nor U4485 (N_4485,N_3524,N_3948);
nand U4486 (N_4486,N_3679,N_3953);
xor U4487 (N_4487,N_3685,N_3600);
nor U4488 (N_4488,N_3548,N_3917);
and U4489 (N_4489,N_3783,N_3856);
nand U4490 (N_4490,N_3831,N_3770);
or U4491 (N_4491,N_3887,N_3778);
xnor U4492 (N_4492,N_3785,N_3721);
xor U4493 (N_4493,N_3999,N_3587);
and U4494 (N_4494,N_3515,N_3972);
or U4495 (N_4495,N_3860,N_3814);
and U4496 (N_4496,N_3865,N_3576);
nand U4497 (N_4497,N_3559,N_3687);
and U4498 (N_4498,N_3502,N_3832);
or U4499 (N_4499,N_3636,N_3743);
and U4500 (N_4500,N_4033,N_4179);
xnor U4501 (N_4501,N_4194,N_4083);
and U4502 (N_4502,N_4116,N_4017);
xnor U4503 (N_4503,N_4485,N_4322);
xor U4504 (N_4504,N_4391,N_4195);
nand U4505 (N_4505,N_4229,N_4117);
nor U4506 (N_4506,N_4041,N_4400);
xor U4507 (N_4507,N_4104,N_4458);
nand U4508 (N_4508,N_4442,N_4415);
and U4509 (N_4509,N_4008,N_4167);
and U4510 (N_4510,N_4106,N_4368);
nor U4511 (N_4511,N_4172,N_4143);
nor U4512 (N_4512,N_4219,N_4363);
nand U4513 (N_4513,N_4005,N_4152);
xor U4514 (N_4514,N_4096,N_4217);
nor U4515 (N_4515,N_4136,N_4147);
xnor U4516 (N_4516,N_4191,N_4207);
xnor U4517 (N_4517,N_4085,N_4262);
nor U4518 (N_4518,N_4252,N_4182);
nor U4519 (N_4519,N_4263,N_4407);
xnor U4520 (N_4520,N_4283,N_4410);
nor U4521 (N_4521,N_4145,N_4066);
or U4522 (N_4522,N_4333,N_4094);
nor U4523 (N_4523,N_4231,N_4393);
nand U4524 (N_4524,N_4251,N_4032);
and U4525 (N_4525,N_4255,N_4111);
nand U4526 (N_4526,N_4164,N_4493);
or U4527 (N_4527,N_4009,N_4277);
nor U4528 (N_4528,N_4370,N_4282);
nand U4529 (N_4529,N_4380,N_4245);
xnor U4530 (N_4530,N_4324,N_4451);
nand U4531 (N_4531,N_4343,N_4284);
and U4532 (N_4532,N_4254,N_4409);
nand U4533 (N_4533,N_4151,N_4062);
nor U4534 (N_4534,N_4134,N_4144);
or U4535 (N_4535,N_4318,N_4181);
nand U4536 (N_4536,N_4024,N_4115);
xor U4537 (N_4537,N_4241,N_4440);
and U4538 (N_4538,N_4259,N_4052);
nor U4539 (N_4539,N_4260,N_4031);
and U4540 (N_4540,N_4108,N_4004);
nor U4541 (N_4541,N_4137,N_4481);
or U4542 (N_4542,N_4430,N_4193);
nor U4543 (N_4543,N_4056,N_4471);
and U4544 (N_4544,N_4023,N_4434);
xnor U4545 (N_4545,N_4296,N_4457);
nor U4546 (N_4546,N_4086,N_4226);
nand U4547 (N_4547,N_4436,N_4265);
and U4548 (N_4548,N_4344,N_4081);
and U4549 (N_4549,N_4311,N_4470);
nor U4550 (N_4550,N_4468,N_4073);
and U4551 (N_4551,N_4015,N_4077);
nand U4552 (N_4552,N_4029,N_4000);
or U4553 (N_4553,N_4315,N_4406);
nor U4554 (N_4554,N_4479,N_4051);
nand U4555 (N_4555,N_4490,N_4121);
nor U4556 (N_4556,N_4221,N_4428);
nor U4557 (N_4557,N_4411,N_4297);
nand U4558 (N_4558,N_4379,N_4261);
or U4559 (N_4559,N_4348,N_4356);
nand U4560 (N_4560,N_4280,N_4359);
and U4561 (N_4561,N_4487,N_4087);
and U4562 (N_4562,N_4088,N_4264);
nand U4563 (N_4563,N_4270,N_4427);
or U4564 (N_4564,N_4466,N_4107);
and U4565 (N_4565,N_4294,N_4192);
nor U4566 (N_4566,N_4090,N_4184);
xor U4567 (N_4567,N_4268,N_4486);
xnor U4568 (N_4568,N_4313,N_4337);
nor U4569 (N_4569,N_4250,N_4199);
or U4570 (N_4570,N_4385,N_4465);
nor U4571 (N_4571,N_4141,N_4330);
and U4572 (N_4572,N_4460,N_4495);
and U4573 (N_4573,N_4446,N_4175);
nand U4574 (N_4574,N_4109,N_4401);
nor U4575 (N_4575,N_4196,N_4371);
nor U4576 (N_4576,N_4257,N_4341);
nand U4577 (N_4577,N_4467,N_4012);
nor U4578 (N_4578,N_4354,N_4010);
or U4579 (N_4579,N_4435,N_4036);
nor U4580 (N_4580,N_4075,N_4156);
and U4581 (N_4581,N_4497,N_4028);
nand U4582 (N_4582,N_4154,N_4477);
xor U4583 (N_4583,N_4149,N_4227);
xor U4584 (N_4584,N_4119,N_4204);
or U4585 (N_4585,N_4059,N_4247);
nand U4586 (N_4586,N_4346,N_4285);
or U4587 (N_4587,N_4068,N_4352);
nand U4588 (N_4588,N_4105,N_4053);
xnor U4589 (N_4589,N_4482,N_4146);
nor U4590 (N_4590,N_4365,N_4367);
and U4591 (N_4591,N_4070,N_4233);
or U4592 (N_4592,N_4431,N_4014);
nand U4593 (N_4593,N_4168,N_4057);
and U4594 (N_4594,N_4473,N_4065);
nor U4595 (N_4595,N_4288,N_4358);
xor U4596 (N_4596,N_4092,N_4441);
or U4597 (N_4597,N_4273,N_4114);
nand U4598 (N_4598,N_4395,N_4040);
xor U4599 (N_4599,N_4498,N_4291);
nand U4600 (N_4600,N_4044,N_4098);
nand U4601 (N_4601,N_4235,N_4128);
xnor U4602 (N_4602,N_4123,N_4148);
and U4603 (N_4603,N_4357,N_4405);
nor U4604 (N_4604,N_4027,N_4491);
and U4605 (N_4605,N_4190,N_4126);
xnor U4606 (N_4606,N_4003,N_4376);
xnor U4607 (N_4607,N_4211,N_4310);
or U4608 (N_4608,N_4183,N_4317);
or U4609 (N_4609,N_4178,N_4323);
nor U4610 (N_4610,N_4278,N_4237);
and U4611 (N_4611,N_4412,N_4418);
xor U4612 (N_4612,N_4054,N_4061);
xor U4613 (N_4613,N_4404,N_4042);
nand U4614 (N_4614,N_4499,N_4093);
or U4615 (N_4615,N_4492,N_4206);
nand U4616 (N_4616,N_4069,N_4214);
nand U4617 (N_4617,N_4329,N_4021);
nor U4618 (N_4618,N_4099,N_4389);
nor U4619 (N_4619,N_4080,N_4048);
or U4620 (N_4620,N_4013,N_4279);
and U4621 (N_4621,N_4290,N_4381);
and U4622 (N_4622,N_4342,N_4177);
and U4623 (N_4623,N_4139,N_4113);
nand U4624 (N_4624,N_4464,N_4131);
or U4625 (N_4625,N_4443,N_4338);
xor U4626 (N_4626,N_4159,N_4225);
nand U4627 (N_4627,N_4349,N_4271);
and U4628 (N_4628,N_4394,N_4138);
or U4629 (N_4629,N_4063,N_4198);
nor U4630 (N_4630,N_4421,N_4266);
and U4631 (N_4631,N_4319,N_4174);
or U4632 (N_4632,N_4132,N_4300);
and U4633 (N_4633,N_4244,N_4034);
xnor U4634 (N_4634,N_4447,N_4292);
or U4635 (N_4635,N_4474,N_4478);
nand U4636 (N_4636,N_4102,N_4320);
xnor U4637 (N_4637,N_4429,N_4223);
xnor U4638 (N_4638,N_4305,N_4176);
nand U4639 (N_4639,N_4188,N_4325);
xor U4640 (N_4640,N_4364,N_4018);
and U4641 (N_4641,N_4150,N_4011);
nor U4642 (N_4642,N_4072,N_4417);
and U4643 (N_4643,N_4459,N_4375);
xnor U4644 (N_4644,N_4450,N_4082);
xnor U4645 (N_4645,N_4396,N_4208);
xnor U4646 (N_4646,N_4216,N_4448);
and U4647 (N_4647,N_4129,N_4248);
nor U4648 (N_4648,N_4307,N_4456);
and U4649 (N_4649,N_4408,N_4373);
nand U4650 (N_4650,N_4162,N_4374);
and U4651 (N_4651,N_4050,N_4331);
nor U4652 (N_4652,N_4202,N_4035);
xor U4653 (N_4653,N_4372,N_4240);
nor U4654 (N_4654,N_4019,N_4232);
xor U4655 (N_4655,N_4392,N_4239);
xnor U4656 (N_4656,N_4045,N_4327);
xor U4657 (N_4657,N_4475,N_4185);
xnor U4658 (N_4658,N_4228,N_4390);
or U4659 (N_4659,N_4306,N_4006);
nand U4660 (N_4660,N_4016,N_4127);
nand U4661 (N_4661,N_4274,N_4308);
or U4662 (N_4662,N_4462,N_4230);
and U4663 (N_4663,N_4142,N_4002);
and U4664 (N_4664,N_4186,N_4432);
nand U4665 (N_4665,N_4347,N_4298);
or U4666 (N_4666,N_4091,N_4449);
and U4667 (N_4667,N_4339,N_4100);
nand U4668 (N_4668,N_4161,N_4488);
nand U4669 (N_4669,N_4334,N_4483);
and U4670 (N_4670,N_4038,N_4416);
and U4671 (N_4671,N_4118,N_4439);
nor U4672 (N_4672,N_4422,N_4209);
xor U4673 (N_4673,N_4160,N_4353);
or U4674 (N_4674,N_4304,N_4419);
and U4675 (N_4675,N_4007,N_4071);
nor U4676 (N_4676,N_4095,N_4130);
nand U4677 (N_4677,N_4494,N_4423);
nor U4678 (N_4678,N_4414,N_4166);
xnor U4679 (N_4679,N_4340,N_4454);
or U4680 (N_4680,N_4078,N_4360);
and U4681 (N_4681,N_4084,N_4079);
and U4682 (N_4682,N_4133,N_4180);
and U4683 (N_4683,N_4246,N_4135);
nor U4684 (N_4684,N_4224,N_4484);
nor U4685 (N_4685,N_4351,N_4426);
nand U4686 (N_4686,N_4218,N_4158);
nand U4687 (N_4687,N_4125,N_4067);
xor U4688 (N_4688,N_4201,N_4043);
and U4689 (N_4689,N_4189,N_4037);
nand U4690 (N_4690,N_4489,N_4321);
and U4691 (N_4691,N_4382,N_4220);
or U4692 (N_4692,N_4171,N_4438);
and U4693 (N_4693,N_4452,N_4328);
and U4694 (N_4694,N_4402,N_4362);
xor U4695 (N_4695,N_4303,N_4295);
nand U4696 (N_4696,N_4089,N_4433);
nand U4697 (N_4697,N_4124,N_4424);
xor U4698 (N_4698,N_4155,N_4302);
or U4699 (N_4699,N_4336,N_4197);
nor U4700 (N_4700,N_4377,N_4074);
or U4701 (N_4701,N_4293,N_4437);
nand U4702 (N_4702,N_4049,N_4165);
xnor U4703 (N_4703,N_4215,N_4378);
nor U4704 (N_4704,N_4163,N_4110);
and U4705 (N_4705,N_4238,N_4205);
and U4706 (N_4706,N_4212,N_4326);
nor U4707 (N_4707,N_4210,N_4420);
xor U4708 (N_4708,N_4272,N_4469);
xnor U4709 (N_4709,N_4361,N_4369);
nor U4710 (N_4710,N_4299,N_4398);
nand U4711 (N_4711,N_4269,N_4383);
xor U4712 (N_4712,N_4076,N_4480);
or U4713 (N_4713,N_4122,N_4289);
xnor U4714 (N_4714,N_4267,N_4097);
nand U4715 (N_4715,N_4169,N_4055);
and U4716 (N_4716,N_4039,N_4397);
nor U4717 (N_4717,N_4234,N_4187);
xnor U4718 (N_4718,N_4287,N_4249);
and U4719 (N_4719,N_4275,N_4025);
xnor U4720 (N_4720,N_4200,N_4345);
nand U4721 (N_4721,N_4476,N_4153);
nand U4722 (N_4722,N_4463,N_4461);
nand U4723 (N_4723,N_4047,N_4455);
nor U4724 (N_4724,N_4258,N_4173);
or U4725 (N_4725,N_4213,N_4103);
xnor U4726 (N_4726,N_4170,N_4332);
and U4727 (N_4727,N_4301,N_4350);
or U4728 (N_4728,N_4286,N_4001);
nor U4729 (N_4729,N_4276,N_4120);
xnor U4730 (N_4730,N_4413,N_4242);
or U4731 (N_4731,N_4281,N_4046);
and U4732 (N_4732,N_4425,N_4020);
nor U4733 (N_4733,N_4384,N_4312);
xor U4734 (N_4734,N_4403,N_4203);
nand U4735 (N_4735,N_4140,N_4496);
or U4736 (N_4736,N_4314,N_4058);
nand U4737 (N_4737,N_4026,N_4388);
nor U4738 (N_4738,N_4366,N_4253);
xnor U4739 (N_4739,N_4335,N_4309);
nor U4740 (N_4740,N_4060,N_4445);
and U4741 (N_4741,N_4222,N_4236);
nand U4742 (N_4742,N_4112,N_4453);
or U4743 (N_4743,N_4386,N_4387);
xor U4744 (N_4744,N_4064,N_4256);
nor U4745 (N_4745,N_4444,N_4157);
nand U4746 (N_4746,N_4243,N_4030);
nand U4747 (N_4747,N_4316,N_4472);
nor U4748 (N_4748,N_4355,N_4399);
and U4749 (N_4749,N_4101,N_4022);
nand U4750 (N_4750,N_4021,N_4109);
xor U4751 (N_4751,N_4168,N_4245);
or U4752 (N_4752,N_4367,N_4052);
xnor U4753 (N_4753,N_4444,N_4488);
xor U4754 (N_4754,N_4027,N_4397);
nand U4755 (N_4755,N_4168,N_4008);
or U4756 (N_4756,N_4021,N_4261);
and U4757 (N_4757,N_4143,N_4454);
nand U4758 (N_4758,N_4096,N_4393);
nand U4759 (N_4759,N_4096,N_4366);
xor U4760 (N_4760,N_4151,N_4192);
nor U4761 (N_4761,N_4094,N_4001);
and U4762 (N_4762,N_4304,N_4251);
and U4763 (N_4763,N_4338,N_4334);
xnor U4764 (N_4764,N_4042,N_4494);
nand U4765 (N_4765,N_4168,N_4446);
or U4766 (N_4766,N_4201,N_4135);
nor U4767 (N_4767,N_4449,N_4139);
or U4768 (N_4768,N_4183,N_4190);
xnor U4769 (N_4769,N_4418,N_4282);
or U4770 (N_4770,N_4028,N_4349);
or U4771 (N_4771,N_4365,N_4495);
nand U4772 (N_4772,N_4154,N_4288);
nand U4773 (N_4773,N_4472,N_4095);
nand U4774 (N_4774,N_4277,N_4052);
and U4775 (N_4775,N_4110,N_4299);
and U4776 (N_4776,N_4369,N_4442);
or U4777 (N_4777,N_4188,N_4080);
and U4778 (N_4778,N_4312,N_4326);
nor U4779 (N_4779,N_4337,N_4215);
nor U4780 (N_4780,N_4224,N_4133);
and U4781 (N_4781,N_4131,N_4323);
and U4782 (N_4782,N_4423,N_4216);
or U4783 (N_4783,N_4291,N_4484);
nor U4784 (N_4784,N_4313,N_4343);
and U4785 (N_4785,N_4337,N_4321);
and U4786 (N_4786,N_4192,N_4300);
and U4787 (N_4787,N_4363,N_4339);
xor U4788 (N_4788,N_4443,N_4047);
and U4789 (N_4789,N_4235,N_4251);
nor U4790 (N_4790,N_4076,N_4164);
and U4791 (N_4791,N_4308,N_4107);
nor U4792 (N_4792,N_4432,N_4153);
nand U4793 (N_4793,N_4183,N_4006);
nor U4794 (N_4794,N_4145,N_4422);
nor U4795 (N_4795,N_4308,N_4151);
and U4796 (N_4796,N_4326,N_4338);
or U4797 (N_4797,N_4456,N_4462);
nor U4798 (N_4798,N_4142,N_4219);
and U4799 (N_4799,N_4176,N_4487);
nand U4800 (N_4800,N_4016,N_4275);
xnor U4801 (N_4801,N_4067,N_4249);
and U4802 (N_4802,N_4318,N_4435);
or U4803 (N_4803,N_4307,N_4421);
and U4804 (N_4804,N_4083,N_4058);
nor U4805 (N_4805,N_4428,N_4145);
or U4806 (N_4806,N_4267,N_4459);
nor U4807 (N_4807,N_4061,N_4228);
xor U4808 (N_4808,N_4084,N_4343);
or U4809 (N_4809,N_4396,N_4240);
nor U4810 (N_4810,N_4135,N_4086);
xnor U4811 (N_4811,N_4202,N_4303);
nand U4812 (N_4812,N_4395,N_4111);
nor U4813 (N_4813,N_4486,N_4303);
xor U4814 (N_4814,N_4406,N_4244);
or U4815 (N_4815,N_4179,N_4292);
nor U4816 (N_4816,N_4338,N_4362);
and U4817 (N_4817,N_4384,N_4316);
or U4818 (N_4818,N_4143,N_4323);
xnor U4819 (N_4819,N_4035,N_4226);
nand U4820 (N_4820,N_4342,N_4219);
nand U4821 (N_4821,N_4419,N_4346);
or U4822 (N_4822,N_4443,N_4218);
xnor U4823 (N_4823,N_4366,N_4377);
and U4824 (N_4824,N_4149,N_4331);
or U4825 (N_4825,N_4320,N_4284);
nand U4826 (N_4826,N_4147,N_4022);
xnor U4827 (N_4827,N_4294,N_4063);
or U4828 (N_4828,N_4196,N_4437);
and U4829 (N_4829,N_4066,N_4253);
and U4830 (N_4830,N_4269,N_4112);
and U4831 (N_4831,N_4044,N_4241);
nor U4832 (N_4832,N_4186,N_4352);
xnor U4833 (N_4833,N_4282,N_4381);
xor U4834 (N_4834,N_4489,N_4082);
xor U4835 (N_4835,N_4388,N_4335);
and U4836 (N_4836,N_4301,N_4211);
xnor U4837 (N_4837,N_4295,N_4260);
xnor U4838 (N_4838,N_4028,N_4388);
nand U4839 (N_4839,N_4246,N_4497);
and U4840 (N_4840,N_4078,N_4310);
nand U4841 (N_4841,N_4405,N_4138);
nor U4842 (N_4842,N_4397,N_4085);
nor U4843 (N_4843,N_4220,N_4210);
nand U4844 (N_4844,N_4307,N_4101);
and U4845 (N_4845,N_4450,N_4315);
nor U4846 (N_4846,N_4224,N_4138);
and U4847 (N_4847,N_4054,N_4330);
and U4848 (N_4848,N_4062,N_4259);
nor U4849 (N_4849,N_4213,N_4128);
nand U4850 (N_4850,N_4164,N_4043);
nand U4851 (N_4851,N_4405,N_4092);
nand U4852 (N_4852,N_4415,N_4328);
xnor U4853 (N_4853,N_4252,N_4250);
xor U4854 (N_4854,N_4225,N_4346);
nor U4855 (N_4855,N_4003,N_4030);
or U4856 (N_4856,N_4021,N_4404);
nor U4857 (N_4857,N_4011,N_4269);
nor U4858 (N_4858,N_4267,N_4039);
xor U4859 (N_4859,N_4045,N_4382);
and U4860 (N_4860,N_4249,N_4051);
or U4861 (N_4861,N_4182,N_4130);
or U4862 (N_4862,N_4234,N_4270);
xnor U4863 (N_4863,N_4185,N_4454);
nand U4864 (N_4864,N_4132,N_4136);
or U4865 (N_4865,N_4051,N_4321);
nand U4866 (N_4866,N_4373,N_4150);
or U4867 (N_4867,N_4437,N_4316);
or U4868 (N_4868,N_4170,N_4014);
nand U4869 (N_4869,N_4448,N_4313);
xor U4870 (N_4870,N_4372,N_4452);
xor U4871 (N_4871,N_4434,N_4025);
or U4872 (N_4872,N_4081,N_4490);
nor U4873 (N_4873,N_4143,N_4403);
xnor U4874 (N_4874,N_4285,N_4484);
nor U4875 (N_4875,N_4124,N_4073);
nand U4876 (N_4876,N_4367,N_4205);
nor U4877 (N_4877,N_4266,N_4318);
and U4878 (N_4878,N_4420,N_4193);
nand U4879 (N_4879,N_4262,N_4485);
or U4880 (N_4880,N_4459,N_4030);
and U4881 (N_4881,N_4159,N_4235);
nand U4882 (N_4882,N_4062,N_4098);
nor U4883 (N_4883,N_4325,N_4406);
nand U4884 (N_4884,N_4475,N_4160);
xor U4885 (N_4885,N_4169,N_4214);
or U4886 (N_4886,N_4311,N_4244);
nor U4887 (N_4887,N_4380,N_4155);
nand U4888 (N_4888,N_4350,N_4249);
nor U4889 (N_4889,N_4024,N_4350);
nor U4890 (N_4890,N_4078,N_4160);
or U4891 (N_4891,N_4459,N_4124);
nand U4892 (N_4892,N_4348,N_4175);
nand U4893 (N_4893,N_4298,N_4414);
nor U4894 (N_4894,N_4404,N_4448);
and U4895 (N_4895,N_4387,N_4457);
nand U4896 (N_4896,N_4189,N_4489);
nor U4897 (N_4897,N_4024,N_4081);
xnor U4898 (N_4898,N_4485,N_4148);
nor U4899 (N_4899,N_4255,N_4178);
or U4900 (N_4900,N_4386,N_4439);
xnor U4901 (N_4901,N_4430,N_4467);
or U4902 (N_4902,N_4122,N_4277);
nand U4903 (N_4903,N_4201,N_4143);
nor U4904 (N_4904,N_4118,N_4141);
nand U4905 (N_4905,N_4213,N_4111);
and U4906 (N_4906,N_4355,N_4105);
xnor U4907 (N_4907,N_4053,N_4069);
xnor U4908 (N_4908,N_4060,N_4350);
nor U4909 (N_4909,N_4156,N_4292);
nand U4910 (N_4910,N_4106,N_4446);
nor U4911 (N_4911,N_4461,N_4397);
nand U4912 (N_4912,N_4201,N_4480);
or U4913 (N_4913,N_4291,N_4244);
nor U4914 (N_4914,N_4242,N_4482);
nor U4915 (N_4915,N_4347,N_4033);
nor U4916 (N_4916,N_4347,N_4315);
and U4917 (N_4917,N_4086,N_4143);
nor U4918 (N_4918,N_4105,N_4104);
nor U4919 (N_4919,N_4283,N_4050);
and U4920 (N_4920,N_4018,N_4408);
nand U4921 (N_4921,N_4190,N_4300);
xnor U4922 (N_4922,N_4449,N_4380);
and U4923 (N_4923,N_4287,N_4173);
and U4924 (N_4924,N_4425,N_4114);
and U4925 (N_4925,N_4286,N_4248);
nand U4926 (N_4926,N_4090,N_4348);
and U4927 (N_4927,N_4449,N_4280);
or U4928 (N_4928,N_4347,N_4195);
nor U4929 (N_4929,N_4261,N_4257);
xnor U4930 (N_4930,N_4301,N_4170);
nand U4931 (N_4931,N_4384,N_4081);
xor U4932 (N_4932,N_4229,N_4219);
nor U4933 (N_4933,N_4332,N_4452);
nor U4934 (N_4934,N_4298,N_4253);
nand U4935 (N_4935,N_4404,N_4060);
xor U4936 (N_4936,N_4166,N_4352);
nand U4937 (N_4937,N_4339,N_4193);
or U4938 (N_4938,N_4206,N_4236);
nor U4939 (N_4939,N_4149,N_4167);
or U4940 (N_4940,N_4156,N_4432);
and U4941 (N_4941,N_4208,N_4276);
and U4942 (N_4942,N_4179,N_4005);
or U4943 (N_4943,N_4270,N_4474);
xor U4944 (N_4944,N_4331,N_4221);
xnor U4945 (N_4945,N_4329,N_4385);
xor U4946 (N_4946,N_4162,N_4121);
xnor U4947 (N_4947,N_4372,N_4130);
nand U4948 (N_4948,N_4309,N_4122);
xor U4949 (N_4949,N_4355,N_4461);
and U4950 (N_4950,N_4072,N_4294);
nor U4951 (N_4951,N_4050,N_4126);
nor U4952 (N_4952,N_4061,N_4264);
nor U4953 (N_4953,N_4192,N_4150);
xnor U4954 (N_4954,N_4173,N_4319);
and U4955 (N_4955,N_4045,N_4039);
nand U4956 (N_4956,N_4305,N_4470);
xor U4957 (N_4957,N_4298,N_4460);
and U4958 (N_4958,N_4437,N_4330);
xor U4959 (N_4959,N_4003,N_4403);
nor U4960 (N_4960,N_4227,N_4064);
xor U4961 (N_4961,N_4191,N_4132);
and U4962 (N_4962,N_4215,N_4356);
nand U4963 (N_4963,N_4113,N_4323);
xnor U4964 (N_4964,N_4300,N_4261);
or U4965 (N_4965,N_4384,N_4206);
nand U4966 (N_4966,N_4315,N_4433);
nor U4967 (N_4967,N_4456,N_4195);
nor U4968 (N_4968,N_4198,N_4118);
xor U4969 (N_4969,N_4364,N_4124);
xnor U4970 (N_4970,N_4249,N_4489);
or U4971 (N_4971,N_4362,N_4363);
or U4972 (N_4972,N_4109,N_4080);
nand U4973 (N_4973,N_4407,N_4473);
xnor U4974 (N_4974,N_4494,N_4145);
or U4975 (N_4975,N_4452,N_4459);
and U4976 (N_4976,N_4048,N_4243);
nand U4977 (N_4977,N_4204,N_4205);
nand U4978 (N_4978,N_4138,N_4468);
and U4979 (N_4979,N_4033,N_4466);
xor U4980 (N_4980,N_4070,N_4415);
nor U4981 (N_4981,N_4289,N_4450);
and U4982 (N_4982,N_4071,N_4377);
and U4983 (N_4983,N_4454,N_4261);
or U4984 (N_4984,N_4335,N_4434);
or U4985 (N_4985,N_4242,N_4338);
and U4986 (N_4986,N_4096,N_4156);
nand U4987 (N_4987,N_4077,N_4253);
xnor U4988 (N_4988,N_4269,N_4473);
xor U4989 (N_4989,N_4066,N_4495);
nor U4990 (N_4990,N_4084,N_4096);
and U4991 (N_4991,N_4460,N_4413);
and U4992 (N_4992,N_4397,N_4373);
nor U4993 (N_4993,N_4406,N_4019);
nor U4994 (N_4994,N_4450,N_4236);
and U4995 (N_4995,N_4339,N_4419);
nor U4996 (N_4996,N_4444,N_4183);
or U4997 (N_4997,N_4118,N_4214);
nand U4998 (N_4998,N_4323,N_4292);
or U4999 (N_4999,N_4263,N_4470);
and U5000 (N_5000,N_4734,N_4837);
or U5001 (N_5001,N_4834,N_4771);
nor U5002 (N_5002,N_4515,N_4849);
or U5003 (N_5003,N_4839,N_4598);
or U5004 (N_5004,N_4966,N_4503);
xnor U5005 (N_5005,N_4955,N_4833);
or U5006 (N_5006,N_4567,N_4888);
or U5007 (N_5007,N_4563,N_4787);
nand U5008 (N_5008,N_4733,N_4809);
and U5009 (N_5009,N_4573,N_4516);
and U5010 (N_5010,N_4933,N_4585);
and U5011 (N_5011,N_4813,N_4824);
and U5012 (N_5012,N_4612,N_4583);
nand U5013 (N_5013,N_4520,N_4924);
nor U5014 (N_5014,N_4670,N_4804);
and U5015 (N_5015,N_4614,N_4697);
xnor U5016 (N_5016,N_4679,N_4694);
xor U5017 (N_5017,N_4609,N_4658);
or U5018 (N_5018,N_4711,N_4810);
nand U5019 (N_5019,N_4847,N_4958);
nor U5020 (N_5020,N_4564,N_4832);
nand U5021 (N_5021,N_4659,N_4501);
nor U5022 (N_5022,N_4651,N_4584);
nor U5023 (N_5023,N_4867,N_4635);
or U5024 (N_5024,N_4764,N_4953);
nand U5025 (N_5025,N_4677,N_4606);
xor U5026 (N_5026,N_4945,N_4518);
xor U5027 (N_5027,N_4591,N_4696);
or U5028 (N_5028,N_4829,N_4715);
or U5029 (N_5029,N_4812,N_4806);
nand U5030 (N_5030,N_4758,N_4765);
nor U5031 (N_5031,N_4714,N_4979);
xnor U5032 (N_5032,N_4961,N_4856);
and U5033 (N_5033,N_4808,N_4992);
and U5034 (N_5034,N_4912,N_4907);
nand U5035 (N_5035,N_4899,N_4700);
nor U5036 (N_5036,N_4865,N_4802);
or U5037 (N_5037,N_4741,N_4746);
and U5038 (N_5038,N_4773,N_4624);
or U5039 (N_5039,N_4820,N_4920);
xnor U5040 (N_5040,N_4536,N_4836);
or U5041 (N_5041,N_4822,N_4892);
nand U5042 (N_5042,N_4960,N_4608);
or U5043 (N_5043,N_4754,N_4618);
xnor U5044 (N_5044,N_4919,N_4649);
xor U5045 (N_5045,N_4556,N_4547);
nand U5046 (N_5046,N_4653,N_4638);
nand U5047 (N_5047,N_4791,N_4757);
nand U5048 (N_5048,N_4623,N_4702);
xor U5049 (N_5049,N_4819,N_4514);
or U5050 (N_5050,N_4718,N_4610);
nand U5051 (N_5051,N_4657,N_4941);
xor U5052 (N_5052,N_4875,N_4852);
xor U5053 (N_5053,N_4579,N_4590);
nor U5054 (N_5054,N_4772,N_4934);
xnor U5055 (N_5055,N_4687,N_4664);
nor U5056 (N_5056,N_4965,N_4707);
nand U5057 (N_5057,N_4735,N_4523);
nand U5058 (N_5058,N_4753,N_4871);
and U5059 (N_5059,N_4723,N_4937);
and U5060 (N_5060,N_4826,N_4835);
and U5061 (N_5061,N_4554,N_4908);
or U5062 (N_5062,N_4825,N_4983);
and U5063 (N_5063,N_4790,N_4628);
or U5064 (N_5064,N_4990,N_4751);
or U5065 (N_5065,N_4781,N_4971);
nor U5066 (N_5066,N_4626,N_4925);
nand U5067 (N_5067,N_4748,N_4782);
xnor U5068 (N_5068,N_4668,N_4534);
nand U5069 (N_5069,N_4922,N_4502);
nand U5070 (N_5070,N_4926,N_4568);
xor U5071 (N_5071,N_4543,N_4974);
nand U5072 (N_5072,N_4749,N_4581);
nand U5073 (N_5073,N_4768,N_4863);
nand U5074 (N_5074,N_4505,N_4603);
and U5075 (N_5075,N_4617,N_4840);
or U5076 (N_5076,N_4654,N_4666);
and U5077 (N_5077,N_4551,N_4507);
nand U5078 (N_5078,N_4594,N_4905);
and U5079 (N_5079,N_4743,N_4732);
xor U5080 (N_5080,N_4795,N_4548);
xor U5081 (N_5081,N_4967,N_4959);
xnor U5082 (N_5082,N_4785,N_4690);
xor U5083 (N_5083,N_4762,N_4900);
and U5084 (N_5084,N_4616,N_4942);
and U5085 (N_5085,N_4607,N_4513);
nor U5086 (N_5086,N_4755,N_4823);
and U5087 (N_5087,N_4525,N_4986);
or U5088 (N_5088,N_4977,N_4948);
and U5089 (N_5089,N_4589,N_4910);
and U5090 (N_5090,N_4917,N_4797);
xnor U5091 (N_5091,N_4662,N_4636);
xor U5092 (N_5092,N_4683,N_4987);
xnor U5093 (N_5093,N_4864,N_4645);
and U5094 (N_5094,N_4538,N_4691);
nor U5095 (N_5095,N_4783,N_4774);
xnor U5096 (N_5096,N_4582,N_4970);
nor U5097 (N_5097,N_4519,N_4600);
or U5098 (N_5098,N_4704,N_4995);
nor U5099 (N_5099,N_4828,N_4855);
xnor U5100 (N_5100,N_4510,N_4681);
nand U5101 (N_5101,N_4593,N_4529);
nand U5102 (N_5102,N_4602,N_4909);
nand U5103 (N_5103,N_4973,N_4817);
or U5104 (N_5104,N_4742,N_4642);
or U5105 (N_5105,N_4876,N_4509);
nand U5106 (N_5106,N_4578,N_4553);
nor U5107 (N_5107,N_4760,N_4844);
nand U5108 (N_5108,N_4857,N_4798);
nand U5109 (N_5109,N_4946,N_4560);
nor U5110 (N_5110,N_4730,N_4969);
xor U5111 (N_5111,N_4821,N_4650);
or U5112 (N_5112,N_4587,N_4663);
xor U5113 (N_5113,N_4994,N_4897);
xor U5114 (N_5114,N_4964,N_4939);
nor U5115 (N_5115,N_4752,N_4851);
nand U5116 (N_5116,N_4570,N_4859);
nor U5117 (N_5117,N_4877,N_4678);
nor U5118 (N_5118,N_4588,N_4893);
xnor U5119 (N_5119,N_4688,N_4592);
nand U5120 (N_5120,N_4577,N_4745);
xnor U5121 (N_5121,N_4984,N_4631);
and U5122 (N_5122,N_4540,N_4800);
or U5123 (N_5123,N_4862,N_4550);
or U5124 (N_5124,N_4775,N_4527);
or U5125 (N_5125,N_4763,N_4901);
xor U5126 (N_5126,N_4956,N_4738);
and U5127 (N_5127,N_4896,N_4853);
nor U5128 (N_5128,N_4722,N_4918);
xor U5129 (N_5129,N_4838,N_4861);
nand U5130 (N_5130,N_4555,N_4508);
and U5131 (N_5131,N_4906,N_4655);
nor U5132 (N_5132,N_4619,N_4938);
xor U5133 (N_5133,N_4803,N_4737);
nand U5134 (N_5134,N_4770,N_4921);
nor U5135 (N_5135,N_4744,N_4575);
or U5136 (N_5136,N_4846,N_4894);
nand U5137 (N_5137,N_4880,N_4843);
or U5138 (N_5138,N_4978,N_4815);
nand U5139 (N_5139,N_4890,N_4727);
or U5140 (N_5140,N_4981,N_4996);
or U5141 (N_5141,N_4597,N_4885);
or U5142 (N_5142,N_4706,N_4565);
nand U5143 (N_5143,N_4728,N_4627);
xnor U5144 (N_5144,N_4557,N_4930);
nor U5145 (N_5145,N_4976,N_4621);
nor U5146 (N_5146,N_4870,N_4613);
and U5147 (N_5147,N_4850,N_4661);
xor U5148 (N_5148,N_4675,N_4710);
xnor U5149 (N_5149,N_4652,N_4673);
nand U5150 (N_5150,N_4685,N_4689);
or U5151 (N_5151,N_4858,N_4506);
and U5152 (N_5152,N_4927,N_4957);
xor U5153 (N_5153,N_4667,N_4720);
nor U5154 (N_5154,N_4972,N_4993);
nor U5155 (N_5155,N_4801,N_4580);
xor U5156 (N_5156,N_4895,N_4647);
nand U5157 (N_5157,N_4717,N_4999);
or U5158 (N_5158,N_4705,N_4698);
and U5159 (N_5159,N_4914,N_4660);
or U5160 (N_5160,N_4676,N_4947);
nand U5161 (N_5161,N_4796,N_4991);
or U5162 (N_5162,N_4701,N_4827);
xnor U5163 (N_5163,N_4854,N_4805);
xnor U5164 (N_5164,N_4786,N_4750);
nor U5165 (N_5165,N_4630,N_4528);
nor U5166 (N_5166,N_4686,N_4656);
nand U5167 (N_5167,N_4868,N_4788);
xnor U5168 (N_5168,N_4566,N_4767);
and U5169 (N_5169,N_4541,N_4530);
xor U5170 (N_5170,N_4904,N_4869);
or U5171 (N_5171,N_4872,N_4879);
xor U5172 (N_5172,N_4747,N_4963);
or U5173 (N_5173,N_4719,N_4646);
or U5174 (N_5174,N_4873,N_4574);
nor U5175 (N_5175,N_4916,N_4708);
or U5176 (N_5176,N_4545,N_4776);
nand U5177 (N_5177,N_4860,N_4692);
nand U5178 (N_5178,N_4640,N_4985);
xor U5179 (N_5179,N_4671,N_4703);
nand U5180 (N_5180,N_4915,N_4932);
xor U5181 (N_5181,N_4622,N_4968);
nand U5182 (N_5182,N_4569,N_4726);
nor U5183 (N_5183,N_4562,N_4998);
and U5184 (N_5184,N_4644,N_4881);
or U5185 (N_5185,N_4611,N_4542);
or U5186 (N_5186,N_4940,N_4944);
and U5187 (N_5187,N_4595,N_4980);
nor U5188 (N_5188,N_4639,N_4891);
or U5189 (N_5189,N_4533,N_4665);
or U5190 (N_5190,N_4951,N_4586);
xor U5191 (N_5191,N_4522,N_4601);
or U5192 (N_5192,N_4884,N_4779);
xor U5193 (N_5193,N_4643,N_4521);
nor U5194 (N_5194,N_4558,N_4845);
and U5195 (N_5195,N_4721,N_4988);
xor U5196 (N_5196,N_4641,N_4814);
or U5197 (N_5197,N_4713,N_4633);
or U5198 (N_5198,N_4949,N_4634);
or U5199 (N_5199,N_4923,N_4830);
and U5200 (N_5200,N_4954,N_4841);
nor U5201 (N_5201,N_4807,N_4682);
and U5202 (N_5202,N_4778,N_4929);
and U5203 (N_5203,N_4928,N_4725);
and U5204 (N_5204,N_4848,N_4599);
or U5205 (N_5205,N_4878,N_4784);
nor U5206 (N_5206,N_4935,N_4889);
and U5207 (N_5207,N_4769,N_4911);
and U5208 (N_5208,N_4531,N_4780);
nor U5209 (N_5209,N_4517,N_4792);
xnor U5210 (N_5210,N_4739,N_4874);
or U5211 (N_5211,N_4962,N_4716);
and U5212 (N_5212,N_4695,N_4684);
nor U5213 (N_5213,N_4680,N_4842);
nand U5214 (N_5214,N_4931,N_4799);
xnor U5215 (N_5215,N_4982,N_4546);
and U5216 (N_5216,N_4759,N_4552);
nor U5217 (N_5217,N_4561,N_4625);
or U5218 (N_5218,N_4572,N_4898);
and U5219 (N_5219,N_4637,N_4789);
nand U5220 (N_5220,N_4604,N_4724);
and U5221 (N_5221,N_4535,N_4740);
nand U5222 (N_5222,N_4756,N_4512);
or U5223 (N_5223,N_4632,N_4989);
nand U5224 (N_5224,N_4620,N_4615);
nor U5225 (N_5225,N_4544,N_4709);
nand U5226 (N_5226,N_4866,N_4712);
nand U5227 (N_5227,N_4936,N_4672);
or U5228 (N_5228,N_4605,N_4975);
and U5229 (N_5229,N_4818,N_4913);
xor U5230 (N_5230,N_4537,N_4576);
nor U5231 (N_5231,N_4793,N_4596);
nor U5232 (N_5232,N_4729,N_4549);
nand U5233 (N_5233,N_4903,N_4539);
xnor U5234 (N_5234,N_4950,N_4766);
nand U5235 (N_5235,N_4731,N_4674);
or U5236 (N_5236,N_4997,N_4831);
nand U5237 (N_5237,N_4669,N_4811);
nand U5238 (N_5238,N_4882,N_4500);
or U5239 (N_5239,N_4526,N_4886);
nor U5240 (N_5240,N_4511,N_4943);
or U5241 (N_5241,N_4777,N_4524);
nand U5242 (N_5242,N_4504,N_4699);
nand U5243 (N_5243,N_4887,N_4629);
nand U5244 (N_5244,N_4736,N_4794);
or U5245 (N_5245,N_4559,N_4532);
nand U5246 (N_5246,N_4648,N_4761);
and U5247 (N_5247,N_4952,N_4571);
nand U5248 (N_5248,N_4693,N_4816);
or U5249 (N_5249,N_4883,N_4902);
nor U5250 (N_5250,N_4569,N_4686);
nor U5251 (N_5251,N_4986,N_4556);
and U5252 (N_5252,N_4708,N_4943);
and U5253 (N_5253,N_4965,N_4577);
or U5254 (N_5254,N_4516,N_4873);
nor U5255 (N_5255,N_4673,N_4991);
nand U5256 (N_5256,N_4871,N_4756);
nand U5257 (N_5257,N_4961,N_4520);
xor U5258 (N_5258,N_4662,N_4690);
xnor U5259 (N_5259,N_4533,N_4739);
nor U5260 (N_5260,N_4850,N_4915);
nor U5261 (N_5261,N_4982,N_4622);
nand U5262 (N_5262,N_4555,N_4547);
and U5263 (N_5263,N_4689,N_4934);
or U5264 (N_5264,N_4935,N_4552);
xnor U5265 (N_5265,N_4793,N_4659);
xor U5266 (N_5266,N_4713,N_4980);
and U5267 (N_5267,N_4581,N_4663);
and U5268 (N_5268,N_4594,N_4526);
xnor U5269 (N_5269,N_4657,N_4790);
or U5270 (N_5270,N_4627,N_4993);
and U5271 (N_5271,N_4629,N_4527);
or U5272 (N_5272,N_4804,N_4904);
or U5273 (N_5273,N_4554,N_4637);
nand U5274 (N_5274,N_4604,N_4799);
nor U5275 (N_5275,N_4630,N_4636);
nor U5276 (N_5276,N_4959,N_4540);
and U5277 (N_5277,N_4512,N_4575);
or U5278 (N_5278,N_4563,N_4553);
and U5279 (N_5279,N_4936,N_4985);
or U5280 (N_5280,N_4922,N_4862);
nor U5281 (N_5281,N_4715,N_4555);
xor U5282 (N_5282,N_4799,N_4764);
and U5283 (N_5283,N_4917,N_4908);
nor U5284 (N_5284,N_4728,N_4639);
or U5285 (N_5285,N_4859,N_4560);
and U5286 (N_5286,N_4660,N_4829);
nor U5287 (N_5287,N_4955,N_4569);
xnor U5288 (N_5288,N_4718,N_4525);
or U5289 (N_5289,N_4773,N_4651);
xor U5290 (N_5290,N_4836,N_4642);
nor U5291 (N_5291,N_4874,N_4651);
and U5292 (N_5292,N_4997,N_4779);
xor U5293 (N_5293,N_4721,N_4706);
xor U5294 (N_5294,N_4668,N_4576);
xor U5295 (N_5295,N_4958,N_4742);
xnor U5296 (N_5296,N_4924,N_4517);
xnor U5297 (N_5297,N_4563,N_4548);
nand U5298 (N_5298,N_4587,N_4628);
nand U5299 (N_5299,N_4812,N_4887);
xor U5300 (N_5300,N_4623,N_4862);
nor U5301 (N_5301,N_4859,N_4905);
and U5302 (N_5302,N_4540,N_4920);
xor U5303 (N_5303,N_4515,N_4531);
xor U5304 (N_5304,N_4956,N_4576);
or U5305 (N_5305,N_4586,N_4881);
nor U5306 (N_5306,N_4546,N_4511);
and U5307 (N_5307,N_4603,N_4758);
xnor U5308 (N_5308,N_4858,N_4924);
nor U5309 (N_5309,N_4733,N_4739);
nor U5310 (N_5310,N_4542,N_4661);
nor U5311 (N_5311,N_4585,N_4506);
nor U5312 (N_5312,N_4668,N_4501);
or U5313 (N_5313,N_4814,N_4539);
nor U5314 (N_5314,N_4955,N_4651);
and U5315 (N_5315,N_4927,N_4605);
xor U5316 (N_5316,N_4558,N_4589);
xor U5317 (N_5317,N_4977,N_4767);
xor U5318 (N_5318,N_4920,N_4876);
and U5319 (N_5319,N_4778,N_4931);
nand U5320 (N_5320,N_4515,N_4941);
and U5321 (N_5321,N_4892,N_4871);
nor U5322 (N_5322,N_4781,N_4871);
xor U5323 (N_5323,N_4813,N_4875);
nand U5324 (N_5324,N_4831,N_4739);
nor U5325 (N_5325,N_4645,N_4856);
nand U5326 (N_5326,N_4824,N_4791);
nor U5327 (N_5327,N_4583,N_4806);
nand U5328 (N_5328,N_4633,N_4810);
or U5329 (N_5329,N_4561,N_4857);
or U5330 (N_5330,N_4618,N_4744);
xnor U5331 (N_5331,N_4710,N_4701);
and U5332 (N_5332,N_4863,N_4526);
nand U5333 (N_5333,N_4706,N_4975);
nand U5334 (N_5334,N_4613,N_4924);
or U5335 (N_5335,N_4951,N_4991);
or U5336 (N_5336,N_4642,N_4822);
nand U5337 (N_5337,N_4580,N_4976);
and U5338 (N_5338,N_4914,N_4840);
nand U5339 (N_5339,N_4609,N_4757);
xnor U5340 (N_5340,N_4980,N_4749);
and U5341 (N_5341,N_4759,N_4800);
or U5342 (N_5342,N_4539,N_4532);
and U5343 (N_5343,N_4698,N_4887);
nand U5344 (N_5344,N_4944,N_4550);
and U5345 (N_5345,N_4895,N_4701);
nand U5346 (N_5346,N_4712,N_4626);
nand U5347 (N_5347,N_4583,N_4776);
or U5348 (N_5348,N_4904,N_4534);
nand U5349 (N_5349,N_4569,N_4801);
xnor U5350 (N_5350,N_4834,N_4920);
nand U5351 (N_5351,N_4954,N_4859);
and U5352 (N_5352,N_4534,N_4531);
and U5353 (N_5353,N_4505,N_4886);
and U5354 (N_5354,N_4845,N_4563);
nor U5355 (N_5355,N_4767,N_4743);
nor U5356 (N_5356,N_4974,N_4522);
xor U5357 (N_5357,N_4750,N_4830);
nor U5358 (N_5358,N_4742,N_4796);
or U5359 (N_5359,N_4892,N_4786);
or U5360 (N_5360,N_4747,N_4675);
and U5361 (N_5361,N_4648,N_4994);
and U5362 (N_5362,N_4989,N_4616);
xor U5363 (N_5363,N_4919,N_4594);
or U5364 (N_5364,N_4621,N_4831);
and U5365 (N_5365,N_4683,N_4655);
or U5366 (N_5366,N_4991,N_4905);
nand U5367 (N_5367,N_4500,N_4614);
and U5368 (N_5368,N_4778,N_4926);
or U5369 (N_5369,N_4842,N_4957);
and U5370 (N_5370,N_4677,N_4910);
and U5371 (N_5371,N_4789,N_4707);
nor U5372 (N_5372,N_4686,N_4659);
xor U5373 (N_5373,N_4712,N_4538);
nand U5374 (N_5374,N_4878,N_4597);
nand U5375 (N_5375,N_4560,N_4759);
xnor U5376 (N_5376,N_4552,N_4914);
and U5377 (N_5377,N_4964,N_4518);
nor U5378 (N_5378,N_4594,N_4901);
and U5379 (N_5379,N_4553,N_4689);
and U5380 (N_5380,N_4640,N_4801);
and U5381 (N_5381,N_4616,N_4954);
or U5382 (N_5382,N_4527,N_4599);
nand U5383 (N_5383,N_4522,N_4813);
nor U5384 (N_5384,N_4685,N_4656);
nand U5385 (N_5385,N_4539,N_4634);
nor U5386 (N_5386,N_4552,N_4761);
and U5387 (N_5387,N_4919,N_4868);
xor U5388 (N_5388,N_4937,N_4734);
nand U5389 (N_5389,N_4765,N_4979);
nor U5390 (N_5390,N_4892,N_4561);
nor U5391 (N_5391,N_4751,N_4596);
nor U5392 (N_5392,N_4779,N_4840);
and U5393 (N_5393,N_4532,N_4926);
nor U5394 (N_5394,N_4649,N_4535);
and U5395 (N_5395,N_4765,N_4587);
nor U5396 (N_5396,N_4757,N_4567);
or U5397 (N_5397,N_4638,N_4862);
or U5398 (N_5398,N_4902,N_4728);
or U5399 (N_5399,N_4553,N_4951);
and U5400 (N_5400,N_4967,N_4935);
xnor U5401 (N_5401,N_4806,N_4536);
nor U5402 (N_5402,N_4700,N_4998);
xnor U5403 (N_5403,N_4880,N_4972);
and U5404 (N_5404,N_4558,N_4507);
nor U5405 (N_5405,N_4945,N_4998);
and U5406 (N_5406,N_4521,N_4679);
xnor U5407 (N_5407,N_4933,N_4845);
or U5408 (N_5408,N_4617,N_4505);
nor U5409 (N_5409,N_4842,N_4997);
nor U5410 (N_5410,N_4631,N_4991);
nor U5411 (N_5411,N_4963,N_4535);
nor U5412 (N_5412,N_4759,N_4584);
and U5413 (N_5413,N_4768,N_4873);
or U5414 (N_5414,N_4674,N_4810);
and U5415 (N_5415,N_4583,N_4574);
xnor U5416 (N_5416,N_4642,N_4967);
or U5417 (N_5417,N_4698,N_4613);
xor U5418 (N_5418,N_4716,N_4624);
xnor U5419 (N_5419,N_4750,N_4797);
nand U5420 (N_5420,N_4579,N_4629);
and U5421 (N_5421,N_4636,N_4784);
or U5422 (N_5422,N_4876,N_4588);
xor U5423 (N_5423,N_4951,N_4817);
nand U5424 (N_5424,N_4801,N_4513);
or U5425 (N_5425,N_4883,N_4922);
xnor U5426 (N_5426,N_4698,N_4957);
xor U5427 (N_5427,N_4726,N_4882);
and U5428 (N_5428,N_4851,N_4946);
xor U5429 (N_5429,N_4534,N_4648);
nor U5430 (N_5430,N_4947,N_4960);
nor U5431 (N_5431,N_4665,N_4964);
and U5432 (N_5432,N_4654,N_4906);
nand U5433 (N_5433,N_4971,N_4654);
or U5434 (N_5434,N_4953,N_4624);
xor U5435 (N_5435,N_4694,N_4631);
nand U5436 (N_5436,N_4716,N_4640);
or U5437 (N_5437,N_4734,N_4731);
and U5438 (N_5438,N_4721,N_4519);
and U5439 (N_5439,N_4578,N_4970);
xor U5440 (N_5440,N_4680,N_4631);
or U5441 (N_5441,N_4763,N_4993);
xor U5442 (N_5442,N_4745,N_4736);
or U5443 (N_5443,N_4560,N_4732);
nand U5444 (N_5444,N_4506,N_4885);
or U5445 (N_5445,N_4657,N_4802);
nor U5446 (N_5446,N_4816,N_4905);
xor U5447 (N_5447,N_4934,N_4739);
nand U5448 (N_5448,N_4579,N_4994);
nand U5449 (N_5449,N_4507,N_4916);
xor U5450 (N_5450,N_4701,N_4761);
and U5451 (N_5451,N_4852,N_4501);
nor U5452 (N_5452,N_4863,N_4990);
or U5453 (N_5453,N_4532,N_4816);
or U5454 (N_5454,N_4715,N_4898);
or U5455 (N_5455,N_4546,N_4813);
nand U5456 (N_5456,N_4714,N_4601);
nor U5457 (N_5457,N_4874,N_4941);
nand U5458 (N_5458,N_4947,N_4830);
and U5459 (N_5459,N_4578,N_4936);
or U5460 (N_5460,N_4976,N_4688);
nand U5461 (N_5461,N_4628,N_4599);
or U5462 (N_5462,N_4637,N_4565);
nand U5463 (N_5463,N_4648,N_4877);
xor U5464 (N_5464,N_4852,N_4966);
or U5465 (N_5465,N_4943,N_4716);
and U5466 (N_5466,N_4744,N_4647);
and U5467 (N_5467,N_4905,N_4501);
nand U5468 (N_5468,N_4946,N_4732);
xor U5469 (N_5469,N_4727,N_4899);
and U5470 (N_5470,N_4649,N_4652);
and U5471 (N_5471,N_4672,N_4816);
and U5472 (N_5472,N_4727,N_4733);
xnor U5473 (N_5473,N_4690,N_4601);
or U5474 (N_5474,N_4868,N_4805);
nand U5475 (N_5475,N_4763,N_4749);
nor U5476 (N_5476,N_4622,N_4838);
xnor U5477 (N_5477,N_4999,N_4801);
nand U5478 (N_5478,N_4735,N_4716);
or U5479 (N_5479,N_4715,N_4824);
xor U5480 (N_5480,N_4562,N_4544);
nand U5481 (N_5481,N_4989,N_4927);
or U5482 (N_5482,N_4815,N_4596);
xnor U5483 (N_5483,N_4736,N_4983);
or U5484 (N_5484,N_4596,N_4953);
and U5485 (N_5485,N_4634,N_4759);
nand U5486 (N_5486,N_4842,N_4786);
or U5487 (N_5487,N_4636,N_4752);
nor U5488 (N_5488,N_4658,N_4940);
nand U5489 (N_5489,N_4734,N_4582);
nor U5490 (N_5490,N_4871,N_4976);
nand U5491 (N_5491,N_4983,N_4832);
nor U5492 (N_5492,N_4831,N_4678);
nand U5493 (N_5493,N_4848,N_4513);
xor U5494 (N_5494,N_4770,N_4633);
and U5495 (N_5495,N_4973,N_4781);
xnor U5496 (N_5496,N_4648,N_4673);
or U5497 (N_5497,N_4778,N_4588);
xor U5498 (N_5498,N_4522,N_4833);
and U5499 (N_5499,N_4895,N_4616);
or U5500 (N_5500,N_5042,N_5199);
xor U5501 (N_5501,N_5033,N_5023);
or U5502 (N_5502,N_5489,N_5085);
nand U5503 (N_5503,N_5149,N_5152);
nor U5504 (N_5504,N_5467,N_5338);
nor U5505 (N_5505,N_5260,N_5286);
xnor U5506 (N_5506,N_5353,N_5406);
xor U5507 (N_5507,N_5375,N_5093);
and U5508 (N_5508,N_5277,N_5056);
nor U5509 (N_5509,N_5430,N_5455);
nor U5510 (N_5510,N_5411,N_5378);
nand U5511 (N_5511,N_5090,N_5217);
nor U5512 (N_5512,N_5204,N_5313);
nor U5513 (N_5513,N_5321,N_5150);
xor U5514 (N_5514,N_5257,N_5194);
or U5515 (N_5515,N_5483,N_5423);
nor U5516 (N_5516,N_5103,N_5154);
and U5517 (N_5517,N_5071,N_5229);
nor U5518 (N_5518,N_5188,N_5376);
nor U5519 (N_5519,N_5118,N_5458);
xor U5520 (N_5520,N_5379,N_5230);
xor U5521 (N_5521,N_5235,N_5187);
or U5522 (N_5522,N_5245,N_5363);
nor U5523 (N_5523,N_5221,N_5362);
and U5524 (N_5524,N_5479,N_5039);
nand U5525 (N_5525,N_5298,N_5404);
and U5526 (N_5526,N_5481,N_5002);
xnor U5527 (N_5527,N_5328,N_5111);
and U5528 (N_5528,N_5198,N_5314);
and U5529 (N_5529,N_5330,N_5102);
and U5530 (N_5530,N_5143,N_5053);
and U5531 (N_5531,N_5128,N_5388);
and U5532 (N_5532,N_5193,N_5228);
and U5533 (N_5533,N_5209,N_5317);
xnor U5534 (N_5534,N_5097,N_5393);
nand U5535 (N_5535,N_5383,N_5334);
xnor U5536 (N_5536,N_5066,N_5357);
and U5537 (N_5537,N_5164,N_5469);
or U5538 (N_5538,N_5280,N_5231);
nand U5539 (N_5539,N_5471,N_5410);
nor U5540 (N_5540,N_5211,N_5468);
and U5541 (N_5541,N_5202,N_5282);
or U5542 (N_5542,N_5425,N_5315);
nand U5543 (N_5543,N_5266,N_5225);
xor U5544 (N_5544,N_5178,N_5269);
xor U5545 (N_5545,N_5465,N_5121);
and U5546 (N_5546,N_5360,N_5349);
nor U5547 (N_5547,N_5488,N_5215);
nand U5548 (N_5548,N_5496,N_5310);
or U5549 (N_5549,N_5044,N_5001);
xnor U5550 (N_5550,N_5431,N_5241);
nor U5551 (N_5551,N_5180,N_5438);
xor U5552 (N_5552,N_5446,N_5141);
nor U5553 (N_5553,N_5451,N_5478);
or U5554 (N_5554,N_5356,N_5276);
nand U5555 (N_5555,N_5059,N_5181);
or U5556 (N_5556,N_5304,N_5084);
xnor U5557 (N_5557,N_5226,N_5041);
or U5558 (N_5558,N_5473,N_5160);
or U5559 (N_5559,N_5470,N_5380);
or U5560 (N_5560,N_5476,N_5403);
xnor U5561 (N_5561,N_5250,N_5437);
and U5562 (N_5562,N_5267,N_5371);
xnor U5563 (N_5563,N_5030,N_5146);
or U5564 (N_5564,N_5435,N_5457);
nor U5565 (N_5565,N_5132,N_5122);
nand U5566 (N_5566,N_5147,N_5119);
or U5567 (N_5567,N_5350,N_5192);
nand U5568 (N_5568,N_5368,N_5013);
and U5569 (N_5569,N_5072,N_5480);
nor U5570 (N_5570,N_5037,N_5016);
nand U5571 (N_5571,N_5113,N_5264);
and U5572 (N_5572,N_5070,N_5238);
and U5573 (N_5573,N_5005,N_5292);
nor U5574 (N_5574,N_5336,N_5249);
nor U5575 (N_5575,N_5498,N_5104);
nor U5576 (N_5576,N_5026,N_5110);
nor U5577 (N_5577,N_5061,N_5274);
or U5578 (N_5578,N_5244,N_5397);
and U5579 (N_5579,N_5012,N_5327);
xnor U5580 (N_5580,N_5445,N_5220);
and U5581 (N_5581,N_5253,N_5015);
or U5582 (N_5582,N_5216,N_5067);
nand U5583 (N_5583,N_5144,N_5354);
or U5584 (N_5584,N_5052,N_5407);
nor U5585 (N_5585,N_5265,N_5167);
or U5586 (N_5586,N_5299,N_5018);
nand U5587 (N_5587,N_5400,N_5034);
nand U5588 (N_5588,N_5390,N_5134);
or U5589 (N_5589,N_5197,N_5046);
xor U5590 (N_5590,N_5243,N_5055);
nor U5591 (N_5591,N_5342,N_5112);
nor U5592 (N_5592,N_5424,N_5463);
nor U5593 (N_5593,N_5352,N_5232);
nor U5594 (N_5594,N_5011,N_5396);
xor U5595 (N_5595,N_5027,N_5233);
nand U5596 (N_5596,N_5021,N_5224);
and U5597 (N_5597,N_5466,N_5413);
nor U5598 (N_5598,N_5311,N_5019);
nand U5599 (N_5599,N_5444,N_5322);
nand U5600 (N_5600,N_5271,N_5065);
or U5601 (N_5601,N_5326,N_5272);
nand U5602 (N_5602,N_5184,N_5291);
or U5603 (N_5603,N_5125,N_5038);
nand U5604 (N_5604,N_5186,N_5384);
nor U5605 (N_5605,N_5392,N_5242);
xnor U5606 (N_5606,N_5073,N_5462);
nor U5607 (N_5607,N_5252,N_5234);
or U5608 (N_5608,N_5078,N_5340);
nand U5609 (N_5609,N_5323,N_5080);
xnor U5610 (N_5610,N_5218,N_5017);
and U5611 (N_5611,N_5416,N_5227);
nand U5612 (N_5612,N_5214,N_5454);
or U5613 (N_5613,N_5082,N_5283);
nor U5614 (N_5614,N_5247,N_5135);
nor U5615 (N_5615,N_5115,N_5094);
nand U5616 (N_5616,N_5117,N_5421);
xor U5617 (N_5617,N_5475,N_5162);
nand U5618 (N_5618,N_5157,N_5312);
and U5619 (N_5619,N_5083,N_5177);
and U5620 (N_5620,N_5300,N_5418);
and U5621 (N_5621,N_5258,N_5433);
nor U5622 (N_5622,N_5472,N_5248);
and U5623 (N_5623,N_5443,N_5096);
or U5624 (N_5624,N_5040,N_5440);
xnor U5625 (N_5625,N_5048,N_5156);
nand U5626 (N_5626,N_5136,N_5159);
xor U5627 (N_5627,N_5309,N_5414);
xor U5628 (N_5628,N_5341,N_5064);
nand U5629 (N_5629,N_5405,N_5047);
nor U5630 (N_5630,N_5477,N_5297);
xor U5631 (N_5631,N_5486,N_5155);
and U5632 (N_5632,N_5068,N_5295);
xor U5633 (N_5633,N_5212,N_5151);
nor U5634 (N_5634,N_5256,N_5043);
and U5635 (N_5635,N_5306,N_5126);
nand U5636 (N_5636,N_5100,N_5116);
xor U5637 (N_5637,N_5175,N_5205);
and U5638 (N_5638,N_5316,N_5004);
and U5639 (N_5639,N_5449,N_5436);
xnor U5640 (N_5640,N_5259,N_5369);
nand U5641 (N_5641,N_5262,N_5035);
xnor U5642 (N_5642,N_5077,N_5464);
or U5643 (N_5643,N_5163,N_5439);
xor U5644 (N_5644,N_5196,N_5372);
or U5645 (N_5645,N_5367,N_5058);
or U5646 (N_5646,N_5389,N_5255);
or U5647 (N_5647,N_5060,N_5032);
nor U5648 (N_5648,N_5460,N_5394);
and U5649 (N_5649,N_5366,N_5278);
nor U5650 (N_5650,N_5108,N_5029);
nor U5651 (N_5651,N_5288,N_5074);
and U5652 (N_5652,N_5138,N_5107);
nand U5653 (N_5653,N_5484,N_5279);
or U5654 (N_5654,N_5415,N_5182);
or U5655 (N_5655,N_5308,N_5172);
nor U5656 (N_5656,N_5325,N_5398);
xnor U5657 (N_5657,N_5261,N_5050);
nand U5658 (N_5658,N_5263,N_5169);
xnor U5659 (N_5659,N_5361,N_5275);
or U5660 (N_5660,N_5130,N_5203);
and U5661 (N_5661,N_5485,N_5069);
or U5662 (N_5662,N_5237,N_5010);
or U5663 (N_5663,N_5095,N_5296);
nor U5664 (N_5664,N_5101,N_5329);
nand U5665 (N_5665,N_5377,N_5432);
and U5666 (N_5666,N_5179,N_5429);
or U5667 (N_5667,N_5000,N_5076);
xor U5668 (N_5668,N_5007,N_5320);
or U5669 (N_5669,N_5493,N_5219);
xor U5670 (N_5670,N_5124,N_5106);
nor U5671 (N_5671,N_5222,N_5387);
and U5672 (N_5672,N_5370,N_5452);
and U5673 (N_5673,N_5153,N_5246);
nor U5674 (N_5674,N_5402,N_5109);
or U5675 (N_5675,N_5461,N_5098);
xnor U5676 (N_5676,N_5165,N_5206);
or U5677 (N_5677,N_5254,N_5092);
xnor U5678 (N_5678,N_5191,N_5490);
nand U5679 (N_5679,N_5399,N_5062);
xnor U5680 (N_5680,N_5281,N_5207);
nand U5681 (N_5681,N_5020,N_5105);
nor U5682 (N_5682,N_5054,N_5332);
and U5683 (N_5683,N_5409,N_5331);
or U5684 (N_5684,N_5426,N_5365);
nor U5685 (N_5685,N_5079,N_5441);
or U5686 (N_5686,N_5434,N_5131);
nor U5687 (N_5687,N_5448,N_5450);
nand U5688 (N_5688,N_5139,N_5127);
nor U5689 (N_5689,N_5408,N_5022);
nand U5690 (N_5690,N_5137,N_5494);
or U5691 (N_5691,N_5459,N_5285);
or U5692 (N_5692,N_5495,N_5497);
nor U5693 (N_5693,N_5168,N_5339);
and U5694 (N_5694,N_5456,N_5086);
nor U5695 (N_5695,N_5099,N_5359);
or U5696 (N_5696,N_5174,N_5063);
nor U5697 (N_5697,N_5391,N_5087);
nand U5698 (N_5698,N_5381,N_5190);
or U5699 (N_5699,N_5145,N_5351);
nand U5700 (N_5700,N_5417,N_5347);
xnor U5701 (N_5701,N_5324,N_5049);
nand U5702 (N_5702,N_5487,N_5208);
or U5703 (N_5703,N_5031,N_5236);
nand U5704 (N_5704,N_5170,N_5223);
xor U5705 (N_5705,N_5185,N_5294);
xor U5706 (N_5706,N_5422,N_5492);
xnor U5707 (N_5707,N_5176,N_5028);
xnor U5708 (N_5708,N_5009,N_5302);
nand U5709 (N_5709,N_5045,N_5318);
or U5710 (N_5710,N_5364,N_5453);
or U5711 (N_5711,N_5395,N_5158);
nor U5712 (N_5712,N_5091,N_5382);
nor U5713 (N_5713,N_5114,N_5213);
nand U5714 (N_5714,N_5024,N_5343);
nand U5715 (N_5715,N_5419,N_5133);
and U5716 (N_5716,N_5385,N_5482);
nand U5717 (N_5717,N_5088,N_5344);
xor U5718 (N_5718,N_5284,N_5319);
nand U5719 (N_5719,N_5447,N_5401);
and U5720 (N_5720,N_5346,N_5200);
nand U5721 (N_5721,N_5305,N_5251);
nand U5722 (N_5722,N_5358,N_5491);
and U5723 (N_5723,N_5189,N_5386);
or U5724 (N_5724,N_5075,N_5161);
nor U5725 (N_5725,N_5499,N_5355);
nand U5726 (N_5726,N_5420,N_5270);
nand U5727 (N_5727,N_5348,N_5025);
xor U5728 (N_5728,N_5148,N_5442);
nor U5729 (N_5729,N_5374,N_5240);
and U5730 (N_5730,N_5201,N_5081);
nand U5731 (N_5731,N_5036,N_5287);
nor U5732 (N_5732,N_5428,N_5183);
xnor U5733 (N_5733,N_5293,N_5345);
nand U5734 (N_5734,N_5173,N_5166);
or U5735 (N_5735,N_5120,N_5140);
or U5736 (N_5736,N_5089,N_5239);
and U5737 (N_5737,N_5333,N_5412);
xnor U5738 (N_5738,N_5303,N_5289);
or U5739 (N_5739,N_5307,N_5014);
xnor U5740 (N_5740,N_5301,N_5008);
xor U5741 (N_5741,N_5195,N_5474);
xor U5742 (N_5742,N_5427,N_5290);
xor U5743 (N_5743,N_5051,N_5337);
or U5744 (N_5744,N_5142,N_5129);
and U5745 (N_5745,N_5057,N_5273);
nand U5746 (N_5746,N_5210,N_5003);
or U5747 (N_5747,N_5006,N_5268);
and U5748 (N_5748,N_5123,N_5335);
and U5749 (N_5749,N_5171,N_5373);
or U5750 (N_5750,N_5457,N_5208);
and U5751 (N_5751,N_5483,N_5348);
nand U5752 (N_5752,N_5323,N_5364);
or U5753 (N_5753,N_5396,N_5244);
nand U5754 (N_5754,N_5361,N_5384);
xnor U5755 (N_5755,N_5236,N_5380);
nor U5756 (N_5756,N_5022,N_5423);
and U5757 (N_5757,N_5460,N_5008);
nand U5758 (N_5758,N_5262,N_5117);
xnor U5759 (N_5759,N_5028,N_5350);
nand U5760 (N_5760,N_5384,N_5133);
and U5761 (N_5761,N_5090,N_5185);
nand U5762 (N_5762,N_5447,N_5142);
nor U5763 (N_5763,N_5266,N_5341);
nor U5764 (N_5764,N_5144,N_5020);
nand U5765 (N_5765,N_5308,N_5076);
or U5766 (N_5766,N_5326,N_5033);
and U5767 (N_5767,N_5279,N_5034);
nand U5768 (N_5768,N_5329,N_5198);
nor U5769 (N_5769,N_5109,N_5255);
nor U5770 (N_5770,N_5327,N_5225);
or U5771 (N_5771,N_5433,N_5000);
xor U5772 (N_5772,N_5320,N_5468);
xnor U5773 (N_5773,N_5359,N_5113);
or U5774 (N_5774,N_5170,N_5283);
or U5775 (N_5775,N_5260,N_5296);
nand U5776 (N_5776,N_5319,N_5308);
nor U5777 (N_5777,N_5368,N_5288);
xnor U5778 (N_5778,N_5233,N_5323);
nand U5779 (N_5779,N_5299,N_5279);
nand U5780 (N_5780,N_5452,N_5444);
or U5781 (N_5781,N_5220,N_5256);
nand U5782 (N_5782,N_5021,N_5176);
xnor U5783 (N_5783,N_5338,N_5207);
and U5784 (N_5784,N_5485,N_5309);
nor U5785 (N_5785,N_5207,N_5004);
nand U5786 (N_5786,N_5343,N_5410);
nor U5787 (N_5787,N_5474,N_5065);
and U5788 (N_5788,N_5288,N_5292);
or U5789 (N_5789,N_5050,N_5251);
xnor U5790 (N_5790,N_5023,N_5170);
nand U5791 (N_5791,N_5058,N_5009);
xor U5792 (N_5792,N_5334,N_5027);
xor U5793 (N_5793,N_5437,N_5402);
or U5794 (N_5794,N_5176,N_5234);
and U5795 (N_5795,N_5312,N_5262);
or U5796 (N_5796,N_5171,N_5124);
nand U5797 (N_5797,N_5382,N_5400);
nor U5798 (N_5798,N_5292,N_5279);
nor U5799 (N_5799,N_5099,N_5068);
or U5800 (N_5800,N_5259,N_5495);
xnor U5801 (N_5801,N_5374,N_5443);
or U5802 (N_5802,N_5140,N_5119);
nand U5803 (N_5803,N_5191,N_5142);
xor U5804 (N_5804,N_5080,N_5053);
xor U5805 (N_5805,N_5432,N_5109);
xor U5806 (N_5806,N_5164,N_5334);
nand U5807 (N_5807,N_5424,N_5449);
nor U5808 (N_5808,N_5467,N_5136);
or U5809 (N_5809,N_5011,N_5441);
nand U5810 (N_5810,N_5341,N_5025);
xor U5811 (N_5811,N_5067,N_5309);
or U5812 (N_5812,N_5160,N_5044);
and U5813 (N_5813,N_5066,N_5004);
or U5814 (N_5814,N_5149,N_5334);
and U5815 (N_5815,N_5347,N_5458);
xnor U5816 (N_5816,N_5039,N_5204);
or U5817 (N_5817,N_5291,N_5163);
nand U5818 (N_5818,N_5316,N_5360);
or U5819 (N_5819,N_5496,N_5436);
and U5820 (N_5820,N_5217,N_5494);
nor U5821 (N_5821,N_5392,N_5138);
and U5822 (N_5822,N_5355,N_5373);
nand U5823 (N_5823,N_5237,N_5284);
nand U5824 (N_5824,N_5166,N_5408);
or U5825 (N_5825,N_5105,N_5442);
or U5826 (N_5826,N_5028,N_5483);
nor U5827 (N_5827,N_5412,N_5173);
nand U5828 (N_5828,N_5185,N_5472);
xnor U5829 (N_5829,N_5249,N_5200);
xnor U5830 (N_5830,N_5360,N_5382);
nor U5831 (N_5831,N_5319,N_5415);
or U5832 (N_5832,N_5206,N_5084);
nand U5833 (N_5833,N_5487,N_5016);
nor U5834 (N_5834,N_5462,N_5411);
nand U5835 (N_5835,N_5427,N_5298);
nand U5836 (N_5836,N_5415,N_5065);
nor U5837 (N_5837,N_5265,N_5482);
and U5838 (N_5838,N_5159,N_5134);
nor U5839 (N_5839,N_5354,N_5223);
or U5840 (N_5840,N_5264,N_5239);
nand U5841 (N_5841,N_5086,N_5320);
nor U5842 (N_5842,N_5255,N_5272);
or U5843 (N_5843,N_5300,N_5359);
nand U5844 (N_5844,N_5202,N_5052);
nand U5845 (N_5845,N_5364,N_5056);
xor U5846 (N_5846,N_5174,N_5237);
nor U5847 (N_5847,N_5350,N_5195);
nand U5848 (N_5848,N_5013,N_5092);
or U5849 (N_5849,N_5192,N_5148);
and U5850 (N_5850,N_5362,N_5077);
nor U5851 (N_5851,N_5013,N_5455);
xor U5852 (N_5852,N_5138,N_5082);
or U5853 (N_5853,N_5035,N_5145);
xnor U5854 (N_5854,N_5214,N_5254);
nor U5855 (N_5855,N_5149,N_5287);
or U5856 (N_5856,N_5392,N_5285);
nor U5857 (N_5857,N_5364,N_5133);
nor U5858 (N_5858,N_5048,N_5111);
and U5859 (N_5859,N_5386,N_5415);
and U5860 (N_5860,N_5419,N_5422);
or U5861 (N_5861,N_5339,N_5246);
nor U5862 (N_5862,N_5331,N_5068);
nand U5863 (N_5863,N_5466,N_5491);
nand U5864 (N_5864,N_5300,N_5128);
nor U5865 (N_5865,N_5140,N_5071);
and U5866 (N_5866,N_5413,N_5327);
nand U5867 (N_5867,N_5282,N_5178);
nor U5868 (N_5868,N_5349,N_5070);
nor U5869 (N_5869,N_5474,N_5341);
and U5870 (N_5870,N_5349,N_5233);
nand U5871 (N_5871,N_5420,N_5026);
or U5872 (N_5872,N_5419,N_5193);
and U5873 (N_5873,N_5213,N_5363);
nand U5874 (N_5874,N_5215,N_5240);
or U5875 (N_5875,N_5451,N_5225);
or U5876 (N_5876,N_5179,N_5018);
nand U5877 (N_5877,N_5451,N_5205);
and U5878 (N_5878,N_5215,N_5265);
and U5879 (N_5879,N_5262,N_5282);
or U5880 (N_5880,N_5326,N_5336);
nand U5881 (N_5881,N_5029,N_5475);
and U5882 (N_5882,N_5295,N_5039);
and U5883 (N_5883,N_5036,N_5103);
nand U5884 (N_5884,N_5339,N_5412);
or U5885 (N_5885,N_5406,N_5388);
or U5886 (N_5886,N_5326,N_5108);
nor U5887 (N_5887,N_5425,N_5242);
and U5888 (N_5888,N_5170,N_5441);
or U5889 (N_5889,N_5466,N_5047);
nand U5890 (N_5890,N_5391,N_5224);
or U5891 (N_5891,N_5164,N_5462);
or U5892 (N_5892,N_5280,N_5485);
or U5893 (N_5893,N_5034,N_5406);
nor U5894 (N_5894,N_5490,N_5456);
xor U5895 (N_5895,N_5318,N_5085);
or U5896 (N_5896,N_5236,N_5036);
nor U5897 (N_5897,N_5336,N_5098);
or U5898 (N_5898,N_5043,N_5059);
nand U5899 (N_5899,N_5351,N_5302);
or U5900 (N_5900,N_5007,N_5080);
and U5901 (N_5901,N_5114,N_5460);
xnor U5902 (N_5902,N_5119,N_5360);
nand U5903 (N_5903,N_5412,N_5115);
or U5904 (N_5904,N_5205,N_5358);
and U5905 (N_5905,N_5481,N_5451);
or U5906 (N_5906,N_5157,N_5251);
xor U5907 (N_5907,N_5390,N_5036);
and U5908 (N_5908,N_5264,N_5074);
xor U5909 (N_5909,N_5215,N_5449);
xor U5910 (N_5910,N_5218,N_5416);
xnor U5911 (N_5911,N_5034,N_5176);
and U5912 (N_5912,N_5082,N_5440);
nor U5913 (N_5913,N_5456,N_5024);
nor U5914 (N_5914,N_5192,N_5180);
xnor U5915 (N_5915,N_5202,N_5498);
or U5916 (N_5916,N_5380,N_5242);
xor U5917 (N_5917,N_5329,N_5010);
nand U5918 (N_5918,N_5335,N_5385);
or U5919 (N_5919,N_5116,N_5139);
or U5920 (N_5920,N_5165,N_5177);
nand U5921 (N_5921,N_5106,N_5310);
or U5922 (N_5922,N_5321,N_5309);
nor U5923 (N_5923,N_5332,N_5053);
xor U5924 (N_5924,N_5392,N_5308);
nor U5925 (N_5925,N_5168,N_5146);
or U5926 (N_5926,N_5182,N_5301);
xor U5927 (N_5927,N_5242,N_5310);
nand U5928 (N_5928,N_5000,N_5136);
and U5929 (N_5929,N_5041,N_5043);
xor U5930 (N_5930,N_5145,N_5316);
and U5931 (N_5931,N_5135,N_5261);
or U5932 (N_5932,N_5099,N_5006);
nor U5933 (N_5933,N_5125,N_5236);
nand U5934 (N_5934,N_5471,N_5104);
or U5935 (N_5935,N_5031,N_5182);
or U5936 (N_5936,N_5351,N_5380);
or U5937 (N_5937,N_5109,N_5143);
or U5938 (N_5938,N_5397,N_5372);
nor U5939 (N_5939,N_5428,N_5059);
and U5940 (N_5940,N_5323,N_5139);
nor U5941 (N_5941,N_5178,N_5306);
nand U5942 (N_5942,N_5307,N_5008);
or U5943 (N_5943,N_5094,N_5035);
nand U5944 (N_5944,N_5320,N_5405);
or U5945 (N_5945,N_5223,N_5210);
or U5946 (N_5946,N_5240,N_5261);
or U5947 (N_5947,N_5444,N_5122);
or U5948 (N_5948,N_5131,N_5205);
xor U5949 (N_5949,N_5366,N_5419);
xnor U5950 (N_5950,N_5233,N_5287);
xor U5951 (N_5951,N_5021,N_5007);
nand U5952 (N_5952,N_5174,N_5439);
xor U5953 (N_5953,N_5308,N_5361);
xor U5954 (N_5954,N_5061,N_5369);
xnor U5955 (N_5955,N_5015,N_5053);
and U5956 (N_5956,N_5377,N_5391);
nor U5957 (N_5957,N_5143,N_5336);
and U5958 (N_5958,N_5382,N_5324);
nor U5959 (N_5959,N_5177,N_5128);
or U5960 (N_5960,N_5149,N_5244);
nand U5961 (N_5961,N_5237,N_5033);
xor U5962 (N_5962,N_5239,N_5263);
and U5963 (N_5963,N_5234,N_5016);
xor U5964 (N_5964,N_5088,N_5013);
and U5965 (N_5965,N_5160,N_5195);
or U5966 (N_5966,N_5229,N_5118);
nor U5967 (N_5967,N_5364,N_5272);
or U5968 (N_5968,N_5439,N_5331);
or U5969 (N_5969,N_5153,N_5068);
nor U5970 (N_5970,N_5088,N_5409);
xnor U5971 (N_5971,N_5060,N_5329);
or U5972 (N_5972,N_5303,N_5133);
xor U5973 (N_5973,N_5280,N_5299);
nand U5974 (N_5974,N_5413,N_5053);
xnor U5975 (N_5975,N_5392,N_5094);
nand U5976 (N_5976,N_5151,N_5097);
nor U5977 (N_5977,N_5055,N_5205);
nand U5978 (N_5978,N_5296,N_5360);
xor U5979 (N_5979,N_5395,N_5032);
or U5980 (N_5980,N_5218,N_5306);
xor U5981 (N_5981,N_5448,N_5120);
or U5982 (N_5982,N_5036,N_5088);
and U5983 (N_5983,N_5461,N_5275);
or U5984 (N_5984,N_5124,N_5324);
nand U5985 (N_5985,N_5197,N_5452);
nor U5986 (N_5986,N_5109,N_5129);
and U5987 (N_5987,N_5400,N_5296);
nor U5988 (N_5988,N_5150,N_5361);
nor U5989 (N_5989,N_5467,N_5407);
nor U5990 (N_5990,N_5319,N_5265);
and U5991 (N_5991,N_5335,N_5092);
nor U5992 (N_5992,N_5110,N_5123);
or U5993 (N_5993,N_5266,N_5402);
nand U5994 (N_5994,N_5021,N_5422);
or U5995 (N_5995,N_5124,N_5299);
and U5996 (N_5996,N_5490,N_5081);
nor U5997 (N_5997,N_5111,N_5012);
and U5998 (N_5998,N_5215,N_5324);
nand U5999 (N_5999,N_5266,N_5303);
nor U6000 (N_6000,N_5929,N_5726);
nor U6001 (N_6001,N_5764,N_5584);
and U6002 (N_6002,N_5691,N_5760);
xnor U6003 (N_6003,N_5916,N_5632);
xor U6004 (N_6004,N_5544,N_5555);
or U6005 (N_6005,N_5828,N_5517);
and U6006 (N_6006,N_5700,N_5879);
or U6007 (N_6007,N_5933,N_5634);
nand U6008 (N_6008,N_5949,N_5821);
nand U6009 (N_6009,N_5559,N_5848);
xnor U6010 (N_6010,N_5988,N_5731);
nor U6011 (N_6011,N_5610,N_5585);
xor U6012 (N_6012,N_5947,N_5894);
nor U6013 (N_6013,N_5853,N_5950);
nor U6014 (N_6014,N_5506,N_5702);
nor U6015 (N_6015,N_5843,N_5914);
or U6016 (N_6016,N_5866,N_5613);
xnor U6017 (N_6017,N_5786,N_5687);
xor U6018 (N_6018,N_5908,N_5540);
and U6019 (N_6019,N_5653,N_5719);
nand U6020 (N_6020,N_5825,N_5831);
nor U6021 (N_6021,N_5685,N_5553);
nand U6022 (N_6022,N_5713,N_5514);
nand U6023 (N_6023,N_5619,N_5565);
nor U6024 (N_6024,N_5934,N_5795);
or U6025 (N_6025,N_5666,N_5679);
nand U6026 (N_6026,N_5961,N_5952);
nor U6027 (N_6027,N_5567,N_5995);
xnor U6028 (N_6028,N_5937,N_5596);
or U6029 (N_6029,N_5775,N_5510);
nand U6030 (N_6030,N_5751,N_5616);
xor U6031 (N_6031,N_5686,N_5812);
nor U6032 (N_6032,N_5993,N_5745);
xor U6033 (N_6033,N_5939,N_5851);
xor U6034 (N_6034,N_5975,N_5655);
and U6035 (N_6035,N_5829,N_5976);
nand U6036 (N_6036,N_5744,N_5902);
nand U6037 (N_6037,N_5926,N_5723);
and U6038 (N_6038,N_5862,N_5542);
nand U6039 (N_6039,N_5539,N_5991);
and U6040 (N_6040,N_5779,N_5999);
or U6041 (N_6041,N_5641,N_5675);
xnor U6042 (N_6042,N_5913,N_5529);
nand U6043 (N_6043,N_5872,N_5583);
nor U6044 (N_6044,N_5852,N_5622);
nand U6045 (N_6045,N_5919,N_5859);
and U6046 (N_6046,N_5577,N_5878);
nor U6047 (N_6047,N_5868,N_5763);
and U6048 (N_6048,N_5663,N_5614);
or U6049 (N_6049,N_5524,N_5730);
nor U6050 (N_6050,N_5736,N_5766);
nor U6051 (N_6051,N_5516,N_5692);
or U6052 (N_6052,N_5907,N_5773);
and U6053 (N_6053,N_5547,N_5587);
or U6054 (N_6054,N_5667,N_5782);
or U6055 (N_6055,N_5645,N_5841);
nand U6056 (N_6056,N_5912,N_5652);
xor U6057 (N_6057,N_5807,N_5793);
nor U6058 (N_6058,N_5591,N_5860);
xor U6059 (N_6059,N_5518,N_5981);
nand U6060 (N_6060,N_5874,N_5599);
xnor U6061 (N_6061,N_5617,N_5722);
xor U6062 (N_6062,N_5920,N_5800);
nand U6063 (N_6063,N_5978,N_5701);
or U6064 (N_6064,N_5799,N_5531);
xnor U6065 (N_6065,N_5625,N_5754);
xor U6066 (N_6066,N_5770,N_5811);
or U6067 (N_6067,N_5906,N_5562);
nand U6068 (N_6068,N_5564,N_5681);
xnor U6069 (N_6069,N_5966,N_5850);
nand U6070 (N_6070,N_5755,N_5554);
nor U6071 (N_6071,N_5855,N_5956);
xor U6072 (N_6072,N_5582,N_5987);
nor U6073 (N_6073,N_5750,N_5810);
or U6074 (N_6074,N_5758,N_5958);
nand U6075 (N_6075,N_5876,N_5910);
and U6076 (N_6076,N_5814,N_5594);
and U6077 (N_6077,N_5898,N_5818);
xor U6078 (N_6078,N_5572,N_5532);
xnor U6079 (N_6079,N_5636,N_5899);
nor U6080 (N_6080,N_5781,N_5593);
nand U6081 (N_6081,N_5545,N_5595);
nand U6082 (N_6082,N_5560,N_5802);
and U6083 (N_6083,N_5943,N_5541);
nor U6084 (N_6084,N_5832,N_5928);
or U6085 (N_6085,N_5710,N_5602);
nand U6086 (N_6086,N_5787,N_5967);
nor U6087 (N_6087,N_5566,N_5791);
or U6088 (N_6088,N_5670,N_5936);
nand U6089 (N_6089,N_5881,N_5656);
nor U6090 (N_6090,N_5705,N_5556);
and U6091 (N_6091,N_5715,N_5607);
nor U6092 (N_6092,N_5611,N_5671);
and U6093 (N_6093,N_5959,N_5895);
or U6094 (N_6094,N_5528,N_5889);
or U6095 (N_6095,N_5767,N_5930);
xnor U6096 (N_6096,N_5674,N_5873);
nand U6097 (N_6097,N_5627,N_5626);
nor U6098 (N_6098,N_5858,N_5648);
and U6099 (N_6099,N_5659,N_5618);
or U6100 (N_6100,N_5826,N_5985);
xnor U6101 (N_6101,N_5983,N_5523);
nand U6102 (N_6102,N_5884,N_5776);
or U6103 (N_6103,N_5624,N_5660);
or U6104 (N_6104,N_5854,N_5598);
xnor U6105 (N_6105,N_5844,N_5769);
nor U6106 (N_6106,N_5977,N_5921);
or U6107 (N_6107,N_5837,N_5957);
xor U6108 (N_6108,N_5798,N_5732);
xnor U6109 (N_6109,N_5882,N_5903);
nand U6110 (N_6110,N_5892,N_5534);
xnor U6111 (N_6111,N_5911,N_5546);
or U6112 (N_6112,N_5836,N_5570);
or U6113 (N_6113,N_5753,N_5604);
xnor U6114 (N_6114,N_5717,N_5998);
and U6115 (N_6115,N_5830,N_5661);
nor U6116 (N_6116,N_5951,N_5697);
or U6117 (N_6117,N_5849,N_5915);
xor U6118 (N_6118,N_5724,N_5623);
xor U6119 (N_6119,N_5521,N_5935);
nand U6120 (N_6120,N_5603,N_5527);
or U6121 (N_6121,N_5746,N_5606);
and U6122 (N_6122,N_5870,N_5633);
and U6123 (N_6123,N_5808,N_5643);
xor U6124 (N_6124,N_5944,N_5777);
xnor U6125 (N_6125,N_5927,N_5989);
nor U6126 (N_6126,N_5984,N_5561);
xnor U6127 (N_6127,N_5678,N_5945);
and U6128 (N_6128,N_5580,N_5897);
or U6129 (N_6129,N_5706,N_5778);
nor U6130 (N_6130,N_5890,N_5630);
nor U6131 (N_6131,N_5609,N_5846);
or U6132 (N_6132,N_5635,N_5568);
xor U6133 (N_6133,N_5768,N_5507);
and U6134 (N_6134,N_5864,N_5857);
and U6135 (N_6135,N_5709,N_5772);
and U6136 (N_6136,N_5662,N_5942);
and U6137 (N_6137,N_5809,N_5785);
nand U6138 (N_6138,N_5676,N_5941);
xnor U6139 (N_6139,N_5720,N_5824);
nand U6140 (N_6140,N_5579,N_5839);
and U6141 (N_6141,N_5869,N_5590);
and U6142 (N_6142,N_5955,N_5756);
nand U6143 (N_6143,N_5704,N_5718);
nor U6144 (N_6144,N_5642,N_5918);
and U6145 (N_6145,N_5707,N_5512);
or U6146 (N_6146,N_5640,N_5729);
or U6147 (N_6147,N_5789,N_5694);
xnor U6148 (N_6148,N_5924,N_5757);
nor U6149 (N_6149,N_5822,N_5639);
and U6150 (N_6150,N_5578,N_5574);
or U6151 (N_6151,N_5885,N_5817);
nor U6152 (N_6152,N_5628,N_5592);
nor U6153 (N_6153,N_5695,N_5714);
xnor U6154 (N_6154,N_5550,N_5806);
and U6155 (N_6155,N_5875,N_5980);
or U6156 (N_6156,N_5797,N_5522);
and U6157 (N_6157,N_5509,N_5815);
nor U6158 (N_6158,N_5548,N_5823);
nand U6159 (N_6159,N_5601,N_5833);
or U6160 (N_6160,N_5992,N_5699);
nand U6161 (N_6161,N_5552,N_5657);
nor U6162 (N_6162,N_5650,N_5741);
nor U6163 (N_6163,N_5673,N_5649);
nand U6164 (N_6164,N_5505,N_5917);
nand U6165 (N_6165,N_5589,N_5508);
or U6166 (N_6166,N_5813,N_5631);
and U6167 (N_6167,N_5896,N_5904);
or U6168 (N_6168,N_5804,N_5932);
nand U6169 (N_6169,N_5733,N_5549);
and U6170 (N_6170,N_5765,N_5712);
nor U6171 (N_6171,N_5743,N_5788);
or U6172 (N_6172,N_5557,N_5880);
nor U6173 (N_6173,N_5888,N_5996);
or U6174 (N_6174,N_5840,N_5835);
xor U6175 (N_6175,N_5605,N_5819);
nor U6176 (N_6176,N_5863,N_5759);
and U6177 (N_6177,N_5972,N_5997);
nor U6178 (N_6178,N_5971,N_5931);
nand U6179 (N_6179,N_5973,N_5535);
nand U6180 (N_6180,N_5986,N_5742);
nand U6181 (N_6181,N_5569,N_5537);
or U6182 (N_6182,N_5962,N_5734);
nand U6183 (N_6183,N_5612,N_5974);
and U6184 (N_6184,N_5677,N_5502);
nand U6185 (N_6185,N_5504,N_5689);
xor U6186 (N_6186,N_5865,N_5519);
and U6187 (N_6187,N_5615,N_5909);
xor U6188 (N_6188,N_5771,N_5576);
nor U6189 (N_6189,N_5644,N_5703);
nand U6190 (N_6190,N_5646,N_5905);
nand U6191 (N_6191,N_5748,N_5500);
xor U6192 (N_6192,N_5708,N_5965);
xor U6193 (N_6193,N_5842,N_5693);
xnor U6194 (N_6194,N_5827,N_5725);
nand U6195 (N_6195,N_5551,N_5600);
nor U6196 (N_6196,N_5683,N_5690);
xnor U6197 (N_6197,N_5665,N_5696);
or U6198 (N_6198,N_5900,N_5513);
nand U6199 (N_6199,N_5886,N_5739);
and U6200 (N_6200,N_5834,N_5780);
nor U6201 (N_6201,N_5716,N_5893);
nor U6202 (N_6202,N_5698,N_5761);
xnor U6203 (N_6203,N_5538,N_5654);
xor U6204 (N_6204,N_5563,N_5620);
nand U6205 (N_6205,N_5964,N_5536);
nand U6206 (N_6206,N_5515,N_5784);
or U6207 (N_6207,N_5621,N_5856);
and U6208 (N_6208,N_5680,N_5668);
and U6209 (N_6209,N_5588,N_5790);
or U6210 (N_6210,N_5970,N_5608);
nor U6211 (N_6211,N_5747,N_5658);
or U6212 (N_6212,N_5533,N_5586);
nor U6213 (N_6213,N_5525,N_5629);
and U6214 (N_6214,N_5940,N_5526);
xor U6215 (N_6215,N_5953,N_5948);
nor U6216 (N_6216,N_5638,N_5672);
and U6217 (N_6217,N_5573,N_5581);
and U6218 (N_6218,N_5954,N_5805);
nand U6219 (N_6219,N_5801,N_5503);
or U6220 (N_6220,N_5735,N_5543);
nand U6221 (N_6221,N_5922,N_5925);
and U6222 (N_6222,N_5558,N_5979);
or U6223 (N_6223,N_5688,N_5752);
or U6224 (N_6224,N_5575,N_5647);
nor U6225 (N_6225,N_5520,N_5796);
nor U6226 (N_6226,N_5762,N_5867);
nand U6227 (N_6227,N_5684,N_5901);
and U6228 (N_6228,N_5749,N_5721);
xnor U6229 (N_6229,N_5727,N_5820);
xor U6230 (N_6230,N_5923,N_5946);
xnor U6231 (N_6231,N_5845,N_5669);
nor U6232 (N_6232,N_5664,N_5597);
nor U6233 (N_6233,N_5501,N_5571);
nand U6234 (N_6234,N_5803,N_5682);
or U6235 (N_6235,N_5794,N_5728);
nand U6236 (N_6236,N_5838,N_5891);
nand U6237 (N_6237,N_5887,N_5960);
and U6238 (N_6238,N_5738,N_5938);
and U6239 (N_6239,N_5847,N_5740);
or U6240 (N_6240,N_5990,N_5883);
nand U6241 (N_6241,N_5651,N_5969);
nand U6242 (N_6242,N_5994,N_5861);
nor U6243 (N_6243,N_5530,N_5968);
nand U6244 (N_6244,N_5774,N_5982);
or U6245 (N_6245,N_5711,N_5816);
nor U6246 (N_6246,N_5783,N_5792);
or U6247 (N_6247,N_5511,N_5877);
xnor U6248 (N_6248,N_5963,N_5637);
nand U6249 (N_6249,N_5871,N_5737);
xor U6250 (N_6250,N_5524,N_5940);
nor U6251 (N_6251,N_5721,N_5871);
nor U6252 (N_6252,N_5596,N_5974);
and U6253 (N_6253,N_5701,N_5702);
xnor U6254 (N_6254,N_5750,N_5584);
xnor U6255 (N_6255,N_5544,N_5857);
or U6256 (N_6256,N_5626,N_5950);
xnor U6257 (N_6257,N_5981,N_5741);
and U6258 (N_6258,N_5787,N_5859);
xnor U6259 (N_6259,N_5555,N_5610);
xnor U6260 (N_6260,N_5980,N_5987);
nor U6261 (N_6261,N_5784,N_5728);
nor U6262 (N_6262,N_5736,N_5634);
xor U6263 (N_6263,N_5717,N_5678);
or U6264 (N_6264,N_5901,N_5798);
or U6265 (N_6265,N_5707,N_5641);
xor U6266 (N_6266,N_5535,N_5907);
nor U6267 (N_6267,N_5738,N_5860);
xor U6268 (N_6268,N_5611,N_5924);
nor U6269 (N_6269,N_5545,N_5582);
xor U6270 (N_6270,N_5829,N_5534);
or U6271 (N_6271,N_5548,N_5888);
xor U6272 (N_6272,N_5859,N_5576);
or U6273 (N_6273,N_5612,N_5729);
or U6274 (N_6274,N_5946,N_5977);
xor U6275 (N_6275,N_5634,N_5790);
nand U6276 (N_6276,N_5888,N_5950);
and U6277 (N_6277,N_5888,N_5580);
xor U6278 (N_6278,N_5557,N_5563);
xnor U6279 (N_6279,N_5687,N_5927);
or U6280 (N_6280,N_5794,N_5881);
nor U6281 (N_6281,N_5731,N_5605);
xnor U6282 (N_6282,N_5829,N_5888);
xnor U6283 (N_6283,N_5573,N_5789);
nand U6284 (N_6284,N_5606,N_5661);
nor U6285 (N_6285,N_5817,N_5574);
nand U6286 (N_6286,N_5758,N_5723);
and U6287 (N_6287,N_5663,N_5690);
nor U6288 (N_6288,N_5531,N_5951);
xnor U6289 (N_6289,N_5802,N_5623);
xor U6290 (N_6290,N_5934,N_5507);
xnor U6291 (N_6291,N_5703,N_5672);
or U6292 (N_6292,N_5704,N_5592);
nand U6293 (N_6293,N_5570,N_5770);
nor U6294 (N_6294,N_5946,N_5526);
nand U6295 (N_6295,N_5979,N_5807);
nand U6296 (N_6296,N_5939,N_5977);
or U6297 (N_6297,N_5699,N_5525);
nor U6298 (N_6298,N_5935,N_5635);
and U6299 (N_6299,N_5729,N_5859);
or U6300 (N_6300,N_5986,N_5672);
xnor U6301 (N_6301,N_5684,N_5642);
nor U6302 (N_6302,N_5830,N_5767);
or U6303 (N_6303,N_5923,N_5931);
xnor U6304 (N_6304,N_5539,N_5620);
or U6305 (N_6305,N_5638,N_5593);
xor U6306 (N_6306,N_5928,N_5530);
nor U6307 (N_6307,N_5547,N_5640);
and U6308 (N_6308,N_5765,N_5865);
xor U6309 (N_6309,N_5558,N_5843);
nor U6310 (N_6310,N_5799,N_5607);
nand U6311 (N_6311,N_5730,N_5923);
or U6312 (N_6312,N_5885,N_5903);
xor U6313 (N_6313,N_5713,N_5827);
xor U6314 (N_6314,N_5598,N_5569);
or U6315 (N_6315,N_5862,N_5793);
nor U6316 (N_6316,N_5918,N_5659);
xnor U6317 (N_6317,N_5680,N_5582);
xor U6318 (N_6318,N_5769,N_5809);
or U6319 (N_6319,N_5584,N_5524);
or U6320 (N_6320,N_5868,N_5508);
or U6321 (N_6321,N_5852,N_5636);
or U6322 (N_6322,N_5994,N_5744);
nand U6323 (N_6323,N_5953,N_5555);
nor U6324 (N_6324,N_5787,N_5889);
nand U6325 (N_6325,N_5565,N_5889);
or U6326 (N_6326,N_5628,N_5552);
nor U6327 (N_6327,N_5547,N_5907);
xor U6328 (N_6328,N_5829,N_5885);
xor U6329 (N_6329,N_5551,N_5837);
xnor U6330 (N_6330,N_5836,N_5502);
and U6331 (N_6331,N_5709,N_5768);
nand U6332 (N_6332,N_5752,N_5773);
and U6333 (N_6333,N_5683,N_5814);
and U6334 (N_6334,N_5908,N_5725);
nor U6335 (N_6335,N_5751,N_5997);
xnor U6336 (N_6336,N_5925,N_5670);
xnor U6337 (N_6337,N_5753,N_5509);
or U6338 (N_6338,N_5954,N_5730);
and U6339 (N_6339,N_5856,N_5597);
and U6340 (N_6340,N_5745,N_5731);
and U6341 (N_6341,N_5816,N_5787);
and U6342 (N_6342,N_5557,N_5586);
xnor U6343 (N_6343,N_5549,N_5502);
or U6344 (N_6344,N_5867,N_5669);
nand U6345 (N_6345,N_5689,N_5698);
xnor U6346 (N_6346,N_5590,N_5520);
nor U6347 (N_6347,N_5879,N_5685);
nand U6348 (N_6348,N_5545,N_5616);
nand U6349 (N_6349,N_5666,N_5570);
nand U6350 (N_6350,N_5549,N_5942);
nor U6351 (N_6351,N_5541,N_5902);
xor U6352 (N_6352,N_5822,N_5738);
nor U6353 (N_6353,N_5819,N_5767);
and U6354 (N_6354,N_5716,N_5576);
or U6355 (N_6355,N_5789,N_5888);
and U6356 (N_6356,N_5932,N_5957);
or U6357 (N_6357,N_5948,N_5971);
or U6358 (N_6358,N_5518,N_5686);
and U6359 (N_6359,N_5507,N_5839);
and U6360 (N_6360,N_5583,N_5670);
xor U6361 (N_6361,N_5906,N_5782);
nand U6362 (N_6362,N_5886,N_5618);
xnor U6363 (N_6363,N_5549,N_5839);
xnor U6364 (N_6364,N_5625,N_5608);
nand U6365 (N_6365,N_5932,N_5926);
xnor U6366 (N_6366,N_5711,N_5739);
nand U6367 (N_6367,N_5936,N_5769);
nand U6368 (N_6368,N_5890,N_5553);
xnor U6369 (N_6369,N_5533,N_5887);
xnor U6370 (N_6370,N_5678,N_5899);
nor U6371 (N_6371,N_5550,N_5818);
and U6372 (N_6372,N_5659,N_5757);
or U6373 (N_6373,N_5504,N_5926);
xor U6374 (N_6374,N_5967,N_5519);
nor U6375 (N_6375,N_5787,N_5769);
nand U6376 (N_6376,N_5946,N_5685);
xor U6377 (N_6377,N_5798,N_5975);
xnor U6378 (N_6378,N_5772,N_5731);
nand U6379 (N_6379,N_5823,N_5569);
or U6380 (N_6380,N_5788,N_5585);
and U6381 (N_6381,N_5706,N_5887);
and U6382 (N_6382,N_5746,N_5757);
or U6383 (N_6383,N_5892,N_5584);
nand U6384 (N_6384,N_5511,N_5957);
xnor U6385 (N_6385,N_5936,N_5925);
xnor U6386 (N_6386,N_5535,N_5777);
nand U6387 (N_6387,N_5796,N_5618);
nor U6388 (N_6388,N_5947,N_5669);
and U6389 (N_6389,N_5844,N_5765);
nand U6390 (N_6390,N_5914,N_5511);
nor U6391 (N_6391,N_5827,N_5986);
and U6392 (N_6392,N_5872,N_5550);
nand U6393 (N_6393,N_5707,N_5822);
xnor U6394 (N_6394,N_5931,N_5639);
nor U6395 (N_6395,N_5908,N_5889);
xor U6396 (N_6396,N_5737,N_5968);
or U6397 (N_6397,N_5778,N_5696);
nand U6398 (N_6398,N_5998,N_5867);
nand U6399 (N_6399,N_5741,N_5581);
and U6400 (N_6400,N_5717,N_5708);
and U6401 (N_6401,N_5555,N_5862);
nor U6402 (N_6402,N_5892,N_5512);
or U6403 (N_6403,N_5503,N_5923);
nor U6404 (N_6404,N_5914,N_5571);
nand U6405 (N_6405,N_5517,N_5629);
nor U6406 (N_6406,N_5545,N_5751);
and U6407 (N_6407,N_5711,N_5603);
and U6408 (N_6408,N_5686,N_5805);
or U6409 (N_6409,N_5831,N_5707);
or U6410 (N_6410,N_5560,N_5700);
xnor U6411 (N_6411,N_5855,N_5611);
nor U6412 (N_6412,N_5598,N_5581);
or U6413 (N_6413,N_5510,N_5642);
xnor U6414 (N_6414,N_5896,N_5900);
and U6415 (N_6415,N_5748,N_5511);
nand U6416 (N_6416,N_5792,N_5940);
nand U6417 (N_6417,N_5664,N_5862);
nor U6418 (N_6418,N_5551,N_5899);
nand U6419 (N_6419,N_5982,N_5988);
or U6420 (N_6420,N_5576,N_5673);
xnor U6421 (N_6421,N_5792,N_5739);
or U6422 (N_6422,N_5533,N_5710);
or U6423 (N_6423,N_5659,N_5803);
or U6424 (N_6424,N_5589,N_5534);
nor U6425 (N_6425,N_5717,N_5620);
and U6426 (N_6426,N_5612,N_5897);
xnor U6427 (N_6427,N_5633,N_5522);
nor U6428 (N_6428,N_5683,N_5697);
and U6429 (N_6429,N_5587,N_5899);
xnor U6430 (N_6430,N_5786,N_5557);
and U6431 (N_6431,N_5883,N_5828);
nand U6432 (N_6432,N_5788,N_5975);
nor U6433 (N_6433,N_5978,N_5970);
and U6434 (N_6434,N_5991,N_5653);
and U6435 (N_6435,N_5667,N_5731);
xor U6436 (N_6436,N_5538,N_5626);
or U6437 (N_6437,N_5779,N_5927);
nand U6438 (N_6438,N_5576,N_5561);
and U6439 (N_6439,N_5856,N_5941);
nand U6440 (N_6440,N_5752,N_5509);
nor U6441 (N_6441,N_5893,N_5918);
nand U6442 (N_6442,N_5962,N_5765);
xor U6443 (N_6443,N_5919,N_5695);
and U6444 (N_6444,N_5579,N_5793);
nor U6445 (N_6445,N_5780,N_5657);
and U6446 (N_6446,N_5614,N_5621);
or U6447 (N_6447,N_5630,N_5696);
nor U6448 (N_6448,N_5968,N_5588);
nand U6449 (N_6449,N_5684,N_5763);
and U6450 (N_6450,N_5504,N_5974);
and U6451 (N_6451,N_5993,N_5691);
or U6452 (N_6452,N_5894,N_5906);
and U6453 (N_6453,N_5939,N_5850);
nand U6454 (N_6454,N_5676,N_5884);
nand U6455 (N_6455,N_5971,N_5533);
xor U6456 (N_6456,N_5679,N_5544);
and U6457 (N_6457,N_5786,N_5913);
and U6458 (N_6458,N_5778,N_5673);
xnor U6459 (N_6459,N_5991,N_5681);
or U6460 (N_6460,N_5619,N_5709);
xor U6461 (N_6461,N_5967,N_5625);
and U6462 (N_6462,N_5555,N_5899);
xnor U6463 (N_6463,N_5766,N_5542);
nand U6464 (N_6464,N_5949,N_5847);
and U6465 (N_6465,N_5730,N_5529);
or U6466 (N_6466,N_5671,N_5547);
xor U6467 (N_6467,N_5514,N_5791);
xnor U6468 (N_6468,N_5930,N_5954);
xnor U6469 (N_6469,N_5780,N_5970);
nor U6470 (N_6470,N_5980,N_5525);
and U6471 (N_6471,N_5951,N_5514);
and U6472 (N_6472,N_5545,N_5758);
xnor U6473 (N_6473,N_5732,N_5567);
or U6474 (N_6474,N_5882,N_5711);
nor U6475 (N_6475,N_5650,N_5843);
xor U6476 (N_6476,N_5849,N_5622);
and U6477 (N_6477,N_5561,N_5642);
or U6478 (N_6478,N_5704,N_5850);
or U6479 (N_6479,N_5758,N_5740);
xnor U6480 (N_6480,N_5573,N_5513);
nor U6481 (N_6481,N_5944,N_5788);
or U6482 (N_6482,N_5899,N_5963);
and U6483 (N_6483,N_5557,N_5841);
xor U6484 (N_6484,N_5642,N_5606);
nor U6485 (N_6485,N_5787,N_5764);
nor U6486 (N_6486,N_5907,N_5515);
and U6487 (N_6487,N_5873,N_5592);
or U6488 (N_6488,N_5783,N_5758);
nand U6489 (N_6489,N_5962,N_5760);
and U6490 (N_6490,N_5610,N_5668);
nor U6491 (N_6491,N_5514,N_5886);
nor U6492 (N_6492,N_5826,N_5999);
or U6493 (N_6493,N_5568,N_5784);
nand U6494 (N_6494,N_5688,N_5872);
and U6495 (N_6495,N_5564,N_5677);
nand U6496 (N_6496,N_5527,N_5762);
nand U6497 (N_6497,N_5983,N_5504);
nor U6498 (N_6498,N_5847,N_5540);
or U6499 (N_6499,N_5892,N_5948);
or U6500 (N_6500,N_6497,N_6356);
nor U6501 (N_6501,N_6074,N_6431);
and U6502 (N_6502,N_6077,N_6081);
nand U6503 (N_6503,N_6128,N_6309);
nand U6504 (N_6504,N_6275,N_6266);
xnor U6505 (N_6505,N_6348,N_6480);
xnor U6506 (N_6506,N_6486,N_6211);
nor U6507 (N_6507,N_6227,N_6188);
nor U6508 (N_6508,N_6463,N_6137);
nor U6509 (N_6509,N_6132,N_6263);
and U6510 (N_6510,N_6235,N_6057);
nand U6511 (N_6511,N_6114,N_6388);
and U6512 (N_6512,N_6375,N_6103);
and U6513 (N_6513,N_6230,N_6250);
xor U6514 (N_6514,N_6038,N_6201);
nand U6515 (N_6515,N_6018,N_6214);
xor U6516 (N_6516,N_6402,N_6244);
nand U6517 (N_6517,N_6179,N_6198);
and U6518 (N_6518,N_6096,N_6116);
and U6519 (N_6519,N_6156,N_6025);
xor U6520 (N_6520,N_6138,N_6086);
and U6521 (N_6521,N_6424,N_6273);
and U6522 (N_6522,N_6104,N_6499);
and U6523 (N_6523,N_6110,N_6452);
xor U6524 (N_6524,N_6127,N_6233);
xor U6525 (N_6525,N_6400,N_6457);
and U6526 (N_6526,N_6279,N_6195);
or U6527 (N_6527,N_6405,N_6082);
or U6528 (N_6528,N_6395,N_6217);
or U6529 (N_6529,N_6231,N_6146);
and U6530 (N_6530,N_6390,N_6352);
or U6531 (N_6531,N_6428,N_6306);
and U6532 (N_6532,N_6350,N_6097);
nor U6533 (N_6533,N_6087,N_6341);
xnor U6534 (N_6534,N_6307,N_6248);
nand U6535 (N_6535,N_6184,N_6069);
nor U6536 (N_6536,N_6385,N_6041);
or U6537 (N_6537,N_6310,N_6102);
nand U6538 (N_6538,N_6487,N_6076);
nor U6539 (N_6539,N_6362,N_6139);
nand U6540 (N_6540,N_6006,N_6118);
or U6541 (N_6541,N_6247,N_6289);
xor U6542 (N_6542,N_6414,N_6245);
nand U6543 (N_6543,N_6084,N_6320);
nand U6544 (N_6544,N_6048,N_6064);
or U6545 (N_6545,N_6399,N_6010);
nand U6546 (N_6546,N_6040,N_6444);
nor U6547 (N_6547,N_6257,N_6152);
xor U6548 (N_6548,N_6291,N_6148);
or U6549 (N_6549,N_6333,N_6387);
nand U6550 (N_6550,N_6462,N_6197);
or U6551 (N_6551,N_6377,N_6368);
nand U6552 (N_6552,N_6216,N_6080);
nor U6553 (N_6553,N_6191,N_6366);
and U6554 (N_6554,N_6369,N_6353);
and U6555 (N_6555,N_6327,N_6088);
nand U6556 (N_6556,N_6277,N_6408);
or U6557 (N_6557,N_6049,N_6029);
or U6558 (N_6558,N_6060,N_6254);
and U6559 (N_6559,N_6354,N_6446);
and U6560 (N_6560,N_6406,N_6447);
and U6561 (N_6561,N_6202,N_6099);
or U6562 (N_6562,N_6409,N_6240);
nand U6563 (N_6563,N_6459,N_6092);
and U6564 (N_6564,N_6062,N_6160);
xnor U6565 (N_6565,N_6030,N_6458);
or U6566 (N_6566,N_6304,N_6044);
nor U6567 (N_6567,N_6050,N_6416);
and U6568 (N_6568,N_6477,N_6445);
or U6569 (N_6569,N_6219,N_6008);
nor U6570 (N_6570,N_6415,N_6024);
and U6571 (N_6571,N_6465,N_6422);
nor U6572 (N_6572,N_6126,N_6376);
or U6573 (N_6573,N_6013,N_6393);
xor U6574 (N_6574,N_6051,N_6488);
nor U6575 (N_6575,N_6209,N_6281);
or U6576 (N_6576,N_6331,N_6261);
and U6577 (N_6577,N_6164,N_6059);
xnor U6578 (N_6578,N_6206,N_6323);
xor U6579 (N_6579,N_6015,N_6367);
and U6580 (N_6580,N_6176,N_6192);
nand U6581 (N_6581,N_6055,N_6482);
nor U6582 (N_6582,N_6089,N_6267);
nor U6583 (N_6583,N_6251,N_6056);
xnor U6584 (N_6584,N_6265,N_6053);
and U6585 (N_6585,N_6063,N_6221);
and U6586 (N_6586,N_6287,N_6034);
nor U6587 (N_6587,N_6449,N_6259);
or U6588 (N_6588,N_6067,N_6370);
nand U6589 (N_6589,N_6363,N_6210);
nand U6590 (N_6590,N_6299,N_6478);
or U6591 (N_6591,N_6429,N_6154);
nor U6592 (N_6592,N_6145,N_6141);
nand U6593 (N_6593,N_6173,N_6364);
nand U6594 (N_6594,N_6317,N_6434);
nand U6595 (N_6595,N_6213,N_6319);
xor U6596 (N_6596,N_6288,N_6149);
nor U6597 (N_6597,N_6316,N_6218);
nand U6598 (N_6598,N_6335,N_6294);
and U6599 (N_6599,N_6430,N_6091);
nand U6600 (N_6600,N_6283,N_6085);
nor U6601 (N_6601,N_6113,N_6384);
nand U6602 (N_6602,N_6124,N_6303);
nand U6603 (N_6603,N_6404,N_6485);
nand U6604 (N_6604,N_6374,N_6282);
nand U6605 (N_6605,N_6391,N_6318);
nor U6606 (N_6606,N_6474,N_6016);
nand U6607 (N_6607,N_6397,N_6403);
nor U6608 (N_6608,N_6337,N_6125);
nor U6609 (N_6609,N_6361,N_6065);
nor U6610 (N_6610,N_6153,N_6360);
or U6611 (N_6611,N_6225,N_6420);
xor U6612 (N_6612,N_6413,N_6163);
and U6613 (N_6613,N_6302,N_6454);
nand U6614 (N_6614,N_6054,N_6365);
and U6615 (N_6615,N_6421,N_6494);
xnor U6616 (N_6616,N_6472,N_6329);
nand U6617 (N_6617,N_6439,N_6185);
nor U6618 (N_6618,N_6242,N_6491);
or U6619 (N_6619,N_6456,N_6336);
nor U6620 (N_6620,N_6269,N_6020);
xor U6621 (N_6621,N_6204,N_6111);
nand U6622 (N_6622,N_6171,N_6342);
or U6623 (N_6623,N_6070,N_6151);
nand U6624 (N_6624,N_6121,N_6328);
nor U6625 (N_6625,N_6140,N_6433);
xor U6626 (N_6626,N_6432,N_6134);
xnor U6627 (N_6627,N_6107,N_6223);
or U6628 (N_6628,N_6479,N_6078);
or U6629 (N_6629,N_6410,N_6311);
and U6630 (N_6630,N_6483,N_6312);
nand U6631 (N_6631,N_6313,N_6167);
and U6632 (N_6632,N_6386,N_6441);
and U6633 (N_6633,N_6425,N_6004);
xor U6634 (N_6634,N_6464,N_6412);
or U6635 (N_6635,N_6493,N_6372);
nand U6636 (N_6636,N_6448,N_6005);
nor U6637 (N_6637,N_6325,N_6042);
xnor U6638 (N_6638,N_6150,N_6026);
nor U6639 (N_6639,N_6205,N_6243);
or U6640 (N_6640,N_6011,N_6438);
and U6641 (N_6641,N_6298,N_6270);
xor U6642 (N_6642,N_6481,N_6161);
and U6643 (N_6643,N_6268,N_6358);
xnor U6644 (N_6644,N_6398,N_6182);
or U6645 (N_6645,N_6039,N_6133);
xor U6646 (N_6646,N_6093,N_6009);
xor U6647 (N_6647,N_6332,N_6003);
nor U6648 (N_6648,N_6338,N_6278);
and U6649 (N_6649,N_6189,N_6468);
and U6650 (N_6650,N_6083,N_6181);
and U6651 (N_6651,N_6371,N_6061);
and U6652 (N_6652,N_6417,N_6274);
nor U6653 (N_6653,N_6382,N_6471);
xor U6654 (N_6654,N_6271,N_6381);
or U6655 (N_6655,N_6222,N_6224);
nand U6656 (N_6656,N_6120,N_6285);
xnor U6657 (N_6657,N_6451,N_6172);
nand U6658 (N_6658,N_6200,N_6334);
and U6659 (N_6659,N_6105,N_6007);
nor U6660 (N_6660,N_6293,N_6072);
and U6661 (N_6661,N_6258,N_6427);
or U6662 (N_6662,N_6196,N_6476);
nor U6663 (N_6663,N_6071,N_6068);
or U6664 (N_6664,N_6117,N_6455);
nor U6665 (N_6665,N_6359,N_6389);
nand U6666 (N_6666,N_6357,N_6392);
and U6667 (N_6667,N_6495,N_6344);
nor U6668 (N_6668,N_6147,N_6186);
or U6669 (N_6669,N_6058,N_6276);
nor U6670 (N_6670,N_6380,N_6045);
xor U6671 (N_6671,N_6467,N_6119);
xnor U6672 (N_6672,N_6101,N_6453);
nor U6673 (N_6673,N_6321,N_6256);
xor U6674 (N_6674,N_6340,N_6193);
nor U6675 (N_6675,N_6002,N_6158);
nand U6676 (N_6676,N_6295,N_6166);
nor U6677 (N_6677,N_6346,N_6228);
nand U6678 (N_6678,N_6023,N_6489);
or U6679 (N_6679,N_6426,N_6098);
or U6680 (N_6680,N_6203,N_6411);
and U6681 (N_6681,N_6450,N_6212);
and U6682 (N_6682,N_6330,N_6470);
xor U6683 (N_6683,N_6090,N_6165);
or U6684 (N_6684,N_6326,N_6112);
nor U6685 (N_6685,N_6143,N_6052);
xor U6686 (N_6686,N_6496,N_6207);
xnor U6687 (N_6687,N_6178,N_6183);
xor U6688 (N_6688,N_6473,N_6260);
nor U6689 (N_6689,N_6226,N_6234);
nand U6690 (N_6690,N_6347,N_6252);
and U6691 (N_6691,N_6162,N_6168);
and U6692 (N_6692,N_6027,N_6100);
nand U6693 (N_6693,N_6157,N_6000);
or U6694 (N_6694,N_6046,N_6272);
nor U6695 (N_6695,N_6180,N_6075);
nand U6696 (N_6696,N_6440,N_6300);
nand U6697 (N_6697,N_6383,N_6229);
xor U6698 (N_6698,N_6142,N_6407);
or U6699 (N_6699,N_6419,N_6322);
xor U6700 (N_6700,N_6136,N_6094);
or U6701 (N_6701,N_6014,N_6190);
and U6702 (N_6702,N_6033,N_6264);
nand U6703 (N_6703,N_6017,N_6079);
and U6704 (N_6704,N_6296,N_6442);
and U6705 (N_6705,N_6066,N_6253);
or U6706 (N_6706,N_6170,N_6109);
nor U6707 (N_6707,N_6305,N_6423);
nor U6708 (N_6708,N_6394,N_6498);
nand U6709 (N_6709,N_6469,N_6255);
nand U6710 (N_6710,N_6246,N_6418);
nand U6711 (N_6711,N_6355,N_6012);
xor U6712 (N_6712,N_6351,N_6437);
and U6713 (N_6713,N_6108,N_6492);
or U6714 (N_6714,N_6031,N_6290);
xnor U6715 (N_6715,N_6155,N_6106);
and U6716 (N_6716,N_6436,N_6396);
nor U6717 (N_6717,N_6021,N_6194);
or U6718 (N_6718,N_6208,N_6187);
or U6719 (N_6719,N_6199,N_6135);
or U6720 (N_6720,N_6308,N_6324);
xor U6721 (N_6721,N_6175,N_6028);
xnor U6722 (N_6722,N_6460,N_6466);
nand U6723 (N_6723,N_6301,N_6314);
nand U6724 (N_6724,N_6122,N_6236);
xnor U6725 (N_6725,N_6232,N_6032);
xnor U6726 (N_6726,N_6339,N_6095);
or U6727 (N_6727,N_6262,N_6022);
xnor U6728 (N_6728,N_6129,N_6001);
and U6729 (N_6729,N_6284,N_6159);
nand U6730 (N_6730,N_6490,N_6019);
nor U6731 (N_6731,N_6401,N_6349);
nor U6732 (N_6732,N_6315,N_6345);
nor U6733 (N_6733,N_6435,N_6443);
or U6734 (N_6734,N_6373,N_6239);
xor U6735 (N_6735,N_6047,N_6144);
xnor U6736 (N_6736,N_6475,N_6115);
nand U6737 (N_6737,N_6036,N_6379);
nor U6738 (N_6738,N_6073,N_6174);
xor U6739 (N_6739,N_6237,N_6378);
nor U6740 (N_6740,N_6241,N_6037);
nor U6741 (N_6741,N_6220,N_6043);
and U6742 (N_6742,N_6461,N_6238);
nand U6743 (N_6743,N_6280,N_6297);
or U6744 (N_6744,N_6292,N_6286);
nand U6745 (N_6745,N_6484,N_6131);
and U6746 (N_6746,N_6035,N_6343);
and U6747 (N_6747,N_6123,N_6215);
and U6748 (N_6748,N_6249,N_6169);
nor U6749 (N_6749,N_6177,N_6130);
or U6750 (N_6750,N_6055,N_6458);
nor U6751 (N_6751,N_6158,N_6199);
nor U6752 (N_6752,N_6328,N_6367);
xnor U6753 (N_6753,N_6048,N_6115);
nand U6754 (N_6754,N_6110,N_6227);
xor U6755 (N_6755,N_6387,N_6111);
and U6756 (N_6756,N_6357,N_6269);
nor U6757 (N_6757,N_6143,N_6359);
nand U6758 (N_6758,N_6016,N_6082);
nor U6759 (N_6759,N_6246,N_6006);
xnor U6760 (N_6760,N_6087,N_6226);
xnor U6761 (N_6761,N_6067,N_6417);
xor U6762 (N_6762,N_6379,N_6381);
nor U6763 (N_6763,N_6490,N_6401);
and U6764 (N_6764,N_6250,N_6101);
nand U6765 (N_6765,N_6334,N_6247);
xor U6766 (N_6766,N_6178,N_6344);
nor U6767 (N_6767,N_6131,N_6291);
xnor U6768 (N_6768,N_6255,N_6408);
nor U6769 (N_6769,N_6077,N_6382);
nand U6770 (N_6770,N_6305,N_6302);
xor U6771 (N_6771,N_6321,N_6476);
xor U6772 (N_6772,N_6114,N_6381);
and U6773 (N_6773,N_6234,N_6313);
and U6774 (N_6774,N_6167,N_6355);
or U6775 (N_6775,N_6220,N_6323);
nor U6776 (N_6776,N_6186,N_6066);
xnor U6777 (N_6777,N_6078,N_6033);
and U6778 (N_6778,N_6305,N_6065);
or U6779 (N_6779,N_6463,N_6195);
xor U6780 (N_6780,N_6216,N_6227);
or U6781 (N_6781,N_6268,N_6141);
nor U6782 (N_6782,N_6105,N_6419);
and U6783 (N_6783,N_6381,N_6283);
xor U6784 (N_6784,N_6069,N_6238);
xnor U6785 (N_6785,N_6226,N_6175);
xnor U6786 (N_6786,N_6172,N_6218);
xor U6787 (N_6787,N_6058,N_6129);
or U6788 (N_6788,N_6372,N_6120);
xor U6789 (N_6789,N_6111,N_6433);
or U6790 (N_6790,N_6229,N_6196);
nand U6791 (N_6791,N_6421,N_6230);
or U6792 (N_6792,N_6404,N_6026);
or U6793 (N_6793,N_6348,N_6060);
nand U6794 (N_6794,N_6272,N_6186);
and U6795 (N_6795,N_6374,N_6179);
nor U6796 (N_6796,N_6026,N_6104);
nor U6797 (N_6797,N_6375,N_6200);
and U6798 (N_6798,N_6368,N_6307);
and U6799 (N_6799,N_6315,N_6273);
nor U6800 (N_6800,N_6022,N_6065);
nand U6801 (N_6801,N_6285,N_6002);
nor U6802 (N_6802,N_6308,N_6427);
xnor U6803 (N_6803,N_6466,N_6376);
nor U6804 (N_6804,N_6267,N_6439);
nand U6805 (N_6805,N_6286,N_6468);
or U6806 (N_6806,N_6326,N_6336);
xnor U6807 (N_6807,N_6067,N_6274);
nor U6808 (N_6808,N_6327,N_6138);
and U6809 (N_6809,N_6273,N_6290);
nor U6810 (N_6810,N_6084,N_6439);
xor U6811 (N_6811,N_6177,N_6311);
and U6812 (N_6812,N_6073,N_6214);
nor U6813 (N_6813,N_6166,N_6223);
xnor U6814 (N_6814,N_6321,N_6433);
nor U6815 (N_6815,N_6146,N_6082);
or U6816 (N_6816,N_6076,N_6082);
nor U6817 (N_6817,N_6187,N_6413);
nand U6818 (N_6818,N_6319,N_6444);
nand U6819 (N_6819,N_6280,N_6113);
and U6820 (N_6820,N_6001,N_6261);
nand U6821 (N_6821,N_6449,N_6346);
xor U6822 (N_6822,N_6424,N_6019);
or U6823 (N_6823,N_6050,N_6169);
and U6824 (N_6824,N_6052,N_6284);
and U6825 (N_6825,N_6204,N_6206);
and U6826 (N_6826,N_6375,N_6271);
or U6827 (N_6827,N_6193,N_6322);
nand U6828 (N_6828,N_6268,N_6328);
or U6829 (N_6829,N_6188,N_6050);
xnor U6830 (N_6830,N_6455,N_6314);
xor U6831 (N_6831,N_6436,N_6145);
or U6832 (N_6832,N_6102,N_6061);
nand U6833 (N_6833,N_6184,N_6015);
or U6834 (N_6834,N_6344,N_6213);
or U6835 (N_6835,N_6175,N_6150);
xor U6836 (N_6836,N_6497,N_6211);
nor U6837 (N_6837,N_6185,N_6218);
or U6838 (N_6838,N_6370,N_6379);
nor U6839 (N_6839,N_6263,N_6498);
nor U6840 (N_6840,N_6345,N_6239);
nor U6841 (N_6841,N_6485,N_6278);
nor U6842 (N_6842,N_6246,N_6453);
nand U6843 (N_6843,N_6017,N_6346);
xnor U6844 (N_6844,N_6473,N_6058);
xnor U6845 (N_6845,N_6331,N_6035);
xnor U6846 (N_6846,N_6375,N_6355);
nor U6847 (N_6847,N_6263,N_6485);
and U6848 (N_6848,N_6006,N_6031);
nand U6849 (N_6849,N_6289,N_6083);
nor U6850 (N_6850,N_6242,N_6389);
nand U6851 (N_6851,N_6401,N_6005);
xnor U6852 (N_6852,N_6318,N_6327);
xnor U6853 (N_6853,N_6359,N_6062);
nand U6854 (N_6854,N_6111,N_6171);
xor U6855 (N_6855,N_6296,N_6176);
nand U6856 (N_6856,N_6357,N_6141);
xor U6857 (N_6857,N_6236,N_6047);
xor U6858 (N_6858,N_6363,N_6323);
nand U6859 (N_6859,N_6319,N_6279);
nand U6860 (N_6860,N_6366,N_6136);
and U6861 (N_6861,N_6116,N_6006);
and U6862 (N_6862,N_6204,N_6360);
nand U6863 (N_6863,N_6119,N_6491);
xnor U6864 (N_6864,N_6243,N_6418);
and U6865 (N_6865,N_6176,N_6191);
or U6866 (N_6866,N_6409,N_6376);
nor U6867 (N_6867,N_6331,N_6478);
nor U6868 (N_6868,N_6267,N_6284);
and U6869 (N_6869,N_6458,N_6461);
or U6870 (N_6870,N_6074,N_6369);
and U6871 (N_6871,N_6497,N_6328);
nor U6872 (N_6872,N_6008,N_6235);
nor U6873 (N_6873,N_6066,N_6082);
or U6874 (N_6874,N_6265,N_6416);
xor U6875 (N_6875,N_6452,N_6203);
or U6876 (N_6876,N_6486,N_6033);
nand U6877 (N_6877,N_6290,N_6116);
and U6878 (N_6878,N_6179,N_6194);
xnor U6879 (N_6879,N_6151,N_6087);
xnor U6880 (N_6880,N_6283,N_6320);
and U6881 (N_6881,N_6135,N_6327);
nand U6882 (N_6882,N_6497,N_6182);
and U6883 (N_6883,N_6368,N_6116);
nand U6884 (N_6884,N_6287,N_6044);
nor U6885 (N_6885,N_6038,N_6406);
nor U6886 (N_6886,N_6438,N_6234);
nor U6887 (N_6887,N_6298,N_6397);
nand U6888 (N_6888,N_6183,N_6319);
nor U6889 (N_6889,N_6080,N_6449);
nand U6890 (N_6890,N_6131,N_6339);
and U6891 (N_6891,N_6333,N_6081);
or U6892 (N_6892,N_6183,N_6495);
nand U6893 (N_6893,N_6466,N_6294);
nand U6894 (N_6894,N_6034,N_6130);
or U6895 (N_6895,N_6172,N_6018);
nor U6896 (N_6896,N_6447,N_6174);
xor U6897 (N_6897,N_6223,N_6235);
nand U6898 (N_6898,N_6488,N_6111);
and U6899 (N_6899,N_6353,N_6341);
xnor U6900 (N_6900,N_6039,N_6099);
or U6901 (N_6901,N_6303,N_6460);
or U6902 (N_6902,N_6294,N_6118);
nand U6903 (N_6903,N_6182,N_6106);
xnor U6904 (N_6904,N_6100,N_6189);
xor U6905 (N_6905,N_6420,N_6023);
xor U6906 (N_6906,N_6349,N_6231);
nand U6907 (N_6907,N_6066,N_6474);
xor U6908 (N_6908,N_6177,N_6375);
and U6909 (N_6909,N_6430,N_6171);
or U6910 (N_6910,N_6194,N_6135);
and U6911 (N_6911,N_6349,N_6146);
and U6912 (N_6912,N_6068,N_6001);
nand U6913 (N_6913,N_6136,N_6316);
nor U6914 (N_6914,N_6404,N_6133);
nand U6915 (N_6915,N_6241,N_6377);
nand U6916 (N_6916,N_6016,N_6268);
or U6917 (N_6917,N_6026,N_6081);
nor U6918 (N_6918,N_6029,N_6406);
or U6919 (N_6919,N_6090,N_6266);
or U6920 (N_6920,N_6422,N_6007);
and U6921 (N_6921,N_6448,N_6135);
xor U6922 (N_6922,N_6344,N_6050);
or U6923 (N_6923,N_6390,N_6457);
nor U6924 (N_6924,N_6420,N_6300);
xnor U6925 (N_6925,N_6329,N_6417);
or U6926 (N_6926,N_6090,N_6269);
or U6927 (N_6927,N_6088,N_6096);
nand U6928 (N_6928,N_6150,N_6376);
nor U6929 (N_6929,N_6296,N_6209);
or U6930 (N_6930,N_6477,N_6059);
nor U6931 (N_6931,N_6445,N_6047);
xor U6932 (N_6932,N_6315,N_6189);
nand U6933 (N_6933,N_6402,N_6175);
nand U6934 (N_6934,N_6303,N_6213);
and U6935 (N_6935,N_6114,N_6164);
nand U6936 (N_6936,N_6224,N_6280);
nand U6937 (N_6937,N_6326,N_6442);
nand U6938 (N_6938,N_6259,N_6384);
nand U6939 (N_6939,N_6087,N_6344);
or U6940 (N_6940,N_6023,N_6401);
nor U6941 (N_6941,N_6367,N_6397);
or U6942 (N_6942,N_6247,N_6138);
nand U6943 (N_6943,N_6044,N_6251);
nand U6944 (N_6944,N_6263,N_6115);
xor U6945 (N_6945,N_6072,N_6419);
and U6946 (N_6946,N_6391,N_6121);
or U6947 (N_6947,N_6255,N_6224);
or U6948 (N_6948,N_6007,N_6029);
and U6949 (N_6949,N_6214,N_6302);
or U6950 (N_6950,N_6257,N_6171);
nand U6951 (N_6951,N_6402,N_6489);
and U6952 (N_6952,N_6249,N_6465);
nor U6953 (N_6953,N_6452,N_6314);
xor U6954 (N_6954,N_6162,N_6091);
xor U6955 (N_6955,N_6280,N_6055);
xnor U6956 (N_6956,N_6422,N_6025);
and U6957 (N_6957,N_6072,N_6046);
and U6958 (N_6958,N_6241,N_6134);
nor U6959 (N_6959,N_6321,N_6270);
and U6960 (N_6960,N_6488,N_6082);
nor U6961 (N_6961,N_6298,N_6293);
and U6962 (N_6962,N_6007,N_6318);
xnor U6963 (N_6963,N_6055,N_6376);
xnor U6964 (N_6964,N_6472,N_6241);
xor U6965 (N_6965,N_6005,N_6102);
xnor U6966 (N_6966,N_6372,N_6191);
or U6967 (N_6967,N_6482,N_6464);
and U6968 (N_6968,N_6034,N_6028);
nand U6969 (N_6969,N_6030,N_6188);
or U6970 (N_6970,N_6460,N_6166);
nor U6971 (N_6971,N_6124,N_6323);
xor U6972 (N_6972,N_6419,N_6249);
and U6973 (N_6973,N_6324,N_6346);
nand U6974 (N_6974,N_6146,N_6241);
xnor U6975 (N_6975,N_6401,N_6295);
and U6976 (N_6976,N_6338,N_6286);
xor U6977 (N_6977,N_6389,N_6036);
and U6978 (N_6978,N_6173,N_6011);
or U6979 (N_6979,N_6203,N_6019);
nand U6980 (N_6980,N_6144,N_6455);
and U6981 (N_6981,N_6425,N_6093);
xor U6982 (N_6982,N_6433,N_6242);
and U6983 (N_6983,N_6051,N_6467);
nand U6984 (N_6984,N_6124,N_6469);
nand U6985 (N_6985,N_6090,N_6029);
xor U6986 (N_6986,N_6009,N_6421);
and U6987 (N_6987,N_6343,N_6169);
or U6988 (N_6988,N_6035,N_6455);
xor U6989 (N_6989,N_6044,N_6277);
or U6990 (N_6990,N_6270,N_6380);
or U6991 (N_6991,N_6150,N_6449);
xor U6992 (N_6992,N_6238,N_6348);
nand U6993 (N_6993,N_6390,N_6296);
and U6994 (N_6994,N_6498,N_6047);
and U6995 (N_6995,N_6105,N_6410);
or U6996 (N_6996,N_6465,N_6229);
nand U6997 (N_6997,N_6059,N_6299);
nor U6998 (N_6998,N_6049,N_6150);
or U6999 (N_6999,N_6205,N_6237);
and U7000 (N_7000,N_6737,N_6747);
or U7001 (N_7001,N_6553,N_6781);
nor U7002 (N_7002,N_6964,N_6689);
nand U7003 (N_7003,N_6792,N_6874);
nor U7004 (N_7004,N_6534,N_6790);
or U7005 (N_7005,N_6894,N_6925);
nand U7006 (N_7006,N_6782,N_6521);
xor U7007 (N_7007,N_6639,N_6982);
and U7008 (N_7008,N_6569,N_6941);
xor U7009 (N_7009,N_6641,N_6678);
nand U7010 (N_7010,N_6883,N_6738);
nor U7011 (N_7011,N_6680,N_6997);
nor U7012 (N_7012,N_6511,N_6959);
or U7013 (N_7013,N_6596,N_6991);
nand U7014 (N_7014,N_6652,N_6872);
and U7015 (N_7015,N_6528,N_6613);
or U7016 (N_7016,N_6977,N_6881);
xnor U7017 (N_7017,N_6969,N_6983);
or U7018 (N_7018,N_6556,N_6840);
nor U7019 (N_7019,N_6994,N_6812);
xnor U7020 (N_7020,N_6890,N_6674);
or U7021 (N_7021,N_6708,N_6806);
nand U7022 (N_7022,N_6951,N_6931);
nand U7023 (N_7023,N_6697,N_6956);
nor U7024 (N_7024,N_6974,N_6780);
or U7025 (N_7025,N_6990,N_6645);
nand U7026 (N_7026,N_6939,N_6516);
nand U7027 (N_7027,N_6510,N_6763);
nand U7028 (N_7028,N_6808,N_6861);
nor U7029 (N_7029,N_6813,N_6906);
nor U7030 (N_7030,N_6547,N_6594);
nor U7031 (N_7031,N_6744,N_6887);
nand U7032 (N_7032,N_6519,N_6835);
or U7033 (N_7033,N_6989,N_6533);
nor U7034 (N_7034,N_6745,N_6715);
nand U7035 (N_7035,N_6638,N_6949);
xor U7036 (N_7036,N_6686,N_6650);
xor U7037 (N_7037,N_6651,N_6920);
nand U7038 (N_7038,N_6892,N_6502);
nor U7039 (N_7039,N_6953,N_6635);
nand U7040 (N_7040,N_6724,N_6663);
and U7041 (N_7041,N_6520,N_6914);
xnor U7042 (N_7042,N_6506,N_6625);
or U7043 (N_7043,N_6954,N_6620);
nor U7044 (N_7044,N_6814,N_6713);
xor U7045 (N_7045,N_6750,N_6593);
nor U7046 (N_7046,N_6976,N_6616);
and U7047 (N_7047,N_6661,N_6798);
and U7048 (N_7048,N_6501,N_6891);
nor U7049 (N_7049,N_6859,N_6868);
nor U7050 (N_7050,N_6870,N_6725);
nor U7051 (N_7051,N_6801,N_6618);
nor U7052 (N_7052,N_6564,N_6796);
and U7053 (N_7053,N_6797,N_6692);
nand U7054 (N_7054,N_6847,N_6525);
or U7055 (N_7055,N_6843,N_6934);
or U7056 (N_7056,N_6875,N_6961);
nand U7057 (N_7057,N_6807,N_6764);
nor U7058 (N_7058,N_6673,N_6825);
nand U7059 (N_7059,N_6985,N_6581);
or U7060 (N_7060,N_6529,N_6504);
nor U7061 (N_7061,N_6546,N_6975);
nor U7062 (N_7062,N_6555,N_6841);
nand U7063 (N_7063,N_6821,N_6749);
nor U7064 (N_7064,N_6935,N_6769);
nand U7065 (N_7065,N_6784,N_6646);
nand U7066 (N_7066,N_6754,N_6878);
or U7067 (N_7067,N_6598,N_6545);
and U7068 (N_7068,N_6865,N_6615);
xor U7069 (N_7069,N_6828,N_6921);
or U7070 (N_7070,N_6753,N_6815);
xor U7071 (N_7071,N_6880,N_6681);
and U7072 (N_7072,N_6551,N_6653);
and U7073 (N_7073,N_6644,N_6933);
nor U7074 (N_7074,N_6968,N_6853);
nor U7075 (N_7075,N_6911,N_6623);
nor U7076 (N_7076,N_6743,N_6657);
xnor U7077 (N_7077,N_6714,N_6633);
or U7078 (N_7078,N_6675,N_6901);
nand U7079 (N_7079,N_6770,N_6535);
nor U7080 (N_7080,N_6606,N_6945);
nor U7081 (N_7081,N_6728,N_6688);
xor U7082 (N_7082,N_6845,N_6909);
or U7083 (N_7083,N_6926,N_6761);
nor U7084 (N_7084,N_6919,N_6836);
and U7085 (N_7085,N_6775,N_6559);
and U7086 (N_7086,N_6774,N_6946);
or U7087 (N_7087,N_6647,N_6590);
nor U7088 (N_7088,N_6624,N_6703);
or U7089 (N_7089,N_6550,N_6958);
nor U7090 (N_7090,N_6608,N_6793);
nand U7091 (N_7091,N_6972,N_6928);
or U7092 (N_7092,N_6785,N_6566);
nor U7093 (N_7093,N_6563,N_6805);
and U7094 (N_7094,N_6866,N_6950);
and U7095 (N_7095,N_6871,N_6849);
and U7096 (N_7096,N_6733,N_6943);
nor U7097 (N_7097,N_6922,N_6531);
nand U7098 (N_7098,N_6570,N_6595);
and U7099 (N_7099,N_6822,N_6952);
and U7100 (N_7100,N_6777,N_6588);
nand U7101 (N_7101,N_6587,N_6723);
and U7102 (N_7102,N_6572,N_6690);
and U7103 (N_7103,N_6896,N_6831);
or U7104 (N_7104,N_6607,N_6736);
xor U7105 (N_7105,N_6779,N_6695);
or U7106 (N_7106,N_6834,N_6605);
xnor U7107 (N_7107,N_6666,N_6755);
xor U7108 (N_7108,N_6571,N_6739);
nand U7109 (N_7109,N_6691,N_6766);
nand U7110 (N_7110,N_6705,N_6709);
nor U7111 (N_7111,N_6756,N_6729);
xor U7112 (N_7112,N_6508,N_6548);
or U7113 (N_7113,N_6819,N_6817);
xor U7114 (N_7114,N_6698,N_6893);
xnor U7115 (N_7115,N_6971,N_6643);
xor U7116 (N_7116,N_6706,N_6963);
xnor U7117 (N_7117,N_6947,N_6716);
nor U7118 (N_7118,N_6670,N_6536);
and U7119 (N_7119,N_6583,N_6514);
nor U7120 (N_7120,N_6824,N_6526);
or U7121 (N_7121,N_6966,N_6567);
and U7122 (N_7122,N_6575,N_6957);
nand U7123 (N_7123,N_6850,N_6704);
and U7124 (N_7124,N_6549,N_6827);
and U7125 (N_7125,N_6981,N_6560);
nand U7126 (N_7126,N_6602,N_6562);
or U7127 (N_7127,N_6748,N_6540);
or U7128 (N_7128,N_6539,N_6507);
nand U7129 (N_7129,N_6667,N_6513);
or U7130 (N_7130,N_6803,N_6710);
nand U7131 (N_7131,N_6768,N_6965);
nor U7132 (N_7132,N_6542,N_6721);
xor U7133 (N_7133,N_6752,N_6913);
nor U7134 (N_7134,N_6858,N_6979);
nand U7135 (N_7135,N_6885,N_6636);
or U7136 (N_7136,N_6517,N_6654);
or U7137 (N_7137,N_6573,N_6852);
or U7138 (N_7138,N_6627,N_6735);
or U7139 (N_7139,N_6902,N_6523);
and U7140 (N_7140,N_6897,N_6741);
nor U7141 (N_7141,N_6876,N_6809);
nand U7142 (N_7142,N_6856,N_6684);
xnor U7143 (N_7143,N_6936,N_6787);
and U7144 (N_7144,N_6915,N_6672);
nand U7145 (N_7145,N_6776,N_6869);
xnor U7146 (N_7146,N_6524,N_6772);
nor U7147 (N_7147,N_6973,N_6614);
or U7148 (N_7148,N_6863,N_6918);
nor U7149 (N_7149,N_6585,N_6621);
and U7150 (N_7150,N_6732,N_6862);
nor U7151 (N_7151,N_6599,N_6903);
nand U7152 (N_7152,N_6677,N_6617);
xnor U7153 (N_7153,N_6541,N_6669);
and U7154 (N_7154,N_6992,N_6879);
xor U7155 (N_7155,N_6642,N_6842);
nand U7156 (N_7156,N_6582,N_6799);
nand U7157 (N_7157,N_6898,N_6867);
or U7158 (N_7158,N_6631,N_6632);
xor U7159 (N_7159,N_6771,N_6640);
and U7160 (N_7160,N_6655,N_6942);
or U7161 (N_7161,N_6757,N_6586);
nor U7162 (N_7162,N_6882,N_6844);
or U7163 (N_7163,N_6899,N_6751);
nor U7164 (N_7164,N_6682,N_6589);
nand U7165 (N_7165,N_6719,N_6576);
nand U7166 (N_7166,N_6758,N_6543);
xnor U7167 (N_7167,N_6846,N_6693);
nor U7168 (N_7168,N_6577,N_6888);
or U7169 (N_7169,N_6886,N_6530);
nand U7170 (N_7170,N_6760,N_6718);
or U7171 (N_7171,N_6702,N_6660);
xor U7172 (N_7172,N_6905,N_6722);
nor U7173 (N_7173,N_6938,N_6937);
xor U7174 (N_7174,N_6668,N_6561);
xor U7175 (N_7175,N_6940,N_6515);
nand U7176 (N_7176,N_6610,N_6948);
nor U7177 (N_7177,N_6854,N_6700);
xnor U7178 (N_7178,N_6912,N_6648);
or U7179 (N_7179,N_6707,N_6685);
or U7180 (N_7180,N_6970,N_6823);
or U7181 (N_7181,N_6634,N_6727);
xor U7182 (N_7182,N_6786,N_6699);
and U7183 (N_7183,N_6591,N_6619);
nor U7184 (N_7184,N_6829,N_6838);
nor U7185 (N_7185,N_6765,N_6980);
nand U7186 (N_7186,N_6518,N_6999);
or U7187 (N_7187,N_6503,N_6955);
nor U7188 (N_7188,N_6742,N_6544);
nand U7189 (N_7189,N_6794,N_6960);
and U7190 (N_7190,N_6804,N_6683);
nand U7191 (N_7191,N_6662,N_6537);
xnor U7192 (N_7192,N_6679,N_6726);
or U7193 (N_7193,N_6832,N_6604);
xnor U7194 (N_7194,N_6759,N_6687);
or U7195 (N_7195,N_6851,N_6622);
nand U7196 (N_7196,N_6986,N_6554);
nor U7197 (N_7197,N_6826,N_6565);
nor U7198 (N_7198,N_6578,N_6802);
nor U7199 (N_7199,N_6512,N_6904);
and U7200 (N_7200,N_6712,N_6923);
xor U7201 (N_7201,N_6864,N_6500);
xor U7202 (N_7202,N_6665,N_6731);
or U7203 (N_7203,N_6839,N_6944);
xnor U7204 (N_7204,N_6538,N_6580);
nand U7205 (N_7205,N_6696,N_6649);
nor U7206 (N_7206,N_6527,N_6609);
or U7207 (N_7207,N_6637,N_6818);
and U7208 (N_7208,N_6995,N_6584);
nand U7209 (N_7209,N_6717,N_6579);
or U7210 (N_7210,N_6910,N_6916);
nand U7211 (N_7211,N_6597,N_6962);
nor U7212 (N_7212,N_6773,N_6532);
and U7213 (N_7213,N_6855,N_6626);
or U7214 (N_7214,N_6929,N_6833);
xnor U7215 (N_7215,N_6557,N_6720);
nand U7216 (N_7216,N_6701,N_6600);
nor U7217 (N_7217,N_6789,N_6746);
or U7218 (N_7218,N_6884,N_6998);
or U7219 (N_7219,N_6917,N_6522);
nor U7220 (N_7220,N_6612,N_6628);
xor U7221 (N_7221,N_6788,N_6800);
nand U7222 (N_7222,N_6810,N_6791);
nor U7223 (N_7223,N_6592,N_6907);
nand U7224 (N_7224,N_6900,N_6895);
and U7225 (N_7225,N_6795,N_6984);
xor U7226 (N_7226,N_6574,N_6927);
xor U7227 (N_7227,N_6988,N_6932);
xor U7228 (N_7228,N_6816,N_6630);
nor U7229 (N_7229,N_6767,N_6694);
or U7230 (N_7230,N_6908,N_6778);
nor U7231 (N_7231,N_6930,N_6629);
nand U7232 (N_7232,N_6873,N_6711);
nor U7233 (N_7233,N_6671,N_6509);
and U7234 (N_7234,N_6664,N_6603);
and U7235 (N_7235,N_6505,N_6730);
xnor U7236 (N_7236,N_6568,N_6740);
nand U7237 (N_7237,N_6656,N_6857);
nor U7238 (N_7238,N_6967,N_6811);
nand U7239 (N_7239,N_6762,N_6611);
or U7240 (N_7240,N_6552,N_6783);
or U7241 (N_7241,N_6734,N_6658);
and U7242 (N_7242,N_6978,N_6924);
xor U7243 (N_7243,N_6676,N_6987);
and U7244 (N_7244,N_6889,N_6601);
nand U7245 (N_7245,N_6877,N_6837);
nor U7246 (N_7246,N_6993,N_6848);
nor U7247 (N_7247,N_6860,N_6659);
or U7248 (N_7248,N_6830,N_6820);
and U7249 (N_7249,N_6996,N_6558);
nor U7250 (N_7250,N_6532,N_6910);
or U7251 (N_7251,N_6992,N_6829);
and U7252 (N_7252,N_6998,N_6532);
or U7253 (N_7253,N_6687,N_6637);
and U7254 (N_7254,N_6955,N_6721);
or U7255 (N_7255,N_6841,N_6701);
xnor U7256 (N_7256,N_6946,N_6735);
xor U7257 (N_7257,N_6707,N_6538);
xor U7258 (N_7258,N_6846,N_6776);
nor U7259 (N_7259,N_6829,N_6984);
xnor U7260 (N_7260,N_6566,N_6915);
nor U7261 (N_7261,N_6736,N_6714);
or U7262 (N_7262,N_6684,N_6988);
nor U7263 (N_7263,N_6855,N_6704);
nand U7264 (N_7264,N_6804,N_6851);
xor U7265 (N_7265,N_6698,N_6960);
and U7266 (N_7266,N_6670,N_6615);
or U7267 (N_7267,N_6935,N_6746);
or U7268 (N_7268,N_6555,N_6643);
nand U7269 (N_7269,N_6933,N_6521);
nor U7270 (N_7270,N_6950,N_6574);
xnor U7271 (N_7271,N_6941,N_6607);
and U7272 (N_7272,N_6883,N_6838);
nand U7273 (N_7273,N_6716,N_6585);
or U7274 (N_7274,N_6799,N_6858);
nand U7275 (N_7275,N_6511,N_6980);
nor U7276 (N_7276,N_6804,N_6515);
and U7277 (N_7277,N_6656,N_6884);
xnor U7278 (N_7278,N_6572,N_6576);
nor U7279 (N_7279,N_6720,N_6990);
or U7280 (N_7280,N_6542,N_6705);
and U7281 (N_7281,N_6753,N_6527);
xor U7282 (N_7282,N_6851,N_6712);
or U7283 (N_7283,N_6924,N_6800);
or U7284 (N_7284,N_6646,N_6973);
and U7285 (N_7285,N_6577,N_6781);
or U7286 (N_7286,N_6619,N_6531);
or U7287 (N_7287,N_6831,N_6699);
or U7288 (N_7288,N_6762,N_6721);
xor U7289 (N_7289,N_6621,N_6701);
nor U7290 (N_7290,N_6703,N_6843);
xor U7291 (N_7291,N_6788,N_6723);
and U7292 (N_7292,N_6626,N_6691);
nor U7293 (N_7293,N_6631,N_6667);
and U7294 (N_7294,N_6839,N_6893);
xnor U7295 (N_7295,N_6878,N_6683);
xor U7296 (N_7296,N_6919,N_6780);
and U7297 (N_7297,N_6824,N_6893);
and U7298 (N_7298,N_6858,N_6870);
xor U7299 (N_7299,N_6935,N_6698);
nor U7300 (N_7300,N_6821,N_6985);
or U7301 (N_7301,N_6696,N_6773);
or U7302 (N_7302,N_6797,N_6815);
or U7303 (N_7303,N_6938,N_6785);
and U7304 (N_7304,N_6684,N_6662);
nor U7305 (N_7305,N_6661,N_6895);
and U7306 (N_7306,N_6812,N_6976);
or U7307 (N_7307,N_6614,N_6938);
and U7308 (N_7308,N_6862,N_6520);
xor U7309 (N_7309,N_6726,N_6561);
xor U7310 (N_7310,N_6827,N_6731);
nand U7311 (N_7311,N_6893,N_6933);
nand U7312 (N_7312,N_6793,N_6683);
nor U7313 (N_7313,N_6568,N_6781);
nand U7314 (N_7314,N_6718,N_6528);
and U7315 (N_7315,N_6991,N_6543);
nor U7316 (N_7316,N_6799,N_6840);
or U7317 (N_7317,N_6913,N_6742);
nand U7318 (N_7318,N_6756,N_6693);
nor U7319 (N_7319,N_6563,N_6542);
and U7320 (N_7320,N_6891,N_6777);
xnor U7321 (N_7321,N_6866,N_6615);
xor U7322 (N_7322,N_6848,N_6973);
or U7323 (N_7323,N_6601,N_6731);
nor U7324 (N_7324,N_6911,N_6781);
and U7325 (N_7325,N_6780,N_6928);
or U7326 (N_7326,N_6556,N_6584);
or U7327 (N_7327,N_6964,N_6790);
and U7328 (N_7328,N_6563,N_6703);
nand U7329 (N_7329,N_6761,N_6666);
nor U7330 (N_7330,N_6827,N_6824);
nand U7331 (N_7331,N_6594,N_6952);
xnor U7332 (N_7332,N_6656,N_6965);
nand U7333 (N_7333,N_6564,N_6984);
nand U7334 (N_7334,N_6676,N_6544);
and U7335 (N_7335,N_6631,N_6927);
nand U7336 (N_7336,N_6552,N_6727);
nor U7337 (N_7337,N_6613,N_6550);
and U7338 (N_7338,N_6800,N_6762);
and U7339 (N_7339,N_6675,N_6729);
nor U7340 (N_7340,N_6973,N_6917);
nand U7341 (N_7341,N_6799,N_6997);
nor U7342 (N_7342,N_6518,N_6971);
and U7343 (N_7343,N_6723,N_6516);
and U7344 (N_7344,N_6514,N_6885);
nand U7345 (N_7345,N_6876,N_6918);
xor U7346 (N_7346,N_6690,N_6568);
nand U7347 (N_7347,N_6642,N_6580);
nand U7348 (N_7348,N_6843,N_6560);
xor U7349 (N_7349,N_6916,N_6930);
xnor U7350 (N_7350,N_6507,N_6583);
and U7351 (N_7351,N_6966,N_6606);
nand U7352 (N_7352,N_6632,N_6931);
nor U7353 (N_7353,N_6902,N_6966);
xnor U7354 (N_7354,N_6723,N_6639);
nor U7355 (N_7355,N_6656,N_6913);
nor U7356 (N_7356,N_6947,N_6833);
and U7357 (N_7357,N_6901,N_6713);
nor U7358 (N_7358,N_6538,N_6913);
xor U7359 (N_7359,N_6849,N_6878);
or U7360 (N_7360,N_6927,N_6882);
nor U7361 (N_7361,N_6703,N_6817);
and U7362 (N_7362,N_6939,N_6716);
nor U7363 (N_7363,N_6825,N_6748);
xnor U7364 (N_7364,N_6936,N_6731);
nand U7365 (N_7365,N_6798,N_6788);
nor U7366 (N_7366,N_6535,N_6970);
and U7367 (N_7367,N_6579,N_6588);
or U7368 (N_7368,N_6985,N_6702);
or U7369 (N_7369,N_6979,N_6955);
and U7370 (N_7370,N_6575,N_6651);
and U7371 (N_7371,N_6538,N_6803);
nand U7372 (N_7372,N_6930,N_6732);
and U7373 (N_7373,N_6609,N_6629);
nand U7374 (N_7374,N_6837,N_6960);
and U7375 (N_7375,N_6837,N_6932);
xnor U7376 (N_7376,N_6987,N_6709);
and U7377 (N_7377,N_6598,N_6987);
and U7378 (N_7378,N_6820,N_6628);
or U7379 (N_7379,N_6642,N_6581);
nor U7380 (N_7380,N_6729,N_6785);
xor U7381 (N_7381,N_6913,N_6771);
nor U7382 (N_7382,N_6909,N_6563);
nand U7383 (N_7383,N_6586,N_6895);
and U7384 (N_7384,N_6831,N_6815);
or U7385 (N_7385,N_6588,N_6563);
xor U7386 (N_7386,N_6836,N_6605);
nor U7387 (N_7387,N_6679,N_6824);
nor U7388 (N_7388,N_6617,N_6905);
nand U7389 (N_7389,N_6587,N_6986);
nand U7390 (N_7390,N_6562,N_6621);
xnor U7391 (N_7391,N_6872,N_6734);
or U7392 (N_7392,N_6864,N_6784);
or U7393 (N_7393,N_6687,N_6997);
and U7394 (N_7394,N_6872,N_6775);
xnor U7395 (N_7395,N_6818,N_6901);
or U7396 (N_7396,N_6942,N_6829);
xor U7397 (N_7397,N_6836,N_6524);
nor U7398 (N_7398,N_6900,N_6915);
and U7399 (N_7399,N_6661,N_6530);
xor U7400 (N_7400,N_6512,N_6877);
nor U7401 (N_7401,N_6515,N_6926);
nand U7402 (N_7402,N_6780,N_6940);
and U7403 (N_7403,N_6962,N_6833);
nand U7404 (N_7404,N_6728,N_6950);
nor U7405 (N_7405,N_6913,N_6559);
xnor U7406 (N_7406,N_6660,N_6882);
nand U7407 (N_7407,N_6875,N_6864);
nand U7408 (N_7408,N_6562,N_6811);
and U7409 (N_7409,N_6567,N_6994);
xor U7410 (N_7410,N_6570,N_6543);
and U7411 (N_7411,N_6790,N_6945);
xnor U7412 (N_7412,N_6591,N_6969);
xnor U7413 (N_7413,N_6510,N_6801);
nor U7414 (N_7414,N_6627,N_6536);
xor U7415 (N_7415,N_6607,N_6899);
nand U7416 (N_7416,N_6686,N_6794);
xor U7417 (N_7417,N_6589,N_6526);
nand U7418 (N_7418,N_6652,N_6506);
nor U7419 (N_7419,N_6729,N_6501);
nand U7420 (N_7420,N_6873,N_6767);
or U7421 (N_7421,N_6675,N_6513);
nor U7422 (N_7422,N_6847,N_6973);
nand U7423 (N_7423,N_6651,N_6675);
xor U7424 (N_7424,N_6705,N_6771);
and U7425 (N_7425,N_6506,N_6872);
nor U7426 (N_7426,N_6779,N_6560);
or U7427 (N_7427,N_6757,N_6566);
or U7428 (N_7428,N_6541,N_6654);
nand U7429 (N_7429,N_6777,N_6606);
or U7430 (N_7430,N_6835,N_6576);
nor U7431 (N_7431,N_6942,N_6673);
nand U7432 (N_7432,N_6686,N_6944);
and U7433 (N_7433,N_6712,N_6718);
nor U7434 (N_7434,N_6701,N_6786);
or U7435 (N_7435,N_6573,N_6551);
or U7436 (N_7436,N_6555,N_6684);
xnor U7437 (N_7437,N_6519,N_6500);
and U7438 (N_7438,N_6763,N_6554);
xnor U7439 (N_7439,N_6573,N_6641);
nor U7440 (N_7440,N_6857,N_6718);
nor U7441 (N_7441,N_6536,N_6692);
nor U7442 (N_7442,N_6619,N_6908);
xor U7443 (N_7443,N_6654,N_6683);
or U7444 (N_7444,N_6765,N_6609);
or U7445 (N_7445,N_6583,N_6888);
and U7446 (N_7446,N_6763,N_6758);
nand U7447 (N_7447,N_6547,N_6855);
or U7448 (N_7448,N_6923,N_6845);
nand U7449 (N_7449,N_6851,N_6834);
nor U7450 (N_7450,N_6737,N_6798);
nor U7451 (N_7451,N_6591,N_6661);
nor U7452 (N_7452,N_6823,N_6812);
and U7453 (N_7453,N_6679,N_6689);
nor U7454 (N_7454,N_6928,N_6946);
or U7455 (N_7455,N_6642,N_6967);
xor U7456 (N_7456,N_6663,N_6533);
and U7457 (N_7457,N_6630,N_6729);
or U7458 (N_7458,N_6851,N_6545);
and U7459 (N_7459,N_6741,N_6830);
xor U7460 (N_7460,N_6820,N_6521);
and U7461 (N_7461,N_6696,N_6644);
nand U7462 (N_7462,N_6673,N_6990);
nor U7463 (N_7463,N_6982,N_6515);
and U7464 (N_7464,N_6949,N_6805);
or U7465 (N_7465,N_6798,N_6656);
nand U7466 (N_7466,N_6745,N_6909);
or U7467 (N_7467,N_6512,N_6952);
and U7468 (N_7468,N_6709,N_6833);
and U7469 (N_7469,N_6515,N_6901);
or U7470 (N_7470,N_6602,N_6681);
nand U7471 (N_7471,N_6552,N_6617);
nor U7472 (N_7472,N_6860,N_6644);
and U7473 (N_7473,N_6577,N_6506);
nor U7474 (N_7474,N_6523,N_6934);
xnor U7475 (N_7475,N_6894,N_6578);
or U7476 (N_7476,N_6606,N_6882);
and U7477 (N_7477,N_6527,N_6654);
nor U7478 (N_7478,N_6750,N_6572);
or U7479 (N_7479,N_6984,N_6949);
xnor U7480 (N_7480,N_6852,N_6533);
and U7481 (N_7481,N_6929,N_6625);
or U7482 (N_7482,N_6951,N_6865);
xnor U7483 (N_7483,N_6962,N_6678);
nor U7484 (N_7484,N_6945,N_6652);
or U7485 (N_7485,N_6672,N_6661);
nand U7486 (N_7486,N_6605,N_6844);
xnor U7487 (N_7487,N_6983,N_6920);
nor U7488 (N_7488,N_6959,N_6579);
or U7489 (N_7489,N_6576,N_6905);
nand U7490 (N_7490,N_6752,N_6821);
nor U7491 (N_7491,N_6814,N_6897);
and U7492 (N_7492,N_6616,N_6706);
nor U7493 (N_7493,N_6772,N_6732);
and U7494 (N_7494,N_6854,N_6510);
xnor U7495 (N_7495,N_6837,N_6586);
xor U7496 (N_7496,N_6838,N_6810);
nor U7497 (N_7497,N_6847,N_6763);
or U7498 (N_7498,N_6752,N_6517);
nand U7499 (N_7499,N_6819,N_6637);
nor U7500 (N_7500,N_7174,N_7324);
xnor U7501 (N_7501,N_7131,N_7411);
nand U7502 (N_7502,N_7102,N_7307);
xor U7503 (N_7503,N_7068,N_7031);
xnor U7504 (N_7504,N_7367,N_7327);
xnor U7505 (N_7505,N_7357,N_7227);
nor U7506 (N_7506,N_7389,N_7302);
nand U7507 (N_7507,N_7257,N_7139);
nor U7508 (N_7508,N_7026,N_7467);
nand U7509 (N_7509,N_7124,N_7234);
nand U7510 (N_7510,N_7188,N_7310);
or U7511 (N_7511,N_7431,N_7228);
nand U7512 (N_7512,N_7496,N_7086);
xnor U7513 (N_7513,N_7195,N_7469);
xnor U7514 (N_7514,N_7413,N_7323);
xnor U7515 (N_7515,N_7082,N_7128);
nor U7516 (N_7516,N_7450,N_7463);
xnor U7517 (N_7517,N_7064,N_7447);
and U7518 (N_7518,N_7027,N_7080);
and U7519 (N_7519,N_7308,N_7244);
nand U7520 (N_7520,N_7189,N_7043);
or U7521 (N_7521,N_7300,N_7474);
or U7522 (N_7522,N_7329,N_7415);
nand U7523 (N_7523,N_7019,N_7083);
nand U7524 (N_7524,N_7059,N_7309);
or U7525 (N_7525,N_7279,N_7408);
and U7526 (N_7526,N_7473,N_7073);
and U7527 (N_7527,N_7110,N_7380);
nand U7528 (N_7528,N_7140,N_7490);
or U7529 (N_7529,N_7097,N_7481);
or U7530 (N_7530,N_7299,N_7079);
nor U7531 (N_7531,N_7109,N_7401);
xor U7532 (N_7532,N_7283,N_7185);
xnor U7533 (N_7533,N_7253,N_7468);
or U7534 (N_7534,N_7479,N_7211);
and U7535 (N_7535,N_7275,N_7282);
or U7536 (N_7536,N_7480,N_7176);
nand U7537 (N_7537,N_7397,N_7364);
nand U7538 (N_7538,N_7280,N_7391);
nor U7539 (N_7539,N_7210,N_7049);
xnor U7540 (N_7540,N_7246,N_7351);
nand U7541 (N_7541,N_7296,N_7233);
nand U7542 (N_7542,N_7156,N_7138);
nor U7543 (N_7543,N_7243,N_7444);
nor U7544 (N_7544,N_7038,N_7338);
nor U7545 (N_7545,N_7004,N_7151);
or U7546 (N_7546,N_7165,N_7432);
or U7547 (N_7547,N_7184,N_7120);
nand U7548 (N_7548,N_7428,N_7331);
or U7549 (N_7549,N_7122,N_7266);
nor U7550 (N_7550,N_7149,N_7426);
nor U7551 (N_7551,N_7350,N_7457);
nor U7552 (N_7552,N_7093,N_7088);
or U7553 (N_7553,N_7263,N_7284);
xnor U7554 (N_7554,N_7335,N_7084);
nor U7555 (N_7555,N_7333,N_7392);
nand U7556 (N_7556,N_7325,N_7262);
and U7557 (N_7557,N_7123,N_7191);
nand U7558 (N_7558,N_7424,N_7314);
xor U7559 (N_7559,N_7106,N_7281);
or U7560 (N_7560,N_7409,N_7154);
and U7561 (N_7561,N_7090,N_7342);
or U7562 (N_7562,N_7236,N_7256);
xnor U7563 (N_7563,N_7039,N_7204);
xnor U7564 (N_7564,N_7250,N_7194);
nand U7565 (N_7565,N_7462,N_7241);
xor U7566 (N_7566,N_7277,N_7180);
nor U7567 (N_7567,N_7359,N_7247);
and U7568 (N_7568,N_7404,N_7321);
xnor U7569 (N_7569,N_7037,N_7183);
nand U7570 (N_7570,N_7453,N_7157);
xnor U7571 (N_7571,N_7330,N_7438);
nand U7572 (N_7572,N_7293,N_7044);
or U7573 (N_7573,N_7024,N_7416);
xnor U7574 (N_7574,N_7425,N_7203);
nor U7575 (N_7575,N_7214,N_7197);
nand U7576 (N_7576,N_7472,N_7458);
and U7577 (N_7577,N_7094,N_7100);
or U7578 (N_7578,N_7013,N_7274);
and U7579 (N_7579,N_7287,N_7187);
xor U7580 (N_7580,N_7245,N_7406);
xnor U7581 (N_7581,N_7301,N_7051);
nor U7582 (N_7582,N_7200,N_7028);
and U7583 (N_7583,N_7229,N_7419);
xnor U7584 (N_7584,N_7119,N_7407);
or U7585 (N_7585,N_7476,N_7053);
nand U7586 (N_7586,N_7202,N_7178);
nand U7587 (N_7587,N_7395,N_7213);
nand U7588 (N_7588,N_7379,N_7014);
or U7589 (N_7589,N_7316,N_7441);
nor U7590 (N_7590,N_7252,N_7378);
nand U7591 (N_7591,N_7159,N_7060);
nor U7592 (N_7592,N_7354,N_7251);
or U7593 (N_7593,N_7141,N_7482);
and U7594 (N_7594,N_7226,N_7326);
or U7595 (N_7595,N_7108,N_7368);
or U7596 (N_7596,N_7217,N_7173);
and U7597 (N_7597,N_7341,N_7095);
nand U7598 (N_7598,N_7319,N_7248);
nand U7599 (N_7599,N_7050,N_7315);
xor U7600 (N_7600,N_7096,N_7105);
and U7601 (N_7601,N_7112,N_7345);
nor U7602 (N_7602,N_7448,N_7232);
nand U7603 (N_7603,N_7360,N_7091);
or U7604 (N_7604,N_7132,N_7443);
xor U7605 (N_7605,N_7423,N_7207);
nand U7606 (N_7606,N_7313,N_7040);
or U7607 (N_7607,N_7451,N_7168);
or U7608 (N_7608,N_7058,N_7161);
or U7609 (N_7609,N_7454,N_7172);
nor U7610 (N_7610,N_7117,N_7158);
and U7611 (N_7611,N_7393,N_7466);
nand U7612 (N_7612,N_7491,N_7322);
nor U7613 (N_7613,N_7125,N_7276);
nor U7614 (N_7614,N_7270,N_7373);
nor U7615 (N_7615,N_7362,N_7489);
nand U7616 (N_7616,N_7237,N_7446);
nor U7617 (N_7617,N_7056,N_7355);
xnor U7618 (N_7618,N_7147,N_7460);
nor U7619 (N_7619,N_7025,N_7437);
and U7620 (N_7620,N_7388,N_7212);
xnor U7621 (N_7621,N_7286,N_7418);
and U7622 (N_7622,N_7186,N_7427);
or U7623 (N_7623,N_7487,N_7081);
xnor U7624 (N_7624,N_7118,N_7224);
xor U7625 (N_7625,N_7346,N_7278);
and U7626 (N_7626,N_7259,N_7041);
nor U7627 (N_7627,N_7340,N_7459);
nand U7628 (N_7628,N_7008,N_7255);
nor U7629 (N_7629,N_7494,N_7449);
or U7630 (N_7630,N_7272,N_7107);
or U7631 (N_7631,N_7261,N_7304);
or U7632 (N_7632,N_7209,N_7386);
nand U7633 (N_7633,N_7181,N_7042);
nand U7634 (N_7634,N_7070,N_7442);
nor U7635 (N_7635,N_7126,N_7371);
xnor U7636 (N_7636,N_7052,N_7303);
xor U7637 (N_7637,N_7394,N_7206);
xnor U7638 (N_7638,N_7336,N_7492);
nand U7639 (N_7639,N_7167,N_7020);
nand U7640 (N_7640,N_7223,N_7000);
xnor U7641 (N_7641,N_7493,N_7366);
nand U7642 (N_7642,N_7190,N_7023);
nor U7643 (N_7643,N_7072,N_7320);
nand U7644 (N_7644,N_7115,N_7290);
and U7645 (N_7645,N_7445,N_7047);
nand U7646 (N_7646,N_7375,N_7225);
nand U7647 (N_7647,N_7046,N_7349);
nand U7648 (N_7648,N_7057,N_7018);
xnor U7649 (N_7649,N_7478,N_7221);
xor U7650 (N_7650,N_7376,N_7498);
xnor U7651 (N_7651,N_7436,N_7067);
nor U7652 (N_7652,N_7348,N_7218);
or U7653 (N_7653,N_7182,N_7148);
xor U7654 (N_7654,N_7033,N_7101);
nor U7655 (N_7655,N_7430,N_7129);
nand U7656 (N_7656,N_7077,N_7265);
nor U7657 (N_7657,N_7098,N_7435);
nand U7658 (N_7658,N_7477,N_7001);
and U7659 (N_7659,N_7162,N_7412);
nor U7660 (N_7660,N_7150,N_7153);
nand U7661 (N_7661,N_7127,N_7216);
xnor U7662 (N_7662,N_7170,N_7334);
xnor U7663 (N_7663,N_7240,N_7075);
and U7664 (N_7664,N_7143,N_7420);
xor U7665 (N_7665,N_7422,N_7339);
nand U7666 (N_7666,N_7483,N_7358);
nand U7667 (N_7667,N_7365,N_7017);
or U7668 (N_7668,N_7273,N_7306);
xor U7669 (N_7669,N_7145,N_7269);
nor U7670 (N_7670,N_7405,N_7439);
nor U7671 (N_7671,N_7328,N_7297);
nand U7672 (N_7672,N_7344,N_7005);
xnor U7673 (N_7673,N_7009,N_7074);
xor U7674 (N_7674,N_7231,N_7136);
nor U7675 (N_7675,N_7434,N_7169);
nand U7676 (N_7676,N_7220,N_7470);
or U7677 (N_7677,N_7114,N_7160);
or U7678 (N_7678,N_7011,N_7164);
xor U7679 (N_7679,N_7130,N_7030);
xnor U7680 (N_7680,N_7012,N_7010);
and U7681 (N_7681,N_7363,N_7045);
nor U7682 (N_7682,N_7134,N_7193);
nand U7683 (N_7683,N_7295,N_7343);
nand U7684 (N_7684,N_7163,N_7078);
nand U7685 (N_7685,N_7452,N_7455);
and U7686 (N_7686,N_7374,N_7133);
nor U7687 (N_7687,N_7369,N_7387);
xnor U7688 (N_7688,N_7288,N_7135);
nor U7689 (N_7689,N_7103,N_7337);
xor U7690 (N_7690,N_7015,N_7402);
and U7691 (N_7691,N_7222,N_7264);
nand U7692 (N_7692,N_7456,N_7497);
or U7693 (N_7693,N_7111,N_7034);
and U7694 (N_7694,N_7166,N_7486);
nor U7695 (N_7695,N_7006,N_7016);
xnor U7696 (N_7696,N_7347,N_7032);
and U7697 (N_7697,N_7317,N_7076);
xor U7698 (N_7698,N_7137,N_7219);
and U7699 (N_7699,N_7242,N_7087);
xnor U7700 (N_7700,N_7356,N_7258);
and U7701 (N_7701,N_7179,N_7488);
or U7702 (N_7702,N_7292,N_7298);
and U7703 (N_7703,N_7239,N_7305);
nor U7704 (N_7704,N_7036,N_7440);
nand U7705 (N_7705,N_7069,N_7235);
and U7706 (N_7706,N_7370,N_7155);
xnor U7707 (N_7707,N_7361,N_7289);
and U7708 (N_7708,N_7383,N_7285);
or U7709 (N_7709,N_7113,N_7352);
xnor U7710 (N_7710,N_7116,N_7238);
nor U7711 (N_7711,N_7205,N_7152);
and U7712 (N_7712,N_7433,N_7065);
xor U7713 (N_7713,N_7267,N_7063);
nand U7714 (N_7714,N_7429,N_7485);
or U7715 (N_7715,N_7230,N_7066);
nand U7716 (N_7716,N_7054,N_7071);
xor U7717 (N_7717,N_7002,N_7171);
and U7718 (N_7718,N_7085,N_7092);
or U7719 (N_7719,N_7390,N_7144);
or U7720 (N_7720,N_7385,N_7377);
nor U7721 (N_7721,N_7414,N_7400);
nand U7722 (N_7722,N_7215,N_7099);
nor U7723 (N_7723,N_7399,N_7294);
or U7724 (N_7724,N_7410,N_7484);
and U7725 (N_7725,N_7461,N_7196);
xnor U7726 (N_7726,N_7104,N_7121);
or U7727 (N_7727,N_7464,N_7291);
nand U7728 (N_7728,N_7495,N_7146);
nor U7729 (N_7729,N_7035,N_7372);
xor U7730 (N_7730,N_7417,N_7177);
nor U7731 (N_7731,N_7421,N_7142);
nand U7732 (N_7732,N_7007,N_7029);
and U7733 (N_7733,N_7353,N_7260);
nor U7734 (N_7734,N_7398,N_7021);
or U7735 (N_7735,N_7471,N_7318);
nand U7736 (N_7736,N_7249,N_7198);
nor U7737 (N_7737,N_7201,N_7271);
nor U7738 (N_7738,N_7208,N_7089);
and U7739 (N_7739,N_7061,N_7396);
and U7740 (N_7740,N_7499,N_7175);
and U7741 (N_7741,N_7062,N_7332);
or U7742 (N_7742,N_7381,N_7022);
or U7743 (N_7743,N_7311,N_7384);
nand U7744 (N_7744,N_7003,N_7268);
and U7745 (N_7745,N_7048,N_7312);
or U7746 (N_7746,N_7465,N_7192);
xnor U7747 (N_7747,N_7403,N_7254);
or U7748 (N_7748,N_7199,N_7055);
nor U7749 (N_7749,N_7382,N_7475);
and U7750 (N_7750,N_7480,N_7369);
and U7751 (N_7751,N_7170,N_7231);
xor U7752 (N_7752,N_7333,N_7205);
or U7753 (N_7753,N_7325,N_7299);
or U7754 (N_7754,N_7370,N_7467);
nand U7755 (N_7755,N_7388,N_7225);
nand U7756 (N_7756,N_7303,N_7062);
xor U7757 (N_7757,N_7129,N_7328);
nand U7758 (N_7758,N_7272,N_7425);
and U7759 (N_7759,N_7398,N_7142);
xnor U7760 (N_7760,N_7087,N_7360);
xnor U7761 (N_7761,N_7181,N_7294);
xor U7762 (N_7762,N_7289,N_7157);
nor U7763 (N_7763,N_7309,N_7162);
or U7764 (N_7764,N_7406,N_7044);
or U7765 (N_7765,N_7492,N_7495);
or U7766 (N_7766,N_7124,N_7175);
or U7767 (N_7767,N_7494,N_7440);
nor U7768 (N_7768,N_7038,N_7335);
nor U7769 (N_7769,N_7183,N_7369);
xor U7770 (N_7770,N_7434,N_7067);
nand U7771 (N_7771,N_7475,N_7319);
nand U7772 (N_7772,N_7191,N_7444);
or U7773 (N_7773,N_7091,N_7287);
and U7774 (N_7774,N_7387,N_7366);
xnor U7775 (N_7775,N_7257,N_7249);
and U7776 (N_7776,N_7407,N_7301);
nand U7777 (N_7777,N_7000,N_7325);
nor U7778 (N_7778,N_7369,N_7263);
and U7779 (N_7779,N_7168,N_7210);
and U7780 (N_7780,N_7008,N_7411);
nand U7781 (N_7781,N_7245,N_7308);
and U7782 (N_7782,N_7432,N_7147);
nand U7783 (N_7783,N_7357,N_7452);
xor U7784 (N_7784,N_7095,N_7164);
nor U7785 (N_7785,N_7232,N_7440);
and U7786 (N_7786,N_7409,N_7118);
nor U7787 (N_7787,N_7310,N_7268);
nor U7788 (N_7788,N_7482,N_7469);
nor U7789 (N_7789,N_7261,N_7218);
or U7790 (N_7790,N_7454,N_7338);
and U7791 (N_7791,N_7394,N_7154);
xor U7792 (N_7792,N_7038,N_7361);
nor U7793 (N_7793,N_7394,N_7221);
or U7794 (N_7794,N_7424,N_7283);
and U7795 (N_7795,N_7425,N_7239);
nor U7796 (N_7796,N_7211,N_7417);
nor U7797 (N_7797,N_7319,N_7348);
or U7798 (N_7798,N_7393,N_7237);
nor U7799 (N_7799,N_7188,N_7287);
and U7800 (N_7800,N_7413,N_7061);
or U7801 (N_7801,N_7106,N_7309);
xnor U7802 (N_7802,N_7153,N_7268);
and U7803 (N_7803,N_7090,N_7061);
xor U7804 (N_7804,N_7463,N_7137);
nand U7805 (N_7805,N_7212,N_7127);
nor U7806 (N_7806,N_7439,N_7032);
nor U7807 (N_7807,N_7255,N_7481);
nor U7808 (N_7808,N_7083,N_7106);
nor U7809 (N_7809,N_7194,N_7499);
nor U7810 (N_7810,N_7075,N_7148);
xnor U7811 (N_7811,N_7329,N_7197);
xor U7812 (N_7812,N_7238,N_7251);
nand U7813 (N_7813,N_7116,N_7449);
xnor U7814 (N_7814,N_7215,N_7210);
xnor U7815 (N_7815,N_7200,N_7005);
xnor U7816 (N_7816,N_7101,N_7166);
xnor U7817 (N_7817,N_7316,N_7002);
xnor U7818 (N_7818,N_7218,N_7184);
xnor U7819 (N_7819,N_7264,N_7015);
or U7820 (N_7820,N_7262,N_7429);
xnor U7821 (N_7821,N_7089,N_7389);
and U7822 (N_7822,N_7033,N_7234);
and U7823 (N_7823,N_7263,N_7115);
and U7824 (N_7824,N_7460,N_7278);
and U7825 (N_7825,N_7175,N_7028);
nor U7826 (N_7826,N_7306,N_7085);
and U7827 (N_7827,N_7486,N_7305);
or U7828 (N_7828,N_7155,N_7200);
nand U7829 (N_7829,N_7167,N_7030);
xor U7830 (N_7830,N_7247,N_7045);
and U7831 (N_7831,N_7190,N_7314);
or U7832 (N_7832,N_7216,N_7132);
nand U7833 (N_7833,N_7147,N_7385);
and U7834 (N_7834,N_7336,N_7120);
or U7835 (N_7835,N_7452,N_7207);
nor U7836 (N_7836,N_7368,N_7119);
or U7837 (N_7837,N_7125,N_7188);
or U7838 (N_7838,N_7345,N_7215);
nand U7839 (N_7839,N_7126,N_7378);
nand U7840 (N_7840,N_7257,N_7266);
xnor U7841 (N_7841,N_7257,N_7381);
nand U7842 (N_7842,N_7244,N_7213);
or U7843 (N_7843,N_7449,N_7041);
nand U7844 (N_7844,N_7390,N_7496);
nand U7845 (N_7845,N_7263,N_7313);
nor U7846 (N_7846,N_7245,N_7410);
and U7847 (N_7847,N_7259,N_7275);
nor U7848 (N_7848,N_7427,N_7060);
nor U7849 (N_7849,N_7364,N_7248);
nand U7850 (N_7850,N_7057,N_7292);
xnor U7851 (N_7851,N_7314,N_7281);
or U7852 (N_7852,N_7275,N_7123);
xor U7853 (N_7853,N_7141,N_7017);
nand U7854 (N_7854,N_7488,N_7280);
or U7855 (N_7855,N_7337,N_7236);
and U7856 (N_7856,N_7316,N_7310);
or U7857 (N_7857,N_7266,N_7153);
nand U7858 (N_7858,N_7479,N_7436);
nor U7859 (N_7859,N_7453,N_7135);
nor U7860 (N_7860,N_7302,N_7342);
and U7861 (N_7861,N_7229,N_7073);
xor U7862 (N_7862,N_7197,N_7428);
xnor U7863 (N_7863,N_7103,N_7197);
nor U7864 (N_7864,N_7090,N_7477);
and U7865 (N_7865,N_7392,N_7238);
xor U7866 (N_7866,N_7123,N_7339);
and U7867 (N_7867,N_7402,N_7257);
xnor U7868 (N_7868,N_7029,N_7321);
or U7869 (N_7869,N_7213,N_7372);
xnor U7870 (N_7870,N_7441,N_7252);
nor U7871 (N_7871,N_7283,N_7242);
and U7872 (N_7872,N_7128,N_7077);
xor U7873 (N_7873,N_7016,N_7082);
or U7874 (N_7874,N_7493,N_7473);
nor U7875 (N_7875,N_7487,N_7299);
nand U7876 (N_7876,N_7142,N_7188);
nor U7877 (N_7877,N_7429,N_7224);
nor U7878 (N_7878,N_7498,N_7246);
and U7879 (N_7879,N_7174,N_7448);
xnor U7880 (N_7880,N_7156,N_7119);
nand U7881 (N_7881,N_7416,N_7286);
nor U7882 (N_7882,N_7283,N_7304);
xnor U7883 (N_7883,N_7286,N_7094);
nor U7884 (N_7884,N_7287,N_7458);
xor U7885 (N_7885,N_7086,N_7405);
or U7886 (N_7886,N_7463,N_7216);
or U7887 (N_7887,N_7258,N_7251);
and U7888 (N_7888,N_7424,N_7174);
or U7889 (N_7889,N_7461,N_7153);
nor U7890 (N_7890,N_7442,N_7170);
nor U7891 (N_7891,N_7469,N_7398);
nand U7892 (N_7892,N_7285,N_7041);
nor U7893 (N_7893,N_7258,N_7095);
or U7894 (N_7894,N_7188,N_7180);
or U7895 (N_7895,N_7112,N_7396);
xnor U7896 (N_7896,N_7219,N_7025);
nand U7897 (N_7897,N_7220,N_7367);
xor U7898 (N_7898,N_7073,N_7209);
or U7899 (N_7899,N_7312,N_7046);
xnor U7900 (N_7900,N_7281,N_7451);
or U7901 (N_7901,N_7055,N_7343);
and U7902 (N_7902,N_7231,N_7102);
nand U7903 (N_7903,N_7289,N_7253);
or U7904 (N_7904,N_7471,N_7047);
xnor U7905 (N_7905,N_7456,N_7122);
or U7906 (N_7906,N_7281,N_7178);
xor U7907 (N_7907,N_7297,N_7194);
xor U7908 (N_7908,N_7125,N_7399);
and U7909 (N_7909,N_7090,N_7050);
or U7910 (N_7910,N_7129,N_7445);
nand U7911 (N_7911,N_7263,N_7179);
or U7912 (N_7912,N_7366,N_7031);
nand U7913 (N_7913,N_7382,N_7191);
nand U7914 (N_7914,N_7279,N_7191);
nand U7915 (N_7915,N_7340,N_7332);
nor U7916 (N_7916,N_7333,N_7038);
nor U7917 (N_7917,N_7475,N_7401);
or U7918 (N_7918,N_7449,N_7018);
or U7919 (N_7919,N_7420,N_7352);
and U7920 (N_7920,N_7300,N_7421);
and U7921 (N_7921,N_7159,N_7417);
nor U7922 (N_7922,N_7046,N_7141);
and U7923 (N_7923,N_7473,N_7139);
nor U7924 (N_7924,N_7259,N_7231);
xor U7925 (N_7925,N_7192,N_7029);
xnor U7926 (N_7926,N_7446,N_7246);
xnor U7927 (N_7927,N_7239,N_7468);
nand U7928 (N_7928,N_7248,N_7222);
or U7929 (N_7929,N_7394,N_7177);
xnor U7930 (N_7930,N_7369,N_7422);
nand U7931 (N_7931,N_7257,N_7222);
and U7932 (N_7932,N_7265,N_7128);
and U7933 (N_7933,N_7015,N_7190);
nor U7934 (N_7934,N_7446,N_7088);
or U7935 (N_7935,N_7187,N_7214);
and U7936 (N_7936,N_7435,N_7097);
or U7937 (N_7937,N_7281,N_7124);
or U7938 (N_7938,N_7012,N_7211);
nand U7939 (N_7939,N_7340,N_7254);
and U7940 (N_7940,N_7056,N_7357);
nor U7941 (N_7941,N_7456,N_7085);
nand U7942 (N_7942,N_7143,N_7142);
and U7943 (N_7943,N_7023,N_7196);
nor U7944 (N_7944,N_7215,N_7256);
nand U7945 (N_7945,N_7041,N_7314);
and U7946 (N_7946,N_7403,N_7068);
or U7947 (N_7947,N_7363,N_7113);
nand U7948 (N_7948,N_7444,N_7003);
or U7949 (N_7949,N_7272,N_7240);
xor U7950 (N_7950,N_7224,N_7441);
nor U7951 (N_7951,N_7318,N_7266);
nand U7952 (N_7952,N_7115,N_7027);
and U7953 (N_7953,N_7022,N_7400);
nor U7954 (N_7954,N_7182,N_7144);
or U7955 (N_7955,N_7435,N_7301);
xor U7956 (N_7956,N_7427,N_7283);
nand U7957 (N_7957,N_7339,N_7190);
and U7958 (N_7958,N_7155,N_7021);
or U7959 (N_7959,N_7383,N_7448);
xnor U7960 (N_7960,N_7326,N_7194);
nand U7961 (N_7961,N_7397,N_7251);
and U7962 (N_7962,N_7363,N_7054);
or U7963 (N_7963,N_7360,N_7392);
nor U7964 (N_7964,N_7284,N_7175);
nand U7965 (N_7965,N_7225,N_7151);
xor U7966 (N_7966,N_7331,N_7051);
or U7967 (N_7967,N_7235,N_7128);
or U7968 (N_7968,N_7440,N_7077);
and U7969 (N_7969,N_7062,N_7151);
nand U7970 (N_7970,N_7181,N_7050);
and U7971 (N_7971,N_7117,N_7292);
nand U7972 (N_7972,N_7077,N_7245);
nor U7973 (N_7973,N_7053,N_7019);
xor U7974 (N_7974,N_7003,N_7193);
and U7975 (N_7975,N_7198,N_7475);
or U7976 (N_7976,N_7261,N_7241);
xnor U7977 (N_7977,N_7152,N_7302);
nand U7978 (N_7978,N_7236,N_7494);
nor U7979 (N_7979,N_7411,N_7087);
or U7980 (N_7980,N_7479,N_7269);
xor U7981 (N_7981,N_7377,N_7105);
and U7982 (N_7982,N_7086,N_7054);
xnor U7983 (N_7983,N_7096,N_7081);
xor U7984 (N_7984,N_7089,N_7293);
or U7985 (N_7985,N_7154,N_7346);
or U7986 (N_7986,N_7467,N_7258);
and U7987 (N_7987,N_7102,N_7222);
or U7988 (N_7988,N_7253,N_7089);
and U7989 (N_7989,N_7118,N_7236);
or U7990 (N_7990,N_7136,N_7365);
nand U7991 (N_7991,N_7489,N_7099);
or U7992 (N_7992,N_7025,N_7334);
nand U7993 (N_7993,N_7338,N_7209);
nand U7994 (N_7994,N_7261,N_7008);
and U7995 (N_7995,N_7026,N_7148);
or U7996 (N_7996,N_7438,N_7061);
nor U7997 (N_7997,N_7009,N_7240);
or U7998 (N_7998,N_7341,N_7471);
or U7999 (N_7999,N_7246,N_7363);
or U8000 (N_8000,N_7751,N_7542);
and U8001 (N_8001,N_7870,N_7895);
or U8002 (N_8002,N_7748,N_7889);
nor U8003 (N_8003,N_7684,N_7908);
nand U8004 (N_8004,N_7814,N_7567);
and U8005 (N_8005,N_7711,N_7916);
and U8006 (N_8006,N_7672,N_7742);
and U8007 (N_8007,N_7901,N_7918);
or U8008 (N_8008,N_7877,N_7668);
xor U8009 (N_8009,N_7595,N_7647);
or U8010 (N_8010,N_7949,N_7944);
or U8011 (N_8011,N_7630,N_7846);
or U8012 (N_8012,N_7864,N_7701);
nor U8013 (N_8013,N_7927,N_7580);
nand U8014 (N_8014,N_7521,N_7839);
or U8015 (N_8015,N_7764,N_7696);
nor U8016 (N_8016,N_7854,N_7692);
nor U8017 (N_8017,N_7719,N_7603);
and U8018 (N_8018,N_7900,N_7859);
and U8019 (N_8019,N_7744,N_7606);
or U8020 (N_8020,N_7938,N_7737);
and U8021 (N_8021,N_7828,N_7669);
xor U8022 (N_8022,N_7851,N_7589);
and U8023 (N_8023,N_7991,N_7952);
nand U8024 (N_8024,N_7602,N_7718);
nor U8025 (N_8025,N_7934,N_7945);
nand U8026 (N_8026,N_7735,N_7967);
nor U8027 (N_8027,N_7882,N_7765);
and U8028 (N_8028,N_7906,N_7811);
nor U8029 (N_8029,N_7679,N_7646);
nor U8030 (N_8030,N_7999,N_7734);
or U8031 (N_8031,N_7946,N_7831);
nor U8032 (N_8032,N_7809,N_7709);
or U8033 (N_8033,N_7667,N_7503);
xor U8034 (N_8034,N_7577,N_7691);
nand U8035 (N_8035,N_7573,N_7540);
or U8036 (N_8036,N_7535,N_7849);
nand U8037 (N_8037,N_7759,N_7773);
or U8038 (N_8038,N_7836,N_7555);
nor U8039 (N_8039,N_7896,N_7827);
or U8040 (N_8040,N_7779,N_7749);
xnor U8041 (N_8041,N_7951,N_7825);
xor U8042 (N_8042,N_7775,N_7845);
and U8043 (N_8043,N_7997,N_7625);
or U8044 (N_8044,N_7605,N_7898);
xor U8045 (N_8045,N_7887,N_7880);
nand U8046 (N_8046,N_7941,N_7541);
or U8047 (N_8047,N_7850,N_7995);
and U8048 (N_8048,N_7597,N_7826);
xor U8049 (N_8049,N_7863,N_7641);
nor U8050 (N_8050,N_7879,N_7914);
or U8051 (N_8051,N_7682,N_7717);
nand U8052 (N_8052,N_7788,N_7614);
or U8053 (N_8053,N_7958,N_7659);
or U8054 (N_8054,N_7925,N_7917);
or U8055 (N_8055,N_7816,N_7835);
xor U8056 (N_8056,N_7922,N_7984);
and U8057 (N_8057,N_7693,N_7968);
xor U8058 (N_8058,N_7664,N_7907);
nand U8059 (N_8059,N_7897,N_7969);
or U8060 (N_8060,N_7937,N_7506);
xnor U8061 (N_8061,N_7558,N_7818);
nor U8062 (N_8062,N_7593,N_7830);
nor U8063 (N_8063,N_7913,N_7725);
nor U8064 (N_8064,N_7700,N_7634);
or U8065 (N_8065,N_7753,N_7862);
and U8066 (N_8066,N_7578,N_7566);
and U8067 (N_8067,N_7635,N_7987);
nand U8068 (N_8068,N_7621,N_7784);
xnor U8069 (N_8069,N_7572,N_7754);
xor U8070 (N_8070,N_7674,N_7729);
xor U8071 (N_8071,N_7727,N_7758);
and U8072 (N_8072,N_7965,N_7515);
xnor U8073 (N_8073,N_7675,N_7961);
or U8074 (N_8074,N_7955,N_7721);
xor U8075 (N_8075,N_7800,N_7723);
nand U8076 (N_8076,N_7990,N_7837);
xnor U8077 (N_8077,N_7716,N_7663);
or U8078 (N_8078,N_7732,N_7988);
nand U8079 (N_8079,N_7881,N_7770);
xnor U8080 (N_8080,N_7998,N_7601);
nor U8081 (N_8081,N_7598,N_7776);
nor U8082 (N_8082,N_7591,N_7645);
or U8083 (N_8083,N_7553,N_7867);
and U8084 (N_8084,N_7752,N_7611);
and U8085 (N_8085,N_7575,N_7694);
or U8086 (N_8086,N_7584,N_7661);
or U8087 (N_8087,N_7795,N_7713);
or U8088 (N_8088,N_7974,N_7912);
or U8089 (N_8089,N_7791,N_7655);
nor U8090 (N_8090,N_7824,N_7511);
and U8091 (N_8091,N_7627,N_7648);
or U8092 (N_8092,N_7690,N_7981);
nand U8093 (N_8093,N_7763,N_7571);
nand U8094 (N_8094,N_7929,N_7983);
or U8095 (N_8095,N_7893,N_7801);
xnor U8096 (N_8096,N_7528,N_7670);
or U8097 (N_8097,N_7815,N_7502);
or U8098 (N_8098,N_7842,N_7857);
nor U8099 (N_8099,N_7799,N_7794);
and U8100 (N_8100,N_7689,N_7569);
and U8101 (N_8101,N_7631,N_7736);
and U8102 (N_8102,N_7852,N_7620);
and U8103 (N_8103,N_7531,N_7676);
nand U8104 (N_8104,N_7564,N_7552);
xnor U8105 (N_8105,N_7878,N_7899);
xor U8106 (N_8106,N_7747,N_7960);
nor U8107 (N_8107,N_7891,N_7774);
or U8108 (N_8108,N_7804,N_7964);
nor U8109 (N_8109,N_7819,N_7726);
nand U8110 (N_8110,N_7890,N_7714);
or U8111 (N_8111,N_7756,N_7802);
nor U8112 (N_8112,N_7996,N_7728);
nand U8113 (N_8113,N_7833,N_7532);
nand U8114 (N_8114,N_7640,N_7978);
or U8115 (N_8115,N_7894,N_7868);
or U8116 (N_8116,N_7649,N_7563);
or U8117 (N_8117,N_7657,N_7834);
and U8118 (N_8118,N_7582,N_7508);
nand U8119 (N_8119,N_7847,N_7789);
xor U8120 (N_8120,N_7778,N_7673);
xor U8121 (N_8121,N_7545,N_7841);
and U8122 (N_8122,N_7704,N_7588);
or U8123 (N_8123,N_7660,N_7554);
nor U8124 (N_8124,N_7524,N_7685);
and U8125 (N_8125,N_7607,N_7688);
nor U8126 (N_8126,N_7931,N_7810);
xnor U8127 (N_8127,N_7514,N_7579);
and U8128 (N_8128,N_7643,N_7757);
nor U8129 (N_8129,N_7613,N_7807);
or U8130 (N_8130,N_7618,N_7838);
or U8131 (N_8131,N_7534,N_7708);
and U8132 (N_8132,N_7808,N_7947);
xor U8133 (N_8133,N_7680,N_7817);
xnor U8134 (N_8134,N_7972,N_7509);
nand U8135 (N_8135,N_7512,N_7982);
xor U8136 (N_8136,N_7755,N_7740);
or U8137 (N_8137,N_7823,N_7651);
xor U8138 (N_8138,N_7548,N_7963);
xnor U8139 (N_8139,N_7518,N_7743);
and U8140 (N_8140,N_7932,N_7662);
and U8141 (N_8141,N_7962,N_7604);
nor U8142 (N_8142,N_7581,N_7544);
xnor U8143 (N_8143,N_7761,N_7724);
or U8144 (N_8144,N_7550,N_7892);
xnor U8145 (N_8145,N_7562,N_7950);
or U8146 (N_8146,N_7869,N_7608);
or U8147 (N_8147,N_7762,N_7678);
xnor U8148 (N_8148,N_7596,N_7919);
and U8149 (N_8149,N_7574,N_7903);
nor U8150 (N_8150,N_7533,N_7970);
nor U8151 (N_8151,N_7953,N_7796);
nor U8152 (N_8152,N_7586,N_7905);
nor U8153 (N_8153,N_7538,N_7760);
nand U8154 (N_8154,N_7860,N_7741);
and U8155 (N_8155,N_7650,N_7510);
nor U8156 (N_8156,N_7858,N_7629);
xnor U8157 (N_8157,N_7576,N_7710);
and U8158 (N_8158,N_7520,N_7658);
or U8159 (N_8159,N_7720,N_7599);
and U8160 (N_8160,N_7956,N_7805);
nor U8161 (N_8161,N_7557,N_7695);
xnor U8162 (N_8162,N_7873,N_7654);
and U8163 (N_8163,N_7626,N_7565);
nor U8164 (N_8164,N_7633,N_7653);
and U8165 (N_8165,N_7832,N_7939);
nor U8166 (N_8166,N_7875,N_7786);
and U8167 (N_8167,N_7766,N_7888);
and U8168 (N_8168,N_7876,N_7666);
xnor U8169 (N_8169,N_7942,N_7568);
and U8170 (N_8170,N_7971,N_7624);
nor U8171 (N_8171,N_7855,N_7853);
nand U8172 (N_8172,N_7522,N_7677);
or U8173 (N_8173,N_7517,N_7821);
nor U8174 (N_8174,N_7639,N_7687);
or U8175 (N_8175,N_7902,N_7915);
nor U8176 (N_8176,N_7556,N_7785);
or U8177 (N_8177,N_7780,N_7686);
and U8178 (N_8178,N_7585,N_7943);
or U8179 (N_8179,N_7772,N_7976);
or U8180 (N_8180,N_7872,N_7609);
nand U8181 (N_8181,N_7536,N_7911);
xnor U8182 (N_8182,N_7948,N_7986);
xnor U8183 (N_8183,N_7530,N_7697);
xor U8184 (N_8184,N_7681,N_7745);
nor U8185 (N_8185,N_7928,N_7871);
nand U8186 (N_8186,N_7957,N_7703);
nand U8187 (N_8187,N_7547,N_7782);
nor U8188 (N_8188,N_7707,N_7977);
nor U8189 (N_8189,N_7840,N_7856);
or U8190 (N_8190,N_7638,N_7739);
xor U8191 (N_8191,N_7738,N_7702);
and U8192 (N_8192,N_7781,N_7500);
and U8193 (N_8193,N_7583,N_7886);
and U8194 (N_8194,N_7549,N_7926);
nor U8195 (N_8195,N_7787,N_7592);
xnor U8196 (N_8196,N_7612,N_7623);
nand U8197 (N_8197,N_7993,N_7722);
nand U8198 (N_8198,N_7570,N_7767);
nand U8199 (N_8199,N_7513,N_7940);
xor U8200 (N_8200,N_7806,N_7813);
or U8201 (N_8201,N_7930,N_7798);
or U8202 (N_8202,N_7966,N_7671);
and U8203 (N_8203,N_7731,N_7848);
or U8204 (N_8204,N_7652,N_7989);
xnor U8205 (N_8205,N_7730,N_7610);
nand U8206 (N_8206,N_7587,N_7959);
xor U8207 (N_8207,N_7844,N_7885);
xor U8208 (N_8208,N_7921,N_7560);
nand U8209 (N_8209,N_7622,N_7539);
xnor U8210 (N_8210,N_7519,N_7628);
xor U8211 (N_8211,N_7910,N_7637);
nand U8212 (N_8212,N_7768,N_7769);
nor U8213 (N_8213,N_7642,N_7994);
or U8214 (N_8214,N_7504,N_7559);
xor U8215 (N_8215,N_7636,N_7884);
or U8216 (N_8216,N_7822,N_7883);
nand U8217 (N_8217,N_7683,N_7590);
nor U8218 (N_8218,N_7526,N_7985);
xor U8219 (N_8219,N_7561,N_7803);
nand U8220 (N_8220,N_7861,N_7935);
xor U8221 (N_8221,N_7537,N_7616);
nor U8222 (N_8222,N_7705,N_7656);
nand U8223 (N_8223,N_7516,N_7865);
nand U8224 (N_8224,N_7792,N_7746);
nor U8225 (N_8225,N_7644,N_7594);
and U8226 (N_8226,N_7980,N_7619);
and U8227 (N_8227,N_7924,N_7750);
or U8228 (N_8228,N_7699,N_7501);
xnor U8229 (N_8229,N_7527,N_7505);
and U8230 (N_8230,N_7615,N_7933);
xnor U8231 (N_8231,N_7909,N_7954);
or U8232 (N_8232,N_7507,N_7904);
and U8233 (N_8233,N_7790,N_7829);
nand U8234 (N_8234,N_7992,N_7600);
or U8235 (N_8235,N_7632,N_7923);
nor U8236 (N_8236,N_7529,N_7979);
or U8237 (N_8237,N_7525,N_7920);
or U8238 (N_8238,N_7812,N_7843);
nor U8239 (N_8239,N_7698,N_7771);
nand U8240 (N_8240,N_7936,N_7715);
nor U8241 (N_8241,N_7543,N_7820);
nand U8242 (N_8242,N_7665,N_7733);
xor U8243 (N_8243,N_7797,N_7973);
xnor U8244 (N_8244,N_7866,N_7975);
nand U8245 (N_8245,N_7706,N_7793);
xor U8246 (N_8246,N_7617,N_7523);
and U8247 (N_8247,N_7874,N_7712);
xnor U8248 (N_8248,N_7551,N_7783);
nor U8249 (N_8249,N_7546,N_7777);
and U8250 (N_8250,N_7685,N_7691);
nor U8251 (N_8251,N_7638,N_7970);
nor U8252 (N_8252,N_7661,N_7869);
nor U8253 (N_8253,N_7528,N_7895);
xnor U8254 (N_8254,N_7527,N_7618);
and U8255 (N_8255,N_7942,N_7860);
or U8256 (N_8256,N_7574,N_7523);
nand U8257 (N_8257,N_7814,N_7657);
xnor U8258 (N_8258,N_7639,N_7996);
xnor U8259 (N_8259,N_7804,N_7559);
nor U8260 (N_8260,N_7953,N_7708);
xor U8261 (N_8261,N_7994,N_7870);
and U8262 (N_8262,N_7704,N_7620);
and U8263 (N_8263,N_7509,N_7845);
and U8264 (N_8264,N_7895,N_7644);
and U8265 (N_8265,N_7667,N_7621);
xnor U8266 (N_8266,N_7581,N_7887);
and U8267 (N_8267,N_7804,N_7915);
xor U8268 (N_8268,N_7504,N_7575);
xor U8269 (N_8269,N_7627,N_7644);
nand U8270 (N_8270,N_7683,N_7922);
nor U8271 (N_8271,N_7942,N_7802);
or U8272 (N_8272,N_7549,N_7680);
nand U8273 (N_8273,N_7671,N_7868);
or U8274 (N_8274,N_7696,N_7941);
and U8275 (N_8275,N_7808,N_7806);
nand U8276 (N_8276,N_7712,N_7625);
xor U8277 (N_8277,N_7595,N_7768);
xnor U8278 (N_8278,N_7643,N_7549);
nor U8279 (N_8279,N_7846,N_7873);
nand U8280 (N_8280,N_7569,N_7714);
and U8281 (N_8281,N_7732,N_7716);
or U8282 (N_8282,N_7933,N_7650);
and U8283 (N_8283,N_7861,N_7895);
xor U8284 (N_8284,N_7900,N_7664);
or U8285 (N_8285,N_7735,N_7580);
nor U8286 (N_8286,N_7637,N_7846);
xnor U8287 (N_8287,N_7786,N_7682);
or U8288 (N_8288,N_7689,N_7861);
nor U8289 (N_8289,N_7884,N_7694);
xor U8290 (N_8290,N_7996,N_7787);
xnor U8291 (N_8291,N_7982,N_7717);
and U8292 (N_8292,N_7955,N_7657);
nand U8293 (N_8293,N_7819,N_7716);
nor U8294 (N_8294,N_7745,N_7992);
and U8295 (N_8295,N_7672,N_7822);
nor U8296 (N_8296,N_7890,N_7706);
or U8297 (N_8297,N_7639,N_7817);
nor U8298 (N_8298,N_7705,N_7975);
nor U8299 (N_8299,N_7918,N_7687);
nand U8300 (N_8300,N_7972,N_7758);
xnor U8301 (N_8301,N_7563,N_7745);
xnor U8302 (N_8302,N_7976,N_7857);
nor U8303 (N_8303,N_7924,N_7832);
or U8304 (N_8304,N_7752,N_7988);
or U8305 (N_8305,N_7654,N_7724);
nand U8306 (N_8306,N_7717,N_7738);
nand U8307 (N_8307,N_7660,N_7670);
or U8308 (N_8308,N_7793,N_7805);
xor U8309 (N_8309,N_7528,N_7745);
nor U8310 (N_8310,N_7670,N_7574);
or U8311 (N_8311,N_7604,N_7643);
and U8312 (N_8312,N_7891,N_7643);
xor U8313 (N_8313,N_7759,N_7839);
xor U8314 (N_8314,N_7612,N_7992);
or U8315 (N_8315,N_7765,N_7803);
xor U8316 (N_8316,N_7843,N_7907);
nor U8317 (N_8317,N_7654,N_7867);
xnor U8318 (N_8318,N_7550,N_7856);
nor U8319 (N_8319,N_7647,N_7766);
and U8320 (N_8320,N_7966,N_7544);
or U8321 (N_8321,N_7810,N_7847);
or U8322 (N_8322,N_7933,N_7807);
and U8323 (N_8323,N_7928,N_7712);
or U8324 (N_8324,N_7666,N_7624);
or U8325 (N_8325,N_7768,N_7866);
nor U8326 (N_8326,N_7861,N_7894);
nor U8327 (N_8327,N_7578,N_7851);
or U8328 (N_8328,N_7978,N_7902);
xor U8329 (N_8329,N_7936,N_7535);
xor U8330 (N_8330,N_7722,N_7639);
nand U8331 (N_8331,N_7649,N_7503);
nor U8332 (N_8332,N_7965,N_7572);
xnor U8333 (N_8333,N_7638,N_7987);
and U8334 (N_8334,N_7668,N_7926);
xor U8335 (N_8335,N_7731,N_7645);
or U8336 (N_8336,N_7768,N_7814);
xnor U8337 (N_8337,N_7748,N_7743);
or U8338 (N_8338,N_7751,N_7548);
xnor U8339 (N_8339,N_7896,N_7892);
or U8340 (N_8340,N_7754,N_7947);
nor U8341 (N_8341,N_7967,N_7900);
or U8342 (N_8342,N_7797,N_7578);
nor U8343 (N_8343,N_7612,N_7901);
and U8344 (N_8344,N_7819,N_7526);
xor U8345 (N_8345,N_7663,N_7904);
xnor U8346 (N_8346,N_7830,N_7661);
nor U8347 (N_8347,N_7865,N_7639);
or U8348 (N_8348,N_7731,N_7568);
xnor U8349 (N_8349,N_7779,N_7953);
nor U8350 (N_8350,N_7503,N_7750);
xnor U8351 (N_8351,N_7771,N_7510);
xnor U8352 (N_8352,N_7943,N_7565);
and U8353 (N_8353,N_7742,N_7971);
nor U8354 (N_8354,N_7686,N_7798);
or U8355 (N_8355,N_7994,N_7892);
xnor U8356 (N_8356,N_7831,N_7695);
nand U8357 (N_8357,N_7979,N_7974);
nand U8358 (N_8358,N_7736,N_7667);
and U8359 (N_8359,N_7920,N_7850);
nor U8360 (N_8360,N_7506,N_7978);
or U8361 (N_8361,N_7633,N_7843);
and U8362 (N_8362,N_7590,N_7707);
nor U8363 (N_8363,N_7666,N_7789);
or U8364 (N_8364,N_7740,N_7700);
xor U8365 (N_8365,N_7562,N_7551);
or U8366 (N_8366,N_7943,N_7909);
or U8367 (N_8367,N_7790,N_7603);
xor U8368 (N_8368,N_7510,N_7890);
and U8369 (N_8369,N_7821,N_7854);
or U8370 (N_8370,N_7604,N_7803);
nor U8371 (N_8371,N_7891,N_7908);
or U8372 (N_8372,N_7935,N_7538);
and U8373 (N_8373,N_7604,N_7947);
or U8374 (N_8374,N_7676,N_7703);
nor U8375 (N_8375,N_7528,N_7971);
or U8376 (N_8376,N_7526,N_7505);
or U8377 (N_8377,N_7788,N_7523);
xor U8378 (N_8378,N_7883,N_7741);
and U8379 (N_8379,N_7645,N_7810);
nand U8380 (N_8380,N_7632,N_7666);
nor U8381 (N_8381,N_7557,N_7615);
nand U8382 (N_8382,N_7647,N_7987);
xnor U8383 (N_8383,N_7668,N_7734);
xnor U8384 (N_8384,N_7899,N_7963);
and U8385 (N_8385,N_7935,N_7697);
or U8386 (N_8386,N_7998,N_7988);
xnor U8387 (N_8387,N_7916,N_7956);
and U8388 (N_8388,N_7886,N_7958);
nor U8389 (N_8389,N_7983,N_7805);
or U8390 (N_8390,N_7863,N_7966);
or U8391 (N_8391,N_7505,N_7890);
nor U8392 (N_8392,N_7729,N_7775);
xor U8393 (N_8393,N_7535,N_7773);
xor U8394 (N_8394,N_7833,N_7715);
xor U8395 (N_8395,N_7545,N_7814);
or U8396 (N_8396,N_7627,N_7750);
nor U8397 (N_8397,N_7574,N_7774);
or U8398 (N_8398,N_7518,N_7702);
nor U8399 (N_8399,N_7589,N_7997);
nor U8400 (N_8400,N_7649,N_7817);
or U8401 (N_8401,N_7507,N_7849);
nand U8402 (N_8402,N_7503,N_7862);
nand U8403 (N_8403,N_7531,N_7606);
xor U8404 (N_8404,N_7528,N_7964);
or U8405 (N_8405,N_7979,N_7853);
xor U8406 (N_8406,N_7801,N_7994);
xnor U8407 (N_8407,N_7721,N_7674);
or U8408 (N_8408,N_7638,N_7835);
nor U8409 (N_8409,N_7849,N_7819);
nor U8410 (N_8410,N_7561,N_7788);
or U8411 (N_8411,N_7816,N_7564);
xnor U8412 (N_8412,N_7931,N_7842);
xnor U8413 (N_8413,N_7825,N_7772);
or U8414 (N_8414,N_7541,N_7698);
nor U8415 (N_8415,N_7725,N_7884);
nor U8416 (N_8416,N_7643,N_7940);
xor U8417 (N_8417,N_7969,N_7884);
nand U8418 (N_8418,N_7737,N_7672);
xor U8419 (N_8419,N_7946,N_7562);
xnor U8420 (N_8420,N_7856,N_7822);
nand U8421 (N_8421,N_7602,N_7819);
and U8422 (N_8422,N_7726,N_7609);
nand U8423 (N_8423,N_7940,N_7834);
or U8424 (N_8424,N_7902,N_7993);
xnor U8425 (N_8425,N_7581,N_7903);
nor U8426 (N_8426,N_7676,N_7791);
xor U8427 (N_8427,N_7576,N_7946);
and U8428 (N_8428,N_7646,N_7667);
nor U8429 (N_8429,N_7585,N_7729);
xnor U8430 (N_8430,N_7652,N_7743);
and U8431 (N_8431,N_7929,N_7937);
or U8432 (N_8432,N_7570,N_7895);
and U8433 (N_8433,N_7875,N_7938);
nor U8434 (N_8434,N_7766,N_7508);
xor U8435 (N_8435,N_7773,N_7874);
nand U8436 (N_8436,N_7925,N_7756);
or U8437 (N_8437,N_7514,N_7706);
nand U8438 (N_8438,N_7886,N_7631);
nand U8439 (N_8439,N_7503,N_7523);
and U8440 (N_8440,N_7816,N_7993);
and U8441 (N_8441,N_7825,N_7846);
nand U8442 (N_8442,N_7997,N_7921);
nor U8443 (N_8443,N_7958,N_7868);
or U8444 (N_8444,N_7584,N_7656);
and U8445 (N_8445,N_7600,N_7638);
nor U8446 (N_8446,N_7873,N_7561);
or U8447 (N_8447,N_7914,N_7651);
nand U8448 (N_8448,N_7875,N_7867);
nor U8449 (N_8449,N_7814,N_7929);
nand U8450 (N_8450,N_7570,N_7530);
and U8451 (N_8451,N_7866,N_7832);
and U8452 (N_8452,N_7879,N_7512);
nand U8453 (N_8453,N_7610,N_7674);
or U8454 (N_8454,N_7999,N_7852);
xnor U8455 (N_8455,N_7807,N_7829);
nor U8456 (N_8456,N_7691,N_7625);
and U8457 (N_8457,N_7918,N_7836);
nor U8458 (N_8458,N_7809,N_7837);
or U8459 (N_8459,N_7757,N_7702);
or U8460 (N_8460,N_7508,N_7932);
nor U8461 (N_8461,N_7764,N_7943);
or U8462 (N_8462,N_7970,N_7607);
nor U8463 (N_8463,N_7724,N_7776);
nor U8464 (N_8464,N_7870,N_7763);
or U8465 (N_8465,N_7777,N_7909);
and U8466 (N_8466,N_7566,N_7512);
or U8467 (N_8467,N_7547,N_7813);
and U8468 (N_8468,N_7954,N_7911);
xnor U8469 (N_8469,N_7799,N_7826);
nor U8470 (N_8470,N_7819,N_7898);
or U8471 (N_8471,N_7644,N_7715);
or U8472 (N_8472,N_7910,N_7734);
nor U8473 (N_8473,N_7990,N_7948);
and U8474 (N_8474,N_7770,N_7877);
nor U8475 (N_8475,N_7957,N_7776);
or U8476 (N_8476,N_7715,N_7548);
xor U8477 (N_8477,N_7539,N_7773);
nor U8478 (N_8478,N_7705,N_7660);
nand U8479 (N_8479,N_7915,N_7633);
or U8480 (N_8480,N_7826,N_7584);
or U8481 (N_8481,N_7866,N_7522);
or U8482 (N_8482,N_7777,N_7522);
nor U8483 (N_8483,N_7692,N_7810);
or U8484 (N_8484,N_7528,N_7501);
nand U8485 (N_8485,N_7679,N_7774);
nor U8486 (N_8486,N_7511,N_7553);
xor U8487 (N_8487,N_7606,N_7622);
nand U8488 (N_8488,N_7783,N_7671);
or U8489 (N_8489,N_7570,N_7705);
nor U8490 (N_8490,N_7668,N_7882);
xnor U8491 (N_8491,N_7834,N_7822);
nand U8492 (N_8492,N_7913,N_7800);
xor U8493 (N_8493,N_7618,N_7871);
nor U8494 (N_8494,N_7984,N_7588);
or U8495 (N_8495,N_7632,N_7784);
xor U8496 (N_8496,N_7750,N_7802);
nor U8497 (N_8497,N_7524,N_7786);
xor U8498 (N_8498,N_7825,N_7676);
xnor U8499 (N_8499,N_7921,N_7840);
or U8500 (N_8500,N_8257,N_8391);
and U8501 (N_8501,N_8221,N_8052);
nor U8502 (N_8502,N_8328,N_8403);
xor U8503 (N_8503,N_8115,N_8423);
xor U8504 (N_8504,N_8459,N_8167);
nand U8505 (N_8505,N_8264,N_8353);
nor U8506 (N_8506,N_8348,N_8412);
or U8507 (N_8507,N_8346,N_8079);
and U8508 (N_8508,N_8213,N_8483);
nor U8509 (N_8509,N_8121,N_8496);
and U8510 (N_8510,N_8226,N_8380);
xor U8511 (N_8511,N_8061,N_8015);
nand U8512 (N_8512,N_8267,N_8057);
xor U8513 (N_8513,N_8302,N_8143);
xor U8514 (N_8514,N_8426,N_8023);
and U8515 (N_8515,N_8244,N_8070);
and U8516 (N_8516,N_8365,N_8261);
nand U8517 (N_8517,N_8487,N_8104);
and U8518 (N_8518,N_8164,N_8235);
xor U8519 (N_8519,N_8214,N_8080);
or U8520 (N_8520,N_8227,N_8435);
and U8521 (N_8521,N_8316,N_8005);
xnor U8522 (N_8522,N_8140,N_8461);
nor U8523 (N_8523,N_8108,N_8427);
xor U8524 (N_8524,N_8107,N_8277);
and U8525 (N_8525,N_8037,N_8351);
nor U8526 (N_8526,N_8374,N_8249);
nor U8527 (N_8527,N_8083,N_8046);
nor U8528 (N_8528,N_8364,N_8418);
and U8529 (N_8529,N_8132,N_8480);
nand U8530 (N_8530,N_8398,N_8479);
nor U8531 (N_8531,N_8066,N_8169);
nand U8532 (N_8532,N_8361,N_8338);
nor U8533 (N_8533,N_8481,N_8147);
and U8534 (N_8534,N_8040,N_8254);
or U8535 (N_8535,N_8295,N_8332);
or U8536 (N_8536,N_8285,N_8102);
nor U8537 (N_8537,N_8417,N_8032);
or U8538 (N_8538,N_8135,N_8002);
nand U8539 (N_8539,N_8125,N_8401);
nand U8540 (N_8540,N_8175,N_8333);
xor U8541 (N_8541,N_8047,N_8034);
nand U8542 (N_8542,N_8149,N_8283);
nand U8543 (N_8543,N_8001,N_8345);
xnor U8544 (N_8544,N_8280,N_8356);
nand U8545 (N_8545,N_8337,N_8242);
or U8546 (N_8546,N_8059,N_8297);
nand U8547 (N_8547,N_8062,N_8373);
nand U8548 (N_8548,N_8237,N_8068);
nor U8549 (N_8549,N_8464,N_8484);
nor U8550 (N_8550,N_8336,N_8263);
xor U8551 (N_8551,N_8449,N_8259);
or U8552 (N_8552,N_8076,N_8072);
xor U8553 (N_8553,N_8156,N_8308);
or U8554 (N_8554,N_8446,N_8362);
or U8555 (N_8555,N_8021,N_8093);
and U8556 (N_8556,N_8182,N_8489);
or U8557 (N_8557,N_8476,N_8067);
and U8558 (N_8558,N_8084,N_8177);
nor U8559 (N_8559,N_8320,N_8019);
or U8560 (N_8560,N_8103,N_8424);
nor U8561 (N_8561,N_8245,N_8395);
nand U8562 (N_8562,N_8016,N_8270);
xor U8563 (N_8563,N_8180,N_8128);
xnor U8564 (N_8564,N_8318,N_8344);
xor U8565 (N_8565,N_8168,N_8036);
and U8566 (N_8566,N_8445,N_8131);
xor U8567 (N_8567,N_8136,N_8405);
nand U8568 (N_8568,N_8187,N_8311);
nor U8569 (N_8569,N_8394,N_8251);
nand U8570 (N_8570,N_8051,N_8219);
or U8571 (N_8571,N_8491,N_8069);
xnor U8572 (N_8572,N_8443,N_8408);
and U8573 (N_8573,N_8279,N_8312);
and U8574 (N_8574,N_8410,N_8207);
nor U8575 (N_8575,N_8266,N_8114);
or U8576 (N_8576,N_8262,N_8444);
nand U8577 (N_8577,N_8185,N_8497);
xor U8578 (N_8578,N_8363,N_8048);
xor U8579 (N_8579,N_8247,N_8350);
nor U8580 (N_8580,N_8465,N_8276);
nand U8581 (N_8581,N_8379,N_8367);
and U8582 (N_8582,N_8335,N_8269);
or U8583 (N_8583,N_8196,N_8421);
nand U8584 (N_8584,N_8392,N_8310);
or U8585 (N_8585,N_8229,N_8290);
and U8586 (N_8586,N_8305,N_8171);
or U8587 (N_8587,N_8087,N_8122);
xnor U8588 (N_8588,N_8321,N_8499);
xor U8589 (N_8589,N_8455,N_8378);
xnor U8590 (N_8590,N_8409,N_8217);
nor U8591 (N_8591,N_8203,N_8357);
xnor U8592 (N_8592,N_8330,N_8215);
nand U8593 (N_8593,N_8039,N_8381);
and U8594 (N_8594,N_8442,N_8457);
and U8595 (N_8595,N_8293,N_8212);
or U8596 (N_8596,N_8097,N_8054);
or U8597 (N_8597,N_8233,N_8129);
nor U8598 (N_8598,N_8466,N_8492);
or U8599 (N_8599,N_8360,N_8201);
nand U8600 (N_8600,N_8225,N_8091);
xnor U8601 (N_8601,N_8377,N_8299);
and U8602 (N_8602,N_8399,N_8400);
or U8603 (N_8603,N_8073,N_8438);
nand U8604 (N_8604,N_8390,N_8090);
nor U8605 (N_8605,N_8393,N_8460);
nor U8606 (N_8606,N_8292,N_8155);
xor U8607 (N_8607,N_8241,N_8017);
nor U8608 (N_8608,N_8202,N_8240);
and U8609 (N_8609,N_8060,N_8077);
nand U8610 (N_8610,N_8272,N_8138);
and U8611 (N_8611,N_8192,N_8243);
and U8612 (N_8612,N_8056,N_8472);
or U8613 (N_8613,N_8411,N_8208);
or U8614 (N_8614,N_8453,N_8458);
xnor U8615 (N_8615,N_8078,N_8291);
and U8616 (N_8616,N_8003,N_8146);
and U8617 (N_8617,N_8000,N_8317);
nor U8618 (N_8618,N_8281,N_8428);
nand U8619 (N_8619,N_8313,N_8158);
and U8620 (N_8620,N_8368,N_8041);
or U8621 (N_8621,N_8139,N_8488);
or U8622 (N_8622,N_8152,N_8064);
nand U8623 (N_8623,N_8425,N_8007);
nand U8624 (N_8624,N_8162,N_8074);
or U8625 (N_8625,N_8210,N_8404);
or U8626 (N_8626,N_8439,N_8256);
xnor U8627 (N_8627,N_8137,N_8450);
xnor U8628 (N_8628,N_8329,N_8284);
or U8629 (N_8629,N_8331,N_8117);
nand U8630 (N_8630,N_8151,N_8173);
or U8631 (N_8631,N_8211,N_8275);
and U8632 (N_8632,N_8315,N_8452);
or U8633 (N_8633,N_8199,N_8018);
nor U8634 (N_8634,N_8089,N_8440);
or U8635 (N_8635,N_8309,N_8209);
xnor U8636 (N_8636,N_8050,N_8216);
xnor U8637 (N_8637,N_8286,N_8033);
xnor U8638 (N_8638,N_8150,N_8282);
nand U8639 (N_8639,N_8198,N_8075);
xnor U8640 (N_8640,N_8416,N_8273);
nand U8641 (N_8641,N_8013,N_8341);
or U8642 (N_8642,N_8342,N_8011);
and U8643 (N_8643,N_8294,N_8239);
or U8644 (N_8644,N_8038,N_8396);
nand U8645 (N_8645,N_8231,N_8144);
or U8646 (N_8646,N_8278,N_8230);
or U8647 (N_8647,N_8397,N_8106);
xnor U8648 (N_8648,N_8385,N_8025);
xor U8649 (N_8649,N_8133,N_8008);
nand U8650 (N_8650,N_8448,N_8268);
nor U8651 (N_8651,N_8478,N_8183);
or U8652 (N_8652,N_8323,N_8288);
or U8653 (N_8653,N_8407,N_8327);
nand U8654 (N_8654,N_8375,N_8485);
and U8655 (N_8655,N_8027,N_8271);
or U8656 (N_8656,N_8101,N_8454);
nor U8657 (N_8657,N_8126,N_8094);
nand U8658 (N_8658,N_8172,N_8406);
nand U8659 (N_8659,N_8303,N_8339);
nor U8660 (N_8660,N_8238,N_8206);
xnor U8661 (N_8661,N_8186,N_8223);
and U8662 (N_8662,N_8366,N_8200);
nor U8663 (N_8663,N_8402,N_8145);
nand U8664 (N_8664,N_8307,N_8370);
nor U8665 (N_8665,N_8470,N_8109);
nor U8666 (N_8666,N_8420,N_8447);
or U8667 (N_8667,N_8088,N_8436);
xor U8668 (N_8668,N_8298,N_8142);
nor U8669 (N_8669,N_8154,N_8190);
xor U8670 (N_8670,N_8358,N_8413);
and U8671 (N_8671,N_8165,N_8477);
xnor U8672 (N_8672,N_8274,N_8159);
nor U8673 (N_8673,N_8176,N_8092);
xor U8674 (N_8674,N_8347,N_8042);
nand U8675 (N_8675,N_8236,N_8471);
nand U8676 (N_8676,N_8301,N_8498);
nor U8677 (N_8677,N_8194,N_8248);
xor U8678 (N_8678,N_8174,N_8388);
nor U8679 (N_8679,N_8228,N_8071);
or U8680 (N_8680,N_8468,N_8127);
nor U8681 (N_8681,N_8118,N_8099);
nand U8682 (N_8682,N_8009,N_8422);
xnor U8683 (N_8683,N_8255,N_8343);
xnor U8684 (N_8684,N_8014,N_8319);
or U8685 (N_8685,N_8157,N_8352);
and U8686 (N_8686,N_8389,N_8045);
and U8687 (N_8687,N_8431,N_8296);
nor U8688 (N_8688,N_8384,N_8495);
or U8689 (N_8689,N_8082,N_8434);
and U8690 (N_8690,N_8220,N_8467);
nor U8691 (N_8691,N_8232,N_8258);
nor U8692 (N_8692,N_8197,N_8325);
and U8693 (N_8693,N_8010,N_8081);
and U8694 (N_8694,N_8195,N_8095);
nor U8695 (N_8695,N_8306,N_8304);
nor U8696 (N_8696,N_8124,N_8494);
xor U8697 (N_8697,N_8322,N_8065);
nand U8698 (N_8698,N_8252,N_8463);
or U8699 (N_8699,N_8086,N_8130);
or U8700 (N_8700,N_8031,N_8161);
xnor U8701 (N_8701,N_8326,N_8287);
xor U8702 (N_8702,N_8355,N_8372);
nand U8703 (N_8703,N_8191,N_8112);
and U8704 (N_8704,N_8340,N_8166);
nor U8705 (N_8705,N_8030,N_8265);
xor U8706 (N_8706,N_8163,N_8004);
nor U8707 (N_8707,N_8055,N_8441);
xnor U8708 (N_8708,N_8024,N_8178);
or U8709 (N_8709,N_8386,N_8189);
nor U8710 (N_8710,N_8029,N_8359);
nand U8711 (N_8711,N_8096,N_8179);
or U8712 (N_8712,N_8113,N_8012);
xor U8713 (N_8713,N_8035,N_8026);
nor U8714 (N_8714,N_8204,N_8063);
nand U8715 (N_8715,N_8486,N_8193);
nor U8716 (N_8716,N_8049,N_8058);
and U8717 (N_8717,N_8433,N_8205);
xor U8718 (N_8718,N_8382,N_8170);
and U8719 (N_8719,N_8224,N_8119);
nor U8720 (N_8720,N_8437,N_8141);
or U8721 (N_8721,N_8120,N_8098);
or U8722 (N_8722,N_8387,N_8250);
nand U8723 (N_8723,N_8188,N_8475);
or U8724 (N_8724,N_8116,N_8022);
nand U8725 (N_8725,N_8246,N_8349);
and U8726 (N_8726,N_8028,N_8289);
xnor U8727 (N_8727,N_8469,N_8105);
nor U8728 (N_8728,N_8134,N_8354);
nand U8729 (N_8729,N_8253,N_8123);
or U8730 (N_8730,N_8456,N_8218);
nand U8731 (N_8731,N_8419,N_8429);
nand U8732 (N_8732,N_8006,N_8334);
and U8733 (N_8733,N_8043,N_8260);
nand U8734 (N_8734,N_8222,N_8053);
xnor U8735 (N_8735,N_8324,N_8181);
and U8736 (N_8736,N_8300,N_8369);
or U8737 (N_8737,N_8451,N_8314);
xnor U8738 (N_8738,N_8376,N_8430);
nand U8739 (N_8739,N_8110,N_8234);
nor U8740 (N_8740,N_8493,N_8111);
or U8741 (N_8741,N_8415,N_8371);
nor U8742 (N_8742,N_8473,N_8085);
nand U8743 (N_8743,N_8490,N_8100);
nand U8744 (N_8744,N_8153,N_8044);
nand U8745 (N_8745,N_8482,N_8383);
xor U8746 (N_8746,N_8020,N_8184);
nand U8747 (N_8747,N_8432,N_8462);
or U8748 (N_8748,N_8414,N_8160);
nand U8749 (N_8749,N_8474,N_8148);
and U8750 (N_8750,N_8190,N_8223);
xnor U8751 (N_8751,N_8468,N_8109);
or U8752 (N_8752,N_8159,N_8078);
nand U8753 (N_8753,N_8270,N_8094);
or U8754 (N_8754,N_8033,N_8060);
nand U8755 (N_8755,N_8063,N_8301);
nand U8756 (N_8756,N_8328,N_8133);
and U8757 (N_8757,N_8261,N_8078);
or U8758 (N_8758,N_8385,N_8140);
nand U8759 (N_8759,N_8331,N_8256);
xnor U8760 (N_8760,N_8450,N_8399);
and U8761 (N_8761,N_8210,N_8097);
nand U8762 (N_8762,N_8321,N_8240);
xor U8763 (N_8763,N_8018,N_8060);
nor U8764 (N_8764,N_8334,N_8356);
xor U8765 (N_8765,N_8486,N_8147);
and U8766 (N_8766,N_8036,N_8157);
nor U8767 (N_8767,N_8016,N_8190);
and U8768 (N_8768,N_8099,N_8148);
nand U8769 (N_8769,N_8297,N_8131);
xor U8770 (N_8770,N_8192,N_8072);
xnor U8771 (N_8771,N_8489,N_8377);
nand U8772 (N_8772,N_8298,N_8040);
xnor U8773 (N_8773,N_8357,N_8373);
or U8774 (N_8774,N_8133,N_8215);
and U8775 (N_8775,N_8149,N_8202);
and U8776 (N_8776,N_8415,N_8374);
nor U8777 (N_8777,N_8301,N_8371);
and U8778 (N_8778,N_8288,N_8388);
nand U8779 (N_8779,N_8358,N_8112);
nand U8780 (N_8780,N_8443,N_8363);
and U8781 (N_8781,N_8110,N_8100);
or U8782 (N_8782,N_8498,N_8163);
or U8783 (N_8783,N_8346,N_8310);
or U8784 (N_8784,N_8419,N_8427);
xnor U8785 (N_8785,N_8312,N_8108);
and U8786 (N_8786,N_8087,N_8143);
xnor U8787 (N_8787,N_8340,N_8161);
and U8788 (N_8788,N_8259,N_8491);
nand U8789 (N_8789,N_8419,N_8102);
nor U8790 (N_8790,N_8165,N_8238);
nor U8791 (N_8791,N_8246,N_8198);
nand U8792 (N_8792,N_8125,N_8136);
or U8793 (N_8793,N_8181,N_8299);
nand U8794 (N_8794,N_8332,N_8053);
nand U8795 (N_8795,N_8170,N_8153);
nor U8796 (N_8796,N_8135,N_8109);
and U8797 (N_8797,N_8154,N_8010);
xor U8798 (N_8798,N_8398,N_8010);
and U8799 (N_8799,N_8073,N_8123);
and U8800 (N_8800,N_8082,N_8333);
nor U8801 (N_8801,N_8413,N_8442);
or U8802 (N_8802,N_8113,N_8483);
nor U8803 (N_8803,N_8183,N_8107);
or U8804 (N_8804,N_8463,N_8398);
xor U8805 (N_8805,N_8063,N_8229);
nand U8806 (N_8806,N_8378,N_8272);
and U8807 (N_8807,N_8291,N_8249);
nand U8808 (N_8808,N_8304,N_8443);
and U8809 (N_8809,N_8102,N_8071);
nand U8810 (N_8810,N_8373,N_8127);
and U8811 (N_8811,N_8224,N_8208);
xnor U8812 (N_8812,N_8323,N_8404);
and U8813 (N_8813,N_8201,N_8159);
xnor U8814 (N_8814,N_8385,N_8355);
nand U8815 (N_8815,N_8231,N_8286);
nor U8816 (N_8816,N_8284,N_8150);
nor U8817 (N_8817,N_8296,N_8259);
nor U8818 (N_8818,N_8431,N_8276);
xnor U8819 (N_8819,N_8319,N_8145);
xor U8820 (N_8820,N_8301,N_8073);
nand U8821 (N_8821,N_8187,N_8154);
nand U8822 (N_8822,N_8011,N_8366);
nand U8823 (N_8823,N_8215,N_8006);
nand U8824 (N_8824,N_8438,N_8024);
nand U8825 (N_8825,N_8375,N_8441);
nor U8826 (N_8826,N_8196,N_8141);
or U8827 (N_8827,N_8121,N_8054);
nor U8828 (N_8828,N_8484,N_8268);
and U8829 (N_8829,N_8225,N_8231);
nand U8830 (N_8830,N_8241,N_8413);
nand U8831 (N_8831,N_8063,N_8010);
nand U8832 (N_8832,N_8109,N_8045);
or U8833 (N_8833,N_8234,N_8478);
and U8834 (N_8834,N_8075,N_8136);
or U8835 (N_8835,N_8145,N_8388);
nand U8836 (N_8836,N_8397,N_8409);
and U8837 (N_8837,N_8055,N_8261);
and U8838 (N_8838,N_8470,N_8128);
nor U8839 (N_8839,N_8352,N_8395);
and U8840 (N_8840,N_8284,N_8247);
and U8841 (N_8841,N_8214,N_8057);
nor U8842 (N_8842,N_8346,N_8102);
xor U8843 (N_8843,N_8261,N_8408);
or U8844 (N_8844,N_8284,N_8198);
xor U8845 (N_8845,N_8202,N_8215);
nor U8846 (N_8846,N_8241,N_8381);
xnor U8847 (N_8847,N_8137,N_8489);
nand U8848 (N_8848,N_8199,N_8063);
nor U8849 (N_8849,N_8005,N_8118);
or U8850 (N_8850,N_8400,N_8194);
nor U8851 (N_8851,N_8059,N_8454);
nand U8852 (N_8852,N_8426,N_8211);
nor U8853 (N_8853,N_8485,N_8376);
or U8854 (N_8854,N_8048,N_8284);
nor U8855 (N_8855,N_8303,N_8353);
xnor U8856 (N_8856,N_8051,N_8266);
or U8857 (N_8857,N_8416,N_8118);
nor U8858 (N_8858,N_8449,N_8470);
or U8859 (N_8859,N_8049,N_8372);
xor U8860 (N_8860,N_8086,N_8324);
nand U8861 (N_8861,N_8169,N_8195);
or U8862 (N_8862,N_8417,N_8340);
or U8863 (N_8863,N_8401,N_8215);
nor U8864 (N_8864,N_8023,N_8167);
nand U8865 (N_8865,N_8489,N_8361);
and U8866 (N_8866,N_8296,N_8225);
xnor U8867 (N_8867,N_8127,N_8154);
nor U8868 (N_8868,N_8049,N_8385);
nor U8869 (N_8869,N_8282,N_8104);
xor U8870 (N_8870,N_8377,N_8016);
nor U8871 (N_8871,N_8184,N_8022);
xor U8872 (N_8872,N_8442,N_8385);
xor U8873 (N_8873,N_8126,N_8257);
nand U8874 (N_8874,N_8159,N_8150);
nor U8875 (N_8875,N_8425,N_8409);
and U8876 (N_8876,N_8389,N_8261);
xnor U8877 (N_8877,N_8086,N_8422);
xor U8878 (N_8878,N_8214,N_8327);
xnor U8879 (N_8879,N_8395,N_8268);
nor U8880 (N_8880,N_8398,N_8026);
and U8881 (N_8881,N_8392,N_8400);
nor U8882 (N_8882,N_8275,N_8242);
nor U8883 (N_8883,N_8368,N_8257);
nor U8884 (N_8884,N_8059,N_8109);
xnor U8885 (N_8885,N_8178,N_8428);
nand U8886 (N_8886,N_8305,N_8451);
xnor U8887 (N_8887,N_8138,N_8220);
nand U8888 (N_8888,N_8060,N_8015);
nand U8889 (N_8889,N_8148,N_8220);
or U8890 (N_8890,N_8249,N_8001);
and U8891 (N_8891,N_8429,N_8244);
nand U8892 (N_8892,N_8331,N_8222);
xor U8893 (N_8893,N_8230,N_8257);
and U8894 (N_8894,N_8469,N_8038);
nor U8895 (N_8895,N_8373,N_8406);
nand U8896 (N_8896,N_8218,N_8480);
or U8897 (N_8897,N_8220,N_8124);
or U8898 (N_8898,N_8449,N_8157);
xnor U8899 (N_8899,N_8382,N_8205);
nand U8900 (N_8900,N_8034,N_8321);
nand U8901 (N_8901,N_8405,N_8270);
nand U8902 (N_8902,N_8161,N_8203);
nand U8903 (N_8903,N_8063,N_8169);
xnor U8904 (N_8904,N_8463,N_8271);
xor U8905 (N_8905,N_8344,N_8486);
nand U8906 (N_8906,N_8391,N_8332);
or U8907 (N_8907,N_8050,N_8220);
and U8908 (N_8908,N_8074,N_8283);
or U8909 (N_8909,N_8060,N_8147);
nor U8910 (N_8910,N_8317,N_8025);
nor U8911 (N_8911,N_8040,N_8220);
or U8912 (N_8912,N_8160,N_8117);
xor U8913 (N_8913,N_8465,N_8171);
nor U8914 (N_8914,N_8478,N_8278);
or U8915 (N_8915,N_8313,N_8166);
nand U8916 (N_8916,N_8151,N_8279);
and U8917 (N_8917,N_8431,N_8114);
nand U8918 (N_8918,N_8363,N_8455);
xnor U8919 (N_8919,N_8469,N_8085);
xor U8920 (N_8920,N_8452,N_8210);
xnor U8921 (N_8921,N_8193,N_8213);
xor U8922 (N_8922,N_8009,N_8219);
or U8923 (N_8923,N_8139,N_8258);
nor U8924 (N_8924,N_8023,N_8034);
xnor U8925 (N_8925,N_8256,N_8492);
nor U8926 (N_8926,N_8142,N_8254);
xnor U8927 (N_8927,N_8107,N_8268);
xor U8928 (N_8928,N_8390,N_8092);
or U8929 (N_8929,N_8028,N_8264);
xnor U8930 (N_8930,N_8336,N_8355);
xor U8931 (N_8931,N_8209,N_8032);
nand U8932 (N_8932,N_8028,N_8062);
nor U8933 (N_8933,N_8390,N_8446);
nand U8934 (N_8934,N_8341,N_8081);
nor U8935 (N_8935,N_8051,N_8449);
and U8936 (N_8936,N_8246,N_8027);
nand U8937 (N_8937,N_8492,N_8059);
xnor U8938 (N_8938,N_8209,N_8348);
nand U8939 (N_8939,N_8056,N_8458);
or U8940 (N_8940,N_8036,N_8479);
xor U8941 (N_8941,N_8136,N_8271);
nand U8942 (N_8942,N_8164,N_8185);
nor U8943 (N_8943,N_8143,N_8118);
xor U8944 (N_8944,N_8055,N_8314);
or U8945 (N_8945,N_8387,N_8085);
nor U8946 (N_8946,N_8428,N_8467);
and U8947 (N_8947,N_8426,N_8292);
nand U8948 (N_8948,N_8079,N_8021);
nand U8949 (N_8949,N_8048,N_8312);
and U8950 (N_8950,N_8345,N_8417);
and U8951 (N_8951,N_8378,N_8437);
xor U8952 (N_8952,N_8030,N_8049);
nand U8953 (N_8953,N_8415,N_8047);
xor U8954 (N_8954,N_8474,N_8457);
xor U8955 (N_8955,N_8104,N_8449);
nor U8956 (N_8956,N_8260,N_8082);
nand U8957 (N_8957,N_8396,N_8165);
nor U8958 (N_8958,N_8209,N_8265);
and U8959 (N_8959,N_8011,N_8451);
nand U8960 (N_8960,N_8135,N_8466);
nand U8961 (N_8961,N_8259,N_8435);
and U8962 (N_8962,N_8463,N_8003);
nand U8963 (N_8963,N_8158,N_8297);
or U8964 (N_8964,N_8177,N_8166);
and U8965 (N_8965,N_8117,N_8206);
nor U8966 (N_8966,N_8294,N_8271);
nand U8967 (N_8967,N_8022,N_8261);
nand U8968 (N_8968,N_8305,N_8467);
nand U8969 (N_8969,N_8034,N_8126);
xor U8970 (N_8970,N_8029,N_8048);
nand U8971 (N_8971,N_8475,N_8022);
xor U8972 (N_8972,N_8199,N_8468);
or U8973 (N_8973,N_8053,N_8415);
xor U8974 (N_8974,N_8388,N_8373);
xnor U8975 (N_8975,N_8358,N_8285);
xnor U8976 (N_8976,N_8297,N_8140);
nand U8977 (N_8977,N_8386,N_8028);
or U8978 (N_8978,N_8363,N_8465);
nand U8979 (N_8979,N_8100,N_8357);
or U8980 (N_8980,N_8295,N_8290);
nor U8981 (N_8981,N_8004,N_8251);
nor U8982 (N_8982,N_8051,N_8088);
and U8983 (N_8983,N_8269,N_8353);
or U8984 (N_8984,N_8460,N_8289);
xor U8985 (N_8985,N_8116,N_8257);
and U8986 (N_8986,N_8035,N_8411);
xor U8987 (N_8987,N_8192,N_8038);
nand U8988 (N_8988,N_8086,N_8141);
and U8989 (N_8989,N_8050,N_8424);
nand U8990 (N_8990,N_8350,N_8330);
or U8991 (N_8991,N_8231,N_8380);
or U8992 (N_8992,N_8201,N_8396);
and U8993 (N_8993,N_8462,N_8235);
and U8994 (N_8994,N_8075,N_8195);
xnor U8995 (N_8995,N_8430,N_8126);
nor U8996 (N_8996,N_8425,N_8352);
and U8997 (N_8997,N_8284,N_8405);
nor U8998 (N_8998,N_8487,N_8081);
xnor U8999 (N_8999,N_8149,N_8094);
and U9000 (N_9000,N_8662,N_8766);
or U9001 (N_9001,N_8628,N_8619);
xor U9002 (N_9002,N_8796,N_8891);
xor U9003 (N_9003,N_8977,N_8643);
nand U9004 (N_9004,N_8874,N_8747);
nand U9005 (N_9005,N_8799,N_8802);
xnor U9006 (N_9006,N_8877,N_8566);
nor U9007 (N_9007,N_8688,N_8551);
and U9008 (N_9008,N_8851,N_8961);
nand U9009 (N_9009,N_8920,N_8943);
and U9010 (N_9010,N_8950,N_8785);
nor U9011 (N_9011,N_8758,N_8743);
or U9012 (N_9012,N_8817,N_8836);
nand U9013 (N_9013,N_8801,N_8520);
nor U9014 (N_9014,N_8532,N_8821);
or U9015 (N_9015,N_8718,N_8938);
nand U9016 (N_9016,N_8672,N_8592);
or U9017 (N_9017,N_8835,N_8966);
nand U9018 (N_9018,N_8948,N_8702);
xnor U9019 (N_9019,N_8694,N_8812);
or U9020 (N_9020,N_8654,N_8599);
nor U9021 (N_9021,N_8514,N_8728);
xor U9022 (N_9022,N_8971,N_8924);
nand U9023 (N_9023,N_8954,N_8589);
nand U9024 (N_9024,N_8915,N_8717);
xnor U9025 (N_9025,N_8648,N_8623);
and U9026 (N_9026,N_8576,N_8746);
xnor U9027 (N_9027,N_8893,N_8585);
nor U9028 (N_9028,N_8511,N_8951);
xnor U9029 (N_9029,N_8981,N_8539);
nand U9030 (N_9030,N_8856,N_8629);
nand U9031 (N_9031,N_8755,N_8650);
nand U9032 (N_9032,N_8637,N_8507);
and U9033 (N_9033,N_8724,N_8522);
nor U9034 (N_9034,N_8556,N_8770);
nor U9035 (N_9035,N_8934,N_8897);
and U9036 (N_9036,N_8984,N_8982);
xor U9037 (N_9037,N_8818,N_8940);
nand U9038 (N_9038,N_8819,N_8779);
nor U9039 (N_9039,N_8669,N_8942);
and U9040 (N_9040,N_8614,N_8579);
nor U9041 (N_9041,N_8886,N_8910);
and U9042 (N_9042,N_8871,N_8786);
nor U9043 (N_9043,N_8945,N_8853);
and U9044 (N_9044,N_8793,N_8823);
or U9045 (N_9045,N_8596,N_8881);
xnor U9046 (N_9046,N_8732,N_8882);
xnor U9047 (N_9047,N_8653,N_8788);
and U9048 (N_9048,N_8761,N_8700);
nor U9049 (N_9049,N_8660,N_8610);
nor U9050 (N_9050,N_8635,N_8734);
and U9051 (N_9051,N_8894,N_8537);
nor U9052 (N_9052,N_8754,N_8735);
and U9053 (N_9053,N_8742,N_8565);
nand U9054 (N_9054,N_8800,N_8560);
nor U9055 (N_9055,N_8983,N_8727);
nor U9056 (N_9056,N_8976,N_8606);
or U9057 (N_9057,N_8771,N_8626);
nand U9058 (N_9058,N_8932,N_8768);
and U9059 (N_9059,N_8974,N_8553);
and U9060 (N_9060,N_8816,N_8548);
nor U9061 (N_9061,N_8958,N_8620);
xnor U9062 (N_9062,N_8852,N_8639);
or U9063 (N_9063,N_8839,N_8611);
xor U9064 (N_9064,N_8506,N_8922);
nand U9065 (N_9065,N_8850,N_8904);
nand U9066 (N_9066,N_8921,N_8730);
nand U9067 (N_9067,N_8841,N_8960);
or U9068 (N_9068,N_8757,N_8590);
or U9069 (N_9069,N_8593,N_8760);
or U9070 (N_9070,N_8645,N_8638);
nor U9071 (N_9071,N_8583,N_8925);
nor U9072 (N_9072,N_8655,N_8798);
or U9073 (N_9073,N_8778,N_8965);
and U9074 (N_9074,N_8741,N_8666);
and U9075 (N_9075,N_8518,N_8665);
and U9076 (N_9076,N_8602,N_8545);
xnor U9077 (N_9077,N_8646,N_8946);
and U9078 (N_9078,N_8644,N_8875);
and U9079 (N_9079,N_8573,N_8870);
or U9080 (N_9080,N_8794,N_8753);
nand U9081 (N_9081,N_8675,N_8681);
xnor U9082 (N_9082,N_8918,N_8615);
and U9083 (N_9083,N_8510,N_8519);
or U9084 (N_9084,N_8618,N_8726);
nor U9085 (N_9085,N_8985,N_8538);
nand U9086 (N_9086,N_8873,N_8919);
and U9087 (N_9087,N_8956,N_8616);
nand U9088 (N_9088,N_8679,N_8964);
xnor U9089 (N_9089,N_8909,N_8572);
nand U9090 (N_9090,N_8720,N_8612);
or U9091 (N_9091,N_8561,N_8703);
nor U9092 (N_9092,N_8745,N_8825);
nor U9093 (N_9093,N_8869,N_8959);
and U9094 (N_9094,N_8782,N_8953);
nand U9095 (N_9095,N_8931,N_8831);
xor U9096 (N_9096,N_8708,N_8854);
nand U9097 (N_9097,N_8582,N_8664);
and U9098 (N_9098,N_8670,N_8797);
nor U9099 (N_9099,N_8591,N_8804);
nand U9100 (N_9100,N_8855,N_8863);
or U9101 (N_9101,N_8992,N_8687);
or U9102 (N_9102,N_8697,N_8574);
xnor U9103 (N_9103,N_8916,N_8824);
xor U9104 (N_9104,N_8895,N_8595);
or U9105 (N_9105,N_8581,N_8725);
xnor U9106 (N_9106,N_8883,N_8927);
xor U9107 (N_9107,N_8526,N_8990);
nand U9108 (N_9108,N_8923,N_8947);
xor U9109 (N_9109,N_8994,N_8557);
or U9110 (N_9110,N_8807,N_8563);
and U9111 (N_9111,N_8723,N_8667);
xor U9112 (N_9112,N_8775,N_8978);
nor U9113 (N_9113,N_8685,N_8714);
and U9114 (N_9114,N_8684,N_8903);
or U9115 (N_9115,N_8691,N_8795);
and U9116 (N_9116,N_8791,N_8699);
or U9117 (N_9117,N_8555,N_8827);
or U9118 (N_9118,N_8609,N_8975);
nor U9119 (N_9119,N_8554,N_8955);
nor U9120 (N_9120,N_8762,N_8504);
and U9121 (N_9121,N_8584,N_8859);
xor U9122 (N_9122,N_8907,N_8929);
nor U9123 (N_9123,N_8604,N_8997);
xor U9124 (N_9124,N_8517,N_8678);
nand U9125 (N_9125,N_8858,N_8630);
or U9126 (N_9126,N_8502,N_8968);
nor U9127 (N_9127,N_8868,N_8970);
xnor U9128 (N_9128,N_8764,N_8647);
or U9129 (N_9129,N_8674,N_8663);
and U9130 (N_9130,N_8733,N_8876);
and U9131 (N_9131,N_8657,N_8711);
xnor U9132 (N_9132,N_8826,N_8884);
xor U9133 (N_9133,N_8815,N_8926);
or U9134 (N_9134,N_8906,N_8833);
and U9135 (N_9135,N_8790,N_8568);
and U9136 (N_9136,N_8803,N_8842);
nor U9137 (N_9137,N_8600,N_8999);
and U9138 (N_9138,N_8979,N_8888);
or U9139 (N_9139,N_8658,N_8806);
or U9140 (N_9140,N_8844,N_8707);
nand U9141 (N_9141,N_8696,N_8719);
nand U9142 (N_9142,N_8624,N_8944);
xor U9143 (N_9143,N_8515,N_8750);
or U9144 (N_9144,N_8957,N_8535);
nand U9145 (N_9145,N_8880,N_8721);
nand U9146 (N_9146,N_8503,N_8577);
or U9147 (N_9147,N_8973,N_8636);
and U9148 (N_9148,N_8998,N_8890);
and U9149 (N_9149,N_8748,N_8704);
nor U9150 (N_9150,N_8847,N_8530);
and U9151 (N_9151,N_8980,N_8531);
nor U9152 (N_9152,N_8722,N_8949);
and U9153 (N_9153,N_8731,N_8605);
nand U9154 (N_9154,N_8905,N_8680);
and U9155 (N_9155,N_8772,N_8642);
and U9156 (N_9156,N_8682,N_8969);
and U9157 (N_9157,N_8889,N_8558);
or U9158 (N_9158,N_8587,N_8622);
nand U9159 (N_9159,N_8668,N_8879);
and U9160 (N_9160,N_8617,N_8900);
or U9161 (N_9161,N_8580,N_8784);
nor U9162 (N_9162,N_8987,N_8546);
and U9163 (N_9163,N_8967,N_8513);
nand U9164 (N_9164,N_8578,N_8671);
and U9165 (N_9165,N_8840,N_8763);
or U9166 (N_9166,N_8570,N_8729);
nor U9167 (N_9167,N_8542,N_8597);
or U9168 (N_9168,N_8575,N_8529);
nand U9169 (N_9169,N_8972,N_8509);
xnor U9170 (N_9170,N_8928,N_8834);
nand U9171 (N_9171,N_8547,N_8822);
nor U9172 (N_9172,N_8739,N_8829);
and U9173 (N_9173,N_8941,N_8676);
and U9174 (N_9174,N_8524,N_8712);
nand U9175 (N_9175,N_8810,N_8652);
or U9176 (N_9176,N_8911,N_8588);
nand U9177 (N_9177,N_8751,N_8683);
nor U9178 (N_9178,N_8774,N_8936);
xor U9179 (N_9179,N_8661,N_8773);
or U9180 (N_9180,N_8899,N_8740);
and U9181 (N_9181,N_8536,N_8783);
nor U9182 (N_9182,N_8634,N_8963);
xnor U9183 (N_9183,N_8845,N_8693);
xor U9184 (N_9184,N_8914,N_8861);
xnor U9185 (N_9185,N_8820,N_8737);
nand U9186 (N_9186,N_8843,N_8995);
xor U9187 (N_9187,N_8549,N_8640);
or U9188 (N_9188,N_8902,N_8598);
xnor U9189 (N_9189,N_8986,N_8695);
nor U9190 (N_9190,N_8885,N_8908);
xnor U9191 (N_9191,N_8896,N_8544);
and U9192 (N_9192,N_8705,N_8534);
xnor U9193 (N_9193,N_8659,N_8552);
xnor U9194 (N_9194,N_8550,N_8715);
nor U9195 (N_9195,N_8607,N_8789);
and U9196 (N_9196,N_8736,N_8848);
xor U9197 (N_9197,N_8586,N_8814);
xnor U9198 (N_9198,N_8501,N_8709);
or U9199 (N_9199,N_8787,N_8698);
nand U9200 (N_9200,N_8756,N_8633);
nor U9201 (N_9201,N_8862,N_8866);
nand U9202 (N_9202,N_8769,N_8649);
and U9203 (N_9203,N_8562,N_8792);
nand U9204 (N_9204,N_8752,N_8828);
xor U9205 (N_9205,N_8571,N_8621);
or U9206 (N_9206,N_8878,N_8777);
and U9207 (N_9207,N_8749,N_8867);
nor U9208 (N_9208,N_8838,N_8613);
xnor U9209 (N_9209,N_8543,N_8738);
nor U9210 (N_9210,N_8521,N_8989);
or U9211 (N_9211,N_8701,N_8988);
nor U9212 (N_9212,N_8811,N_8887);
and U9213 (N_9213,N_8860,N_8991);
or U9214 (N_9214,N_8632,N_8809);
and U9215 (N_9215,N_8872,N_8677);
and U9216 (N_9216,N_8559,N_8780);
or U9217 (N_9217,N_8716,N_8690);
nor U9218 (N_9218,N_8781,N_8917);
xnor U9219 (N_9219,N_8505,N_8912);
or U9220 (N_9220,N_8930,N_8641);
nand U9221 (N_9221,N_8837,N_8508);
nor U9222 (N_9222,N_8759,N_8512);
nor U9223 (N_9223,N_8625,N_8656);
xor U9224 (N_9224,N_8525,N_8933);
nand U9225 (N_9225,N_8608,N_8996);
or U9226 (N_9226,N_8937,N_8776);
nor U9227 (N_9227,N_8830,N_8528);
nor U9228 (N_9228,N_8805,N_8686);
xnor U9229 (N_9229,N_8849,N_8857);
and U9230 (N_9230,N_8541,N_8864);
nand U9231 (N_9231,N_8865,N_8962);
and U9232 (N_9232,N_8898,N_8913);
nand U9233 (N_9233,N_8540,N_8692);
nor U9234 (N_9234,N_8808,N_8892);
nor U9235 (N_9235,N_8567,N_8603);
xnor U9236 (N_9236,N_8767,N_8564);
nand U9237 (N_9237,N_8500,N_8744);
xor U9238 (N_9238,N_8689,N_8901);
xnor U9239 (N_9239,N_8713,N_8832);
nand U9240 (N_9240,N_8673,N_8765);
nor U9241 (N_9241,N_8631,N_8706);
nand U9242 (N_9242,N_8846,N_8523);
nor U9243 (N_9243,N_8813,N_8993);
xor U9244 (N_9244,N_8710,N_8527);
nor U9245 (N_9245,N_8627,N_8601);
xnor U9246 (N_9246,N_8569,N_8935);
nor U9247 (N_9247,N_8594,N_8516);
or U9248 (N_9248,N_8952,N_8651);
and U9249 (N_9249,N_8939,N_8533);
or U9250 (N_9250,N_8579,N_8785);
or U9251 (N_9251,N_8996,N_8712);
nand U9252 (N_9252,N_8648,N_8877);
nand U9253 (N_9253,N_8877,N_8908);
nor U9254 (N_9254,N_8945,N_8935);
and U9255 (N_9255,N_8654,N_8922);
or U9256 (N_9256,N_8780,N_8560);
nand U9257 (N_9257,N_8585,N_8511);
nor U9258 (N_9258,N_8993,N_8724);
or U9259 (N_9259,N_8503,N_8709);
nand U9260 (N_9260,N_8594,N_8532);
xnor U9261 (N_9261,N_8946,N_8957);
xnor U9262 (N_9262,N_8507,N_8664);
nand U9263 (N_9263,N_8710,N_8655);
or U9264 (N_9264,N_8754,N_8559);
or U9265 (N_9265,N_8660,N_8981);
or U9266 (N_9266,N_8747,N_8924);
nor U9267 (N_9267,N_8715,N_8767);
nor U9268 (N_9268,N_8504,N_8999);
nor U9269 (N_9269,N_8722,N_8867);
nand U9270 (N_9270,N_8747,N_8616);
nor U9271 (N_9271,N_8905,N_8607);
xnor U9272 (N_9272,N_8950,N_8763);
nor U9273 (N_9273,N_8955,N_8714);
xor U9274 (N_9274,N_8664,N_8915);
or U9275 (N_9275,N_8885,N_8545);
xnor U9276 (N_9276,N_8927,N_8518);
nand U9277 (N_9277,N_8770,N_8866);
xnor U9278 (N_9278,N_8721,N_8719);
or U9279 (N_9279,N_8765,N_8954);
xor U9280 (N_9280,N_8883,N_8921);
and U9281 (N_9281,N_8896,N_8828);
and U9282 (N_9282,N_8743,N_8683);
xnor U9283 (N_9283,N_8665,N_8507);
nand U9284 (N_9284,N_8697,N_8837);
nor U9285 (N_9285,N_8857,N_8654);
nor U9286 (N_9286,N_8745,N_8766);
nand U9287 (N_9287,N_8623,N_8968);
xor U9288 (N_9288,N_8936,N_8517);
and U9289 (N_9289,N_8758,N_8755);
or U9290 (N_9290,N_8591,N_8770);
xnor U9291 (N_9291,N_8965,N_8793);
and U9292 (N_9292,N_8821,N_8717);
xnor U9293 (N_9293,N_8745,N_8536);
or U9294 (N_9294,N_8939,N_8559);
and U9295 (N_9295,N_8715,N_8651);
nor U9296 (N_9296,N_8516,N_8780);
nand U9297 (N_9297,N_8603,N_8659);
or U9298 (N_9298,N_8972,N_8860);
xor U9299 (N_9299,N_8675,N_8551);
nor U9300 (N_9300,N_8622,N_8596);
and U9301 (N_9301,N_8871,N_8647);
nand U9302 (N_9302,N_8823,N_8634);
or U9303 (N_9303,N_8623,N_8888);
xnor U9304 (N_9304,N_8555,N_8595);
nor U9305 (N_9305,N_8515,N_8855);
and U9306 (N_9306,N_8872,N_8753);
nor U9307 (N_9307,N_8866,N_8878);
xor U9308 (N_9308,N_8956,N_8536);
and U9309 (N_9309,N_8778,N_8997);
nor U9310 (N_9310,N_8776,N_8535);
nand U9311 (N_9311,N_8586,N_8901);
and U9312 (N_9312,N_8536,N_8585);
nand U9313 (N_9313,N_8543,N_8802);
and U9314 (N_9314,N_8997,N_8921);
or U9315 (N_9315,N_8680,N_8544);
nand U9316 (N_9316,N_8851,N_8991);
and U9317 (N_9317,N_8818,N_8777);
nor U9318 (N_9318,N_8861,N_8675);
nand U9319 (N_9319,N_8576,N_8719);
and U9320 (N_9320,N_8887,N_8621);
and U9321 (N_9321,N_8990,N_8668);
and U9322 (N_9322,N_8623,N_8539);
xnor U9323 (N_9323,N_8646,N_8809);
xor U9324 (N_9324,N_8530,N_8893);
nor U9325 (N_9325,N_8734,N_8581);
xnor U9326 (N_9326,N_8855,N_8856);
or U9327 (N_9327,N_8583,N_8681);
nor U9328 (N_9328,N_8738,N_8733);
xnor U9329 (N_9329,N_8899,N_8684);
xor U9330 (N_9330,N_8738,N_8892);
or U9331 (N_9331,N_8988,N_8851);
or U9332 (N_9332,N_8634,N_8870);
or U9333 (N_9333,N_8713,N_8642);
and U9334 (N_9334,N_8892,N_8911);
nand U9335 (N_9335,N_8832,N_8837);
nand U9336 (N_9336,N_8957,N_8716);
nor U9337 (N_9337,N_8966,N_8946);
xor U9338 (N_9338,N_8504,N_8960);
xnor U9339 (N_9339,N_8791,N_8883);
or U9340 (N_9340,N_8772,N_8695);
nor U9341 (N_9341,N_8909,N_8886);
and U9342 (N_9342,N_8533,N_8538);
and U9343 (N_9343,N_8665,N_8887);
xnor U9344 (N_9344,N_8660,N_8570);
nor U9345 (N_9345,N_8794,N_8860);
nor U9346 (N_9346,N_8840,N_8853);
or U9347 (N_9347,N_8810,N_8989);
nor U9348 (N_9348,N_8621,N_8811);
or U9349 (N_9349,N_8635,N_8780);
nand U9350 (N_9350,N_8620,N_8643);
and U9351 (N_9351,N_8708,N_8772);
nand U9352 (N_9352,N_8626,N_8534);
nor U9353 (N_9353,N_8686,N_8713);
or U9354 (N_9354,N_8971,N_8807);
or U9355 (N_9355,N_8978,N_8965);
xor U9356 (N_9356,N_8756,N_8881);
nor U9357 (N_9357,N_8541,N_8973);
nor U9358 (N_9358,N_8917,N_8552);
nand U9359 (N_9359,N_8516,N_8990);
and U9360 (N_9360,N_8692,N_8775);
nor U9361 (N_9361,N_8838,N_8588);
nor U9362 (N_9362,N_8730,N_8994);
nand U9363 (N_9363,N_8752,N_8528);
or U9364 (N_9364,N_8926,N_8848);
and U9365 (N_9365,N_8803,N_8548);
or U9366 (N_9366,N_8895,N_8764);
xnor U9367 (N_9367,N_8695,N_8797);
nor U9368 (N_9368,N_8565,N_8893);
nor U9369 (N_9369,N_8701,N_8605);
nand U9370 (N_9370,N_8598,N_8790);
and U9371 (N_9371,N_8630,N_8843);
and U9372 (N_9372,N_8996,N_8603);
nand U9373 (N_9373,N_8918,N_8539);
xnor U9374 (N_9374,N_8887,N_8637);
xnor U9375 (N_9375,N_8947,N_8613);
or U9376 (N_9376,N_8896,N_8954);
and U9377 (N_9377,N_8633,N_8551);
nor U9378 (N_9378,N_8644,N_8566);
and U9379 (N_9379,N_8745,N_8658);
and U9380 (N_9380,N_8819,N_8739);
and U9381 (N_9381,N_8985,N_8924);
or U9382 (N_9382,N_8701,N_8774);
and U9383 (N_9383,N_8527,N_8743);
nand U9384 (N_9384,N_8817,N_8871);
or U9385 (N_9385,N_8891,N_8977);
and U9386 (N_9386,N_8878,N_8644);
and U9387 (N_9387,N_8505,N_8883);
xnor U9388 (N_9388,N_8974,N_8994);
nor U9389 (N_9389,N_8610,N_8612);
nor U9390 (N_9390,N_8745,N_8604);
nand U9391 (N_9391,N_8947,N_8710);
nand U9392 (N_9392,N_8603,N_8717);
nand U9393 (N_9393,N_8555,N_8737);
nand U9394 (N_9394,N_8866,N_8829);
nor U9395 (N_9395,N_8751,N_8509);
and U9396 (N_9396,N_8673,N_8503);
xor U9397 (N_9397,N_8786,N_8633);
xor U9398 (N_9398,N_8851,N_8514);
and U9399 (N_9399,N_8852,N_8624);
nor U9400 (N_9400,N_8933,N_8764);
nor U9401 (N_9401,N_8763,N_8630);
nand U9402 (N_9402,N_8900,N_8514);
or U9403 (N_9403,N_8557,N_8880);
xnor U9404 (N_9404,N_8563,N_8928);
nand U9405 (N_9405,N_8842,N_8812);
and U9406 (N_9406,N_8742,N_8991);
or U9407 (N_9407,N_8978,N_8564);
nand U9408 (N_9408,N_8579,N_8750);
nand U9409 (N_9409,N_8969,N_8519);
nor U9410 (N_9410,N_8548,N_8818);
or U9411 (N_9411,N_8590,N_8639);
and U9412 (N_9412,N_8579,N_8968);
and U9413 (N_9413,N_8959,N_8978);
xnor U9414 (N_9414,N_8983,N_8515);
and U9415 (N_9415,N_8701,N_8576);
nor U9416 (N_9416,N_8587,N_8591);
and U9417 (N_9417,N_8941,N_8729);
nand U9418 (N_9418,N_8664,N_8761);
nor U9419 (N_9419,N_8629,N_8579);
nand U9420 (N_9420,N_8940,N_8639);
nor U9421 (N_9421,N_8803,N_8764);
xnor U9422 (N_9422,N_8887,N_8886);
xor U9423 (N_9423,N_8968,N_8937);
and U9424 (N_9424,N_8628,N_8574);
or U9425 (N_9425,N_8847,N_8998);
xnor U9426 (N_9426,N_8604,N_8807);
nand U9427 (N_9427,N_8903,N_8547);
and U9428 (N_9428,N_8519,N_8950);
nand U9429 (N_9429,N_8780,N_8813);
and U9430 (N_9430,N_8702,N_8990);
xor U9431 (N_9431,N_8950,N_8898);
nand U9432 (N_9432,N_8585,N_8924);
nand U9433 (N_9433,N_8818,N_8963);
or U9434 (N_9434,N_8574,N_8732);
nor U9435 (N_9435,N_8625,N_8592);
xnor U9436 (N_9436,N_8679,N_8821);
and U9437 (N_9437,N_8933,N_8683);
and U9438 (N_9438,N_8911,N_8803);
nand U9439 (N_9439,N_8819,N_8932);
nor U9440 (N_9440,N_8608,N_8958);
nand U9441 (N_9441,N_8851,N_8751);
and U9442 (N_9442,N_8834,N_8515);
xnor U9443 (N_9443,N_8777,N_8571);
nor U9444 (N_9444,N_8613,N_8819);
xnor U9445 (N_9445,N_8900,N_8905);
xnor U9446 (N_9446,N_8625,N_8804);
nor U9447 (N_9447,N_8804,N_8687);
xor U9448 (N_9448,N_8912,N_8828);
xor U9449 (N_9449,N_8874,N_8687);
nand U9450 (N_9450,N_8642,N_8765);
and U9451 (N_9451,N_8628,N_8662);
or U9452 (N_9452,N_8677,N_8834);
or U9453 (N_9453,N_8973,N_8808);
xor U9454 (N_9454,N_8621,N_8858);
nor U9455 (N_9455,N_8728,N_8804);
nand U9456 (N_9456,N_8536,N_8558);
nor U9457 (N_9457,N_8869,N_8584);
xor U9458 (N_9458,N_8848,N_8725);
or U9459 (N_9459,N_8605,N_8834);
and U9460 (N_9460,N_8884,N_8698);
nand U9461 (N_9461,N_8660,N_8885);
nand U9462 (N_9462,N_8953,N_8789);
nor U9463 (N_9463,N_8719,N_8713);
xor U9464 (N_9464,N_8542,N_8611);
xnor U9465 (N_9465,N_8802,N_8879);
nor U9466 (N_9466,N_8765,N_8538);
or U9467 (N_9467,N_8908,N_8748);
or U9468 (N_9468,N_8796,N_8574);
xnor U9469 (N_9469,N_8514,N_8903);
or U9470 (N_9470,N_8759,N_8788);
and U9471 (N_9471,N_8515,N_8959);
nand U9472 (N_9472,N_8897,N_8917);
and U9473 (N_9473,N_8949,N_8950);
nand U9474 (N_9474,N_8985,N_8665);
nand U9475 (N_9475,N_8524,N_8782);
or U9476 (N_9476,N_8639,N_8860);
nand U9477 (N_9477,N_8701,N_8835);
or U9478 (N_9478,N_8839,N_8938);
and U9479 (N_9479,N_8971,N_8545);
or U9480 (N_9480,N_8897,N_8548);
or U9481 (N_9481,N_8529,N_8820);
nor U9482 (N_9482,N_8586,N_8836);
nand U9483 (N_9483,N_8797,N_8976);
xnor U9484 (N_9484,N_8663,N_8666);
and U9485 (N_9485,N_8620,N_8883);
xor U9486 (N_9486,N_8863,N_8953);
nand U9487 (N_9487,N_8760,N_8670);
or U9488 (N_9488,N_8536,N_8772);
nand U9489 (N_9489,N_8834,N_8821);
and U9490 (N_9490,N_8828,N_8550);
and U9491 (N_9491,N_8565,N_8843);
and U9492 (N_9492,N_8509,N_8539);
and U9493 (N_9493,N_8853,N_8520);
nor U9494 (N_9494,N_8809,N_8957);
nor U9495 (N_9495,N_8711,N_8742);
xor U9496 (N_9496,N_8841,N_8971);
or U9497 (N_9497,N_8939,N_8683);
xnor U9498 (N_9498,N_8785,N_8693);
or U9499 (N_9499,N_8685,N_8674);
and U9500 (N_9500,N_9428,N_9477);
nand U9501 (N_9501,N_9124,N_9416);
and U9502 (N_9502,N_9326,N_9373);
nor U9503 (N_9503,N_9492,N_9417);
nor U9504 (N_9504,N_9365,N_9331);
nor U9505 (N_9505,N_9362,N_9069);
nor U9506 (N_9506,N_9142,N_9367);
nor U9507 (N_9507,N_9241,N_9052);
and U9508 (N_9508,N_9121,N_9449);
xor U9509 (N_9509,N_9419,N_9473);
nor U9510 (N_9510,N_9036,N_9329);
nor U9511 (N_9511,N_9466,N_9354);
xor U9512 (N_9512,N_9455,N_9337);
or U9513 (N_9513,N_9424,N_9258);
nand U9514 (N_9514,N_9087,N_9441);
xor U9515 (N_9515,N_9300,N_9443);
nor U9516 (N_9516,N_9135,N_9015);
or U9517 (N_9517,N_9144,N_9308);
and U9518 (N_9518,N_9173,N_9325);
nand U9519 (N_9519,N_9474,N_9030);
xor U9520 (N_9520,N_9145,N_9041);
nand U9521 (N_9521,N_9029,N_9486);
nand U9522 (N_9522,N_9371,N_9407);
xnor U9523 (N_9523,N_9001,N_9249);
or U9524 (N_9524,N_9336,N_9000);
or U9525 (N_9525,N_9434,N_9275);
or U9526 (N_9526,N_9155,N_9463);
and U9527 (N_9527,N_9237,N_9430);
nand U9528 (N_9528,N_9094,N_9098);
and U9529 (N_9529,N_9229,N_9292);
nor U9530 (N_9530,N_9074,N_9127);
xnor U9531 (N_9531,N_9208,N_9277);
nor U9532 (N_9532,N_9396,N_9402);
or U9533 (N_9533,N_9032,N_9202);
or U9534 (N_9534,N_9390,N_9279);
nand U9535 (N_9535,N_9273,N_9255);
nand U9536 (N_9536,N_9060,N_9066);
nor U9537 (N_9537,N_9392,N_9487);
or U9538 (N_9538,N_9379,N_9083);
nand U9539 (N_9539,N_9147,N_9479);
nor U9540 (N_9540,N_9148,N_9011);
or U9541 (N_9541,N_9187,N_9086);
and U9542 (N_9542,N_9388,N_9150);
or U9543 (N_9543,N_9374,N_9276);
xnor U9544 (N_9544,N_9489,N_9157);
and U9545 (N_9545,N_9037,N_9451);
nor U9546 (N_9546,N_9178,N_9028);
nor U9547 (N_9547,N_9395,N_9248);
and U9548 (N_9548,N_9498,N_9118);
or U9549 (N_9549,N_9339,N_9034);
xor U9550 (N_9550,N_9251,N_9188);
nor U9551 (N_9551,N_9038,N_9107);
nand U9552 (N_9552,N_9170,N_9169);
nor U9553 (N_9553,N_9132,N_9432);
nor U9554 (N_9554,N_9447,N_9317);
nand U9555 (N_9555,N_9422,N_9033);
and U9556 (N_9556,N_9082,N_9270);
nor U9557 (N_9557,N_9141,N_9387);
and U9558 (N_9558,N_9024,N_9198);
and U9559 (N_9559,N_9213,N_9008);
and U9560 (N_9560,N_9210,N_9484);
and U9561 (N_9561,N_9233,N_9261);
or U9562 (N_9562,N_9471,N_9195);
xnor U9563 (N_9563,N_9189,N_9214);
and U9564 (N_9564,N_9497,N_9031);
nand U9565 (N_9565,N_9280,N_9151);
nor U9566 (N_9566,N_9257,N_9103);
nor U9567 (N_9567,N_9380,N_9352);
and U9568 (N_9568,N_9359,N_9475);
and U9569 (N_9569,N_9122,N_9081);
or U9570 (N_9570,N_9057,N_9294);
and U9571 (N_9571,N_9154,N_9059);
xor U9572 (N_9572,N_9462,N_9406);
and U9573 (N_9573,N_9223,N_9109);
xnor U9574 (N_9574,N_9310,N_9281);
or U9575 (N_9575,N_9005,N_9482);
nor U9576 (N_9576,N_9491,N_9200);
or U9577 (N_9577,N_9468,N_9146);
nand U9578 (N_9578,N_9334,N_9226);
nor U9579 (N_9579,N_9285,N_9092);
or U9580 (N_9580,N_9314,N_9348);
xnor U9581 (N_9581,N_9481,N_9306);
nand U9582 (N_9582,N_9050,N_9347);
xnor U9583 (N_9583,N_9100,N_9172);
xor U9584 (N_9584,N_9211,N_9240);
nor U9585 (N_9585,N_9408,N_9217);
xor U9586 (N_9586,N_9397,N_9427);
and U9587 (N_9587,N_9368,N_9341);
or U9588 (N_9588,N_9399,N_9168);
and U9589 (N_9589,N_9453,N_9244);
and U9590 (N_9590,N_9360,N_9377);
nand U9591 (N_9591,N_9049,N_9376);
or U9592 (N_9592,N_9420,N_9105);
nor U9593 (N_9593,N_9017,N_9137);
nand U9594 (N_9594,N_9322,N_9394);
and U9595 (N_9595,N_9311,N_9139);
or U9596 (N_9596,N_9070,N_9206);
or U9597 (N_9597,N_9062,N_9435);
or U9598 (N_9598,N_9344,N_9196);
nand U9599 (N_9599,N_9393,N_9126);
xor U9600 (N_9600,N_9176,N_9156);
and U9601 (N_9601,N_9293,N_9400);
and U9602 (N_9602,N_9485,N_9246);
nand U9603 (N_9603,N_9296,N_9180);
xor U9604 (N_9604,N_9191,N_9415);
nor U9605 (N_9605,N_9209,N_9316);
nand U9606 (N_9606,N_9044,N_9287);
and U9607 (N_9607,N_9464,N_9452);
xor U9608 (N_9608,N_9335,N_9426);
nor U9609 (N_9609,N_9253,N_9047);
xor U9610 (N_9610,N_9478,N_9375);
xnor U9611 (N_9611,N_9458,N_9386);
nor U9612 (N_9612,N_9439,N_9252);
nand U9613 (N_9613,N_9013,N_9099);
nor U9614 (N_9614,N_9055,N_9192);
nand U9615 (N_9615,N_9078,N_9265);
nor U9616 (N_9616,N_9269,N_9299);
nand U9617 (N_9617,N_9327,N_9190);
and U9618 (N_9618,N_9174,N_9186);
or U9619 (N_9619,N_9093,N_9051);
xnor U9620 (N_9620,N_9019,N_9429);
or U9621 (N_9621,N_9027,N_9320);
nor U9622 (N_9622,N_9129,N_9490);
or U9623 (N_9623,N_9219,N_9340);
or U9624 (N_9624,N_9254,N_9446);
nand U9625 (N_9625,N_9457,N_9023);
xnor U9626 (N_9626,N_9215,N_9138);
or U9627 (N_9627,N_9260,N_9315);
xnor U9628 (N_9628,N_9267,N_9073);
nor U9629 (N_9629,N_9004,N_9288);
and U9630 (N_9630,N_9425,N_9216);
nor U9631 (N_9631,N_9351,N_9197);
nor U9632 (N_9632,N_9106,N_9222);
nand U9633 (N_9633,N_9134,N_9143);
xnor U9634 (N_9634,N_9480,N_9342);
or U9635 (N_9635,N_9035,N_9193);
and U9636 (N_9636,N_9289,N_9303);
nor U9637 (N_9637,N_9166,N_9469);
nand U9638 (N_9638,N_9467,N_9231);
xor U9639 (N_9639,N_9048,N_9366);
xor U9640 (N_9640,N_9324,N_9112);
xnor U9641 (N_9641,N_9204,N_9272);
and U9642 (N_9642,N_9108,N_9445);
and U9643 (N_9643,N_9496,N_9323);
xnor U9644 (N_9644,N_9101,N_9104);
xnor U9645 (N_9645,N_9307,N_9088);
nor U9646 (N_9646,N_9184,N_9465);
or U9647 (N_9647,N_9022,N_9053);
and U9648 (N_9648,N_9045,N_9181);
xor U9649 (N_9649,N_9330,N_9018);
nor U9650 (N_9650,N_9133,N_9068);
nor U9651 (N_9651,N_9256,N_9403);
and U9652 (N_9652,N_9363,N_9438);
nor U9653 (N_9653,N_9391,N_9221);
and U9654 (N_9654,N_9372,N_9065);
and U9655 (N_9655,N_9071,N_9114);
and U9656 (N_9656,N_9476,N_9321);
and U9657 (N_9657,N_9309,N_9454);
or U9658 (N_9658,N_9056,N_9456);
and U9659 (N_9659,N_9077,N_9021);
or U9660 (N_9660,N_9370,N_9110);
or U9661 (N_9661,N_9115,N_9378);
nand U9662 (N_9662,N_9224,N_9239);
or U9663 (N_9663,N_9123,N_9164);
or U9664 (N_9664,N_9421,N_9385);
and U9665 (N_9665,N_9472,N_9250);
xor U9666 (N_9666,N_9020,N_9167);
or U9667 (N_9667,N_9091,N_9343);
nor U9668 (N_9668,N_9163,N_9194);
nand U9669 (N_9669,N_9383,N_9268);
nor U9670 (N_9670,N_9436,N_9297);
xnor U9671 (N_9671,N_9009,N_9130);
nor U9672 (N_9672,N_9412,N_9042);
nand U9673 (N_9673,N_9437,N_9153);
nand U9674 (N_9674,N_9271,N_9266);
and U9675 (N_9675,N_9090,N_9025);
nor U9676 (N_9676,N_9284,N_9355);
and U9677 (N_9677,N_9274,N_9301);
nor U9678 (N_9678,N_9358,N_9433);
nand U9679 (N_9679,N_9319,N_9003);
or U9680 (N_9680,N_9450,N_9113);
nand U9681 (N_9681,N_9067,N_9460);
nand U9682 (N_9682,N_9085,N_9313);
and U9683 (N_9683,N_9158,N_9201);
and U9684 (N_9684,N_9043,N_9096);
nand U9685 (N_9685,N_9061,N_9054);
xnor U9686 (N_9686,N_9338,N_9010);
nand U9687 (N_9687,N_9409,N_9136);
nor U9688 (N_9688,N_9381,N_9075);
nand U9689 (N_9689,N_9398,N_9072);
xor U9690 (N_9690,N_9389,N_9423);
or U9691 (N_9691,N_9304,N_9161);
or U9692 (N_9692,N_9218,N_9404);
nand U9693 (N_9693,N_9182,N_9076);
or U9694 (N_9694,N_9461,N_9212);
or U9695 (N_9695,N_9418,N_9199);
xor U9696 (N_9696,N_9353,N_9414);
nor U9697 (N_9697,N_9357,N_9230);
xor U9698 (N_9698,N_9245,N_9149);
and U9699 (N_9699,N_9295,N_9384);
xnor U9700 (N_9700,N_9064,N_9236);
nand U9701 (N_9701,N_9159,N_9401);
or U9702 (N_9702,N_9332,N_9058);
xnor U9703 (N_9703,N_9356,N_9470);
and U9704 (N_9704,N_9111,N_9286);
xor U9705 (N_9705,N_9262,N_9203);
nand U9706 (N_9706,N_9350,N_9012);
nor U9707 (N_9707,N_9220,N_9007);
nor U9708 (N_9708,N_9063,N_9278);
xor U9709 (N_9709,N_9312,N_9228);
nand U9710 (N_9710,N_9282,N_9247);
nand U9711 (N_9711,N_9002,N_9459);
xnor U9712 (N_9712,N_9205,N_9227);
or U9713 (N_9713,N_9442,N_9225);
xor U9714 (N_9714,N_9046,N_9345);
and U9715 (N_9715,N_9444,N_9014);
xnor U9716 (N_9716,N_9349,N_9264);
xnor U9717 (N_9717,N_9493,N_9131);
nand U9718 (N_9718,N_9152,N_9207);
or U9719 (N_9719,N_9382,N_9080);
and U9720 (N_9720,N_9243,N_9290);
nor U9721 (N_9721,N_9185,N_9318);
nor U9722 (N_9722,N_9175,N_9305);
nor U9723 (N_9723,N_9302,N_9016);
nand U9724 (N_9724,N_9259,N_9431);
or U9725 (N_9725,N_9183,N_9084);
xor U9726 (N_9726,N_9232,N_9298);
and U9727 (N_9727,N_9039,N_9079);
or U9728 (N_9728,N_9179,N_9488);
nor U9729 (N_9729,N_9160,N_9040);
nor U9730 (N_9730,N_9140,N_9361);
xnor U9731 (N_9731,N_9333,N_9117);
and U9732 (N_9732,N_9125,N_9405);
or U9733 (N_9733,N_9177,N_9369);
and U9734 (N_9734,N_9119,N_9128);
or U9735 (N_9735,N_9364,N_9499);
and U9736 (N_9736,N_9234,N_9291);
xor U9737 (N_9737,N_9162,N_9171);
or U9738 (N_9738,N_9495,N_9006);
nand U9739 (N_9739,N_9102,N_9411);
and U9740 (N_9740,N_9448,N_9346);
xnor U9741 (N_9741,N_9026,N_9120);
nor U9742 (N_9742,N_9413,N_9483);
or U9743 (N_9743,N_9089,N_9263);
or U9744 (N_9744,N_9410,N_9095);
or U9745 (N_9745,N_9097,N_9283);
xnor U9746 (N_9746,N_9440,N_9165);
xor U9747 (N_9747,N_9328,N_9494);
nand U9748 (N_9748,N_9116,N_9235);
nand U9749 (N_9749,N_9242,N_9238);
and U9750 (N_9750,N_9089,N_9435);
and U9751 (N_9751,N_9407,N_9012);
or U9752 (N_9752,N_9103,N_9407);
or U9753 (N_9753,N_9239,N_9328);
nand U9754 (N_9754,N_9063,N_9091);
and U9755 (N_9755,N_9074,N_9201);
nand U9756 (N_9756,N_9379,N_9263);
or U9757 (N_9757,N_9229,N_9373);
or U9758 (N_9758,N_9404,N_9075);
nor U9759 (N_9759,N_9036,N_9219);
nand U9760 (N_9760,N_9388,N_9376);
xnor U9761 (N_9761,N_9347,N_9322);
xor U9762 (N_9762,N_9026,N_9403);
nor U9763 (N_9763,N_9161,N_9259);
nand U9764 (N_9764,N_9446,N_9190);
nor U9765 (N_9765,N_9460,N_9237);
nand U9766 (N_9766,N_9082,N_9334);
and U9767 (N_9767,N_9045,N_9419);
xor U9768 (N_9768,N_9019,N_9196);
nor U9769 (N_9769,N_9176,N_9129);
and U9770 (N_9770,N_9410,N_9478);
or U9771 (N_9771,N_9442,N_9131);
nor U9772 (N_9772,N_9437,N_9321);
nor U9773 (N_9773,N_9298,N_9010);
or U9774 (N_9774,N_9463,N_9065);
and U9775 (N_9775,N_9213,N_9488);
xor U9776 (N_9776,N_9453,N_9407);
or U9777 (N_9777,N_9058,N_9417);
nor U9778 (N_9778,N_9460,N_9003);
and U9779 (N_9779,N_9022,N_9219);
nor U9780 (N_9780,N_9039,N_9350);
or U9781 (N_9781,N_9242,N_9174);
nand U9782 (N_9782,N_9474,N_9177);
nand U9783 (N_9783,N_9149,N_9321);
nor U9784 (N_9784,N_9396,N_9497);
nor U9785 (N_9785,N_9304,N_9011);
xnor U9786 (N_9786,N_9314,N_9373);
or U9787 (N_9787,N_9333,N_9223);
or U9788 (N_9788,N_9454,N_9063);
xor U9789 (N_9789,N_9128,N_9039);
xor U9790 (N_9790,N_9282,N_9221);
xor U9791 (N_9791,N_9195,N_9019);
xor U9792 (N_9792,N_9121,N_9322);
xor U9793 (N_9793,N_9270,N_9132);
nand U9794 (N_9794,N_9267,N_9070);
and U9795 (N_9795,N_9366,N_9164);
or U9796 (N_9796,N_9083,N_9099);
nor U9797 (N_9797,N_9337,N_9418);
or U9798 (N_9798,N_9417,N_9486);
or U9799 (N_9799,N_9000,N_9424);
or U9800 (N_9800,N_9099,N_9332);
nand U9801 (N_9801,N_9105,N_9464);
xor U9802 (N_9802,N_9284,N_9162);
nor U9803 (N_9803,N_9069,N_9275);
xnor U9804 (N_9804,N_9065,N_9019);
nor U9805 (N_9805,N_9418,N_9151);
or U9806 (N_9806,N_9085,N_9068);
and U9807 (N_9807,N_9262,N_9140);
xor U9808 (N_9808,N_9376,N_9063);
nand U9809 (N_9809,N_9124,N_9032);
nor U9810 (N_9810,N_9444,N_9178);
and U9811 (N_9811,N_9053,N_9322);
nand U9812 (N_9812,N_9020,N_9340);
or U9813 (N_9813,N_9386,N_9232);
nand U9814 (N_9814,N_9364,N_9222);
or U9815 (N_9815,N_9490,N_9109);
xor U9816 (N_9816,N_9381,N_9337);
xnor U9817 (N_9817,N_9035,N_9137);
or U9818 (N_9818,N_9252,N_9271);
nor U9819 (N_9819,N_9099,N_9022);
nand U9820 (N_9820,N_9053,N_9287);
or U9821 (N_9821,N_9090,N_9471);
and U9822 (N_9822,N_9242,N_9244);
nand U9823 (N_9823,N_9101,N_9030);
nand U9824 (N_9824,N_9137,N_9222);
or U9825 (N_9825,N_9011,N_9067);
xnor U9826 (N_9826,N_9495,N_9202);
and U9827 (N_9827,N_9045,N_9327);
nor U9828 (N_9828,N_9365,N_9238);
xnor U9829 (N_9829,N_9335,N_9283);
and U9830 (N_9830,N_9478,N_9143);
nand U9831 (N_9831,N_9419,N_9243);
xor U9832 (N_9832,N_9129,N_9287);
and U9833 (N_9833,N_9267,N_9321);
or U9834 (N_9834,N_9344,N_9153);
and U9835 (N_9835,N_9130,N_9100);
and U9836 (N_9836,N_9461,N_9419);
xnor U9837 (N_9837,N_9407,N_9210);
xnor U9838 (N_9838,N_9481,N_9023);
nor U9839 (N_9839,N_9424,N_9458);
and U9840 (N_9840,N_9103,N_9118);
nand U9841 (N_9841,N_9139,N_9039);
nor U9842 (N_9842,N_9404,N_9469);
or U9843 (N_9843,N_9353,N_9459);
nor U9844 (N_9844,N_9298,N_9043);
nor U9845 (N_9845,N_9141,N_9235);
xnor U9846 (N_9846,N_9082,N_9198);
nand U9847 (N_9847,N_9098,N_9328);
and U9848 (N_9848,N_9384,N_9101);
nand U9849 (N_9849,N_9372,N_9133);
xnor U9850 (N_9850,N_9306,N_9186);
nand U9851 (N_9851,N_9403,N_9029);
nor U9852 (N_9852,N_9343,N_9376);
and U9853 (N_9853,N_9117,N_9345);
nor U9854 (N_9854,N_9265,N_9440);
nand U9855 (N_9855,N_9167,N_9271);
xor U9856 (N_9856,N_9056,N_9015);
nor U9857 (N_9857,N_9361,N_9069);
and U9858 (N_9858,N_9481,N_9210);
xnor U9859 (N_9859,N_9335,N_9307);
nand U9860 (N_9860,N_9138,N_9051);
nand U9861 (N_9861,N_9026,N_9459);
nor U9862 (N_9862,N_9111,N_9070);
and U9863 (N_9863,N_9284,N_9051);
nand U9864 (N_9864,N_9327,N_9068);
or U9865 (N_9865,N_9467,N_9177);
xnor U9866 (N_9866,N_9279,N_9169);
nand U9867 (N_9867,N_9237,N_9105);
or U9868 (N_9868,N_9314,N_9128);
or U9869 (N_9869,N_9178,N_9300);
or U9870 (N_9870,N_9235,N_9341);
and U9871 (N_9871,N_9455,N_9476);
and U9872 (N_9872,N_9213,N_9073);
or U9873 (N_9873,N_9016,N_9194);
xor U9874 (N_9874,N_9401,N_9205);
and U9875 (N_9875,N_9444,N_9350);
nand U9876 (N_9876,N_9341,N_9385);
nand U9877 (N_9877,N_9336,N_9249);
or U9878 (N_9878,N_9292,N_9264);
nand U9879 (N_9879,N_9373,N_9125);
or U9880 (N_9880,N_9256,N_9148);
and U9881 (N_9881,N_9346,N_9050);
nor U9882 (N_9882,N_9456,N_9162);
and U9883 (N_9883,N_9191,N_9002);
xor U9884 (N_9884,N_9234,N_9355);
nor U9885 (N_9885,N_9391,N_9412);
nand U9886 (N_9886,N_9372,N_9442);
nor U9887 (N_9887,N_9033,N_9183);
nor U9888 (N_9888,N_9478,N_9416);
or U9889 (N_9889,N_9032,N_9030);
xnor U9890 (N_9890,N_9150,N_9473);
xor U9891 (N_9891,N_9111,N_9200);
xor U9892 (N_9892,N_9319,N_9391);
nand U9893 (N_9893,N_9097,N_9365);
nor U9894 (N_9894,N_9062,N_9197);
nor U9895 (N_9895,N_9103,N_9068);
xnor U9896 (N_9896,N_9261,N_9006);
nor U9897 (N_9897,N_9458,N_9394);
and U9898 (N_9898,N_9496,N_9033);
and U9899 (N_9899,N_9418,N_9049);
xor U9900 (N_9900,N_9383,N_9344);
nor U9901 (N_9901,N_9424,N_9322);
nor U9902 (N_9902,N_9445,N_9251);
xnor U9903 (N_9903,N_9297,N_9243);
or U9904 (N_9904,N_9044,N_9087);
nor U9905 (N_9905,N_9076,N_9409);
nor U9906 (N_9906,N_9197,N_9404);
xnor U9907 (N_9907,N_9486,N_9438);
xor U9908 (N_9908,N_9462,N_9409);
xor U9909 (N_9909,N_9227,N_9414);
or U9910 (N_9910,N_9055,N_9057);
nand U9911 (N_9911,N_9026,N_9390);
nand U9912 (N_9912,N_9037,N_9252);
nand U9913 (N_9913,N_9293,N_9152);
or U9914 (N_9914,N_9342,N_9180);
or U9915 (N_9915,N_9009,N_9393);
nand U9916 (N_9916,N_9043,N_9463);
nand U9917 (N_9917,N_9482,N_9432);
xor U9918 (N_9918,N_9289,N_9232);
or U9919 (N_9919,N_9417,N_9267);
xnor U9920 (N_9920,N_9239,N_9000);
xor U9921 (N_9921,N_9469,N_9144);
nor U9922 (N_9922,N_9106,N_9462);
nor U9923 (N_9923,N_9105,N_9073);
and U9924 (N_9924,N_9448,N_9200);
and U9925 (N_9925,N_9176,N_9428);
nand U9926 (N_9926,N_9142,N_9055);
and U9927 (N_9927,N_9127,N_9482);
nor U9928 (N_9928,N_9381,N_9385);
nor U9929 (N_9929,N_9138,N_9182);
nor U9930 (N_9930,N_9355,N_9335);
xnor U9931 (N_9931,N_9361,N_9342);
nand U9932 (N_9932,N_9415,N_9098);
or U9933 (N_9933,N_9259,N_9277);
or U9934 (N_9934,N_9118,N_9486);
xnor U9935 (N_9935,N_9246,N_9442);
nor U9936 (N_9936,N_9113,N_9332);
nor U9937 (N_9937,N_9210,N_9101);
xor U9938 (N_9938,N_9049,N_9321);
nor U9939 (N_9939,N_9410,N_9184);
or U9940 (N_9940,N_9295,N_9400);
or U9941 (N_9941,N_9300,N_9324);
nand U9942 (N_9942,N_9381,N_9215);
or U9943 (N_9943,N_9062,N_9307);
or U9944 (N_9944,N_9327,N_9424);
and U9945 (N_9945,N_9411,N_9283);
nor U9946 (N_9946,N_9464,N_9213);
nand U9947 (N_9947,N_9241,N_9313);
nand U9948 (N_9948,N_9146,N_9236);
nand U9949 (N_9949,N_9076,N_9324);
nand U9950 (N_9950,N_9355,N_9161);
and U9951 (N_9951,N_9371,N_9459);
nand U9952 (N_9952,N_9335,N_9471);
xor U9953 (N_9953,N_9315,N_9022);
and U9954 (N_9954,N_9034,N_9132);
nor U9955 (N_9955,N_9489,N_9256);
nand U9956 (N_9956,N_9253,N_9011);
nand U9957 (N_9957,N_9258,N_9354);
or U9958 (N_9958,N_9139,N_9288);
and U9959 (N_9959,N_9497,N_9128);
nand U9960 (N_9960,N_9300,N_9320);
nand U9961 (N_9961,N_9412,N_9487);
xnor U9962 (N_9962,N_9378,N_9250);
and U9963 (N_9963,N_9293,N_9131);
and U9964 (N_9964,N_9117,N_9401);
or U9965 (N_9965,N_9111,N_9273);
nand U9966 (N_9966,N_9232,N_9265);
xnor U9967 (N_9967,N_9113,N_9368);
nor U9968 (N_9968,N_9132,N_9382);
xor U9969 (N_9969,N_9227,N_9106);
xor U9970 (N_9970,N_9117,N_9356);
nand U9971 (N_9971,N_9175,N_9126);
or U9972 (N_9972,N_9036,N_9276);
xnor U9973 (N_9973,N_9370,N_9426);
or U9974 (N_9974,N_9183,N_9224);
nand U9975 (N_9975,N_9482,N_9083);
nand U9976 (N_9976,N_9209,N_9281);
and U9977 (N_9977,N_9319,N_9177);
nor U9978 (N_9978,N_9252,N_9176);
or U9979 (N_9979,N_9075,N_9326);
or U9980 (N_9980,N_9041,N_9286);
nand U9981 (N_9981,N_9225,N_9197);
and U9982 (N_9982,N_9427,N_9237);
xnor U9983 (N_9983,N_9207,N_9300);
or U9984 (N_9984,N_9296,N_9139);
nor U9985 (N_9985,N_9021,N_9324);
nand U9986 (N_9986,N_9491,N_9000);
nand U9987 (N_9987,N_9438,N_9493);
xnor U9988 (N_9988,N_9366,N_9097);
nor U9989 (N_9989,N_9358,N_9360);
xor U9990 (N_9990,N_9499,N_9304);
or U9991 (N_9991,N_9176,N_9136);
or U9992 (N_9992,N_9055,N_9416);
or U9993 (N_9993,N_9392,N_9021);
or U9994 (N_9994,N_9413,N_9031);
xor U9995 (N_9995,N_9329,N_9131);
and U9996 (N_9996,N_9243,N_9209);
nand U9997 (N_9997,N_9456,N_9340);
xnor U9998 (N_9998,N_9200,N_9171);
xnor U9999 (N_9999,N_9003,N_9077);
xor U10000 (N_10000,N_9528,N_9819);
and U10001 (N_10001,N_9527,N_9577);
xnor U10002 (N_10002,N_9739,N_9617);
and U10003 (N_10003,N_9638,N_9817);
xor U10004 (N_10004,N_9595,N_9635);
xor U10005 (N_10005,N_9984,N_9969);
or U10006 (N_10006,N_9601,N_9772);
and U10007 (N_10007,N_9594,N_9636);
nor U10008 (N_10008,N_9782,N_9626);
xor U10009 (N_10009,N_9725,N_9987);
or U10010 (N_10010,N_9812,N_9986);
nor U10011 (N_10011,N_9976,N_9671);
and U10012 (N_10012,N_9608,N_9687);
or U10013 (N_10013,N_9643,N_9702);
xnor U10014 (N_10014,N_9700,N_9720);
and U10015 (N_10015,N_9914,N_9569);
xor U10016 (N_10016,N_9688,N_9717);
and U10017 (N_10017,N_9565,N_9933);
and U10018 (N_10018,N_9654,N_9848);
and U10019 (N_10019,N_9691,N_9925);
and U10020 (N_10020,N_9821,N_9514);
and U10021 (N_10021,N_9830,N_9781);
nor U10022 (N_10022,N_9934,N_9652);
and U10023 (N_10023,N_9982,N_9944);
nor U10024 (N_10024,N_9784,N_9723);
nand U10025 (N_10025,N_9795,N_9731);
nand U10026 (N_10026,N_9815,N_9680);
nand U10027 (N_10027,N_9648,N_9946);
and U10028 (N_10028,N_9997,N_9697);
and U10029 (N_10029,N_9615,N_9568);
nand U10030 (N_10030,N_9541,N_9765);
or U10031 (N_10031,N_9742,N_9502);
and U10032 (N_10032,N_9573,N_9834);
or U10033 (N_10033,N_9836,N_9869);
or U10034 (N_10034,N_9953,N_9837);
or U10035 (N_10035,N_9898,N_9983);
nand U10036 (N_10036,N_9818,N_9543);
nor U10037 (N_10037,N_9508,N_9651);
nor U10038 (N_10038,N_9631,N_9597);
nand U10039 (N_10039,N_9932,N_9961);
nor U10040 (N_10040,N_9531,N_9604);
nand U10041 (N_10041,N_9832,N_9753);
xnor U10042 (N_10042,N_9999,N_9586);
xor U10043 (N_10043,N_9920,N_9589);
or U10044 (N_10044,N_9909,N_9672);
xor U10045 (N_10045,N_9555,N_9979);
xor U10046 (N_10046,N_9730,N_9800);
nor U10047 (N_10047,N_9655,N_9596);
or U10048 (N_10048,N_9995,N_9501);
nor U10049 (N_10049,N_9685,N_9590);
nand U10050 (N_10050,N_9851,N_9978);
or U10051 (N_10051,N_9841,N_9805);
and U10052 (N_10052,N_9644,N_9534);
nor U10053 (N_10053,N_9574,N_9560);
and U10054 (N_10054,N_9828,N_9770);
nand U10055 (N_10055,N_9639,N_9811);
and U10056 (N_10056,N_9764,N_9535);
or U10057 (N_10057,N_9599,N_9799);
nor U10058 (N_10058,N_9657,N_9509);
or U10059 (N_10059,N_9939,N_9642);
and U10060 (N_10060,N_9632,N_9647);
nand U10061 (N_10061,N_9641,N_9855);
or U10062 (N_10062,N_9542,N_9558);
nand U10063 (N_10063,N_9940,N_9669);
xor U10064 (N_10064,N_9780,N_9945);
nor U10065 (N_10065,N_9516,N_9899);
nand U10066 (N_10066,N_9876,N_9549);
or U10067 (N_10067,N_9538,N_9689);
or U10068 (N_10068,N_9958,N_9751);
and U10069 (N_10069,N_9718,N_9522);
and U10070 (N_10070,N_9695,N_9658);
nand U10071 (N_10071,N_9826,N_9930);
xor U10072 (N_10072,N_9552,N_9889);
and U10073 (N_10073,N_9845,N_9884);
xnor U10074 (N_10074,N_9910,N_9735);
nand U10075 (N_10075,N_9518,N_9745);
xnor U10076 (N_10076,N_9532,N_9778);
nand U10077 (N_10077,N_9622,N_9992);
or U10078 (N_10078,N_9544,N_9540);
xnor U10079 (N_10079,N_9551,N_9686);
and U10080 (N_10080,N_9754,N_9748);
and U10081 (N_10081,N_9653,N_9500);
or U10082 (N_10082,N_9714,N_9874);
xor U10083 (N_10083,N_9867,N_9530);
nor U10084 (N_10084,N_9853,N_9504);
and U10085 (N_10085,N_9775,N_9791);
nor U10086 (N_10086,N_9667,N_9557);
xor U10087 (N_10087,N_9768,N_9779);
nand U10088 (N_10088,N_9873,N_9980);
or U10089 (N_10089,N_9835,N_9734);
xor U10090 (N_10090,N_9513,N_9825);
and U10091 (N_10091,N_9762,N_9690);
or U10092 (N_10092,N_9776,N_9715);
or U10093 (N_10093,N_9550,N_9561);
nand U10094 (N_10094,N_9892,N_9810);
xor U10095 (N_10095,N_9807,N_9760);
nor U10096 (N_10096,N_9875,N_9916);
or U10097 (N_10097,N_9526,N_9600);
and U10098 (N_10098,N_9750,N_9882);
and U10099 (N_10099,N_9693,N_9843);
nand U10100 (N_10100,N_9554,N_9582);
nor U10101 (N_10101,N_9736,N_9732);
nor U10102 (N_10102,N_9880,N_9763);
xnor U10103 (N_10103,N_9571,N_9709);
and U10104 (N_10104,N_9957,N_9840);
xor U10105 (N_10105,N_9860,N_9621);
xor U10106 (N_10106,N_9793,N_9878);
or U10107 (N_10107,N_9895,N_9623);
or U10108 (N_10108,N_9668,N_9646);
and U10109 (N_10109,N_9996,N_9525);
xor U10110 (N_10110,N_9801,N_9786);
or U10111 (N_10111,N_9578,N_9808);
nand U10112 (N_10112,N_9896,N_9728);
nand U10113 (N_10113,N_9906,N_9517);
xor U10114 (N_10114,N_9673,N_9656);
and U10115 (N_10115,N_9719,N_9607);
and U10116 (N_10116,N_9816,N_9902);
or U10117 (N_10117,N_9507,N_9901);
xnor U10118 (N_10118,N_9907,N_9703);
or U10119 (N_10119,N_9881,N_9602);
nand U10120 (N_10120,N_9804,N_9798);
nor U10121 (N_10121,N_9698,N_9660);
xnor U10122 (N_10122,N_9955,N_9774);
nor U10123 (N_10123,N_9822,N_9645);
nand U10124 (N_10124,N_9633,N_9994);
and U10125 (N_10125,N_9659,N_9975);
xor U10126 (N_10126,N_9894,N_9966);
nand U10127 (N_10127,N_9827,N_9905);
nor U10128 (N_10128,N_9721,N_9640);
and U10129 (N_10129,N_9971,N_9759);
and U10130 (N_10130,N_9922,N_9985);
and U10131 (N_10131,N_9972,N_9785);
nor U10132 (N_10132,N_9846,N_9575);
nand U10133 (N_10133,N_9796,N_9942);
nor U10134 (N_10134,N_9701,N_9548);
nand U10135 (N_10135,N_9831,N_9842);
nand U10136 (N_10136,N_9684,N_9885);
nand U10137 (N_10137,N_9929,N_9564);
nor U10138 (N_10138,N_9960,N_9908);
and U10139 (N_10139,N_9973,N_9663);
nand U10140 (N_10140,N_9611,N_9954);
or U10141 (N_10141,N_9588,N_9592);
nor U10142 (N_10142,N_9861,N_9612);
nor U10143 (N_10143,N_9678,N_9625);
or U10144 (N_10144,N_9814,N_9959);
and U10145 (N_10145,N_9707,N_9512);
and U10146 (N_10146,N_9727,N_9917);
nand U10147 (N_10147,N_9566,N_9886);
and U10148 (N_10148,N_9950,N_9809);
or U10149 (N_10149,N_9912,N_9806);
nor U10150 (N_10150,N_9743,N_9729);
or U10151 (N_10151,N_9533,N_9813);
xor U10152 (N_10152,N_9724,N_9581);
xnor U10153 (N_10153,N_9563,N_9579);
nor U10154 (N_10154,N_9794,N_9593);
xor U10155 (N_10155,N_9505,N_9629);
nand U10156 (N_10156,N_9562,N_9769);
xor U10157 (N_10157,N_9918,N_9584);
nor U10158 (N_10158,N_9741,N_9503);
nor U10159 (N_10159,N_9890,N_9587);
or U10160 (N_10160,N_9737,N_9649);
xnor U10161 (N_10161,N_9928,N_9948);
or U10162 (N_10162,N_9974,N_9967);
and U10163 (N_10163,N_9936,N_9692);
xnor U10164 (N_10164,N_9598,N_9802);
nand U10165 (N_10165,N_9634,N_9650);
nor U10166 (N_10166,N_9758,N_9704);
and U10167 (N_10167,N_9941,N_9537);
and U10168 (N_10168,N_9977,N_9773);
and U10169 (N_10169,N_9877,N_9547);
and U10170 (N_10170,N_9570,N_9792);
nor U10171 (N_10171,N_9591,N_9897);
nand U10172 (N_10172,N_9937,N_9614);
xor U10173 (N_10173,N_9755,N_9767);
nor U10174 (N_10174,N_9850,N_9964);
nand U10175 (N_10175,N_9887,N_9858);
nor U10176 (N_10176,N_9662,N_9998);
or U10177 (N_10177,N_9713,N_9520);
nor U10178 (N_10178,N_9722,N_9519);
xnor U10179 (N_10179,N_9556,N_9833);
and U10180 (N_10180,N_9740,N_9852);
and U10181 (N_10181,N_9871,N_9610);
nand U10182 (N_10182,N_9866,N_9824);
xor U10183 (N_10183,N_9787,N_9536);
or U10184 (N_10184,N_9803,N_9864);
nor U10185 (N_10185,N_9696,N_9956);
xor U10186 (N_10186,N_9847,N_9854);
xnor U10187 (N_10187,N_9926,N_9559);
xnor U10188 (N_10188,N_9583,N_9738);
nor U10189 (N_10189,N_9529,N_9524);
or U10190 (N_10190,N_9628,N_9756);
and U10191 (N_10191,N_9726,N_9771);
nand U10192 (N_10192,N_9844,N_9988);
xor U10193 (N_10193,N_9893,N_9790);
xor U10194 (N_10194,N_9572,N_9951);
nor U10195 (N_10195,N_9619,N_9747);
xnor U10196 (N_10196,N_9924,N_9708);
nor U10197 (N_10197,N_9839,N_9921);
and U10198 (N_10198,N_9888,N_9510);
or U10199 (N_10199,N_9838,N_9911);
nand U10200 (N_10200,N_9661,N_9706);
nor U10201 (N_10201,N_9609,N_9947);
nor U10202 (N_10202,N_9968,N_9938);
xor U10203 (N_10203,N_9935,N_9630);
nor U10204 (N_10204,N_9823,N_9949);
or U10205 (N_10205,N_9757,N_9962);
xor U10206 (N_10206,N_9923,N_9675);
and U10207 (N_10207,N_9506,N_9670);
or U10208 (N_10208,N_9783,N_9683);
xor U10209 (N_10209,N_9679,N_9789);
nor U10210 (N_10210,N_9865,N_9863);
nor U10211 (N_10211,N_9970,N_9637);
nor U10212 (N_10212,N_9576,N_9931);
or U10213 (N_10213,N_9712,N_9943);
nand U10214 (N_10214,N_9511,N_9963);
nand U10215 (N_10215,N_9915,N_9539);
and U10216 (N_10216,N_9681,N_9857);
nor U10217 (N_10217,N_9676,N_9952);
or U10218 (N_10218,N_9618,N_9515);
or U10219 (N_10219,N_9989,N_9677);
nand U10220 (N_10220,N_9616,N_9891);
xnor U10221 (N_10221,N_9927,N_9605);
nor U10222 (N_10222,N_9900,N_9746);
and U10223 (N_10223,N_9761,N_9521);
and U10224 (N_10224,N_9859,N_9919);
or U10225 (N_10225,N_9879,N_9870);
nor U10226 (N_10226,N_9567,N_9913);
nand U10227 (N_10227,N_9553,N_9777);
xor U10228 (N_10228,N_9990,N_9624);
nor U10229 (N_10229,N_9749,N_9705);
and U10230 (N_10230,N_9849,N_9883);
or U10231 (N_10231,N_9716,N_9620);
nand U10232 (N_10232,N_9991,N_9856);
or U10233 (N_10233,N_9694,N_9904);
nor U10234 (N_10234,N_9711,N_9788);
or U10235 (N_10235,N_9674,N_9613);
nand U10236 (N_10236,N_9981,N_9820);
and U10237 (N_10237,N_9829,N_9682);
nor U10238 (N_10238,N_9903,N_9699);
or U10239 (N_10239,N_9580,N_9862);
nand U10240 (N_10240,N_9993,N_9797);
nor U10241 (N_10241,N_9666,N_9606);
nor U10242 (N_10242,N_9710,N_9766);
and U10243 (N_10243,N_9872,N_9627);
xor U10244 (N_10244,N_9664,N_9665);
or U10245 (N_10245,N_9523,N_9585);
or U10246 (N_10246,N_9744,N_9603);
or U10247 (N_10247,N_9545,N_9965);
and U10248 (N_10248,N_9546,N_9752);
or U10249 (N_10249,N_9733,N_9868);
nor U10250 (N_10250,N_9654,N_9897);
xnor U10251 (N_10251,N_9553,N_9767);
nand U10252 (N_10252,N_9790,N_9560);
or U10253 (N_10253,N_9839,N_9844);
or U10254 (N_10254,N_9558,N_9817);
and U10255 (N_10255,N_9698,N_9886);
and U10256 (N_10256,N_9555,N_9675);
or U10257 (N_10257,N_9742,N_9761);
or U10258 (N_10258,N_9524,N_9883);
nor U10259 (N_10259,N_9931,N_9731);
nand U10260 (N_10260,N_9827,N_9919);
or U10261 (N_10261,N_9674,N_9956);
nand U10262 (N_10262,N_9880,N_9551);
or U10263 (N_10263,N_9666,N_9677);
xor U10264 (N_10264,N_9767,N_9682);
xor U10265 (N_10265,N_9669,N_9630);
or U10266 (N_10266,N_9558,N_9546);
nor U10267 (N_10267,N_9611,N_9913);
or U10268 (N_10268,N_9741,N_9719);
nor U10269 (N_10269,N_9832,N_9715);
and U10270 (N_10270,N_9682,N_9868);
and U10271 (N_10271,N_9767,N_9544);
or U10272 (N_10272,N_9550,N_9723);
or U10273 (N_10273,N_9734,N_9967);
or U10274 (N_10274,N_9531,N_9789);
nand U10275 (N_10275,N_9910,N_9600);
nand U10276 (N_10276,N_9885,N_9890);
xnor U10277 (N_10277,N_9866,N_9741);
or U10278 (N_10278,N_9742,N_9895);
nand U10279 (N_10279,N_9876,N_9620);
or U10280 (N_10280,N_9673,N_9756);
nand U10281 (N_10281,N_9514,N_9840);
nand U10282 (N_10282,N_9711,N_9538);
and U10283 (N_10283,N_9711,N_9592);
nand U10284 (N_10284,N_9981,N_9530);
nor U10285 (N_10285,N_9766,N_9595);
nand U10286 (N_10286,N_9972,N_9997);
nand U10287 (N_10287,N_9630,N_9603);
and U10288 (N_10288,N_9661,N_9974);
nand U10289 (N_10289,N_9501,N_9779);
and U10290 (N_10290,N_9651,N_9564);
xor U10291 (N_10291,N_9663,N_9608);
nor U10292 (N_10292,N_9737,N_9972);
xor U10293 (N_10293,N_9521,N_9817);
xnor U10294 (N_10294,N_9855,N_9967);
nand U10295 (N_10295,N_9589,N_9918);
xnor U10296 (N_10296,N_9763,N_9601);
nor U10297 (N_10297,N_9582,N_9913);
nand U10298 (N_10298,N_9628,N_9867);
nor U10299 (N_10299,N_9728,N_9983);
and U10300 (N_10300,N_9521,N_9795);
xor U10301 (N_10301,N_9705,N_9967);
and U10302 (N_10302,N_9748,N_9575);
and U10303 (N_10303,N_9851,N_9764);
or U10304 (N_10304,N_9563,N_9928);
and U10305 (N_10305,N_9562,N_9547);
nand U10306 (N_10306,N_9878,N_9593);
xor U10307 (N_10307,N_9988,N_9950);
nand U10308 (N_10308,N_9719,N_9656);
nand U10309 (N_10309,N_9897,N_9684);
and U10310 (N_10310,N_9628,N_9826);
nor U10311 (N_10311,N_9882,N_9814);
nand U10312 (N_10312,N_9589,N_9657);
and U10313 (N_10313,N_9996,N_9756);
and U10314 (N_10314,N_9725,N_9719);
or U10315 (N_10315,N_9911,N_9763);
or U10316 (N_10316,N_9644,N_9849);
nor U10317 (N_10317,N_9691,N_9684);
and U10318 (N_10318,N_9684,N_9878);
nor U10319 (N_10319,N_9959,N_9791);
or U10320 (N_10320,N_9911,N_9624);
xnor U10321 (N_10321,N_9801,N_9535);
or U10322 (N_10322,N_9513,N_9774);
or U10323 (N_10323,N_9783,N_9602);
nand U10324 (N_10324,N_9635,N_9928);
or U10325 (N_10325,N_9687,N_9618);
nor U10326 (N_10326,N_9658,N_9861);
xor U10327 (N_10327,N_9983,N_9677);
nor U10328 (N_10328,N_9650,N_9707);
or U10329 (N_10329,N_9981,N_9892);
xnor U10330 (N_10330,N_9673,N_9882);
nand U10331 (N_10331,N_9855,N_9730);
nand U10332 (N_10332,N_9590,N_9887);
nand U10333 (N_10333,N_9976,N_9831);
or U10334 (N_10334,N_9746,N_9541);
and U10335 (N_10335,N_9609,N_9840);
and U10336 (N_10336,N_9518,N_9785);
nor U10337 (N_10337,N_9569,N_9574);
xnor U10338 (N_10338,N_9625,N_9519);
and U10339 (N_10339,N_9734,N_9818);
xor U10340 (N_10340,N_9845,N_9927);
xnor U10341 (N_10341,N_9834,N_9633);
xor U10342 (N_10342,N_9779,N_9598);
nand U10343 (N_10343,N_9846,N_9541);
or U10344 (N_10344,N_9744,N_9801);
or U10345 (N_10345,N_9699,N_9997);
nor U10346 (N_10346,N_9774,N_9791);
xor U10347 (N_10347,N_9683,N_9909);
or U10348 (N_10348,N_9635,N_9958);
nand U10349 (N_10349,N_9634,N_9995);
and U10350 (N_10350,N_9620,N_9596);
nor U10351 (N_10351,N_9601,N_9895);
or U10352 (N_10352,N_9737,N_9901);
nor U10353 (N_10353,N_9886,N_9974);
nand U10354 (N_10354,N_9746,N_9919);
nand U10355 (N_10355,N_9943,N_9884);
nand U10356 (N_10356,N_9595,N_9610);
nand U10357 (N_10357,N_9682,N_9970);
xnor U10358 (N_10358,N_9842,N_9610);
xnor U10359 (N_10359,N_9947,N_9723);
xnor U10360 (N_10360,N_9947,N_9640);
and U10361 (N_10361,N_9815,N_9774);
nand U10362 (N_10362,N_9868,N_9896);
nor U10363 (N_10363,N_9819,N_9652);
or U10364 (N_10364,N_9813,N_9550);
or U10365 (N_10365,N_9752,N_9665);
and U10366 (N_10366,N_9898,N_9535);
nor U10367 (N_10367,N_9784,N_9988);
xnor U10368 (N_10368,N_9705,N_9618);
xor U10369 (N_10369,N_9854,N_9635);
nor U10370 (N_10370,N_9993,N_9827);
and U10371 (N_10371,N_9645,N_9807);
nor U10372 (N_10372,N_9727,N_9516);
and U10373 (N_10373,N_9892,N_9944);
nand U10374 (N_10374,N_9738,N_9753);
and U10375 (N_10375,N_9631,N_9676);
and U10376 (N_10376,N_9555,N_9740);
nand U10377 (N_10377,N_9657,N_9901);
and U10378 (N_10378,N_9737,N_9665);
or U10379 (N_10379,N_9547,N_9835);
nor U10380 (N_10380,N_9531,N_9597);
and U10381 (N_10381,N_9986,N_9729);
xor U10382 (N_10382,N_9969,N_9780);
nand U10383 (N_10383,N_9891,N_9531);
nor U10384 (N_10384,N_9570,N_9780);
nor U10385 (N_10385,N_9788,N_9565);
or U10386 (N_10386,N_9653,N_9929);
nand U10387 (N_10387,N_9919,N_9698);
xor U10388 (N_10388,N_9722,N_9505);
nand U10389 (N_10389,N_9594,N_9679);
and U10390 (N_10390,N_9981,N_9927);
nand U10391 (N_10391,N_9638,N_9688);
nor U10392 (N_10392,N_9661,N_9522);
nand U10393 (N_10393,N_9809,N_9615);
nor U10394 (N_10394,N_9650,N_9866);
nand U10395 (N_10395,N_9589,N_9635);
or U10396 (N_10396,N_9808,N_9933);
xnor U10397 (N_10397,N_9571,N_9707);
xor U10398 (N_10398,N_9979,N_9956);
nand U10399 (N_10399,N_9817,N_9793);
or U10400 (N_10400,N_9655,N_9519);
xor U10401 (N_10401,N_9984,N_9866);
nand U10402 (N_10402,N_9536,N_9765);
xnor U10403 (N_10403,N_9906,N_9723);
nor U10404 (N_10404,N_9783,N_9820);
or U10405 (N_10405,N_9907,N_9553);
nor U10406 (N_10406,N_9613,N_9519);
xor U10407 (N_10407,N_9652,N_9999);
and U10408 (N_10408,N_9834,N_9978);
or U10409 (N_10409,N_9836,N_9993);
nand U10410 (N_10410,N_9610,N_9879);
xnor U10411 (N_10411,N_9905,N_9972);
and U10412 (N_10412,N_9604,N_9805);
xnor U10413 (N_10413,N_9940,N_9820);
and U10414 (N_10414,N_9650,N_9841);
nand U10415 (N_10415,N_9715,N_9678);
and U10416 (N_10416,N_9630,N_9898);
nor U10417 (N_10417,N_9751,N_9959);
and U10418 (N_10418,N_9578,N_9912);
nor U10419 (N_10419,N_9593,N_9684);
nor U10420 (N_10420,N_9803,N_9852);
and U10421 (N_10421,N_9972,N_9832);
or U10422 (N_10422,N_9933,N_9711);
or U10423 (N_10423,N_9693,N_9509);
xor U10424 (N_10424,N_9909,N_9942);
nor U10425 (N_10425,N_9558,N_9758);
nand U10426 (N_10426,N_9932,N_9663);
nor U10427 (N_10427,N_9688,N_9912);
and U10428 (N_10428,N_9942,N_9548);
nand U10429 (N_10429,N_9640,N_9925);
xor U10430 (N_10430,N_9553,N_9892);
or U10431 (N_10431,N_9526,N_9960);
xor U10432 (N_10432,N_9545,N_9587);
and U10433 (N_10433,N_9993,N_9612);
xnor U10434 (N_10434,N_9933,N_9602);
nor U10435 (N_10435,N_9527,N_9580);
nor U10436 (N_10436,N_9634,N_9977);
or U10437 (N_10437,N_9514,N_9662);
nor U10438 (N_10438,N_9544,N_9525);
xor U10439 (N_10439,N_9629,N_9840);
or U10440 (N_10440,N_9995,N_9521);
nand U10441 (N_10441,N_9922,N_9909);
nor U10442 (N_10442,N_9713,N_9677);
and U10443 (N_10443,N_9662,N_9726);
nand U10444 (N_10444,N_9843,N_9774);
nand U10445 (N_10445,N_9785,N_9633);
and U10446 (N_10446,N_9830,N_9730);
xor U10447 (N_10447,N_9644,N_9669);
xor U10448 (N_10448,N_9813,N_9884);
nor U10449 (N_10449,N_9654,N_9653);
xor U10450 (N_10450,N_9622,N_9918);
nor U10451 (N_10451,N_9620,N_9785);
nand U10452 (N_10452,N_9980,N_9567);
nand U10453 (N_10453,N_9666,N_9852);
nand U10454 (N_10454,N_9576,N_9811);
and U10455 (N_10455,N_9689,N_9840);
or U10456 (N_10456,N_9719,N_9806);
xnor U10457 (N_10457,N_9882,N_9538);
or U10458 (N_10458,N_9597,N_9857);
and U10459 (N_10459,N_9976,N_9541);
nand U10460 (N_10460,N_9853,N_9890);
nor U10461 (N_10461,N_9907,N_9916);
nor U10462 (N_10462,N_9957,N_9747);
nand U10463 (N_10463,N_9879,N_9944);
or U10464 (N_10464,N_9623,N_9749);
or U10465 (N_10465,N_9623,N_9581);
or U10466 (N_10466,N_9815,N_9552);
xnor U10467 (N_10467,N_9662,N_9641);
nor U10468 (N_10468,N_9500,N_9824);
nand U10469 (N_10469,N_9553,N_9711);
xnor U10470 (N_10470,N_9786,N_9993);
and U10471 (N_10471,N_9789,N_9521);
or U10472 (N_10472,N_9936,N_9923);
or U10473 (N_10473,N_9720,N_9765);
or U10474 (N_10474,N_9640,N_9888);
or U10475 (N_10475,N_9683,N_9695);
and U10476 (N_10476,N_9873,N_9992);
or U10477 (N_10477,N_9601,N_9624);
or U10478 (N_10478,N_9918,N_9776);
or U10479 (N_10479,N_9628,N_9602);
nor U10480 (N_10480,N_9772,N_9684);
xor U10481 (N_10481,N_9735,N_9867);
nor U10482 (N_10482,N_9547,N_9777);
nand U10483 (N_10483,N_9723,N_9736);
nand U10484 (N_10484,N_9760,N_9572);
nor U10485 (N_10485,N_9636,N_9626);
or U10486 (N_10486,N_9518,N_9641);
xor U10487 (N_10487,N_9692,N_9959);
xor U10488 (N_10488,N_9879,N_9775);
nand U10489 (N_10489,N_9990,N_9852);
nand U10490 (N_10490,N_9564,N_9871);
nand U10491 (N_10491,N_9578,N_9941);
xor U10492 (N_10492,N_9897,N_9584);
and U10493 (N_10493,N_9884,N_9648);
or U10494 (N_10494,N_9503,N_9801);
nand U10495 (N_10495,N_9682,N_9720);
nor U10496 (N_10496,N_9652,N_9562);
nand U10497 (N_10497,N_9770,N_9672);
nand U10498 (N_10498,N_9541,N_9908);
or U10499 (N_10499,N_9772,N_9755);
nand U10500 (N_10500,N_10205,N_10176);
nor U10501 (N_10501,N_10479,N_10024);
and U10502 (N_10502,N_10227,N_10251);
and U10503 (N_10503,N_10337,N_10464);
or U10504 (N_10504,N_10491,N_10015);
and U10505 (N_10505,N_10173,N_10234);
or U10506 (N_10506,N_10013,N_10331);
or U10507 (N_10507,N_10177,N_10070);
nand U10508 (N_10508,N_10079,N_10091);
nand U10509 (N_10509,N_10436,N_10489);
xor U10510 (N_10510,N_10414,N_10295);
or U10511 (N_10511,N_10154,N_10165);
or U10512 (N_10512,N_10032,N_10223);
nor U10513 (N_10513,N_10408,N_10190);
and U10514 (N_10514,N_10422,N_10049);
and U10515 (N_10515,N_10369,N_10439);
nand U10516 (N_10516,N_10306,N_10314);
nand U10517 (N_10517,N_10022,N_10143);
and U10518 (N_10518,N_10092,N_10344);
and U10519 (N_10519,N_10480,N_10304);
xnor U10520 (N_10520,N_10420,N_10158);
xnor U10521 (N_10521,N_10048,N_10267);
nor U10522 (N_10522,N_10229,N_10359);
nand U10523 (N_10523,N_10381,N_10351);
nor U10524 (N_10524,N_10276,N_10279);
nand U10525 (N_10525,N_10488,N_10492);
nand U10526 (N_10526,N_10148,N_10121);
nand U10527 (N_10527,N_10493,N_10478);
nor U10528 (N_10528,N_10313,N_10191);
nor U10529 (N_10529,N_10224,N_10084);
nor U10530 (N_10530,N_10060,N_10250);
and U10531 (N_10531,N_10253,N_10130);
and U10532 (N_10532,N_10243,N_10118);
nor U10533 (N_10533,N_10355,N_10244);
and U10534 (N_10534,N_10090,N_10261);
and U10535 (N_10535,N_10281,N_10147);
nor U10536 (N_10536,N_10323,N_10058);
xnor U10537 (N_10537,N_10256,N_10135);
nor U10538 (N_10538,N_10132,N_10394);
or U10539 (N_10539,N_10160,N_10405);
and U10540 (N_10540,N_10000,N_10496);
and U10541 (N_10541,N_10425,N_10172);
xnor U10542 (N_10542,N_10231,N_10141);
and U10543 (N_10543,N_10477,N_10003);
nor U10544 (N_10544,N_10164,N_10076);
and U10545 (N_10545,N_10282,N_10393);
or U10546 (N_10546,N_10499,N_10124);
nor U10547 (N_10547,N_10265,N_10109);
or U10548 (N_10548,N_10202,N_10389);
and U10549 (N_10549,N_10407,N_10081);
nand U10550 (N_10550,N_10221,N_10378);
or U10551 (N_10551,N_10290,N_10072);
or U10552 (N_10552,N_10459,N_10482);
or U10553 (N_10553,N_10208,N_10150);
nor U10554 (N_10554,N_10106,N_10370);
and U10555 (N_10555,N_10009,N_10317);
and U10556 (N_10556,N_10367,N_10028);
xor U10557 (N_10557,N_10428,N_10174);
and U10558 (N_10558,N_10366,N_10376);
and U10559 (N_10559,N_10123,N_10430);
nor U10560 (N_10560,N_10192,N_10495);
and U10561 (N_10561,N_10036,N_10194);
and U10562 (N_10562,N_10320,N_10324);
and U10563 (N_10563,N_10001,N_10211);
xor U10564 (N_10564,N_10062,N_10218);
or U10565 (N_10565,N_10181,N_10475);
xnor U10566 (N_10566,N_10441,N_10128);
xnor U10567 (N_10567,N_10247,N_10263);
nand U10568 (N_10568,N_10305,N_10277);
and U10569 (N_10569,N_10350,N_10102);
and U10570 (N_10570,N_10008,N_10392);
xnor U10571 (N_10571,N_10063,N_10472);
or U10572 (N_10572,N_10122,N_10451);
nor U10573 (N_10573,N_10363,N_10240);
nor U10574 (N_10574,N_10438,N_10080);
nor U10575 (N_10575,N_10075,N_10326);
nand U10576 (N_10576,N_10409,N_10110);
or U10577 (N_10577,N_10435,N_10384);
or U10578 (N_10578,N_10342,N_10108);
nand U10579 (N_10579,N_10179,N_10166);
or U10580 (N_10580,N_10497,N_10415);
or U10581 (N_10581,N_10364,N_10426);
or U10582 (N_10582,N_10115,N_10171);
xor U10583 (N_10583,N_10259,N_10198);
and U10584 (N_10584,N_10039,N_10440);
and U10585 (N_10585,N_10446,N_10292);
or U10586 (N_10586,N_10054,N_10453);
or U10587 (N_10587,N_10059,N_10434);
or U10588 (N_10588,N_10483,N_10269);
nand U10589 (N_10589,N_10383,N_10225);
nand U10590 (N_10590,N_10254,N_10200);
nand U10591 (N_10591,N_10026,N_10053);
nand U10592 (N_10592,N_10233,N_10466);
or U10593 (N_10593,N_10377,N_10444);
nor U10594 (N_10594,N_10429,N_10449);
or U10595 (N_10595,N_10380,N_10236);
nand U10596 (N_10596,N_10155,N_10016);
and U10597 (N_10597,N_10352,N_10066);
or U10598 (N_10598,N_10291,N_10460);
nand U10599 (N_10599,N_10338,N_10113);
xnor U10600 (N_10600,N_10268,N_10417);
and U10601 (N_10601,N_10458,N_10461);
nand U10602 (N_10602,N_10217,N_10385);
nand U10603 (N_10603,N_10086,N_10206);
xor U10604 (N_10604,N_10213,N_10073);
or U10605 (N_10605,N_10368,N_10178);
xor U10606 (N_10606,N_10120,N_10209);
nand U10607 (N_10607,N_10180,N_10140);
nand U10608 (N_10608,N_10283,N_10195);
and U10609 (N_10609,N_10159,N_10299);
or U10610 (N_10610,N_10294,N_10356);
or U10611 (N_10611,N_10322,N_10134);
or U10612 (N_10612,N_10144,N_10035);
and U10613 (N_10613,N_10149,N_10327);
nor U10614 (N_10614,N_10427,N_10406);
nand U10615 (N_10615,N_10288,N_10196);
nor U10616 (N_10616,N_10473,N_10471);
nand U10617 (N_10617,N_10232,N_10151);
xnor U10618 (N_10618,N_10249,N_10457);
nor U10619 (N_10619,N_10278,N_10310);
xnor U10620 (N_10620,N_10474,N_10127);
or U10621 (N_10621,N_10280,N_10012);
and U10622 (N_10622,N_10333,N_10235);
xnor U10623 (N_10623,N_10052,N_10416);
or U10624 (N_10624,N_10152,N_10345);
nand U10625 (N_10625,N_10004,N_10002);
xnor U10626 (N_10626,N_10237,N_10145);
nand U10627 (N_10627,N_10442,N_10131);
nand U10628 (N_10628,N_10038,N_10047);
nand U10629 (N_10629,N_10014,N_10271);
xnor U10630 (N_10630,N_10321,N_10498);
nand U10631 (N_10631,N_10481,N_10252);
xor U10632 (N_10632,N_10034,N_10401);
nand U10633 (N_10633,N_10199,N_10193);
nor U10634 (N_10634,N_10156,N_10297);
or U10635 (N_10635,N_10167,N_10273);
nor U10636 (N_10636,N_10094,N_10411);
and U10637 (N_10637,N_10400,N_10228);
nor U10638 (N_10638,N_10107,N_10117);
or U10639 (N_10639,N_10007,N_10289);
and U10640 (N_10640,N_10391,N_10074);
xor U10641 (N_10641,N_10037,N_10216);
nor U10642 (N_10642,N_10431,N_10387);
nand U10643 (N_10643,N_10349,N_10095);
nand U10644 (N_10644,N_10332,N_10146);
nor U10645 (N_10645,N_10089,N_10258);
or U10646 (N_10646,N_10319,N_10085);
nor U10647 (N_10647,N_10046,N_10067);
or U10648 (N_10648,N_10051,N_10129);
and U10649 (N_10649,N_10412,N_10230);
nand U10650 (N_10650,N_10097,N_10125);
and U10651 (N_10651,N_10114,N_10303);
xor U10652 (N_10652,N_10104,N_10403);
nand U10653 (N_10653,N_10215,N_10182);
and U10654 (N_10654,N_10043,N_10365);
or U10655 (N_10655,N_10347,N_10287);
nor U10656 (N_10656,N_10162,N_10111);
xnor U10657 (N_10657,N_10126,N_10161);
or U10658 (N_10658,N_10203,N_10274);
nor U10659 (N_10659,N_10087,N_10424);
and U10660 (N_10660,N_10284,N_10465);
or U10661 (N_10661,N_10476,N_10248);
or U10662 (N_10662,N_10470,N_10157);
nand U10663 (N_10663,N_10329,N_10204);
nand U10664 (N_10664,N_10357,N_10302);
xor U10665 (N_10665,N_10241,N_10170);
nand U10666 (N_10666,N_10005,N_10098);
nand U10667 (N_10667,N_10031,N_10375);
nand U10668 (N_10668,N_10336,N_10023);
and U10669 (N_10669,N_10116,N_10275);
nor U10670 (N_10670,N_10340,N_10325);
or U10671 (N_10671,N_10018,N_10398);
nor U10672 (N_10672,N_10348,N_10169);
xnor U10673 (N_10673,N_10040,N_10207);
or U10674 (N_10674,N_10186,N_10119);
nand U10675 (N_10675,N_10112,N_10335);
nand U10676 (N_10676,N_10137,N_10272);
or U10677 (N_10677,N_10021,N_10153);
and U10678 (N_10678,N_10055,N_10133);
nand U10679 (N_10679,N_10316,N_10242);
and U10680 (N_10680,N_10006,N_10168);
nand U10681 (N_10681,N_10358,N_10450);
xor U10682 (N_10682,N_10390,N_10360);
nand U10683 (N_10683,N_10270,N_10136);
nand U10684 (N_10684,N_10257,N_10219);
nand U10685 (N_10685,N_10455,N_10262);
xnor U10686 (N_10686,N_10056,N_10373);
xor U10687 (N_10687,N_10068,N_10078);
xnor U10688 (N_10688,N_10309,N_10293);
and U10689 (N_10689,N_10286,N_10315);
nand U10690 (N_10690,N_10341,N_10307);
xor U10691 (N_10691,N_10064,N_10372);
nand U10692 (N_10692,N_10183,N_10246);
nand U10693 (N_10693,N_10020,N_10044);
xnor U10694 (N_10694,N_10027,N_10017);
nor U10695 (N_10695,N_10395,N_10041);
xor U10696 (N_10696,N_10245,N_10445);
nand U10697 (N_10697,N_10421,N_10197);
nor U10698 (N_10698,N_10462,N_10402);
or U10699 (N_10699,N_10328,N_10099);
or U10700 (N_10700,N_10486,N_10346);
or U10701 (N_10701,N_10362,N_10033);
or U10702 (N_10702,N_10030,N_10071);
xor U10703 (N_10703,N_10399,N_10065);
nand U10704 (N_10704,N_10404,N_10184);
nor U10705 (N_10705,N_10238,N_10410);
nand U10706 (N_10706,N_10214,N_10226);
and U10707 (N_10707,N_10494,N_10388);
or U10708 (N_10708,N_10485,N_10361);
or U10709 (N_10709,N_10487,N_10308);
or U10710 (N_10710,N_10334,N_10469);
and U10711 (N_10711,N_10300,N_10083);
or U10712 (N_10712,N_10201,N_10019);
and U10713 (N_10713,N_10452,N_10266);
nand U10714 (N_10714,N_10057,N_10011);
nand U10715 (N_10715,N_10354,N_10285);
nand U10716 (N_10716,N_10353,N_10301);
xnor U10717 (N_10717,N_10396,N_10382);
or U10718 (N_10718,N_10330,N_10397);
nor U10719 (N_10719,N_10210,N_10189);
or U10720 (N_10720,N_10082,N_10413);
xor U10721 (N_10721,N_10433,N_10318);
nand U10722 (N_10722,N_10448,N_10418);
or U10723 (N_10723,N_10490,N_10185);
or U10724 (N_10724,N_10222,N_10187);
and U10725 (N_10725,N_10042,N_10386);
nor U10726 (N_10726,N_10220,N_10175);
or U10727 (N_10727,N_10103,N_10050);
and U10728 (N_10728,N_10463,N_10096);
nor U10729 (N_10729,N_10025,N_10105);
nand U10730 (N_10730,N_10010,N_10454);
and U10731 (N_10731,N_10077,N_10423);
nor U10732 (N_10732,N_10100,N_10069);
or U10733 (N_10733,N_10374,N_10142);
xnor U10734 (N_10734,N_10061,N_10468);
nand U10735 (N_10735,N_10371,N_10264);
nand U10736 (N_10736,N_10379,N_10296);
nor U10737 (N_10737,N_10484,N_10212);
or U10738 (N_10738,N_10447,N_10312);
xor U10739 (N_10739,N_10139,N_10432);
nor U10740 (N_10740,N_10443,N_10101);
nand U10741 (N_10741,N_10188,N_10255);
and U10742 (N_10742,N_10088,N_10260);
or U10743 (N_10743,N_10298,N_10343);
and U10744 (N_10744,N_10419,N_10239);
or U10745 (N_10745,N_10029,N_10311);
nor U10746 (N_10746,N_10456,N_10339);
xnor U10747 (N_10747,N_10163,N_10138);
nand U10748 (N_10748,N_10437,N_10093);
and U10749 (N_10749,N_10467,N_10045);
and U10750 (N_10750,N_10127,N_10115);
nand U10751 (N_10751,N_10398,N_10145);
xnor U10752 (N_10752,N_10424,N_10097);
and U10753 (N_10753,N_10006,N_10128);
and U10754 (N_10754,N_10198,N_10081);
nand U10755 (N_10755,N_10385,N_10303);
nor U10756 (N_10756,N_10163,N_10207);
and U10757 (N_10757,N_10437,N_10046);
or U10758 (N_10758,N_10457,N_10221);
nor U10759 (N_10759,N_10194,N_10046);
nand U10760 (N_10760,N_10305,N_10002);
xnor U10761 (N_10761,N_10008,N_10290);
and U10762 (N_10762,N_10164,N_10252);
or U10763 (N_10763,N_10076,N_10248);
nand U10764 (N_10764,N_10289,N_10301);
xor U10765 (N_10765,N_10032,N_10194);
or U10766 (N_10766,N_10295,N_10175);
nor U10767 (N_10767,N_10233,N_10442);
nor U10768 (N_10768,N_10089,N_10493);
nand U10769 (N_10769,N_10161,N_10281);
nor U10770 (N_10770,N_10414,N_10109);
xor U10771 (N_10771,N_10447,N_10477);
nor U10772 (N_10772,N_10479,N_10125);
nor U10773 (N_10773,N_10342,N_10493);
nor U10774 (N_10774,N_10018,N_10277);
nor U10775 (N_10775,N_10373,N_10396);
nor U10776 (N_10776,N_10033,N_10480);
nor U10777 (N_10777,N_10075,N_10486);
xnor U10778 (N_10778,N_10488,N_10155);
or U10779 (N_10779,N_10389,N_10310);
or U10780 (N_10780,N_10322,N_10395);
nor U10781 (N_10781,N_10187,N_10435);
nor U10782 (N_10782,N_10000,N_10350);
and U10783 (N_10783,N_10253,N_10128);
xor U10784 (N_10784,N_10031,N_10477);
or U10785 (N_10785,N_10196,N_10119);
and U10786 (N_10786,N_10111,N_10074);
nor U10787 (N_10787,N_10109,N_10471);
nand U10788 (N_10788,N_10454,N_10175);
and U10789 (N_10789,N_10432,N_10023);
and U10790 (N_10790,N_10292,N_10040);
or U10791 (N_10791,N_10343,N_10112);
or U10792 (N_10792,N_10236,N_10353);
nor U10793 (N_10793,N_10045,N_10143);
xnor U10794 (N_10794,N_10474,N_10441);
or U10795 (N_10795,N_10381,N_10086);
nand U10796 (N_10796,N_10039,N_10400);
and U10797 (N_10797,N_10036,N_10380);
nor U10798 (N_10798,N_10304,N_10351);
nand U10799 (N_10799,N_10075,N_10372);
or U10800 (N_10800,N_10093,N_10385);
xnor U10801 (N_10801,N_10418,N_10447);
nand U10802 (N_10802,N_10141,N_10117);
xnor U10803 (N_10803,N_10137,N_10250);
and U10804 (N_10804,N_10101,N_10099);
or U10805 (N_10805,N_10433,N_10443);
nor U10806 (N_10806,N_10378,N_10184);
nor U10807 (N_10807,N_10209,N_10499);
and U10808 (N_10808,N_10305,N_10061);
nand U10809 (N_10809,N_10074,N_10394);
xnor U10810 (N_10810,N_10035,N_10354);
nand U10811 (N_10811,N_10468,N_10461);
nand U10812 (N_10812,N_10040,N_10271);
and U10813 (N_10813,N_10425,N_10473);
nor U10814 (N_10814,N_10407,N_10360);
nor U10815 (N_10815,N_10242,N_10473);
or U10816 (N_10816,N_10158,N_10099);
nor U10817 (N_10817,N_10401,N_10022);
nand U10818 (N_10818,N_10378,N_10413);
nor U10819 (N_10819,N_10180,N_10470);
nor U10820 (N_10820,N_10112,N_10472);
or U10821 (N_10821,N_10291,N_10002);
nand U10822 (N_10822,N_10125,N_10293);
or U10823 (N_10823,N_10077,N_10185);
and U10824 (N_10824,N_10451,N_10358);
nand U10825 (N_10825,N_10263,N_10077);
nand U10826 (N_10826,N_10069,N_10348);
xnor U10827 (N_10827,N_10328,N_10348);
nand U10828 (N_10828,N_10312,N_10162);
and U10829 (N_10829,N_10446,N_10209);
nor U10830 (N_10830,N_10142,N_10047);
nand U10831 (N_10831,N_10200,N_10327);
nand U10832 (N_10832,N_10015,N_10149);
or U10833 (N_10833,N_10129,N_10126);
nor U10834 (N_10834,N_10396,N_10175);
xnor U10835 (N_10835,N_10225,N_10388);
xor U10836 (N_10836,N_10033,N_10355);
xor U10837 (N_10837,N_10135,N_10163);
nor U10838 (N_10838,N_10276,N_10351);
nand U10839 (N_10839,N_10060,N_10195);
or U10840 (N_10840,N_10387,N_10269);
nand U10841 (N_10841,N_10079,N_10430);
or U10842 (N_10842,N_10477,N_10259);
xnor U10843 (N_10843,N_10460,N_10177);
and U10844 (N_10844,N_10100,N_10320);
nand U10845 (N_10845,N_10495,N_10247);
and U10846 (N_10846,N_10051,N_10029);
nand U10847 (N_10847,N_10280,N_10141);
or U10848 (N_10848,N_10370,N_10250);
nand U10849 (N_10849,N_10451,N_10391);
or U10850 (N_10850,N_10017,N_10107);
or U10851 (N_10851,N_10198,N_10327);
and U10852 (N_10852,N_10140,N_10488);
xnor U10853 (N_10853,N_10349,N_10007);
xor U10854 (N_10854,N_10163,N_10489);
nor U10855 (N_10855,N_10262,N_10001);
nor U10856 (N_10856,N_10153,N_10395);
nor U10857 (N_10857,N_10329,N_10317);
xnor U10858 (N_10858,N_10152,N_10491);
nand U10859 (N_10859,N_10485,N_10120);
nor U10860 (N_10860,N_10386,N_10388);
nand U10861 (N_10861,N_10169,N_10223);
nand U10862 (N_10862,N_10361,N_10304);
nand U10863 (N_10863,N_10408,N_10102);
and U10864 (N_10864,N_10112,N_10236);
or U10865 (N_10865,N_10047,N_10318);
xor U10866 (N_10866,N_10130,N_10254);
or U10867 (N_10867,N_10160,N_10318);
xnor U10868 (N_10868,N_10072,N_10111);
xor U10869 (N_10869,N_10090,N_10294);
or U10870 (N_10870,N_10031,N_10460);
nand U10871 (N_10871,N_10262,N_10263);
nor U10872 (N_10872,N_10449,N_10210);
or U10873 (N_10873,N_10415,N_10466);
nand U10874 (N_10874,N_10213,N_10390);
or U10875 (N_10875,N_10431,N_10446);
or U10876 (N_10876,N_10335,N_10411);
xnor U10877 (N_10877,N_10165,N_10484);
or U10878 (N_10878,N_10238,N_10439);
nor U10879 (N_10879,N_10382,N_10471);
or U10880 (N_10880,N_10144,N_10118);
or U10881 (N_10881,N_10072,N_10115);
or U10882 (N_10882,N_10199,N_10198);
nor U10883 (N_10883,N_10351,N_10355);
xnor U10884 (N_10884,N_10088,N_10183);
and U10885 (N_10885,N_10079,N_10152);
xor U10886 (N_10886,N_10426,N_10448);
or U10887 (N_10887,N_10041,N_10106);
nand U10888 (N_10888,N_10404,N_10357);
or U10889 (N_10889,N_10271,N_10155);
nand U10890 (N_10890,N_10201,N_10054);
nor U10891 (N_10891,N_10077,N_10252);
and U10892 (N_10892,N_10187,N_10328);
and U10893 (N_10893,N_10455,N_10147);
or U10894 (N_10894,N_10114,N_10283);
and U10895 (N_10895,N_10296,N_10396);
nor U10896 (N_10896,N_10308,N_10115);
xor U10897 (N_10897,N_10076,N_10433);
nand U10898 (N_10898,N_10385,N_10201);
nor U10899 (N_10899,N_10270,N_10382);
or U10900 (N_10900,N_10038,N_10049);
or U10901 (N_10901,N_10253,N_10313);
or U10902 (N_10902,N_10206,N_10088);
xnor U10903 (N_10903,N_10061,N_10183);
xnor U10904 (N_10904,N_10239,N_10411);
xnor U10905 (N_10905,N_10274,N_10128);
xor U10906 (N_10906,N_10239,N_10499);
nor U10907 (N_10907,N_10024,N_10068);
nor U10908 (N_10908,N_10199,N_10105);
nor U10909 (N_10909,N_10096,N_10012);
and U10910 (N_10910,N_10130,N_10121);
or U10911 (N_10911,N_10401,N_10172);
nand U10912 (N_10912,N_10182,N_10061);
nand U10913 (N_10913,N_10448,N_10052);
nor U10914 (N_10914,N_10194,N_10429);
xor U10915 (N_10915,N_10121,N_10232);
and U10916 (N_10916,N_10361,N_10034);
and U10917 (N_10917,N_10018,N_10427);
xnor U10918 (N_10918,N_10146,N_10461);
and U10919 (N_10919,N_10238,N_10296);
nand U10920 (N_10920,N_10416,N_10073);
or U10921 (N_10921,N_10202,N_10217);
or U10922 (N_10922,N_10350,N_10065);
or U10923 (N_10923,N_10021,N_10299);
nand U10924 (N_10924,N_10116,N_10394);
nand U10925 (N_10925,N_10170,N_10223);
xor U10926 (N_10926,N_10240,N_10274);
and U10927 (N_10927,N_10248,N_10466);
or U10928 (N_10928,N_10289,N_10356);
nand U10929 (N_10929,N_10470,N_10256);
nand U10930 (N_10930,N_10363,N_10277);
or U10931 (N_10931,N_10376,N_10170);
nand U10932 (N_10932,N_10444,N_10358);
and U10933 (N_10933,N_10401,N_10390);
nand U10934 (N_10934,N_10267,N_10123);
nand U10935 (N_10935,N_10368,N_10061);
nand U10936 (N_10936,N_10006,N_10218);
nand U10937 (N_10937,N_10060,N_10238);
nand U10938 (N_10938,N_10229,N_10141);
or U10939 (N_10939,N_10165,N_10285);
nand U10940 (N_10940,N_10243,N_10472);
and U10941 (N_10941,N_10312,N_10029);
nor U10942 (N_10942,N_10212,N_10060);
or U10943 (N_10943,N_10272,N_10453);
xor U10944 (N_10944,N_10200,N_10090);
nor U10945 (N_10945,N_10328,N_10135);
xnor U10946 (N_10946,N_10423,N_10195);
nand U10947 (N_10947,N_10476,N_10034);
nor U10948 (N_10948,N_10042,N_10058);
or U10949 (N_10949,N_10363,N_10294);
and U10950 (N_10950,N_10263,N_10469);
nor U10951 (N_10951,N_10448,N_10331);
nor U10952 (N_10952,N_10038,N_10445);
xnor U10953 (N_10953,N_10245,N_10144);
nand U10954 (N_10954,N_10380,N_10213);
or U10955 (N_10955,N_10351,N_10280);
and U10956 (N_10956,N_10333,N_10307);
and U10957 (N_10957,N_10028,N_10426);
nor U10958 (N_10958,N_10057,N_10063);
xnor U10959 (N_10959,N_10269,N_10337);
nor U10960 (N_10960,N_10184,N_10097);
and U10961 (N_10961,N_10288,N_10247);
nor U10962 (N_10962,N_10498,N_10276);
xnor U10963 (N_10963,N_10407,N_10153);
nor U10964 (N_10964,N_10498,N_10135);
nand U10965 (N_10965,N_10474,N_10480);
nor U10966 (N_10966,N_10018,N_10013);
nor U10967 (N_10967,N_10336,N_10382);
or U10968 (N_10968,N_10065,N_10024);
nand U10969 (N_10969,N_10434,N_10020);
and U10970 (N_10970,N_10429,N_10264);
nand U10971 (N_10971,N_10235,N_10200);
nand U10972 (N_10972,N_10403,N_10329);
and U10973 (N_10973,N_10241,N_10050);
nor U10974 (N_10974,N_10398,N_10058);
nor U10975 (N_10975,N_10040,N_10416);
nor U10976 (N_10976,N_10138,N_10489);
and U10977 (N_10977,N_10142,N_10144);
xnor U10978 (N_10978,N_10173,N_10190);
xor U10979 (N_10979,N_10162,N_10358);
nor U10980 (N_10980,N_10042,N_10471);
nand U10981 (N_10981,N_10293,N_10181);
xor U10982 (N_10982,N_10023,N_10266);
or U10983 (N_10983,N_10395,N_10212);
and U10984 (N_10984,N_10179,N_10312);
nor U10985 (N_10985,N_10385,N_10143);
and U10986 (N_10986,N_10317,N_10453);
or U10987 (N_10987,N_10297,N_10180);
and U10988 (N_10988,N_10236,N_10436);
nand U10989 (N_10989,N_10432,N_10143);
and U10990 (N_10990,N_10001,N_10269);
nand U10991 (N_10991,N_10421,N_10166);
nor U10992 (N_10992,N_10247,N_10173);
nor U10993 (N_10993,N_10467,N_10112);
or U10994 (N_10994,N_10444,N_10282);
xnor U10995 (N_10995,N_10358,N_10280);
nand U10996 (N_10996,N_10373,N_10077);
and U10997 (N_10997,N_10167,N_10469);
xnor U10998 (N_10998,N_10418,N_10280);
nor U10999 (N_10999,N_10287,N_10349);
xor U11000 (N_11000,N_10723,N_10581);
nor U11001 (N_11001,N_10923,N_10588);
nand U11002 (N_11002,N_10727,N_10880);
nand U11003 (N_11003,N_10770,N_10792);
xor U11004 (N_11004,N_10867,N_10715);
nand U11005 (N_11005,N_10992,N_10692);
nand U11006 (N_11006,N_10550,N_10736);
xnor U11007 (N_11007,N_10962,N_10531);
nor U11008 (N_11008,N_10985,N_10644);
and U11009 (N_11009,N_10946,N_10660);
nand U11010 (N_11010,N_10640,N_10824);
or U11011 (N_11011,N_10786,N_10895);
or U11012 (N_11012,N_10828,N_10500);
or U11013 (N_11013,N_10721,N_10939);
xnor U11014 (N_11014,N_10774,N_10998);
and U11015 (N_11015,N_10646,N_10604);
or U11016 (N_11016,N_10707,N_10822);
nor U11017 (N_11017,N_10871,N_10607);
nor U11018 (N_11018,N_10870,N_10806);
xnor U11019 (N_11019,N_10567,N_10613);
or U11020 (N_11020,N_10653,N_10526);
nor U11021 (N_11021,N_10893,N_10733);
and U11022 (N_11022,N_10502,N_10560);
nand U11023 (N_11023,N_10699,N_10573);
and U11024 (N_11024,N_10948,N_10817);
xnor U11025 (N_11025,N_10963,N_10790);
and U11026 (N_11026,N_10927,N_10802);
or U11027 (N_11027,N_10971,N_10685);
nand U11028 (N_11028,N_10979,N_10791);
nor U11029 (N_11029,N_10850,N_10695);
or U11030 (N_11030,N_10801,N_10796);
or U11031 (N_11031,N_10805,N_10689);
or U11032 (N_11032,N_10658,N_10576);
and U11033 (N_11033,N_10760,N_10600);
and U11034 (N_11034,N_10919,N_10914);
and U11035 (N_11035,N_10928,N_10631);
nand U11036 (N_11036,N_10930,N_10599);
and U11037 (N_11037,N_10512,N_10997);
nand U11038 (N_11038,N_10759,N_10652);
nor U11039 (N_11039,N_10524,N_10632);
nor U11040 (N_11040,N_10575,N_10837);
or U11041 (N_11041,N_10889,N_10712);
and U11042 (N_11042,N_10840,N_10857);
or U11043 (N_11043,N_10855,N_10702);
or U11044 (N_11044,N_10545,N_10908);
and U11045 (N_11045,N_10616,N_10982);
xnor U11046 (N_11046,N_10903,N_10884);
or U11047 (N_11047,N_10746,N_10785);
nor U11048 (N_11048,N_10834,N_10793);
or U11049 (N_11049,N_10947,N_10776);
nand U11050 (N_11050,N_10825,N_10700);
or U11051 (N_11051,N_10995,N_10758);
xnor U11052 (N_11052,N_10691,N_10964);
or U11053 (N_11053,N_10654,N_10641);
nor U11054 (N_11054,N_10735,N_10552);
nand U11055 (N_11055,N_10974,N_10940);
or U11056 (N_11056,N_10729,N_10628);
or U11057 (N_11057,N_10905,N_10566);
or U11058 (N_11058,N_10929,N_10590);
xor U11059 (N_11059,N_10909,N_10624);
or U11060 (N_11060,N_10858,N_10528);
nor U11061 (N_11061,N_10651,N_10775);
nor U11062 (N_11062,N_10559,N_10984);
xor U11063 (N_11063,N_10683,N_10856);
and U11064 (N_11064,N_10864,N_10745);
nand U11065 (N_11065,N_10619,N_10623);
nand U11066 (N_11066,N_10626,N_10782);
and U11067 (N_11067,N_10783,N_10584);
or U11068 (N_11068,N_10606,N_10541);
xor U11069 (N_11069,N_10739,N_10525);
xnor U11070 (N_11070,N_10708,N_10841);
or U11071 (N_11071,N_10907,N_10516);
nand U11072 (N_11072,N_10868,N_10517);
and U11073 (N_11073,N_10876,N_10612);
and U11074 (N_11074,N_10642,N_10961);
nor U11075 (N_11075,N_10582,N_10762);
xor U11076 (N_11076,N_10921,N_10682);
and U11077 (N_11077,N_10661,N_10798);
xor U11078 (N_11078,N_10922,N_10521);
nand U11079 (N_11079,N_10911,N_10593);
nand U11080 (N_11080,N_10953,N_10852);
nand U11081 (N_11081,N_10764,N_10788);
nand U11082 (N_11082,N_10585,N_10767);
xor U11083 (N_11083,N_10975,N_10527);
nand U11084 (N_11084,N_10650,N_10748);
xor U11085 (N_11085,N_10509,N_10618);
nor U11086 (N_11086,N_10558,N_10999);
nor U11087 (N_11087,N_10669,N_10950);
or U11088 (N_11088,N_10771,N_10981);
nor U11089 (N_11089,N_10565,N_10645);
xor U11090 (N_11090,N_10508,N_10711);
nand U11091 (N_11091,N_10554,N_10784);
nand U11092 (N_11092,N_10924,N_10693);
xor U11093 (N_11093,N_10761,N_10901);
or U11094 (N_11094,N_10752,N_10709);
nand U11095 (N_11095,N_10656,N_10958);
or U11096 (N_11096,N_10900,N_10842);
xor U11097 (N_11097,N_10913,N_10941);
and U11098 (N_11098,N_10781,N_10676);
nor U11099 (N_11099,N_10568,N_10863);
nand U11100 (N_11100,N_10996,N_10755);
xor U11101 (N_11101,N_10595,N_10569);
and U11102 (N_11102,N_10986,N_10978);
nor U11103 (N_11103,N_10869,N_10917);
or U11104 (N_11104,N_10583,N_10538);
nand U11105 (N_11105,N_10537,N_10637);
or U11106 (N_11106,N_10505,N_10865);
and U11107 (N_11107,N_10993,N_10605);
or U11108 (N_11108,N_10898,N_10885);
nand U11109 (N_11109,N_10714,N_10659);
and U11110 (N_11110,N_10534,N_10672);
nand U11111 (N_11111,N_10955,N_10926);
xnor U11112 (N_11112,N_10960,N_10813);
nor U11113 (N_11113,N_10596,N_10763);
nand U11114 (N_11114,N_10737,N_10747);
nand U11115 (N_11115,N_10899,N_10610);
and U11116 (N_11116,N_10779,N_10915);
nand U11117 (N_11117,N_10894,N_10906);
xor U11118 (N_11118,N_10670,N_10561);
or U11119 (N_11119,N_10777,N_10860);
nor U11120 (N_11120,N_10608,N_10601);
xor U11121 (N_11121,N_10831,N_10620);
xor U11122 (N_11122,N_10722,N_10968);
nand U11123 (N_11123,N_10592,N_10872);
nor U11124 (N_11124,N_10976,N_10814);
and U11125 (N_11125,N_10787,N_10598);
nor U11126 (N_11126,N_10826,N_10627);
nor U11127 (N_11127,N_10625,N_10875);
and U11128 (N_11128,N_10536,N_10851);
xnor U11129 (N_11129,N_10804,N_10674);
nor U11130 (N_11130,N_10757,N_10942);
and U11131 (N_11131,N_10795,N_10734);
or U11132 (N_11132,N_10819,N_10719);
nand U11133 (N_11133,N_10730,N_10551);
xor U11134 (N_11134,N_10529,N_10861);
xor U11135 (N_11135,N_10562,N_10713);
nor U11136 (N_11136,N_10935,N_10990);
or U11137 (N_11137,N_10701,N_10688);
nand U11138 (N_11138,N_10936,N_10879);
or U11139 (N_11139,N_10938,N_10706);
nand U11140 (N_11140,N_10543,N_10916);
xor U11141 (N_11141,N_10829,N_10518);
xor U11142 (N_11142,N_10987,N_10991);
xor U11143 (N_11143,N_10918,N_10671);
or U11144 (N_11144,N_10966,N_10769);
and U11145 (N_11145,N_10845,N_10920);
nor U11146 (N_11146,N_10535,N_10847);
nand U11147 (N_11147,N_10731,N_10718);
nand U11148 (N_11148,N_10883,N_10967);
xor U11149 (N_11149,N_10647,N_10952);
nor U11150 (N_11150,N_10836,N_10548);
or U11151 (N_11151,N_10511,N_10983);
or U11152 (N_11152,N_10663,N_10891);
xnor U11153 (N_11153,N_10902,N_10629);
and U11154 (N_11154,N_10820,N_10944);
nor U11155 (N_11155,N_10579,N_10896);
xor U11156 (N_11156,N_10611,N_10989);
and U11157 (N_11157,N_10556,N_10811);
nor U11158 (N_11158,N_10603,N_10680);
xor U11159 (N_11159,N_10705,N_10778);
xnor U11160 (N_11160,N_10725,N_10530);
nor U11161 (N_11161,N_10675,N_10686);
or U11162 (N_11162,N_10615,N_10533);
nor U11163 (N_11163,N_10614,N_10597);
xor U11164 (N_11164,N_10972,N_10666);
or U11165 (N_11165,N_10578,N_10827);
and U11166 (N_11166,N_10704,N_10980);
and U11167 (N_11167,N_10756,N_10807);
and U11168 (N_11168,N_10662,N_10882);
or U11169 (N_11169,N_10931,N_10854);
or U11170 (N_11170,N_10848,N_10766);
nand U11171 (N_11171,N_10667,N_10507);
nand U11172 (N_11172,N_10959,N_10513);
nor U11173 (N_11173,N_10504,N_10818);
nand U11174 (N_11174,N_10720,N_10639);
nor U11175 (N_11175,N_10634,N_10539);
and U11176 (N_11176,N_10749,N_10728);
nand U11177 (N_11177,N_10520,N_10859);
xor U11178 (N_11178,N_10553,N_10890);
nand U11179 (N_11179,N_10810,N_10892);
nand U11180 (N_11180,N_10910,N_10514);
and U11181 (N_11181,N_10542,N_10994);
xor U11182 (N_11182,N_10673,N_10503);
and U11183 (N_11183,N_10602,N_10874);
and U11184 (N_11184,N_10572,N_10949);
or U11185 (N_11185,N_10633,N_10717);
nand U11186 (N_11186,N_10988,N_10741);
and U11187 (N_11187,N_10544,N_10591);
and U11188 (N_11188,N_10594,N_10710);
nor U11189 (N_11189,N_10753,N_10951);
or U11190 (N_11190,N_10549,N_10956);
nand U11191 (N_11191,N_10933,N_10519);
nor U11192 (N_11192,N_10772,N_10510);
nor U11193 (N_11193,N_10703,N_10925);
nand U11194 (N_11194,N_10945,N_10580);
nor U11195 (N_11195,N_10934,N_10823);
or U11196 (N_11196,N_10743,N_10523);
or U11197 (N_11197,N_10977,N_10738);
nand U11198 (N_11198,N_10803,N_10835);
nand U11199 (N_11199,N_10833,N_10587);
xnor U11200 (N_11200,N_10904,N_10794);
nand U11201 (N_11201,N_10866,N_10888);
and U11202 (N_11202,N_10609,N_10522);
nor U11203 (N_11203,N_10873,N_10821);
xor U11204 (N_11204,N_10768,N_10638);
or U11205 (N_11205,N_10684,N_10844);
nor U11206 (N_11206,N_10532,N_10677);
xnor U11207 (N_11207,N_10809,N_10589);
or U11208 (N_11208,N_10577,N_10564);
nand U11209 (N_11209,N_10937,N_10681);
xor U11210 (N_11210,N_10732,N_10555);
and U11211 (N_11211,N_10954,N_10643);
and U11212 (N_11212,N_10546,N_10750);
nand U11213 (N_11213,N_10897,N_10832);
or U11214 (N_11214,N_10557,N_10698);
and U11215 (N_11215,N_10973,N_10797);
or U11216 (N_11216,N_10678,N_10815);
or U11217 (N_11217,N_10687,N_10515);
xor U11218 (N_11218,N_10586,N_10943);
or U11219 (N_11219,N_10696,N_10635);
nor U11220 (N_11220,N_10649,N_10657);
or U11221 (N_11221,N_10636,N_10780);
xor U11222 (N_11222,N_10668,N_10617);
nand U11223 (N_11223,N_10694,N_10800);
or U11224 (N_11224,N_10808,N_10970);
nand U11225 (N_11225,N_10740,N_10886);
nor U11226 (N_11226,N_10697,N_10839);
or U11227 (N_11227,N_10622,N_10690);
and U11228 (N_11228,N_10846,N_10816);
and U11229 (N_11229,N_10679,N_10773);
xnor U11230 (N_11230,N_10570,N_10621);
or U11231 (N_11231,N_10799,N_10754);
xnor U11232 (N_11232,N_10630,N_10665);
xnor U11233 (N_11233,N_10563,N_10838);
nand U11234 (N_11234,N_10969,N_10571);
nand U11235 (N_11235,N_10716,N_10932);
nand U11236 (N_11236,N_10843,N_10765);
nand U11237 (N_11237,N_10648,N_10878);
nand U11238 (N_11238,N_10506,N_10726);
or U11239 (N_11239,N_10830,N_10501);
nor U11240 (N_11240,N_10724,N_10812);
or U11241 (N_11241,N_10912,N_10965);
or U11242 (N_11242,N_10881,N_10664);
nand U11243 (N_11243,N_10849,N_10789);
nand U11244 (N_11244,N_10887,N_10862);
or U11245 (N_11245,N_10877,N_10540);
xnor U11246 (N_11246,N_10853,N_10957);
or U11247 (N_11247,N_10574,N_10655);
nor U11248 (N_11248,N_10744,N_10742);
xnor U11249 (N_11249,N_10751,N_10547);
or U11250 (N_11250,N_10904,N_10888);
nand U11251 (N_11251,N_10595,N_10870);
or U11252 (N_11252,N_10535,N_10667);
nor U11253 (N_11253,N_10764,N_10760);
xor U11254 (N_11254,N_10944,N_10881);
nand U11255 (N_11255,N_10671,N_10510);
nand U11256 (N_11256,N_10874,N_10768);
or U11257 (N_11257,N_10766,N_10715);
xor U11258 (N_11258,N_10607,N_10843);
xor U11259 (N_11259,N_10746,N_10591);
xor U11260 (N_11260,N_10954,N_10624);
xnor U11261 (N_11261,N_10657,N_10538);
nand U11262 (N_11262,N_10725,N_10976);
nand U11263 (N_11263,N_10804,N_10930);
nor U11264 (N_11264,N_10922,N_10749);
or U11265 (N_11265,N_10962,N_10663);
nor U11266 (N_11266,N_10936,N_10771);
or U11267 (N_11267,N_10523,N_10849);
or U11268 (N_11268,N_10823,N_10658);
nor U11269 (N_11269,N_10918,N_10667);
nand U11270 (N_11270,N_10589,N_10776);
and U11271 (N_11271,N_10630,N_10835);
or U11272 (N_11272,N_10701,N_10921);
xor U11273 (N_11273,N_10957,N_10997);
nand U11274 (N_11274,N_10723,N_10592);
nor U11275 (N_11275,N_10513,N_10835);
nand U11276 (N_11276,N_10796,N_10735);
nand U11277 (N_11277,N_10835,N_10677);
xor U11278 (N_11278,N_10524,N_10531);
xnor U11279 (N_11279,N_10574,N_10908);
xor U11280 (N_11280,N_10554,N_10856);
nand U11281 (N_11281,N_10791,N_10814);
nor U11282 (N_11282,N_10982,N_10952);
nor U11283 (N_11283,N_10721,N_10877);
nand U11284 (N_11284,N_10860,N_10993);
and U11285 (N_11285,N_10719,N_10588);
xnor U11286 (N_11286,N_10894,N_10540);
nor U11287 (N_11287,N_10839,N_10817);
xor U11288 (N_11288,N_10635,N_10585);
nand U11289 (N_11289,N_10861,N_10835);
or U11290 (N_11290,N_10646,N_10744);
or U11291 (N_11291,N_10825,N_10869);
and U11292 (N_11292,N_10985,N_10845);
and U11293 (N_11293,N_10842,N_10669);
nor U11294 (N_11294,N_10628,N_10603);
and U11295 (N_11295,N_10608,N_10849);
or U11296 (N_11296,N_10578,N_10597);
xnor U11297 (N_11297,N_10635,N_10623);
xor U11298 (N_11298,N_10649,N_10981);
nand U11299 (N_11299,N_10547,N_10629);
and U11300 (N_11300,N_10574,N_10703);
nand U11301 (N_11301,N_10682,N_10697);
nor U11302 (N_11302,N_10772,N_10737);
nand U11303 (N_11303,N_10938,N_10917);
or U11304 (N_11304,N_10568,N_10966);
or U11305 (N_11305,N_10986,N_10862);
nor U11306 (N_11306,N_10837,N_10565);
xnor U11307 (N_11307,N_10821,N_10871);
or U11308 (N_11308,N_10575,N_10689);
nand U11309 (N_11309,N_10543,N_10886);
nor U11310 (N_11310,N_10871,N_10635);
or U11311 (N_11311,N_10592,N_10704);
nand U11312 (N_11312,N_10835,N_10789);
xnor U11313 (N_11313,N_10660,N_10937);
or U11314 (N_11314,N_10960,N_10874);
or U11315 (N_11315,N_10502,N_10975);
nor U11316 (N_11316,N_10647,N_10887);
xnor U11317 (N_11317,N_10538,N_10706);
or U11318 (N_11318,N_10816,N_10533);
or U11319 (N_11319,N_10964,N_10954);
xnor U11320 (N_11320,N_10536,N_10935);
xor U11321 (N_11321,N_10961,N_10778);
nor U11322 (N_11322,N_10888,N_10846);
nor U11323 (N_11323,N_10786,N_10822);
xor U11324 (N_11324,N_10788,N_10666);
nor U11325 (N_11325,N_10756,N_10647);
xor U11326 (N_11326,N_10505,N_10746);
or U11327 (N_11327,N_10917,N_10748);
xor U11328 (N_11328,N_10889,N_10579);
and U11329 (N_11329,N_10906,N_10571);
xor U11330 (N_11330,N_10658,N_10565);
nand U11331 (N_11331,N_10753,N_10857);
nor U11332 (N_11332,N_10697,N_10773);
nand U11333 (N_11333,N_10880,N_10601);
nand U11334 (N_11334,N_10925,N_10798);
nand U11335 (N_11335,N_10796,N_10535);
xor U11336 (N_11336,N_10666,N_10505);
nor U11337 (N_11337,N_10947,N_10584);
nand U11338 (N_11338,N_10550,N_10693);
nor U11339 (N_11339,N_10513,N_10699);
and U11340 (N_11340,N_10586,N_10621);
xnor U11341 (N_11341,N_10578,N_10972);
nor U11342 (N_11342,N_10893,N_10615);
and U11343 (N_11343,N_10614,N_10609);
nand U11344 (N_11344,N_10951,N_10713);
nand U11345 (N_11345,N_10898,N_10671);
xor U11346 (N_11346,N_10824,N_10904);
xnor U11347 (N_11347,N_10783,N_10905);
xor U11348 (N_11348,N_10761,N_10887);
xnor U11349 (N_11349,N_10815,N_10997);
nand U11350 (N_11350,N_10889,N_10904);
xnor U11351 (N_11351,N_10814,N_10568);
nor U11352 (N_11352,N_10658,N_10680);
and U11353 (N_11353,N_10605,N_10558);
nor U11354 (N_11354,N_10953,N_10561);
or U11355 (N_11355,N_10792,N_10953);
xor U11356 (N_11356,N_10765,N_10925);
and U11357 (N_11357,N_10531,N_10750);
nor U11358 (N_11358,N_10955,N_10835);
xnor U11359 (N_11359,N_10823,N_10844);
and U11360 (N_11360,N_10926,N_10798);
and U11361 (N_11361,N_10657,N_10743);
or U11362 (N_11362,N_10585,N_10911);
nand U11363 (N_11363,N_10610,N_10557);
nand U11364 (N_11364,N_10945,N_10655);
xor U11365 (N_11365,N_10783,N_10990);
or U11366 (N_11366,N_10708,N_10797);
nand U11367 (N_11367,N_10717,N_10584);
nor U11368 (N_11368,N_10680,N_10760);
nand U11369 (N_11369,N_10911,N_10952);
or U11370 (N_11370,N_10720,N_10577);
nand U11371 (N_11371,N_10655,N_10949);
and U11372 (N_11372,N_10829,N_10689);
or U11373 (N_11373,N_10762,N_10502);
or U11374 (N_11374,N_10851,N_10773);
and U11375 (N_11375,N_10633,N_10991);
xor U11376 (N_11376,N_10884,N_10787);
nor U11377 (N_11377,N_10932,N_10809);
nor U11378 (N_11378,N_10770,N_10814);
nor U11379 (N_11379,N_10759,N_10626);
or U11380 (N_11380,N_10595,N_10901);
or U11381 (N_11381,N_10992,N_10578);
nor U11382 (N_11382,N_10520,N_10892);
and U11383 (N_11383,N_10961,N_10522);
and U11384 (N_11384,N_10955,N_10976);
nor U11385 (N_11385,N_10638,N_10797);
nand U11386 (N_11386,N_10943,N_10616);
xor U11387 (N_11387,N_10868,N_10900);
and U11388 (N_11388,N_10922,N_10907);
and U11389 (N_11389,N_10964,N_10712);
or U11390 (N_11390,N_10834,N_10812);
nor U11391 (N_11391,N_10851,N_10513);
or U11392 (N_11392,N_10526,N_10848);
and U11393 (N_11393,N_10684,N_10819);
or U11394 (N_11394,N_10515,N_10915);
xnor U11395 (N_11395,N_10752,N_10616);
nor U11396 (N_11396,N_10899,N_10575);
nand U11397 (N_11397,N_10955,N_10880);
nor U11398 (N_11398,N_10833,N_10980);
xnor U11399 (N_11399,N_10775,N_10541);
nor U11400 (N_11400,N_10638,N_10694);
nand U11401 (N_11401,N_10890,N_10793);
nand U11402 (N_11402,N_10626,N_10914);
or U11403 (N_11403,N_10786,N_10517);
nor U11404 (N_11404,N_10904,N_10705);
and U11405 (N_11405,N_10853,N_10812);
nor U11406 (N_11406,N_10692,N_10711);
nand U11407 (N_11407,N_10521,N_10657);
nor U11408 (N_11408,N_10708,N_10752);
xnor U11409 (N_11409,N_10679,N_10772);
xor U11410 (N_11410,N_10908,N_10919);
nor U11411 (N_11411,N_10998,N_10728);
and U11412 (N_11412,N_10505,N_10522);
or U11413 (N_11413,N_10573,N_10921);
nor U11414 (N_11414,N_10801,N_10569);
and U11415 (N_11415,N_10996,N_10760);
xnor U11416 (N_11416,N_10853,N_10884);
nand U11417 (N_11417,N_10537,N_10550);
xor U11418 (N_11418,N_10883,N_10975);
nor U11419 (N_11419,N_10966,N_10671);
nand U11420 (N_11420,N_10983,N_10903);
nor U11421 (N_11421,N_10645,N_10850);
nor U11422 (N_11422,N_10891,N_10744);
nand U11423 (N_11423,N_10852,N_10596);
nor U11424 (N_11424,N_10800,N_10940);
or U11425 (N_11425,N_10918,N_10710);
nor U11426 (N_11426,N_10569,N_10637);
and U11427 (N_11427,N_10878,N_10779);
nor U11428 (N_11428,N_10984,N_10747);
or U11429 (N_11429,N_10640,N_10531);
and U11430 (N_11430,N_10787,N_10928);
nor U11431 (N_11431,N_10814,N_10832);
or U11432 (N_11432,N_10646,N_10512);
and U11433 (N_11433,N_10573,N_10747);
or U11434 (N_11434,N_10683,N_10523);
and U11435 (N_11435,N_10971,N_10938);
and U11436 (N_11436,N_10849,N_10912);
and U11437 (N_11437,N_10739,N_10991);
or U11438 (N_11438,N_10936,N_10761);
or U11439 (N_11439,N_10627,N_10678);
nor U11440 (N_11440,N_10502,N_10601);
xnor U11441 (N_11441,N_10888,N_10829);
xnor U11442 (N_11442,N_10912,N_10580);
nand U11443 (N_11443,N_10862,N_10863);
or U11444 (N_11444,N_10966,N_10679);
and U11445 (N_11445,N_10534,N_10738);
xor U11446 (N_11446,N_10628,N_10572);
xor U11447 (N_11447,N_10590,N_10813);
and U11448 (N_11448,N_10872,N_10849);
or U11449 (N_11449,N_10903,N_10766);
or U11450 (N_11450,N_10651,N_10599);
nand U11451 (N_11451,N_10519,N_10662);
and U11452 (N_11452,N_10578,N_10698);
xnor U11453 (N_11453,N_10816,N_10564);
xor U11454 (N_11454,N_10666,N_10907);
nor U11455 (N_11455,N_10547,N_10768);
nand U11456 (N_11456,N_10636,N_10868);
nor U11457 (N_11457,N_10914,N_10694);
or U11458 (N_11458,N_10505,N_10754);
nor U11459 (N_11459,N_10835,N_10967);
nor U11460 (N_11460,N_10991,N_10839);
nand U11461 (N_11461,N_10534,N_10553);
nor U11462 (N_11462,N_10882,N_10909);
and U11463 (N_11463,N_10992,N_10655);
xor U11464 (N_11464,N_10624,N_10895);
and U11465 (N_11465,N_10690,N_10812);
xnor U11466 (N_11466,N_10677,N_10564);
nand U11467 (N_11467,N_10993,N_10777);
nand U11468 (N_11468,N_10868,N_10596);
nand U11469 (N_11469,N_10982,N_10578);
nand U11470 (N_11470,N_10630,N_10903);
nor U11471 (N_11471,N_10920,N_10804);
and U11472 (N_11472,N_10790,N_10856);
or U11473 (N_11473,N_10551,N_10546);
nor U11474 (N_11474,N_10629,N_10814);
nand U11475 (N_11475,N_10758,N_10597);
and U11476 (N_11476,N_10980,N_10664);
xnor U11477 (N_11477,N_10595,N_10621);
and U11478 (N_11478,N_10816,N_10587);
nor U11479 (N_11479,N_10844,N_10878);
and U11480 (N_11480,N_10899,N_10875);
and U11481 (N_11481,N_10756,N_10804);
or U11482 (N_11482,N_10962,N_10725);
nor U11483 (N_11483,N_10869,N_10759);
xnor U11484 (N_11484,N_10596,N_10863);
xor U11485 (N_11485,N_10589,N_10711);
and U11486 (N_11486,N_10505,N_10727);
or U11487 (N_11487,N_10992,N_10688);
nand U11488 (N_11488,N_10845,N_10939);
xnor U11489 (N_11489,N_10531,N_10952);
xor U11490 (N_11490,N_10793,N_10771);
or U11491 (N_11491,N_10545,N_10708);
nor U11492 (N_11492,N_10599,N_10761);
nand U11493 (N_11493,N_10525,N_10550);
xnor U11494 (N_11494,N_10753,N_10829);
nand U11495 (N_11495,N_10664,N_10720);
nand U11496 (N_11496,N_10646,N_10608);
nand U11497 (N_11497,N_10804,N_10729);
or U11498 (N_11498,N_10525,N_10601);
nand U11499 (N_11499,N_10774,N_10576);
nand U11500 (N_11500,N_11314,N_11218);
xor U11501 (N_11501,N_11379,N_11120);
xor U11502 (N_11502,N_11066,N_11170);
xor U11503 (N_11503,N_11094,N_11315);
nand U11504 (N_11504,N_11406,N_11029);
xor U11505 (N_11505,N_11189,N_11125);
nand U11506 (N_11506,N_11443,N_11147);
and U11507 (N_11507,N_11131,N_11168);
and U11508 (N_11508,N_11145,N_11467);
nand U11509 (N_11509,N_11446,N_11305);
or U11510 (N_11510,N_11191,N_11181);
nand U11511 (N_11511,N_11038,N_11163);
nand U11512 (N_11512,N_11090,N_11475);
nand U11513 (N_11513,N_11386,N_11450);
nand U11514 (N_11514,N_11052,N_11018);
nor U11515 (N_11515,N_11167,N_11397);
xnor U11516 (N_11516,N_11266,N_11077);
xnor U11517 (N_11517,N_11150,N_11425);
or U11518 (N_11518,N_11025,N_11304);
nand U11519 (N_11519,N_11206,N_11358);
nor U11520 (N_11520,N_11354,N_11098);
or U11521 (N_11521,N_11008,N_11026);
nand U11522 (N_11522,N_11208,N_11123);
and U11523 (N_11523,N_11159,N_11117);
or U11524 (N_11524,N_11148,N_11111);
or U11525 (N_11525,N_11118,N_11031);
xnor U11526 (N_11526,N_11114,N_11325);
nor U11527 (N_11527,N_11065,N_11192);
and U11528 (N_11528,N_11233,N_11087);
nand U11529 (N_11529,N_11193,N_11011);
and U11530 (N_11530,N_11432,N_11010);
nor U11531 (N_11531,N_11422,N_11494);
nor U11532 (N_11532,N_11166,N_11198);
xor U11533 (N_11533,N_11368,N_11486);
nor U11534 (N_11534,N_11057,N_11230);
and U11535 (N_11535,N_11106,N_11030);
or U11536 (N_11536,N_11171,N_11319);
nand U11537 (N_11537,N_11188,N_11149);
or U11538 (N_11538,N_11477,N_11037);
nand U11539 (N_11539,N_11427,N_11258);
nor U11540 (N_11540,N_11219,N_11023);
or U11541 (N_11541,N_11491,N_11240);
and U11542 (N_11542,N_11341,N_11134);
xnor U11543 (N_11543,N_11400,N_11330);
nand U11544 (N_11544,N_11212,N_11173);
nand U11545 (N_11545,N_11271,N_11039);
nand U11546 (N_11546,N_11311,N_11448);
xor U11547 (N_11547,N_11115,N_11210);
and U11548 (N_11548,N_11403,N_11441);
and U11549 (N_11549,N_11299,N_11091);
nor U11550 (N_11550,N_11069,N_11370);
or U11551 (N_11551,N_11267,N_11468);
and U11552 (N_11552,N_11202,N_11339);
nand U11553 (N_11553,N_11490,N_11155);
nand U11554 (N_11554,N_11074,N_11351);
nand U11555 (N_11555,N_11433,N_11156);
or U11556 (N_11556,N_11084,N_11485);
and U11557 (N_11557,N_11287,N_11479);
nor U11558 (N_11558,N_11059,N_11333);
and U11559 (N_11559,N_11332,N_11153);
and U11560 (N_11560,N_11020,N_11234);
nor U11561 (N_11561,N_11036,N_11488);
nand U11562 (N_11562,N_11042,N_11334);
xnor U11563 (N_11563,N_11337,N_11264);
xnor U11564 (N_11564,N_11353,N_11110);
nand U11565 (N_11565,N_11027,N_11205);
and U11566 (N_11566,N_11024,N_11127);
or U11567 (N_11567,N_11412,N_11157);
xor U11568 (N_11568,N_11273,N_11423);
xnor U11569 (N_11569,N_11165,N_11478);
xnor U11570 (N_11570,N_11275,N_11414);
xnor U11571 (N_11571,N_11146,N_11225);
nor U11572 (N_11572,N_11221,N_11396);
nand U11573 (N_11573,N_11277,N_11142);
nand U11574 (N_11574,N_11032,N_11420);
nor U11575 (N_11575,N_11338,N_11112);
nor U11576 (N_11576,N_11001,N_11250);
nand U11577 (N_11577,N_11308,N_11133);
xor U11578 (N_11578,N_11194,N_11092);
nand U11579 (N_11579,N_11228,N_11238);
or U11580 (N_11580,N_11377,N_11384);
and U11581 (N_11581,N_11435,N_11487);
or U11582 (N_11582,N_11140,N_11455);
and U11583 (N_11583,N_11005,N_11324);
nand U11584 (N_11584,N_11312,N_11051);
xor U11585 (N_11585,N_11348,N_11257);
nor U11586 (N_11586,N_11043,N_11089);
and U11587 (N_11587,N_11070,N_11461);
or U11588 (N_11588,N_11410,N_11232);
nor U11589 (N_11589,N_11045,N_11101);
and U11590 (N_11590,N_11430,N_11012);
xor U11591 (N_11591,N_11434,N_11498);
or U11592 (N_11592,N_11102,N_11096);
nand U11593 (N_11593,N_11457,N_11454);
nor U11594 (N_11594,N_11175,N_11122);
or U11595 (N_11595,N_11076,N_11345);
and U11596 (N_11596,N_11442,N_11280);
nor U11597 (N_11597,N_11174,N_11383);
or U11598 (N_11598,N_11121,N_11183);
nor U11599 (N_11599,N_11137,N_11364);
or U11600 (N_11600,N_11391,N_11374);
nand U11601 (N_11601,N_11048,N_11180);
and U11602 (N_11602,N_11399,N_11429);
nor U11603 (N_11603,N_11046,N_11285);
and U11604 (N_11604,N_11007,N_11003);
or U11605 (N_11605,N_11313,N_11317);
xnor U11606 (N_11606,N_11154,N_11099);
xnor U11607 (N_11607,N_11318,N_11215);
or U11608 (N_11608,N_11229,N_11058);
xor U11609 (N_11609,N_11022,N_11371);
xor U11610 (N_11610,N_11105,N_11224);
or U11611 (N_11611,N_11081,N_11458);
nand U11612 (N_11612,N_11116,N_11331);
and U11613 (N_11613,N_11108,N_11342);
xor U11614 (N_11614,N_11244,N_11359);
or U11615 (N_11615,N_11404,N_11248);
and U11616 (N_11616,N_11416,N_11109);
nand U11617 (N_11617,N_11204,N_11056);
nand U11618 (N_11618,N_11428,N_11437);
nand U11619 (N_11619,N_11344,N_11247);
xor U11620 (N_11620,N_11255,N_11365);
or U11621 (N_11621,N_11360,N_11392);
xor U11622 (N_11622,N_11409,N_11380);
or U11623 (N_11623,N_11436,N_11418);
or U11624 (N_11624,N_11469,N_11214);
xor U11625 (N_11625,N_11246,N_11292);
nand U11626 (N_11626,N_11297,N_11073);
nand U11627 (N_11627,N_11213,N_11449);
or U11628 (N_11628,N_11444,N_11465);
or U11629 (N_11629,N_11295,N_11274);
and U11630 (N_11630,N_11321,N_11323);
and U11631 (N_11631,N_11265,N_11211);
or U11632 (N_11632,N_11000,N_11252);
and U11633 (N_11633,N_11417,N_11268);
xor U11634 (N_11634,N_11367,N_11472);
nand U11635 (N_11635,N_11340,N_11372);
or U11636 (N_11636,N_11398,N_11347);
or U11637 (N_11637,N_11289,N_11326);
or U11638 (N_11638,N_11049,N_11316);
or U11639 (N_11639,N_11482,N_11216);
xor U11640 (N_11640,N_11373,N_11253);
nand U11641 (N_11641,N_11261,N_11044);
or U11642 (N_11642,N_11064,N_11055);
xor U11643 (N_11643,N_11471,N_11207);
nor U11644 (N_11644,N_11484,N_11186);
xnor U11645 (N_11645,N_11050,N_11242);
nor U11646 (N_11646,N_11381,N_11415);
xor U11647 (N_11647,N_11178,N_11119);
or U11648 (N_11648,N_11141,N_11306);
xnor U11649 (N_11649,N_11093,N_11493);
nor U11650 (N_11650,N_11424,N_11002);
xnor U11651 (N_11651,N_11236,N_11209);
nand U11652 (N_11652,N_11300,N_11309);
nand U11653 (N_11653,N_11172,N_11335);
or U11654 (N_11654,N_11041,N_11237);
nor U11655 (N_11655,N_11245,N_11426);
and U11656 (N_11656,N_11097,N_11389);
nand U11657 (N_11657,N_11307,N_11222);
nand U11658 (N_11658,N_11382,N_11362);
nor U11659 (N_11659,N_11480,N_11203);
xor U11660 (N_11660,N_11408,N_11256);
nand U11661 (N_11661,N_11489,N_11294);
and U11662 (N_11662,N_11466,N_11013);
nor U11663 (N_11663,N_11162,N_11366);
and U11664 (N_11664,N_11462,N_11394);
xnor U11665 (N_11665,N_11495,N_11067);
and U11666 (N_11666,N_11390,N_11113);
xor U11667 (N_11667,N_11459,N_11496);
nand U11668 (N_11668,N_11452,N_11009);
and U11669 (N_11669,N_11251,N_11291);
xnor U11670 (N_11670,N_11034,N_11243);
nand U11671 (N_11671,N_11078,N_11260);
and U11672 (N_11672,N_11082,N_11464);
nor U11673 (N_11673,N_11278,N_11016);
xnor U11674 (N_11674,N_11103,N_11343);
nor U11675 (N_11675,N_11035,N_11350);
or U11676 (N_11676,N_11336,N_11470);
xor U11677 (N_11677,N_11355,N_11231);
or U11678 (N_11678,N_11176,N_11499);
xnor U11679 (N_11679,N_11376,N_11182);
and U11680 (N_11680,N_11259,N_11328);
nand U11681 (N_11681,N_11402,N_11438);
and U11682 (N_11682,N_11405,N_11160);
xnor U11683 (N_11683,N_11262,N_11021);
nand U11684 (N_11684,N_11144,N_11130);
nand U11685 (N_11685,N_11138,N_11196);
and U11686 (N_11686,N_11015,N_11227);
nand U11687 (N_11687,N_11124,N_11393);
nor U11688 (N_11688,N_11068,N_11378);
xnor U11689 (N_11689,N_11346,N_11047);
xnor U11690 (N_11690,N_11290,N_11263);
nand U11691 (N_11691,N_11169,N_11282);
or U11692 (N_11692,N_11132,N_11473);
nand U11693 (N_11693,N_11476,N_11184);
nand U11694 (N_11694,N_11497,N_11288);
nor U11695 (N_11695,N_11445,N_11440);
xor U11696 (N_11696,N_11320,N_11302);
nand U11697 (N_11697,N_11135,N_11270);
nand U11698 (N_11698,N_11357,N_11195);
or U11699 (N_11699,N_11028,N_11387);
or U11700 (N_11700,N_11327,N_11136);
or U11701 (N_11701,N_11283,N_11293);
nand U11702 (N_11702,N_11152,N_11126);
or U11703 (N_11703,N_11086,N_11421);
nor U11704 (N_11704,N_11481,N_11411);
nor U11705 (N_11705,N_11158,N_11419);
or U11706 (N_11706,N_11492,N_11201);
xnor U11707 (N_11707,N_11128,N_11298);
xor U11708 (N_11708,N_11447,N_11281);
xor U11709 (N_11709,N_11104,N_11017);
or U11710 (N_11710,N_11272,N_11033);
xnor U11711 (N_11711,N_11303,N_11407);
and U11712 (N_11712,N_11356,N_11269);
nor U11713 (N_11713,N_11296,N_11040);
nand U11714 (N_11714,N_11284,N_11185);
or U11715 (N_11715,N_11019,N_11004);
xnor U11716 (N_11716,N_11187,N_11385);
xnor U11717 (N_11717,N_11431,N_11451);
or U11718 (N_11718,N_11235,N_11054);
or U11719 (N_11719,N_11075,N_11088);
or U11720 (N_11720,N_11463,N_11279);
xnor U11721 (N_11721,N_11197,N_11301);
and U11722 (N_11722,N_11080,N_11329);
nand U11723 (N_11723,N_11363,N_11352);
or U11724 (N_11724,N_11375,N_11177);
nand U11725 (N_11725,N_11095,N_11060);
or U11726 (N_11726,N_11062,N_11226);
xnor U11727 (N_11727,N_11063,N_11053);
nand U11728 (N_11728,N_11061,N_11161);
and U11729 (N_11729,N_11079,N_11223);
and U11730 (N_11730,N_11100,N_11164);
nand U11731 (N_11731,N_11129,N_11286);
or U11732 (N_11732,N_11456,N_11369);
or U11733 (N_11733,N_11254,N_11453);
xnor U11734 (N_11734,N_11249,N_11190);
or U11735 (N_11735,N_11474,N_11239);
nor U11736 (N_11736,N_11083,N_11014);
nand U11737 (N_11737,N_11200,N_11199);
nand U11738 (N_11738,N_11220,N_11439);
or U11739 (N_11739,N_11388,N_11151);
nand U11740 (N_11740,N_11072,N_11085);
and U11741 (N_11741,N_11401,N_11361);
or U11742 (N_11742,N_11143,N_11322);
or U11743 (N_11743,N_11241,N_11310);
and U11744 (N_11744,N_11483,N_11460);
or U11745 (N_11745,N_11071,N_11349);
nor U11746 (N_11746,N_11006,N_11179);
and U11747 (N_11747,N_11276,N_11413);
and U11748 (N_11748,N_11139,N_11217);
or U11749 (N_11749,N_11395,N_11107);
or U11750 (N_11750,N_11184,N_11444);
xor U11751 (N_11751,N_11395,N_11479);
xor U11752 (N_11752,N_11331,N_11254);
xnor U11753 (N_11753,N_11396,N_11044);
or U11754 (N_11754,N_11447,N_11269);
nand U11755 (N_11755,N_11349,N_11130);
nor U11756 (N_11756,N_11353,N_11257);
or U11757 (N_11757,N_11153,N_11453);
nand U11758 (N_11758,N_11399,N_11306);
nand U11759 (N_11759,N_11182,N_11256);
or U11760 (N_11760,N_11480,N_11238);
xnor U11761 (N_11761,N_11387,N_11094);
xor U11762 (N_11762,N_11328,N_11104);
nor U11763 (N_11763,N_11055,N_11143);
nand U11764 (N_11764,N_11386,N_11358);
and U11765 (N_11765,N_11406,N_11181);
or U11766 (N_11766,N_11330,N_11269);
or U11767 (N_11767,N_11294,N_11179);
and U11768 (N_11768,N_11251,N_11444);
or U11769 (N_11769,N_11258,N_11422);
nor U11770 (N_11770,N_11140,N_11075);
and U11771 (N_11771,N_11459,N_11325);
or U11772 (N_11772,N_11071,N_11328);
and U11773 (N_11773,N_11387,N_11473);
nand U11774 (N_11774,N_11163,N_11040);
nor U11775 (N_11775,N_11223,N_11007);
or U11776 (N_11776,N_11103,N_11067);
and U11777 (N_11777,N_11467,N_11414);
nand U11778 (N_11778,N_11097,N_11066);
and U11779 (N_11779,N_11469,N_11220);
or U11780 (N_11780,N_11425,N_11326);
and U11781 (N_11781,N_11326,N_11342);
or U11782 (N_11782,N_11286,N_11375);
xnor U11783 (N_11783,N_11113,N_11369);
nor U11784 (N_11784,N_11006,N_11141);
nand U11785 (N_11785,N_11373,N_11181);
nand U11786 (N_11786,N_11356,N_11146);
nand U11787 (N_11787,N_11404,N_11253);
or U11788 (N_11788,N_11377,N_11338);
nor U11789 (N_11789,N_11059,N_11117);
or U11790 (N_11790,N_11212,N_11416);
xor U11791 (N_11791,N_11113,N_11349);
nand U11792 (N_11792,N_11269,N_11215);
nor U11793 (N_11793,N_11435,N_11472);
or U11794 (N_11794,N_11304,N_11225);
nand U11795 (N_11795,N_11397,N_11321);
or U11796 (N_11796,N_11208,N_11404);
nor U11797 (N_11797,N_11023,N_11144);
xor U11798 (N_11798,N_11141,N_11296);
nand U11799 (N_11799,N_11486,N_11333);
nor U11800 (N_11800,N_11034,N_11004);
nand U11801 (N_11801,N_11170,N_11394);
xnor U11802 (N_11802,N_11305,N_11302);
and U11803 (N_11803,N_11153,N_11204);
or U11804 (N_11804,N_11329,N_11066);
nand U11805 (N_11805,N_11239,N_11487);
or U11806 (N_11806,N_11176,N_11293);
nor U11807 (N_11807,N_11314,N_11169);
or U11808 (N_11808,N_11006,N_11090);
or U11809 (N_11809,N_11250,N_11018);
or U11810 (N_11810,N_11145,N_11322);
and U11811 (N_11811,N_11181,N_11157);
or U11812 (N_11812,N_11007,N_11313);
xor U11813 (N_11813,N_11013,N_11463);
nand U11814 (N_11814,N_11236,N_11482);
xor U11815 (N_11815,N_11048,N_11086);
xnor U11816 (N_11816,N_11004,N_11279);
xnor U11817 (N_11817,N_11465,N_11473);
xnor U11818 (N_11818,N_11238,N_11155);
nand U11819 (N_11819,N_11447,N_11338);
nor U11820 (N_11820,N_11440,N_11423);
or U11821 (N_11821,N_11260,N_11462);
nor U11822 (N_11822,N_11202,N_11376);
nor U11823 (N_11823,N_11234,N_11041);
xor U11824 (N_11824,N_11403,N_11453);
and U11825 (N_11825,N_11067,N_11265);
and U11826 (N_11826,N_11228,N_11397);
xnor U11827 (N_11827,N_11468,N_11125);
xnor U11828 (N_11828,N_11198,N_11205);
or U11829 (N_11829,N_11448,N_11050);
nand U11830 (N_11830,N_11038,N_11439);
and U11831 (N_11831,N_11494,N_11049);
and U11832 (N_11832,N_11288,N_11281);
and U11833 (N_11833,N_11083,N_11103);
nand U11834 (N_11834,N_11308,N_11166);
or U11835 (N_11835,N_11102,N_11118);
or U11836 (N_11836,N_11317,N_11420);
and U11837 (N_11837,N_11334,N_11366);
nor U11838 (N_11838,N_11317,N_11476);
nor U11839 (N_11839,N_11489,N_11099);
or U11840 (N_11840,N_11043,N_11261);
xor U11841 (N_11841,N_11321,N_11496);
nor U11842 (N_11842,N_11168,N_11040);
nand U11843 (N_11843,N_11318,N_11092);
and U11844 (N_11844,N_11045,N_11108);
or U11845 (N_11845,N_11309,N_11431);
and U11846 (N_11846,N_11490,N_11081);
or U11847 (N_11847,N_11317,N_11188);
xor U11848 (N_11848,N_11242,N_11370);
nor U11849 (N_11849,N_11017,N_11286);
and U11850 (N_11850,N_11091,N_11167);
nor U11851 (N_11851,N_11459,N_11389);
xnor U11852 (N_11852,N_11333,N_11018);
or U11853 (N_11853,N_11437,N_11186);
and U11854 (N_11854,N_11209,N_11219);
xor U11855 (N_11855,N_11226,N_11213);
and U11856 (N_11856,N_11355,N_11202);
or U11857 (N_11857,N_11100,N_11427);
nand U11858 (N_11858,N_11013,N_11462);
nand U11859 (N_11859,N_11419,N_11136);
xnor U11860 (N_11860,N_11341,N_11142);
and U11861 (N_11861,N_11143,N_11231);
xnor U11862 (N_11862,N_11445,N_11303);
nor U11863 (N_11863,N_11388,N_11027);
nor U11864 (N_11864,N_11018,N_11485);
or U11865 (N_11865,N_11117,N_11440);
nor U11866 (N_11866,N_11305,N_11397);
or U11867 (N_11867,N_11398,N_11037);
and U11868 (N_11868,N_11221,N_11313);
and U11869 (N_11869,N_11158,N_11159);
and U11870 (N_11870,N_11453,N_11031);
and U11871 (N_11871,N_11229,N_11419);
xor U11872 (N_11872,N_11312,N_11443);
xor U11873 (N_11873,N_11029,N_11174);
nor U11874 (N_11874,N_11267,N_11394);
nand U11875 (N_11875,N_11322,N_11151);
nor U11876 (N_11876,N_11427,N_11321);
and U11877 (N_11877,N_11412,N_11078);
or U11878 (N_11878,N_11285,N_11414);
xor U11879 (N_11879,N_11367,N_11069);
nand U11880 (N_11880,N_11412,N_11338);
nor U11881 (N_11881,N_11325,N_11066);
nand U11882 (N_11882,N_11272,N_11139);
nor U11883 (N_11883,N_11321,N_11141);
xnor U11884 (N_11884,N_11201,N_11224);
or U11885 (N_11885,N_11283,N_11188);
xor U11886 (N_11886,N_11176,N_11110);
and U11887 (N_11887,N_11294,N_11094);
xnor U11888 (N_11888,N_11201,N_11264);
nand U11889 (N_11889,N_11048,N_11096);
or U11890 (N_11890,N_11272,N_11167);
or U11891 (N_11891,N_11483,N_11058);
nand U11892 (N_11892,N_11378,N_11380);
nand U11893 (N_11893,N_11287,N_11231);
or U11894 (N_11894,N_11230,N_11320);
and U11895 (N_11895,N_11318,N_11168);
xor U11896 (N_11896,N_11339,N_11348);
nand U11897 (N_11897,N_11279,N_11477);
or U11898 (N_11898,N_11300,N_11215);
xnor U11899 (N_11899,N_11418,N_11049);
nand U11900 (N_11900,N_11431,N_11404);
nand U11901 (N_11901,N_11439,N_11159);
xor U11902 (N_11902,N_11388,N_11229);
and U11903 (N_11903,N_11042,N_11414);
xnor U11904 (N_11904,N_11199,N_11031);
or U11905 (N_11905,N_11388,N_11186);
xnor U11906 (N_11906,N_11274,N_11009);
xnor U11907 (N_11907,N_11487,N_11381);
or U11908 (N_11908,N_11479,N_11396);
nor U11909 (N_11909,N_11256,N_11134);
xnor U11910 (N_11910,N_11039,N_11336);
nand U11911 (N_11911,N_11202,N_11485);
nand U11912 (N_11912,N_11111,N_11185);
xnor U11913 (N_11913,N_11240,N_11123);
or U11914 (N_11914,N_11227,N_11072);
nor U11915 (N_11915,N_11073,N_11392);
or U11916 (N_11916,N_11023,N_11283);
and U11917 (N_11917,N_11318,N_11359);
nor U11918 (N_11918,N_11167,N_11140);
xnor U11919 (N_11919,N_11443,N_11383);
nor U11920 (N_11920,N_11450,N_11155);
and U11921 (N_11921,N_11032,N_11311);
xor U11922 (N_11922,N_11025,N_11104);
nand U11923 (N_11923,N_11247,N_11094);
or U11924 (N_11924,N_11012,N_11486);
nor U11925 (N_11925,N_11388,N_11440);
and U11926 (N_11926,N_11391,N_11103);
xor U11927 (N_11927,N_11464,N_11056);
or U11928 (N_11928,N_11487,N_11392);
and U11929 (N_11929,N_11497,N_11498);
nor U11930 (N_11930,N_11254,N_11440);
xor U11931 (N_11931,N_11313,N_11443);
nor U11932 (N_11932,N_11421,N_11293);
or U11933 (N_11933,N_11166,N_11415);
nand U11934 (N_11934,N_11112,N_11364);
and U11935 (N_11935,N_11065,N_11275);
xor U11936 (N_11936,N_11121,N_11368);
xor U11937 (N_11937,N_11036,N_11205);
or U11938 (N_11938,N_11120,N_11206);
or U11939 (N_11939,N_11119,N_11346);
nor U11940 (N_11940,N_11323,N_11374);
nand U11941 (N_11941,N_11079,N_11029);
nor U11942 (N_11942,N_11068,N_11437);
nor U11943 (N_11943,N_11197,N_11317);
and U11944 (N_11944,N_11201,N_11165);
nor U11945 (N_11945,N_11413,N_11263);
nor U11946 (N_11946,N_11037,N_11281);
or U11947 (N_11947,N_11474,N_11078);
nand U11948 (N_11948,N_11297,N_11125);
nand U11949 (N_11949,N_11422,N_11483);
or U11950 (N_11950,N_11461,N_11126);
xor U11951 (N_11951,N_11188,N_11193);
xnor U11952 (N_11952,N_11375,N_11018);
nor U11953 (N_11953,N_11116,N_11234);
and U11954 (N_11954,N_11309,N_11070);
nand U11955 (N_11955,N_11065,N_11368);
and U11956 (N_11956,N_11158,N_11493);
nor U11957 (N_11957,N_11192,N_11027);
xnor U11958 (N_11958,N_11217,N_11105);
nor U11959 (N_11959,N_11372,N_11001);
and U11960 (N_11960,N_11134,N_11171);
xor U11961 (N_11961,N_11163,N_11274);
and U11962 (N_11962,N_11314,N_11258);
xor U11963 (N_11963,N_11423,N_11367);
nand U11964 (N_11964,N_11166,N_11201);
xnor U11965 (N_11965,N_11448,N_11003);
and U11966 (N_11966,N_11004,N_11431);
xnor U11967 (N_11967,N_11292,N_11085);
xor U11968 (N_11968,N_11236,N_11346);
nor U11969 (N_11969,N_11048,N_11274);
nor U11970 (N_11970,N_11459,N_11429);
nand U11971 (N_11971,N_11432,N_11129);
xnor U11972 (N_11972,N_11262,N_11181);
or U11973 (N_11973,N_11339,N_11183);
or U11974 (N_11974,N_11008,N_11425);
or U11975 (N_11975,N_11369,N_11226);
nand U11976 (N_11976,N_11190,N_11363);
nor U11977 (N_11977,N_11402,N_11129);
nand U11978 (N_11978,N_11180,N_11005);
nor U11979 (N_11979,N_11130,N_11170);
nand U11980 (N_11980,N_11178,N_11485);
xor U11981 (N_11981,N_11140,N_11396);
and U11982 (N_11982,N_11083,N_11299);
and U11983 (N_11983,N_11463,N_11362);
nor U11984 (N_11984,N_11385,N_11463);
and U11985 (N_11985,N_11333,N_11134);
nor U11986 (N_11986,N_11163,N_11045);
nand U11987 (N_11987,N_11324,N_11221);
xor U11988 (N_11988,N_11483,N_11362);
nor U11989 (N_11989,N_11013,N_11243);
and U11990 (N_11990,N_11443,N_11467);
and U11991 (N_11991,N_11266,N_11057);
nor U11992 (N_11992,N_11388,N_11334);
nand U11993 (N_11993,N_11375,N_11045);
nand U11994 (N_11994,N_11243,N_11075);
nand U11995 (N_11995,N_11303,N_11218);
xnor U11996 (N_11996,N_11363,N_11065);
and U11997 (N_11997,N_11488,N_11072);
or U11998 (N_11998,N_11048,N_11418);
xor U11999 (N_11999,N_11141,N_11232);
xor U12000 (N_12000,N_11564,N_11833);
nand U12001 (N_12001,N_11814,N_11985);
and U12002 (N_12002,N_11509,N_11531);
nand U12003 (N_12003,N_11544,N_11717);
or U12004 (N_12004,N_11958,N_11730);
xnor U12005 (N_12005,N_11984,N_11608);
nand U12006 (N_12006,N_11554,N_11806);
and U12007 (N_12007,N_11713,N_11714);
or U12008 (N_12008,N_11828,N_11522);
xor U12009 (N_12009,N_11679,N_11678);
nor U12010 (N_12010,N_11595,N_11987);
nand U12011 (N_12011,N_11941,N_11621);
nor U12012 (N_12012,N_11942,N_11964);
xor U12013 (N_12013,N_11562,N_11688);
nor U12014 (N_12014,N_11890,N_11517);
or U12015 (N_12015,N_11909,N_11514);
nor U12016 (N_12016,N_11691,N_11537);
nand U12017 (N_12017,N_11755,N_11983);
xnor U12018 (N_12018,N_11644,N_11732);
and U12019 (N_12019,N_11830,N_11752);
or U12020 (N_12020,N_11640,N_11816);
xor U12021 (N_12021,N_11797,N_11846);
nand U12022 (N_12022,N_11706,N_11799);
nor U12023 (N_12023,N_11515,N_11609);
or U12024 (N_12024,N_11548,N_11617);
and U12025 (N_12025,N_11520,N_11792);
nand U12026 (N_12026,N_11694,N_11980);
nor U12027 (N_12027,N_11920,N_11534);
or U12028 (N_12028,N_11676,N_11708);
nand U12029 (N_12029,N_11782,N_11989);
or U12030 (N_12030,N_11992,N_11769);
nand U12031 (N_12031,N_11986,N_11976);
nor U12032 (N_12032,N_11604,N_11669);
and U12033 (N_12033,N_11998,N_11837);
nor U12034 (N_12034,N_11930,N_11990);
nor U12035 (N_12035,N_11926,N_11660);
nand U12036 (N_12036,N_11583,N_11551);
or U12037 (N_12037,N_11800,N_11711);
nor U12038 (N_12038,N_11900,N_11695);
or U12039 (N_12039,N_11675,N_11826);
and U12040 (N_12040,N_11745,N_11581);
and U12041 (N_12041,N_11950,N_11911);
or U12042 (N_12042,N_11882,N_11994);
and U12043 (N_12043,N_11635,N_11997);
nor U12044 (N_12044,N_11703,N_11529);
xor U12045 (N_12045,N_11668,N_11663);
or U12046 (N_12046,N_11957,N_11982);
and U12047 (N_12047,N_11933,N_11588);
or U12048 (N_12048,N_11786,N_11892);
xnor U12049 (N_12049,N_11611,N_11569);
xnor U12050 (N_12050,N_11841,N_11666);
xnor U12051 (N_12051,N_11775,N_11712);
xor U12052 (N_12052,N_11507,N_11637);
and U12053 (N_12053,N_11704,N_11757);
xnor U12054 (N_12054,N_11856,N_11838);
or U12055 (N_12055,N_11571,N_11683);
nor U12056 (N_12056,N_11527,N_11824);
or U12057 (N_12057,N_11690,N_11705);
xnor U12058 (N_12058,N_11570,N_11511);
or U12059 (N_12059,N_11685,N_11863);
nand U12060 (N_12060,N_11988,N_11662);
xor U12061 (N_12061,N_11633,N_11532);
xor U12062 (N_12062,N_11650,N_11540);
nor U12063 (N_12063,N_11884,N_11839);
and U12064 (N_12064,N_11682,N_11654);
or U12065 (N_12065,N_11738,N_11724);
xor U12066 (N_12066,N_11916,N_11802);
and U12067 (N_12067,N_11613,N_11739);
xor U12068 (N_12068,N_11935,N_11743);
and U12069 (N_12069,N_11788,N_11567);
or U12070 (N_12070,N_11949,N_11969);
nand U12071 (N_12071,N_11879,N_11861);
and U12072 (N_12072,N_11908,N_11615);
nand U12073 (N_12073,N_11746,N_11995);
and U12074 (N_12074,N_11823,N_11598);
nand U12075 (N_12075,N_11597,N_11897);
or U12076 (N_12076,N_11963,N_11510);
or U12077 (N_12077,N_11525,N_11655);
or U12078 (N_12078,N_11643,N_11697);
nand U12079 (N_12079,N_11904,N_11818);
xor U12080 (N_12080,N_11565,N_11937);
or U12081 (N_12081,N_11710,N_11545);
or U12082 (N_12082,N_11812,N_11901);
xnor U12083 (N_12083,N_11751,N_11555);
nand U12084 (N_12084,N_11639,N_11991);
xnor U12085 (N_12085,N_11891,N_11858);
and U12086 (N_12086,N_11967,N_11898);
nand U12087 (N_12087,N_11822,N_11749);
or U12088 (N_12088,N_11726,N_11918);
or U12089 (N_12089,N_11894,N_11651);
nor U12090 (N_12090,N_11864,N_11912);
nor U12091 (N_12091,N_11731,N_11931);
or U12092 (N_12092,N_11886,N_11770);
nand U12093 (N_12093,N_11764,N_11878);
or U12094 (N_12094,N_11665,N_11850);
or U12095 (N_12095,N_11975,N_11533);
and U12096 (N_12096,N_11844,N_11560);
and U12097 (N_12097,N_11872,N_11512);
nor U12098 (N_12098,N_11725,N_11889);
or U12099 (N_12099,N_11981,N_11578);
xnor U12100 (N_12100,N_11780,N_11767);
nand U12101 (N_12101,N_11718,N_11526);
xnor U12102 (N_12102,N_11783,N_11915);
or U12103 (N_12103,N_11945,N_11661);
nor U12104 (N_12104,N_11993,N_11664);
nor U12105 (N_12105,N_11793,N_11747);
and U12106 (N_12106,N_11720,N_11550);
xor U12107 (N_12107,N_11952,N_11922);
or U12108 (N_12108,N_11847,N_11895);
nor U12109 (N_12109,N_11584,N_11760);
and U12110 (N_12110,N_11859,N_11519);
and U12111 (N_12111,N_11542,N_11681);
nor U12112 (N_12112,N_11524,N_11677);
or U12113 (N_12113,N_11590,N_11921);
xnor U12114 (N_12114,N_11836,N_11811);
xnor U12115 (N_12115,N_11742,N_11785);
xnor U12116 (N_12116,N_11728,N_11702);
or U12117 (N_12117,N_11721,N_11813);
nand U12118 (N_12118,N_11804,N_11899);
and U12119 (N_12119,N_11888,N_11781);
or U12120 (N_12120,N_11819,N_11636);
nor U12121 (N_12121,N_11734,N_11798);
and U12122 (N_12122,N_11599,N_11763);
or U12123 (N_12123,N_11853,N_11883);
nand U12124 (N_12124,N_11871,N_11947);
or U12125 (N_12125,N_11521,N_11500);
and U12126 (N_12126,N_11698,N_11996);
and U12127 (N_12127,N_11809,N_11924);
xor U12128 (N_12128,N_11848,N_11791);
nor U12129 (N_12129,N_11910,N_11808);
nor U12130 (N_12130,N_11552,N_11727);
and U12131 (N_12131,N_11541,N_11765);
xor U12132 (N_12132,N_11978,N_11652);
and U12133 (N_12133,N_11946,N_11936);
nand U12134 (N_12134,N_11502,N_11622);
nor U12135 (N_12135,N_11955,N_11960);
and U12136 (N_12136,N_11553,N_11586);
and U12137 (N_12137,N_11753,N_11944);
and U12138 (N_12138,N_11907,N_11956);
and U12139 (N_12139,N_11642,N_11674);
xor U12140 (N_12140,N_11647,N_11954);
and U12141 (N_12141,N_11672,N_11624);
nor U12142 (N_12142,N_11735,N_11687);
and U12143 (N_12143,N_11815,N_11953);
nand U12144 (N_12144,N_11641,N_11601);
or U12145 (N_12145,N_11585,N_11592);
xnor U12146 (N_12146,N_11972,N_11501);
or U12147 (N_12147,N_11868,N_11591);
nand U12148 (N_12148,N_11670,N_11699);
nand U12149 (N_12149,N_11539,N_11795);
and U12150 (N_12150,N_11754,N_11866);
and U12151 (N_12151,N_11787,N_11961);
and U12152 (N_12152,N_11602,N_11630);
nor U12153 (N_12153,N_11593,N_11938);
nand U12154 (N_12154,N_11543,N_11605);
or U12155 (N_12155,N_11736,N_11629);
and U12156 (N_12156,N_11845,N_11733);
nor U12157 (N_12157,N_11614,N_11729);
and U12158 (N_12158,N_11925,N_11707);
xnor U12159 (N_12159,N_11612,N_11790);
xnor U12160 (N_12160,N_11805,N_11865);
nor U12161 (N_12161,N_11905,N_11616);
xor U12162 (N_12162,N_11772,N_11744);
xnor U12163 (N_12163,N_11880,N_11842);
nand U12164 (N_12164,N_11796,N_11831);
nand U12165 (N_12165,N_11563,N_11914);
nor U12166 (N_12166,N_11821,N_11820);
or U12167 (N_12167,N_11577,N_11934);
and U12168 (N_12168,N_11758,N_11870);
xor U12169 (N_12169,N_11558,N_11832);
nand U12170 (N_12170,N_11874,N_11549);
or U12171 (N_12171,N_11970,N_11840);
or U12172 (N_12172,N_11885,N_11784);
or U12173 (N_12173,N_11761,N_11627);
xnor U12174 (N_12174,N_11535,N_11959);
xnor U12175 (N_12175,N_11771,N_11632);
or U12176 (N_12176,N_11580,N_11759);
nand U12177 (N_12177,N_11506,N_11919);
nand U12178 (N_12178,N_11851,N_11881);
nand U12179 (N_12179,N_11692,N_11530);
xnor U12180 (N_12180,N_11862,N_11538);
nor U12181 (N_12181,N_11631,N_11715);
xor U12182 (N_12182,N_11741,N_11620);
nor U12183 (N_12183,N_11834,N_11508);
and U12184 (N_12184,N_11547,N_11857);
xnor U12185 (N_12185,N_11927,N_11740);
xnor U12186 (N_12186,N_11594,N_11876);
nor U12187 (N_12187,N_11607,N_11877);
and U12188 (N_12188,N_11929,N_11855);
nand U12189 (N_12189,N_11778,N_11557);
nand U12190 (N_12190,N_11849,N_11977);
and U12191 (N_12191,N_11973,N_11928);
nor U12192 (N_12192,N_11825,N_11686);
nor U12193 (N_12193,N_11860,N_11566);
and U12194 (N_12194,N_11689,N_11902);
xnor U12195 (N_12195,N_11653,N_11579);
and U12196 (N_12196,N_11638,N_11582);
or U12197 (N_12197,N_11867,N_11893);
or U12198 (N_12198,N_11829,N_11854);
xnor U12199 (N_12199,N_11999,N_11574);
or U12200 (N_12200,N_11673,N_11974);
nand U12201 (N_12201,N_11794,N_11737);
and U12202 (N_12202,N_11873,N_11762);
or U12203 (N_12203,N_11965,N_11750);
xor U12204 (N_12204,N_11659,N_11768);
or U12205 (N_12205,N_11777,N_11923);
nand U12206 (N_12206,N_11896,N_11875);
or U12207 (N_12207,N_11835,N_11505);
xor U12208 (N_12208,N_11573,N_11966);
and U12209 (N_12209,N_11556,N_11932);
nand U12210 (N_12210,N_11700,N_11606);
nand U12211 (N_12211,N_11667,N_11716);
and U12212 (N_12212,N_11649,N_11684);
or U12213 (N_12213,N_11623,N_11701);
and U12214 (N_12214,N_11523,N_11801);
xnor U12215 (N_12215,N_11869,N_11968);
or U12216 (N_12216,N_11789,N_11568);
and U12217 (N_12217,N_11906,N_11723);
nand U12218 (N_12218,N_11766,N_11589);
xor U12219 (N_12219,N_11528,N_11939);
or U12220 (N_12220,N_11803,N_11576);
and U12221 (N_12221,N_11657,N_11951);
nand U12222 (N_12222,N_11913,N_11587);
and U12223 (N_12223,N_11546,N_11917);
and U12224 (N_12224,N_11852,N_11503);
and U12225 (N_12225,N_11618,N_11843);
nor U12226 (N_12226,N_11518,N_11513);
and U12227 (N_12227,N_11656,N_11709);
nand U12228 (N_12228,N_11756,N_11807);
and U12229 (N_12229,N_11625,N_11680);
and U12230 (N_12230,N_11773,N_11516);
nand U12231 (N_12231,N_11626,N_11693);
and U12232 (N_12232,N_11648,N_11810);
xnor U12233 (N_12233,N_11600,N_11504);
or U12234 (N_12234,N_11596,N_11610);
xor U12235 (N_12235,N_11817,N_11603);
nor U12236 (N_12236,N_11645,N_11722);
nor U12237 (N_12237,N_11943,N_11719);
or U12238 (N_12238,N_11779,N_11619);
nand U12239 (N_12239,N_11696,N_11774);
nor U12240 (N_12240,N_11536,N_11940);
or U12241 (N_12241,N_11646,N_11628);
nand U12242 (N_12242,N_11971,N_11887);
or U12243 (N_12243,N_11962,N_11658);
nor U12244 (N_12244,N_11575,N_11634);
nand U12245 (N_12245,N_11827,N_11559);
and U12246 (N_12246,N_11948,N_11572);
nand U12247 (N_12247,N_11979,N_11671);
and U12248 (N_12248,N_11561,N_11903);
nor U12249 (N_12249,N_11748,N_11776);
nand U12250 (N_12250,N_11773,N_11588);
and U12251 (N_12251,N_11561,N_11810);
xor U12252 (N_12252,N_11843,N_11637);
nor U12253 (N_12253,N_11828,N_11690);
xnor U12254 (N_12254,N_11510,N_11511);
xor U12255 (N_12255,N_11718,N_11761);
nand U12256 (N_12256,N_11901,N_11820);
and U12257 (N_12257,N_11534,N_11736);
nand U12258 (N_12258,N_11867,N_11921);
xor U12259 (N_12259,N_11614,N_11769);
and U12260 (N_12260,N_11613,N_11728);
nand U12261 (N_12261,N_11783,N_11856);
nor U12262 (N_12262,N_11870,N_11834);
nor U12263 (N_12263,N_11726,N_11684);
and U12264 (N_12264,N_11732,N_11736);
nand U12265 (N_12265,N_11536,N_11541);
nand U12266 (N_12266,N_11666,N_11953);
or U12267 (N_12267,N_11754,N_11794);
nand U12268 (N_12268,N_11580,N_11522);
nor U12269 (N_12269,N_11926,N_11595);
nor U12270 (N_12270,N_11708,N_11625);
nand U12271 (N_12271,N_11884,N_11711);
xnor U12272 (N_12272,N_11950,N_11747);
or U12273 (N_12273,N_11670,N_11945);
or U12274 (N_12274,N_11962,N_11765);
nand U12275 (N_12275,N_11581,N_11611);
nand U12276 (N_12276,N_11863,N_11941);
and U12277 (N_12277,N_11873,N_11805);
xor U12278 (N_12278,N_11950,N_11843);
or U12279 (N_12279,N_11940,N_11803);
nor U12280 (N_12280,N_11776,N_11963);
nor U12281 (N_12281,N_11980,N_11967);
nand U12282 (N_12282,N_11507,N_11948);
nor U12283 (N_12283,N_11675,N_11704);
xnor U12284 (N_12284,N_11838,N_11521);
nor U12285 (N_12285,N_11968,N_11855);
or U12286 (N_12286,N_11655,N_11530);
or U12287 (N_12287,N_11837,N_11596);
xor U12288 (N_12288,N_11549,N_11890);
nor U12289 (N_12289,N_11537,N_11656);
nand U12290 (N_12290,N_11630,N_11526);
xnor U12291 (N_12291,N_11694,N_11708);
xnor U12292 (N_12292,N_11699,N_11826);
or U12293 (N_12293,N_11514,N_11717);
nand U12294 (N_12294,N_11519,N_11576);
or U12295 (N_12295,N_11641,N_11571);
nand U12296 (N_12296,N_11953,N_11593);
nand U12297 (N_12297,N_11878,N_11881);
nand U12298 (N_12298,N_11950,N_11641);
or U12299 (N_12299,N_11638,N_11926);
or U12300 (N_12300,N_11978,N_11673);
nand U12301 (N_12301,N_11653,N_11560);
nor U12302 (N_12302,N_11623,N_11656);
or U12303 (N_12303,N_11984,N_11975);
nor U12304 (N_12304,N_11696,N_11723);
nand U12305 (N_12305,N_11619,N_11842);
xor U12306 (N_12306,N_11576,N_11536);
nand U12307 (N_12307,N_11508,N_11605);
nand U12308 (N_12308,N_11872,N_11580);
nand U12309 (N_12309,N_11557,N_11771);
nor U12310 (N_12310,N_11589,N_11677);
nor U12311 (N_12311,N_11660,N_11980);
nand U12312 (N_12312,N_11548,N_11619);
or U12313 (N_12313,N_11657,N_11796);
nor U12314 (N_12314,N_11524,N_11991);
nand U12315 (N_12315,N_11513,N_11692);
or U12316 (N_12316,N_11927,N_11807);
nand U12317 (N_12317,N_11829,N_11573);
nor U12318 (N_12318,N_11515,N_11651);
xnor U12319 (N_12319,N_11746,N_11542);
nand U12320 (N_12320,N_11779,N_11976);
nor U12321 (N_12321,N_11743,N_11671);
nand U12322 (N_12322,N_11938,N_11882);
xor U12323 (N_12323,N_11973,N_11975);
and U12324 (N_12324,N_11699,N_11509);
nor U12325 (N_12325,N_11645,N_11650);
nand U12326 (N_12326,N_11657,N_11952);
and U12327 (N_12327,N_11958,N_11615);
xnor U12328 (N_12328,N_11674,N_11672);
xor U12329 (N_12329,N_11571,N_11545);
nand U12330 (N_12330,N_11639,N_11936);
or U12331 (N_12331,N_11542,N_11799);
or U12332 (N_12332,N_11661,N_11949);
xor U12333 (N_12333,N_11631,N_11611);
nand U12334 (N_12334,N_11839,N_11552);
nor U12335 (N_12335,N_11512,N_11522);
and U12336 (N_12336,N_11858,N_11768);
nand U12337 (N_12337,N_11502,N_11907);
nor U12338 (N_12338,N_11669,N_11969);
and U12339 (N_12339,N_11986,N_11947);
or U12340 (N_12340,N_11708,N_11587);
nand U12341 (N_12341,N_11701,N_11566);
or U12342 (N_12342,N_11745,N_11621);
xor U12343 (N_12343,N_11813,N_11530);
xor U12344 (N_12344,N_11539,N_11623);
and U12345 (N_12345,N_11908,N_11828);
xnor U12346 (N_12346,N_11936,N_11724);
nand U12347 (N_12347,N_11827,N_11816);
nor U12348 (N_12348,N_11811,N_11715);
nor U12349 (N_12349,N_11509,N_11748);
and U12350 (N_12350,N_11570,N_11573);
xnor U12351 (N_12351,N_11628,N_11991);
nand U12352 (N_12352,N_11708,N_11942);
or U12353 (N_12353,N_11651,N_11906);
nand U12354 (N_12354,N_11635,N_11507);
nand U12355 (N_12355,N_11908,N_11533);
nor U12356 (N_12356,N_11690,N_11939);
and U12357 (N_12357,N_11877,N_11516);
nand U12358 (N_12358,N_11802,N_11647);
nand U12359 (N_12359,N_11551,N_11575);
or U12360 (N_12360,N_11956,N_11707);
xnor U12361 (N_12361,N_11688,N_11599);
nor U12362 (N_12362,N_11598,N_11652);
or U12363 (N_12363,N_11662,N_11943);
nor U12364 (N_12364,N_11678,N_11858);
nor U12365 (N_12365,N_11744,N_11692);
and U12366 (N_12366,N_11598,N_11802);
and U12367 (N_12367,N_11923,N_11694);
xor U12368 (N_12368,N_11918,N_11681);
xor U12369 (N_12369,N_11743,N_11697);
nor U12370 (N_12370,N_11575,N_11638);
nand U12371 (N_12371,N_11578,N_11561);
xnor U12372 (N_12372,N_11762,N_11904);
xor U12373 (N_12373,N_11771,N_11831);
or U12374 (N_12374,N_11646,N_11742);
and U12375 (N_12375,N_11904,N_11547);
and U12376 (N_12376,N_11551,N_11610);
nor U12377 (N_12377,N_11575,N_11935);
or U12378 (N_12378,N_11528,N_11966);
nor U12379 (N_12379,N_11837,N_11896);
or U12380 (N_12380,N_11683,N_11535);
or U12381 (N_12381,N_11860,N_11702);
and U12382 (N_12382,N_11504,N_11556);
nor U12383 (N_12383,N_11933,N_11609);
or U12384 (N_12384,N_11806,N_11656);
nand U12385 (N_12385,N_11955,N_11655);
xnor U12386 (N_12386,N_11681,N_11582);
nor U12387 (N_12387,N_11578,N_11725);
and U12388 (N_12388,N_11969,N_11854);
and U12389 (N_12389,N_11674,N_11715);
nor U12390 (N_12390,N_11769,N_11925);
nand U12391 (N_12391,N_11882,N_11934);
xnor U12392 (N_12392,N_11664,N_11736);
nor U12393 (N_12393,N_11775,N_11825);
xnor U12394 (N_12394,N_11648,N_11670);
nor U12395 (N_12395,N_11807,N_11739);
xor U12396 (N_12396,N_11684,N_11897);
or U12397 (N_12397,N_11878,N_11793);
nand U12398 (N_12398,N_11999,N_11716);
xor U12399 (N_12399,N_11697,N_11679);
xor U12400 (N_12400,N_11880,N_11894);
or U12401 (N_12401,N_11599,N_11684);
nor U12402 (N_12402,N_11806,N_11874);
xnor U12403 (N_12403,N_11847,N_11540);
and U12404 (N_12404,N_11754,N_11750);
or U12405 (N_12405,N_11942,N_11783);
and U12406 (N_12406,N_11944,N_11779);
or U12407 (N_12407,N_11643,N_11508);
nor U12408 (N_12408,N_11833,N_11602);
and U12409 (N_12409,N_11593,N_11963);
and U12410 (N_12410,N_11907,N_11906);
xor U12411 (N_12411,N_11913,N_11918);
and U12412 (N_12412,N_11816,N_11738);
and U12413 (N_12413,N_11560,N_11524);
and U12414 (N_12414,N_11858,N_11762);
nor U12415 (N_12415,N_11766,N_11963);
nor U12416 (N_12416,N_11990,N_11886);
xor U12417 (N_12417,N_11760,N_11518);
or U12418 (N_12418,N_11675,N_11598);
or U12419 (N_12419,N_11940,N_11735);
nand U12420 (N_12420,N_11561,N_11545);
nand U12421 (N_12421,N_11900,N_11895);
or U12422 (N_12422,N_11882,N_11988);
and U12423 (N_12423,N_11793,N_11515);
and U12424 (N_12424,N_11734,N_11732);
and U12425 (N_12425,N_11608,N_11540);
nor U12426 (N_12426,N_11671,N_11770);
nand U12427 (N_12427,N_11761,N_11650);
nand U12428 (N_12428,N_11734,N_11962);
and U12429 (N_12429,N_11664,N_11923);
nand U12430 (N_12430,N_11651,N_11956);
xnor U12431 (N_12431,N_11715,N_11575);
or U12432 (N_12432,N_11886,N_11759);
nand U12433 (N_12433,N_11597,N_11950);
and U12434 (N_12434,N_11667,N_11982);
and U12435 (N_12435,N_11582,N_11949);
or U12436 (N_12436,N_11647,N_11537);
nand U12437 (N_12437,N_11606,N_11544);
nor U12438 (N_12438,N_11762,N_11818);
and U12439 (N_12439,N_11983,N_11849);
and U12440 (N_12440,N_11968,N_11540);
xor U12441 (N_12441,N_11642,N_11872);
nor U12442 (N_12442,N_11524,N_11564);
xnor U12443 (N_12443,N_11689,N_11741);
xnor U12444 (N_12444,N_11629,N_11839);
nor U12445 (N_12445,N_11526,N_11694);
and U12446 (N_12446,N_11756,N_11698);
and U12447 (N_12447,N_11737,N_11621);
or U12448 (N_12448,N_11962,N_11762);
xor U12449 (N_12449,N_11853,N_11744);
or U12450 (N_12450,N_11690,N_11604);
nor U12451 (N_12451,N_11673,N_11629);
and U12452 (N_12452,N_11769,N_11627);
xor U12453 (N_12453,N_11554,N_11630);
and U12454 (N_12454,N_11780,N_11808);
and U12455 (N_12455,N_11767,N_11546);
xor U12456 (N_12456,N_11830,N_11551);
xnor U12457 (N_12457,N_11573,N_11696);
and U12458 (N_12458,N_11907,N_11635);
or U12459 (N_12459,N_11714,N_11891);
xor U12460 (N_12460,N_11736,N_11652);
and U12461 (N_12461,N_11644,N_11642);
xor U12462 (N_12462,N_11506,N_11795);
nor U12463 (N_12463,N_11589,N_11956);
nor U12464 (N_12464,N_11784,N_11909);
nor U12465 (N_12465,N_11552,N_11687);
and U12466 (N_12466,N_11920,N_11700);
and U12467 (N_12467,N_11942,N_11642);
nand U12468 (N_12468,N_11583,N_11913);
nand U12469 (N_12469,N_11988,N_11846);
xnor U12470 (N_12470,N_11831,N_11979);
or U12471 (N_12471,N_11921,N_11699);
xnor U12472 (N_12472,N_11877,N_11914);
and U12473 (N_12473,N_11854,N_11769);
xnor U12474 (N_12474,N_11663,N_11569);
nand U12475 (N_12475,N_11870,N_11913);
or U12476 (N_12476,N_11960,N_11968);
nand U12477 (N_12477,N_11605,N_11801);
xnor U12478 (N_12478,N_11563,N_11724);
xor U12479 (N_12479,N_11847,N_11528);
xnor U12480 (N_12480,N_11901,N_11684);
nor U12481 (N_12481,N_11609,N_11903);
and U12482 (N_12482,N_11890,N_11649);
xor U12483 (N_12483,N_11640,N_11542);
nand U12484 (N_12484,N_11587,N_11648);
nand U12485 (N_12485,N_11839,N_11966);
nor U12486 (N_12486,N_11545,N_11749);
nand U12487 (N_12487,N_11708,N_11915);
xnor U12488 (N_12488,N_11589,N_11779);
nor U12489 (N_12489,N_11519,N_11714);
nor U12490 (N_12490,N_11864,N_11752);
xnor U12491 (N_12491,N_11640,N_11841);
nor U12492 (N_12492,N_11800,N_11989);
and U12493 (N_12493,N_11853,N_11612);
xor U12494 (N_12494,N_11563,N_11575);
and U12495 (N_12495,N_11787,N_11928);
nand U12496 (N_12496,N_11556,N_11790);
xnor U12497 (N_12497,N_11767,N_11544);
nand U12498 (N_12498,N_11629,N_11907);
nand U12499 (N_12499,N_11714,N_11643);
or U12500 (N_12500,N_12249,N_12244);
nor U12501 (N_12501,N_12356,N_12002);
or U12502 (N_12502,N_12323,N_12490);
nand U12503 (N_12503,N_12303,N_12499);
xor U12504 (N_12504,N_12487,N_12101);
nand U12505 (N_12505,N_12191,N_12429);
nand U12506 (N_12506,N_12325,N_12371);
nand U12507 (N_12507,N_12478,N_12098);
xor U12508 (N_12508,N_12354,N_12068);
or U12509 (N_12509,N_12165,N_12364);
nor U12510 (N_12510,N_12352,N_12294);
xnor U12511 (N_12511,N_12351,N_12146);
or U12512 (N_12512,N_12015,N_12187);
nor U12513 (N_12513,N_12466,N_12105);
or U12514 (N_12514,N_12327,N_12476);
nand U12515 (N_12515,N_12344,N_12275);
nor U12516 (N_12516,N_12086,N_12217);
xor U12517 (N_12517,N_12047,N_12407);
xnor U12518 (N_12518,N_12130,N_12374);
nand U12519 (N_12519,N_12291,N_12247);
xor U12520 (N_12520,N_12106,N_12180);
xor U12521 (N_12521,N_12234,N_12428);
or U12522 (N_12522,N_12363,N_12329);
and U12523 (N_12523,N_12052,N_12111);
or U12524 (N_12524,N_12056,N_12383);
nor U12525 (N_12525,N_12050,N_12391);
and U12526 (N_12526,N_12142,N_12007);
nor U12527 (N_12527,N_12459,N_12250);
xor U12528 (N_12528,N_12456,N_12141);
or U12529 (N_12529,N_12372,N_12257);
and U12530 (N_12530,N_12253,N_12474);
or U12531 (N_12531,N_12166,N_12308);
or U12532 (N_12532,N_12122,N_12230);
xnor U12533 (N_12533,N_12023,N_12379);
nand U12534 (N_12534,N_12151,N_12183);
xor U12535 (N_12535,N_12337,N_12335);
xnor U12536 (N_12536,N_12302,N_12232);
nor U12537 (N_12537,N_12212,N_12132);
and U12538 (N_12538,N_12357,N_12353);
xnor U12539 (N_12539,N_12158,N_12013);
and U12540 (N_12540,N_12346,N_12081);
nor U12541 (N_12541,N_12279,N_12358);
xor U12542 (N_12542,N_12274,N_12286);
nor U12543 (N_12543,N_12322,N_12037);
or U12544 (N_12544,N_12376,N_12091);
and U12545 (N_12545,N_12173,N_12485);
nand U12546 (N_12546,N_12160,N_12243);
nand U12547 (N_12547,N_12398,N_12450);
xnor U12548 (N_12548,N_12432,N_12215);
and U12549 (N_12549,N_12276,N_12287);
xnor U12550 (N_12550,N_12318,N_12320);
or U12551 (N_12551,N_12139,N_12186);
nor U12552 (N_12552,N_12126,N_12107);
xnor U12553 (N_12553,N_12345,N_12155);
or U12554 (N_12554,N_12316,N_12467);
and U12555 (N_12555,N_12197,N_12266);
nand U12556 (N_12556,N_12283,N_12022);
nor U12557 (N_12557,N_12159,N_12133);
nand U12558 (N_12558,N_12334,N_12076);
nor U12559 (N_12559,N_12468,N_12348);
or U12560 (N_12560,N_12156,N_12324);
nand U12561 (N_12561,N_12462,N_12451);
nand U12562 (N_12562,N_12410,N_12072);
xor U12563 (N_12563,N_12425,N_12472);
and U12564 (N_12564,N_12099,N_12486);
xnor U12565 (N_12565,N_12108,N_12009);
and U12566 (N_12566,N_12365,N_12268);
or U12567 (N_12567,N_12033,N_12110);
nor U12568 (N_12568,N_12413,N_12393);
nor U12569 (N_12569,N_12220,N_12092);
xor U12570 (N_12570,N_12058,N_12078);
or U12571 (N_12571,N_12103,N_12304);
and U12572 (N_12572,N_12359,N_12039);
or U12573 (N_12573,N_12347,N_12460);
or U12574 (N_12574,N_12241,N_12458);
or U12575 (N_12575,N_12027,N_12182);
nand U12576 (N_12576,N_12388,N_12259);
nand U12577 (N_12577,N_12066,N_12470);
nand U12578 (N_12578,N_12043,N_12317);
nor U12579 (N_12579,N_12307,N_12190);
nand U12580 (N_12580,N_12069,N_12455);
nor U12581 (N_12581,N_12404,N_12332);
nor U12582 (N_12582,N_12164,N_12201);
xnor U12583 (N_12583,N_12127,N_12427);
and U12584 (N_12584,N_12284,N_12071);
xor U12585 (N_12585,N_12349,N_12040);
and U12586 (N_12586,N_12477,N_12178);
nand U12587 (N_12587,N_12029,N_12239);
and U12588 (N_12588,N_12342,N_12436);
xor U12589 (N_12589,N_12113,N_12447);
nand U12590 (N_12590,N_12479,N_12157);
nand U12591 (N_12591,N_12063,N_12445);
nor U12592 (N_12592,N_12385,N_12480);
xnor U12593 (N_12593,N_12100,N_12331);
xnor U12594 (N_12594,N_12211,N_12179);
or U12595 (N_12595,N_12090,N_12340);
nand U12596 (N_12596,N_12366,N_12134);
nand U12597 (N_12597,N_12369,N_12226);
nand U12598 (N_12598,N_12281,N_12395);
nor U12599 (N_12599,N_12278,N_12489);
or U12600 (N_12600,N_12271,N_12300);
and U12601 (N_12601,N_12321,N_12272);
nor U12602 (N_12602,N_12403,N_12394);
nor U12603 (N_12603,N_12494,N_12319);
nand U12604 (N_12604,N_12198,N_12038);
nor U12605 (N_12605,N_12204,N_12292);
xnor U12606 (N_12606,N_12075,N_12073);
xnor U12607 (N_12607,N_12061,N_12418);
and U12608 (N_12608,N_12210,N_12030);
xor U12609 (N_12609,N_12233,N_12341);
or U12610 (N_12610,N_12434,N_12207);
xor U12611 (N_12611,N_12355,N_12282);
nor U12612 (N_12612,N_12012,N_12417);
nand U12613 (N_12613,N_12227,N_12299);
or U12614 (N_12614,N_12054,N_12312);
nor U12615 (N_12615,N_12188,N_12154);
and U12616 (N_12616,N_12016,N_12412);
nor U12617 (N_12617,N_12229,N_12449);
and U12618 (N_12618,N_12017,N_12021);
or U12619 (N_12619,N_12116,N_12301);
or U12620 (N_12620,N_12441,N_12121);
or U12621 (N_12621,N_12044,N_12175);
nor U12622 (N_12622,N_12392,N_12454);
nand U12623 (N_12623,N_12004,N_12491);
nor U12624 (N_12624,N_12032,N_12067);
and U12625 (N_12625,N_12419,N_12048);
nor U12626 (N_12626,N_12095,N_12083);
xnor U12627 (N_12627,N_12438,N_12123);
and U12628 (N_12628,N_12034,N_12085);
or U12629 (N_12629,N_12255,N_12059);
nand U12630 (N_12630,N_12203,N_12473);
or U12631 (N_12631,N_12254,N_12339);
nor U12632 (N_12632,N_12435,N_12138);
nand U12633 (N_12633,N_12416,N_12382);
or U12634 (N_12634,N_12296,N_12350);
or U12635 (N_12635,N_12326,N_12084);
nand U12636 (N_12636,N_12010,N_12036);
or U12637 (N_12637,N_12446,N_12169);
or U12638 (N_12638,N_12225,N_12192);
nor U12639 (N_12639,N_12137,N_12181);
nand U12640 (N_12640,N_12368,N_12475);
and U12641 (N_12641,N_12170,N_12439);
nor U12642 (N_12642,N_12080,N_12492);
and U12643 (N_12643,N_12177,N_12338);
nand U12644 (N_12644,N_12430,N_12252);
nor U12645 (N_12645,N_12117,N_12223);
xor U12646 (N_12646,N_12094,N_12251);
nor U12647 (N_12647,N_12129,N_12104);
and U12648 (N_12648,N_12461,N_12463);
nor U12649 (N_12649,N_12415,N_12144);
xnor U12650 (N_12650,N_12168,N_12024);
xnor U12651 (N_12651,N_12031,N_12314);
nor U12652 (N_12652,N_12102,N_12196);
and U12653 (N_12653,N_12262,N_12049);
nor U12654 (N_12654,N_12114,N_12235);
nor U12655 (N_12655,N_12424,N_12184);
nor U12656 (N_12656,N_12045,N_12484);
nand U12657 (N_12657,N_12057,N_12008);
or U12658 (N_12658,N_12026,N_12493);
nor U12659 (N_12659,N_12495,N_12402);
nand U12660 (N_12660,N_12443,N_12444);
nand U12661 (N_12661,N_12246,N_12228);
and U12662 (N_12662,N_12360,N_12224);
xor U12663 (N_12663,N_12497,N_12200);
nor U12664 (N_12664,N_12280,N_12150);
nand U12665 (N_12665,N_12258,N_12149);
or U12666 (N_12666,N_12311,N_12136);
or U12667 (N_12667,N_12310,N_12315);
and U12668 (N_12668,N_12119,N_12089);
nor U12669 (N_12669,N_12199,N_12448);
or U12670 (N_12670,N_12167,N_12483);
and U12671 (N_12671,N_12336,N_12264);
xor U12672 (N_12672,N_12361,N_12375);
or U12673 (N_12673,N_12147,N_12112);
and U12674 (N_12674,N_12028,N_12140);
xnor U12675 (N_12675,N_12285,N_12118);
nand U12676 (N_12676,N_12143,N_12426);
nand U12677 (N_12677,N_12409,N_12163);
nand U12678 (N_12678,N_12390,N_12482);
xor U12679 (N_12679,N_12011,N_12380);
xor U12680 (N_12680,N_12437,N_12452);
nor U12681 (N_12681,N_12263,N_12219);
and U12682 (N_12682,N_12189,N_12305);
or U12683 (N_12683,N_12046,N_12373);
and U12684 (N_12684,N_12384,N_12408);
nor U12685 (N_12685,N_12270,N_12135);
and U12686 (N_12686,N_12464,N_12306);
xor U12687 (N_12687,N_12465,N_12120);
xnor U12688 (N_12688,N_12498,N_12025);
nand U12689 (N_12689,N_12273,N_12422);
xor U12690 (N_12690,N_12269,N_12381);
nand U12691 (N_12691,N_12209,N_12145);
nor U12692 (N_12692,N_12218,N_12148);
xnor U12693 (N_12693,N_12289,N_12205);
xor U12694 (N_12694,N_12064,N_12313);
xor U12695 (N_12695,N_12041,N_12193);
nand U12696 (N_12696,N_12256,N_12082);
and U12697 (N_12697,N_12236,N_12242);
nand U12698 (N_12698,N_12330,N_12496);
nand U12699 (N_12699,N_12265,N_12411);
or U12700 (N_12700,N_12221,N_12488);
nand U12701 (N_12701,N_12020,N_12077);
and U12702 (N_12702,N_12387,N_12000);
and U12703 (N_12703,N_12328,N_12096);
nor U12704 (N_12704,N_12019,N_12214);
and U12705 (N_12705,N_12288,N_12295);
nor U12706 (N_12706,N_12062,N_12290);
nand U12707 (N_12707,N_12124,N_12400);
or U12708 (N_12708,N_12362,N_12001);
or U12709 (N_12709,N_12471,N_12006);
and U12710 (N_12710,N_12277,N_12005);
xnor U12711 (N_12711,N_12297,N_12261);
nor U12712 (N_12712,N_12216,N_12237);
and U12713 (N_12713,N_12042,N_12298);
nand U12714 (N_12714,N_12405,N_12240);
and U12715 (N_12715,N_12213,N_12194);
and U12716 (N_12716,N_12195,N_12453);
and U12717 (N_12717,N_12293,N_12386);
nand U12718 (N_12718,N_12065,N_12389);
nand U12719 (N_12719,N_12333,N_12035);
nand U12720 (N_12720,N_12079,N_12014);
and U12721 (N_12721,N_12469,N_12172);
xnor U12722 (N_12722,N_12442,N_12431);
and U12723 (N_12723,N_12399,N_12185);
or U12724 (N_12724,N_12003,N_12074);
nor U12725 (N_12725,N_12208,N_12267);
nor U12726 (N_12726,N_12051,N_12171);
nand U12727 (N_12727,N_12421,N_12433);
nand U12728 (N_12728,N_12131,N_12174);
nand U12729 (N_12729,N_12162,N_12070);
or U12730 (N_12730,N_12245,N_12088);
or U12731 (N_12731,N_12440,N_12396);
and U12732 (N_12732,N_12238,N_12053);
nor U12733 (N_12733,N_12377,N_12260);
and U12734 (N_12734,N_12343,N_12367);
xor U12735 (N_12735,N_12378,N_12153);
nor U12736 (N_12736,N_12093,N_12097);
and U12737 (N_12737,N_12152,N_12125);
xor U12738 (N_12738,N_12206,N_12231);
xor U12739 (N_12739,N_12420,N_12414);
or U12740 (N_12740,N_12018,N_12161);
or U12741 (N_12741,N_12406,N_12055);
and U12742 (N_12742,N_12401,N_12397);
nor U12743 (N_12743,N_12370,N_12309);
and U12744 (N_12744,N_12457,N_12115);
nor U12745 (N_12745,N_12248,N_12087);
xnor U12746 (N_12746,N_12176,N_12423);
or U12747 (N_12747,N_12222,N_12109);
nand U12748 (N_12748,N_12060,N_12202);
or U12749 (N_12749,N_12128,N_12481);
and U12750 (N_12750,N_12476,N_12368);
xor U12751 (N_12751,N_12336,N_12212);
nand U12752 (N_12752,N_12457,N_12316);
or U12753 (N_12753,N_12006,N_12161);
and U12754 (N_12754,N_12253,N_12048);
and U12755 (N_12755,N_12431,N_12481);
xor U12756 (N_12756,N_12142,N_12259);
nor U12757 (N_12757,N_12215,N_12048);
or U12758 (N_12758,N_12392,N_12396);
and U12759 (N_12759,N_12100,N_12181);
or U12760 (N_12760,N_12080,N_12153);
and U12761 (N_12761,N_12202,N_12270);
and U12762 (N_12762,N_12265,N_12447);
xor U12763 (N_12763,N_12260,N_12152);
or U12764 (N_12764,N_12125,N_12433);
or U12765 (N_12765,N_12108,N_12432);
and U12766 (N_12766,N_12402,N_12162);
and U12767 (N_12767,N_12015,N_12196);
xnor U12768 (N_12768,N_12351,N_12482);
and U12769 (N_12769,N_12281,N_12292);
and U12770 (N_12770,N_12117,N_12013);
nand U12771 (N_12771,N_12050,N_12133);
or U12772 (N_12772,N_12344,N_12166);
or U12773 (N_12773,N_12179,N_12101);
nand U12774 (N_12774,N_12234,N_12009);
xnor U12775 (N_12775,N_12406,N_12209);
xnor U12776 (N_12776,N_12231,N_12033);
xnor U12777 (N_12777,N_12451,N_12198);
and U12778 (N_12778,N_12093,N_12460);
nand U12779 (N_12779,N_12167,N_12349);
nor U12780 (N_12780,N_12160,N_12335);
and U12781 (N_12781,N_12316,N_12232);
nand U12782 (N_12782,N_12452,N_12314);
xnor U12783 (N_12783,N_12076,N_12034);
nor U12784 (N_12784,N_12273,N_12050);
or U12785 (N_12785,N_12297,N_12136);
nor U12786 (N_12786,N_12422,N_12203);
nand U12787 (N_12787,N_12498,N_12326);
or U12788 (N_12788,N_12170,N_12036);
xor U12789 (N_12789,N_12312,N_12300);
xnor U12790 (N_12790,N_12271,N_12422);
nand U12791 (N_12791,N_12482,N_12326);
nand U12792 (N_12792,N_12188,N_12255);
xnor U12793 (N_12793,N_12266,N_12078);
nand U12794 (N_12794,N_12261,N_12018);
nor U12795 (N_12795,N_12370,N_12431);
and U12796 (N_12796,N_12009,N_12485);
nor U12797 (N_12797,N_12245,N_12432);
nor U12798 (N_12798,N_12294,N_12213);
and U12799 (N_12799,N_12311,N_12280);
and U12800 (N_12800,N_12030,N_12397);
nor U12801 (N_12801,N_12007,N_12185);
xnor U12802 (N_12802,N_12263,N_12010);
or U12803 (N_12803,N_12304,N_12261);
xor U12804 (N_12804,N_12367,N_12100);
nor U12805 (N_12805,N_12401,N_12366);
nand U12806 (N_12806,N_12048,N_12272);
nand U12807 (N_12807,N_12034,N_12154);
or U12808 (N_12808,N_12330,N_12294);
and U12809 (N_12809,N_12437,N_12315);
nand U12810 (N_12810,N_12140,N_12023);
xnor U12811 (N_12811,N_12166,N_12316);
and U12812 (N_12812,N_12385,N_12075);
nor U12813 (N_12813,N_12322,N_12052);
or U12814 (N_12814,N_12419,N_12154);
nand U12815 (N_12815,N_12297,N_12087);
xnor U12816 (N_12816,N_12071,N_12156);
or U12817 (N_12817,N_12293,N_12328);
nand U12818 (N_12818,N_12303,N_12401);
or U12819 (N_12819,N_12102,N_12084);
nand U12820 (N_12820,N_12402,N_12249);
and U12821 (N_12821,N_12154,N_12128);
xnor U12822 (N_12822,N_12040,N_12167);
xnor U12823 (N_12823,N_12468,N_12077);
nor U12824 (N_12824,N_12209,N_12480);
xor U12825 (N_12825,N_12029,N_12418);
and U12826 (N_12826,N_12216,N_12103);
nand U12827 (N_12827,N_12340,N_12326);
xnor U12828 (N_12828,N_12189,N_12149);
xnor U12829 (N_12829,N_12031,N_12470);
xnor U12830 (N_12830,N_12179,N_12425);
or U12831 (N_12831,N_12279,N_12168);
nand U12832 (N_12832,N_12208,N_12426);
nor U12833 (N_12833,N_12179,N_12111);
xor U12834 (N_12834,N_12197,N_12409);
and U12835 (N_12835,N_12472,N_12298);
nand U12836 (N_12836,N_12347,N_12080);
or U12837 (N_12837,N_12470,N_12239);
nor U12838 (N_12838,N_12075,N_12405);
and U12839 (N_12839,N_12242,N_12469);
xnor U12840 (N_12840,N_12227,N_12201);
nand U12841 (N_12841,N_12475,N_12434);
xnor U12842 (N_12842,N_12099,N_12004);
xor U12843 (N_12843,N_12125,N_12495);
nor U12844 (N_12844,N_12012,N_12066);
nand U12845 (N_12845,N_12071,N_12197);
xor U12846 (N_12846,N_12496,N_12368);
and U12847 (N_12847,N_12492,N_12232);
and U12848 (N_12848,N_12279,N_12310);
nand U12849 (N_12849,N_12385,N_12177);
or U12850 (N_12850,N_12184,N_12445);
xor U12851 (N_12851,N_12037,N_12162);
nor U12852 (N_12852,N_12426,N_12021);
xnor U12853 (N_12853,N_12138,N_12475);
nand U12854 (N_12854,N_12088,N_12427);
or U12855 (N_12855,N_12466,N_12149);
or U12856 (N_12856,N_12488,N_12405);
and U12857 (N_12857,N_12233,N_12122);
nand U12858 (N_12858,N_12141,N_12239);
nand U12859 (N_12859,N_12350,N_12266);
nor U12860 (N_12860,N_12058,N_12157);
or U12861 (N_12861,N_12496,N_12143);
and U12862 (N_12862,N_12441,N_12183);
or U12863 (N_12863,N_12466,N_12498);
xnor U12864 (N_12864,N_12235,N_12243);
nand U12865 (N_12865,N_12048,N_12324);
or U12866 (N_12866,N_12429,N_12023);
or U12867 (N_12867,N_12111,N_12010);
xor U12868 (N_12868,N_12057,N_12193);
or U12869 (N_12869,N_12332,N_12097);
nand U12870 (N_12870,N_12356,N_12474);
xor U12871 (N_12871,N_12437,N_12081);
or U12872 (N_12872,N_12175,N_12204);
xnor U12873 (N_12873,N_12293,N_12167);
nor U12874 (N_12874,N_12493,N_12451);
and U12875 (N_12875,N_12337,N_12039);
xor U12876 (N_12876,N_12170,N_12133);
nand U12877 (N_12877,N_12348,N_12177);
or U12878 (N_12878,N_12004,N_12459);
nand U12879 (N_12879,N_12067,N_12147);
nand U12880 (N_12880,N_12247,N_12064);
and U12881 (N_12881,N_12164,N_12002);
xor U12882 (N_12882,N_12497,N_12392);
or U12883 (N_12883,N_12053,N_12477);
and U12884 (N_12884,N_12179,N_12149);
or U12885 (N_12885,N_12154,N_12088);
or U12886 (N_12886,N_12317,N_12420);
nand U12887 (N_12887,N_12341,N_12149);
or U12888 (N_12888,N_12410,N_12157);
and U12889 (N_12889,N_12402,N_12481);
nand U12890 (N_12890,N_12041,N_12149);
and U12891 (N_12891,N_12295,N_12055);
xnor U12892 (N_12892,N_12137,N_12209);
and U12893 (N_12893,N_12188,N_12014);
or U12894 (N_12894,N_12223,N_12193);
nand U12895 (N_12895,N_12135,N_12304);
nand U12896 (N_12896,N_12231,N_12273);
xor U12897 (N_12897,N_12174,N_12217);
nor U12898 (N_12898,N_12227,N_12166);
and U12899 (N_12899,N_12339,N_12186);
nand U12900 (N_12900,N_12083,N_12446);
xor U12901 (N_12901,N_12116,N_12059);
xor U12902 (N_12902,N_12152,N_12205);
or U12903 (N_12903,N_12233,N_12443);
or U12904 (N_12904,N_12298,N_12476);
xnor U12905 (N_12905,N_12155,N_12460);
xor U12906 (N_12906,N_12368,N_12115);
nand U12907 (N_12907,N_12397,N_12456);
and U12908 (N_12908,N_12432,N_12420);
xor U12909 (N_12909,N_12420,N_12154);
and U12910 (N_12910,N_12134,N_12494);
and U12911 (N_12911,N_12390,N_12408);
xor U12912 (N_12912,N_12286,N_12235);
xor U12913 (N_12913,N_12357,N_12467);
nor U12914 (N_12914,N_12386,N_12172);
nand U12915 (N_12915,N_12241,N_12486);
or U12916 (N_12916,N_12295,N_12106);
nor U12917 (N_12917,N_12192,N_12074);
nor U12918 (N_12918,N_12066,N_12017);
or U12919 (N_12919,N_12217,N_12322);
nand U12920 (N_12920,N_12115,N_12159);
and U12921 (N_12921,N_12444,N_12009);
or U12922 (N_12922,N_12045,N_12039);
nand U12923 (N_12923,N_12457,N_12409);
and U12924 (N_12924,N_12457,N_12490);
nand U12925 (N_12925,N_12352,N_12416);
or U12926 (N_12926,N_12238,N_12082);
xnor U12927 (N_12927,N_12356,N_12042);
xnor U12928 (N_12928,N_12429,N_12368);
and U12929 (N_12929,N_12269,N_12480);
and U12930 (N_12930,N_12044,N_12012);
nor U12931 (N_12931,N_12456,N_12457);
xor U12932 (N_12932,N_12134,N_12354);
and U12933 (N_12933,N_12142,N_12398);
and U12934 (N_12934,N_12230,N_12326);
or U12935 (N_12935,N_12358,N_12382);
or U12936 (N_12936,N_12476,N_12145);
and U12937 (N_12937,N_12291,N_12060);
xor U12938 (N_12938,N_12348,N_12322);
nor U12939 (N_12939,N_12077,N_12314);
nor U12940 (N_12940,N_12020,N_12424);
nand U12941 (N_12941,N_12129,N_12469);
nand U12942 (N_12942,N_12144,N_12457);
xnor U12943 (N_12943,N_12003,N_12015);
xnor U12944 (N_12944,N_12485,N_12291);
xnor U12945 (N_12945,N_12437,N_12174);
xnor U12946 (N_12946,N_12279,N_12192);
nand U12947 (N_12947,N_12113,N_12230);
xnor U12948 (N_12948,N_12007,N_12421);
or U12949 (N_12949,N_12336,N_12318);
nand U12950 (N_12950,N_12322,N_12116);
xor U12951 (N_12951,N_12410,N_12053);
or U12952 (N_12952,N_12029,N_12460);
or U12953 (N_12953,N_12208,N_12049);
nand U12954 (N_12954,N_12069,N_12358);
nor U12955 (N_12955,N_12267,N_12456);
and U12956 (N_12956,N_12122,N_12021);
nor U12957 (N_12957,N_12448,N_12369);
and U12958 (N_12958,N_12445,N_12457);
nor U12959 (N_12959,N_12400,N_12380);
or U12960 (N_12960,N_12423,N_12432);
nor U12961 (N_12961,N_12426,N_12489);
xor U12962 (N_12962,N_12371,N_12488);
and U12963 (N_12963,N_12254,N_12353);
nand U12964 (N_12964,N_12111,N_12349);
nand U12965 (N_12965,N_12197,N_12239);
or U12966 (N_12966,N_12182,N_12332);
and U12967 (N_12967,N_12319,N_12364);
and U12968 (N_12968,N_12327,N_12458);
xnor U12969 (N_12969,N_12296,N_12329);
xnor U12970 (N_12970,N_12066,N_12249);
nor U12971 (N_12971,N_12223,N_12189);
xor U12972 (N_12972,N_12133,N_12181);
and U12973 (N_12973,N_12336,N_12324);
nand U12974 (N_12974,N_12475,N_12272);
xnor U12975 (N_12975,N_12411,N_12431);
or U12976 (N_12976,N_12211,N_12021);
or U12977 (N_12977,N_12059,N_12433);
nand U12978 (N_12978,N_12182,N_12266);
or U12979 (N_12979,N_12273,N_12355);
xnor U12980 (N_12980,N_12380,N_12194);
nor U12981 (N_12981,N_12307,N_12213);
xor U12982 (N_12982,N_12234,N_12034);
or U12983 (N_12983,N_12157,N_12084);
xor U12984 (N_12984,N_12141,N_12303);
and U12985 (N_12985,N_12324,N_12190);
nand U12986 (N_12986,N_12196,N_12066);
and U12987 (N_12987,N_12226,N_12100);
or U12988 (N_12988,N_12337,N_12393);
or U12989 (N_12989,N_12438,N_12406);
nor U12990 (N_12990,N_12318,N_12490);
xor U12991 (N_12991,N_12102,N_12466);
xor U12992 (N_12992,N_12354,N_12214);
and U12993 (N_12993,N_12030,N_12410);
or U12994 (N_12994,N_12009,N_12174);
nor U12995 (N_12995,N_12318,N_12334);
or U12996 (N_12996,N_12059,N_12079);
and U12997 (N_12997,N_12084,N_12266);
nor U12998 (N_12998,N_12087,N_12183);
and U12999 (N_12999,N_12456,N_12059);
nand U13000 (N_13000,N_12816,N_12667);
xnor U13001 (N_13001,N_12807,N_12805);
nand U13002 (N_13002,N_12826,N_12878);
or U13003 (N_13003,N_12517,N_12556);
or U13004 (N_13004,N_12579,N_12853);
nor U13005 (N_13005,N_12776,N_12561);
nor U13006 (N_13006,N_12958,N_12673);
and U13007 (N_13007,N_12934,N_12830);
and U13008 (N_13008,N_12941,N_12914);
and U13009 (N_13009,N_12856,N_12912);
nor U13010 (N_13010,N_12584,N_12529);
nor U13011 (N_13011,N_12705,N_12753);
nor U13012 (N_13012,N_12626,N_12659);
nor U13013 (N_13013,N_12769,N_12749);
nand U13014 (N_13014,N_12965,N_12552);
and U13015 (N_13015,N_12835,N_12797);
nand U13016 (N_13016,N_12932,N_12515);
nor U13017 (N_13017,N_12735,N_12635);
or U13018 (N_13018,N_12988,N_12569);
and U13019 (N_13019,N_12600,N_12869);
xnor U13020 (N_13020,N_12520,N_12633);
xnor U13021 (N_13021,N_12980,N_12876);
nor U13022 (N_13022,N_12512,N_12647);
xnor U13023 (N_13023,N_12592,N_12799);
and U13024 (N_13024,N_12855,N_12658);
nand U13025 (N_13025,N_12583,N_12939);
or U13026 (N_13026,N_12759,N_12565);
nor U13027 (N_13027,N_12949,N_12974);
nand U13028 (N_13028,N_12792,N_12793);
xor U13029 (N_13029,N_12587,N_12657);
or U13030 (N_13030,N_12846,N_12957);
or U13031 (N_13031,N_12930,N_12896);
nand U13032 (N_13032,N_12977,N_12599);
or U13033 (N_13033,N_12683,N_12841);
or U13034 (N_13034,N_12973,N_12865);
xor U13035 (N_13035,N_12984,N_12688);
or U13036 (N_13036,N_12595,N_12636);
xnor U13037 (N_13037,N_12811,N_12573);
or U13038 (N_13038,N_12628,N_12831);
and U13039 (N_13039,N_12610,N_12863);
and U13040 (N_13040,N_12728,N_12894);
or U13041 (N_13041,N_12603,N_12605);
or U13042 (N_13042,N_12882,N_12630);
nor U13043 (N_13043,N_12644,N_12889);
and U13044 (N_13044,N_12761,N_12677);
and U13045 (N_13045,N_12567,N_12755);
nor U13046 (N_13046,N_12666,N_12551);
or U13047 (N_13047,N_12656,N_12913);
or U13048 (N_13048,N_12664,N_12685);
or U13049 (N_13049,N_12982,N_12507);
and U13050 (N_13050,N_12686,N_12942);
and U13051 (N_13051,N_12526,N_12820);
nor U13052 (N_13052,N_12819,N_12554);
nand U13053 (N_13053,N_12506,N_12773);
nor U13054 (N_13054,N_12992,N_12682);
or U13055 (N_13055,N_12919,N_12993);
or U13056 (N_13056,N_12615,N_12585);
and U13057 (N_13057,N_12707,N_12722);
and U13058 (N_13058,N_12622,N_12589);
nand U13059 (N_13059,N_12593,N_12983);
or U13060 (N_13060,N_12618,N_12777);
and U13061 (N_13061,N_12774,N_12521);
and U13062 (N_13062,N_12756,N_12772);
and U13063 (N_13063,N_12901,N_12588);
xnor U13064 (N_13064,N_12732,N_12947);
xnor U13065 (N_13065,N_12525,N_12779);
or U13066 (N_13066,N_12864,N_12842);
or U13067 (N_13067,N_12668,N_12539);
and U13068 (N_13068,N_12638,N_12900);
xor U13069 (N_13069,N_12994,N_12717);
nand U13070 (N_13070,N_12812,N_12911);
and U13071 (N_13071,N_12870,N_12832);
or U13072 (N_13072,N_12535,N_12810);
nor U13073 (N_13073,N_12568,N_12572);
or U13074 (N_13074,N_12617,N_12940);
nor U13075 (N_13075,N_12696,N_12724);
xnor U13076 (N_13076,N_12893,N_12654);
nor U13077 (N_13077,N_12851,N_12899);
nand U13078 (N_13078,N_12933,N_12623);
xor U13079 (N_13079,N_12718,N_12743);
or U13080 (N_13080,N_12787,N_12655);
nand U13081 (N_13081,N_12500,N_12719);
or U13082 (N_13082,N_12577,N_12582);
or U13083 (N_13083,N_12680,N_12821);
nor U13084 (N_13084,N_12527,N_12996);
nand U13085 (N_13085,N_12563,N_12857);
or U13086 (N_13086,N_12860,N_12627);
and U13087 (N_13087,N_12836,N_12702);
and U13088 (N_13088,N_12604,N_12738);
or U13089 (N_13089,N_12516,N_12897);
nor U13090 (N_13090,N_12989,N_12833);
xnor U13091 (N_13091,N_12884,N_12523);
or U13092 (N_13092,N_12502,N_12642);
xnor U13093 (N_13093,N_12954,N_12736);
nand U13094 (N_13094,N_12766,N_12663);
and U13095 (N_13095,N_12951,N_12981);
and U13096 (N_13096,N_12534,N_12524);
nand U13097 (N_13097,N_12923,N_12625);
nor U13098 (N_13098,N_12910,N_12519);
nand U13099 (N_13099,N_12794,N_12538);
xnor U13100 (N_13100,N_12829,N_12621);
or U13101 (N_13101,N_12676,N_12557);
xnor U13102 (N_13102,N_12956,N_12886);
or U13103 (N_13103,N_12854,N_12731);
or U13104 (N_13104,N_12924,N_12640);
nor U13105 (N_13105,N_12990,N_12601);
nand U13106 (N_13106,N_12639,N_12918);
nor U13107 (N_13107,N_12672,N_12837);
or U13108 (N_13108,N_12687,N_12975);
nand U13109 (N_13109,N_12955,N_12745);
or U13110 (N_13110,N_12715,N_12945);
nand U13111 (N_13111,N_12750,N_12959);
nand U13112 (N_13112,N_12915,N_12969);
and U13113 (N_13113,N_12771,N_12720);
nand U13114 (N_13114,N_12818,N_12783);
nor U13115 (N_13115,N_12671,N_12691);
nor U13116 (N_13116,N_12608,N_12867);
xor U13117 (N_13117,N_12723,N_12742);
nand U13118 (N_13118,N_12961,N_12530);
xor U13119 (N_13119,N_12679,N_12948);
nor U13120 (N_13120,N_12960,N_12637);
and U13121 (N_13121,N_12692,N_12651);
nor U13122 (N_13122,N_12952,N_12727);
or U13123 (N_13123,N_12710,N_12566);
or U13124 (N_13124,N_12698,N_12646);
nor U13125 (N_13125,N_12859,N_12553);
nand U13126 (N_13126,N_12734,N_12542);
xnor U13127 (N_13127,N_12858,N_12689);
nor U13128 (N_13128,N_12614,N_12976);
or U13129 (N_13129,N_12748,N_12697);
nor U13130 (N_13130,N_12866,N_12877);
xnor U13131 (N_13131,N_12985,N_12550);
nand U13132 (N_13132,N_12574,N_12967);
or U13133 (N_13133,N_12744,N_12775);
and U13134 (N_13134,N_12536,N_12765);
or U13135 (N_13135,N_12760,N_12972);
or U13136 (N_13136,N_12558,N_12596);
nor U13137 (N_13137,N_12662,N_12547);
nand U13138 (N_13138,N_12518,N_12849);
nand U13139 (N_13139,N_12768,N_12571);
or U13140 (N_13140,N_12845,N_12806);
or U13141 (N_13141,N_12619,N_12790);
nor U13142 (N_13142,N_12950,N_12712);
xor U13143 (N_13143,N_12620,N_12559);
or U13144 (N_13144,N_12861,N_12575);
and U13145 (N_13145,N_12508,N_12580);
and U13146 (N_13146,N_12549,N_12681);
and U13147 (N_13147,N_12632,N_12704);
xnor U13148 (N_13148,N_12629,N_12796);
and U13149 (N_13149,N_12741,N_12721);
xor U13150 (N_13150,N_12645,N_12813);
nand U13151 (N_13151,N_12908,N_12822);
or U13152 (N_13152,N_12709,N_12504);
nor U13153 (N_13153,N_12528,N_12935);
or U13154 (N_13154,N_12757,N_12979);
or U13155 (N_13155,N_12986,N_12785);
and U13156 (N_13156,N_12828,N_12802);
nand U13157 (N_13157,N_12739,N_12920);
and U13158 (N_13158,N_12648,N_12544);
or U13159 (N_13159,N_12825,N_12560);
nor U13160 (N_13160,N_12888,N_12533);
or U13161 (N_13161,N_12746,N_12546);
nor U13162 (N_13162,N_12747,N_12838);
nand U13163 (N_13163,N_12781,N_12540);
or U13164 (N_13164,N_12548,N_12782);
or U13165 (N_13165,N_12740,N_12562);
xor U13166 (N_13166,N_12780,N_12624);
or U13167 (N_13167,N_12844,N_12987);
or U13168 (N_13168,N_12834,N_12902);
or U13169 (N_13169,N_12823,N_12729);
and U13170 (N_13170,N_12581,N_12602);
nor U13171 (N_13171,N_12578,N_12926);
or U13172 (N_13172,N_12611,N_12824);
nand U13173 (N_13173,N_12598,N_12670);
and U13174 (N_13174,N_12970,N_12809);
xnor U13175 (N_13175,N_12694,N_12814);
xnor U13176 (N_13176,N_12963,N_12968);
or U13177 (N_13177,N_12713,N_12532);
and U13178 (N_13178,N_12778,N_12937);
xor U13179 (N_13179,N_12669,N_12726);
nor U13180 (N_13180,N_12700,N_12762);
xnor U13181 (N_13181,N_12999,N_12883);
and U13182 (N_13182,N_12953,N_12788);
nor U13183 (N_13183,N_12699,N_12890);
nor U13184 (N_13184,N_12801,N_12752);
xor U13185 (N_13185,N_12922,N_12531);
or U13186 (N_13186,N_12716,N_12885);
nor U13187 (N_13187,N_12616,N_12800);
nand U13188 (N_13188,N_12827,N_12879);
xor U13189 (N_13189,N_12678,N_12997);
and U13190 (N_13190,N_12675,N_12652);
or U13191 (N_13191,N_12660,N_12665);
nor U13192 (N_13192,N_12505,N_12929);
or U13193 (N_13193,N_12555,N_12631);
nand U13194 (N_13194,N_12925,N_12995);
and U13195 (N_13195,N_12928,N_12962);
nand U13196 (N_13196,N_12905,N_12840);
nor U13197 (N_13197,N_12891,N_12511);
and U13198 (N_13198,N_12594,N_12541);
nor U13199 (N_13199,N_12880,N_12978);
and U13200 (N_13200,N_12971,N_12684);
and U13201 (N_13201,N_12916,N_12751);
xnor U13202 (N_13202,N_12789,N_12708);
nor U13203 (N_13203,N_12725,N_12501);
and U13204 (N_13204,N_12871,N_12808);
nor U13205 (N_13205,N_12921,N_12643);
nand U13206 (N_13206,N_12570,N_12898);
nand U13207 (N_13207,N_12873,N_12904);
nor U13208 (N_13208,N_12909,N_12703);
nor U13209 (N_13209,N_12649,N_12927);
and U13210 (N_13210,N_12695,N_12862);
and U13211 (N_13211,N_12641,N_12537);
and U13212 (N_13212,N_12804,N_12590);
nor U13213 (N_13213,N_12784,N_12564);
or U13214 (N_13214,N_12606,N_12892);
and U13215 (N_13215,N_12730,N_12881);
nor U13216 (N_13216,N_12767,N_12895);
xor U13217 (N_13217,N_12795,N_12714);
or U13218 (N_13218,N_12543,N_12903);
nand U13219 (N_13219,N_12576,N_12653);
nor U13220 (N_13220,N_12514,N_12650);
nand U13221 (N_13221,N_12907,N_12966);
xor U13222 (N_13222,N_12791,N_12938);
or U13223 (N_13223,N_12848,N_12711);
and U13224 (N_13224,N_12875,N_12868);
xnor U13225 (N_13225,N_12733,N_12764);
or U13226 (N_13226,N_12964,N_12693);
and U13227 (N_13227,N_12545,N_12998);
xor U13228 (N_13228,N_12786,N_12803);
and U13229 (N_13229,N_12763,N_12661);
nand U13230 (N_13230,N_12706,N_12850);
or U13231 (N_13231,N_12509,N_12839);
or U13232 (N_13232,N_12991,N_12591);
nor U13233 (N_13233,N_12737,N_12852);
or U13234 (N_13234,N_12815,N_12607);
nor U13235 (N_13235,N_12872,N_12931);
and U13236 (N_13236,N_12690,N_12847);
xor U13237 (N_13237,N_12887,N_12503);
nor U13238 (N_13238,N_12513,N_12674);
nor U13239 (N_13239,N_12613,N_12943);
or U13240 (N_13240,N_12946,N_12754);
or U13241 (N_13241,N_12874,N_12817);
xnor U13242 (N_13242,N_12609,N_12522);
or U13243 (N_13243,N_12597,N_12944);
or U13244 (N_13244,N_12936,N_12758);
nand U13245 (N_13245,N_12586,N_12770);
nand U13246 (N_13246,N_12906,N_12917);
nor U13247 (N_13247,N_12798,N_12510);
xnor U13248 (N_13248,N_12634,N_12843);
nor U13249 (N_13249,N_12701,N_12612);
nand U13250 (N_13250,N_12931,N_12804);
and U13251 (N_13251,N_12978,N_12563);
or U13252 (N_13252,N_12505,N_12825);
or U13253 (N_13253,N_12520,N_12674);
nand U13254 (N_13254,N_12516,N_12560);
xor U13255 (N_13255,N_12647,N_12595);
nand U13256 (N_13256,N_12911,N_12905);
xnor U13257 (N_13257,N_12524,N_12567);
or U13258 (N_13258,N_12748,N_12700);
xor U13259 (N_13259,N_12645,N_12821);
nand U13260 (N_13260,N_12587,N_12739);
or U13261 (N_13261,N_12616,N_12523);
xor U13262 (N_13262,N_12689,N_12626);
xor U13263 (N_13263,N_12809,N_12559);
and U13264 (N_13264,N_12819,N_12940);
xor U13265 (N_13265,N_12656,N_12993);
nor U13266 (N_13266,N_12918,N_12930);
xnor U13267 (N_13267,N_12629,N_12652);
nand U13268 (N_13268,N_12811,N_12601);
and U13269 (N_13269,N_12924,N_12523);
xor U13270 (N_13270,N_12559,N_12838);
xnor U13271 (N_13271,N_12900,N_12614);
nand U13272 (N_13272,N_12922,N_12540);
or U13273 (N_13273,N_12560,N_12599);
nor U13274 (N_13274,N_12610,N_12976);
xor U13275 (N_13275,N_12592,N_12594);
and U13276 (N_13276,N_12757,N_12794);
nand U13277 (N_13277,N_12883,N_12974);
nor U13278 (N_13278,N_12683,N_12553);
nand U13279 (N_13279,N_12997,N_12505);
nand U13280 (N_13280,N_12837,N_12592);
nor U13281 (N_13281,N_12898,N_12819);
nand U13282 (N_13282,N_12841,N_12549);
or U13283 (N_13283,N_12683,N_12532);
nand U13284 (N_13284,N_12555,N_12679);
or U13285 (N_13285,N_12875,N_12962);
nand U13286 (N_13286,N_12641,N_12622);
or U13287 (N_13287,N_12562,N_12948);
or U13288 (N_13288,N_12845,N_12778);
xor U13289 (N_13289,N_12537,N_12944);
xnor U13290 (N_13290,N_12662,N_12846);
nor U13291 (N_13291,N_12947,N_12789);
xor U13292 (N_13292,N_12627,N_12889);
or U13293 (N_13293,N_12651,N_12961);
and U13294 (N_13294,N_12831,N_12501);
and U13295 (N_13295,N_12573,N_12582);
nor U13296 (N_13296,N_12781,N_12538);
nand U13297 (N_13297,N_12615,N_12536);
xor U13298 (N_13298,N_12692,N_12946);
nand U13299 (N_13299,N_12715,N_12799);
nand U13300 (N_13300,N_12778,N_12575);
and U13301 (N_13301,N_12991,N_12546);
nand U13302 (N_13302,N_12783,N_12955);
or U13303 (N_13303,N_12880,N_12760);
nand U13304 (N_13304,N_12633,N_12718);
nor U13305 (N_13305,N_12567,N_12841);
nor U13306 (N_13306,N_12712,N_12864);
and U13307 (N_13307,N_12722,N_12935);
or U13308 (N_13308,N_12575,N_12968);
nor U13309 (N_13309,N_12585,N_12952);
or U13310 (N_13310,N_12679,N_12577);
and U13311 (N_13311,N_12574,N_12881);
xor U13312 (N_13312,N_12801,N_12525);
xnor U13313 (N_13313,N_12976,N_12668);
and U13314 (N_13314,N_12997,N_12739);
xnor U13315 (N_13315,N_12860,N_12760);
nand U13316 (N_13316,N_12821,N_12918);
nor U13317 (N_13317,N_12549,N_12788);
nand U13318 (N_13318,N_12675,N_12869);
xnor U13319 (N_13319,N_12859,N_12652);
or U13320 (N_13320,N_12508,N_12761);
or U13321 (N_13321,N_12567,N_12820);
nand U13322 (N_13322,N_12730,N_12867);
nand U13323 (N_13323,N_12540,N_12952);
and U13324 (N_13324,N_12764,N_12722);
xor U13325 (N_13325,N_12950,N_12549);
nor U13326 (N_13326,N_12981,N_12755);
xnor U13327 (N_13327,N_12549,N_12633);
nand U13328 (N_13328,N_12623,N_12881);
or U13329 (N_13329,N_12985,N_12980);
nor U13330 (N_13330,N_12768,N_12502);
nor U13331 (N_13331,N_12920,N_12825);
or U13332 (N_13332,N_12893,N_12569);
nand U13333 (N_13333,N_12854,N_12867);
and U13334 (N_13334,N_12645,N_12701);
xor U13335 (N_13335,N_12568,N_12593);
and U13336 (N_13336,N_12964,N_12568);
nor U13337 (N_13337,N_12994,N_12710);
xnor U13338 (N_13338,N_12909,N_12618);
or U13339 (N_13339,N_12585,N_12953);
nand U13340 (N_13340,N_12841,N_12747);
and U13341 (N_13341,N_12626,N_12516);
nand U13342 (N_13342,N_12728,N_12850);
nand U13343 (N_13343,N_12896,N_12513);
nor U13344 (N_13344,N_12857,N_12853);
and U13345 (N_13345,N_12530,N_12554);
nor U13346 (N_13346,N_12649,N_12861);
or U13347 (N_13347,N_12588,N_12581);
nor U13348 (N_13348,N_12939,N_12514);
or U13349 (N_13349,N_12525,N_12952);
nand U13350 (N_13350,N_12866,N_12819);
nor U13351 (N_13351,N_12945,N_12680);
xor U13352 (N_13352,N_12624,N_12945);
xor U13353 (N_13353,N_12540,N_12756);
xor U13354 (N_13354,N_12736,N_12878);
nand U13355 (N_13355,N_12850,N_12681);
nand U13356 (N_13356,N_12670,N_12751);
and U13357 (N_13357,N_12926,N_12987);
nor U13358 (N_13358,N_12634,N_12562);
and U13359 (N_13359,N_12728,N_12840);
nor U13360 (N_13360,N_12611,N_12638);
nand U13361 (N_13361,N_12585,N_12899);
xnor U13362 (N_13362,N_12702,N_12573);
nand U13363 (N_13363,N_12821,N_12837);
or U13364 (N_13364,N_12617,N_12934);
nor U13365 (N_13365,N_12960,N_12717);
nor U13366 (N_13366,N_12507,N_12724);
or U13367 (N_13367,N_12618,N_12517);
nor U13368 (N_13368,N_12731,N_12645);
nand U13369 (N_13369,N_12511,N_12555);
xnor U13370 (N_13370,N_12596,N_12510);
or U13371 (N_13371,N_12507,N_12510);
xnor U13372 (N_13372,N_12604,N_12695);
or U13373 (N_13373,N_12634,N_12874);
and U13374 (N_13374,N_12996,N_12760);
and U13375 (N_13375,N_12963,N_12528);
xor U13376 (N_13376,N_12701,N_12644);
and U13377 (N_13377,N_12503,N_12582);
xor U13378 (N_13378,N_12837,N_12558);
and U13379 (N_13379,N_12750,N_12914);
nand U13380 (N_13380,N_12896,N_12690);
nand U13381 (N_13381,N_12833,N_12760);
xor U13382 (N_13382,N_12907,N_12773);
and U13383 (N_13383,N_12956,N_12619);
xnor U13384 (N_13384,N_12997,N_12976);
nand U13385 (N_13385,N_12600,N_12928);
and U13386 (N_13386,N_12643,N_12507);
and U13387 (N_13387,N_12794,N_12958);
or U13388 (N_13388,N_12523,N_12658);
and U13389 (N_13389,N_12653,N_12591);
nand U13390 (N_13390,N_12800,N_12538);
or U13391 (N_13391,N_12800,N_12946);
xor U13392 (N_13392,N_12766,N_12593);
xnor U13393 (N_13393,N_12666,N_12778);
or U13394 (N_13394,N_12570,N_12880);
and U13395 (N_13395,N_12606,N_12512);
nor U13396 (N_13396,N_12636,N_12985);
or U13397 (N_13397,N_12987,N_12681);
or U13398 (N_13398,N_12592,N_12542);
nor U13399 (N_13399,N_12794,N_12701);
or U13400 (N_13400,N_12504,N_12693);
nor U13401 (N_13401,N_12609,N_12871);
and U13402 (N_13402,N_12948,N_12837);
nor U13403 (N_13403,N_12741,N_12769);
xnor U13404 (N_13404,N_12814,N_12516);
or U13405 (N_13405,N_12610,N_12885);
nand U13406 (N_13406,N_12517,N_12678);
nand U13407 (N_13407,N_12649,N_12997);
and U13408 (N_13408,N_12677,N_12853);
nand U13409 (N_13409,N_12897,N_12693);
or U13410 (N_13410,N_12714,N_12943);
nand U13411 (N_13411,N_12691,N_12603);
xnor U13412 (N_13412,N_12782,N_12891);
or U13413 (N_13413,N_12982,N_12523);
and U13414 (N_13414,N_12606,N_12761);
or U13415 (N_13415,N_12938,N_12823);
nand U13416 (N_13416,N_12852,N_12593);
xor U13417 (N_13417,N_12965,N_12686);
xor U13418 (N_13418,N_12926,N_12727);
xnor U13419 (N_13419,N_12745,N_12536);
xor U13420 (N_13420,N_12909,N_12538);
or U13421 (N_13421,N_12845,N_12769);
or U13422 (N_13422,N_12934,N_12879);
nor U13423 (N_13423,N_12795,N_12842);
xor U13424 (N_13424,N_12700,N_12786);
nor U13425 (N_13425,N_12713,N_12655);
and U13426 (N_13426,N_12896,N_12723);
or U13427 (N_13427,N_12832,N_12936);
nand U13428 (N_13428,N_12866,N_12584);
nand U13429 (N_13429,N_12907,N_12950);
or U13430 (N_13430,N_12748,N_12869);
or U13431 (N_13431,N_12749,N_12514);
and U13432 (N_13432,N_12735,N_12904);
xnor U13433 (N_13433,N_12841,N_12606);
and U13434 (N_13434,N_12833,N_12561);
xor U13435 (N_13435,N_12551,N_12837);
nor U13436 (N_13436,N_12610,N_12959);
or U13437 (N_13437,N_12570,N_12508);
nand U13438 (N_13438,N_12544,N_12677);
nor U13439 (N_13439,N_12557,N_12734);
and U13440 (N_13440,N_12892,N_12854);
or U13441 (N_13441,N_12589,N_12618);
nor U13442 (N_13442,N_12554,N_12827);
xnor U13443 (N_13443,N_12796,N_12926);
nor U13444 (N_13444,N_12565,N_12856);
nand U13445 (N_13445,N_12719,N_12835);
and U13446 (N_13446,N_12903,N_12605);
nor U13447 (N_13447,N_12997,N_12651);
xor U13448 (N_13448,N_12874,N_12826);
and U13449 (N_13449,N_12642,N_12937);
xnor U13450 (N_13450,N_12537,N_12504);
and U13451 (N_13451,N_12686,N_12937);
nor U13452 (N_13452,N_12976,N_12747);
xor U13453 (N_13453,N_12839,N_12955);
or U13454 (N_13454,N_12770,N_12937);
nor U13455 (N_13455,N_12670,N_12752);
or U13456 (N_13456,N_12913,N_12678);
nand U13457 (N_13457,N_12758,N_12832);
nand U13458 (N_13458,N_12614,N_12650);
or U13459 (N_13459,N_12957,N_12742);
nand U13460 (N_13460,N_12626,N_12770);
xnor U13461 (N_13461,N_12838,N_12542);
and U13462 (N_13462,N_12907,N_12659);
nor U13463 (N_13463,N_12794,N_12745);
nor U13464 (N_13464,N_12786,N_12562);
nand U13465 (N_13465,N_12582,N_12671);
and U13466 (N_13466,N_12543,N_12770);
or U13467 (N_13467,N_12997,N_12740);
nand U13468 (N_13468,N_12733,N_12623);
or U13469 (N_13469,N_12523,N_12713);
and U13470 (N_13470,N_12819,N_12965);
or U13471 (N_13471,N_12587,N_12862);
and U13472 (N_13472,N_12725,N_12920);
nor U13473 (N_13473,N_12649,N_12578);
or U13474 (N_13474,N_12621,N_12679);
nand U13475 (N_13475,N_12785,N_12606);
xor U13476 (N_13476,N_12945,N_12682);
and U13477 (N_13477,N_12626,N_12793);
nor U13478 (N_13478,N_12850,N_12969);
xor U13479 (N_13479,N_12929,N_12931);
or U13480 (N_13480,N_12675,N_12990);
nor U13481 (N_13481,N_12703,N_12555);
and U13482 (N_13482,N_12965,N_12723);
nor U13483 (N_13483,N_12510,N_12520);
xor U13484 (N_13484,N_12642,N_12573);
or U13485 (N_13485,N_12615,N_12898);
and U13486 (N_13486,N_12593,N_12807);
nand U13487 (N_13487,N_12634,N_12876);
nor U13488 (N_13488,N_12543,N_12687);
and U13489 (N_13489,N_12736,N_12598);
nor U13490 (N_13490,N_12724,N_12833);
nor U13491 (N_13491,N_12566,N_12987);
and U13492 (N_13492,N_12865,N_12792);
xor U13493 (N_13493,N_12858,N_12802);
and U13494 (N_13494,N_12535,N_12790);
nand U13495 (N_13495,N_12705,N_12692);
and U13496 (N_13496,N_12648,N_12742);
nand U13497 (N_13497,N_12614,N_12846);
nand U13498 (N_13498,N_12689,N_12798);
nand U13499 (N_13499,N_12602,N_12928);
and U13500 (N_13500,N_13013,N_13073);
and U13501 (N_13501,N_13192,N_13471);
xnor U13502 (N_13502,N_13110,N_13119);
and U13503 (N_13503,N_13054,N_13261);
or U13504 (N_13504,N_13216,N_13333);
and U13505 (N_13505,N_13231,N_13461);
and U13506 (N_13506,N_13227,N_13037);
nor U13507 (N_13507,N_13141,N_13277);
or U13508 (N_13508,N_13423,N_13284);
and U13509 (N_13509,N_13418,N_13036);
nand U13510 (N_13510,N_13030,N_13003);
nand U13511 (N_13511,N_13462,N_13487);
nor U13512 (N_13512,N_13228,N_13479);
and U13513 (N_13513,N_13397,N_13352);
or U13514 (N_13514,N_13497,N_13004);
and U13515 (N_13515,N_13485,N_13409);
nor U13516 (N_13516,N_13388,N_13172);
or U13517 (N_13517,N_13079,N_13304);
xnor U13518 (N_13518,N_13392,N_13134);
and U13519 (N_13519,N_13191,N_13088);
and U13520 (N_13520,N_13140,N_13345);
and U13521 (N_13521,N_13321,N_13325);
and U13522 (N_13522,N_13414,N_13308);
nand U13523 (N_13523,N_13106,N_13326);
or U13524 (N_13524,N_13449,N_13302);
and U13525 (N_13525,N_13393,N_13419);
and U13526 (N_13526,N_13052,N_13235);
nand U13527 (N_13527,N_13203,N_13437);
nand U13528 (N_13528,N_13039,N_13383);
nor U13529 (N_13529,N_13221,N_13441);
nand U13530 (N_13530,N_13456,N_13122);
nor U13531 (N_13531,N_13102,N_13319);
xor U13532 (N_13532,N_13185,N_13042);
and U13533 (N_13533,N_13044,N_13247);
nand U13534 (N_13534,N_13432,N_13226);
and U13535 (N_13535,N_13447,N_13041);
nand U13536 (N_13536,N_13468,N_13253);
or U13537 (N_13537,N_13202,N_13312);
nand U13538 (N_13538,N_13257,N_13022);
nor U13539 (N_13539,N_13223,N_13454);
and U13540 (N_13540,N_13421,N_13299);
or U13541 (N_13541,N_13293,N_13165);
nand U13542 (N_13542,N_13362,N_13180);
and U13543 (N_13543,N_13427,N_13371);
xnor U13544 (N_13544,N_13071,N_13472);
nand U13545 (N_13545,N_13217,N_13033);
xnor U13546 (N_13546,N_13107,N_13210);
nor U13547 (N_13547,N_13368,N_13194);
nor U13548 (N_13548,N_13098,N_13364);
or U13549 (N_13549,N_13114,N_13380);
nand U13550 (N_13550,N_13330,N_13096);
and U13551 (N_13551,N_13002,N_13117);
and U13552 (N_13552,N_13199,N_13459);
or U13553 (N_13553,N_13011,N_13045);
or U13554 (N_13554,N_13076,N_13327);
xnor U13555 (N_13555,N_13491,N_13336);
nor U13556 (N_13556,N_13297,N_13341);
nor U13557 (N_13557,N_13047,N_13183);
nor U13558 (N_13558,N_13328,N_13438);
xor U13559 (N_13559,N_13389,N_13422);
xor U13560 (N_13560,N_13279,N_13120);
xnor U13561 (N_13561,N_13104,N_13118);
and U13562 (N_13562,N_13271,N_13258);
nor U13563 (N_13563,N_13386,N_13281);
xnor U13564 (N_13564,N_13061,N_13094);
nand U13565 (N_13565,N_13373,N_13143);
xor U13566 (N_13566,N_13315,N_13245);
nand U13567 (N_13567,N_13081,N_13062);
nand U13568 (N_13568,N_13178,N_13264);
and U13569 (N_13569,N_13023,N_13077);
xnor U13570 (N_13570,N_13382,N_13286);
or U13571 (N_13571,N_13375,N_13402);
nor U13572 (N_13572,N_13353,N_13145);
or U13573 (N_13573,N_13085,N_13265);
xor U13574 (N_13574,N_13137,N_13478);
or U13575 (N_13575,N_13429,N_13323);
nand U13576 (N_13576,N_13316,N_13209);
nand U13577 (N_13577,N_13480,N_13473);
nor U13578 (N_13578,N_13405,N_13334);
or U13579 (N_13579,N_13310,N_13055);
nor U13580 (N_13580,N_13218,N_13057);
and U13581 (N_13581,N_13072,N_13208);
and U13582 (N_13582,N_13469,N_13492);
xor U13583 (N_13583,N_13006,N_13347);
nand U13584 (N_13584,N_13095,N_13488);
and U13585 (N_13585,N_13028,N_13354);
xnor U13586 (N_13586,N_13018,N_13394);
nor U13587 (N_13587,N_13099,N_13356);
and U13588 (N_13588,N_13266,N_13464);
and U13589 (N_13589,N_13015,N_13442);
nand U13590 (N_13590,N_13320,N_13463);
and U13591 (N_13591,N_13411,N_13474);
xnor U13592 (N_13592,N_13189,N_13433);
nor U13593 (N_13593,N_13278,N_13309);
nor U13594 (N_13594,N_13046,N_13243);
or U13595 (N_13595,N_13358,N_13395);
or U13596 (N_13596,N_13126,N_13369);
xor U13597 (N_13597,N_13313,N_13444);
or U13598 (N_13598,N_13059,N_13434);
and U13599 (N_13599,N_13273,N_13484);
nand U13600 (N_13600,N_13372,N_13108);
nor U13601 (N_13601,N_13241,N_13049);
or U13602 (N_13602,N_13187,N_13166);
or U13603 (N_13603,N_13063,N_13360);
nand U13604 (N_13604,N_13244,N_13458);
nand U13605 (N_13605,N_13056,N_13417);
or U13606 (N_13606,N_13246,N_13379);
or U13607 (N_13607,N_13340,N_13019);
nand U13608 (N_13608,N_13374,N_13387);
nor U13609 (N_13609,N_13025,N_13342);
nand U13610 (N_13610,N_13406,N_13038);
nor U13611 (N_13611,N_13142,N_13162);
or U13612 (N_13612,N_13322,N_13020);
xnor U13613 (N_13613,N_13008,N_13317);
and U13614 (N_13614,N_13470,N_13301);
nor U13615 (N_13615,N_13158,N_13343);
nor U13616 (N_13616,N_13215,N_13251);
nor U13617 (N_13617,N_13270,N_13408);
xnor U13618 (N_13618,N_13450,N_13031);
and U13619 (N_13619,N_13365,N_13069);
nor U13620 (N_13620,N_13282,N_13465);
nor U13621 (N_13621,N_13436,N_13200);
nor U13622 (N_13622,N_13176,N_13481);
nand U13623 (N_13623,N_13300,N_13186);
nor U13624 (N_13624,N_13445,N_13133);
xnor U13625 (N_13625,N_13242,N_13359);
and U13626 (N_13626,N_13448,N_13475);
and U13627 (N_13627,N_13324,N_13381);
nand U13628 (N_13628,N_13425,N_13483);
nand U13629 (N_13629,N_13080,N_13138);
xnor U13630 (N_13630,N_13151,N_13311);
xor U13631 (N_13631,N_13065,N_13439);
nor U13632 (N_13632,N_13291,N_13109);
or U13633 (N_13633,N_13066,N_13152);
xor U13634 (N_13634,N_13154,N_13136);
nand U13635 (N_13635,N_13466,N_13026);
nand U13636 (N_13636,N_13260,N_13197);
or U13637 (N_13637,N_13115,N_13225);
nor U13638 (N_13638,N_13149,N_13053);
nand U13639 (N_13639,N_13346,N_13283);
xnor U13640 (N_13640,N_13111,N_13285);
xor U13641 (N_13641,N_13263,N_13498);
nor U13642 (N_13642,N_13024,N_13074);
and U13643 (N_13643,N_13196,N_13043);
or U13644 (N_13644,N_13295,N_13084);
xor U13645 (N_13645,N_13494,N_13089);
xor U13646 (N_13646,N_13146,N_13351);
nor U13647 (N_13647,N_13174,N_13410);
xnor U13648 (N_13648,N_13105,N_13170);
xnor U13649 (N_13649,N_13355,N_13307);
or U13650 (N_13650,N_13254,N_13125);
nand U13651 (N_13651,N_13428,N_13173);
nand U13652 (N_13652,N_13400,N_13193);
nor U13653 (N_13653,N_13268,N_13378);
or U13654 (N_13654,N_13135,N_13361);
nand U13655 (N_13655,N_13112,N_13083);
or U13656 (N_13656,N_13082,N_13179);
nor U13657 (N_13657,N_13060,N_13211);
xnor U13658 (N_13658,N_13440,N_13156);
nand U13659 (N_13659,N_13467,N_13403);
nand U13660 (N_13660,N_13415,N_13452);
nor U13661 (N_13661,N_13177,N_13219);
xor U13662 (N_13662,N_13391,N_13103);
nor U13663 (N_13663,N_13222,N_13198);
and U13664 (N_13664,N_13132,N_13490);
or U13665 (N_13665,N_13250,N_13298);
nor U13666 (N_13666,N_13236,N_13384);
xor U13667 (N_13667,N_13029,N_13007);
or U13668 (N_13668,N_13234,N_13413);
nor U13669 (N_13669,N_13303,N_13276);
nand U13670 (N_13670,N_13318,N_13237);
nand U13671 (N_13671,N_13067,N_13092);
or U13672 (N_13672,N_13129,N_13460);
xor U13673 (N_13673,N_13093,N_13249);
nand U13674 (N_13674,N_13240,N_13147);
and U13675 (N_13675,N_13288,N_13139);
and U13676 (N_13676,N_13123,N_13087);
xnor U13677 (N_13677,N_13367,N_13399);
and U13678 (N_13678,N_13090,N_13314);
or U13679 (N_13679,N_13296,N_13404);
or U13680 (N_13680,N_13280,N_13167);
nand U13681 (N_13681,N_13121,N_13213);
xnor U13682 (N_13682,N_13363,N_13124);
xnor U13683 (N_13683,N_13163,N_13262);
xor U13684 (N_13684,N_13290,N_13034);
xor U13685 (N_13685,N_13493,N_13188);
nand U13686 (N_13686,N_13477,N_13339);
or U13687 (N_13687,N_13416,N_13420);
and U13688 (N_13688,N_13160,N_13032);
and U13689 (N_13689,N_13329,N_13169);
xor U13690 (N_13690,N_13269,N_13287);
or U13691 (N_13691,N_13144,N_13184);
nand U13692 (N_13692,N_13159,N_13068);
nor U13693 (N_13693,N_13349,N_13256);
xnor U13694 (N_13694,N_13274,N_13292);
nand U13695 (N_13695,N_13001,N_13086);
and U13696 (N_13696,N_13155,N_13412);
xor U13697 (N_13697,N_13267,N_13214);
xor U13698 (N_13698,N_13335,N_13206);
or U13699 (N_13699,N_13332,N_13455);
nor U13700 (N_13700,N_13426,N_13161);
or U13701 (N_13701,N_13035,N_13229);
nand U13702 (N_13702,N_13050,N_13201);
xnor U13703 (N_13703,N_13148,N_13091);
nand U13704 (N_13704,N_13113,N_13259);
xnor U13705 (N_13705,N_13331,N_13294);
nor U13706 (N_13706,N_13014,N_13012);
or U13707 (N_13707,N_13350,N_13252);
or U13708 (N_13708,N_13212,N_13130);
nor U13709 (N_13709,N_13499,N_13116);
and U13710 (N_13710,N_13128,N_13131);
xor U13711 (N_13711,N_13100,N_13064);
nand U13712 (N_13712,N_13366,N_13181);
and U13713 (N_13713,N_13027,N_13370);
nor U13714 (N_13714,N_13435,N_13058);
xor U13715 (N_13715,N_13248,N_13010);
nand U13716 (N_13716,N_13451,N_13097);
nor U13717 (N_13717,N_13476,N_13168);
or U13718 (N_13718,N_13070,N_13376);
nor U13719 (N_13719,N_13446,N_13255);
and U13720 (N_13720,N_13407,N_13443);
nor U13721 (N_13721,N_13289,N_13398);
xnor U13722 (N_13722,N_13150,N_13431);
or U13723 (N_13723,N_13239,N_13207);
xor U13724 (N_13724,N_13305,N_13338);
nand U13725 (N_13725,N_13021,N_13005);
nand U13726 (N_13726,N_13075,N_13348);
xnor U13727 (N_13727,N_13051,N_13182);
xnor U13728 (N_13728,N_13127,N_13000);
nor U13729 (N_13729,N_13171,N_13495);
nor U13730 (N_13730,N_13205,N_13175);
xnor U13731 (N_13731,N_13453,N_13486);
nand U13732 (N_13732,N_13233,N_13306);
xor U13733 (N_13733,N_13164,N_13220);
and U13734 (N_13734,N_13401,N_13048);
and U13735 (N_13735,N_13390,N_13424);
nor U13736 (N_13736,N_13230,N_13396);
and U13737 (N_13737,N_13496,N_13238);
or U13738 (N_13738,N_13357,N_13337);
and U13739 (N_13739,N_13157,N_13232);
nand U13740 (N_13740,N_13153,N_13009);
xor U13741 (N_13741,N_13344,N_13224);
xnor U13742 (N_13742,N_13101,N_13482);
and U13743 (N_13743,N_13204,N_13272);
and U13744 (N_13744,N_13195,N_13017);
or U13745 (N_13745,N_13457,N_13377);
xor U13746 (N_13746,N_13385,N_13040);
and U13747 (N_13747,N_13016,N_13430);
nand U13748 (N_13748,N_13078,N_13190);
nand U13749 (N_13749,N_13275,N_13489);
xnor U13750 (N_13750,N_13054,N_13149);
nand U13751 (N_13751,N_13352,N_13159);
and U13752 (N_13752,N_13237,N_13155);
or U13753 (N_13753,N_13411,N_13003);
nor U13754 (N_13754,N_13365,N_13029);
nand U13755 (N_13755,N_13187,N_13243);
and U13756 (N_13756,N_13498,N_13190);
nor U13757 (N_13757,N_13353,N_13014);
nand U13758 (N_13758,N_13064,N_13401);
and U13759 (N_13759,N_13013,N_13342);
xnor U13760 (N_13760,N_13007,N_13233);
nor U13761 (N_13761,N_13347,N_13285);
nand U13762 (N_13762,N_13260,N_13473);
nand U13763 (N_13763,N_13247,N_13130);
or U13764 (N_13764,N_13408,N_13054);
xor U13765 (N_13765,N_13090,N_13235);
nand U13766 (N_13766,N_13377,N_13192);
xnor U13767 (N_13767,N_13085,N_13404);
nor U13768 (N_13768,N_13054,N_13465);
nor U13769 (N_13769,N_13092,N_13296);
and U13770 (N_13770,N_13160,N_13257);
and U13771 (N_13771,N_13453,N_13246);
and U13772 (N_13772,N_13183,N_13367);
nor U13773 (N_13773,N_13219,N_13280);
or U13774 (N_13774,N_13422,N_13437);
or U13775 (N_13775,N_13321,N_13304);
or U13776 (N_13776,N_13278,N_13340);
or U13777 (N_13777,N_13174,N_13011);
or U13778 (N_13778,N_13477,N_13202);
nor U13779 (N_13779,N_13278,N_13426);
or U13780 (N_13780,N_13299,N_13482);
or U13781 (N_13781,N_13186,N_13356);
nor U13782 (N_13782,N_13136,N_13128);
or U13783 (N_13783,N_13317,N_13027);
and U13784 (N_13784,N_13162,N_13496);
nor U13785 (N_13785,N_13268,N_13223);
and U13786 (N_13786,N_13446,N_13308);
and U13787 (N_13787,N_13137,N_13232);
nor U13788 (N_13788,N_13339,N_13409);
and U13789 (N_13789,N_13336,N_13015);
nor U13790 (N_13790,N_13368,N_13350);
nor U13791 (N_13791,N_13098,N_13441);
nor U13792 (N_13792,N_13477,N_13461);
xor U13793 (N_13793,N_13315,N_13050);
nor U13794 (N_13794,N_13258,N_13314);
nand U13795 (N_13795,N_13460,N_13437);
nor U13796 (N_13796,N_13175,N_13412);
nand U13797 (N_13797,N_13429,N_13220);
or U13798 (N_13798,N_13086,N_13376);
and U13799 (N_13799,N_13482,N_13049);
nand U13800 (N_13800,N_13494,N_13130);
or U13801 (N_13801,N_13307,N_13013);
nor U13802 (N_13802,N_13178,N_13233);
or U13803 (N_13803,N_13191,N_13009);
xnor U13804 (N_13804,N_13417,N_13016);
xnor U13805 (N_13805,N_13130,N_13390);
or U13806 (N_13806,N_13144,N_13268);
nor U13807 (N_13807,N_13072,N_13327);
nand U13808 (N_13808,N_13055,N_13409);
xnor U13809 (N_13809,N_13025,N_13473);
nand U13810 (N_13810,N_13483,N_13437);
nand U13811 (N_13811,N_13197,N_13403);
nor U13812 (N_13812,N_13291,N_13474);
or U13813 (N_13813,N_13181,N_13272);
xor U13814 (N_13814,N_13260,N_13268);
nand U13815 (N_13815,N_13075,N_13252);
and U13816 (N_13816,N_13374,N_13498);
or U13817 (N_13817,N_13230,N_13357);
xnor U13818 (N_13818,N_13120,N_13012);
or U13819 (N_13819,N_13218,N_13369);
xnor U13820 (N_13820,N_13035,N_13094);
nand U13821 (N_13821,N_13049,N_13016);
or U13822 (N_13822,N_13286,N_13069);
and U13823 (N_13823,N_13251,N_13354);
xnor U13824 (N_13824,N_13230,N_13298);
xnor U13825 (N_13825,N_13310,N_13213);
nor U13826 (N_13826,N_13495,N_13223);
nor U13827 (N_13827,N_13208,N_13215);
and U13828 (N_13828,N_13024,N_13415);
xnor U13829 (N_13829,N_13432,N_13066);
nor U13830 (N_13830,N_13487,N_13326);
nand U13831 (N_13831,N_13260,N_13129);
nand U13832 (N_13832,N_13297,N_13201);
and U13833 (N_13833,N_13428,N_13008);
or U13834 (N_13834,N_13245,N_13102);
nand U13835 (N_13835,N_13242,N_13222);
nand U13836 (N_13836,N_13224,N_13252);
or U13837 (N_13837,N_13096,N_13196);
nand U13838 (N_13838,N_13044,N_13068);
nand U13839 (N_13839,N_13129,N_13184);
nand U13840 (N_13840,N_13343,N_13333);
nor U13841 (N_13841,N_13266,N_13062);
nor U13842 (N_13842,N_13346,N_13178);
or U13843 (N_13843,N_13097,N_13446);
nand U13844 (N_13844,N_13095,N_13022);
and U13845 (N_13845,N_13324,N_13426);
xor U13846 (N_13846,N_13404,N_13339);
nor U13847 (N_13847,N_13193,N_13131);
xnor U13848 (N_13848,N_13090,N_13488);
and U13849 (N_13849,N_13418,N_13106);
nor U13850 (N_13850,N_13374,N_13071);
and U13851 (N_13851,N_13073,N_13259);
nand U13852 (N_13852,N_13406,N_13129);
xnor U13853 (N_13853,N_13306,N_13098);
nor U13854 (N_13854,N_13012,N_13129);
and U13855 (N_13855,N_13157,N_13054);
xnor U13856 (N_13856,N_13488,N_13311);
or U13857 (N_13857,N_13127,N_13126);
and U13858 (N_13858,N_13148,N_13062);
nand U13859 (N_13859,N_13264,N_13099);
nand U13860 (N_13860,N_13155,N_13199);
nor U13861 (N_13861,N_13175,N_13030);
xnor U13862 (N_13862,N_13266,N_13354);
xor U13863 (N_13863,N_13005,N_13128);
nor U13864 (N_13864,N_13450,N_13161);
xor U13865 (N_13865,N_13458,N_13058);
nor U13866 (N_13866,N_13273,N_13120);
xnor U13867 (N_13867,N_13179,N_13469);
nor U13868 (N_13868,N_13355,N_13040);
xnor U13869 (N_13869,N_13332,N_13166);
or U13870 (N_13870,N_13386,N_13197);
xnor U13871 (N_13871,N_13339,N_13364);
and U13872 (N_13872,N_13217,N_13425);
nor U13873 (N_13873,N_13088,N_13256);
nand U13874 (N_13874,N_13098,N_13423);
nor U13875 (N_13875,N_13406,N_13372);
nor U13876 (N_13876,N_13146,N_13193);
nor U13877 (N_13877,N_13054,N_13235);
xnor U13878 (N_13878,N_13361,N_13056);
or U13879 (N_13879,N_13370,N_13197);
xnor U13880 (N_13880,N_13396,N_13364);
nand U13881 (N_13881,N_13385,N_13281);
xnor U13882 (N_13882,N_13273,N_13052);
or U13883 (N_13883,N_13224,N_13354);
nor U13884 (N_13884,N_13091,N_13089);
nand U13885 (N_13885,N_13316,N_13378);
or U13886 (N_13886,N_13209,N_13119);
nand U13887 (N_13887,N_13181,N_13196);
xnor U13888 (N_13888,N_13158,N_13241);
xnor U13889 (N_13889,N_13275,N_13248);
nand U13890 (N_13890,N_13098,N_13470);
or U13891 (N_13891,N_13297,N_13037);
and U13892 (N_13892,N_13468,N_13174);
or U13893 (N_13893,N_13212,N_13303);
and U13894 (N_13894,N_13061,N_13044);
nand U13895 (N_13895,N_13327,N_13154);
nor U13896 (N_13896,N_13046,N_13392);
nor U13897 (N_13897,N_13464,N_13180);
or U13898 (N_13898,N_13199,N_13307);
or U13899 (N_13899,N_13345,N_13016);
xor U13900 (N_13900,N_13251,N_13192);
or U13901 (N_13901,N_13257,N_13013);
nor U13902 (N_13902,N_13201,N_13100);
nor U13903 (N_13903,N_13134,N_13040);
or U13904 (N_13904,N_13478,N_13477);
nor U13905 (N_13905,N_13002,N_13328);
nor U13906 (N_13906,N_13180,N_13239);
nor U13907 (N_13907,N_13288,N_13326);
xnor U13908 (N_13908,N_13100,N_13016);
or U13909 (N_13909,N_13275,N_13418);
and U13910 (N_13910,N_13107,N_13383);
xnor U13911 (N_13911,N_13372,N_13362);
xor U13912 (N_13912,N_13203,N_13390);
and U13913 (N_13913,N_13363,N_13262);
nor U13914 (N_13914,N_13036,N_13498);
or U13915 (N_13915,N_13063,N_13489);
or U13916 (N_13916,N_13450,N_13010);
xor U13917 (N_13917,N_13155,N_13414);
nor U13918 (N_13918,N_13047,N_13184);
nand U13919 (N_13919,N_13025,N_13121);
xor U13920 (N_13920,N_13408,N_13330);
and U13921 (N_13921,N_13072,N_13322);
and U13922 (N_13922,N_13494,N_13284);
nor U13923 (N_13923,N_13173,N_13160);
nand U13924 (N_13924,N_13035,N_13207);
and U13925 (N_13925,N_13370,N_13312);
nor U13926 (N_13926,N_13347,N_13033);
or U13927 (N_13927,N_13178,N_13477);
xnor U13928 (N_13928,N_13454,N_13339);
or U13929 (N_13929,N_13211,N_13364);
xor U13930 (N_13930,N_13097,N_13260);
or U13931 (N_13931,N_13180,N_13156);
nor U13932 (N_13932,N_13340,N_13436);
or U13933 (N_13933,N_13267,N_13180);
nand U13934 (N_13934,N_13152,N_13219);
and U13935 (N_13935,N_13189,N_13117);
nand U13936 (N_13936,N_13381,N_13103);
nor U13937 (N_13937,N_13479,N_13075);
or U13938 (N_13938,N_13486,N_13080);
nor U13939 (N_13939,N_13422,N_13264);
xnor U13940 (N_13940,N_13170,N_13098);
and U13941 (N_13941,N_13140,N_13339);
nor U13942 (N_13942,N_13054,N_13401);
or U13943 (N_13943,N_13266,N_13438);
xor U13944 (N_13944,N_13274,N_13336);
nand U13945 (N_13945,N_13246,N_13342);
nor U13946 (N_13946,N_13064,N_13442);
and U13947 (N_13947,N_13073,N_13481);
xor U13948 (N_13948,N_13015,N_13499);
or U13949 (N_13949,N_13359,N_13393);
nand U13950 (N_13950,N_13164,N_13059);
nor U13951 (N_13951,N_13232,N_13283);
xnor U13952 (N_13952,N_13145,N_13338);
or U13953 (N_13953,N_13134,N_13058);
nor U13954 (N_13954,N_13117,N_13003);
and U13955 (N_13955,N_13042,N_13286);
xor U13956 (N_13956,N_13316,N_13139);
nor U13957 (N_13957,N_13140,N_13103);
nor U13958 (N_13958,N_13337,N_13008);
and U13959 (N_13959,N_13351,N_13184);
nand U13960 (N_13960,N_13252,N_13282);
nand U13961 (N_13961,N_13472,N_13285);
nor U13962 (N_13962,N_13474,N_13127);
nor U13963 (N_13963,N_13377,N_13188);
nor U13964 (N_13964,N_13001,N_13300);
nand U13965 (N_13965,N_13018,N_13112);
or U13966 (N_13966,N_13199,N_13439);
xnor U13967 (N_13967,N_13023,N_13052);
or U13968 (N_13968,N_13196,N_13222);
nor U13969 (N_13969,N_13214,N_13280);
xor U13970 (N_13970,N_13359,N_13415);
or U13971 (N_13971,N_13370,N_13032);
nand U13972 (N_13972,N_13098,N_13358);
nor U13973 (N_13973,N_13468,N_13372);
nand U13974 (N_13974,N_13221,N_13211);
nand U13975 (N_13975,N_13385,N_13060);
and U13976 (N_13976,N_13476,N_13023);
or U13977 (N_13977,N_13425,N_13104);
nand U13978 (N_13978,N_13324,N_13362);
xor U13979 (N_13979,N_13163,N_13420);
or U13980 (N_13980,N_13488,N_13075);
and U13981 (N_13981,N_13192,N_13284);
nand U13982 (N_13982,N_13155,N_13114);
or U13983 (N_13983,N_13217,N_13358);
nand U13984 (N_13984,N_13032,N_13124);
or U13985 (N_13985,N_13198,N_13459);
or U13986 (N_13986,N_13437,N_13458);
and U13987 (N_13987,N_13097,N_13389);
and U13988 (N_13988,N_13496,N_13294);
or U13989 (N_13989,N_13408,N_13274);
nand U13990 (N_13990,N_13430,N_13321);
and U13991 (N_13991,N_13031,N_13006);
xnor U13992 (N_13992,N_13021,N_13090);
nor U13993 (N_13993,N_13206,N_13289);
or U13994 (N_13994,N_13035,N_13183);
or U13995 (N_13995,N_13342,N_13272);
nand U13996 (N_13996,N_13101,N_13229);
nor U13997 (N_13997,N_13160,N_13190);
nand U13998 (N_13998,N_13062,N_13111);
and U13999 (N_13999,N_13461,N_13232);
nand U14000 (N_14000,N_13925,N_13619);
or U14001 (N_14001,N_13641,N_13706);
nand U14002 (N_14002,N_13874,N_13620);
nand U14003 (N_14003,N_13767,N_13687);
nand U14004 (N_14004,N_13914,N_13541);
xor U14005 (N_14005,N_13899,N_13606);
nor U14006 (N_14006,N_13944,N_13537);
nand U14007 (N_14007,N_13857,N_13754);
or U14008 (N_14008,N_13546,N_13793);
nor U14009 (N_14009,N_13600,N_13926);
nor U14010 (N_14010,N_13545,N_13552);
or U14011 (N_14011,N_13603,N_13681);
nor U14012 (N_14012,N_13562,N_13918);
or U14013 (N_14013,N_13916,N_13710);
xnor U14014 (N_14014,N_13745,N_13594);
or U14015 (N_14015,N_13882,N_13580);
nand U14016 (N_14016,N_13997,N_13883);
nand U14017 (N_14017,N_13579,N_13954);
or U14018 (N_14018,N_13516,N_13787);
nor U14019 (N_14019,N_13674,N_13842);
xnor U14020 (N_14020,N_13662,N_13604);
nand U14021 (N_14021,N_13952,N_13500);
or U14022 (N_14022,N_13707,N_13703);
or U14023 (N_14023,N_13559,N_13844);
xor U14024 (N_14024,N_13575,N_13515);
or U14025 (N_14025,N_13624,N_13752);
or U14026 (N_14026,N_13930,N_13869);
nor U14027 (N_14027,N_13790,N_13525);
or U14028 (N_14028,N_13742,N_13753);
nor U14029 (N_14029,N_13549,N_13766);
xor U14030 (N_14030,N_13659,N_13621);
nand U14031 (N_14031,N_13775,N_13556);
or U14032 (N_14032,N_13543,N_13760);
or U14033 (N_14033,N_13743,N_13596);
or U14034 (N_14034,N_13784,N_13726);
xnor U14035 (N_14035,N_13675,N_13506);
or U14036 (N_14036,N_13840,N_13599);
and U14037 (N_14037,N_13908,N_13632);
xor U14038 (N_14038,N_13833,N_13670);
and U14039 (N_14039,N_13507,N_13544);
nor U14040 (N_14040,N_13656,N_13613);
nor U14041 (N_14041,N_13848,N_13649);
xnor U14042 (N_14042,N_13705,N_13586);
or U14043 (N_14043,N_13934,N_13886);
and U14044 (N_14044,N_13845,N_13979);
xor U14045 (N_14045,N_13563,N_13984);
nor U14046 (N_14046,N_13861,N_13587);
and U14047 (N_14047,N_13936,N_13969);
nor U14048 (N_14048,N_13666,N_13947);
or U14049 (N_14049,N_13783,N_13521);
nand U14050 (N_14050,N_13737,N_13965);
xor U14051 (N_14051,N_13591,N_13985);
nor U14052 (N_14052,N_13803,N_13609);
and U14053 (N_14053,N_13709,N_13770);
and U14054 (N_14054,N_13825,N_13827);
nor U14055 (N_14055,N_13851,N_13922);
and U14056 (N_14056,N_13906,N_13815);
or U14057 (N_14057,N_13957,N_13838);
or U14058 (N_14058,N_13530,N_13650);
or U14059 (N_14059,N_13638,N_13786);
xor U14060 (N_14060,N_13729,N_13730);
and U14061 (N_14061,N_13721,N_13762);
or U14062 (N_14062,N_13514,N_13990);
or U14063 (N_14063,N_13668,N_13776);
and U14064 (N_14064,N_13807,N_13768);
nor U14065 (N_14065,N_13592,N_13777);
nor U14066 (N_14066,N_13532,N_13690);
nor U14067 (N_14067,N_13841,N_13715);
nand U14068 (N_14068,N_13505,N_13865);
xor U14069 (N_14069,N_13871,N_13856);
nand U14070 (N_14070,N_13771,N_13864);
xor U14071 (N_14071,N_13629,N_13903);
nand U14072 (N_14072,N_13757,N_13896);
nand U14073 (N_14073,N_13900,N_13878);
or U14074 (N_14074,N_13764,N_13608);
and U14075 (N_14075,N_13810,N_13567);
nand U14076 (N_14076,N_13610,N_13590);
nand U14077 (N_14077,N_13512,N_13876);
and U14078 (N_14078,N_13818,N_13716);
and U14079 (N_14079,N_13931,N_13643);
xnor U14080 (N_14080,N_13894,N_13653);
xor U14081 (N_14081,N_13607,N_13870);
or U14082 (N_14082,N_13588,N_13695);
xor U14083 (N_14083,N_13655,N_13692);
or U14084 (N_14084,N_13879,N_13704);
xor U14085 (N_14085,N_13673,N_13948);
nand U14086 (N_14086,N_13572,N_13982);
nand U14087 (N_14087,N_13582,N_13774);
and U14088 (N_14088,N_13738,N_13701);
xnor U14089 (N_14089,N_13791,N_13828);
xor U14090 (N_14090,N_13664,N_13780);
nor U14091 (N_14091,N_13699,N_13975);
or U14092 (N_14092,N_13955,N_13538);
nand U14093 (N_14093,N_13511,N_13824);
and U14094 (N_14094,N_13831,N_13678);
and U14095 (N_14095,N_13904,N_13533);
nand U14096 (N_14096,N_13785,N_13553);
and U14097 (N_14097,N_13884,N_13826);
and U14098 (N_14098,N_13712,N_13583);
xnor U14099 (N_14099,N_13688,N_13637);
xor U14100 (N_14100,N_13999,N_13855);
and U14101 (N_14101,N_13635,N_13928);
xnor U14102 (N_14102,N_13667,N_13526);
xor U14103 (N_14103,N_13685,N_13817);
nor U14104 (N_14104,N_13773,N_13593);
xnor U14105 (N_14105,N_13551,N_13581);
and U14106 (N_14106,N_13565,N_13960);
nand U14107 (N_14107,N_13866,N_13501);
or U14108 (N_14108,N_13569,N_13750);
and U14109 (N_14109,N_13973,N_13995);
nand U14110 (N_14110,N_13510,N_13809);
or U14111 (N_14111,N_13834,N_13920);
xor U14112 (N_14112,N_13779,N_13676);
and U14113 (N_14113,N_13555,N_13763);
xnor U14114 (N_14114,N_13802,N_13814);
and U14115 (N_14115,N_13746,N_13504);
xnor U14116 (N_14116,N_13679,N_13540);
nand U14117 (N_14117,N_13765,N_13626);
or U14118 (N_14118,N_13863,N_13937);
and U14119 (N_14119,N_13912,N_13816);
or U14120 (N_14120,N_13548,N_13938);
nor U14121 (N_14121,N_13539,N_13798);
or U14122 (N_14122,N_13837,N_13823);
xor U14123 (N_14123,N_13658,N_13713);
and U14124 (N_14124,N_13945,N_13911);
or U14125 (N_14125,N_13509,N_13598);
and U14126 (N_14126,N_13949,N_13782);
nand U14127 (N_14127,N_13518,N_13958);
nor U14128 (N_14128,N_13756,N_13939);
nor U14129 (N_14129,N_13860,N_13564);
xor U14130 (N_14130,N_13808,N_13634);
nand U14131 (N_14131,N_13996,N_13648);
nor U14132 (N_14132,N_13942,N_13987);
nand U14133 (N_14133,N_13797,N_13633);
nand U14134 (N_14134,N_13988,N_13835);
and U14135 (N_14135,N_13998,N_13616);
and U14136 (N_14136,N_13630,N_13571);
or U14137 (N_14137,N_13927,N_13714);
xnor U14138 (N_14138,N_13910,N_13820);
and U14139 (N_14139,N_13672,N_13953);
xnor U14140 (N_14140,N_13751,N_13811);
nor U14141 (N_14141,N_13689,N_13740);
xor U14142 (N_14142,N_13964,N_13535);
xor U14143 (N_14143,N_13519,N_13718);
nand U14144 (N_14144,N_13524,N_13962);
nand U14145 (N_14145,N_13561,N_13758);
or U14146 (N_14146,N_13566,N_13536);
or U14147 (N_14147,N_13986,N_13578);
and U14148 (N_14148,N_13966,N_13932);
xnor U14149 (N_14149,N_13614,N_13612);
nor U14150 (N_14150,N_13854,N_13890);
or U14151 (N_14151,N_13940,N_13684);
xor U14152 (N_14152,N_13829,N_13749);
nand U14153 (N_14153,N_13992,N_13605);
and U14154 (N_14154,N_13623,N_13909);
nand U14155 (N_14155,N_13800,N_13733);
or U14156 (N_14156,N_13769,N_13941);
nand U14157 (N_14157,N_13993,N_13839);
nand U14158 (N_14158,N_13636,N_13888);
xnor U14159 (N_14159,N_13795,N_13921);
and U14160 (N_14160,N_13905,N_13935);
nand U14161 (N_14161,N_13822,N_13568);
nor U14162 (N_14162,N_13924,N_13994);
nand U14163 (N_14163,N_13700,N_13875);
nand U14164 (N_14164,N_13872,N_13560);
nand U14165 (N_14165,N_13880,N_13907);
nand U14166 (N_14166,N_13723,N_13615);
nand U14167 (N_14167,N_13625,N_13852);
nor U14168 (N_14168,N_13885,N_13669);
and U14169 (N_14169,N_13528,N_13671);
nor U14170 (N_14170,N_13702,N_13686);
nor U14171 (N_14171,N_13584,N_13895);
nand U14172 (N_14172,N_13796,N_13917);
nand U14173 (N_14173,N_13933,N_13527);
nand U14174 (N_14174,N_13887,N_13739);
or U14175 (N_14175,N_13748,N_13736);
and U14176 (N_14176,N_13889,N_13628);
xnor U14177 (N_14177,N_13682,N_13963);
and U14178 (N_14178,N_13617,N_13873);
xnor U14179 (N_14179,N_13503,N_13639);
xnor U14180 (N_14180,N_13868,N_13970);
nand U14181 (N_14181,N_13574,N_13977);
nor U14182 (N_14182,N_13627,N_13741);
and U14183 (N_14183,N_13967,N_13696);
xnor U14184 (N_14184,N_13644,N_13722);
and U14185 (N_14185,N_13735,N_13859);
and U14186 (N_14186,N_13761,N_13642);
xor U14187 (N_14187,N_13812,N_13792);
nand U14188 (N_14188,N_13663,N_13806);
xor U14189 (N_14189,N_13819,N_13508);
nand U14190 (N_14190,N_13755,N_13520);
xor U14191 (N_14191,N_13747,N_13577);
and U14192 (N_14192,N_13640,N_13711);
and U14193 (N_14193,N_13956,N_13725);
nand U14194 (N_14194,N_13727,N_13959);
nor U14195 (N_14195,N_13821,N_13980);
nor U14196 (N_14196,N_13646,N_13772);
and U14197 (N_14197,N_13677,N_13651);
xor U14198 (N_14198,N_13877,N_13554);
and U14199 (N_14199,N_13622,N_13968);
nor U14200 (N_14200,N_13813,N_13846);
or U14201 (N_14201,N_13595,N_13732);
or U14202 (N_14202,N_13665,N_13972);
xor U14203 (N_14203,N_13660,N_13843);
or U14204 (N_14204,N_13794,N_13585);
nand U14205 (N_14205,N_13847,N_13717);
xnor U14206 (N_14206,N_13801,N_13778);
nor U14207 (N_14207,N_13691,N_13719);
nor U14208 (N_14208,N_13781,N_13915);
xnor U14209 (N_14209,N_13597,N_13542);
nor U14210 (N_14210,N_13759,N_13708);
or U14211 (N_14211,N_13654,N_13570);
and U14212 (N_14212,N_13943,N_13720);
nor U14213 (N_14213,N_13913,N_13576);
xnor U14214 (N_14214,N_13589,N_13680);
nor U14215 (N_14215,N_13849,N_13693);
nor U14216 (N_14216,N_13517,N_13789);
nand U14217 (N_14217,N_13694,N_13731);
nand U14218 (N_14218,N_13523,N_13862);
xnor U14219 (N_14219,N_13502,N_13631);
or U14220 (N_14220,N_13601,N_13804);
nor U14221 (N_14221,N_13573,N_13836);
xor U14222 (N_14222,N_13557,N_13901);
nand U14223 (N_14223,N_13547,N_13534);
or U14224 (N_14224,N_13919,N_13946);
nor U14225 (N_14225,N_13832,N_13799);
nor U14226 (N_14226,N_13698,N_13976);
and U14227 (N_14227,N_13558,N_13950);
and U14228 (N_14228,N_13892,N_13830);
or U14229 (N_14229,N_13513,N_13645);
and U14230 (N_14230,N_13602,N_13697);
nand U14231 (N_14231,N_13991,N_13971);
xnor U14232 (N_14232,N_13897,N_13652);
nor U14233 (N_14233,N_13983,N_13951);
xnor U14234 (N_14234,N_13657,N_13981);
xor U14235 (N_14235,N_13858,N_13902);
nand U14236 (N_14236,N_13724,N_13647);
nand U14237 (N_14237,N_13853,N_13529);
and U14238 (N_14238,N_13850,N_13978);
xnor U14239 (N_14239,N_13891,N_13923);
xor U14240 (N_14240,N_13522,N_13867);
nand U14241 (N_14241,N_13961,N_13893);
or U14242 (N_14242,N_13683,N_13661);
or U14243 (N_14243,N_13929,N_13788);
xor U14244 (N_14244,N_13881,N_13618);
xnor U14245 (N_14245,N_13805,N_13728);
nor U14246 (N_14246,N_13550,N_13734);
nand U14247 (N_14247,N_13898,N_13989);
nor U14248 (N_14248,N_13974,N_13744);
xnor U14249 (N_14249,N_13611,N_13531);
xor U14250 (N_14250,N_13635,N_13976);
nand U14251 (N_14251,N_13607,N_13843);
nor U14252 (N_14252,N_13799,N_13666);
nand U14253 (N_14253,N_13634,N_13919);
or U14254 (N_14254,N_13500,N_13939);
xor U14255 (N_14255,N_13877,N_13706);
nand U14256 (N_14256,N_13794,N_13872);
nand U14257 (N_14257,N_13566,N_13953);
nand U14258 (N_14258,N_13616,N_13976);
nand U14259 (N_14259,N_13532,N_13755);
xor U14260 (N_14260,N_13934,N_13511);
or U14261 (N_14261,N_13742,N_13938);
or U14262 (N_14262,N_13692,N_13796);
and U14263 (N_14263,N_13699,N_13859);
nor U14264 (N_14264,N_13560,N_13925);
or U14265 (N_14265,N_13733,N_13767);
nand U14266 (N_14266,N_13586,N_13673);
xnor U14267 (N_14267,N_13790,N_13787);
nor U14268 (N_14268,N_13538,N_13647);
or U14269 (N_14269,N_13916,N_13764);
nand U14270 (N_14270,N_13602,N_13722);
xnor U14271 (N_14271,N_13968,N_13678);
nor U14272 (N_14272,N_13865,N_13869);
and U14273 (N_14273,N_13609,N_13946);
and U14274 (N_14274,N_13954,N_13985);
and U14275 (N_14275,N_13876,N_13793);
xor U14276 (N_14276,N_13686,N_13760);
and U14277 (N_14277,N_13591,N_13851);
xor U14278 (N_14278,N_13527,N_13632);
nor U14279 (N_14279,N_13667,N_13700);
nor U14280 (N_14280,N_13579,N_13738);
or U14281 (N_14281,N_13541,N_13825);
nand U14282 (N_14282,N_13568,N_13757);
nor U14283 (N_14283,N_13660,N_13709);
nor U14284 (N_14284,N_13509,N_13710);
xnor U14285 (N_14285,N_13664,N_13722);
nor U14286 (N_14286,N_13529,N_13579);
xnor U14287 (N_14287,N_13830,N_13513);
xor U14288 (N_14288,N_13750,N_13936);
or U14289 (N_14289,N_13835,N_13725);
nand U14290 (N_14290,N_13731,N_13737);
nor U14291 (N_14291,N_13882,N_13577);
nand U14292 (N_14292,N_13674,N_13981);
or U14293 (N_14293,N_13847,N_13772);
or U14294 (N_14294,N_13520,N_13950);
nor U14295 (N_14295,N_13671,N_13667);
nor U14296 (N_14296,N_13774,N_13835);
and U14297 (N_14297,N_13756,N_13684);
xnor U14298 (N_14298,N_13965,N_13552);
nor U14299 (N_14299,N_13783,N_13775);
nor U14300 (N_14300,N_13579,N_13997);
and U14301 (N_14301,N_13753,N_13767);
or U14302 (N_14302,N_13633,N_13762);
or U14303 (N_14303,N_13779,N_13858);
xnor U14304 (N_14304,N_13873,N_13672);
xor U14305 (N_14305,N_13925,N_13639);
xor U14306 (N_14306,N_13986,N_13778);
xor U14307 (N_14307,N_13723,N_13692);
xor U14308 (N_14308,N_13590,N_13871);
nor U14309 (N_14309,N_13995,N_13842);
nand U14310 (N_14310,N_13515,N_13581);
xnor U14311 (N_14311,N_13915,N_13998);
xor U14312 (N_14312,N_13544,N_13564);
or U14313 (N_14313,N_13570,N_13685);
nor U14314 (N_14314,N_13725,N_13543);
and U14315 (N_14315,N_13524,N_13699);
nor U14316 (N_14316,N_13946,N_13898);
xnor U14317 (N_14317,N_13912,N_13867);
or U14318 (N_14318,N_13604,N_13784);
and U14319 (N_14319,N_13809,N_13729);
or U14320 (N_14320,N_13502,N_13632);
or U14321 (N_14321,N_13772,N_13512);
or U14322 (N_14322,N_13887,N_13857);
or U14323 (N_14323,N_13523,N_13517);
and U14324 (N_14324,N_13539,N_13748);
or U14325 (N_14325,N_13945,N_13923);
nand U14326 (N_14326,N_13684,N_13762);
or U14327 (N_14327,N_13687,N_13523);
nor U14328 (N_14328,N_13791,N_13573);
xor U14329 (N_14329,N_13543,N_13666);
or U14330 (N_14330,N_13809,N_13788);
nand U14331 (N_14331,N_13606,N_13585);
and U14332 (N_14332,N_13635,N_13820);
nor U14333 (N_14333,N_13792,N_13768);
nand U14334 (N_14334,N_13762,N_13883);
xnor U14335 (N_14335,N_13788,N_13575);
xnor U14336 (N_14336,N_13744,N_13679);
nand U14337 (N_14337,N_13699,N_13969);
nor U14338 (N_14338,N_13500,N_13978);
nor U14339 (N_14339,N_13877,N_13874);
xor U14340 (N_14340,N_13961,N_13785);
and U14341 (N_14341,N_13776,N_13746);
xor U14342 (N_14342,N_13705,N_13854);
xnor U14343 (N_14343,N_13826,N_13623);
or U14344 (N_14344,N_13907,N_13971);
nor U14345 (N_14345,N_13754,N_13732);
xor U14346 (N_14346,N_13791,N_13604);
or U14347 (N_14347,N_13931,N_13823);
nand U14348 (N_14348,N_13901,N_13694);
nor U14349 (N_14349,N_13637,N_13693);
or U14350 (N_14350,N_13747,N_13991);
nor U14351 (N_14351,N_13749,N_13800);
nor U14352 (N_14352,N_13542,N_13538);
nor U14353 (N_14353,N_13967,N_13854);
and U14354 (N_14354,N_13998,N_13948);
nand U14355 (N_14355,N_13797,N_13695);
xnor U14356 (N_14356,N_13812,N_13537);
nand U14357 (N_14357,N_13587,N_13905);
xnor U14358 (N_14358,N_13589,N_13853);
nor U14359 (N_14359,N_13691,N_13662);
xnor U14360 (N_14360,N_13639,N_13527);
xnor U14361 (N_14361,N_13714,N_13579);
nor U14362 (N_14362,N_13737,N_13626);
nor U14363 (N_14363,N_13734,N_13637);
nor U14364 (N_14364,N_13829,N_13680);
nand U14365 (N_14365,N_13889,N_13917);
xor U14366 (N_14366,N_13503,N_13567);
nand U14367 (N_14367,N_13505,N_13939);
nand U14368 (N_14368,N_13516,N_13741);
or U14369 (N_14369,N_13528,N_13706);
or U14370 (N_14370,N_13510,N_13802);
nand U14371 (N_14371,N_13563,N_13549);
xnor U14372 (N_14372,N_13921,N_13640);
nand U14373 (N_14373,N_13604,N_13900);
or U14374 (N_14374,N_13895,N_13817);
or U14375 (N_14375,N_13761,N_13612);
nand U14376 (N_14376,N_13803,N_13780);
and U14377 (N_14377,N_13603,N_13679);
and U14378 (N_14378,N_13800,N_13867);
xor U14379 (N_14379,N_13740,N_13625);
nor U14380 (N_14380,N_13991,N_13558);
xor U14381 (N_14381,N_13948,N_13960);
nand U14382 (N_14382,N_13718,N_13929);
xor U14383 (N_14383,N_13992,N_13904);
xnor U14384 (N_14384,N_13876,N_13671);
nand U14385 (N_14385,N_13662,N_13693);
nand U14386 (N_14386,N_13682,N_13505);
and U14387 (N_14387,N_13853,N_13972);
and U14388 (N_14388,N_13569,N_13787);
nor U14389 (N_14389,N_13749,N_13776);
and U14390 (N_14390,N_13644,N_13932);
or U14391 (N_14391,N_13508,N_13864);
or U14392 (N_14392,N_13698,N_13898);
nor U14393 (N_14393,N_13608,N_13910);
or U14394 (N_14394,N_13893,N_13994);
nand U14395 (N_14395,N_13636,N_13922);
and U14396 (N_14396,N_13509,N_13811);
nor U14397 (N_14397,N_13687,N_13707);
and U14398 (N_14398,N_13719,N_13657);
nor U14399 (N_14399,N_13946,N_13501);
nor U14400 (N_14400,N_13629,N_13622);
nand U14401 (N_14401,N_13591,N_13976);
xnor U14402 (N_14402,N_13663,N_13630);
and U14403 (N_14403,N_13557,N_13770);
nand U14404 (N_14404,N_13887,N_13803);
or U14405 (N_14405,N_13629,N_13511);
nand U14406 (N_14406,N_13594,N_13619);
or U14407 (N_14407,N_13972,N_13804);
and U14408 (N_14408,N_13960,N_13805);
nor U14409 (N_14409,N_13832,N_13830);
or U14410 (N_14410,N_13914,N_13515);
and U14411 (N_14411,N_13866,N_13594);
and U14412 (N_14412,N_13963,N_13721);
or U14413 (N_14413,N_13838,N_13576);
nand U14414 (N_14414,N_13991,N_13819);
and U14415 (N_14415,N_13776,N_13847);
nand U14416 (N_14416,N_13851,N_13751);
or U14417 (N_14417,N_13684,N_13693);
nand U14418 (N_14418,N_13892,N_13629);
nor U14419 (N_14419,N_13721,N_13857);
and U14420 (N_14420,N_13502,N_13920);
and U14421 (N_14421,N_13945,N_13722);
nor U14422 (N_14422,N_13609,N_13893);
xnor U14423 (N_14423,N_13924,N_13967);
nand U14424 (N_14424,N_13775,N_13916);
or U14425 (N_14425,N_13584,N_13779);
and U14426 (N_14426,N_13707,N_13512);
nor U14427 (N_14427,N_13754,N_13959);
nor U14428 (N_14428,N_13922,N_13928);
or U14429 (N_14429,N_13530,N_13525);
and U14430 (N_14430,N_13507,N_13628);
or U14431 (N_14431,N_13979,N_13636);
nand U14432 (N_14432,N_13841,N_13997);
xor U14433 (N_14433,N_13974,N_13976);
nand U14434 (N_14434,N_13883,N_13998);
nor U14435 (N_14435,N_13838,N_13923);
nand U14436 (N_14436,N_13911,N_13925);
xnor U14437 (N_14437,N_13516,N_13532);
and U14438 (N_14438,N_13670,N_13879);
and U14439 (N_14439,N_13747,N_13918);
and U14440 (N_14440,N_13928,N_13965);
xor U14441 (N_14441,N_13794,N_13840);
xor U14442 (N_14442,N_13534,N_13578);
nand U14443 (N_14443,N_13964,N_13748);
nand U14444 (N_14444,N_13517,N_13647);
xor U14445 (N_14445,N_13613,N_13501);
or U14446 (N_14446,N_13591,N_13775);
and U14447 (N_14447,N_13982,N_13806);
xor U14448 (N_14448,N_13989,N_13877);
or U14449 (N_14449,N_13810,N_13651);
xor U14450 (N_14450,N_13644,N_13624);
and U14451 (N_14451,N_13743,N_13508);
xor U14452 (N_14452,N_13843,N_13566);
nor U14453 (N_14453,N_13658,N_13502);
nor U14454 (N_14454,N_13978,N_13957);
xnor U14455 (N_14455,N_13972,N_13703);
xor U14456 (N_14456,N_13952,N_13906);
or U14457 (N_14457,N_13656,N_13851);
xnor U14458 (N_14458,N_13665,N_13868);
and U14459 (N_14459,N_13890,N_13881);
nand U14460 (N_14460,N_13788,N_13995);
nand U14461 (N_14461,N_13649,N_13901);
xor U14462 (N_14462,N_13780,N_13965);
and U14463 (N_14463,N_13714,N_13600);
nand U14464 (N_14464,N_13577,N_13677);
nand U14465 (N_14465,N_13635,N_13550);
nand U14466 (N_14466,N_13605,N_13827);
nand U14467 (N_14467,N_13506,N_13818);
nand U14468 (N_14468,N_13708,N_13922);
xor U14469 (N_14469,N_13556,N_13971);
and U14470 (N_14470,N_13849,N_13904);
xnor U14471 (N_14471,N_13638,N_13820);
nor U14472 (N_14472,N_13593,N_13761);
nand U14473 (N_14473,N_13941,N_13942);
or U14474 (N_14474,N_13925,N_13531);
or U14475 (N_14475,N_13881,N_13664);
or U14476 (N_14476,N_13982,N_13585);
nor U14477 (N_14477,N_13866,N_13654);
nor U14478 (N_14478,N_13658,N_13923);
and U14479 (N_14479,N_13563,N_13833);
nand U14480 (N_14480,N_13825,N_13886);
xnor U14481 (N_14481,N_13986,N_13548);
or U14482 (N_14482,N_13521,N_13870);
or U14483 (N_14483,N_13957,N_13557);
and U14484 (N_14484,N_13863,N_13793);
nor U14485 (N_14485,N_13560,N_13991);
xor U14486 (N_14486,N_13722,N_13652);
nor U14487 (N_14487,N_13791,N_13519);
xnor U14488 (N_14488,N_13890,N_13849);
or U14489 (N_14489,N_13864,N_13551);
xnor U14490 (N_14490,N_13947,N_13851);
or U14491 (N_14491,N_13922,N_13703);
and U14492 (N_14492,N_13601,N_13508);
nor U14493 (N_14493,N_13958,N_13974);
xnor U14494 (N_14494,N_13961,N_13971);
xnor U14495 (N_14495,N_13713,N_13770);
nor U14496 (N_14496,N_13546,N_13828);
nand U14497 (N_14497,N_13553,N_13569);
nor U14498 (N_14498,N_13505,N_13747);
or U14499 (N_14499,N_13959,N_13960);
and U14500 (N_14500,N_14092,N_14108);
and U14501 (N_14501,N_14120,N_14280);
nand U14502 (N_14502,N_14078,N_14281);
nand U14503 (N_14503,N_14005,N_14492);
nand U14504 (N_14504,N_14329,N_14252);
or U14505 (N_14505,N_14469,N_14466);
nor U14506 (N_14506,N_14449,N_14380);
xor U14507 (N_14507,N_14285,N_14230);
and U14508 (N_14508,N_14071,N_14400);
xnor U14509 (N_14509,N_14464,N_14495);
nand U14510 (N_14510,N_14003,N_14373);
nor U14511 (N_14511,N_14235,N_14127);
or U14512 (N_14512,N_14448,N_14227);
and U14513 (N_14513,N_14037,N_14497);
nor U14514 (N_14514,N_14477,N_14263);
or U14515 (N_14515,N_14017,N_14052);
and U14516 (N_14516,N_14129,N_14045);
nand U14517 (N_14517,N_14236,N_14275);
and U14518 (N_14518,N_14197,N_14441);
nand U14519 (N_14519,N_14090,N_14375);
nor U14520 (N_14520,N_14066,N_14257);
and U14521 (N_14521,N_14075,N_14204);
xnor U14522 (N_14522,N_14138,N_14216);
or U14523 (N_14523,N_14165,N_14198);
nand U14524 (N_14524,N_14151,N_14085);
nand U14525 (N_14525,N_14041,N_14385);
nand U14526 (N_14526,N_14047,N_14026);
and U14527 (N_14527,N_14083,N_14012);
and U14528 (N_14528,N_14038,N_14303);
and U14529 (N_14529,N_14308,N_14137);
nor U14530 (N_14530,N_14399,N_14314);
xnor U14531 (N_14531,N_14491,N_14018);
nor U14532 (N_14532,N_14261,N_14111);
nor U14533 (N_14533,N_14091,N_14228);
and U14534 (N_14534,N_14086,N_14374);
nand U14535 (N_14535,N_14069,N_14337);
nor U14536 (N_14536,N_14136,N_14435);
and U14537 (N_14537,N_14057,N_14175);
xnor U14538 (N_14538,N_14429,N_14110);
xor U14539 (N_14539,N_14403,N_14070);
xor U14540 (N_14540,N_14406,N_14382);
or U14541 (N_14541,N_14209,N_14033);
nor U14542 (N_14542,N_14221,N_14233);
xnor U14543 (N_14543,N_14426,N_14418);
nand U14544 (N_14544,N_14032,N_14455);
nand U14545 (N_14545,N_14055,N_14390);
or U14546 (N_14546,N_14008,N_14183);
or U14547 (N_14547,N_14482,N_14489);
xnor U14548 (N_14548,N_14443,N_14343);
nor U14549 (N_14549,N_14126,N_14474);
and U14550 (N_14550,N_14042,N_14299);
or U14551 (N_14551,N_14076,N_14162);
nand U14552 (N_14552,N_14142,N_14192);
xnor U14553 (N_14553,N_14199,N_14412);
or U14554 (N_14554,N_14481,N_14488);
or U14555 (N_14555,N_14457,N_14363);
nand U14556 (N_14556,N_14378,N_14498);
xor U14557 (N_14557,N_14413,N_14294);
xnor U14558 (N_14558,N_14254,N_14278);
or U14559 (N_14559,N_14333,N_14224);
nand U14560 (N_14560,N_14479,N_14191);
and U14561 (N_14561,N_14117,N_14348);
xor U14562 (N_14562,N_14048,N_14015);
nor U14563 (N_14563,N_14411,N_14408);
nor U14564 (N_14564,N_14011,N_14475);
or U14565 (N_14565,N_14249,N_14472);
or U14566 (N_14566,N_14270,N_14177);
nor U14567 (N_14567,N_14365,N_14058);
or U14568 (N_14568,N_14065,N_14040);
nand U14569 (N_14569,N_14319,N_14367);
nand U14570 (N_14570,N_14476,N_14148);
nand U14571 (N_14571,N_14259,N_14125);
xor U14572 (N_14572,N_14201,N_14462);
and U14573 (N_14573,N_14023,N_14007);
or U14574 (N_14574,N_14339,N_14493);
and U14575 (N_14575,N_14215,N_14107);
and U14576 (N_14576,N_14427,N_14140);
xor U14577 (N_14577,N_14437,N_14158);
nor U14578 (N_14578,N_14219,N_14445);
nor U14579 (N_14579,N_14231,N_14340);
and U14580 (N_14580,N_14346,N_14434);
and U14581 (N_14581,N_14438,N_14483);
nor U14582 (N_14582,N_14327,N_14381);
and U14583 (N_14583,N_14490,N_14321);
nand U14584 (N_14584,N_14356,N_14456);
and U14585 (N_14585,N_14415,N_14376);
xor U14586 (N_14586,N_14205,N_14453);
nor U14587 (N_14587,N_14031,N_14122);
nand U14588 (N_14588,N_14310,N_14164);
nand U14589 (N_14589,N_14282,N_14218);
and U14590 (N_14590,N_14402,N_14250);
xnor U14591 (N_14591,N_14384,N_14077);
or U14592 (N_14592,N_14487,N_14422);
and U14593 (N_14593,N_14022,N_14368);
nand U14594 (N_14594,N_14262,N_14347);
xor U14595 (N_14595,N_14392,N_14465);
or U14596 (N_14596,N_14433,N_14112);
and U14597 (N_14597,N_14034,N_14087);
nand U14598 (N_14598,N_14307,N_14121);
nand U14599 (N_14599,N_14298,N_14103);
or U14600 (N_14600,N_14362,N_14229);
xor U14601 (N_14601,N_14064,N_14234);
nand U14602 (N_14602,N_14253,N_14349);
xnor U14603 (N_14603,N_14371,N_14161);
nor U14604 (N_14604,N_14393,N_14044);
and U14605 (N_14605,N_14440,N_14116);
nand U14606 (N_14606,N_14132,N_14145);
and U14607 (N_14607,N_14217,N_14067);
xor U14608 (N_14608,N_14470,N_14207);
nor U14609 (N_14609,N_14387,N_14266);
nor U14610 (N_14610,N_14370,N_14159);
nor U14611 (N_14611,N_14154,N_14315);
and U14612 (N_14612,N_14106,N_14248);
and U14613 (N_14613,N_14289,N_14147);
and U14614 (N_14614,N_14113,N_14451);
nand U14615 (N_14615,N_14063,N_14265);
or U14616 (N_14616,N_14296,N_14369);
and U14617 (N_14617,N_14332,N_14246);
and U14618 (N_14618,N_14407,N_14267);
or U14619 (N_14619,N_14295,N_14019);
nor U14620 (N_14620,N_14398,N_14212);
nor U14621 (N_14621,N_14173,N_14225);
nor U14622 (N_14622,N_14002,N_14345);
nor U14623 (N_14623,N_14245,N_14035);
nand U14624 (N_14624,N_14021,N_14096);
and U14625 (N_14625,N_14152,N_14222);
nor U14626 (N_14626,N_14170,N_14341);
or U14627 (N_14627,N_14350,N_14318);
or U14628 (N_14628,N_14351,N_14188);
and U14629 (N_14629,N_14279,N_14214);
and U14630 (N_14630,N_14444,N_14478);
nor U14631 (N_14631,N_14238,N_14396);
nor U14632 (N_14632,N_14013,N_14068);
nand U14633 (N_14633,N_14336,N_14467);
and U14634 (N_14634,N_14088,N_14386);
nand U14635 (N_14635,N_14251,N_14283);
xnor U14636 (N_14636,N_14330,N_14352);
nor U14637 (N_14637,N_14020,N_14016);
or U14638 (N_14638,N_14424,N_14028);
nor U14639 (N_14639,N_14157,N_14050);
nand U14640 (N_14640,N_14101,N_14181);
nand U14641 (N_14641,N_14073,N_14485);
nand U14642 (N_14642,N_14202,N_14271);
xor U14643 (N_14643,N_14242,N_14049);
and U14644 (N_14644,N_14179,N_14237);
and U14645 (N_14645,N_14244,N_14043);
nand U14646 (N_14646,N_14405,N_14014);
xor U14647 (N_14647,N_14354,N_14001);
and U14648 (N_14648,N_14284,N_14496);
and U14649 (N_14649,N_14397,N_14105);
xnor U14650 (N_14650,N_14342,N_14211);
xor U14651 (N_14651,N_14160,N_14320);
xor U14652 (N_14652,N_14410,N_14141);
nand U14653 (N_14653,N_14213,N_14134);
or U14654 (N_14654,N_14059,N_14051);
nand U14655 (N_14655,N_14061,N_14499);
nand U14656 (N_14656,N_14223,N_14344);
xor U14657 (N_14657,N_14389,N_14452);
and U14658 (N_14658,N_14442,N_14184);
xor U14659 (N_14659,N_14240,N_14094);
and U14660 (N_14660,N_14287,N_14419);
and U14661 (N_14661,N_14109,N_14316);
or U14662 (N_14662,N_14080,N_14394);
or U14663 (N_14663,N_14036,N_14093);
nand U14664 (N_14664,N_14135,N_14312);
or U14665 (N_14665,N_14232,N_14072);
or U14666 (N_14666,N_14423,N_14364);
and U14667 (N_14667,N_14494,N_14430);
and U14668 (N_14668,N_14473,N_14458);
nand U14669 (N_14669,N_14186,N_14097);
or U14670 (N_14670,N_14004,N_14084);
nor U14671 (N_14671,N_14428,N_14060);
nor U14672 (N_14672,N_14391,N_14420);
and U14673 (N_14673,N_14471,N_14293);
or U14674 (N_14674,N_14178,N_14130);
nand U14675 (N_14675,N_14149,N_14190);
nor U14676 (N_14676,N_14388,N_14133);
and U14677 (N_14677,N_14404,N_14313);
xor U14678 (N_14678,N_14377,N_14432);
nand U14679 (N_14679,N_14417,N_14189);
nor U14680 (N_14680,N_14243,N_14074);
or U14681 (N_14681,N_14169,N_14409);
xnor U14682 (N_14682,N_14166,N_14255);
xnor U14683 (N_14683,N_14300,N_14025);
and U14684 (N_14684,N_14010,N_14335);
or U14685 (N_14685,N_14292,N_14029);
or U14686 (N_14686,N_14273,N_14286);
and U14687 (N_14687,N_14098,N_14102);
nand U14688 (N_14688,N_14104,N_14447);
nand U14689 (N_14689,N_14431,N_14326);
and U14690 (N_14690,N_14325,N_14171);
nor U14691 (N_14691,N_14358,N_14030);
xnor U14692 (N_14692,N_14119,N_14256);
nand U14693 (N_14693,N_14172,N_14421);
nor U14694 (N_14694,N_14174,N_14439);
nor U14695 (N_14695,N_14366,N_14009);
or U14696 (N_14696,N_14311,N_14099);
and U14697 (N_14697,N_14486,N_14291);
and U14698 (N_14698,N_14144,N_14309);
nand U14699 (N_14699,N_14276,N_14463);
nor U14700 (N_14700,N_14053,N_14446);
nor U14701 (N_14701,N_14039,N_14302);
and U14702 (N_14702,N_14206,N_14290);
and U14703 (N_14703,N_14118,N_14180);
and U14704 (N_14704,N_14247,N_14277);
nor U14705 (N_14705,N_14450,N_14131);
or U14706 (N_14706,N_14081,N_14079);
and U14707 (N_14707,N_14304,N_14383);
and U14708 (N_14708,N_14054,N_14167);
and U14709 (N_14709,N_14046,N_14460);
and U14710 (N_14710,N_14194,N_14357);
and U14711 (N_14711,N_14258,N_14226);
and U14712 (N_14712,N_14128,N_14322);
nand U14713 (N_14713,N_14195,N_14239);
nor U14714 (N_14714,N_14454,N_14461);
nand U14715 (N_14715,N_14210,N_14139);
nor U14716 (N_14716,N_14024,N_14241);
nor U14717 (N_14717,N_14089,N_14328);
nor U14718 (N_14718,N_14182,N_14395);
and U14719 (N_14719,N_14401,N_14331);
or U14720 (N_14720,N_14115,N_14459);
xor U14721 (N_14721,N_14297,N_14274);
and U14722 (N_14722,N_14155,N_14288);
or U14723 (N_14723,N_14208,N_14268);
nand U14724 (N_14724,N_14143,N_14163);
nor U14725 (N_14725,N_14379,N_14114);
or U14726 (N_14726,N_14484,N_14264);
nand U14727 (N_14727,N_14124,N_14203);
or U14728 (N_14728,N_14359,N_14334);
nor U14729 (N_14729,N_14006,N_14306);
xor U14730 (N_14730,N_14200,N_14360);
nand U14731 (N_14731,N_14416,N_14305);
or U14732 (N_14732,N_14480,N_14468);
and U14733 (N_14733,N_14027,N_14272);
xnor U14734 (N_14734,N_14260,N_14317);
or U14735 (N_14735,N_14056,N_14353);
nand U14736 (N_14736,N_14176,N_14361);
xor U14737 (N_14737,N_14000,N_14153);
or U14738 (N_14738,N_14372,N_14425);
or U14739 (N_14739,N_14414,N_14095);
xnor U14740 (N_14740,N_14146,N_14301);
and U14741 (N_14741,N_14436,N_14324);
and U14742 (N_14742,N_14355,N_14062);
nand U14743 (N_14743,N_14323,N_14123);
nor U14744 (N_14744,N_14187,N_14100);
and U14745 (N_14745,N_14082,N_14185);
xor U14746 (N_14746,N_14168,N_14269);
and U14747 (N_14747,N_14193,N_14196);
xor U14748 (N_14748,N_14220,N_14156);
or U14749 (N_14749,N_14338,N_14150);
and U14750 (N_14750,N_14258,N_14352);
nand U14751 (N_14751,N_14437,N_14371);
and U14752 (N_14752,N_14470,N_14190);
xor U14753 (N_14753,N_14055,N_14240);
xnor U14754 (N_14754,N_14151,N_14238);
nor U14755 (N_14755,N_14369,N_14039);
and U14756 (N_14756,N_14383,N_14062);
nand U14757 (N_14757,N_14390,N_14064);
xor U14758 (N_14758,N_14042,N_14151);
nor U14759 (N_14759,N_14249,N_14191);
and U14760 (N_14760,N_14048,N_14235);
nand U14761 (N_14761,N_14193,N_14135);
nand U14762 (N_14762,N_14315,N_14172);
nor U14763 (N_14763,N_14347,N_14186);
xnor U14764 (N_14764,N_14122,N_14372);
nand U14765 (N_14765,N_14091,N_14049);
nand U14766 (N_14766,N_14040,N_14245);
or U14767 (N_14767,N_14149,N_14104);
nor U14768 (N_14768,N_14035,N_14340);
or U14769 (N_14769,N_14298,N_14251);
xnor U14770 (N_14770,N_14009,N_14147);
nand U14771 (N_14771,N_14372,N_14177);
xor U14772 (N_14772,N_14313,N_14433);
nand U14773 (N_14773,N_14361,N_14321);
nand U14774 (N_14774,N_14021,N_14059);
nand U14775 (N_14775,N_14042,N_14429);
and U14776 (N_14776,N_14042,N_14442);
xnor U14777 (N_14777,N_14272,N_14331);
nand U14778 (N_14778,N_14421,N_14164);
xor U14779 (N_14779,N_14248,N_14445);
nor U14780 (N_14780,N_14354,N_14133);
nand U14781 (N_14781,N_14052,N_14396);
xnor U14782 (N_14782,N_14300,N_14303);
nor U14783 (N_14783,N_14240,N_14217);
xnor U14784 (N_14784,N_14010,N_14206);
nor U14785 (N_14785,N_14475,N_14466);
nor U14786 (N_14786,N_14415,N_14262);
and U14787 (N_14787,N_14404,N_14499);
or U14788 (N_14788,N_14061,N_14329);
nor U14789 (N_14789,N_14234,N_14238);
and U14790 (N_14790,N_14290,N_14382);
xor U14791 (N_14791,N_14400,N_14151);
and U14792 (N_14792,N_14084,N_14083);
nand U14793 (N_14793,N_14298,N_14307);
xnor U14794 (N_14794,N_14388,N_14268);
and U14795 (N_14795,N_14488,N_14277);
xnor U14796 (N_14796,N_14016,N_14004);
nor U14797 (N_14797,N_14273,N_14071);
nor U14798 (N_14798,N_14408,N_14387);
nor U14799 (N_14799,N_14437,N_14318);
nand U14800 (N_14800,N_14499,N_14168);
or U14801 (N_14801,N_14370,N_14363);
and U14802 (N_14802,N_14337,N_14081);
xor U14803 (N_14803,N_14011,N_14385);
xor U14804 (N_14804,N_14490,N_14468);
nand U14805 (N_14805,N_14414,N_14128);
nor U14806 (N_14806,N_14280,N_14134);
nand U14807 (N_14807,N_14039,N_14151);
nand U14808 (N_14808,N_14492,N_14144);
and U14809 (N_14809,N_14006,N_14370);
nor U14810 (N_14810,N_14285,N_14279);
nand U14811 (N_14811,N_14157,N_14022);
or U14812 (N_14812,N_14072,N_14318);
and U14813 (N_14813,N_14291,N_14285);
nor U14814 (N_14814,N_14285,N_14403);
nor U14815 (N_14815,N_14492,N_14133);
or U14816 (N_14816,N_14269,N_14429);
nand U14817 (N_14817,N_14170,N_14020);
nor U14818 (N_14818,N_14449,N_14403);
xnor U14819 (N_14819,N_14115,N_14085);
nor U14820 (N_14820,N_14329,N_14175);
nand U14821 (N_14821,N_14195,N_14130);
nor U14822 (N_14822,N_14367,N_14086);
and U14823 (N_14823,N_14357,N_14371);
or U14824 (N_14824,N_14337,N_14328);
xor U14825 (N_14825,N_14232,N_14261);
nand U14826 (N_14826,N_14122,N_14117);
nand U14827 (N_14827,N_14372,N_14068);
and U14828 (N_14828,N_14173,N_14288);
nand U14829 (N_14829,N_14164,N_14018);
and U14830 (N_14830,N_14044,N_14020);
xor U14831 (N_14831,N_14240,N_14210);
and U14832 (N_14832,N_14158,N_14167);
xor U14833 (N_14833,N_14137,N_14306);
nand U14834 (N_14834,N_14285,N_14396);
and U14835 (N_14835,N_14243,N_14147);
nor U14836 (N_14836,N_14175,N_14181);
nor U14837 (N_14837,N_14074,N_14400);
nor U14838 (N_14838,N_14331,N_14474);
and U14839 (N_14839,N_14001,N_14456);
and U14840 (N_14840,N_14190,N_14367);
nand U14841 (N_14841,N_14224,N_14209);
nor U14842 (N_14842,N_14135,N_14055);
and U14843 (N_14843,N_14245,N_14187);
nor U14844 (N_14844,N_14087,N_14080);
xnor U14845 (N_14845,N_14389,N_14293);
or U14846 (N_14846,N_14052,N_14310);
xor U14847 (N_14847,N_14449,N_14445);
or U14848 (N_14848,N_14184,N_14225);
xor U14849 (N_14849,N_14350,N_14338);
nand U14850 (N_14850,N_14182,N_14178);
and U14851 (N_14851,N_14406,N_14363);
nand U14852 (N_14852,N_14212,N_14497);
and U14853 (N_14853,N_14256,N_14461);
or U14854 (N_14854,N_14275,N_14041);
xnor U14855 (N_14855,N_14477,N_14319);
or U14856 (N_14856,N_14075,N_14375);
nor U14857 (N_14857,N_14347,N_14020);
or U14858 (N_14858,N_14052,N_14391);
nand U14859 (N_14859,N_14315,N_14473);
or U14860 (N_14860,N_14174,N_14064);
xor U14861 (N_14861,N_14172,N_14133);
nor U14862 (N_14862,N_14244,N_14084);
and U14863 (N_14863,N_14001,N_14068);
nand U14864 (N_14864,N_14106,N_14154);
and U14865 (N_14865,N_14109,N_14088);
xor U14866 (N_14866,N_14336,N_14127);
xnor U14867 (N_14867,N_14301,N_14361);
nand U14868 (N_14868,N_14432,N_14040);
nor U14869 (N_14869,N_14034,N_14348);
or U14870 (N_14870,N_14326,N_14120);
nor U14871 (N_14871,N_14247,N_14152);
nor U14872 (N_14872,N_14026,N_14316);
and U14873 (N_14873,N_14108,N_14247);
or U14874 (N_14874,N_14277,N_14309);
or U14875 (N_14875,N_14434,N_14047);
and U14876 (N_14876,N_14332,N_14249);
and U14877 (N_14877,N_14112,N_14103);
xor U14878 (N_14878,N_14081,N_14459);
nand U14879 (N_14879,N_14295,N_14141);
nand U14880 (N_14880,N_14472,N_14109);
or U14881 (N_14881,N_14158,N_14306);
xnor U14882 (N_14882,N_14202,N_14205);
and U14883 (N_14883,N_14411,N_14438);
and U14884 (N_14884,N_14062,N_14450);
xor U14885 (N_14885,N_14093,N_14447);
xor U14886 (N_14886,N_14407,N_14295);
xor U14887 (N_14887,N_14011,N_14412);
or U14888 (N_14888,N_14231,N_14107);
and U14889 (N_14889,N_14341,N_14366);
nor U14890 (N_14890,N_14353,N_14396);
xor U14891 (N_14891,N_14484,N_14458);
or U14892 (N_14892,N_14215,N_14253);
and U14893 (N_14893,N_14355,N_14353);
and U14894 (N_14894,N_14424,N_14238);
nand U14895 (N_14895,N_14141,N_14451);
xnor U14896 (N_14896,N_14269,N_14019);
nor U14897 (N_14897,N_14248,N_14448);
nor U14898 (N_14898,N_14459,N_14349);
xor U14899 (N_14899,N_14335,N_14448);
and U14900 (N_14900,N_14465,N_14224);
and U14901 (N_14901,N_14430,N_14401);
nor U14902 (N_14902,N_14381,N_14009);
nor U14903 (N_14903,N_14301,N_14447);
or U14904 (N_14904,N_14152,N_14345);
or U14905 (N_14905,N_14262,N_14260);
nor U14906 (N_14906,N_14313,N_14119);
xor U14907 (N_14907,N_14447,N_14266);
or U14908 (N_14908,N_14192,N_14445);
nand U14909 (N_14909,N_14281,N_14023);
xor U14910 (N_14910,N_14355,N_14270);
nand U14911 (N_14911,N_14346,N_14323);
or U14912 (N_14912,N_14375,N_14480);
and U14913 (N_14913,N_14188,N_14237);
nor U14914 (N_14914,N_14342,N_14281);
or U14915 (N_14915,N_14224,N_14204);
nor U14916 (N_14916,N_14268,N_14284);
nor U14917 (N_14917,N_14346,N_14208);
and U14918 (N_14918,N_14082,N_14419);
nand U14919 (N_14919,N_14278,N_14302);
or U14920 (N_14920,N_14191,N_14309);
and U14921 (N_14921,N_14066,N_14043);
xnor U14922 (N_14922,N_14140,N_14178);
and U14923 (N_14923,N_14004,N_14172);
nand U14924 (N_14924,N_14398,N_14303);
nand U14925 (N_14925,N_14296,N_14176);
nand U14926 (N_14926,N_14191,N_14039);
or U14927 (N_14927,N_14213,N_14420);
xnor U14928 (N_14928,N_14191,N_14437);
xnor U14929 (N_14929,N_14062,N_14448);
or U14930 (N_14930,N_14290,N_14384);
or U14931 (N_14931,N_14384,N_14005);
or U14932 (N_14932,N_14004,N_14280);
or U14933 (N_14933,N_14329,N_14020);
and U14934 (N_14934,N_14231,N_14042);
or U14935 (N_14935,N_14403,N_14326);
nor U14936 (N_14936,N_14377,N_14373);
xnor U14937 (N_14937,N_14045,N_14067);
or U14938 (N_14938,N_14418,N_14281);
nand U14939 (N_14939,N_14212,N_14325);
xor U14940 (N_14940,N_14376,N_14416);
xor U14941 (N_14941,N_14009,N_14482);
nor U14942 (N_14942,N_14119,N_14205);
and U14943 (N_14943,N_14475,N_14202);
or U14944 (N_14944,N_14275,N_14490);
nand U14945 (N_14945,N_14434,N_14404);
or U14946 (N_14946,N_14383,N_14391);
and U14947 (N_14947,N_14041,N_14047);
xor U14948 (N_14948,N_14352,N_14101);
xnor U14949 (N_14949,N_14162,N_14279);
or U14950 (N_14950,N_14283,N_14046);
xnor U14951 (N_14951,N_14346,N_14276);
and U14952 (N_14952,N_14278,N_14093);
or U14953 (N_14953,N_14387,N_14219);
nor U14954 (N_14954,N_14127,N_14358);
and U14955 (N_14955,N_14005,N_14403);
xnor U14956 (N_14956,N_14010,N_14211);
and U14957 (N_14957,N_14275,N_14005);
nand U14958 (N_14958,N_14255,N_14104);
nor U14959 (N_14959,N_14190,N_14189);
nand U14960 (N_14960,N_14461,N_14135);
xor U14961 (N_14961,N_14024,N_14162);
nand U14962 (N_14962,N_14056,N_14089);
and U14963 (N_14963,N_14432,N_14364);
xor U14964 (N_14964,N_14415,N_14486);
xor U14965 (N_14965,N_14418,N_14127);
nand U14966 (N_14966,N_14386,N_14225);
or U14967 (N_14967,N_14456,N_14076);
and U14968 (N_14968,N_14235,N_14067);
or U14969 (N_14969,N_14489,N_14041);
xor U14970 (N_14970,N_14053,N_14147);
or U14971 (N_14971,N_14102,N_14241);
or U14972 (N_14972,N_14042,N_14405);
or U14973 (N_14973,N_14389,N_14301);
nand U14974 (N_14974,N_14218,N_14068);
nor U14975 (N_14975,N_14176,N_14171);
or U14976 (N_14976,N_14361,N_14331);
and U14977 (N_14977,N_14108,N_14130);
or U14978 (N_14978,N_14376,N_14218);
nand U14979 (N_14979,N_14301,N_14476);
and U14980 (N_14980,N_14000,N_14019);
nand U14981 (N_14981,N_14015,N_14240);
nor U14982 (N_14982,N_14213,N_14250);
nand U14983 (N_14983,N_14436,N_14421);
nor U14984 (N_14984,N_14145,N_14058);
nor U14985 (N_14985,N_14025,N_14217);
nor U14986 (N_14986,N_14118,N_14427);
nand U14987 (N_14987,N_14075,N_14436);
nor U14988 (N_14988,N_14097,N_14336);
or U14989 (N_14989,N_14212,N_14492);
xnor U14990 (N_14990,N_14211,N_14180);
xnor U14991 (N_14991,N_14000,N_14295);
xor U14992 (N_14992,N_14309,N_14267);
nor U14993 (N_14993,N_14451,N_14175);
nor U14994 (N_14994,N_14302,N_14474);
or U14995 (N_14995,N_14389,N_14203);
nor U14996 (N_14996,N_14032,N_14108);
nor U14997 (N_14997,N_14418,N_14463);
or U14998 (N_14998,N_14346,N_14231);
xnor U14999 (N_14999,N_14163,N_14192);
nand UO_0 (O_0,N_14747,N_14826);
and UO_1 (O_1,N_14631,N_14982);
nor UO_2 (O_2,N_14539,N_14564);
nand UO_3 (O_3,N_14624,N_14940);
and UO_4 (O_4,N_14570,N_14941);
and UO_5 (O_5,N_14620,N_14887);
or UO_6 (O_6,N_14724,N_14851);
nor UO_7 (O_7,N_14989,N_14864);
and UO_8 (O_8,N_14918,N_14518);
nand UO_9 (O_9,N_14521,N_14931);
and UO_10 (O_10,N_14576,N_14929);
nand UO_11 (O_11,N_14902,N_14811);
or UO_12 (O_12,N_14981,N_14711);
and UO_13 (O_13,N_14571,N_14799);
nand UO_14 (O_14,N_14590,N_14823);
and UO_15 (O_15,N_14833,N_14861);
nor UO_16 (O_16,N_14978,N_14646);
nor UO_17 (O_17,N_14947,N_14731);
nor UO_18 (O_18,N_14578,N_14917);
xnor UO_19 (O_19,N_14537,N_14775);
nor UO_20 (O_20,N_14808,N_14996);
and UO_21 (O_21,N_14769,N_14938);
or UO_22 (O_22,N_14785,N_14660);
xor UO_23 (O_23,N_14639,N_14707);
nor UO_24 (O_24,N_14859,N_14547);
xnor UO_25 (O_25,N_14640,N_14950);
and UO_26 (O_26,N_14574,N_14882);
or UO_27 (O_27,N_14734,N_14780);
and UO_28 (O_28,N_14832,N_14655);
nand UO_29 (O_29,N_14802,N_14884);
nor UO_30 (O_30,N_14736,N_14999);
xor UO_31 (O_31,N_14680,N_14916);
xor UO_32 (O_32,N_14820,N_14695);
xnor UO_33 (O_33,N_14732,N_14670);
or UO_34 (O_34,N_14567,N_14636);
and UO_35 (O_35,N_14987,N_14649);
and UO_36 (O_36,N_14662,N_14761);
or UO_37 (O_37,N_14922,N_14794);
and UO_38 (O_38,N_14910,N_14566);
nand UO_39 (O_39,N_14653,N_14877);
nand UO_40 (O_40,N_14990,N_14729);
xnor UO_41 (O_41,N_14562,N_14790);
xor UO_42 (O_42,N_14921,N_14524);
or UO_43 (O_43,N_14946,N_14677);
nor UO_44 (O_44,N_14565,N_14579);
or UO_45 (O_45,N_14984,N_14657);
or UO_46 (O_46,N_14771,N_14824);
nor UO_47 (O_47,N_14621,N_14512);
nand UO_48 (O_48,N_14671,N_14821);
nor UO_49 (O_49,N_14853,N_14651);
or UO_50 (O_50,N_14750,N_14502);
nor UO_51 (O_51,N_14805,N_14791);
and UO_52 (O_52,N_14960,N_14954);
xnor UO_53 (O_53,N_14935,N_14956);
xor UO_54 (O_54,N_14842,N_14798);
and UO_55 (O_55,N_14932,N_14980);
nand UO_56 (O_56,N_14652,N_14756);
and UO_57 (O_57,N_14880,N_14903);
nor UO_58 (O_58,N_14949,N_14638);
nor UO_59 (O_59,N_14614,N_14831);
or UO_60 (O_60,N_14948,N_14597);
xor UO_61 (O_61,N_14866,N_14792);
and UO_62 (O_62,N_14992,N_14913);
and UO_63 (O_63,N_14585,N_14608);
nor UO_64 (O_64,N_14737,N_14767);
nor UO_65 (O_65,N_14899,N_14905);
or UO_66 (O_66,N_14699,N_14971);
nor UO_67 (O_67,N_14860,N_14688);
and UO_68 (O_68,N_14540,N_14745);
nand UO_69 (O_69,N_14828,N_14856);
xnor UO_70 (O_70,N_14559,N_14507);
or UO_71 (O_71,N_14985,N_14676);
and UO_72 (O_72,N_14538,N_14556);
or UO_73 (O_73,N_14613,N_14728);
nand UO_74 (O_74,N_14517,N_14598);
xor UO_75 (O_75,N_14986,N_14872);
or UO_76 (O_76,N_14925,N_14976);
nor UO_77 (O_77,N_14716,N_14901);
nor UO_78 (O_78,N_14584,N_14782);
or UO_79 (O_79,N_14604,N_14546);
xnor UO_80 (O_80,N_14587,N_14839);
nor UO_81 (O_81,N_14615,N_14519);
xnor UO_82 (O_82,N_14541,N_14898);
nor UO_83 (O_83,N_14630,N_14534);
nand UO_84 (O_84,N_14886,N_14829);
xnor UO_85 (O_85,N_14997,N_14702);
nand UO_86 (O_86,N_14983,N_14865);
and UO_87 (O_87,N_14961,N_14966);
nor UO_88 (O_88,N_14911,N_14806);
nor UO_89 (O_89,N_14606,N_14951);
and UO_90 (O_90,N_14772,N_14643);
and UO_91 (O_91,N_14625,N_14758);
or UO_92 (O_92,N_14542,N_14722);
or UO_93 (O_93,N_14689,N_14503);
nand UO_94 (O_94,N_14953,N_14658);
or UO_95 (O_95,N_14843,N_14573);
and UO_96 (O_96,N_14942,N_14786);
and UO_97 (O_97,N_14637,N_14656);
or UO_98 (O_98,N_14763,N_14675);
and UO_99 (O_99,N_14969,N_14553);
or UO_100 (O_100,N_14551,N_14970);
nand UO_101 (O_101,N_14629,N_14810);
xnor UO_102 (O_102,N_14549,N_14569);
and UO_103 (O_103,N_14719,N_14834);
or UO_104 (O_104,N_14558,N_14723);
xor UO_105 (O_105,N_14583,N_14907);
or UO_106 (O_106,N_14659,N_14908);
xor UO_107 (O_107,N_14852,N_14784);
and UO_108 (O_108,N_14513,N_14871);
xor UO_109 (O_109,N_14622,N_14754);
and UO_110 (O_110,N_14691,N_14628);
or UO_111 (O_111,N_14748,N_14881);
nand UO_112 (O_112,N_14744,N_14504);
and UO_113 (O_113,N_14550,N_14588);
xor UO_114 (O_114,N_14577,N_14878);
nand UO_115 (O_115,N_14603,N_14616);
nand UO_116 (O_116,N_14870,N_14777);
nand UO_117 (O_117,N_14706,N_14867);
xnor UO_118 (O_118,N_14891,N_14704);
or UO_119 (O_119,N_14863,N_14525);
and UO_120 (O_120,N_14514,N_14968);
or UO_121 (O_121,N_14818,N_14591);
nor UO_122 (O_122,N_14572,N_14909);
or UO_123 (O_123,N_14965,N_14869);
nand UO_124 (O_124,N_14561,N_14962);
nor UO_125 (O_125,N_14669,N_14876);
nor UO_126 (O_126,N_14885,N_14692);
and UO_127 (O_127,N_14741,N_14850);
or UO_128 (O_128,N_14581,N_14752);
xor UO_129 (O_129,N_14602,N_14623);
and UO_130 (O_130,N_14530,N_14510);
nor UO_131 (O_131,N_14520,N_14690);
or UO_132 (O_132,N_14618,N_14708);
or UO_133 (O_133,N_14827,N_14505);
or UO_134 (O_134,N_14678,N_14617);
nand UO_135 (O_135,N_14648,N_14944);
nor UO_136 (O_136,N_14845,N_14730);
nand UO_137 (O_137,N_14533,N_14720);
and UO_138 (O_138,N_14890,N_14667);
nand UO_139 (O_139,N_14789,N_14764);
nor UO_140 (O_140,N_14554,N_14595);
nand UO_141 (O_141,N_14920,N_14557);
and UO_142 (O_142,N_14847,N_14879);
nor UO_143 (O_143,N_14762,N_14645);
nor UO_144 (O_144,N_14830,N_14906);
and UO_145 (O_145,N_14757,N_14717);
xor UO_146 (O_146,N_14900,N_14500);
nand UO_147 (O_147,N_14710,N_14586);
nor UO_148 (O_148,N_14641,N_14545);
xor UO_149 (O_149,N_14964,N_14812);
and UO_150 (O_150,N_14612,N_14967);
xnor UO_151 (O_151,N_14749,N_14633);
nand UO_152 (O_152,N_14888,N_14679);
nor UO_153 (O_153,N_14816,N_14894);
nand UO_154 (O_154,N_14933,N_14753);
nor UO_155 (O_155,N_14714,N_14846);
nand UO_156 (O_156,N_14819,N_14937);
and UO_157 (O_157,N_14883,N_14698);
or UO_158 (O_158,N_14915,N_14605);
and UO_159 (O_159,N_14596,N_14822);
nor UO_160 (O_160,N_14770,N_14543);
nand UO_161 (O_161,N_14854,N_14664);
and UO_162 (O_162,N_14644,N_14560);
and UO_163 (O_163,N_14840,N_14788);
nand UO_164 (O_164,N_14727,N_14759);
nand UO_165 (O_165,N_14979,N_14774);
or UO_166 (O_166,N_14779,N_14508);
and UO_167 (O_167,N_14528,N_14607);
nand UO_168 (O_168,N_14686,N_14563);
nand UO_169 (O_169,N_14995,N_14582);
xnor UO_170 (O_170,N_14634,N_14778);
and UO_171 (O_171,N_14666,N_14661);
or UO_172 (O_172,N_14804,N_14781);
nand UO_173 (O_173,N_14793,N_14751);
xor UO_174 (O_174,N_14912,N_14536);
nand UO_175 (O_175,N_14776,N_14738);
nand UO_176 (O_176,N_14797,N_14975);
nor UO_177 (O_177,N_14814,N_14855);
and UO_178 (O_178,N_14889,N_14895);
nand UO_179 (O_179,N_14897,N_14632);
nand UO_180 (O_180,N_14681,N_14531);
or UO_181 (O_181,N_14934,N_14725);
nor UO_182 (O_182,N_14957,N_14904);
nor UO_183 (O_183,N_14974,N_14849);
and UO_184 (O_184,N_14610,N_14939);
and UO_185 (O_185,N_14930,N_14693);
nor UO_186 (O_186,N_14665,N_14836);
nand UO_187 (O_187,N_14694,N_14926);
nor UO_188 (O_188,N_14892,N_14773);
xor UO_189 (O_189,N_14787,N_14509);
and UO_190 (O_190,N_14800,N_14796);
and UO_191 (O_191,N_14589,N_14552);
and UO_192 (O_192,N_14746,N_14914);
xor UO_193 (O_193,N_14700,N_14893);
or UO_194 (O_194,N_14919,N_14715);
xnor UO_195 (O_195,N_14568,N_14735);
or UO_196 (O_196,N_14768,N_14783);
xor UO_197 (O_197,N_14532,N_14998);
or UO_198 (O_198,N_14709,N_14743);
or UO_199 (O_199,N_14873,N_14611);
or UO_200 (O_200,N_14994,N_14740);
or UO_201 (O_201,N_14801,N_14682);
and UO_202 (O_202,N_14672,N_14544);
nor UO_203 (O_203,N_14924,N_14712);
nand UO_204 (O_204,N_14627,N_14501);
and UO_205 (O_205,N_14599,N_14896);
nand UO_206 (O_206,N_14683,N_14844);
or UO_207 (O_207,N_14815,N_14642);
xnor UO_208 (O_208,N_14943,N_14526);
and UO_209 (O_209,N_14650,N_14837);
nor UO_210 (O_210,N_14857,N_14713);
xnor UO_211 (O_211,N_14817,N_14647);
nand UO_212 (O_212,N_14959,N_14663);
and UO_213 (O_213,N_14696,N_14580);
nor UO_214 (O_214,N_14874,N_14988);
xor UO_215 (O_215,N_14936,N_14765);
or UO_216 (O_216,N_14527,N_14673);
nor UO_217 (O_217,N_14594,N_14838);
xor UO_218 (O_218,N_14529,N_14795);
or UO_219 (O_219,N_14825,N_14593);
or UO_220 (O_220,N_14506,N_14626);
xnor UO_221 (O_221,N_14522,N_14755);
and UO_222 (O_222,N_14592,N_14928);
xor UO_223 (O_223,N_14760,N_14993);
nor UO_224 (O_224,N_14862,N_14697);
and UO_225 (O_225,N_14803,N_14973);
nor UO_226 (O_226,N_14548,N_14685);
nor UO_227 (O_227,N_14955,N_14958);
xnor UO_228 (O_228,N_14609,N_14963);
or UO_229 (O_229,N_14516,N_14739);
xnor UO_230 (O_230,N_14813,N_14726);
or UO_231 (O_231,N_14654,N_14945);
or UO_232 (O_232,N_14668,N_14701);
and UO_233 (O_233,N_14600,N_14923);
and UO_234 (O_234,N_14684,N_14835);
and UO_235 (O_235,N_14742,N_14635);
or UO_236 (O_236,N_14766,N_14555);
and UO_237 (O_237,N_14952,N_14848);
or UO_238 (O_238,N_14977,N_14972);
xnor UO_239 (O_239,N_14535,N_14927);
nand UO_240 (O_240,N_14601,N_14991);
nor UO_241 (O_241,N_14733,N_14705);
nand UO_242 (O_242,N_14703,N_14718);
nor UO_243 (O_243,N_14674,N_14511);
and UO_244 (O_244,N_14575,N_14807);
or UO_245 (O_245,N_14809,N_14841);
nor UO_246 (O_246,N_14721,N_14619);
xor UO_247 (O_247,N_14875,N_14687);
and UO_248 (O_248,N_14868,N_14515);
nand UO_249 (O_249,N_14523,N_14858);
xor UO_250 (O_250,N_14773,N_14763);
and UO_251 (O_251,N_14672,N_14867);
xor UO_252 (O_252,N_14941,N_14972);
and UO_253 (O_253,N_14669,N_14614);
nand UO_254 (O_254,N_14736,N_14670);
xnor UO_255 (O_255,N_14514,N_14981);
and UO_256 (O_256,N_14651,N_14922);
nor UO_257 (O_257,N_14840,N_14889);
and UO_258 (O_258,N_14727,N_14898);
or UO_259 (O_259,N_14927,N_14817);
nand UO_260 (O_260,N_14977,N_14560);
and UO_261 (O_261,N_14685,N_14954);
nor UO_262 (O_262,N_14683,N_14689);
nand UO_263 (O_263,N_14911,N_14509);
nor UO_264 (O_264,N_14752,N_14661);
nor UO_265 (O_265,N_14958,N_14804);
nor UO_266 (O_266,N_14801,N_14799);
nand UO_267 (O_267,N_14581,N_14825);
nor UO_268 (O_268,N_14738,N_14767);
or UO_269 (O_269,N_14969,N_14855);
or UO_270 (O_270,N_14745,N_14601);
nor UO_271 (O_271,N_14724,N_14571);
xor UO_272 (O_272,N_14720,N_14542);
nor UO_273 (O_273,N_14657,N_14909);
and UO_274 (O_274,N_14516,N_14685);
nor UO_275 (O_275,N_14748,N_14581);
nand UO_276 (O_276,N_14754,N_14706);
or UO_277 (O_277,N_14874,N_14699);
nor UO_278 (O_278,N_14931,N_14888);
xor UO_279 (O_279,N_14817,N_14692);
nand UO_280 (O_280,N_14544,N_14547);
and UO_281 (O_281,N_14513,N_14501);
and UO_282 (O_282,N_14586,N_14765);
and UO_283 (O_283,N_14622,N_14918);
xnor UO_284 (O_284,N_14910,N_14969);
nand UO_285 (O_285,N_14825,N_14686);
nand UO_286 (O_286,N_14985,N_14837);
xnor UO_287 (O_287,N_14541,N_14678);
and UO_288 (O_288,N_14564,N_14523);
nor UO_289 (O_289,N_14869,N_14849);
and UO_290 (O_290,N_14691,N_14843);
nor UO_291 (O_291,N_14987,N_14867);
xor UO_292 (O_292,N_14940,N_14518);
xor UO_293 (O_293,N_14941,N_14586);
nor UO_294 (O_294,N_14756,N_14679);
nor UO_295 (O_295,N_14596,N_14969);
xnor UO_296 (O_296,N_14714,N_14847);
and UO_297 (O_297,N_14759,N_14927);
nand UO_298 (O_298,N_14920,N_14922);
or UO_299 (O_299,N_14779,N_14960);
xnor UO_300 (O_300,N_14713,N_14638);
xor UO_301 (O_301,N_14656,N_14618);
or UO_302 (O_302,N_14603,N_14956);
xnor UO_303 (O_303,N_14846,N_14809);
nor UO_304 (O_304,N_14926,N_14712);
or UO_305 (O_305,N_14974,N_14741);
nand UO_306 (O_306,N_14987,N_14736);
nand UO_307 (O_307,N_14766,N_14575);
or UO_308 (O_308,N_14809,N_14676);
or UO_309 (O_309,N_14776,N_14510);
nor UO_310 (O_310,N_14640,N_14674);
nand UO_311 (O_311,N_14683,N_14750);
or UO_312 (O_312,N_14626,N_14620);
and UO_313 (O_313,N_14872,N_14998);
or UO_314 (O_314,N_14969,N_14912);
nor UO_315 (O_315,N_14572,N_14654);
nor UO_316 (O_316,N_14618,N_14823);
and UO_317 (O_317,N_14571,N_14696);
and UO_318 (O_318,N_14629,N_14664);
and UO_319 (O_319,N_14718,N_14700);
and UO_320 (O_320,N_14777,N_14703);
or UO_321 (O_321,N_14847,N_14644);
xnor UO_322 (O_322,N_14558,N_14682);
xor UO_323 (O_323,N_14632,N_14768);
nand UO_324 (O_324,N_14940,N_14936);
nand UO_325 (O_325,N_14588,N_14662);
xor UO_326 (O_326,N_14656,N_14678);
xnor UO_327 (O_327,N_14515,N_14735);
or UO_328 (O_328,N_14519,N_14528);
nand UO_329 (O_329,N_14902,N_14865);
and UO_330 (O_330,N_14620,N_14632);
and UO_331 (O_331,N_14673,N_14546);
and UO_332 (O_332,N_14646,N_14961);
and UO_333 (O_333,N_14582,N_14571);
nand UO_334 (O_334,N_14743,N_14601);
and UO_335 (O_335,N_14724,N_14731);
nor UO_336 (O_336,N_14766,N_14903);
and UO_337 (O_337,N_14991,N_14845);
nor UO_338 (O_338,N_14546,N_14736);
xnor UO_339 (O_339,N_14639,N_14901);
xnor UO_340 (O_340,N_14899,N_14982);
or UO_341 (O_341,N_14593,N_14694);
and UO_342 (O_342,N_14867,N_14692);
xnor UO_343 (O_343,N_14651,N_14799);
and UO_344 (O_344,N_14622,N_14671);
xnor UO_345 (O_345,N_14997,N_14555);
or UO_346 (O_346,N_14683,N_14558);
or UO_347 (O_347,N_14984,N_14816);
and UO_348 (O_348,N_14626,N_14921);
nor UO_349 (O_349,N_14614,N_14924);
nand UO_350 (O_350,N_14626,N_14962);
nand UO_351 (O_351,N_14813,N_14502);
or UO_352 (O_352,N_14618,N_14518);
nor UO_353 (O_353,N_14961,N_14904);
nand UO_354 (O_354,N_14955,N_14587);
xor UO_355 (O_355,N_14825,N_14534);
nand UO_356 (O_356,N_14500,N_14820);
nor UO_357 (O_357,N_14649,N_14601);
or UO_358 (O_358,N_14930,N_14542);
or UO_359 (O_359,N_14898,N_14803);
or UO_360 (O_360,N_14578,N_14742);
and UO_361 (O_361,N_14897,N_14691);
nand UO_362 (O_362,N_14709,N_14890);
nand UO_363 (O_363,N_14824,N_14865);
and UO_364 (O_364,N_14538,N_14974);
and UO_365 (O_365,N_14631,N_14686);
and UO_366 (O_366,N_14665,N_14856);
or UO_367 (O_367,N_14746,N_14753);
or UO_368 (O_368,N_14961,N_14840);
or UO_369 (O_369,N_14686,N_14649);
nand UO_370 (O_370,N_14578,N_14984);
xnor UO_371 (O_371,N_14703,N_14705);
xor UO_372 (O_372,N_14629,N_14599);
xor UO_373 (O_373,N_14700,N_14812);
nand UO_374 (O_374,N_14691,N_14518);
nor UO_375 (O_375,N_14502,N_14763);
nand UO_376 (O_376,N_14572,N_14992);
nor UO_377 (O_377,N_14816,N_14641);
nor UO_378 (O_378,N_14743,N_14971);
nand UO_379 (O_379,N_14638,N_14974);
and UO_380 (O_380,N_14991,N_14613);
or UO_381 (O_381,N_14936,N_14608);
nand UO_382 (O_382,N_14612,N_14962);
nor UO_383 (O_383,N_14684,N_14523);
nor UO_384 (O_384,N_14768,N_14822);
xor UO_385 (O_385,N_14967,N_14973);
or UO_386 (O_386,N_14886,N_14550);
nor UO_387 (O_387,N_14510,N_14761);
or UO_388 (O_388,N_14790,N_14588);
and UO_389 (O_389,N_14644,N_14746);
and UO_390 (O_390,N_14629,N_14748);
and UO_391 (O_391,N_14993,N_14633);
or UO_392 (O_392,N_14913,N_14795);
xnor UO_393 (O_393,N_14814,N_14522);
nor UO_394 (O_394,N_14631,N_14523);
and UO_395 (O_395,N_14592,N_14965);
or UO_396 (O_396,N_14658,N_14731);
or UO_397 (O_397,N_14891,N_14741);
xor UO_398 (O_398,N_14509,N_14673);
nand UO_399 (O_399,N_14928,N_14839);
or UO_400 (O_400,N_14953,N_14541);
nor UO_401 (O_401,N_14829,N_14983);
and UO_402 (O_402,N_14733,N_14679);
and UO_403 (O_403,N_14592,N_14859);
and UO_404 (O_404,N_14593,N_14826);
xor UO_405 (O_405,N_14998,N_14764);
or UO_406 (O_406,N_14831,N_14846);
nor UO_407 (O_407,N_14510,N_14746);
and UO_408 (O_408,N_14655,N_14840);
or UO_409 (O_409,N_14798,N_14575);
xnor UO_410 (O_410,N_14883,N_14548);
or UO_411 (O_411,N_14800,N_14505);
and UO_412 (O_412,N_14829,N_14814);
nor UO_413 (O_413,N_14986,N_14708);
xnor UO_414 (O_414,N_14609,N_14889);
nand UO_415 (O_415,N_14853,N_14996);
or UO_416 (O_416,N_14950,N_14599);
xnor UO_417 (O_417,N_14624,N_14647);
and UO_418 (O_418,N_14511,N_14548);
or UO_419 (O_419,N_14830,N_14741);
and UO_420 (O_420,N_14725,N_14792);
or UO_421 (O_421,N_14585,N_14554);
or UO_422 (O_422,N_14919,N_14852);
or UO_423 (O_423,N_14529,N_14700);
nand UO_424 (O_424,N_14935,N_14555);
nand UO_425 (O_425,N_14747,N_14715);
or UO_426 (O_426,N_14850,N_14966);
nand UO_427 (O_427,N_14767,N_14757);
nand UO_428 (O_428,N_14773,N_14920);
and UO_429 (O_429,N_14695,N_14670);
and UO_430 (O_430,N_14893,N_14520);
nor UO_431 (O_431,N_14771,N_14690);
or UO_432 (O_432,N_14972,N_14678);
nor UO_433 (O_433,N_14583,N_14804);
and UO_434 (O_434,N_14569,N_14672);
or UO_435 (O_435,N_14789,N_14573);
nand UO_436 (O_436,N_14972,N_14651);
xnor UO_437 (O_437,N_14942,N_14978);
and UO_438 (O_438,N_14867,N_14804);
xor UO_439 (O_439,N_14919,N_14778);
and UO_440 (O_440,N_14509,N_14777);
nand UO_441 (O_441,N_14789,N_14788);
and UO_442 (O_442,N_14657,N_14584);
or UO_443 (O_443,N_14586,N_14876);
xnor UO_444 (O_444,N_14987,N_14878);
and UO_445 (O_445,N_14597,N_14525);
nand UO_446 (O_446,N_14915,N_14730);
xor UO_447 (O_447,N_14635,N_14714);
nand UO_448 (O_448,N_14942,N_14532);
nor UO_449 (O_449,N_14655,N_14505);
and UO_450 (O_450,N_14963,N_14622);
nand UO_451 (O_451,N_14979,N_14699);
xnor UO_452 (O_452,N_14952,N_14629);
nand UO_453 (O_453,N_14598,N_14701);
and UO_454 (O_454,N_14527,N_14500);
nor UO_455 (O_455,N_14508,N_14589);
or UO_456 (O_456,N_14778,N_14557);
nor UO_457 (O_457,N_14522,N_14593);
and UO_458 (O_458,N_14628,N_14805);
nor UO_459 (O_459,N_14978,N_14962);
nor UO_460 (O_460,N_14872,N_14716);
or UO_461 (O_461,N_14855,N_14941);
xor UO_462 (O_462,N_14719,N_14827);
or UO_463 (O_463,N_14987,N_14504);
xor UO_464 (O_464,N_14919,N_14578);
xor UO_465 (O_465,N_14993,N_14968);
and UO_466 (O_466,N_14709,N_14829);
or UO_467 (O_467,N_14622,N_14953);
nor UO_468 (O_468,N_14805,N_14877);
nand UO_469 (O_469,N_14744,N_14640);
nor UO_470 (O_470,N_14816,N_14599);
nor UO_471 (O_471,N_14774,N_14673);
or UO_472 (O_472,N_14732,N_14596);
and UO_473 (O_473,N_14547,N_14796);
nor UO_474 (O_474,N_14899,N_14516);
nor UO_475 (O_475,N_14824,N_14861);
nor UO_476 (O_476,N_14620,N_14968);
nand UO_477 (O_477,N_14597,N_14979);
xnor UO_478 (O_478,N_14699,N_14789);
or UO_479 (O_479,N_14756,N_14678);
nor UO_480 (O_480,N_14736,N_14994);
or UO_481 (O_481,N_14581,N_14522);
nor UO_482 (O_482,N_14652,N_14939);
nor UO_483 (O_483,N_14927,N_14860);
or UO_484 (O_484,N_14767,N_14549);
nand UO_485 (O_485,N_14650,N_14832);
nand UO_486 (O_486,N_14939,N_14881);
and UO_487 (O_487,N_14981,N_14584);
and UO_488 (O_488,N_14901,N_14693);
xnor UO_489 (O_489,N_14647,N_14710);
nor UO_490 (O_490,N_14824,N_14960);
xor UO_491 (O_491,N_14632,N_14521);
or UO_492 (O_492,N_14895,N_14690);
xor UO_493 (O_493,N_14922,N_14749);
nand UO_494 (O_494,N_14575,N_14806);
and UO_495 (O_495,N_14551,N_14749);
nand UO_496 (O_496,N_14762,N_14872);
and UO_497 (O_497,N_14655,N_14924);
and UO_498 (O_498,N_14619,N_14894);
and UO_499 (O_499,N_14610,N_14722);
nand UO_500 (O_500,N_14883,N_14745);
nand UO_501 (O_501,N_14705,N_14744);
and UO_502 (O_502,N_14725,N_14745);
or UO_503 (O_503,N_14546,N_14818);
nand UO_504 (O_504,N_14966,N_14858);
nor UO_505 (O_505,N_14676,N_14599);
and UO_506 (O_506,N_14834,N_14648);
xnor UO_507 (O_507,N_14512,N_14931);
xor UO_508 (O_508,N_14652,N_14826);
xnor UO_509 (O_509,N_14908,N_14504);
nand UO_510 (O_510,N_14756,N_14625);
nand UO_511 (O_511,N_14700,N_14907);
and UO_512 (O_512,N_14524,N_14545);
nand UO_513 (O_513,N_14589,N_14726);
xor UO_514 (O_514,N_14535,N_14529);
nand UO_515 (O_515,N_14661,N_14941);
xor UO_516 (O_516,N_14588,N_14545);
or UO_517 (O_517,N_14885,N_14816);
nor UO_518 (O_518,N_14950,N_14834);
nand UO_519 (O_519,N_14752,N_14672);
or UO_520 (O_520,N_14970,N_14871);
xnor UO_521 (O_521,N_14938,N_14981);
xnor UO_522 (O_522,N_14513,N_14884);
xor UO_523 (O_523,N_14811,N_14932);
nor UO_524 (O_524,N_14793,N_14763);
nand UO_525 (O_525,N_14778,N_14510);
and UO_526 (O_526,N_14502,N_14666);
and UO_527 (O_527,N_14859,N_14901);
or UO_528 (O_528,N_14756,N_14570);
nor UO_529 (O_529,N_14802,N_14711);
and UO_530 (O_530,N_14814,N_14590);
nand UO_531 (O_531,N_14777,N_14563);
nand UO_532 (O_532,N_14816,N_14980);
nor UO_533 (O_533,N_14595,N_14544);
nand UO_534 (O_534,N_14827,N_14924);
nor UO_535 (O_535,N_14731,N_14763);
xnor UO_536 (O_536,N_14594,N_14931);
nand UO_537 (O_537,N_14993,N_14782);
nor UO_538 (O_538,N_14562,N_14612);
xnor UO_539 (O_539,N_14924,N_14553);
xnor UO_540 (O_540,N_14628,N_14853);
xor UO_541 (O_541,N_14794,N_14702);
nand UO_542 (O_542,N_14726,N_14709);
and UO_543 (O_543,N_14737,N_14902);
and UO_544 (O_544,N_14913,N_14841);
xnor UO_545 (O_545,N_14934,N_14824);
and UO_546 (O_546,N_14652,N_14616);
or UO_547 (O_547,N_14558,N_14892);
or UO_548 (O_548,N_14585,N_14654);
nand UO_549 (O_549,N_14921,N_14713);
nor UO_550 (O_550,N_14868,N_14524);
nand UO_551 (O_551,N_14904,N_14978);
xnor UO_552 (O_552,N_14772,N_14892);
and UO_553 (O_553,N_14829,N_14555);
nand UO_554 (O_554,N_14773,N_14754);
nand UO_555 (O_555,N_14966,N_14628);
nor UO_556 (O_556,N_14866,N_14934);
and UO_557 (O_557,N_14870,N_14892);
nor UO_558 (O_558,N_14676,N_14548);
nor UO_559 (O_559,N_14870,N_14941);
or UO_560 (O_560,N_14924,N_14564);
nor UO_561 (O_561,N_14842,N_14919);
and UO_562 (O_562,N_14534,N_14996);
and UO_563 (O_563,N_14723,N_14947);
xor UO_564 (O_564,N_14773,N_14847);
nand UO_565 (O_565,N_14504,N_14500);
xor UO_566 (O_566,N_14798,N_14502);
xor UO_567 (O_567,N_14627,N_14567);
nor UO_568 (O_568,N_14683,N_14705);
and UO_569 (O_569,N_14869,N_14862);
and UO_570 (O_570,N_14747,N_14550);
nand UO_571 (O_571,N_14864,N_14687);
or UO_572 (O_572,N_14815,N_14774);
and UO_573 (O_573,N_14898,N_14874);
nand UO_574 (O_574,N_14844,N_14573);
or UO_575 (O_575,N_14574,N_14682);
and UO_576 (O_576,N_14748,N_14513);
and UO_577 (O_577,N_14793,N_14783);
nand UO_578 (O_578,N_14693,N_14922);
and UO_579 (O_579,N_14500,N_14526);
or UO_580 (O_580,N_14971,N_14992);
nor UO_581 (O_581,N_14950,N_14916);
nand UO_582 (O_582,N_14758,N_14668);
or UO_583 (O_583,N_14868,N_14946);
nor UO_584 (O_584,N_14528,N_14931);
xor UO_585 (O_585,N_14967,N_14894);
or UO_586 (O_586,N_14527,N_14773);
and UO_587 (O_587,N_14894,N_14805);
or UO_588 (O_588,N_14688,N_14633);
xor UO_589 (O_589,N_14536,N_14784);
or UO_590 (O_590,N_14565,N_14557);
nor UO_591 (O_591,N_14730,N_14581);
nand UO_592 (O_592,N_14531,N_14702);
and UO_593 (O_593,N_14796,N_14911);
and UO_594 (O_594,N_14503,N_14554);
nor UO_595 (O_595,N_14778,N_14843);
or UO_596 (O_596,N_14557,N_14891);
xor UO_597 (O_597,N_14810,N_14500);
xnor UO_598 (O_598,N_14735,N_14891);
xnor UO_599 (O_599,N_14654,N_14662);
xor UO_600 (O_600,N_14720,N_14925);
nor UO_601 (O_601,N_14507,N_14789);
xor UO_602 (O_602,N_14827,N_14969);
and UO_603 (O_603,N_14985,N_14987);
xor UO_604 (O_604,N_14667,N_14724);
and UO_605 (O_605,N_14605,N_14694);
or UO_606 (O_606,N_14744,N_14571);
nand UO_607 (O_607,N_14904,N_14768);
nand UO_608 (O_608,N_14622,N_14799);
and UO_609 (O_609,N_14874,N_14633);
or UO_610 (O_610,N_14872,N_14880);
nor UO_611 (O_611,N_14697,N_14892);
xor UO_612 (O_612,N_14769,N_14978);
or UO_613 (O_613,N_14659,N_14962);
and UO_614 (O_614,N_14987,N_14881);
xor UO_615 (O_615,N_14504,N_14923);
nand UO_616 (O_616,N_14977,N_14646);
or UO_617 (O_617,N_14553,N_14560);
xnor UO_618 (O_618,N_14589,N_14867);
or UO_619 (O_619,N_14996,N_14856);
nor UO_620 (O_620,N_14967,N_14712);
or UO_621 (O_621,N_14537,N_14751);
and UO_622 (O_622,N_14940,N_14629);
and UO_623 (O_623,N_14901,N_14705);
or UO_624 (O_624,N_14852,N_14921);
and UO_625 (O_625,N_14559,N_14590);
xnor UO_626 (O_626,N_14882,N_14595);
or UO_627 (O_627,N_14646,N_14925);
or UO_628 (O_628,N_14655,N_14856);
and UO_629 (O_629,N_14768,N_14635);
nand UO_630 (O_630,N_14606,N_14962);
xor UO_631 (O_631,N_14585,N_14790);
nand UO_632 (O_632,N_14569,N_14757);
nor UO_633 (O_633,N_14712,N_14598);
or UO_634 (O_634,N_14666,N_14804);
or UO_635 (O_635,N_14879,N_14751);
or UO_636 (O_636,N_14560,N_14801);
xor UO_637 (O_637,N_14763,N_14609);
xnor UO_638 (O_638,N_14647,N_14941);
and UO_639 (O_639,N_14721,N_14837);
and UO_640 (O_640,N_14579,N_14538);
or UO_641 (O_641,N_14512,N_14949);
nor UO_642 (O_642,N_14545,N_14748);
and UO_643 (O_643,N_14820,N_14674);
and UO_644 (O_644,N_14927,N_14763);
nand UO_645 (O_645,N_14951,N_14748);
nor UO_646 (O_646,N_14641,N_14833);
xnor UO_647 (O_647,N_14808,N_14605);
nand UO_648 (O_648,N_14656,N_14747);
nor UO_649 (O_649,N_14972,N_14859);
xor UO_650 (O_650,N_14932,N_14797);
xor UO_651 (O_651,N_14837,N_14501);
or UO_652 (O_652,N_14839,N_14599);
nor UO_653 (O_653,N_14581,N_14766);
nand UO_654 (O_654,N_14637,N_14576);
or UO_655 (O_655,N_14515,N_14933);
nor UO_656 (O_656,N_14766,N_14865);
or UO_657 (O_657,N_14733,N_14678);
nor UO_658 (O_658,N_14727,N_14805);
and UO_659 (O_659,N_14714,N_14699);
nor UO_660 (O_660,N_14632,N_14654);
nor UO_661 (O_661,N_14564,N_14518);
and UO_662 (O_662,N_14768,N_14603);
nor UO_663 (O_663,N_14968,N_14609);
xor UO_664 (O_664,N_14650,N_14857);
nor UO_665 (O_665,N_14641,N_14910);
or UO_666 (O_666,N_14919,N_14872);
nor UO_667 (O_667,N_14804,N_14635);
and UO_668 (O_668,N_14500,N_14958);
or UO_669 (O_669,N_14638,N_14642);
and UO_670 (O_670,N_14843,N_14859);
nor UO_671 (O_671,N_14800,N_14929);
nand UO_672 (O_672,N_14713,N_14841);
nor UO_673 (O_673,N_14796,N_14745);
nand UO_674 (O_674,N_14630,N_14776);
xor UO_675 (O_675,N_14954,N_14665);
or UO_676 (O_676,N_14907,N_14932);
xnor UO_677 (O_677,N_14600,N_14766);
nand UO_678 (O_678,N_14822,N_14626);
xnor UO_679 (O_679,N_14710,N_14768);
nand UO_680 (O_680,N_14537,N_14824);
and UO_681 (O_681,N_14790,N_14633);
and UO_682 (O_682,N_14865,N_14617);
or UO_683 (O_683,N_14828,N_14875);
xor UO_684 (O_684,N_14621,N_14898);
nor UO_685 (O_685,N_14798,N_14649);
or UO_686 (O_686,N_14600,N_14750);
nor UO_687 (O_687,N_14783,N_14830);
xnor UO_688 (O_688,N_14913,N_14685);
nand UO_689 (O_689,N_14598,N_14511);
xnor UO_690 (O_690,N_14973,N_14623);
nor UO_691 (O_691,N_14605,N_14700);
nor UO_692 (O_692,N_14528,N_14705);
and UO_693 (O_693,N_14834,N_14758);
or UO_694 (O_694,N_14610,N_14832);
nor UO_695 (O_695,N_14861,N_14920);
nand UO_696 (O_696,N_14570,N_14751);
and UO_697 (O_697,N_14888,N_14504);
or UO_698 (O_698,N_14883,N_14987);
or UO_699 (O_699,N_14695,N_14594);
or UO_700 (O_700,N_14672,N_14649);
and UO_701 (O_701,N_14630,N_14869);
nand UO_702 (O_702,N_14813,N_14943);
xor UO_703 (O_703,N_14689,N_14637);
and UO_704 (O_704,N_14729,N_14773);
nor UO_705 (O_705,N_14647,N_14503);
nor UO_706 (O_706,N_14757,N_14999);
nor UO_707 (O_707,N_14792,N_14526);
nand UO_708 (O_708,N_14629,N_14930);
and UO_709 (O_709,N_14936,N_14848);
or UO_710 (O_710,N_14917,N_14672);
nand UO_711 (O_711,N_14994,N_14617);
or UO_712 (O_712,N_14732,N_14504);
nor UO_713 (O_713,N_14657,N_14986);
and UO_714 (O_714,N_14973,N_14838);
nor UO_715 (O_715,N_14721,N_14930);
xnor UO_716 (O_716,N_14939,N_14523);
and UO_717 (O_717,N_14828,N_14841);
xnor UO_718 (O_718,N_14924,N_14539);
and UO_719 (O_719,N_14606,N_14657);
xnor UO_720 (O_720,N_14903,N_14698);
xnor UO_721 (O_721,N_14521,N_14872);
or UO_722 (O_722,N_14520,N_14598);
or UO_723 (O_723,N_14824,N_14850);
and UO_724 (O_724,N_14921,N_14623);
nand UO_725 (O_725,N_14899,N_14936);
nand UO_726 (O_726,N_14593,N_14838);
and UO_727 (O_727,N_14762,N_14787);
and UO_728 (O_728,N_14622,N_14657);
nor UO_729 (O_729,N_14721,N_14525);
or UO_730 (O_730,N_14854,N_14798);
nand UO_731 (O_731,N_14998,N_14706);
nand UO_732 (O_732,N_14955,N_14548);
and UO_733 (O_733,N_14828,N_14866);
or UO_734 (O_734,N_14765,N_14887);
and UO_735 (O_735,N_14646,N_14850);
nand UO_736 (O_736,N_14906,N_14916);
or UO_737 (O_737,N_14580,N_14720);
nand UO_738 (O_738,N_14783,N_14671);
nor UO_739 (O_739,N_14973,N_14752);
nor UO_740 (O_740,N_14983,N_14620);
nand UO_741 (O_741,N_14891,N_14626);
or UO_742 (O_742,N_14589,N_14523);
nand UO_743 (O_743,N_14687,N_14668);
nor UO_744 (O_744,N_14546,N_14566);
nand UO_745 (O_745,N_14671,N_14990);
nor UO_746 (O_746,N_14945,N_14789);
or UO_747 (O_747,N_14727,N_14624);
or UO_748 (O_748,N_14508,N_14720);
or UO_749 (O_749,N_14920,N_14814);
xor UO_750 (O_750,N_14825,N_14971);
and UO_751 (O_751,N_14848,N_14512);
or UO_752 (O_752,N_14582,N_14627);
nor UO_753 (O_753,N_14864,N_14833);
nor UO_754 (O_754,N_14850,N_14829);
or UO_755 (O_755,N_14709,N_14620);
or UO_756 (O_756,N_14561,N_14862);
xor UO_757 (O_757,N_14974,N_14960);
xnor UO_758 (O_758,N_14565,N_14684);
xor UO_759 (O_759,N_14542,N_14589);
nor UO_760 (O_760,N_14709,N_14634);
nand UO_761 (O_761,N_14749,N_14523);
nand UO_762 (O_762,N_14877,N_14913);
and UO_763 (O_763,N_14684,N_14783);
or UO_764 (O_764,N_14622,N_14555);
or UO_765 (O_765,N_14835,N_14512);
xor UO_766 (O_766,N_14963,N_14852);
xnor UO_767 (O_767,N_14640,N_14835);
nand UO_768 (O_768,N_14878,N_14934);
and UO_769 (O_769,N_14578,N_14545);
xor UO_770 (O_770,N_14592,N_14612);
and UO_771 (O_771,N_14838,N_14891);
xor UO_772 (O_772,N_14506,N_14525);
or UO_773 (O_773,N_14528,N_14865);
nand UO_774 (O_774,N_14849,N_14939);
and UO_775 (O_775,N_14609,N_14715);
nand UO_776 (O_776,N_14869,N_14973);
and UO_777 (O_777,N_14798,N_14937);
xnor UO_778 (O_778,N_14907,N_14546);
nand UO_779 (O_779,N_14948,N_14879);
and UO_780 (O_780,N_14629,N_14958);
nand UO_781 (O_781,N_14985,N_14558);
xor UO_782 (O_782,N_14874,N_14544);
or UO_783 (O_783,N_14889,N_14564);
and UO_784 (O_784,N_14873,N_14661);
or UO_785 (O_785,N_14561,N_14868);
and UO_786 (O_786,N_14970,N_14797);
or UO_787 (O_787,N_14876,N_14521);
nor UO_788 (O_788,N_14618,N_14950);
xor UO_789 (O_789,N_14735,N_14812);
nand UO_790 (O_790,N_14845,N_14655);
and UO_791 (O_791,N_14724,N_14585);
or UO_792 (O_792,N_14510,N_14894);
nand UO_793 (O_793,N_14757,N_14894);
nand UO_794 (O_794,N_14863,N_14991);
xnor UO_795 (O_795,N_14626,N_14849);
xor UO_796 (O_796,N_14808,N_14784);
and UO_797 (O_797,N_14653,N_14801);
nand UO_798 (O_798,N_14780,N_14504);
xnor UO_799 (O_799,N_14628,N_14857);
xor UO_800 (O_800,N_14554,N_14828);
nand UO_801 (O_801,N_14793,N_14604);
xnor UO_802 (O_802,N_14781,N_14547);
nand UO_803 (O_803,N_14504,N_14710);
xor UO_804 (O_804,N_14614,N_14822);
nor UO_805 (O_805,N_14741,N_14820);
and UO_806 (O_806,N_14799,N_14564);
and UO_807 (O_807,N_14670,N_14677);
xor UO_808 (O_808,N_14836,N_14828);
xor UO_809 (O_809,N_14772,N_14537);
nand UO_810 (O_810,N_14581,N_14801);
nand UO_811 (O_811,N_14785,N_14837);
xor UO_812 (O_812,N_14992,N_14726);
xnor UO_813 (O_813,N_14544,N_14947);
xor UO_814 (O_814,N_14882,N_14522);
and UO_815 (O_815,N_14806,N_14757);
nand UO_816 (O_816,N_14756,N_14533);
nand UO_817 (O_817,N_14510,N_14512);
nand UO_818 (O_818,N_14650,N_14927);
or UO_819 (O_819,N_14821,N_14712);
and UO_820 (O_820,N_14854,N_14735);
or UO_821 (O_821,N_14998,N_14630);
nand UO_822 (O_822,N_14563,N_14759);
and UO_823 (O_823,N_14822,N_14703);
xor UO_824 (O_824,N_14960,N_14901);
xnor UO_825 (O_825,N_14554,N_14565);
or UO_826 (O_826,N_14939,N_14574);
nor UO_827 (O_827,N_14891,N_14856);
xnor UO_828 (O_828,N_14846,N_14975);
nor UO_829 (O_829,N_14743,N_14567);
and UO_830 (O_830,N_14513,N_14598);
xnor UO_831 (O_831,N_14926,N_14763);
nand UO_832 (O_832,N_14869,N_14963);
and UO_833 (O_833,N_14639,N_14961);
nand UO_834 (O_834,N_14648,N_14970);
xnor UO_835 (O_835,N_14648,N_14659);
and UO_836 (O_836,N_14903,N_14979);
and UO_837 (O_837,N_14717,N_14834);
nand UO_838 (O_838,N_14900,N_14648);
or UO_839 (O_839,N_14533,N_14687);
nand UO_840 (O_840,N_14726,N_14920);
and UO_841 (O_841,N_14661,N_14569);
nor UO_842 (O_842,N_14792,N_14816);
or UO_843 (O_843,N_14509,N_14589);
or UO_844 (O_844,N_14561,N_14960);
or UO_845 (O_845,N_14594,N_14863);
and UO_846 (O_846,N_14958,N_14772);
xor UO_847 (O_847,N_14667,N_14670);
xnor UO_848 (O_848,N_14537,N_14799);
nand UO_849 (O_849,N_14949,N_14813);
xor UO_850 (O_850,N_14967,N_14520);
nor UO_851 (O_851,N_14656,N_14872);
or UO_852 (O_852,N_14752,N_14709);
nor UO_853 (O_853,N_14835,N_14535);
xnor UO_854 (O_854,N_14989,N_14627);
or UO_855 (O_855,N_14639,N_14719);
xor UO_856 (O_856,N_14603,N_14952);
and UO_857 (O_857,N_14552,N_14941);
xor UO_858 (O_858,N_14543,N_14580);
nor UO_859 (O_859,N_14769,N_14830);
nor UO_860 (O_860,N_14755,N_14915);
or UO_861 (O_861,N_14832,N_14725);
nand UO_862 (O_862,N_14607,N_14659);
xor UO_863 (O_863,N_14662,N_14634);
nand UO_864 (O_864,N_14504,N_14619);
nand UO_865 (O_865,N_14876,N_14967);
and UO_866 (O_866,N_14571,N_14790);
and UO_867 (O_867,N_14588,N_14838);
xnor UO_868 (O_868,N_14679,N_14757);
or UO_869 (O_869,N_14608,N_14697);
or UO_870 (O_870,N_14799,N_14739);
nand UO_871 (O_871,N_14523,N_14960);
and UO_872 (O_872,N_14865,N_14699);
and UO_873 (O_873,N_14609,N_14965);
nor UO_874 (O_874,N_14514,N_14503);
and UO_875 (O_875,N_14743,N_14578);
or UO_876 (O_876,N_14519,N_14836);
xor UO_877 (O_877,N_14862,N_14851);
xnor UO_878 (O_878,N_14812,N_14842);
or UO_879 (O_879,N_14659,N_14718);
nand UO_880 (O_880,N_14742,N_14780);
xor UO_881 (O_881,N_14913,N_14630);
xnor UO_882 (O_882,N_14724,N_14866);
nor UO_883 (O_883,N_14803,N_14641);
and UO_884 (O_884,N_14817,N_14855);
or UO_885 (O_885,N_14928,N_14932);
xor UO_886 (O_886,N_14661,N_14845);
and UO_887 (O_887,N_14900,N_14715);
and UO_888 (O_888,N_14855,N_14943);
nor UO_889 (O_889,N_14892,N_14610);
and UO_890 (O_890,N_14562,N_14826);
or UO_891 (O_891,N_14780,N_14776);
or UO_892 (O_892,N_14695,N_14736);
nand UO_893 (O_893,N_14679,N_14829);
nor UO_894 (O_894,N_14759,N_14728);
xor UO_895 (O_895,N_14763,N_14749);
or UO_896 (O_896,N_14856,N_14725);
nor UO_897 (O_897,N_14589,N_14931);
nand UO_898 (O_898,N_14914,N_14648);
and UO_899 (O_899,N_14563,N_14699);
or UO_900 (O_900,N_14948,N_14947);
xor UO_901 (O_901,N_14858,N_14632);
and UO_902 (O_902,N_14790,N_14603);
and UO_903 (O_903,N_14713,N_14938);
xor UO_904 (O_904,N_14635,N_14753);
and UO_905 (O_905,N_14541,N_14511);
nor UO_906 (O_906,N_14573,N_14868);
xnor UO_907 (O_907,N_14853,N_14801);
nor UO_908 (O_908,N_14557,N_14874);
xnor UO_909 (O_909,N_14812,N_14698);
and UO_910 (O_910,N_14757,N_14821);
xnor UO_911 (O_911,N_14919,N_14690);
and UO_912 (O_912,N_14732,N_14623);
or UO_913 (O_913,N_14813,N_14870);
nor UO_914 (O_914,N_14985,N_14808);
nor UO_915 (O_915,N_14825,N_14906);
and UO_916 (O_916,N_14920,N_14673);
nand UO_917 (O_917,N_14909,N_14798);
or UO_918 (O_918,N_14929,N_14610);
nand UO_919 (O_919,N_14624,N_14902);
nand UO_920 (O_920,N_14809,N_14532);
and UO_921 (O_921,N_14826,N_14775);
nand UO_922 (O_922,N_14795,N_14791);
nor UO_923 (O_923,N_14567,N_14935);
nand UO_924 (O_924,N_14728,N_14962);
and UO_925 (O_925,N_14898,N_14682);
xnor UO_926 (O_926,N_14922,N_14691);
nor UO_927 (O_927,N_14805,N_14828);
or UO_928 (O_928,N_14573,N_14879);
or UO_929 (O_929,N_14522,N_14966);
xor UO_930 (O_930,N_14823,N_14567);
xor UO_931 (O_931,N_14866,N_14915);
nand UO_932 (O_932,N_14504,N_14925);
xnor UO_933 (O_933,N_14950,N_14852);
nor UO_934 (O_934,N_14751,N_14534);
xor UO_935 (O_935,N_14660,N_14939);
xnor UO_936 (O_936,N_14695,N_14597);
xor UO_937 (O_937,N_14633,N_14558);
nor UO_938 (O_938,N_14925,N_14793);
xor UO_939 (O_939,N_14735,N_14721);
xor UO_940 (O_940,N_14918,N_14598);
nand UO_941 (O_941,N_14673,N_14916);
xnor UO_942 (O_942,N_14543,N_14515);
nand UO_943 (O_943,N_14777,N_14846);
nand UO_944 (O_944,N_14885,N_14969);
xnor UO_945 (O_945,N_14970,N_14880);
and UO_946 (O_946,N_14847,N_14525);
nor UO_947 (O_947,N_14991,N_14557);
nor UO_948 (O_948,N_14900,N_14807);
nand UO_949 (O_949,N_14709,N_14536);
nand UO_950 (O_950,N_14650,N_14822);
xnor UO_951 (O_951,N_14539,N_14920);
xor UO_952 (O_952,N_14601,N_14640);
nand UO_953 (O_953,N_14766,N_14726);
nand UO_954 (O_954,N_14671,N_14757);
xnor UO_955 (O_955,N_14752,N_14734);
and UO_956 (O_956,N_14763,N_14753);
nor UO_957 (O_957,N_14967,N_14683);
and UO_958 (O_958,N_14907,N_14918);
and UO_959 (O_959,N_14629,N_14734);
nand UO_960 (O_960,N_14806,N_14926);
and UO_961 (O_961,N_14927,N_14615);
or UO_962 (O_962,N_14775,N_14637);
nand UO_963 (O_963,N_14700,N_14579);
nand UO_964 (O_964,N_14785,N_14779);
and UO_965 (O_965,N_14674,N_14530);
nor UO_966 (O_966,N_14995,N_14552);
and UO_967 (O_967,N_14929,N_14821);
nor UO_968 (O_968,N_14795,N_14861);
nor UO_969 (O_969,N_14860,N_14972);
xor UO_970 (O_970,N_14536,N_14967);
nand UO_971 (O_971,N_14542,N_14831);
nor UO_972 (O_972,N_14588,N_14751);
and UO_973 (O_973,N_14740,N_14559);
or UO_974 (O_974,N_14972,N_14776);
and UO_975 (O_975,N_14758,N_14997);
nor UO_976 (O_976,N_14639,N_14630);
or UO_977 (O_977,N_14954,N_14507);
nand UO_978 (O_978,N_14710,N_14524);
xor UO_979 (O_979,N_14834,N_14739);
nor UO_980 (O_980,N_14923,N_14698);
nor UO_981 (O_981,N_14720,N_14858);
nand UO_982 (O_982,N_14516,N_14698);
nand UO_983 (O_983,N_14761,N_14882);
nor UO_984 (O_984,N_14937,N_14885);
nor UO_985 (O_985,N_14832,N_14847);
and UO_986 (O_986,N_14799,N_14956);
xor UO_987 (O_987,N_14779,N_14941);
or UO_988 (O_988,N_14575,N_14591);
nand UO_989 (O_989,N_14910,N_14544);
or UO_990 (O_990,N_14853,N_14812);
or UO_991 (O_991,N_14718,N_14607);
xor UO_992 (O_992,N_14520,N_14711);
and UO_993 (O_993,N_14968,N_14879);
xnor UO_994 (O_994,N_14708,N_14751);
nand UO_995 (O_995,N_14772,N_14669);
and UO_996 (O_996,N_14509,N_14907);
and UO_997 (O_997,N_14688,N_14521);
nor UO_998 (O_998,N_14853,N_14566);
nor UO_999 (O_999,N_14520,N_14820);
xor UO_1000 (O_1000,N_14720,N_14625);
and UO_1001 (O_1001,N_14808,N_14869);
nand UO_1002 (O_1002,N_14996,N_14510);
xor UO_1003 (O_1003,N_14523,N_14772);
nor UO_1004 (O_1004,N_14969,N_14633);
or UO_1005 (O_1005,N_14716,N_14889);
xor UO_1006 (O_1006,N_14876,N_14741);
nor UO_1007 (O_1007,N_14743,N_14964);
or UO_1008 (O_1008,N_14532,N_14501);
nand UO_1009 (O_1009,N_14699,N_14564);
nand UO_1010 (O_1010,N_14945,N_14804);
nand UO_1011 (O_1011,N_14749,N_14825);
nor UO_1012 (O_1012,N_14844,N_14703);
and UO_1013 (O_1013,N_14507,N_14930);
or UO_1014 (O_1014,N_14886,N_14720);
nor UO_1015 (O_1015,N_14697,N_14617);
xnor UO_1016 (O_1016,N_14734,N_14641);
nand UO_1017 (O_1017,N_14511,N_14568);
and UO_1018 (O_1018,N_14698,N_14795);
or UO_1019 (O_1019,N_14540,N_14609);
nand UO_1020 (O_1020,N_14523,N_14660);
xor UO_1021 (O_1021,N_14834,N_14725);
nand UO_1022 (O_1022,N_14601,N_14568);
and UO_1023 (O_1023,N_14608,N_14976);
and UO_1024 (O_1024,N_14748,N_14894);
or UO_1025 (O_1025,N_14920,N_14596);
nand UO_1026 (O_1026,N_14826,N_14564);
and UO_1027 (O_1027,N_14812,N_14591);
or UO_1028 (O_1028,N_14749,N_14833);
nand UO_1029 (O_1029,N_14738,N_14634);
nand UO_1030 (O_1030,N_14594,N_14786);
nand UO_1031 (O_1031,N_14571,N_14817);
nor UO_1032 (O_1032,N_14706,N_14505);
xnor UO_1033 (O_1033,N_14885,N_14580);
nand UO_1034 (O_1034,N_14847,N_14636);
or UO_1035 (O_1035,N_14973,N_14597);
and UO_1036 (O_1036,N_14636,N_14605);
xor UO_1037 (O_1037,N_14741,N_14736);
nor UO_1038 (O_1038,N_14917,N_14913);
nand UO_1039 (O_1039,N_14659,N_14989);
and UO_1040 (O_1040,N_14834,N_14978);
nor UO_1041 (O_1041,N_14942,N_14666);
xor UO_1042 (O_1042,N_14562,N_14683);
nor UO_1043 (O_1043,N_14814,N_14662);
nand UO_1044 (O_1044,N_14870,N_14539);
and UO_1045 (O_1045,N_14680,N_14618);
nor UO_1046 (O_1046,N_14957,N_14565);
xor UO_1047 (O_1047,N_14950,N_14580);
nand UO_1048 (O_1048,N_14685,N_14898);
xnor UO_1049 (O_1049,N_14747,N_14630);
xnor UO_1050 (O_1050,N_14988,N_14958);
nand UO_1051 (O_1051,N_14859,N_14629);
xor UO_1052 (O_1052,N_14555,N_14618);
nand UO_1053 (O_1053,N_14698,N_14908);
or UO_1054 (O_1054,N_14604,N_14548);
or UO_1055 (O_1055,N_14711,N_14838);
nand UO_1056 (O_1056,N_14864,N_14875);
and UO_1057 (O_1057,N_14589,N_14899);
nand UO_1058 (O_1058,N_14887,N_14877);
or UO_1059 (O_1059,N_14892,N_14853);
nor UO_1060 (O_1060,N_14810,N_14881);
nand UO_1061 (O_1061,N_14807,N_14693);
nor UO_1062 (O_1062,N_14612,N_14936);
and UO_1063 (O_1063,N_14515,N_14572);
nand UO_1064 (O_1064,N_14583,N_14647);
nand UO_1065 (O_1065,N_14531,N_14669);
and UO_1066 (O_1066,N_14702,N_14705);
or UO_1067 (O_1067,N_14811,N_14645);
or UO_1068 (O_1068,N_14727,N_14976);
nor UO_1069 (O_1069,N_14905,N_14614);
nor UO_1070 (O_1070,N_14971,N_14594);
xor UO_1071 (O_1071,N_14909,N_14655);
and UO_1072 (O_1072,N_14676,N_14555);
xor UO_1073 (O_1073,N_14883,N_14839);
and UO_1074 (O_1074,N_14563,N_14672);
nand UO_1075 (O_1075,N_14692,N_14902);
nor UO_1076 (O_1076,N_14812,N_14820);
or UO_1077 (O_1077,N_14757,N_14873);
nor UO_1078 (O_1078,N_14704,N_14982);
or UO_1079 (O_1079,N_14900,N_14918);
xor UO_1080 (O_1080,N_14739,N_14861);
and UO_1081 (O_1081,N_14618,N_14972);
or UO_1082 (O_1082,N_14503,N_14807);
or UO_1083 (O_1083,N_14730,N_14537);
and UO_1084 (O_1084,N_14788,N_14675);
nor UO_1085 (O_1085,N_14864,N_14662);
xor UO_1086 (O_1086,N_14533,N_14761);
and UO_1087 (O_1087,N_14594,N_14842);
nor UO_1088 (O_1088,N_14718,N_14529);
nand UO_1089 (O_1089,N_14503,N_14930);
nor UO_1090 (O_1090,N_14532,N_14541);
xor UO_1091 (O_1091,N_14605,N_14596);
xor UO_1092 (O_1092,N_14631,N_14799);
and UO_1093 (O_1093,N_14518,N_14894);
nor UO_1094 (O_1094,N_14538,N_14850);
or UO_1095 (O_1095,N_14998,N_14987);
and UO_1096 (O_1096,N_14649,N_14743);
nor UO_1097 (O_1097,N_14830,N_14516);
and UO_1098 (O_1098,N_14897,N_14812);
or UO_1099 (O_1099,N_14591,N_14821);
xor UO_1100 (O_1100,N_14787,N_14576);
xor UO_1101 (O_1101,N_14751,N_14977);
nor UO_1102 (O_1102,N_14516,N_14699);
or UO_1103 (O_1103,N_14873,N_14994);
xnor UO_1104 (O_1104,N_14597,N_14805);
xnor UO_1105 (O_1105,N_14621,N_14773);
and UO_1106 (O_1106,N_14945,N_14608);
and UO_1107 (O_1107,N_14945,N_14710);
and UO_1108 (O_1108,N_14719,N_14850);
nor UO_1109 (O_1109,N_14548,N_14854);
xor UO_1110 (O_1110,N_14547,N_14579);
and UO_1111 (O_1111,N_14659,N_14874);
xor UO_1112 (O_1112,N_14511,N_14530);
and UO_1113 (O_1113,N_14751,N_14539);
nand UO_1114 (O_1114,N_14691,N_14532);
nand UO_1115 (O_1115,N_14748,N_14719);
and UO_1116 (O_1116,N_14890,N_14637);
or UO_1117 (O_1117,N_14771,N_14692);
xor UO_1118 (O_1118,N_14899,N_14538);
nor UO_1119 (O_1119,N_14582,N_14886);
nor UO_1120 (O_1120,N_14577,N_14615);
and UO_1121 (O_1121,N_14649,N_14535);
nand UO_1122 (O_1122,N_14906,N_14963);
nand UO_1123 (O_1123,N_14536,N_14753);
nor UO_1124 (O_1124,N_14853,N_14608);
xor UO_1125 (O_1125,N_14725,N_14586);
nand UO_1126 (O_1126,N_14671,N_14833);
and UO_1127 (O_1127,N_14950,N_14609);
and UO_1128 (O_1128,N_14998,N_14782);
and UO_1129 (O_1129,N_14573,N_14910);
nand UO_1130 (O_1130,N_14730,N_14797);
nor UO_1131 (O_1131,N_14829,N_14702);
and UO_1132 (O_1132,N_14545,N_14770);
and UO_1133 (O_1133,N_14641,N_14696);
nor UO_1134 (O_1134,N_14814,N_14633);
or UO_1135 (O_1135,N_14576,N_14592);
nand UO_1136 (O_1136,N_14753,N_14834);
or UO_1137 (O_1137,N_14664,N_14810);
or UO_1138 (O_1138,N_14503,N_14830);
nand UO_1139 (O_1139,N_14914,N_14675);
xnor UO_1140 (O_1140,N_14659,N_14634);
or UO_1141 (O_1141,N_14808,N_14500);
or UO_1142 (O_1142,N_14977,N_14844);
and UO_1143 (O_1143,N_14715,N_14746);
nor UO_1144 (O_1144,N_14620,N_14553);
nor UO_1145 (O_1145,N_14903,N_14774);
nor UO_1146 (O_1146,N_14617,N_14528);
and UO_1147 (O_1147,N_14969,N_14750);
and UO_1148 (O_1148,N_14825,N_14812);
or UO_1149 (O_1149,N_14561,N_14535);
nand UO_1150 (O_1150,N_14824,N_14874);
and UO_1151 (O_1151,N_14945,N_14920);
and UO_1152 (O_1152,N_14972,N_14751);
nor UO_1153 (O_1153,N_14964,N_14643);
and UO_1154 (O_1154,N_14886,N_14706);
and UO_1155 (O_1155,N_14681,N_14713);
and UO_1156 (O_1156,N_14974,N_14848);
and UO_1157 (O_1157,N_14964,N_14851);
nand UO_1158 (O_1158,N_14570,N_14880);
nor UO_1159 (O_1159,N_14947,N_14819);
nor UO_1160 (O_1160,N_14565,N_14511);
xor UO_1161 (O_1161,N_14683,N_14695);
or UO_1162 (O_1162,N_14673,N_14776);
nor UO_1163 (O_1163,N_14747,N_14872);
nor UO_1164 (O_1164,N_14631,N_14785);
nand UO_1165 (O_1165,N_14772,N_14757);
and UO_1166 (O_1166,N_14781,N_14870);
or UO_1167 (O_1167,N_14786,N_14807);
xor UO_1168 (O_1168,N_14922,N_14740);
and UO_1169 (O_1169,N_14910,N_14978);
xnor UO_1170 (O_1170,N_14615,N_14701);
nor UO_1171 (O_1171,N_14858,N_14863);
nor UO_1172 (O_1172,N_14783,N_14988);
xor UO_1173 (O_1173,N_14878,N_14991);
nor UO_1174 (O_1174,N_14537,N_14531);
and UO_1175 (O_1175,N_14929,N_14904);
or UO_1176 (O_1176,N_14946,N_14573);
nor UO_1177 (O_1177,N_14679,N_14891);
and UO_1178 (O_1178,N_14707,N_14506);
and UO_1179 (O_1179,N_14703,N_14830);
xor UO_1180 (O_1180,N_14967,N_14868);
nand UO_1181 (O_1181,N_14713,N_14821);
and UO_1182 (O_1182,N_14825,N_14508);
or UO_1183 (O_1183,N_14545,N_14517);
and UO_1184 (O_1184,N_14971,N_14917);
or UO_1185 (O_1185,N_14547,N_14631);
xor UO_1186 (O_1186,N_14561,N_14922);
or UO_1187 (O_1187,N_14918,N_14748);
and UO_1188 (O_1188,N_14616,N_14961);
nor UO_1189 (O_1189,N_14762,N_14960);
or UO_1190 (O_1190,N_14783,N_14947);
and UO_1191 (O_1191,N_14711,N_14726);
or UO_1192 (O_1192,N_14928,N_14655);
nor UO_1193 (O_1193,N_14929,N_14868);
xnor UO_1194 (O_1194,N_14793,N_14784);
nor UO_1195 (O_1195,N_14774,N_14821);
nand UO_1196 (O_1196,N_14790,N_14647);
nand UO_1197 (O_1197,N_14845,N_14683);
nor UO_1198 (O_1198,N_14518,N_14586);
nand UO_1199 (O_1199,N_14637,N_14558);
and UO_1200 (O_1200,N_14566,N_14596);
xnor UO_1201 (O_1201,N_14759,N_14979);
nor UO_1202 (O_1202,N_14994,N_14641);
and UO_1203 (O_1203,N_14508,N_14710);
nor UO_1204 (O_1204,N_14629,N_14906);
or UO_1205 (O_1205,N_14830,N_14857);
xnor UO_1206 (O_1206,N_14767,N_14662);
nor UO_1207 (O_1207,N_14969,N_14940);
nor UO_1208 (O_1208,N_14687,N_14581);
or UO_1209 (O_1209,N_14761,N_14970);
or UO_1210 (O_1210,N_14531,N_14905);
xnor UO_1211 (O_1211,N_14650,N_14500);
and UO_1212 (O_1212,N_14646,N_14872);
nor UO_1213 (O_1213,N_14539,N_14543);
nand UO_1214 (O_1214,N_14584,N_14970);
and UO_1215 (O_1215,N_14901,N_14616);
xor UO_1216 (O_1216,N_14642,N_14964);
or UO_1217 (O_1217,N_14708,N_14522);
xnor UO_1218 (O_1218,N_14965,N_14964);
or UO_1219 (O_1219,N_14655,N_14648);
or UO_1220 (O_1220,N_14642,N_14942);
or UO_1221 (O_1221,N_14983,N_14711);
and UO_1222 (O_1222,N_14645,N_14805);
xnor UO_1223 (O_1223,N_14645,N_14722);
or UO_1224 (O_1224,N_14873,N_14758);
or UO_1225 (O_1225,N_14513,N_14509);
xnor UO_1226 (O_1226,N_14993,N_14635);
and UO_1227 (O_1227,N_14613,N_14504);
and UO_1228 (O_1228,N_14881,N_14533);
and UO_1229 (O_1229,N_14712,N_14795);
and UO_1230 (O_1230,N_14573,N_14508);
nor UO_1231 (O_1231,N_14719,N_14645);
nor UO_1232 (O_1232,N_14857,N_14939);
and UO_1233 (O_1233,N_14859,N_14872);
or UO_1234 (O_1234,N_14624,N_14719);
xnor UO_1235 (O_1235,N_14803,N_14791);
nand UO_1236 (O_1236,N_14570,N_14929);
nor UO_1237 (O_1237,N_14837,N_14697);
nand UO_1238 (O_1238,N_14991,N_14783);
nand UO_1239 (O_1239,N_14685,N_14931);
nor UO_1240 (O_1240,N_14656,N_14748);
or UO_1241 (O_1241,N_14667,N_14815);
and UO_1242 (O_1242,N_14853,N_14513);
and UO_1243 (O_1243,N_14621,N_14928);
xnor UO_1244 (O_1244,N_14781,N_14590);
xor UO_1245 (O_1245,N_14757,N_14516);
xor UO_1246 (O_1246,N_14551,N_14764);
and UO_1247 (O_1247,N_14850,N_14985);
nor UO_1248 (O_1248,N_14961,N_14949);
nand UO_1249 (O_1249,N_14983,N_14876);
and UO_1250 (O_1250,N_14556,N_14805);
or UO_1251 (O_1251,N_14967,N_14851);
nor UO_1252 (O_1252,N_14621,N_14807);
nand UO_1253 (O_1253,N_14903,N_14818);
nor UO_1254 (O_1254,N_14837,N_14711);
nand UO_1255 (O_1255,N_14966,N_14520);
and UO_1256 (O_1256,N_14949,N_14544);
xor UO_1257 (O_1257,N_14613,N_14529);
or UO_1258 (O_1258,N_14544,N_14901);
nor UO_1259 (O_1259,N_14994,N_14579);
nand UO_1260 (O_1260,N_14687,N_14587);
or UO_1261 (O_1261,N_14968,N_14871);
nor UO_1262 (O_1262,N_14726,N_14968);
and UO_1263 (O_1263,N_14937,N_14976);
nand UO_1264 (O_1264,N_14702,N_14522);
and UO_1265 (O_1265,N_14848,N_14705);
and UO_1266 (O_1266,N_14665,N_14939);
or UO_1267 (O_1267,N_14965,N_14533);
and UO_1268 (O_1268,N_14742,N_14530);
or UO_1269 (O_1269,N_14601,N_14848);
nand UO_1270 (O_1270,N_14627,N_14790);
or UO_1271 (O_1271,N_14701,N_14564);
nand UO_1272 (O_1272,N_14933,N_14921);
nor UO_1273 (O_1273,N_14564,N_14602);
or UO_1274 (O_1274,N_14857,N_14849);
and UO_1275 (O_1275,N_14841,N_14627);
xor UO_1276 (O_1276,N_14715,N_14806);
or UO_1277 (O_1277,N_14852,N_14895);
or UO_1278 (O_1278,N_14778,N_14543);
xor UO_1279 (O_1279,N_14772,N_14844);
or UO_1280 (O_1280,N_14797,N_14882);
nor UO_1281 (O_1281,N_14502,N_14994);
nor UO_1282 (O_1282,N_14696,N_14524);
nand UO_1283 (O_1283,N_14556,N_14639);
xor UO_1284 (O_1284,N_14653,N_14611);
nand UO_1285 (O_1285,N_14700,N_14671);
or UO_1286 (O_1286,N_14541,N_14564);
nand UO_1287 (O_1287,N_14729,N_14684);
or UO_1288 (O_1288,N_14622,N_14980);
nand UO_1289 (O_1289,N_14829,N_14996);
or UO_1290 (O_1290,N_14594,N_14623);
or UO_1291 (O_1291,N_14983,N_14807);
nand UO_1292 (O_1292,N_14771,N_14705);
and UO_1293 (O_1293,N_14581,N_14976);
nor UO_1294 (O_1294,N_14940,N_14698);
nand UO_1295 (O_1295,N_14900,N_14621);
nor UO_1296 (O_1296,N_14528,N_14757);
xor UO_1297 (O_1297,N_14660,N_14876);
nand UO_1298 (O_1298,N_14964,N_14860);
nor UO_1299 (O_1299,N_14888,N_14781);
and UO_1300 (O_1300,N_14853,N_14656);
nand UO_1301 (O_1301,N_14568,N_14789);
or UO_1302 (O_1302,N_14749,N_14971);
xor UO_1303 (O_1303,N_14707,N_14943);
xnor UO_1304 (O_1304,N_14872,N_14643);
nand UO_1305 (O_1305,N_14682,N_14944);
and UO_1306 (O_1306,N_14674,N_14946);
or UO_1307 (O_1307,N_14631,N_14915);
nor UO_1308 (O_1308,N_14507,N_14613);
nand UO_1309 (O_1309,N_14752,N_14547);
or UO_1310 (O_1310,N_14842,N_14889);
nand UO_1311 (O_1311,N_14752,N_14776);
xor UO_1312 (O_1312,N_14707,N_14722);
xnor UO_1313 (O_1313,N_14591,N_14942);
or UO_1314 (O_1314,N_14700,N_14771);
nand UO_1315 (O_1315,N_14735,N_14577);
or UO_1316 (O_1316,N_14868,N_14898);
xnor UO_1317 (O_1317,N_14976,N_14684);
nor UO_1318 (O_1318,N_14620,N_14935);
nor UO_1319 (O_1319,N_14568,N_14911);
nand UO_1320 (O_1320,N_14806,N_14951);
nor UO_1321 (O_1321,N_14675,N_14753);
or UO_1322 (O_1322,N_14873,N_14917);
nor UO_1323 (O_1323,N_14796,N_14955);
nor UO_1324 (O_1324,N_14925,N_14871);
nor UO_1325 (O_1325,N_14991,N_14996);
nand UO_1326 (O_1326,N_14760,N_14703);
nor UO_1327 (O_1327,N_14814,N_14651);
nor UO_1328 (O_1328,N_14868,N_14873);
or UO_1329 (O_1329,N_14919,N_14812);
nor UO_1330 (O_1330,N_14808,N_14872);
and UO_1331 (O_1331,N_14634,N_14930);
nand UO_1332 (O_1332,N_14941,N_14719);
and UO_1333 (O_1333,N_14882,N_14623);
and UO_1334 (O_1334,N_14727,N_14606);
and UO_1335 (O_1335,N_14863,N_14932);
and UO_1336 (O_1336,N_14643,N_14529);
and UO_1337 (O_1337,N_14757,N_14877);
nand UO_1338 (O_1338,N_14585,N_14548);
xnor UO_1339 (O_1339,N_14583,N_14887);
nand UO_1340 (O_1340,N_14785,N_14650);
or UO_1341 (O_1341,N_14555,N_14617);
nand UO_1342 (O_1342,N_14576,N_14988);
nand UO_1343 (O_1343,N_14798,N_14666);
or UO_1344 (O_1344,N_14691,N_14740);
and UO_1345 (O_1345,N_14679,N_14894);
nand UO_1346 (O_1346,N_14685,N_14779);
nand UO_1347 (O_1347,N_14668,N_14648);
xnor UO_1348 (O_1348,N_14954,N_14617);
xnor UO_1349 (O_1349,N_14687,N_14849);
and UO_1350 (O_1350,N_14574,N_14922);
and UO_1351 (O_1351,N_14806,N_14907);
and UO_1352 (O_1352,N_14709,N_14844);
nand UO_1353 (O_1353,N_14627,N_14504);
nand UO_1354 (O_1354,N_14900,N_14673);
nand UO_1355 (O_1355,N_14540,N_14544);
nor UO_1356 (O_1356,N_14904,N_14588);
nand UO_1357 (O_1357,N_14832,N_14603);
nor UO_1358 (O_1358,N_14838,N_14979);
nand UO_1359 (O_1359,N_14729,N_14825);
nand UO_1360 (O_1360,N_14531,N_14558);
nor UO_1361 (O_1361,N_14540,N_14926);
xnor UO_1362 (O_1362,N_14740,N_14810);
nor UO_1363 (O_1363,N_14626,N_14637);
and UO_1364 (O_1364,N_14624,N_14878);
xor UO_1365 (O_1365,N_14948,N_14688);
and UO_1366 (O_1366,N_14620,N_14824);
xor UO_1367 (O_1367,N_14759,N_14938);
nor UO_1368 (O_1368,N_14575,N_14505);
or UO_1369 (O_1369,N_14995,N_14955);
and UO_1370 (O_1370,N_14670,N_14994);
nand UO_1371 (O_1371,N_14691,N_14990);
and UO_1372 (O_1372,N_14652,N_14733);
nor UO_1373 (O_1373,N_14981,N_14982);
nand UO_1374 (O_1374,N_14749,N_14981);
nor UO_1375 (O_1375,N_14714,N_14878);
and UO_1376 (O_1376,N_14571,N_14942);
nor UO_1377 (O_1377,N_14558,N_14720);
xor UO_1378 (O_1378,N_14863,N_14859);
nor UO_1379 (O_1379,N_14602,N_14821);
nand UO_1380 (O_1380,N_14691,N_14711);
nand UO_1381 (O_1381,N_14594,N_14779);
nor UO_1382 (O_1382,N_14996,N_14803);
nor UO_1383 (O_1383,N_14792,N_14991);
nor UO_1384 (O_1384,N_14677,N_14782);
nor UO_1385 (O_1385,N_14756,N_14620);
nor UO_1386 (O_1386,N_14777,N_14758);
and UO_1387 (O_1387,N_14836,N_14590);
or UO_1388 (O_1388,N_14548,N_14678);
and UO_1389 (O_1389,N_14780,N_14530);
or UO_1390 (O_1390,N_14522,N_14687);
and UO_1391 (O_1391,N_14633,N_14924);
or UO_1392 (O_1392,N_14860,N_14631);
xnor UO_1393 (O_1393,N_14608,N_14549);
nor UO_1394 (O_1394,N_14814,N_14626);
nand UO_1395 (O_1395,N_14992,N_14576);
or UO_1396 (O_1396,N_14697,N_14881);
nand UO_1397 (O_1397,N_14567,N_14696);
and UO_1398 (O_1398,N_14696,N_14703);
and UO_1399 (O_1399,N_14692,N_14823);
and UO_1400 (O_1400,N_14539,N_14884);
and UO_1401 (O_1401,N_14522,N_14603);
nand UO_1402 (O_1402,N_14639,N_14962);
xnor UO_1403 (O_1403,N_14587,N_14812);
xnor UO_1404 (O_1404,N_14832,N_14952);
xnor UO_1405 (O_1405,N_14759,N_14838);
and UO_1406 (O_1406,N_14674,N_14600);
or UO_1407 (O_1407,N_14554,N_14677);
nand UO_1408 (O_1408,N_14745,N_14785);
nand UO_1409 (O_1409,N_14840,N_14824);
nand UO_1410 (O_1410,N_14717,N_14847);
nand UO_1411 (O_1411,N_14600,N_14816);
and UO_1412 (O_1412,N_14837,N_14975);
nand UO_1413 (O_1413,N_14775,N_14701);
and UO_1414 (O_1414,N_14949,N_14507);
or UO_1415 (O_1415,N_14552,N_14863);
nor UO_1416 (O_1416,N_14782,N_14546);
xor UO_1417 (O_1417,N_14975,N_14729);
or UO_1418 (O_1418,N_14507,N_14812);
or UO_1419 (O_1419,N_14519,N_14917);
or UO_1420 (O_1420,N_14839,N_14758);
or UO_1421 (O_1421,N_14998,N_14645);
xnor UO_1422 (O_1422,N_14793,N_14504);
nor UO_1423 (O_1423,N_14759,N_14758);
nor UO_1424 (O_1424,N_14740,N_14549);
and UO_1425 (O_1425,N_14620,N_14936);
or UO_1426 (O_1426,N_14784,N_14851);
or UO_1427 (O_1427,N_14839,N_14524);
xor UO_1428 (O_1428,N_14665,N_14517);
or UO_1429 (O_1429,N_14964,N_14597);
or UO_1430 (O_1430,N_14800,N_14999);
or UO_1431 (O_1431,N_14804,N_14860);
nand UO_1432 (O_1432,N_14883,N_14788);
nor UO_1433 (O_1433,N_14743,N_14657);
or UO_1434 (O_1434,N_14611,N_14721);
nand UO_1435 (O_1435,N_14804,N_14676);
or UO_1436 (O_1436,N_14955,N_14559);
nand UO_1437 (O_1437,N_14970,N_14923);
nand UO_1438 (O_1438,N_14675,N_14772);
or UO_1439 (O_1439,N_14969,N_14752);
and UO_1440 (O_1440,N_14543,N_14922);
nand UO_1441 (O_1441,N_14574,N_14826);
and UO_1442 (O_1442,N_14608,N_14710);
nand UO_1443 (O_1443,N_14787,N_14591);
xor UO_1444 (O_1444,N_14699,N_14588);
nand UO_1445 (O_1445,N_14849,N_14514);
or UO_1446 (O_1446,N_14685,N_14514);
nand UO_1447 (O_1447,N_14803,N_14571);
or UO_1448 (O_1448,N_14589,N_14538);
and UO_1449 (O_1449,N_14505,N_14597);
nand UO_1450 (O_1450,N_14833,N_14920);
and UO_1451 (O_1451,N_14537,N_14735);
and UO_1452 (O_1452,N_14968,N_14965);
or UO_1453 (O_1453,N_14504,N_14988);
nand UO_1454 (O_1454,N_14762,N_14906);
xor UO_1455 (O_1455,N_14982,N_14977);
and UO_1456 (O_1456,N_14633,N_14820);
and UO_1457 (O_1457,N_14886,N_14913);
xor UO_1458 (O_1458,N_14791,N_14588);
and UO_1459 (O_1459,N_14688,N_14963);
or UO_1460 (O_1460,N_14652,N_14840);
nor UO_1461 (O_1461,N_14584,N_14880);
nor UO_1462 (O_1462,N_14507,N_14573);
and UO_1463 (O_1463,N_14520,N_14620);
or UO_1464 (O_1464,N_14963,N_14805);
xnor UO_1465 (O_1465,N_14609,N_14720);
xor UO_1466 (O_1466,N_14911,N_14703);
nand UO_1467 (O_1467,N_14555,N_14769);
nand UO_1468 (O_1468,N_14602,N_14816);
nand UO_1469 (O_1469,N_14726,N_14894);
nor UO_1470 (O_1470,N_14825,N_14712);
nor UO_1471 (O_1471,N_14881,N_14756);
or UO_1472 (O_1472,N_14567,N_14864);
or UO_1473 (O_1473,N_14587,N_14898);
or UO_1474 (O_1474,N_14838,N_14787);
nand UO_1475 (O_1475,N_14953,N_14927);
nand UO_1476 (O_1476,N_14548,N_14852);
nor UO_1477 (O_1477,N_14725,N_14918);
xor UO_1478 (O_1478,N_14767,N_14591);
and UO_1479 (O_1479,N_14889,N_14927);
or UO_1480 (O_1480,N_14559,N_14599);
nand UO_1481 (O_1481,N_14646,N_14986);
or UO_1482 (O_1482,N_14704,N_14990);
xor UO_1483 (O_1483,N_14882,N_14733);
and UO_1484 (O_1484,N_14836,N_14535);
xnor UO_1485 (O_1485,N_14615,N_14503);
or UO_1486 (O_1486,N_14864,N_14582);
xnor UO_1487 (O_1487,N_14765,N_14612);
nor UO_1488 (O_1488,N_14904,N_14749);
or UO_1489 (O_1489,N_14691,N_14713);
nor UO_1490 (O_1490,N_14898,N_14877);
and UO_1491 (O_1491,N_14610,N_14659);
xor UO_1492 (O_1492,N_14960,N_14624);
nor UO_1493 (O_1493,N_14535,N_14774);
and UO_1494 (O_1494,N_14552,N_14620);
nor UO_1495 (O_1495,N_14590,N_14623);
and UO_1496 (O_1496,N_14654,N_14942);
and UO_1497 (O_1497,N_14614,N_14972);
xor UO_1498 (O_1498,N_14663,N_14764);
and UO_1499 (O_1499,N_14997,N_14946);
xor UO_1500 (O_1500,N_14716,N_14885);
xor UO_1501 (O_1501,N_14958,N_14666);
and UO_1502 (O_1502,N_14734,N_14729);
xnor UO_1503 (O_1503,N_14535,N_14792);
or UO_1504 (O_1504,N_14741,N_14838);
nor UO_1505 (O_1505,N_14755,N_14575);
nand UO_1506 (O_1506,N_14887,N_14813);
xnor UO_1507 (O_1507,N_14621,N_14665);
or UO_1508 (O_1508,N_14646,N_14723);
nor UO_1509 (O_1509,N_14925,N_14956);
or UO_1510 (O_1510,N_14791,N_14815);
nand UO_1511 (O_1511,N_14957,N_14846);
nor UO_1512 (O_1512,N_14884,N_14981);
nand UO_1513 (O_1513,N_14661,N_14906);
or UO_1514 (O_1514,N_14921,N_14615);
xnor UO_1515 (O_1515,N_14720,N_14797);
xor UO_1516 (O_1516,N_14948,N_14612);
xor UO_1517 (O_1517,N_14555,N_14554);
nand UO_1518 (O_1518,N_14817,N_14772);
or UO_1519 (O_1519,N_14889,N_14527);
and UO_1520 (O_1520,N_14567,N_14865);
and UO_1521 (O_1521,N_14880,N_14628);
or UO_1522 (O_1522,N_14564,N_14800);
nand UO_1523 (O_1523,N_14850,N_14695);
xor UO_1524 (O_1524,N_14725,N_14502);
nand UO_1525 (O_1525,N_14674,N_14810);
or UO_1526 (O_1526,N_14922,N_14831);
or UO_1527 (O_1527,N_14754,N_14929);
or UO_1528 (O_1528,N_14569,N_14694);
nor UO_1529 (O_1529,N_14643,N_14830);
nor UO_1530 (O_1530,N_14718,N_14753);
xnor UO_1531 (O_1531,N_14939,N_14880);
or UO_1532 (O_1532,N_14823,N_14536);
and UO_1533 (O_1533,N_14717,N_14883);
xnor UO_1534 (O_1534,N_14617,N_14933);
nand UO_1535 (O_1535,N_14910,N_14997);
nand UO_1536 (O_1536,N_14517,N_14979);
nor UO_1537 (O_1537,N_14889,N_14775);
xnor UO_1538 (O_1538,N_14663,N_14800);
nand UO_1539 (O_1539,N_14636,N_14899);
nand UO_1540 (O_1540,N_14861,N_14564);
nor UO_1541 (O_1541,N_14549,N_14694);
nor UO_1542 (O_1542,N_14985,N_14738);
or UO_1543 (O_1543,N_14848,N_14681);
or UO_1544 (O_1544,N_14615,N_14913);
nor UO_1545 (O_1545,N_14797,N_14795);
nand UO_1546 (O_1546,N_14500,N_14574);
nand UO_1547 (O_1547,N_14976,N_14899);
xnor UO_1548 (O_1548,N_14724,N_14929);
and UO_1549 (O_1549,N_14589,N_14695);
or UO_1550 (O_1550,N_14567,N_14820);
and UO_1551 (O_1551,N_14716,N_14530);
nor UO_1552 (O_1552,N_14750,N_14883);
or UO_1553 (O_1553,N_14558,N_14664);
nor UO_1554 (O_1554,N_14746,N_14995);
and UO_1555 (O_1555,N_14708,N_14587);
and UO_1556 (O_1556,N_14679,N_14874);
and UO_1557 (O_1557,N_14955,N_14655);
nand UO_1558 (O_1558,N_14571,N_14852);
and UO_1559 (O_1559,N_14819,N_14912);
nand UO_1560 (O_1560,N_14873,N_14542);
and UO_1561 (O_1561,N_14786,N_14673);
or UO_1562 (O_1562,N_14725,N_14854);
xnor UO_1563 (O_1563,N_14566,N_14509);
xnor UO_1564 (O_1564,N_14619,N_14729);
xor UO_1565 (O_1565,N_14969,N_14793);
nand UO_1566 (O_1566,N_14803,N_14907);
nand UO_1567 (O_1567,N_14982,N_14676);
or UO_1568 (O_1568,N_14552,N_14726);
nor UO_1569 (O_1569,N_14538,N_14834);
xnor UO_1570 (O_1570,N_14671,N_14928);
and UO_1571 (O_1571,N_14799,N_14731);
xor UO_1572 (O_1572,N_14878,N_14818);
nand UO_1573 (O_1573,N_14577,N_14558);
or UO_1574 (O_1574,N_14915,N_14759);
xor UO_1575 (O_1575,N_14797,N_14650);
and UO_1576 (O_1576,N_14895,N_14773);
or UO_1577 (O_1577,N_14644,N_14642);
nand UO_1578 (O_1578,N_14502,N_14703);
nor UO_1579 (O_1579,N_14723,N_14603);
nand UO_1580 (O_1580,N_14910,N_14520);
nor UO_1581 (O_1581,N_14963,N_14984);
nor UO_1582 (O_1582,N_14925,N_14633);
or UO_1583 (O_1583,N_14532,N_14673);
nor UO_1584 (O_1584,N_14871,N_14616);
xor UO_1585 (O_1585,N_14571,N_14533);
nor UO_1586 (O_1586,N_14599,N_14913);
nor UO_1587 (O_1587,N_14629,N_14877);
nor UO_1588 (O_1588,N_14861,N_14961);
xnor UO_1589 (O_1589,N_14533,N_14980);
xnor UO_1590 (O_1590,N_14988,N_14818);
nand UO_1591 (O_1591,N_14587,N_14633);
nor UO_1592 (O_1592,N_14591,N_14890);
and UO_1593 (O_1593,N_14832,N_14566);
and UO_1594 (O_1594,N_14933,N_14642);
nor UO_1595 (O_1595,N_14850,N_14971);
or UO_1596 (O_1596,N_14525,N_14711);
xor UO_1597 (O_1597,N_14704,N_14848);
nand UO_1598 (O_1598,N_14697,N_14581);
or UO_1599 (O_1599,N_14850,N_14505);
nor UO_1600 (O_1600,N_14990,N_14721);
nor UO_1601 (O_1601,N_14653,N_14933);
nand UO_1602 (O_1602,N_14976,N_14803);
nor UO_1603 (O_1603,N_14751,N_14571);
and UO_1604 (O_1604,N_14974,N_14962);
nand UO_1605 (O_1605,N_14680,N_14807);
nand UO_1606 (O_1606,N_14719,N_14751);
and UO_1607 (O_1607,N_14592,N_14744);
nor UO_1608 (O_1608,N_14689,N_14730);
and UO_1609 (O_1609,N_14926,N_14936);
nand UO_1610 (O_1610,N_14918,N_14876);
or UO_1611 (O_1611,N_14710,N_14928);
or UO_1612 (O_1612,N_14690,N_14887);
xnor UO_1613 (O_1613,N_14686,N_14598);
and UO_1614 (O_1614,N_14566,N_14909);
nor UO_1615 (O_1615,N_14501,N_14860);
and UO_1616 (O_1616,N_14620,N_14866);
or UO_1617 (O_1617,N_14799,N_14998);
nor UO_1618 (O_1618,N_14685,N_14718);
and UO_1619 (O_1619,N_14698,N_14631);
xnor UO_1620 (O_1620,N_14823,N_14678);
xor UO_1621 (O_1621,N_14567,N_14785);
nor UO_1622 (O_1622,N_14828,N_14605);
xnor UO_1623 (O_1623,N_14635,N_14778);
nor UO_1624 (O_1624,N_14530,N_14591);
nand UO_1625 (O_1625,N_14999,N_14665);
or UO_1626 (O_1626,N_14532,N_14861);
or UO_1627 (O_1627,N_14678,N_14564);
and UO_1628 (O_1628,N_14908,N_14875);
and UO_1629 (O_1629,N_14947,N_14946);
xor UO_1630 (O_1630,N_14581,N_14508);
xnor UO_1631 (O_1631,N_14734,N_14615);
or UO_1632 (O_1632,N_14992,N_14933);
or UO_1633 (O_1633,N_14731,N_14681);
nand UO_1634 (O_1634,N_14945,N_14934);
nand UO_1635 (O_1635,N_14642,N_14975);
and UO_1636 (O_1636,N_14651,N_14779);
or UO_1637 (O_1637,N_14675,N_14832);
nor UO_1638 (O_1638,N_14720,N_14815);
xor UO_1639 (O_1639,N_14964,N_14960);
nand UO_1640 (O_1640,N_14737,N_14756);
and UO_1641 (O_1641,N_14990,N_14957);
or UO_1642 (O_1642,N_14620,N_14718);
or UO_1643 (O_1643,N_14986,N_14597);
nor UO_1644 (O_1644,N_14703,N_14740);
xor UO_1645 (O_1645,N_14825,N_14898);
nor UO_1646 (O_1646,N_14959,N_14591);
xor UO_1647 (O_1647,N_14650,N_14620);
nor UO_1648 (O_1648,N_14633,N_14504);
or UO_1649 (O_1649,N_14946,N_14784);
xor UO_1650 (O_1650,N_14719,N_14712);
xor UO_1651 (O_1651,N_14766,N_14904);
or UO_1652 (O_1652,N_14647,N_14541);
or UO_1653 (O_1653,N_14866,N_14871);
nand UO_1654 (O_1654,N_14888,N_14954);
and UO_1655 (O_1655,N_14622,N_14759);
nor UO_1656 (O_1656,N_14606,N_14796);
and UO_1657 (O_1657,N_14777,N_14920);
and UO_1658 (O_1658,N_14796,N_14933);
xnor UO_1659 (O_1659,N_14792,N_14841);
or UO_1660 (O_1660,N_14598,N_14527);
nor UO_1661 (O_1661,N_14529,N_14815);
and UO_1662 (O_1662,N_14615,N_14991);
or UO_1663 (O_1663,N_14868,N_14889);
xnor UO_1664 (O_1664,N_14975,N_14885);
xnor UO_1665 (O_1665,N_14531,N_14614);
xnor UO_1666 (O_1666,N_14650,N_14993);
xor UO_1667 (O_1667,N_14542,N_14805);
or UO_1668 (O_1668,N_14933,N_14726);
xor UO_1669 (O_1669,N_14946,N_14702);
xor UO_1670 (O_1670,N_14810,N_14701);
and UO_1671 (O_1671,N_14938,N_14984);
xor UO_1672 (O_1672,N_14785,N_14767);
nand UO_1673 (O_1673,N_14703,N_14853);
and UO_1674 (O_1674,N_14608,N_14564);
and UO_1675 (O_1675,N_14805,N_14705);
or UO_1676 (O_1676,N_14812,N_14635);
nor UO_1677 (O_1677,N_14548,N_14909);
or UO_1678 (O_1678,N_14699,N_14565);
xor UO_1679 (O_1679,N_14761,N_14830);
nor UO_1680 (O_1680,N_14996,N_14548);
or UO_1681 (O_1681,N_14836,N_14917);
xnor UO_1682 (O_1682,N_14797,N_14826);
xnor UO_1683 (O_1683,N_14797,N_14561);
nor UO_1684 (O_1684,N_14677,N_14734);
nor UO_1685 (O_1685,N_14827,N_14856);
nor UO_1686 (O_1686,N_14733,N_14665);
and UO_1687 (O_1687,N_14790,N_14966);
nor UO_1688 (O_1688,N_14961,N_14579);
or UO_1689 (O_1689,N_14954,N_14650);
nor UO_1690 (O_1690,N_14576,N_14746);
nor UO_1691 (O_1691,N_14504,N_14570);
nor UO_1692 (O_1692,N_14660,N_14716);
nand UO_1693 (O_1693,N_14766,N_14532);
nor UO_1694 (O_1694,N_14863,N_14919);
nor UO_1695 (O_1695,N_14897,N_14804);
or UO_1696 (O_1696,N_14583,N_14962);
nand UO_1697 (O_1697,N_14741,N_14612);
and UO_1698 (O_1698,N_14624,N_14519);
nor UO_1699 (O_1699,N_14873,N_14589);
and UO_1700 (O_1700,N_14656,N_14996);
and UO_1701 (O_1701,N_14976,N_14580);
or UO_1702 (O_1702,N_14541,N_14893);
nor UO_1703 (O_1703,N_14840,N_14521);
nor UO_1704 (O_1704,N_14644,N_14956);
nor UO_1705 (O_1705,N_14924,N_14725);
or UO_1706 (O_1706,N_14557,N_14511);
and UO_1707 (O_1707,N_14995,N_14557);
or UO_1708 (O_1708,N_14690,N_14502);
or UO_1709 (O_1709,N_14822,N_14632);
xor UO_1710 (O_1710,N_14885,N_14987);
nand UO_1711 (O_1711,N_14865,N_14889);
nor UO_1712 (O_1712,N_14871,N_14666);
nor UO_1713 (O_1713,N_14640,N_14596);
xnor UO_1714 (O_1714,N_14921,N_14594);
or UO_1715 (O_1715,N_14845,N_14740);
or UO_1716 (O_1716,N_14970,N_14651);
nor UO_1717 (O_1717,N_14835,N_14711);
nor UO_1718 (O_1718,N_14517,N_14564);
nand UO_1719 (O_1719,N_14843,N_14781);
xnor UO_1720 (O_1720,N_14706,N_14768);
nor UO_1721 (O_1721,N_14518,N_14598);
nor UO_1722 (O_1722,N_14622,N_14943);
nand UO_1723 (O_1723,N_14840,N_14612);
nor UO_1724 (O_1724,N_14668,N_14797);
nor UO_1725 (O_1725,N_14849,N_14684);
and UO_1726 (O_1726,N_14927,N_14699);
nand UO_1727 (O_1727,N_14529,N_14756);
nor UO_1728 (O_1728,N_14993,N_14523);
xor UO_1729 (O_1729,N_14928,N_14750);
or UO_1730 (O_1730,N_14749,N_14930);
nor UO_1731 (O_1731,N_14688,N_14952);
xor UO_1732 (O_1732,N_14651,N_14901);
xnor UO_1733 (O_1733,N_14702,N_14729);
xor UO_1734 (O_1734,N_14601,N_14831);
and UO_1735 (O_1735,N_14922,N_14617);
and UO_1736 (O_1736,N_14858,N_14709);
or UO_1737 (O_1737,N_14979,N_14687);
and UO_1738 (O_1738,N_14890,N_14561);
xnor UO_1739 (O_1739,N_14691,N_14504);
nor UO_1740 (O_1740,N_14649,N_14654);
or UO_1741 (O_1741,N_14649,N_14930);
xnor UO_1742 (O_1742,N_14632,N_14734);
xor UO_1743 (O_1743,N_14583,N_14789);
or UO_1744 (O_1744,N_14735,N_14777);
xor UO_1745 (O_1745,N_14796,N_14804);
nand UO_1746 (O_1746,N_14796,N_14674);
and UO_1747 (O_1747,N_14532,N_14771);
xnor UO_1748 (O_1748,N_14840,N_14506);
or UO_1749 (O_1749,N_14838,N_14803);
or UO_1750 (O_1750,N_14792,N_14801);
nand UO_1751 (O_1751,N_14991,N_14992);
nand UO_1752 (O_1752,N_14828,N_14944);
xnor UO_1753 (O_1753,N_14633,N_14715);
nand UO_1754 (O_1754,N_14985,N_14789);
and UO_1755 (O_1755,N_14969,N_14742);
nand UO_1756 (O_1756,N_14629,N_14543);
nor UO_1757 (O_1757,N_14506,N_14699);
nand UO_1758 (O_1758,N_14589,N_14716);
or UO_1759 (O_1759,N_14820,N_14661);
nand UO_1760 (O_1760,N_14615,N_14723);
or UO_1761 (O_1761,N_14648,N_14564);
nand UO_1762 (O_1762,N_14534,N_14727);
and UO_1763 (O_1763,N_14598,N_14885);
xnor UO_1764 (O_1764,N_14830,N_14833);
nor UO_1765 (O_1765,N_14589,N_14926);
and UO_1766 (O_1766,N_14829,N_14755);
or UO_1767 (O_1767,N_14766,N_14985);
and UO_1768 (O_1768,N_14702,N_14726);
nand UO_1769 (O_1769,N_14747,N_14762);
xor UO_1770 (O_1770,N_14564,N_14510);
nand UO_1771 (O_1771,N_14529,N_14998);
nand UO_1772 (O_1772,N_14683,N_14674);
and UO_1773 (O_1773,N_14966,N_14607);
nor UO_1774 (O_1774,N_14800,N_14975);
or UO_1775 (O_1775,N_14694,N_14813);
and UO_1776 (O_1776,N_14537,N_14782);
and UO_1777 (O_1777,N_14762,N_14746);
or UO_1778 (O_1778,N_14977,N_14648);
nand UO_1779 (O_1779,N_14617,N_14906);
and UO_1780 (O_1780,N_14712,N_14799);
and UO_1781 (O_1781,N_14768,N_14800);
or UO_1782 (O_1782,N_14640,N_14910);
or UO_1783 (O_1783,N_14763,N_14743);
nand UO_1784 (O_1784,N_14788,N_14821);
xor UO_1785 (O_1785,N_14742,N_14535);
or UO_1786 (O_1786,N_14588,N_14692);
xnor UO_1787 (O_1787,N_14957,N_14681);
xor UO_1788 (O_1788,N_14518,N_14788);
and UO_1789 (O_1789,N_14879,N_14899);
xnor UO_1790 (O_1790,N_14775,N_14664);
or UO_1791 (O_1791,N_14636,N_14635);
xor UO_1792 (O_1792,N_14540,N_14759);
xnor UO_1793 (O_1793,N_14772,N_14809);
nor UO_1794 (O_1794,N_14704,N_14568);
xor UO_1795 (O_1795,N_14936,N_14666);
or UO_1796 (O_1796,N_14982,N_14834);
or UO_1797 (O_1797,N_14574,N_14848);
nor UO_1798 (O_1798,N_14558,N_14894);
and UO_1799 (O_1799,N_14605,N_14612);
and UO_1800 (O_1800,N_14979,N_14763);
or UO_1801 (O_1801,N_14644,N_14527);
nor UO_1802 (O_1802,N_14961,N_14581);
nor UO_1803 (O_1803,N_14838,N_14668);
and UO_1804 (O_1804,N_14999,N_14933);
or UO_1805 (O_1805,N_14915,N_14900);
xnor UO_1806 (O_1806,N_14522,N_14861);
xor UO_1807 (O_1807,N_14736,N_14738);
or UO_1808 (O_1808,N_14932,N_14990);
nand UO_1809 (O_1809,N_14663,N_14825);
nor UO_1810 (O_1810,N_14806,N_14571);
or UO_1811 (O_1811,N_14935,N_14803);
xnor UO_1812 (O_1812,N_14587,N_14806);
nor UO_1813 (O_1813,N_14803,N_14758);
and UO_1814 (O_1814,N_14520,N_14517);
or UO_1815 (O_1815,N_14591,N_14645);
or UO_1816 (O_1816,N_14763,N_14520);
or UO_1817 (O_1817,N_14793,N_14553);
nand UO_1818 (O_1818,N_14691,N_14839);
xnor UO_1819 (O_1819,N_14803,N_14607);
nand UO_1820 (O_1820,N_14780,N_14954);
xnor UO_1821 (O_1821,N_14750,N_14562);
and UO_1822 (O_1822,N_14597,N_14502);
nand UO_1823 (O_1823,N_14506,N_14527);
or UO_1824 (O_1824,N_14875,N_14926);
xor UO_1825 (O_1825,N_14845,N_14623);
nor UO_1826 (O_1826,N_14970,N_14668);
nor UO_1827 (O_1827,N_14939,N_14804);
and UO_1828 (O_1828,N_14686,N_14777);
nand UO_1829 (O_1829,N_14594,N_14537);
nand UO_1830 (O_1830,N_14733,N_14995);
xnor UO_1831 (O_1831,N_14860,N_14577);
xnor UO_1832 (O_1832,N_14552,N_14597);
xnor UO_1833 (O_1833,N_14570,N_14768);
nand UO_1834 (O_1834,N_14951,N_14903);
and UO_1835 (O_1835,N_14902,N_14631);
or UO_1836 (O_1836,N_14584,N_14888);
nand UO_1837 (O_1837,N_14981,N_14700);
or UO_1838 (O_1838,N_14720,N_14762);
nor UO_1839 (O_1839,N_14753,N_14907);
and UO_1840 (O_1840,N_14894,N_14986);
nor UO_1841 (O_1841,N_14770,N_14675);
and UO_1842 (O_1842,N_14785,N_14522);
or UO_1843 (O_1843,N_14874,N_14810);
or UO_1844 (O_1844,N_14768,N_14868);
and UO_1845 (O_1845,N_14661,N_14621);
nand UO_1846 (O_1846,N_14768,N_14653);
or UO_1847 (O_1847,N_14543,N_14954);
or UO_1848 (O_1848,N_14592,N_14952);
and UO_1849 (O_1849,N_14738,N_14983);
xnor UO_1850 (O_1850,N_14735,N_14602);
nand UO_1851 (O_1851,N_14807,N_14982);
nand UO_1852 (O_1852,N_14600,N_14565);
nor UO_1853 (O_1853,N_14522,N_14894);
and UO_1854 (O_1854,N_14566,N_14676);
xor UO_1855 (O_1855,N_14553,N_14506);
and UO_1856 (O_1856,N_14917,N_14856);
and UO_1857 (O_1857,N_14544,N_14615);
xor UO_1858 (O_1858,N_14766,N_14854);
nor UO_1859 (O_1859,N_14777,N_14699);
xnor UO_1860 (O_1860,N_14872,N_14832);
and UO_1861 (O_1861,N_14956,N_14638);
nand UO_1862 (O_1862,N_14637,N_14818);
or UO_1863 (O_1863,N_14715,N_14974);
nor UO_1864 (O_1864,N_14952,N_14806);
xnor UO_1865 (O_1865,N_14751,N_14603);
xor UO_1866 (O_1866,N_14537,N_14875);
and UO_1867 (O_1867,N_14822,N_14529);
xnor UO_1868 (O_1868,N_14583,N_14600);
xor UO_1869 (O_1869,N_14767,N_14798);
or UO_1870 (O_1870,N_14682,N_14676);
and UO_1871 (O_1871,N_14742,N_14939);
and UO_1872 (O_1872,N_14658,N_14743);
nor UO_1873 (O_1873,N_14982,N_14863);
and UO_1874 (O_1874,N_14954,N_14512);
xnor UO_1875 (O_1875,N_14748,N_14822);
or UO_1876 (O_1876,N_14708,N_14957);
nand UO_1877 (O_1877,N_14678,N_14833);
nor UO_1878 (O_1878,N_14641,N_14634);
and UO_1879 (O_1879,N_14640,N_14820);
nor UO_1880 (O_1880,N_14681,N_14507);
nand UO_1881 (O_1881,N_14561,N_14726);
and UO_1882 (O_1882,N_14749,N_14748);
or UO_1883 (O_1883,N_14999,N_14589);
or UO_1884 (O_1884,N_14552,N_14797);
xor UO_1885 (O_1885,N_14844,N_14541);
or UO_1886 (O_1886,N_14663,N_14619);
nand UO_1887 (O_1887,N_14840,N_14518);
and UO_1888 (O_1888,N_14567,N_14990);
nor UO_1889 (O_1889,N_14705,N_14958);
nor UO_1890 (O_1890,N_14859,N_14823);
nand UO_1891 (O_1891,N_14637,N_14754);
or UO_1892 (O_1892,N_14528,N_14712);
nand UO_1893 (O_1893,N_14968,N_14881);
and UO_1894 (O_1894,N_14649,N_14855);
nor UO_1895 (O_1895,N_14528,N_14560);
and UO_1896 (O_1896,N_14664,N_14712);
and UO_1897 (O_1897,N_14774,N_14708);
or UO_1898 (O_1898,N_14638,N_14969);
or UO_1899 (O_1899,N_14787,N_14689);
xnor UO_1900 (O_1900,N_14879,N_14877);
xor UO_1901 (O_1901,N_14568,N_14513);
xor UO_1902 (O_1902,N_14714,N_14924);
or UO_1903 (O_1903,N_14800,N_14981);
or UO_1904 (O_1904,N_14762,N_14816);
nand UO_1905 (O_1905,N_14975,N_14540);
nor UO_1906 (O_1906,N_14727,N_14710);
nand UO_1907 (O_1907,N_14901,N_14840);
nand UO_1908 (O_1908,N_14512,N_14925);
and UO_1909 (O_1909,N_14848,N_14576);
or UO_1910 (O_1910,N_14889,N_14996);
or UO_1911 (O_1911,N_14653,N_14874);
xor UO_1912 (O_1912,N_14862,N_14680);
xnor UO_1913 (O_1913,N_14549,N_14584);
or UO_1914 (O_1914,N_14635,N_14868);
nand UO_1915 (O_1915,N_14687,N_14862);
nor UO_1916 (O_1916,N_14506,N_14728);
xor UO_1917 (O_1917,N_14779,N_14621);
or UO_1918 (O_1918,N_14528,N_14956);
nor UO_1919 (O_1919,N_14878,N_14824);
nor UO_1920 (O_1920,N_14797,N_14680);
or UO_1921 (O_1921,N_14703,N_14757);
and UO_1922 (O_1922,N_14515,N_14648);
nor UO_1923 (O_1923,N_14760,N_14541);
nor UO_1924 (O_1924,N_14725,N_14608);
or UO_1925 (O_1925,N_14958,N_14521);
nand UO_1926 (O_1926,N_14506,N_14755);
or UO_1927 (O_1927,N_14843,N_14561);
and UO_1928 (O_1928,N_14613,N_14709);
nor UO_1929 (O_1929,N_14526,N_14556);
nand UO_1930 (O_1930,N_14709,N_14853);
xnor UO_1931 (O_1931,N_14900,N_14698);
nor UO_1932 (O_1932,N_14939,N_14915);
and UO_1933 (O_1933,N_14966,N_14912);
nand UO_1934 (O_1934,N_14560,N_14845);
and UO_1935 (O_1935,N_14866,N_14887);
nand UO_1936 (O_1936,N_14731,N_14655);
nor UO_1937 (O_1937,N_14772,N_14547);
or UO_1938 (O_1938,N_14846,N_14504);
nor UO_1939 (O_1939,N_14657,N_14781);
nand UO_1940 (O_1940,N_14520,N_14665);
and UO_1941 (O_1941,N_14802,N_14799);
nor UO_1942 (O_1942,N_14994,N_14788);
and UO_1943 (O_1943,N_14716,N_14903);
nor UO_1944 (O_1944,N_14722,N_14813);
nor UO_1945 (O_1945,N_14943,N_14577);
or UO_1946 (O_1946,N_14951,N_14717);
and UO_1947 (O_1947,N_14929,N_14773);
or UO_1948 (O_1948,N_14679,N_14983);
or UO_1949 (O_1949,N_14527,N_14949);
and UO_1950 (O_1950,N_14778,N_14976);
nand UO_1951 (O_1951,N_14598,N_14687);
xor UO_1952 (O_1952,N_14974,N_14889);
and UO_1953 (O_1953,N_14593,N_14554);
nor UO_1954 (O_1954,N_14688,N_14845);
and UO_1955 (O_1955,N_14949,N_14554);
nor UO_1956 (O_1956,N_14653,N_14527);
xnor UO_1957 (O_1957,N_14711,N_14935);
nor UO_1958 (O_1958,N_14536,N_14919);
and UO_1959 (O_1959,N_14620,N_14884);
nand UO_1960 (O_1960,N_14704,N_14577);
and UO_1961 (O_1961,N_14761,N_14867);
or UO_1962 (O_1962,N_14597,N_14810);
nor UO_1963 (O_1963,N_14836,N_14994);
nor UO_1964 (O_1964,N_14578,N_14817);
and UO_1965 (O_1965,N_14803,N_14911);
xor UO_1966 (O_1966,N_14735,N_14579);
nand UO_1967 (O_1967,N_14828,N_14534);
xnor UO_1968 (O_1968,N_14823,N_14659);
xnor UO_1969 (O_1969,N_14550,N_14766);
and UO_1970 (O_1970,N_14860,N_14519);
nor UO_1971 (O_1971,N_14644,N_14891);
nor UO_1972 (O_1972,N_14682,N_14658);
or UO_1973 (O_1973,N_14666,N_14865);
or UO_1974 (O_1974,N_14565,N_14945);
nand UO_1975 (O_1975,N_14526,N_14812);
nor UO_1976 (O_1976,N_14665,N_14993);
nand UO_1977 (O_1977,N_14541,N_14870);
nor UO_1978 (O_1978,N_14553,N_14887);
or UO_1979 (O_1979,N_14909,N_14890);
or UO_1980 (O_1980,N_14815,N_14722);
and UO_1981 (O_1981,N_14503,N_14522);
xor UO_1982 (O_1982,N_14523,N_14856);
xor UO_1983 (O_1983,N_14559,N_14529);
nor UO_1984 (O_1984,N_14724,N_14736);
nand UO_1985 (O_1985,N_14795,N_14648);
xor UO_1986 (O_1986,N_14962,N_14922);
and UO_1987 (O_1987,N_14665,N_14679);
xor UO_1988 (O_1988,N_14546,N_14521);
and UO_1989 (O_1989,N_14873,N_14974);
nor UO_1990 (O_1990,N_14862,N_14900);
xor UO_1991 (O_1991,N_14859,N_14711);
or UO_1992 (O_1992,N_14562,N_14689);
xor UO_1993 (O_1993,N_14652,N_14931);
xor UO_1994 (O_1994,N_14669,N_14844);
or UO_1995 (O_1995,N_14519,N_14741);
xnor UO_1996 (O_1996,N_14782,N_14661);
or UO_1997 (O_1997,N_14551,N_14617);
nand UO_1998 (O_1998,N_14860,N_14955);
nor UO_1999 (O_1999,N_14536,N_14968);
endmodule