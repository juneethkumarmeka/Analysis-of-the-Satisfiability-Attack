module basic_1000_10000_1500_20_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_619,In_766);
and U1 (N_1,In_160,In_471);
xnor U2 (N_2,In_565,In_374);
or U3 (N_3,In_15,In_352);
nor U4 (N_4,In_146,In_249);
nand U5 (N_5,In_654,In_897);
xor U6 (N_6,In_258,In_782);
and U7 (N_7,In_48,In_923);
xnor U8 (N_8,In_981,In_450);
nor U9 (N_9,In_446,In_926);
nand U10 (N_10,In_20,In_773);
xor U11 (N_11,In_898,In_141);
and U12 (N_12,In_761,In_608);
nor U13 (N_13,In_78,In_667);
or U14 (N_14,In_128,In_58);
nor U15 (N_15,In_218,In_712);
xnor U16 (N_16,In_193,In_470);
xnor U17 (N_17,In_809,In_340);
xor U18 (N_18,In_56,In_640);
nand U19 (N_19,In_703,In_333);
and U20 (N_20,In_321,In_747);
or U21 (N_21,In_407,In_704);
nand U22 (N_22,In_464,In_267);
nand U23 (N_23,In_757,In_969);
xor U24 (N_24,In_617,In_400);
nor U25 (N_25,In_403,In_482);
nor U26 (N_26,In_103,In_625);
nand U27 (N_27,In_561,In_974);
or U28 (N_28,In_299,In_736);
nand U29 (N_29,In_768,In_236);
xor U30 (N_30,In_404,In_716);
nor U31 (N_31,In_986,In_723);
xor U32 (N_32,In_551,In_247);
xnor U33 (N_33,In_595,In_724);
xor U34 (N_34,In_882,In_887);
xnor U35 (N_35,In_116,In_980);
nor U36 (N_36,In_652,In_602);
nand U37 (N_37,In_270,In_35);
and U38 (N_38,In_324,In_307);
and U39 (N_39,In_246,In_136);
nand U40 (N_40,In_740,In_499);
or U41 (N_41,In_341,In_455);
xnor U42 (N_42,In_540,In_351);
xor U43 (N_43,In_938,In_702);
xnor U44 (N_44,In_901,In_566);
and U45 (N_45,In_947,In_888);
or U46 (N_46,In_548,In_301);
nor U47 (N_47,In_730,In_275);
and U48 (N_48,In_408,In_693);
xor U49 (N_49,In_84,In_37);
nand U50 (N_50,In_728,In_607);
nor U51 (N_51,In_623,In_738);
nor U52 (N_52,In_239,In_253);
nand U53 (N_53,In_826,In_687);
xnor U54 (N_54,In_90,In_706);
or U55 (N_55,In_711,In_401);
and U56 (N_56,In_588,In_658);
xnor U57 (N_57,In_143,In_131);
or U58 (N_58,In_624,In_461);
nor U59 (N_59,In_422,In_643);
xor U60 (N_60,In_835,In_573);
or U61 (N_61,In_286,In_528);
nor U62 (N_62,In_363,In_362);
and U63 (N_63,In_469,In_463);
xor U64 (N_64,In_390,In_771);
or U65 (N_65,In_281,In_448);
nand U66 (N_66,In_346,In_223);
or U67 (N_67,In_361,In_705);
nor U68 (N_68,In_159,In_36);
or U69 (N_69,In_937,In_525);
and U70 (N_70,In_631,In_170);
or U71 (N_71,In_389,In_88);
or U72 (N_72,In_952,In_251);
and U73 (N_73,In_457,In_715);
and U74 (N_74,In_932,In_296);
xor U75 (N_75,In_857,In_801);
xnor U76 (N_76,In_265,In_543);
and U77 (N_77,In_402,In_886);
nor U78 (N_78,In_38,In_676);
nand U79 (N_79,In_961,In_550);
nor U80 (N_80,In_600,In_793);
nand U81 (N_81,In_685,In_927);
and U82 (N_82,In_443,In_43);
nand U83 (N_83,In_939,In_847);
or U84 (N_84,In_962,In_661);
or U85 (N_85,In_774,In_506);
nor U86 (N_86,In_813,In_65);
xnor U87 (N_87,In_649,In_752);
or U88 (N_88,In_368,In_902);
nor U89 (N_89,In_812,In_183);
xnor U90 (N_90,In_612,In_254);
or U91 (N_91,In_486,In_61);
or U92 (N_92,In_266,In_549);
or U93 (N_93,In_130,In_171);
nor U94 (N_94,In_669,In_154);
xnor U95 (N_95,In_46,In_903);
xnor U96 (N_96,In_230,In_673);
xor U97 (N_97,In_531,In_745);
and U98 (N_98,In_398,In_783);
nand U99 (N_99,In_713,In_929);
nor U100 (N_100,In_741,In_49);
and U101 (N_101,In_794,In_489);
or U102 (N_102,In_66,In_632);
nand U103 (N_103,In_827,In_541);
nand U104 (N_104,In_849,In_662);
xnor U105 (N_105,In_495,In_164);
and U106 (N_106,In_344,In_204);
nand U107 (N_107,In_118,In_92);
xnor U108 (N_108,In_996,In_984);
xnor U109 (N_109,In_411,In_999);
xnor U110 (N_110,In_910,In_796);
nand U111 (N_111,In_399,In_257);
xnor U112 (N_112,In_293,In_726);
nor U113 (N_113,In_315,In_206);
xnor U114 (N_114,In_339,In_964);
and U115 (N_115,In_570,In_298);
and U116 (N_116,In_221,In_795);
and U117 (N_117,In_731,In_587);
nand U118 (N_118,In_988,In_921);
and U119 (N_119,In_678,In_472);
nand U120 (N_120,In_831,In_934);
or U121 (N_121,In_904,In_563);
nand U122 (N_122,In_663,In_16);
nand U123 (N_123,In_1,In_209);
and U124 (N_124,In_682,In_900);
xor U125 (N_125,In_231,In_945);
nand U126 (N_126,In_14,In_606);
xor U127 (N_127,In_837,In_539);
nand U128 (N_128,In_553,In_529);
xnor U129 (N_129,In_176,In_310);
or U130 (N_130,In_917,In_144);
or U131 (N_131,In_918,In_511);
nor U132 (N_132,In_824,In_383);
or U133 (N_133,In_329,In_957);
nand U134 (N_134,In_879,In_4);
nand U135 (N_135,In_274,In_593);
nand U136 (N_136,In_271,In_765);
xnor U137 (N_137,In_727,In_191);
xor U138 (N_138,In_334,In_775);
nand U139 (N_139,In_198,In_153);
or U140 (N_140,In_859,In_107);
nor U141 (N_141,In_852,In_376);
or U142 (N_142,In_839,In_873);
or U143 (N_143,In_364,In_180);
nand U144 (N_144,In_598,In_101);
and U145 (N_145,In_454,In_718);
nand U146 (N_146,In_83,In_323);
nor U147 (N_147,In_884,In_425);
nor U148 (N_148,In_392,In_313);
nand U149 (N_149,In_821,In_535);
and U150 (N_150,In_855,In_650);
nand U151 (N_151,In_743,In_876);
and U152 (N_152,In_629,In_93);
or U153 (N_153,In_559,In_759);
and U154 (N_154,In_211,In_203);
and U155 (N_155,In_729,In_201);
nand U156 (N_156,In_54,In_790);
nand U157 (N_157,In_262,In_9);
or U158 (N_158,In_358,In_73);
nand U159 (N_159,In_686,In_998);
xnor U160 (N_160,In_8,In_21);
or U161 (N_161,In_259,In_737);
nor U162 (N_162,In_708,In_544);
xor U163 (N_163,In_30,In_815);
nor U164 (N_164,In_19,In_263);
nor U165 (N_165,In_322,In_468);
nand U166 (N_166,In_990,In_256);
or U167 (N_167,In_758,In_44);
nor U168 (N_168,In_694,In_520);
nand U169 (N_169,In_615,In_50);
or U170 (N_170,In_175,In_893);
xnor U171 (N_171,In_139,In_200);
or U172 (N_172,In_115,In_336);
and U173 (N_173,In_91,In_577);
nor U174 (N_174,In_722,In_142);
nand U175 (N_175,In_555,In_944);
and U176 (N_176,In_992,In_237);
nor U177 (N_177,In_224,In_935);
and U178 (N_178,In_772,In_347);
nand U179 (N_179,In_972,In_72);
xor U180 (N_180,In_830,In_997);
nor U181 (N_181,In_290,In_763);
nor U182 (N_182,In_121,In_502);
xnor U183 (N_183,In_627,In_621);
nor U184 (N_184,In_844,In_907);
or U185 (N_185,In_210,In_445);
and U186 (N_186,In_696,In_395);
nand U187 (N_187,In_371,In_149);
and U188 (N_188,In_355,In_785);
xor U189 (N_189,In_189,In_199);
nand U190 (N_190,In_172,In_622);
xor U191 (N_191,In_314,In_585);
nor U192 (N_192,In_516,In_80);
or U193 (N_193,In_94,In_594);
nor U194 (N_194,In_449,In_488);
or U195 (N_195,In_697,In_556);
and U196 (N_196,In_409,In_165);
xnor U197 (N_197,In_42,In_382);
and U198 (N_198,In_490,In_74);
nand U199 (N_199,In_441,In_76);
xnor U200 (N_200,In_151,In_332);
nor U201 (N_201,In_574,In_523);
or U202 (N_202,In_280,In_357);
nand U203 (N_203,In_820,In_637);
and U204 (N_204,In_484,In_848);
and U205 (N_205,In_861,In_657);
nor U206 (N_206,In_803,In_393);
nand U207 (N_207,In_503,In_811);
nand U208 (N_208,In_987,In_660);
nand U209 (N_209,In_432,In_960);
nor U210 (N_210,In_959,In_895);
or U211 (N_211,In_973,In_672);
nor U212 (N_212,In_985,In_110);
nand U213 (N_213,In_438,In_905);
xor U214 (N_214,In_581,In_39);
nor U215 (N_215,In_147,In_965);
or U216 (N_216,In_452,In_851);
and U217 (N_217,In_633,In_699);
and U218 (N_218,In_791,In_328);
nand U219 (N_219,In_109,In_381);
or U220 (N_220,In_955,In_487);
or U221 (N_221,In_108,In_122);
nand U222 (N_222,In_580,In_519);
nor U223 (N_223,In_527,In_386);
xor U224 (N_224,In_473,In_348);
nor U225 (N_225,In_991,In_806);
nand U226 (N_226,In_406,In_899);
and U227 (N_227,In_546,In_68);
xor U228 (N_228,In_681,In_721);
xor U229 (N_229,In_679,In_132);
nand U230 (N_230,In_430,In_156);
xnor U231 (N_231,In_916,In_860);
nand U232 (N_232,In_264,In_426);
nand U233 (N_233,In_639,In_651);
and U234 (N_234,In_750,In_890);
and U235 (N_235,In_828,In_22);
nor U236 (N_236,In_181,In_767);
nand U237 (N_237,In_162,In_435);
or U238 (N_238,In_659,In_804);
and U239 (N_239,In_509,In_97);
nor U240 (N_240,In_338,In_305);
xor U241 (N_241,In_628,In_808);
nor U242 (N_242,In_294,In_459);
xor U243 (N_243,In_825,In_885);
or U244 (N_244,In_417,In_196);
xnor U245 (N_245,In_5,In_252);
xor U246 (N_246,In_579,In_925);
or U247 (N_247,In_913,In_863);
and U248 (N_248,In_453,In_946);
or U249 (N_249,In_308,In_883);
nand U250 (N_250,In_787,In_248);
xnor U251 (N_251,In_276,In_232);
and U252 (N_252,In_554,In_560);
xor U253 (N_253,In_45,In_359);
nand U254 (N_254,In_356,In_474);
nor U255 (N_255,In_228,In_725);
or U256 (N_256,In_497,In_919);
and U257 (N_257,In_480,In_735);
xnor U258 (N_258,In_123,In_647);
and U259 (N_259,In_982,In_250);
nor U260 (N_260,In_993,In_942);
nand U261 (N_261,In_148,In_134);
nand U262 (N_262,In_779,In_508);
nand U263 (N_263,In_971,In_13);
or U264 (N_264,In_412,In_547);
or U265 (N_265,In_877,In_420);
nor U266 (N_266,In_467,In_292);
nor U267 (N_267,In_312,In_190);
nand U268 (N_268,In_219,In_304);
nand U269 (N_269,In_373,In_963);
xnor U270 (N_270,In_756,In_89);
or U271 (N_271,In_238,In_194);
nor U272 (N_272,In_610,In_832);
or U273 (N_273,In_800,In_261);
nor U274 (N_274,In_379,In_451);
nand U275 (N_275,In_753,In_397);
nor U276 (N_276,In_47,In_868);
xor U277 (N_277,In_272,In_911);
nor U278 (N_278,In_405,In_7);
nor U279 (N_279,In_739,In_309);
xnor U280 (N_280,In_24,In_291);
or U281 (N_281,In_940,In_227);
xor U282 (N_282,In_157,In_57);
and U283 (N_283,In_616,In_853);
xnor U284 (N_284,In_104,In_842);
nand U285 (N_285,In_184,In_846);
and U286 (N_286,In_119,In_127);
or U287 (N_287,In_179,In_688);
or U288 (N_288,In_229,In_133);
xnor U289 (N_289,In_604,In_507);
and U290 (N_290,In_700,In_319);
or U291 (N_291,In_465,In_102);
and U292 (N_292,In_709,In_609);
nand U293 (N_293,In_605,In_460);
nor U294 (N_294,In_17,In_513);
nor U295 (N_295,In_311,In_233);
nand U296 (N_296,In_552,In_576);
nor U297 (N_297,In_367,In_349);
xnor U298 (N_298,In_135,In_225);
and U299 (N_299,In_675,In_86);
or U300 (N_300,In_777,In_11);
xnor U301 (N_301,In_222,In_977);
nand U302 (N_302,In_245,In_216);
and U303 (N_303,In_754,In_538);
xor U304 (N_304,In_350,In_444);
or U305 (N_305,In_477,In_591);
and U306 (N_306,In_335,In_456);
and U307 (N_307,In_833,In_418);
nor U308 (N_308,In_592,In_424);
or U309 (N_309,In_26,In_79);
xnor U310 (N_310,In_207,In_522);
nand U311 (N_311,In_394,In_896);
nor U312 (N_312,In_684,In_603);
or U313 (N_313,In_933,In_427);
or U314 (N_314,In_958,In_129);
xnor U315 (N_315,In_192,In_173);
or U316 (N_316,In_53,In_85);
and U317 (N_317,In_789,In_187);
nor U318 (N_318,In_174,In_70);
nor U319 (N_319,In_431,In_967);
nor U320 (N_320,In_840,In_205);
nand U321 (N_321,In_370,In_569);
nand U322 (N_322,In_421,In_572);
and U323 (N_323,In_995,In_596);
nand U324 (N_324,In_922,In_494);
nor U325 (N_325,In_515,In_99);
xor U326 (N_326,In_354,In_776);
nor U327 (N_327,In_82,In_642);
and U328 (N_328,In_504,In_114);
and U329 (N_329,In_491,In_226);
nor U330 (N_330,In_664,In_778);
nor U331 (N_331,In_575,In_870);
or U332 (N_332,In_843,In_645);
and U333 (N_333,In_111,In_524);
nor U334 (N_334,In_760,In_648);
nand U335 (N_335,In_260,In_345);
nor U336 (N_336,In_871,In_337);
xor U337 (N_337,In_683,In_646);
nor U338 (N_338,In_814,In_571);
and U339 (N_339,In_668,In_924);
or U340 (N_340,In_158,In_439);
and U341 (N_341,In_268,In_691);
nor U342 (N_342,In_822,In_287);
nand U343 (N_343,In_55,In_186);
or U344 (N_344,In_854,In_161);
or U345 (N_345,In_327,In_695);
nor U346 (N_346,In_816,In_442);
xnor U347 (N_347,In_665,In_568);
nand U348 (N_348,In_909,In_719);
and U349 (N_349,In_564,In_126);
nand U350 (N_350,In_113,In_866);
nor U351 (N_351,In_105,In_163);
xnor U352 (N_352,In_720,In_889);
nor U353 (N_353,In_792,In_786);
or U354 (N_354,In_701,In_188);
nand U355 (N_355,In_976,In_951);
nand U356 (N_356,In_865,In_968);
or U357 (N_357,In_920,In_318);
and U358 (N_358,In_862,In_689);
nand U359 (N_359,In_277,In_87);
and U360 (N_360,In_214,In_557);
xnor U361 (N_361,In_948,In_755);
or U362 (N_362,In_823,In_98);
nand U363 (N_363,In_380,In_295);
or U364 (N_364,In_77,In_762);
or U365 (N_365,In_466,In_635);
nor U366 (N_366,In_912,In_213);
and U367 (N_367,In_278,In_447);
or U368 (N_368,In_655,In_69);
xnor U369 (N_369,In_433,In_51);
or U370 (N_370,In_75,In_117);
or U371 (N_371,In_875,In_353);
nor U372 (N_372,In_428,In_597);
xnor U373 (N_373,In_40,In_152);
nand U374 (N_374,In_975,In_838);
nand U375 (N_375,In_64,In_137);
xor U376 (N_376,In_878,In_235);
xnor U377 (N_377,In_273,In_63);
xor U378 (N_378,In_33,In_526);
and U379 (N_379,In_545,In_493);
or U380 (N_380,In_978,In_67);
nor U381 (N_381,In_666,In_562);
and U382 (N_382,In_242,In_644);
and U383 (N_383,In_2,In_611);
or U384 (N_384,In_734,In_498);
and U385 (N_385,In_279,In_241);
xor U386 (N_386,In_798,In_185);
and U387 (N_387,In_140,In_744);
nand U388 (N_388,In_894,In_748);
nor U389 (N_389,In_377,In_505);
and U390 (N_390,In_601,In_169);
nand U391 (N_391,In_285,In_970);
xor U392 (N_392,In_950,In_989);
nand U393 (N_393,In_620,In_100);
or U394 (N_394,In_936,In_521);
and U395 (N_395,In_536,In_841);
xnor U396 (N_396,In_692,In_582);
nor U397 (N_397,In_829,In_440);
and U398 (N_398,In_306,In_375);
nor U399 (N_399,In_300,In_717);
nor U400 (N_400,In_81,In_71);
nor U401 (N_401,In_856,In_510);
nand U402 (N_402,In_630,In_95);
xnor U403 (N_403,In_698,In_388);
and U404 (N_404,In_636,In_6);
xor U405 (N_405,In_369,In_653);
and U406 (N_406,In_805,In_208);
and U407 (N_407,In_60,In_915);
and U408 (N_408,In_928,In_872);
or U409 (N_409,In_881,In_387);
xnor U410 (N_410,In_864,In_120);
xnor U411 (N_411,In_302,In_365);
xnor U412 (N_412,In_671,In_770);
and U413 (N_413,In_289,In_462);
nand U414 (N_414,In_819,In_514);
xnor U415 (N_415,In_217,In_429);
xor U416 (N_416,In_414,In_500);
xor U417 (N_417,In_195,In_496);
and U418 (N_418,In_867,In_780);
and U419 (N_419,In_634,In_331);
or U420 (N_420,In_733,In_413);
xnor U421 (N_421,In_415,In_416);
nand U422 (N_422,In_956,In_537);
xnor U423 (N_423,In_283,In_583);
xnor U424 (N_424,In_168,In_943);
or U425 (N_425,In_255,In_802);
xnor U426 (N_426,In_360,In_0);
or U427 (N_427,In_475,In_28);
nand U428 (N_428,In_3,In_155);
nand U429 (N_429,In_618,In_680);
or U430 (N_430,In_690,In_234);
nor U431 (N_431,In_385,In_641);
nor U432 (N_432,In_732,In_96);
and U433 (N_433,In_481,In_124);
xnor U434 (N_434,In_892,In_810);
or U435 (N_435,In_807,In_742);
nand U436 (N_436,In_434,In_530);
nand U437 (N_437,In_638,In_994);
nor U438 (N_438,In_626,In_836);
nand U439 (N_439,In_613,In_182);
nand U440 (N_440,In_614,In_784);
or U441 (N_441,In_436,In_41);
and U442 (N_442,In_674,In_150);
nand U443 (N_443,In_850,In_590);
nand U444 (N_444,In_845,In_501);
or U445 (N_445,In_177,In_342);
and U446 (N_446,In_542,In_29);
and U447 (N_447,In_586,In_532);
and U448 (N_448,In_458,In_656);
xnor U449 (N_449,In_112,In_18);
and U450 (N_450,In_512,In_584);
or U451 (N_451,In_781,In_818);
xor U452 (N_452,In_930,In_138);
xnor U453 (N_453,In_518,In_908);
xnor U454 (N_454,In_599,In_297);
nand U455 (N_455,In_166,In_954);
xnor U456 (N_456,In_23,In_479);
xor U457 (N_457,In_410,In_269);
or U458 (N_458,In_534,In_533);
or U459 (N_459,In_914,In_372);
xnor U460 (N_460,In_880,In_303);
xnor U461 (N_461,In_817,In_320);
nor U462 (N_462,In_284,In_769);
or U463 (N_463,In_423,In_492);
and U464 (N_464,In_419,In_167);
xor U465 (N_465,In_343,In_558);
and U466 (N_466,In_483,In_437);
nand U467 (N_467,In_378,In_517);
and U468 (N_468,In_966,In_125);
and U469 (N_469,In_59,In_197);
xnor U470 (N_470,In_25,In_788);
nand U471 (N_471,In_670,In_983);
or U472 (N_472,In_212,In_891);
nor U473 (N_473,In_244,In_941);
and U474 (N_474,In_240,In_858);
or U475 (N_475,In_931,In_31);
nor U476 (N_476,In_476,In_62);
or U477 (N_477,In_797,In_485);
xnor U478 (N_478,In_202,In_567);
nand U479 (N_479,In_330,In_317);
nor U480 (N_480,In_325,In_288);
and U481 (N_481,In_834,In_799);
xnor U482 (N_482,In_178,In_906);
or U483 (N_483,In_396,In_52);
and U484 (N_484,In_746,In_145);
xor U485 (N_485,In_220,In_243);
xor U486 (N_486,In_10,In_32);
xor U487 (N_487,In_749,In_751);
nor U488 (N_488,In_874,In_326);
and U489 (N_489,In_366,In_384);
nand U490 (N_490,In_316,In_953);
nand U491 (N_491,In_949,In_215);
and U492 (N_492,In_707,In_391);
nor U493 (N_493,In_869,In_27);
xnor U494 (N_494,In_677,In_714);
nor U495 (N_495,In_979,In_478);
xnor U496 (N_496,In_34,In_589);
or U497 (N_497,In_764,In_578);
xnor U498 (N_498,In_106,In_710);
and U499 (N_499,In_282,In_12);
and U500 (N_500,N_352,N_170);
nand U501 (N_501,N_39,N_432);
nand U502 (N_502,N_327,N_302);
and U503 (N_503,N_349,N_294);
xor U504 (N_504,N_128,N_47);
and U505 (N_505,N_26,N_472);
nor U506 (N_506,N_225,N_133);
xnor U507 (N_507,N_493,N_371);
and U508 (N_508,N_151,N_42);
and U509 (N_509,N_445,N_2);
xnor U510 (N_510,N_312,N_162);
xor U511 (N_511,N_470,N_89);
and U512 (N_512,N_43,N_118);
nand U513 (N_513,N_298,N_131);
and U514 (N_514,N_33,N_319);
nand U515 (N_515,N_449,N_35);
nand U516 (N_516,N_183,N_280);
or U517 (N_517,N_215,N_172);
or U518 (N_518,N_343,N_85);
xor U519 (N_519,N_50,N_479);
nand U520 (N_520,N_301,N_482);
nand U521 (N_521,N_264,N_334);
or U522 (N_522,N_153,N_20);
xnor U523 (N_523,N_290,N_211);
nand U524 (N_524,N_93,N_465);
nor U525 (N_525,N_72,N_221);
and U526 (N_526,N_333,N_195);
or U527 (N_527,N_487,N_263);
nand U528 (N_528,N_339,N_483);
and U529 (N_529,N_37,N_149);
or U530 (N_530,N_469,N_441);
nor U531 (N_531,N_423,N_431);
and U532 (N_532,N_88,N_275);
nand U533 (N_533,N_176,N_255);
xor U534 (N_534,N_383,N_391);
nor U535 (N_535,N_321,N_359);
and U536 (N_536,N_428,N_1);
and U537 (N_537,N_148,N_242);
or U538 (N_538,N_116,N_323);
nor U539 (N_539,N_184,N_58);
nor U540 (N_540,N_273,N_351);
or U541 (N_541,N_135,N_406);
or U542 (N_542,N_364,N_457);
and U543 (N_543,N_220,N_227);
nand U544 (N_544,N_87,N_120);
nand U545 (N_545,N_99,N_387);
or U546 (N_546,N_380,N_397);
and U547 (N_547,N_475,N_295);
nor U548 (N_548,N_353,N_7);
nor U549 (N_549,N_198,N_59);
nor U550 (N_550,N_234,N_159);
nor U551 (N_551,N_408,N_123);
nor U552 (N_552,N_157,N_17);
nor U553 (N_553,N_212,N_67);
nor U554 (N_554,N_163,N_154);
nand U555 (N_555,N_464,N_287);
nor U556 (N_556,N_139,N_365);
nand U557 (N_557,N_25,N_9);
or U558 (N_558,N_3,N_420);
xor U559 (N_559,N_247,N_15);
and U560 (N_560,N_16,N_21);
nor U561 (N_561,N_106,N_223);
xnor U562 (N_562,N_164,N_55);
nand U563 (N_563,N_488,N_285);
nand U564 (N_564,N_324,N_245);
and U565 (N_565,N_138,N_372);
nor U566 (N_566,N_65,N_354);
or U567 (N_567,N_54,N_370);
xor U568 (N_568,N_405,N_100);
nand U569 (N_569,N_476,N_186);
nor U570 (N_570,N_373,N_494);
xor U571 (N_571,N_474,N_167);
nand U572 (N_572,N_330,N_222);
xnor U573 (N_573,N_450,N_369);
or U574 (N_574,N_291,N_248);
nor U575 (N_575,N_80,N_442);
or U576 (N_576,N_219,N_256);
or U577 (N_577,N_288,N_269);
nand U578 (N_578,N_105,N_393);
nand U579 (N_579,N_68,N_262);
and U580 (N_580,N_4,N_165);
nand U581 (N_581,N_341,N_461);
and U582 (N_582,N_272,N_188);
and U583 (N_583,N_376,N_56);
and U584 (N_584,N_274,N_90);
and U585 (N_585,N_62,N_398);
and U586 (N_586,N_180,N_171);
xnor U587 (N_587,N_30,N_158);
or U588 (N_588,N_458,N_95);
or U589 (N_589,N_433,N_10);
xor U590 (N_590,N_467,N_161);
nor U591 (N_591,N_187,N_111);
nor U592 (N_592,N_96,N_127);
nand U593 (N_593,N_297,N_155);
nand U594 (N_594,N_246,N_218);
nor U595 (N_595,N_388,N_283);
nor U596 (N_596,N_70,N_348);
or U597 (N_597,N_236,N_207);
xor U598 (N_598,N_51,N_407);
xor U599 (N_599,N_326,N_103);
nand U600 (N_600,N_11,N_451);
nor U601 (N_601,N_12,N_205);
nand U602 (N_602,N_136,N_377);
or U603 (N_603,N_328,N_210);
xor U604 (N_604,N_214,N_230);
xnor U605 (N_605,N_232,N_454);
and U606 (N_606,N_202,N_434);
nand U607 (N_607,N_41,N_249);
nor U608 (N_608,N_110,N_299);
or U609 (N_609,N_23,N_145);
and U610 (N_610,N_94,N_335);
and U611 (N_611,N_122,N_32);
nand U612 (N_612,N_378,N_278);
or U613 (N_613,N_84,N_224);
or U614 (N_614,N_481,N_189);
or U615 (N_615,N_453,N_484);
nand U616 (N_616,N_243,N_76);
nor U617 (N_617,N_238,N_115);
and U618 (N_618,N_462,N_395);
and U619 (N_619,N_71,N_430);
or U620 (N_620,N_261,N_347);
nand U621 (N_621,N_60,N_24);
and U622 (N_622,N_424,N_217);
and U623 (N_623,N_208,N_109);
or U624 (N_624,N_417,N_258);
and U625 (N_625,N_322,N_440);
nand U626 (N_626,N_473,N_66);
and U627 (N_627,N_315,N_251);
nand U628 (N_628,N_44,N_429);
nand U629 (N_629,N_310,N_240);
nand U630 (N_630,N_426,N_46);
nor U631 (N_631,N_413,N_300);
nor U632 (N_632,N_156,N_412);
nand U633 (N_633,N_201,N_485);
and U634 (N_634,N_314,N_141);
nor U635 (N_635,N_284,N_5);
nor U636 (N_636,N_69,N_411);
or U637 (N_637,N_38,N_196);
xnor U638 (N_638,N_75,N_182);
nor U639 (N_639,N_0,N_265);
and U640 (N_640,N_229,N_181);
nor U641 (N_641,N_308,N_382);
xnor U642 (N_642,N_346,N_190);
or U643 (N_643,N_204,N_112);
or U644 (N_644,N_98,N_193);
nor U645 (N_645,N_194,N_259);
or U646 (N_646,N_400,N_244);
or U647 (N_647,N_92,N_82);
and U648 (N_648,N_277,N_206);
nand U649 (N_649,N_268,N_375);
nand U650 (N_650,N_356,N_331);
nor U651 (N_651,N_126,N_471);
nand U652 (N_652,N_73,N_40);
nand U653 (N_653,N_480,N_418);
and U654 (N_654,N_266,N_425);
nand U655 (N_655,N_22,N_306);
and U656 (N_656,N_14,N_409);
nor U657 (N_657,N_403,N_228);
nor U658 (N_658,N_468,N_124);
or U659 (N_659,N_402,N_421);
nor U660 (N_660,N_125,N_61);
xnor U661 (N_661,N_29,N_366);
and U662 (N_662,N_355,N_137);
nor U663 (N_663,N_448,N_390);
or U664 (N_664,N_6,N_279);
nand U665 (N_665,N_404,N_152);
nor U666 (N_666,N_410,N_45);
nor U667 (N_667,N_27,N_394);
nor U668 (N_668,N_367,N_419);
xor U669 (N_669,N_199,N_174);
and U670 (N_670,N_197,N_19);
and U671 (N_671,N_117,N_8);
nand U672 (N_672,N_337,N_491);
or U673 (N_673,N_363,N_267);
and U674 (N_674,N_130,N_399);
and U675 (N_675,N_233,N_178);
nor U676 (N_676,N_177,N_316);
nor U677 (N_677,N_231,N_271);
xnor U678 (N_678,N_140,N_160);
nand U679 (N_679,N_86,N_307);
xnor U680 (N_680,N_499,N_336);
or U681 (N_681,N_325,N_144);
or U682 (N_682,N_358,N_114);
nand U683 (N_683,N_313,N_385);
xor U684 (N_684,N_345,N_466);
or U685 (N_685,N_292,N_340);
xor U686 (N_686,N_303,N_304);
xnor U687 (N_687,N_386,N_374);
nand U688 (N_688,N_81,N_150);
xor U689 (N_689,N_460,N_477);
nand U690 (N_690,N_250,N_147);
nor U691 (N_691,N_260,N_381);
or U692 (N_692,N_83,N_132);
nor U693 (N_693,N_446,N_191);
and U694 (N_694,N_185,N_209);
xnor U695 (N_695,N_36,N_142);
nand U696 (N_696,N_63,N_452);
or U697 (N_697,N_309,N_57);
nand U698 (N_698,N_253,N_166);
and U699 (N_699,N_79,N_497);
nor U700 (N_700,N_252,N_362);
nand U701 (N_701,N_134,N_257);
xnor U702 (N_702,N_13,N_401);
nand U703 (N_703,N_329,N_447);
xnor U704 (N_704,N_379,N_49);
nand U705 (N_705,N_270,N_490);
and U706 (N_706,N_357,N_179);
and U707 (N_707,N_289,N_192);
nand U708 (N_708,N_361,N_226);
nand U709 (N_709,N_108,N_318);
xor U710 (N_710,N_350,N_443);
nand U711 (N_711,N_455,N_113);
xor U712 (N_712,N_239,N_444);
nand U713 (N_713,N_296,N_344);
nor U714 (N_714,N_101,N_241);
or U715 (N_715,N_414,N_200);
or U716 (N_716,N_478,N_368);
xnor U717 (N_717,N_64,N_456);
and U718 (N_718,N_305,N_495);
xnor U719 (N_719,N_168,N_435);
xnor U720 (N_720,N_175,N_416);
or U721 (N_721,N_52,N_74);
nand U722 (N_722,N_18,N_389);
or U723 (N_723,N_496,N_463);
and U724 (N_724,N_415,N_34);
xor U725 (N_725,N_119,N_489);
nand U726 (N_726,N_213,N_286);
nand U727 (N_727,N_28,N_360);
or U728 (N_728,N_173,N_48);
nor U729 (N_729,N_143,N_78);
or U730 (N_730,N_129,N_91);
xor U731 (N_731,N_498,N_169);
nor U732 (N_732,N_427,N_254);
xnor U733 (N_733,N_439,N_203);
and U734 (N_734,N_492,N_282);
xnor U735 (N_735,N_281,N_422);
nor U736 (N_736,N_216,N_342);
nand U737 (N_737,N_31,N_235);
and U738 (N_738,N_438,N_311);
xnor U739 (N_739,N_121,N_384);
or U740 (N_740,N_320,N_237);
nand U741 (N_741,N_338,N_436);
nor U742 (N_742,N_317,N_332);
xnor U743 (N_743,N_107,N_459);
or U744 (N_744,N_486,N_396);
nand U745 (N_745,N_102,N_392);
xor U746 (N_746,N_437,N_77);
xnor U747 (N_747,N_97,N_293);
nand U748 (N_748,N_104,N_146);
xor U749 (N_749,N_276,N_53);
and U750 (N_750,N_329,N_209);
xor U751 (N_751,N_81,N_435);
nor U752 (N_752,N_253,N_295);
nor U753 (N_753,N_350,N_186);
xnor U754 (N_754,N_327,N_288);
or U755 (N_755,N_210,N_308);
or U756 (N_756,N_212,N_396);
nor U757 (N_757,N_274,N_297);
xnor U758 (N_758,N_391,N_17);
or U759 (N_759,N_388,N_97);
nand U760 (N_760,N_182,N_432);
nand U761 (N_761,N_100,N_79);
nand U762 (N_762,N_65,N_176);
and U763 (N_763,N_274,N_72);
xnor U764 (N_764,N_180,N_454);
and U765 (N_765,N_277,N_326);
or U766 (N_766,N_481,N_196);
nor U767 (N_767,N_7,N_434);
nand U768 (N_768,N_224,N_429);
or U769 (N_769,N_403,N_24);
and U770 (N_770,N_373,N_116);
xnor U771 (N_771,N_15,N_356);
xor U772 (N_772,N_487,N_73);
xor U773 (N_773,N_489,N_416);
nor U774 (N_774,N_110,N_144);
nand U775 (N_775,N_148,N_413);
or U776 (N_776,N_228,N_187);
or U777 (N_777,N_121,N_189);
or U778 (N_778,N_198,N_255);
nor U779 (N_779,N_447,N_76);
and U780 (N_780,N_221,N_187);
or U781 (N_781,N_46,N_199);
xnor U782 (N_782,N_304,N_171);
or U783 (N_783,N_167,N_82);
nand U784 (N_784,N_119,N_255);
and U785 (N_785,N_472,N_247);
nor U786 (N_786,N_304,N_431);
nand U787 (N_787,N_470,N_175);
nand U788 (N_788,N_328,N_227);
nor U789 (N_789,N_203,N_428);
nor U790 (N_790,N_306,N_429);
and U791 (N_791,N_463,N_151);
or U792 (N_792,N_471,N_122);
nand U793 (N_793,N_119,N_139);
nor U794 (N_794,N_307,N_88);
nand U795 (N_795,N_139,N_82);
and U796 (N_796,N_423,N_170);
and U797 (N_797,N_193,N_444);
nand U798 (N_798,N_117,N_160);
xor U799 (N_799,N_428,N_246);
nor U800 (N_800,N_453,N_205);
nand U801 (N_801,N_365,N_421);
xnor U802 (N_802,N_355,N_193);
or U803 (N_803,N_463,N_153);
nor U804 (N_804,N_402,N_336);
or U805 (N_805,N_44,N_287);
and U806 (N_806,N_23,N_442);
or U807 (N_807,N_334,N_209);
nand U808 (N_808,N_94,N_268);
nand U809 (N_809,N_226,N_319);
nor U810 (N_810,N_218,N_307);
nand U811 (N_811,N_280,N_199);
and U812 (N_812,N_49,N_431);
or U813 (N_813,N_260,N_105);
or U814 (N_814,N_206,N_184);
and U815 (N_815,N_272,N_480);
nand U816 (N_816,N_113,N_125);
nand U817 (N_817,N_293,N_435);
xnor U818 (N_818,N_400,N_227);
nand U819 (N_819,N_118,N_176);
and U820 (N_820,N_220,N_146);
nand U821 (N_821,N_92,N_193);
xnor U822 (N_822,N_132,N_405);
or U823 (N_823,N_198,N_150);
or U824 (N_824,N_92,N_84);
or U825 (N_825,N_294,N_316);
nand U826 (N_826,N_342,N_424);
xnor U827 (N_827,N_173,N_287);
nand U828 (N_828,N_286,N_297);
and U829 (N_829,N_382,N_316);
or U830 (N_830,N_364,N_227);
xnor U831 (N_831,N_54,N_95);
or U832 (N_832,N_39,N_421);
or U833 (N_833,N_186,N_225);
and U834 (N_834,N_262,N_172);
and U835 (N_835,N_37,N_420);
and U836 (N_836,N_250,N_151);
nor U837 (N_837,N_149,N_183);
nand U838 (N_838,N_205,N_222);
or U839 (N_839,N_235,N_296);
nand U840 (N_840,N_401,N_10);
xnor U841 (N_841,N_9,N_307);
or U842 (N_842,N_370,N_209);
nor U843 (N_843,N_223,N_493);
nand U844 (N_844,N_499,N_96);
nand U845 (N_845,N_203,N_290);
and U846 (N_846,N_364,N_365);
nand U847 (N_847,N_151,N_306);
or U848 (N_848,N_355,N_196);
nand U849 (N_849,N_101,N_179);
xor U850 (N_850,N_326,N_381);
nand U851 (N_851,N_445,N_333);
xnor U852 (N_852,N_19,N_388);
or U853 (N_853,N_387,N_444);
nand U854 (N_854,N_219,N_89);
xnor U855 (N_855,N_151,N_251);
nand U856 (N_856,N_359,N_467);
nor U857 (N_857,N_64,N_434);
xor U858 (N_858,N_427,N_428);
nor U859 (N_859,N_218,N_466);
nor U860 (N_860,N_433,N_300);
nor U861 (N_861,N_454,N_93);
nand U862 (N_862,N_390,N_187);
nand U863 (N_863,N_338,N_114);
nand U864 (N_864,N_47,N_13);
nor U865 (N_865,N_370,N_406);
nor U866 (N_866,N_104,N_487);
or U867 (N_867,N_361,N_28);
nand U868 (N_868,N_125,N_249);
or U869 (N_869,N_84,N_33);
xor U870 (N_870,N_45,N_440);
xnor U871 (N_871,N_28,N_328);
and U872 (N_872,N_490,N_244);
xor U873 (N_873,N_102,N_242);
nor U874 (N_874,N_203,N_382);
nand U875 (N_875,N_262,N_152);
nand U876 (N_876,N_484,N_174);
nand U877 (N_877,N_296,N_427);
and U878 (N_878,N_388,N_419);
nand U879 (N_879,N_427,N_167);
xnor U880 (N_880,N_409,N_319);
nor U881 (N_881,N_52,N_225);
nor U882 (N_882,N_369,N_229);
or U883 (N_883,N_324,N_99);
xnor U884 (N_884,N_346,N_474);
nor U885 (N_885,N_49,N_109);
xor U886 (N_886,N_482,N_339);
and U887 (N_887,N_100,N_379);
nand U888 (N_888,N_171,N_476);
nor U889 (N_889,N_401,N_279);
and U890 (N_890,N_274,N_480);
and U891 (N_891,N_182,N_314);
nor U892 (N_892,N_100,N_64);
and U893 (N_893,N_195,N_255);
xor U894 (N_894,N_307,N_80);
xor U895 (N_895,N_141,N_296);
or U896 (N_896,N_305,N_241);
and U897 (N_897,N_417,N_47);
and U898 (N_898,N_86,N_109);
nor U899 (N_899,N_312,N_91);
nor U900 (N_900,N_327,N_343);
and U901 (N_901,N_166,N_184);
nand U902 (N_902,N_378,N_113);
nor U903 (N_903,N_97,N_360);
or U904 (N_904,N_126,N_438);
or U905 (N_905,N_420,N_447);
and U906 (N_906,N_495,N_467);
xnor U907 (N_907,N_296,N_437);
nor U908 (N_908,N_165,N_54);
nand U909 (N_909,N_336,N_212);
nor U910 (N_910,N_443,N_301);
xnor U911 (N_911,N_312,N_311);
xnor U912 (N_912,N_473,N_172);
or U913 (N_913,N_344,N_40);
or U914 (N_914,N_102,N_324);
or U915 (N_915,N_351,N_249);
or U916 (N_916,N_368,N_138);
or U917 (N_917,N_414,N_71);
or U918 (N_918,N_227,N_414);
xnor U919 (N_919,N_171,N_471);
nor U920 (N_920,N_499,N_323);
and U921 (N_921,N_379,N_168);
nand U922 (N_922,N_171,N_59);
xor U923 (N_923,N_439,N_128);
xor U924 (N_924,N_474,N_209);
or U925 (N_925,N_101,N_152);
nand U926 (N_926,N_299,N_268);
or U927 (N_927,N_131,N_213);
xor U928 (N_928,N_451,N_57);
and U929 (N_929,N_265,N_277);
nor U930 (N_930,N_206,N_54);
nor U931 (N_931,N_284,N_137);
xor U932 (N_932,N_475,N_156);
or U933 (N_933,N_24,N_366);
nor U934 (N_934,N_390,N_202);
xor U935 (N_935,N_7,N_241);
and U936 (N_936,N_465,N_371);
nor U937 (N_937,N_357,N_226);
nand U938 (N_938,N_71,N_444);
or U939 (N_939,N_489,N_384);
xnor U940 (N_940,N_95,N_324);
and U941 (N_941,N_37,N_163);
xnor U942 (N_942,N_411,N_22);
or U943 (N_943,N_456,N_78);
or U944 (N_944,N_189,N_64);
xnor U945 (N_945,N_231,N_404);
or U946 (N_946,N_245,N_139);
nand U947 (N_947,N_147,N_390);
xnor U948 (N_948,N_255,N_425);
and U949 (N_949,N_279,N_254);
nor U950 (N_950,N_317,N_71);
nand U951 (N_951,N_369,N_443);
xnor U952 (N_952,N_311,N_62);
nand U953 (N_953,N_74,N_192);
nand U954 (N_954,N_46,N_247);
and U955 (N_955,N_267,N_83);
nand U956 (N_956,N_284,N_437);
or U957 (N_957,N_441,N_429);
and U958 (N_958,N_272,N_12);
xnor U959 (N_959,N_421,N_306);
or U960 (N_960,N_482,N_462);
or U961 (N_961,N_228,N_457);
nand U962 (N_962,N_270,N_484);
nand U963 (N_963,N_233,N_361);
xor U964 (N_964,N_203,N_88);
and U965 (N_965,N_243,N_112);
and U966 (N_966,N_347,N_279);
and U967 (N_967,N_280,N_437);
nor U968 (N_968,N_459,N_236);
nand U969 (N_969,N_439,N_135);
xnor U970 (N_970,N_72,N_283);
or U971 (N_971,N_443,N_13);
nand U972 (N_972,N_479,N_51);
nand U973 (N_973,N_178,N_229);
xor U974 (N_974,N_112,N_238);
nand U975 (N_975,N_215,N_358);
nor U976 (N_976,N_415,N_472);
and U977 (N_977,N_389,N_53);
nor U978 (N_978,N_412,N_261);
nor U979 (N_979,N_168,N_366);
and U980 (N_980,N_292,N_175);
nor U981 (N_981,N_39,N_121);
nand U982 (N_982,N_466,N_189);
nand U983 (N_983,N_108,N_490);
xor U984 (N_984,N_461,N_173);
xnor U985 (N_985,N_298,N_492);
nor U986 (N_986,N_28,N_404);
and U987 (N_987,N_146,N_412);
nand U988 (N_988,N_44,N_103);
xnor U989 (N_989,N_161,N_139);
nor U990 (N_990,N_191,N_396);
xnor U991 (N_991,N_326,N_247);
or U992 (N_992,N_497,N_43);
nor U993 (N_993,N_10,N_268);
xor U994 (N_994,N_190,N_354);
nand U995 (N_995,N_249,N_288);
and U996 (N_996,N_29,N_297);
nand U997 (N_997,N_31,N_295);
and U998 (N_998,N_287,N_31);
nand U999 (N_999,N_305,N_323);
and U1000 (N_1000,N_629,N_699);
xor U1001 (N_1001,N_615,N_714);
xor U1002 (N_1002,N_859,N_634);
nand U1003 (N_1003,N_655,N_858);
nand U1004 (N_1004,N_715,N_816);
or U1005 (N_1005,N_993,N_737);
and U1006 (N_1006,N_955,N_742);
nand U1007 (N_1007,N_566,N_956);
nor U1008 (N_1008,N_710,N_645);
xnor U1009 (N_1009,N_686,N_825);
nand U1010 (N_1010,N_977,N_729);
or U1011 (N_1011,N_631,N_899);
xnor U1012 (N_1012,N_787,N_864);
nand U1013 (N_1013,N_754,N_532);
xnor U1014 (N_1014,N_973,N_670);
and U1015 (N_1015,N_675,N_753);
and U1016 (N_1016,N_893,N_616);
xor U1017 (N_1017,N_649,N_549);
nand U1018 (N_1018,N_589,N_559);
xor U1019 (N_1019,N_954,N_668);
or U1020 (N_1020,N_691,N_917);
nor U1021 (N_1021,N_922,N_530);
or U1022 (N_1022,N_726,N_740);
xor U1023 (N_1023,N_966,N_785);
or U1024 (N_1024,N_995,N_693);
xor U1025 (N_1025,N_799,N_554);
or U1026 (N_1026,N_569,N_635);
nand U1027 (N_1027,N_750,N_997);
nor U1028 (N_1028,N_711,N_915);
or U1029 (N_1029,N_651,N_582);
nand U1030 (N_1030,N_961,N_936);
or U1031 (N_1031,N_602,N_947);
or U1032 (N_1032,N_579,N_950);
nand U1033 (N_1033,N_663,N_806);
nand U1034 (N_1034,N_680,N_801);
and U1035 (N_1035,N_830,N_679);
and U1036 (N_1036,N_617,N_879);
and U1037 (N_1037,N_847,N_882);
and U1038 (N_1038,N_507,N_720);
and U1039 (N_1039,N_842,N_919);
and U1040 (N_1040,N_832,N_914);
or U1041 (N_1041,N_578,N_853);
nand U1042 (N_1042,N_875,N_817);
nand U1043 (N_1043,N_876,N_521);
or U1044 (N_1044,N_805,N_683);
xor U1045 (N_1045,N_959,N_650);
xor U1046 (N_1046,N_611,N_940);
xor U1047 (N_1047,N_888,N_577);
or U1048 (N_1048,N_976,N_938);
nand U1049 (N_1049,N_708,N_503);
or U1050 (N_1050,N_734,N_793);
nor U1051 (N_1051,N_908,N_828);
and U1052 (N_1052,N_562,N_697);
or U1053 (N_1053,N_700,N_748);
nor U1054 (N_1054,N_547,N_502);
nand U1055 (N_1055,N_618,N_972);
or U1056 (N_1056,N_756,N_979);
and U1057 (N_1057,N_584,N_990);
nor U1058 (N_1058,N_820,N_774);
nor U1059 (N_1059,N_813,N_719);
or U1060 (N_1060,N_648,N_925);
and U1061 (N_1061,N_945,N_969);
xor U1062 (N_1062,N_594,N_544);
or U1063 (N_1063,N_778,N_926);
nor U1064 (N_1064,N_810,N_883);
or U1065 (N_1065,N_836,N_627);
nor U1066 (N_1066,N_674,N_656);
nor U1067 (N_1067,N_600,N_570);
nor U1068 (N_1068,N_766,N_855);
and U1069 (N_1069,N_890,N_684);
nand U1070 (N_1070,N_643,N_667);
xor U1071 (N_1071,N_534,N_736);
and U1072 (N_1072,N_593,N_531);
and U1073 (N_1073,N_989,N_580);
and U1074 (N_1074,N_827,N_835);
and U1075 (N_1075,N_854,N_550);
and U1076 (N_1076,N_543,N_669);
nand U1077 (N_1077,N_826,N_741);
and U1078 (N_1078,N_731,N_641);
or U1079 (N_1079,N_844,N_840);
xnor U1080 (N_1080,N_970,N_598);
and U1081 (N_1081,N_818,N_768);
and U1082 (N_1082,N_906,N_506);
and U1083 (N_1083,N_717,N_704);
xnor U1084 (N_1084,N_537,N_839);
nor U1085 (N_1085,N_895,N_770);
xnor U1086 (N_1086,N_533,N_843);
xor U1087 (N_1087,N_613,N_500);
nor U1088 (N_1088,N_776,N_520);
nand U1089 (N_1089,N_894,N_980);
nand U1090 (N_1090,N_581,N_536);
or U1091 (N_1091,N_953,N_690);
or U1092 (N_1092,N_743,N_718);
or U1093 (N_1093,N_501,N_789);
nor U1094 (N_1094,N_671,N_733);
nor U1095 (N_1095,N_659,N_913);
and U1096 (N_1096,N_658,N_783);
nand U1097 (N_1097,N_522,N_588);
xnor U1098 (N_1098,N_934,N_732);
and U1099 (N_1099,N_975,N_705);
xnor U1100 (N_1100,N_621,N_504);
nor U1101 (N_1101,N_749,N_886);
nor U1102 (N_1102,N_924,N_777);
nor U1103 (N_1103,N_996,N_623);
nand U1104 (N_1104,N_505,N_986);
or U1105 (N_1105,N_573,N_660);
xor U1106 (N_1106,N_511,N_921);
and U1107 (N_1107,N_971,N_646);
or U1108 (N_1108,N_512,N_516);
nor U1109 (N_1109,N_861,N_608);
nand U1110 (N_1110,N_790,N_760);
xnor U1111 (N_1111,N_586,N_775);
xnor U1112 (N_1112,N_653,N_898);
or U1113 (N_1113,N_892,N_599);
or U1114 (N_1114,N_662,N_991);
xnor U1115 (N_1115,N_786,N_513);
nor U1116 (N_1116,N_571,N_869);
xor U1117 (N_1117,N_982,N_865);
and U1118 (N_1118,N_916,N_657);
and U1119 (N_1119,N_757,N_601);
and U1120 (N_1120,N_791,N_891);
and U1121 (N_1121,N_951,N_746);
or U1122 (N_1122,N_567,N_707);
nor U1123 (N_1123,N_804,N_630);
xnor U1124 (N_1124,N_610,N_872);
or U1125 (N_1125,N_761,N_735);
nor U1126 (N_1126,N_609,N_837);
and U1127 (N_1127,N_900,N_800);
nor U1128 (N_1128,N_905,N_730);
and U1129 (N_1129,N_860,N_745);
nand U1130 (N_1130,N_713,N_937);
nand U1131 (N_1131,N_862,N_654);
nand U1132 (N_1132,N_563,N_878);
nand U1133 (N_1133,N_565,N_738);
nor U1134 (N_1134,N_931,N_845);
and U1135 (N_1135,N_802,N_901);
or U1136 (N_1136,N_968,N_620);
nand U1137 (N_1137,N_985,N_809);
nor U1138 (N_1138,N_685,N_762);
or U1139 (N_1139,N_927,N_984);
or U1140 (N_1140,N_633,N_612);
nor U1141 (N_1141,N_944,N_772);
or U1142 (N_1142,N_568,N_528);
or U1143 (N_1143,N_846,N_765);
nor U1144 (N_1144,N_822,N_930);
nand U1145 (N_1145,N_923,N_935);
nor U1146 (N_1146,N_639,N_592);
nand U1147 (N_1147,N_603,N_518);
and U1148 (N_1148,N_885,N_852);
nor U1149 (N_1149,N_728,N_628);
and U1150 (N_1150,N_918,N_771);
nor U1151 (N_1151,N_622,N_698);
or U1152 (N_1152,N_625,N_517);
nor U1153 (N_1153,N_721,N_811);
xnor U1154 (N_1154,N_725,N_824);
nand U1155 (N_1155,N_831,N_548);
and U1156 (N_1156,N_540,N_644);
nand U1157 (N_1157,N_958,N_652);
or U1158 (N_1158,N_907,N_838);
nand U1159 (N_1159,N_856,N_692);
or U1160 (N_1160,N_677,N_576);
xnor U1161 (N_1161,N_624,N_561);
xor U1162 (N_1162,N_590,N_988);
or U1163 (N_1163,N_724,N_666);
xor U1164 (N_1164,N_779,N_539);
nand U1165 (N_1165,N_767,N_794);
nand U1166 (N_1166,N_850,N_797);
or U1167 (N_1167,N_759,N_965);
nand U1168 (N_1168,N_902,N_515);
or U1169 (N_1169,N_636,N_535);
or U1170 (N_1170,N_527,N_552);
nor U1171 (N_1171,N_673,N_596);
or U1172 (N_1172,N_591,N_744);
xor U1173 (N_1173,N_987,N_819);
xor U1174 (N_1174,N_933,N_874);
nor U1175 (N_1175,N_782,N_851);
nand U1176 (N_1176,N_815,N_682);
xnor U1177 (N_1177,N_703,N_614);
xor U1178 (N_1178,N_637,N_541);
and U1179 (N_1179,N_877,N_595);
nor U1180 (N_1180,N_585,N_546);
nand U1181 (N_1181,N_739,N_676);
nor U1182 (N_1182,N_689,N_928);
xnor U1183 (N_1183,N_727,N_903);
and U1184 (N_1184,N_857,N_723);
xnor U1185 (N_1185,N_747,N_664);
or U1186 (N_1186,N_694,N_868);
nand U1187 (N_1187,N_803,N_716);
or U1188 (N_1188,N_998,N_632);
or U1189 (N_1189,N_911,N_763);
or U1190 (N_1190,N_796,N_795);
nor U1191 (N_1191,N_808,N_572);
and U1192 (N_1192,N_647,N_963);
xnor U1193 (N_1193,N_722,N_642);
and U1194 (N_1194,N_834,N_701);
nand U1195 (N_1195,N_688,N_798);
nor U1196 (N_1196,N_702,N_665);
nand U1197 (N_1197,N_587,N_709);
nor U1198 (N_1198,N_823,N_897);
or U1199 (N_1199,N_773,N_866);
nand U1200 (N_1200,N_781,N_526);
nor U1201 (N_1201,N_681,N_880);
nor U1202 (N_1202,N_994,N_583);
and U1203 (N_1203,N_514,N_524);
and U1204 (N_1204,N_626,N_560);
nand U1205 (N_1205,N_943,N_525);
or U1206 (N_1206,N_941,N_758);
nand U1207 (N_1207,N_867,N_889);
nor U1208 (N_1208,N_607,N_896);
nor U1209 (N_1209,N_841,N_814);
and U1210 (N_1210,N_821,N_553);
and U1211 (N_1211,N_942,N_992);
or U1212 (N_1212,N_881,N_696);
xor U1213 (N_1213,N_529,N_606);
and U1214 (N_1214,N_640,N_870);
or U1215 (N_1215,N_920,N_769);
nand U1216 (N_1216,N_755,N_849);
xnor U1217 (N_1217,N_983,N_661);
nand U1218 (N_1218,N_912,N_557);
nor U1219 (N_1219,N_946,N_904);
and U1220 (N_1220,N_764,N_929);
or U1221 (N_1221,N_687,N_974);
and U1222 (N_1222,N_932,N_962);
nand U1223 (N_1223,N_555,N_751);
xnor U1224 (N_1224,N_510,N_752);
or U1225 (N_1225,N_784,N_981);
nand U1226 (N_1226,N_957,N_678);
xor U1227 (N_1227,N_910,N_884);
and U1228 (N_1228,N_952,N_863);
nor U1229 (N_1229,N_556,N_523);
and U1230 (N_1230,N_604,N_788);
and U1231 (N_1231,N_960,N_564);
nor U1232 (N_1232,N_967,N_964);
and U1233 (N_1233,N_605,N_873);
and U1234 (N_1234,N_558,N_638);
nor U1235 (N_1235,N_871,N_695);
nand U1236 (N_1236,N_780,N_978);
and U1237 (N_1237,N_949,N_939);
xor U1238 (N_1238,N_887,N_619);
nand U1239 (N_1239,N_948,N_575);
nand U1240 (N_1240,N_833,N_792);
and U1241 (N_1241,N_508,N_509);
nand U1242 (N_1242,N_551,N_574);
xor U1243 (N_1243,N_999,N_712);
nor U1244 (N_1244,N_545,N_829);
nor U1245 (N_1245,N_597,N_538);
nand U1246 (N_1246,N_706,N_542);
xnor U1247 (N_1247,N_807,N_672);
nand U1248 (N_1248,N_519,N_848);
xor U1249 (N_1249,N_909,N_812);
nor U1250 (N_1250,N_657,N_509);
and U1251 (N_1251,N_632,N_728);
xor U1252 (N_1252,N_767,N_811);
nor U1253 (N_1253,N_938,N_795);
nor U1254 (N_1254,N_977,N_786);
nor U1255 (N_1255,N_908,N_793);
and U1256 (N_1256,N_746,N_656);
or U1257 (N_1257,N_622,N_524);
nand U1258 (N_1258,N_955,N_660);
and U1259 (N_1259,N_777,N_782);
xnor U1260 (N_1260,N_756,N_763);
and U1261 (N_1261,N_602,N_974);
or U1262 (N_1262,N_631,N_664);
xor U1263 (N_1263,N_766,N_595);
xor U1264 (N_1264,N_860,N_564);
or U1265 (N_1265,N_606,N_749);
xor U1266 (N_1266,N_927,N_598);
and U1267 (N_1267,N_744,N_502);
nor U1268 (N_1268,N_597,N_887);
nor U1269 (N_1269,N_704,N_630);
and U1270 (N_1270,N_764,N_686);
nor U1271 (N_1271,N_697,N_654);
and U1272 (N_1272,N_996,N_585);
nor U1273 (N_1273,N_875,N_667);
or U1274 (N_1274,N_675,N_622);
xnor U1275 (N_1275,N_531,N_574);
xor U1276 (N_1276,N_764,N_870);
nor U1277 (N_1277,N_998,N_637);
and U1278 (N_1278,N_930,N_922);
xor U1279 (N_1279,N_886,N_756);
nand U1280 (N_1280,N_828,N_801);
or U1281 (N_1281,N_838,N_906);
or U1282 (N_1282,N_778,N_949);
xor U1283 (N_1283,N_772,N_947);
and U1284 (N_1284,N_871,N_722);
xor U1285 (N_1285,N_696,N_951);
nand U1286 (N_1286,N_557,N_781);
or U1287 (N_1287,N_952,N_832);
nand U1288 (N_1288,N_932,N_590);
nand U1289 (N_1289,N_823,N_816);
nor U1290 (N_1290,N_757,N_834);
and U1291 (N_1291,N_760,N_742);
nand U1292 (N_1292,N_763,N_508);
xor U1293 (N_1293,N_830,N_681);
and U1294 (N_1294,N_898,N_528);
xnor U1295 (N_1295,N_706,N_710);
nand U1296 (N_1296,N_739,N_642);
or U1297 (N_1297,N_586,N_745);
nand U1298 (N_1298,N_975,N_551);
or U1299 (N_1299,N_549,N_653);
or U1300 (N_1300,N_606,N_878);
or U1301 (N_1301,N_989,N_709);
nand U1302 (N_1302,N_906,N_515);
xor U1303 (N_1303,N_635,N_786);
nand U1304 (N_1304,N_570,N_551);
nand U1305 (N_1305,N_914,N_607);
xnor U1306 (N_1306,N_888,N_894);
nor U1307 (N_1307,N_996,N_992);
and U1308 (N_1308,N_569,N_940);
xnor U1309 (N_1309,N_549,N_764);
and U1310 (N_1310,N_514,N_829);
xnor U1311 (N_1311,N_539,N_864);
nor U1312 (N_1312,N_897,N_951);
xor U1313 (N_1313,N_675,N_736);
nand U1314 (N_1314,N_670,N_558);
xnor U1315 (N_1315,N_861,N_737);
nor U1316 (N_1316,N_581,N_645);
xnor U1317 (N_1317,N_968,N_881);
and U1318 (N_1318,N_852,N_793);
or U1319 (N_1319,N_829,N_694);
or U1320 (N_1320,N_812,N_510);
and U1321 (N_1321,N_782,N_857);
nand U1322 (N_1322,N_942,N_983);
or U1323 (N_1323,N_795,N_564);
nor U1324 (N_1324,N_913,N_708);
nor U1325 (N_1325,N_856,N_701);
or U1326 (N_1326,N_728,N_561);
nor U1327 (N_1327,N_618,N_571);
and U1328 (N_1328,N_690,N_821);
xnor U1329 (N_1329,N_516,N_633);
nor U1330 (N_1330,N_514,N_613);
nor U1331 (N_1331,N_863,N_502);
and U1332 (N_1332,N_992,N_636);
and U1333 (N_1333,N_788,N_644);
xor U1334 (N_1334,N_987,N_993);
nor U1335 (N_1335,N_506,N_872);
nor U1336 (N_1336,N_900,N_929);
and U1337 (N_1337,N_930,N_830);
nand U1338 (N_1338,N_502,N_818);
xnor U1339 (N_1339,N_996,N_911);
xnor U1340 (N_1340,N_736,N_899);
or U1341 (N_1341,N_598,N_830);
nand U1342 (N_1342,N_784,N_739);
nor U1343 (N_1343,N_734,N_967);
or U1344 (N_1344,N_903,N_603);
and U1345 (N_1345,N_917,N_671);
nand U1346 (N_1346,N_928,N_926);
or U1347 (N_1347,N_581,N_705);
xnor U1348 (N_1348,N_590,N_941);
xor U1349 (N_1349,N_507,N_739);
xnor U1350 (N_1350,N_857,N_660);
and U1351 (N_1351,N_768,N_540);
nor U1352 (N_1352,N_667,N_984);
xor U1353 (N_1353,N_849,N_677);
nor U1354 (N_1354,N_828,N_787);
nand U1355 (N_1355,N_974,N_506);
nand U1356 (N_1356,N_755,N_756);
and U1357 (N_1357,N_754,N_566);
or U1358 (N_1358,N_566,N_896);
xnor U1359 (N_1359,N_525,N_792);
nand U1360 (N_1360,N_926,N_919);
xor U1361 (N_1361,N_515,N_659);
xnor U1362 (N_1362,N_947,N_552);
nor U1363 (N_1363,N_868,N_530);
xor U1364 (N_1364,N_728,N_848);
nand U1365 (N_1365,N_865,N_679);
nand U1366 (N_1366,N_647,N_760);
or U1367 (N_1367,N_922,N_959);
xor U1368 (N_1368,N_796,N_552);
or U1369 (N_1369,N_705,N_879);
and U1370 (N_1370,N_789,N_631);
or U1371 (N_1371,N_715,N_709);
or U1372 (N_1372,N_812,N_648);
nor U1373 (N_1373,N_950,N_679);
and U1374 (N_1374,N_731,N_594);
or U1375 (N_1375,N_514,N_794);
or U1376 (N_1376,N_819,N_749);
or U1377 (N_1377,N_581,N_702);
nor U1378 (N_1378,N_502,N_930);
and U1379 (N_1379,N_739,N_523);
nand U1380 (N_1380,N_515,N_604);
and U1381 (N_1381,N_978,N_683);
nand U1382 (N_1382,N_985,N_553);
nand U1383 (N_1383,N_783,N_714);
xor U1384 (N_1384,N_776,N_924);
or U1385 (N_1385,N_895,N_815);
or U1386 (N_1386,N_652,N_693);
nand U1387 (N_1387,N_660,N_809);
nor U1388 (N_1388,N_583,N_877);
nor U1389 (N_1389,N_972,N_892);
nor U1390 (N_1390,N_995,N_752);
xnor U1391 (N_1391,N_512,N_532);
and U1392 (N_1392,N_533,N_648);
xnor U1393 (N_1393,N_542,N_812);
or U1394 (N_1394,N_572,N_716);
nor U1395 (N_1395,N_703,N_852);
and U1396 (N_1396,N_771,N_886);
nand U1397 (N_1397,N_768,N_726);
and U1398 (N_1398,N_612,N_874);
and U1399 (N_1399,N_690,N_783);
nor U1400 (N_1400,N_688,N_513);
nor U1401 (N_1401,N_715,N_834);
or U1402 (N_1402,N_942,N_756);
nand U1403 (N_1403,N_611,N_520);
and U1404 (N_1404,N_723,N_982);
nand U1405 (N_1405,N_537,N_592);
nand U1406 (N_1406,N_805,N_873);
xor U1407 (N_1407,N_894,N_874);
and U1408 (N_1408,N_971,N_602);
nor U1409 (N_1409,N_533,N_558);
nor U1410 (N_1410,N_748,N_857);
nor U1411 (N_1411,N_989,N_678);
nand U1412 (N_1412,N_957,N_883);
and U1413 (N_1413,N_697,N_680);
xor U1414 (N_1414,N_644,N_725);
and U1415 (N_1415,N_954,N_538);
or U1416 (N_1416,N_691,N_509);
or U1417 (N_1417,N_809,N_698);
and U1418 (N_1418,N_615,N_524);
nor U1419 (N_1419,N_878,N_608);
nor U1420 (N_1420,N_850,N_565);
nand U1421 (N_1421,N_852,N_946);
xor U1422 (N_1422,N_676,N_744);
and U1423 (N_1423,N_731,N_985);
and U1424 (N_1424,N_587,N_688);
and U1425 (N_1425,N_756,N_731);
nand U1426 (N_1426,N_887,N_788);
and U1427 (N_1427,N_830,N_867);
nor U1428 (N_1428,N_682,N_806);
or U1429 (N_1429,N_739,N_572);
nor U1430 (N_1430,N_540,N_555);
xor U1431 (N_1431,N_552,N_561);
nor U1432 (N_1432,N_611,N_610);
and U1433 (N_1433,N_964,N_526);
nor U1434 (N_1434,N_740,N_533);
and U1435 (N_1435,N_705,N_834);
xnor U1436 (N_1436,N_648,N_797);
and U1437 (N_1437,N_631,N_938);
xnor U1438 (N_1438,N_754,N_988);
nand U1439 (N_1439,N_592,N_796);
nor U1440 (N_1440,N_739,N_926);
nor U1441 (N_1441,N_688,N_600);
xnor U1442 (N_1442,N_677,N_564);
or U1443 (N_1443,N_572,N_972);
or U1444 (N_1444,N_810,N_889);
or U1445 (N_1445,N_535,N_966);
nand U1446 (N_1446,N_911,N_779);
and U1447 (N_1447,N_514,N_539);
nor U1448 (N_1448,N_799,N_842);
and U1449 (N_1449,N_879,N_531);
nor U1450 (N_1450,N_701,N_823);
nor U1451 (N_1451,N_633,N_673);
or U1452 (N_1452,N_655,N_724);
nor U1453 (N_1453,N_715,N_794);
xor U1454 (N_1454,N_972,N_935);
and U1455 (N_1455,N_573,N_580);
xor U1456 (N_1456,N_807,N_628);
and U1457 (N_1457,N_768,N_899);
or U1458 (N_1458,N_706,N_997);
nor U1459 (N_1459,N_643,N_820);
nand U1460 (N_1460,N_618,N_788);
xnor U1461 (N_1461,N_973,N_862);
or U1462 (N_1462,N_660,N_939);
xnor U1463 (N_1463,N_728,N_921);
xnor U1464 (N_1464,N_647,N_887);
nand U1465 (N_1465,N_541,N_895);
nand U1466 (N_1466,N_948,N_695);
nand U1467 (N_1467,N_720,N_928);
or U1468 (N_1468,N_739,N_629);
and U1469 (N_1469,N_619,N_909);
xor U1470 (N_1470,N_913,N_651);
xor U1471 (N_1471,N_884,N_943);
xnor U1472 (N_1472,N_679,N_862);
nand U1473 (N_1473,N_861,N_984);
xnor U1474 (N_1474,N_856,N_923);
nand U1475 (N_1475,N_637,N_927);
nor U1476 (N_1476,N_973,N_794);
xor U1477 (N_1477,N_798,N_772);
nand U1478 (N_1478,N_936,N_697);
and U1479 (N_1479,N_913,N_867);
nand U1480 (N_1480,N_632,N_615);
nand U1481 (N_1481,N_945,N_981);
and U1482 (N_1482,N_958,N_604);
and U1483 (N_1483,N_613,N_936);
nand U1484 (N_1484,N_806,N_679);
nand U1485 (N_1485,N_752,N_975);
xor U1486 (N_1486,N_802,N_543);
nand U1487 (N_1487,N_792,N_737);
xnor U1488 (N_1488,N_679,N_878);
or U1489 (N_1489,N_787,N_723);
and U1490 (N_1490,N_942,N_883);
nor U1491 (N_1491,N_646,N_725);
nor U1492 (N_1492,N_675,N_989);
or U1493 (N_1493,N_536,N_959);
or U1494 (N_1494,N_552,N_887);
or U1495 (N_1495,N_806,N_535);
nand U1496 (N_1496,N_881,N_938);
nand U1497 (N_1497,N_767,N_879);
and U1498 (N_1498,N_777,N_614);
nand U1499 (N_1499,N_906,N_691);
nor U1500 (N_1500,N_1000,N_1421);
nor U1501 (N_1501,N_1115,N_1209);
xor U1502 (N_1502,N_1225,N_1346);
nor U1503 (N_1503,N_1074,N_1119);
or U1504 (N_1504,N_1282,N_1254);
nand U1505 (N_1505,N_1499,N_1237);
nand U1506 (N_1506,N_1102,N_1287);
and U1507 (N_1507,N_1351,N_1126);
or U1508 (N_1508,N_1096,N_1312);
xor U1509 (N_1509,N_1370,N_1044);
or U1510 (N_1510,N_1054,N_1272);
and U1511 (N_1511,N_1260,N_1223);
nor U1512 (N_1512,N_1374,N_1334);
or U1513 (N_1513,N_1252,N_1311);
nand U1514 (N_1514,N_1232,N_1073);
nor U1515 (N_1515,N_1195,N_1284);
nand U1516 (N_1516,N_1382,N_1434);
or U1517 (N_1517,N_1161,N_1157);
nor U1518 (N_1518,N_1384,N_1429);
and U1519 (N_1519,N_1385,N_1299);
nand U1520 (N_1520,N_1133,N_1456);
nor U1521 (N_1521,N_1337,N_1250);
xor U1522 (N_1522,N_1248,N_1476);
xor U1523 (N_1523,N_1490,N_1240);
or U1524 (N_1524,N_1274,N_1401);
or U1525 (N_1525,N_1449,N_1051);
xor U1526 (N_1526,N_1121,N_1317);
and U1527 (N_1527,N_1338,N_1256);
and U1528 (N_1528,N_1494,N_1495);
nand U1529 (N_1529,N_1049,N_1194);
and U1530 (N_1530,N_1373,N_1182);
or U1531 (N_1531,N_1345,N_1415);
or U1532 (N_1532,N_1143,N_1417);
nand U1533 (N_1533,N_1149,N_1170);
and U1534 (N_1534,N_1220,N_1164);
or U1535 (N_1535,N_1258,N_1275);
nor U1536 (N_1536,N_1086,N_1367);
xnor U1537 (N_1537,N_1413,N_1156);
or U1538 (N_1538,N_1463,N_1215);
or U1539 (N_1539,N_1171,N_1344);
and U1540 (N_1540,N_1448,N_1280);
xnor U1541 (N_1541,N_1372,N_1309);
and U1542 (N_1542,N_1444,N_1199);
and U1543 (N_1543,N_1188,N_1261);
and U1544 (N_1544,N_1124,N_1276);
nor U1545 (N_1545,N_1196,N_1058);
xor U1546 (N_1546,N_1430,N_1094);
xor U1547 (N_1547,N_1079,N_1389);
xor U1548 (N_1548,N_1439,N_1023);
nor U1549 (N_1549,N_1354,N_1033);
and U1550 (N_1550,N_1349,N_1297);
nor U1551 (N_1551,N_1056,N_1239);
nor U1552 (N_1552,N_1486,N_1048);
or U1553 (N_1553,N_1104,N_1355);
nand U1554 (N_1554,N_1208,N_1021);
xor U1555 (N_1555,N_1197,N_1212);
xnor U1556 (N_1556,N_1247,N_1014);
and U1557 (N_1557,N_1175,N_1036);
nor U1558 (N_1558,N_1085,N_1039);
xor U1559 (N_1559,N_1292,N_1469);
and U1560 (N_1560,N_1362,N_1467);
xnor U1561 (N_1561,N_1342,N_1356);
nand U1562 (N_1562,N_1004,N_1482);
and U1563 (N_1563,N_1146,N_1333);
xnor U1564 (N_1564,N_1003,N_1388);
or U1565 (N_1565,N_1410,N_1375);
nor U1566 (N_1566,N_1271,N_1226);
nand U1567 (N_1567,N_1172,N_1443);
and U1568 (N_1568,N_1452,N_1283);
and U1569 (N_1569,N_1174,N_1211);
nand U1570 (N_1570,N_1315,N_1458);
and U1571 (N_1571,N_1107,N_1268);
xor U1572 (N_1572,N_1160,N_1442);
xor U1573 (N_1573,N_1162,N_1350);
and U1574 (N_1574,N_1399,N_1214);
xor U1575 (N_1575,N_1493,N_1433);
xnor U1576 (N_1576,N_1072,N_1217);
xor U1577 (N_1577,N_1406,N_1113);
and U1578 (N_1578,N_1235,N_1114);
and U1579 (N_1579,N_1066,N_1454);
xor U1580 (N_1580,N_1169,N_1403);
and U1581 (N_1581,N_1358,N_1221);
or U1582 (N_1582,N_1123,N_1435);
or U1583 (N_1583,N_1386,N_1380);
xor U1584 (N_1584,N_1087,N_1378);
nand U1585 (N_1585,N_1077,N_1006);
or U1586 (N_1586,N_1238,N_1179);
and U1587 (N_1587,N_1065,N_1125);
nand U1588 (N_1588,N_1191,N_1219);
nand U1589 (N_1589,N_1100,N_1245);
or U1590 (N_1590,N_1042,N_1498);
nor U1591 (N_1591,N_1277,N_1041);
or U1592 (N_1592,N_1425,N_1178);
and U1593 (N_1593,N_1321,N_1427);
or U1594 (N_1594,N_1353,N_1291);
nor U1595 (N_1595,N_1198,N_1229);
nor U1596 (N_1596,N_1440,N_1141);
and U1597 (N_1597,N_1062,N_1393);
or U1598 (N_1598,N_1461,N_1270);
or U1599 (N_1599,N_1052,N_1336);
and U1600 (N_1600,N_1173,N_1364);
xnor U1601 (N_1601,N_1038,N_1492);
xnor U1602 (N_1602,N_1013,N_1070);
xnor U1603 (N_1603,N_1263,N_1426);
nand U1604 (N_1604,N_1383,N_1228);
nor U1605 (N_1605,N_1002,N_1045);
nor U1606 (N_1606,N_1347,N_1279);
xnor U1607 (N_1607,N_1447,N_1218);
nand U1608 (N_1608,N_1117,N_1488);
nand U1609 (N_1609,N_1255,N_1047);
or U1610 (N_1610,N_1416,N_1243);
nor U1611 (N_1611,N_1097,N_1207);
and U1612 (N_1612,N_1290,N_1071);
xor U1613 (N_1613,N_1091,N_1089);
or U1614 (N_1614,N_1025,N_1365);
nor U1615 (N_1615,N_1360,N_1431);
nor U1616 (N_1616,N_1253,N_1020);
and U1617 (N_1617,N_1293,N_1063);
and U1618 (N_1618,N_1496,N_1184);
xnor U1619 (N_1619,N_1151,N_1093);
xor U1620 (N_1620,N_1008,N_1497);
or U1621 (N_1621,N_1473,N_1110);
xor U1622 (N_1622,N_1475,N_1289);
or U1623 (N_1623,N_1186,N_1269);
and U1624 (N_1624,N_1264,N_1026);
and U1625 (N_1625,N_1230,N_1343);
xor U1626 (N_1626,N_1313,N_1316);
or U1627 (N_1627,N_1371,N_1394);
nor U1628 (N_1628,N_1140,N_1408);
or U1629 (N_1629,N_1428,N_1418);
nor U1630 (N_1630,N_1129,N_1200);
and U1631 (N_1631,N_1154,N_1075);
nor U1632 (N_1632,N_1022,N_1472);
or U1633 (N_1633,N_1001,N_1305);
nor U1634 (N_1634,N_1451,N_1481);
and U1635 (N_1635,N_1404,N_1294);
xor U1636 (N_1636,N_1028,N_1308);
and U1637 (N_1637,N_1328,N_1357);
xor U1638 (N_1638,N_1379,N_1165);
or U1639 (N_1639,N_1166,N_1242);
nor U1640 (N_1640,N_1301,N_1024);
xnor U1641 (N_1641,N_1368,N_1152);
or U1642 (N_1642,N_1470,N_1005);
or U1643 (N_1643,N_1095,N_1407);
or U1644 (N_1644,N_1348,N_1139);
and U1645 (N_1645,N_1148,N_1310);
or U1646 (N_1646,N_1314,N_1285);
xnor U1647 (N_1647,N_1320,N_1331);
or U1648 (N_1648,N_1450,N_1483);
or U1649 (N_1649,N_1017,N_1187);
xnor U1650 (N_1650,N_1414,N_1411);
nand U1651 (N_1651,N_1405,N_1167);
nand U1652 (N_1652,N_1259,N_1067);
and U1653 (N_1653,N_1183,N_1273);
nand U1654 (N_1654,N_1142,N_1474);
and U1655 (N_1655,N_1231,N_1122);
xor U1656 (N_1656,N_1236,N_1037);
nor U1657 (N_1657,N_1319,N_1090);
or U1658 (N_1658,N_1491,N_1078);
or U1659 (N_1659,N_1487,N_1249);
or U1660 (N_1660,N_1144,N_1340);
nand U1661 (N_1661,N_1213,N_1180);
xnor U1662 (N_1662,N_1335,N_1032);
and U1663 (N_1663,N_1359,N_1222);
nand U1664 (N_1664,N_1484,N_1084);
nand U1665 (N_1665,N_1307,N_1466);
nand U1666 (N_1666,N_1112,N_1082);
or U1667 (N_1667,N_1251,N_1131);
xor U1668 (N_1668,N_1332,N_1363);
xor U1669 (N_1669,N_1412,N_1296);
and U1670 (N_1670,N_1323,N_1118);
nor U1671 (N_1671,N_1281,N_1076);
or U1672 (N_1672,N_1424,N_1185);
xor U1673 (N_1673,N_1402,N_1009);
and U1674 (N_1674,N_1081,N_1327);
and U1675 (N_1675,N_1181,N_1192);
nor U1676 (N_1676,N_1019,N_1105);
or U1677 (N_1677,N_1163,N_1387);
nor U1678 (N_1678,N_1391,N_1061);
or U1679 (N_1679,N_1210,N_1304);
nor U1680 (N_1680,N_1127,N_1059);
nor U1681 (N_1681,N_1409,N_1176);
and U1682 (N_1682,N_1478,N_1012);
and U1683 (N_1683,N_1128,N_1457);
nand U1684 (N_1684,N_1135,N_1158);
or U1685 (N_1685,N_1465,N_1278);
or U1686 (N_1686,N_1206,N_1468);
xor U1687 (N_1687,N_1446,N_1397);
and U1688 (N_1688,N_1423,N_1108);
or U1689 (N_1689,N_1189,N_1390);
or U1690 (N_1690,N_1099,N_1203);
and U1691 (N_1691,N_1445,N_1257);
nor U1692 (N_1692,N_1060,N_1007);
xnor U1693 (N_1693,N_1262,N_1267);
nand U1694 (N_1694,N_1132,N_1055);
and U1695 (N_1695,N_1201,N_1341);
xor U1696 (N_1696,N_1453,N_1361);
nor U1697 (N_1697,N_1137,N_1437);
nor U1698 (N_1698,N_1300,N_1030);
nand U1699 (N_1699,N_1080,N_1053);
nor U1700 (N_1700,N_1302,N_1150);
xor U1701 (N_1701,N_1266,N_1029);
nand U1702 (N_1702,N_1088,N_1464);
and U1703 (N_1703,N_1101,N_1462);
nand U1704 (N_1704,N_1057,N_1040);
nor U1705 (N_1705,N_1120,N_1471);
nor U1706 (N_1706,N_1111,N_1241);
and U1707 (N_1707,N_1083,N_1422);
xor U1708 (N_1708,N_1064,N_1177);
and U1709 (N_1709,N_1159,N_1147);
xor U1710 (N_1710,N_1216,N_1031);
xnor U1711 (N_1711,N_1489,N_1395);
and U1712 (N_1712,N_1043,N_1050);
xnor U1713 (N_1713,N_1398,N_1103);
nand U1714 (N_1714,N_1329,N_1298);
and U1715 (N_1715,N_1400,N_1369);
xor U1716 (N_1716,N_1366,N_1441);
and U1717 (N_1717,N_1109,N_1224);
xor U1718 (N_1718,N_1145,N_1330);
nand U1719 (N_1719,N_1069,N_1130);
xor U1720 (N_1720,N_1204,N_1155);
nor U1721 (N_1721,N_1286,N_1046);
nor U1722 (N_1722,N_1419,N_1106);
nand U1723 (N_1723,N_1326,N_1098);
nand U1724 (N_1724,N_1436,N_1303);
nand U1725 (N_1725,N_1011,N_1010);
xnor U1726 (N_1726,N_1432,N_1376);
or U1727 (N_1727,N_1193,N_1034);
nand U1728 (N_1728,N_1153,N_1168);
and U1729 (N_1729,N_1459,N_1485);
and U1730 (N_1730,N_1246,N_1233);
xnor U1731 (N_1731,N_1116,N_1288);
nand U1732 (N_1732,N_1205,N_1295);
or U1733 (N_1733,N_1092,N_1477);
and U1734 (N_1734,N_1136,N_1027);
and U1735 (N_1735,N_1318,N_1392);
nor U1736 (N_1736,N_1381,N_1352);
nor U1737 (N_1737,N_1068,N_1202);
nand U1738 (N_1738,N_1015,N_1306);
and U1739 (N_1739,N_1438,N_1227);
xor U1740 (N_1740,N_1377,N_1265);
xnor U1741 (N_1741,N_1325,N_1460);
or U1742 (N_1742,N_1134,N_1480);
and U1743 (N_1743,N_1339,N_1016);
nand U1744 (N_1744,N_1244,N_1234);
nand U1745 (N_1745,N_1455,N_1018);
nor U1746 (N_1746,N_1396,N_1479);
nand U1747 (N_1747,N_1324,N_1035);
or U1748 (N_1748,N_1190,N_1420);
nand U1749 (N_1749,N_1138,N_1322);
nor U1750 (N_1750,N_1362,N_1062);
or U1751 (N_1751,N_1437,N_1380);
nand U1752 (N_1752,N_1095,N_1421);
nand U1753 (N_1753,N_1103,N_1282);
nand U1754 (N_1754,N_1402,N_1308);
nor U1755 (N_1755,N_1287,N_1174);
nor U1756 (N_1756,N_1283,N_1425);
and U1757 (N_1757,N_1372,N_1175);
and U1758 (N_1758,N_1188,N_1382);
and U1759 (N_1759,N_1441,N_1415);
nor U1760 (N_1760,N_1498,N_1469);
nand U1761 (N_1761,N_1210,N_1481);
xor U1762 (N_1762,N_1183,N_1292);
nor U1763 (N_1763,N_1422,N_1138);
nor U1764 (N_1764,N_1294,N_1385);
xor U1765 (N_1765,N_1449,N_1417);
nor U1766 (N_1766,N_1308,N_1454);
nand U1767 (N_1767,N_1015,N_1093);
nor U1768 (N_1768,N_1403,N_1103);
nand U1769 (N_1769,N_1424,N_1278);
nand U1770 (N_1770,N_1499,N_1314);
and U1771 (N_1771,N_1374,N_1225);
xnor U1772 (N_1772,N_1035,N_1458);
and U1773 (N_1773,N_1221,N_1498);
and U1774 (N_1774,N_1049,N_1416);
nand U1775 (N_1775,N_1275,N_1460);
xnor U1776 (N_1776,N_1162,N_1201);
xnor U1777 (N_1777,N_1343,N_1233);
nor U1778 (N_1778,N_1165,N_1034);
nor U1779 (N_1779,N_1448,N_1274);
and U1780 (N_1780,N_1124,N_1200);
nor U1781 (N_1781,N_1262,N_1013);
xor U1782 (N_1782,N_1040,N_1073);
nand U1783 (N_1783,N_1215,N_1191);
and U1784 (N_1784,N_1184,N_1430);
nand U1785 (N_1785,N_1226,N_1280);
and U1786 (N_1786,N_1128,N_1420);
or U1787 (N_1787,N_1483,N_1096);
and U1788 (N_1788,N_1363,N_1144);
nor U1789 (N_1789,N_1144,N_1045);
nor U1790 (N_1790,N_1138,N_1461);
and U1791 (N_1791,N_1085,N_1462);
nor U1792 (N_1792,N_1366,N_1257);
or U1793 (N_1793,N_1377,N_1472);
or U1794 (N_1794,N_1086,N_1089);
and U1795 (N_1795,N_1004,N_1394);
nand U1796 (N_1796,N_1304,N_1261);
nor U1797 (N_1797,N_1357,N_1242);
nand U1798 (N_1798,N_1352,N_1407);
xnor U1799 (N_1799,N_1034,N_1355);
or U1800 (N_1800,N_1237,N_1057);
nand U1801 (N_1801,N_1358,N_1288);
nor U1802 (N_1802,N_1193,N_1499);
xnor U1803 (N_1803,N_1172,N_1495);
xor U1804 (N_1804,N_1099,N_1360);
or U1805 (N_1805,N_1271,N_1232);
nand U1806 (N_1806,N_1110,N_1060);
or U1807 (N_1807,N_1077,N_1305);
or U1808 (N_1808,N_1262,N_1007);
nor U1809 (N_1809,N_1028,N_1391);
and U1810 (N_1810,N_1296,N_1080);
nand U1811 (N_1811,N_1468,N_1358);
nand U1812 (N_1812,N_1162,N_1420);
xnor U1813 (N_1813,N_1255,N_1356);
nor U1814 (N_1814,N_1101,N_1180);
and U1815 (N_1815,N_1251,N_1135);
and U1816 (N_1816,N_1109,N_1443);
and U1817 (N_1817,N_1329,N_1020);
xnor U1818 (N_1818,N_1259,N_1223);
nand U1819 (N_1819,N_1341,N_1227);
or U1820 (N_1820,N_1469,N_1038);
and U1821 (N_1821,N_1278,N_1499);
nand U1822 (N_1822,N_1112,N_1295);
or U1823 (N_1823,N_1397,N_1047);
xor U1824 (N_1824,N_1021,N_1034);
nand U1825 (N_1825,N_1082,N_1018);
nand U1826 (N_1826,N_1123,N_1467);
xor U1827 (N_1827,N_1284,N_1151);
and U1828 (N_1828,N_1154,N_1187);
and U1829 (N_1829,N_1109,N_1314);
and U1830 (N_1830,N_1408,N_1295);
or U1831 (N_1831,N_1117,N_1296);
or U1832 (N_1832,N_1110,N_1428);
nand U1833 (N_1833,N_1469,N_1035);
nor U1834 (N_1834,N_1447,N_1275);
or U1835 (N_1835,N_1344,N_1169);
and U1836 (N_1836,N_1384,N_1452);
or U1837 (N_1837,N_1256,N_1412);
or U1838 (N_1838,N_1072,N_1452);
nand U1839 (N_1839,N_1399,N_1193);
xnor U1840 (N_1840,N_1118,N_1169);
xor U1841 (N_1841,N_1390,N_1238);
or U1842 (N_1842,N_1383,N_1074);
nand U1843 (N_1843,N_1201,N_1277);
and U1844 (N_1844,N_1213,N_1327);
xnor U1845 (N_1845,N_1208,N_1131);
nor U1846 (N_1846,N_1495,N_1174);
or U1847 (N_1847,N_1087,N_1166);
xnor U1848 (N_1848,N_1209,N_1420);
and U1849 (N_1849,N_1484,N_1113);
nand U1850 (N_1850,N_1307,N_1378);
xnor U1851 (N_1851,N_1462,N_1421);
and U1852 (N_1852,N_1397,N_1110);
nor U1853 (N_1853,N_1488,N_1231);
nor U1854 (N_1854,N_1239,N_1330);
nor U1855 (N_1855,N_1383,N_1055);
nand U1856 (N_1856,N_1485,N_1390);
xor U1857 (N_1857,N_1236,N_1139);
or U1858 (N_1858,N_1247,N_1335);
xnor U1859 (N_1859,N_1328,N_1416);
nor U1860 (N_1860,N_1361,N_1364);
or U1861 (N_1861,N_1473,N_1133);
or U1862 (N_1862,N_1103,N_1007);
or U1863 (N_1863,N_1437,N_1478);
xnor U1864 (N_1864,N_1252,N_1074);
xor U1865 (N_1865,N_1380,N_1314);
nand U1866 (N_1866,N_1182,N_1307);
and U1867 (N_1867,N_1151,N_1388);
and U1868 (N_1868,N_1002,N_1490);
nor U1869 (N_1869,N_1379,N_1237);
xor U1870 (N_1870,N_1072,N_1308);
and U1871 (N_1871,N_1211,N_1388);
and U1872 (N_1872,N_1053,N_1132);
and U1873 (N_1873,N_1326,N_1016);
xor U1874 (N_1874,N_1235,N_1085);
and U1875 (N_1875,N_1290,N_1469);
nor U1876 (N_1876,N_1226,N_1256);
or U1877 (N_1877,N_1169,N_1144);
xnor U1878 (N_1878,N_1260,N_1110);
nand U1879 (N_1879,N_1252,N_1034);
nand U1880 (N_1880,N_1024,N_1340);
xor U1881 (N_1881,N_1439,N_1019);
nand U1882 (N_1882,N_1460,N_1344);
nor U1883 (N_1883,N_1427,N_1265);
or U1884 (N_1884,N_1230,N_1108);
xnor U1885 (N_1885,N_1309,N_1162);
xnor U1886 (N_1886,N_1170,N_1205);
nand U1887 (N_1887,N_1001,N_1197);
nor U1888 (N_1888,N_1315,N_1438);
and U1889 (N_1889,N_1326,N_1341);
nand U1890 (N_1890,N_1246,N_1157);
nor U1891 (N_1891,N_1455,N_1280);
xnor U1892 (N_1892,N_1161,N_1129);
nand U1893 (N_1893,N_1093,N_1487);
nor U1894 (N_1894,N_1116,N_1089);
nor U1895 (N_1895,N_1281,N_1071);
nor U1896 (N_1896,N_1134,N_1013);
xor U1897 (N_1897,N_1392,N_1476);
and U1898 (N_1898,N_1020,N_1220);
or U1899 (N_1899,N_1271,N_1292);
or U1900 (N_1900,N_1223,N_1072);
nand U1901 (N_1901,N_1316,N_1205);
nor U1902 (N_1902,N_1465,N_1041);
and U1903 (N_1903,N_1351,N_1345);
xnor U1904 (N_1904,N_1370,N_1130);
nand U1905 (N_1905,N_1090,N_1330);
nand U1906 (N_1906,N_1321,N_1470);
xnor U1907 (N_1907,N_1437,N_1025);
nor U1908 (N_1908,N_1424,N_1498);
and U1909 (N_1909,N_1015,N_1494);
xnor U1910 (N_1910,N_1082,N_1302);
or U1911 (N_1911,N_1274,N_1333);
and U1912 (N_1912,N_1359,N_1038);
or U1913 (N_1913,N_1493,N_1182);
and U1914 (N_1914,N_1210,N_1234);
nand U1915 (N_1915,N_1094,N_1267);
nand U1916 (N_1916,N_1129,N_1215);
and U1917 (N_1917,N_1336,N_1408);
or U1918 (N_1918,N_1407,N_1134);
nor U1919 (N_1919,N_1183,N_1236);
and U1920 (N_1920,N_1060,N_1127);
or U1921 (N_1921,N_1482,N_1305);
nor U1922 (N_1922,N_1463,N_1227);
or U1923 (N_1923,N_1191,N_1421);
nand U1924 (N_1924,N_1270,N_1433);
xor U1925 (N_1925,N_1487,N_1373);
xnor U1926 (N_1926,N_1091,N_1154);
or U1927 (N_1927,N_1301,N_1324);
nor U1928 (N_1928,N_1407,N_1055);
xor U1929 (N_1929,N_1487,N_1201);
nand U1930 (N_1930,N_1354,N_1175);
nand U1931 (N_1931,N_1479,N_1327);
nand U1932 (N_1932,N_1197,N_1065);
or U1933 (N_1933,N_1241,N_1221);
xor U1934 (N_1934,N_1188,N_1112);
xor U1935 (N_1935,N_1283,N_1144);
nand U1936 (N_1936,N_1121,N_1347);
and U1937 (N_1937,N_1305,N_1172);
xnor U1938 (N_1938,N_1499,N_1445);
or U1939 (N_1939,N_1236,N_1318);
nand U1940 (N_1940,N_1240,N_1188);
or U1941 (N_1941,N_1421,N_1196);
xnor U1942 (N_1942,N_1306,N_1422);
nor U1943 (N_1943,N_1055,N_1482);
and U1944 (N_1944,N_1225,N_1186);
nor U1945 (N_1945,N_1383,N_1416);
nor U1946 (N_1946,N_1367,N_1103);
or U1947 (N_1947,N_1320,N_1051);
nand U1948 (N_1948,N_1368,N_1338);
nand U1949 (N_1949,N_1140,N_1215);
or U1950 (N_1950,N_1307,N_1274);
or U1951 (N_1951,N_1010,N_1205);
nand U1952 (N_1952,N_1322,N_1169);
xnor U1953 (N_1953,N_1447,N_1395);
or U1954 (N_1954,N_1246,N_1448);
or U1955 (N_1955,N_1374,N_1130);
and U1956 (N_1956,N_1192,N_1413);
nand U1957 (N_1957,N_1065,N_1027);
and U1958 (N_1958,N_1273,N_1479);
or U1959 (N_1959,N_1137,N_1212);
and U1960 (N_1960,N_1004,N_1214);
and U1961 (N_1961,N_1180,N_1389);
nand U1962 (N_1962,N_1159,N_1364);
and U1963 (N_1963,N_1488,N_1460);
and U1964 (N_1964,N_1026,N_1190);
and U1965 (N_1965,N_1203,N_1102);
xnor U1966 (N_1966,N_1359,N_1022);
or U1967 (N_1967,N_1452,N_1439);
xor U1968 (N_1968,N_1359,N_1307);
nor U1969 (N_1969,N_1098,N_1280);
xnor U1970 (N_1970,N_1183,N_1261);
and U1971 (N_1971,N_1148,N_1498);
nor U1972 (N_1972,N_1249,N_1111);
xnor U1973 (N_1973,N_1374,N_1099);
xor U1974 (N_1974,N_1066,N_1213);
or U1975 (N_1975,N_1255,N_1142);
nor U1976 (N_1976,N_1469,N_1326);
and U1977 (N_1977,N_1266,N_1298);
or U1978 (N_1978,N_1020,N_1256);
xnor U1979 (N_1979,N_1154,N_1277);
xor U1980 (N_1980,N_1120,N_1025);
nor U1981 (N_1981,N_1082,N_1246);
or U1982 (N_1982,N_1091,N_1015);
nor U1983 (N_1983,N_1339,N_1479);
nand U1984 (N_1984,N_1046,N_1064);
or U1985 (N_1985,N_1289,N_1491);
nand U1986 (N_1986,N_1154,N_1203);
nor U1987 (N_1987,N_1302,N_1309);
or U1988 (N_1988,N_1273,N_1165);
nand U1989 (N_1989,N_1418,N_1125);
nor U1990 (N_1990,N_1419,N_1163);
and U1991 (N_1991,N_1264,N_1134);
xor U1992 (N_1992,N_1405,N_1336);
and U1993 (N_1993,N_1339,N_1336);
xor U1994 (N_1994,N_1125,N_1142);
or U1995 (N_1995,N_1268,N_1033);
and U1996 (N_1996,N_1248,N_1270);
or U1997 (N_1997,N_1187,N_1337);
nand U1998 (N_1998,N_1243,N_1459);
xnor U1999 (N_1999,N_1235,N_1409);
nand U2000 (N_2000,N_1968,N_1581);
nand U2001 (N_2001,N_1669,N_1576);
nor U2002 (N_2002,N_1998,N_1686);
and U2003 (N_2003,N_1894,N_1935);
or U2004 (N_2004,N_1712,N_1947);
and U2005 (N_2005,N_1824,N_1967);
nand U2006 (N_2006,N_1898,N_1795);
and U2007 (N_2007,N_1932,N_1509);
nor U2008 (N_2008,N_1612,N_1508);
nor U2009 (N_2009,N_1610,N_1505);
or U2010 (N_2010,N_1873,N_1806);
or U2011 (N_2011,N_1684,N_1830);
nor U2012 (N_2012,N_1865,N_1924);
and U2013 (N_2013,N_1648,N_1845);
nor U2014 (N_2014,N_1903,N_1628);
and U2015 (N_2015,N_1640,N_1578);
nand U2016 (N_2016,N_1861,N_1737);
or U2017 (N_2017,N_1966,N_1887);
xor U2018 (N_2018,N_1604,N_1811);
nor U2019 (N_2019,N_1881,N_1981);
nand U2020 (N_2020,N_1750,N_1707);
and U2021 (N_2021,N_1674,N_1758);
nand U2022 (N_2022,N_1635,N_1999);
xnor U2023 (N_2023,N_1848,N_1683);
xnor U2024 (N_2024,N_1961,N_1632);
nand U2025 (N_2025,N_1788,N_1697);
nor U2026 (N_2026,N_1975,N_1766);
nand U2027 (N_2027,N_1859,N_1982);
nand U2028 (N_2028,N_1643,N_1516);
nor U2029 (N_2029,N_1700,N_1690);
and U2030 (N_2030,N_1876,N_1936);
nand U2031 (N_2031,N_1971,N_1799);
or U2032 (N_2032,N_1779,N_1759);
or U2033 (N_2033,N_1741,N_1634);
nor U2034 (N_2034,N_1528,N_1921);
or U2035 (N_2035,N_1960,N_1535);
and U2036 (N_2036,N_1626,N_1621);
nand U2037 (N_2037,N_1794,N_1668);
and U2038 (N_2038,N_1980,N_1653);
nand U2039 (N_2039,N_1776,N_1571);
or U2040 (N_2040,N_1720,N_1679);
nor U2041 (N_2041,N_1948,N_1841);
and U2042 (N_2042,N_1711,N_1771);
nor U2043 (N_2043,N_1895,N_1785);
xor U2044 (N_2044,N_1792,N_1600);
or U2045 (N_2045,N_1883,N_1807);
and U2046 (N_2046,N_1905,N_1702);
nor U2047 (N_2047,N_1694,N_1805);
and U2048 (N_2048,N_1959,N_1602);
nand U2049 (N_2049,N_1606,N_1951);
and U2050 (N_2050,N_1540,N_1914);
nand U2051 (N_2051,N_1970,N_1527);
or U2052 (N_2052,N_1793,N_1593);
or U2053 (N_2053,N_1941,N_1732);
and U2054 (N_2054,N_1617,N_1531);
or U2055 (N_2055,N_1662,N_1911);
xnor U2056 (N_2056,N_1767,N_1624);
or U2057 (N_2057,N_1687,N_1716);
or U2058 (N_2058,N_1726,N_1658);
xnor U2059 (N_2059,N_1644,N_1995);
nor U2060 (N_2060,N_1688,N_1676);
nand U2061 (N_2061,N_1820,N_1920);
nand U2062 (N_2062,N_1693,N_1659);
nor U2063 (N_2063,N_1666,N_1570);
or U2064 (N_2064,N_1500,N_1558);
nand U2065 (N_2065,N_1917,N_1762);
xor U2066 (N_2066,N_1844,N_1990);
nor U2067 (N_2067,N_1928,N_1614);
nand U2068 (N_2068,N_1955,N_1543);
nand U2069 (N_2069,N_1577,N_1969);
and U2070 (N_2070,N_1585,N_1681);
and U2071 (N_2071,N_1885,N_1862);
nand U2072 (N_2072,N_1596,N_1986);
nand U2073 (N_2073,N_1850,N_1703);
xor U2074 (N_2074,N_1625,N_1976);
xnor U2075 (N_2075,N_1709,N_1560);
nand U2076 (N_2076,N_1651,N_1934);
and U2077 (N_2077,N_1818,N_1912);
nand U2078 (N_2078,N_1890,N_1782);
xnor U2079 (N_2079,N_1569,N_1812);
or U2080 (N_2080,N_1665,N_1546);
xor U2081 (N_2081,N_1944,N_1773);
or U2082 (N_2082,N_1704,N_1991);
or U2083 (N_2083,N_1564,N_1699);
nor U2084 (N_2084,N_1534,N_1705);
and U2085 (N_2085,N_1708,N_1670);
nand U2086 (N_2086,N_1797,N_1927);
and U2087 (N_2087,N_1598,N_1728);
nor U2088 (N_2088,N_1958,N_1992);
xor U2089 (N_2089,N_1926,N_1591);
nand U2090 (N_2090,N_1838,N_1538);
and U2091 (N_2091,N_1647,N_1733);
xnor U2092 (N_2092,N_1725,N_1754);
or U2093 (N_2093,N_1671,N_1770);
or U2094 (N_2094,N_1846,N_1518);
or U2095 (N_2095,N_1918,N_1520);
xnor U2096 (N_2096,N_1663,N_1553);
nand U2097 (N_2097,N_1816,N_1633);
nor U2098 (N_2098,N_1523,N_1541);
or U2099 (N_2099,N_1855,N_1983);
xor U2100 (N_2100,N_1768,N_1680);
nand U2101 (N_2101,N_1605,N_1871);
and U2102 (N_2102,N_1764,N_1809);
or U2103 (N_2103,N_1719,N_1512);
nor U2104 (N_2104,N_1526,N_1774);
or U2105 (N_2105,N_1965,N_1682);
and U2106 (N_2106,N_1909,N_1837);
or U2107 (N_2107,N_1867,N_1775);
or U2108 (N_2108,N_1532,N_1957);
nor U2109 (N_2109,N_1645,N_1763);
nor U2110 (N_2110,N_1889,N_1777);
and U2111 (N_2111,N_1599,N_1756);
and U2112 (N_2112,N_1563,N_1833);
nand U2113 (N_2113,N_1667,N_1989);
nor U2114 (N_2114,N_1696,N_1575);
nor U2115 (N_2115,N_1622,N_1603);
nand U2116 (N_2116,N_1555,N_1580);
nor U2117 (N_2117,N_1721,N_1650);
xor U2118 (N_2118,N_1620,N_1973);
and U2119 (N_2119,N_1907,N_1502);
xor U2120 (N_2120,N_1521,N_1542);
and U2121 (N_2121,N_1878,N_1790);
nand U2122 (N_2122,N_1778,N_1803);
and U2123 (N_2123,N_1589,N_1977);
nor U2124 (N_2124,N_1748,N_1916);
and U2125 (N_2125,N_1829,N_1601);
xor U2126 (N_2126,N_1590,N_1853);
nand U2127 (N_2127,N_1689,N_1942);
or U2128 (N_2128,N_1910,N_1529);
nand U2129 (N_2129,N_1884,N_1945);
or U2130 (N_2130,N_1565,N_1723);
and U2131 (N_2131,N_1893,N_1616);
xnor U2132 (N_2132,N_1586,N_1828);
and U2133 (N_2133,N_1874,N_1559);
xnor U2134 (N_2134,N_1840,N_1706);
nand U2135 (N_2135,N_1956,N_1677);
or U2136 (N_2136,N_1718,N_1963);
xor U2137 (N_2137,N_1835,N_1537);
and U2138 (N_2138,N_1739,N_1722);
nand U2139 (N_2139,N_1854,N_1557);
xor U2140 (N_2140,N_1937,N_1849);
nor U2141 (N_2141,N_1742,N_1655);
nand U2142 (N_2142,N_1888,N_1801);
xnor U2143 (N_2143,N_1556,N_1631);
and U2144 (N_2144,N_1933,N_1548);
and U2145 (N_2145,N_1673,N_1525);
nor U2146 (N_2146,N_1760,N_1827);
and U2147 (N_2147,N_1734,N_1765);
xnor U2148 (N_2148,N_1636,N_1901);
nor U2149 (N_2149,N_1710,N_1660);
xor U2150 (N_2150,N_1730,N_1925);
xnor U2151 (N_2151,N_1780,N_1875);
or U2152 (N_2152,N_1772,N_1761);
and U2153 (N_2153,N_1781,N_1654);
xnor U2154 (N_2154,N_1988,N_1836);
nor U2155 (N_2155,N_1545,N_1646);
and U2156 (N_2156,N_1698,N_1842);
xor U2157 (N_2157,N_1847,N_1514);
or U2158 (N_2158,N_1630,N_1568);
xor U2159 (N_2159,N_1791,N_1691);
and U2160 (N_2160,N_1996,N_1783);
nor U2161 (N_2161,N_1952,N_1784);
nor U2162 (N_2162,N_1810,N_1607);
nand U2163 (N_2163,N_1796,N_1929);
nand U2164 (N_2164,N_1738,N_1597);
and U2165 (N_2165,N_1856,N_1804);
nor U2166 (N_2166,N_1819,N_1954);
xor U2167 (N_2167,N_1745,N_1552);
nor U2168 (N_2168,N_1979,N_1930);
and U2169 (N_2169,N_1753,N_1611);
nand U2170 (N_2170,N_1735,N_1972);
xnor U2171 (N_2171,N_1997,N_1913);
xnor U2172 (N_2172,N_1870,N_1817);
nor U2173 (N_2173,N_1993,N_1619);
nor U2174 (N_2174,N_1752,N_1579);
nand U2175 (N_2175,N_1949,N_1510);
and U2176 (N_2176,N_1814,N_1714);
or U2177 (N_2177,N_1931,N_1869);
xnor U2178 (N_2178,N_1744,N_1536);
xnor U2179 (N_2179,N_1550,N_1641);
xor U2180 (N_2180,N_1609,N_1615);
nor U2181 (N_2181,N_1573,N_1815);
nand U2182 (N_2182,N_1896,N_1902);
nand U2183 (N_2183,N_1638,N_1897);
nor U2184 (N_2184,N_1715,N_1751);
nand U2185 (N_2185,N_1639,N_1595);
or U2186 (N_2186,N_1839,N_1857);
nor U2187 (N_2187,N_1826,N_1656);
nand U2188 (N_2188,N_1872,N_1922);
nand U2189 (N_2189,N_1623,N_1749);
and U2190 (N_2190,N_1740,N_1900);
nor U2191 (N_2191,N_1747,N_1724);
nand U2192 (N_2192,N_1940,N_1994);
xnor U2193 (N_2193,N_1798,N_1561);
and U2194 (N_2194,N_1892,N_1821);
nand U2195 (N_2195,N_1554,N_1964);
and U2196 (N_2196,N_1562,N_1637);
and U2197 (N_2197,N_1675,N_1915);
nand U2198 (N_2198,N_1822,N_1939);
or U2199 (N_2199,N_1868,N_1904);
and U2200 (N_2200,N_1789,N_1517);
or U2201 (N_2201,N_1544,N_1831);
or U2202 (N_2202,N_1506,N_1962);
nand U2203 (N_2203,N_1880,N_1757);
xor U2204 (N_2204,N_1943,N_1787);
nand U2205 (N_2205,N_1627,N_1974);
nand U2206 (N_2206,N_1701,N_1524);
nor U2207 (N_2207,N_1672,N_1882);
and U2208 (N_2208,N_1608,N_1566);
and U2209 (N_2209,N_1588,N_1522);
and U2210 (N_2210,N_1729,N_1583);
nor U2211 (N_2211,N_1985,N_1551);
nor U2212 (N_2212,N_1825,N_1584);
nand U2213 (N_2213,N_1899,N_1695);
xnor U2214 (N_2214,N_1717,N_1938);
xor U2215 (N_2215,N_1519,N_1755);
nor U2216 (N_2216,N_1727,N_1864);
nor U2217 (N_2217,N_1592,N_1800);
or U2218 (N_2218,N_1919,N_1832);
or U2219 (N_2219,N_1908,N_1978);
or U2220 (N_2220,N_1692,N_1511);
nand U2221 (N_2221,N_1642,N_1731);
and U2222 (N_2222,N_1736,N_1549);
or U2223 (N_2223,N_1906,N_1594);
xnor U2224 (N_2224,N_1504,N_1533);
xor U2225 (N_2225,N_1501,N_1678);
xnor U2226 (N_2226,N_1946,N_1574);
or U2227 (N_2227,N_1743,N_1852);
xor U2228 (N_2228,N_1851,N_1507);
xor U2229 (N_2229,N_1891,N_1572);
or U2230 (N_2230,N_1858,N_1652);
or U2231 (N_2231,N_1713,N_1567);
xnor U2232 (N_2232,N_1834,N_1547);
nand U2233 (N_2233,N_1530,N_1613);
xor U2234 (N_2234,N_1582,N_1587);
nor U2235 (N_2235,N_1813,N_1769);
nor U2236 (N_2236,N_1808,N_1823);
nand U2237 (N_2237,N_1629,N_1860);
nor U2238 (N_2238,N_1984,N_1539);
and U2239 (N_2239,N_1886,N_1802);
nor U2240 (N_2240,N_1661,N_1649);
and U2241 (N_2241,N_1879,N_1877);
and U2242 (N_2242,N_1746,N_1950);
or U2243 (N_2243,N_1863,N_1923);
and U2244 (N_2244,N_1866,N_1513);
and U2245 (N_2245,N_1664,N_1685);
xnor U2246 (N_2246,N_1515,N_1618);
or U2247 (N_2247,N_1786,N_1657);
and U2248 (N_2248,N_1953,N_1843);
nor U2249 (N_2249,N_1503,N_1987);
and U2250 (N_2250,N_1968,N_1660);
nand U2251 (N_2251,N_1651,N_1657);
nor U2252 (N_2252,N_1582,N_1717);
nand U2253 (N_2253,N_1779,N_1693);
nand U2254 (N_2254,N_1744,N_1975);
xor U2255 (N_2255,N_1625,N_1629);
nor U2256 (N_2256,N_1537,N_1729);
nor U2257 (N_2257,N_1960,N_1821);
nand U2258 (N_2258,N_1711,N_1684);
nand U2259 (N_2259,N_1986,N_1676);
nand U2260 (N_2260,N_1603,N_1666);
or U2261 (N_2261,N_1924,N_1601);
nor U2262 (N_2262,N_1663,N_1608);
xor U2263 (N_2263,N_1789,N_1741);
xnor U2264 (N_2264,N_1655,N_1941);
nor U2265 (N_2265,N_1642,N_1563);
and U2266 (N_2266,N_1949,N_1981);
or U2267 (N_2267,N_1592,N_1859);
and U2268 (N_2268,N_1731,N_1734);
or U2269 (N_2269,N_1834,N_1518);
xor U2270 (N_2270,N_1739,N_1617);
and U2271 (N_2271,N_1807,N_1826);
or U2272 (N_2272,N_1553,N_1675);
or U2273 (N_2273,N_1928,N_1545);
or U2274 (N_2274,N_1675,N_1749);
xor U2275 (N_2275,N_1774,N_1569);
nor U2276 (N_2276,N_1502,N_1638);
or U2277 (N_2277,N_1533,N_1923);
and U2278 (N_2278,N_1976,N_1742);
and U2279 (N_2279,N_1528,N_1855);
xnor U2280 (N_2280,N_1718,N_1512);
or U2281 (N_2281,N_1635,N_1551);
xor U2282 (N_2282,N_1607,N_1549);
nor U2283 (N_2283,N_1801,N_1855);
xnor U2284 (N_2284,N_1574,N_1971);
xnor U2285 (N_2285,N_1621,N_1681);
xnor U2286 (N_2286,N_1555,N_1805);
or U2287 (N_2287,N_1933,N_1685);
and U2288 (N_2288,N_1634,N_1942);
nor U2289 (N_2289,N_1548,N_1533);
xor U2290 (N_2290,N_1681,N_1884);
xor U2291 (N_2291,N_1655,N_1991);
xnor U2292 (N_2292,N_1660,N_1618);
and U2293 (N_2293,N_1839,N_1958);
xor U2294 (N_2294,N_1959,N_1983);
nor U2295 (N_2295,N_1998,N_1828);
xor U2296 (N_2296,N_1974,N_1937);
or U2297 (N_2297,N_1638,N_1514);
and U2298 (N_2298,N_1734,N_1538);
nor U2299 (N_2299,N_1945,N_1709);
or U2300 (N_2300,N_1960,N_1766);
nor U2301 (N_2301,N_1997,N_1971);
or U2302 (N_2302,N_1846,N_1702);
and U2303 (N_2303,N_1749,N_1621);
and U2304 (N_2304,N_1786,N_1573);
nand U2305 (N_2305,N_1709,N_1881);
and U2306 (N_2306,N_1818,N_1655);
or U2307 (N_2307,N_1871,N_1683);
or U2308 (N_2308,N_1599,N_1881);
or U2309 (N_2309,N_1586,N_1917);
xnor U2310 (N_2310,N_1930,N_1847);
or U2311 (N_2311,N_1962,N_1635);
and U2312 (N_2312,N_1971,N_1916);
or U2313 (N_2313,N_1911,N_1539);
or U2314 (N_2314,N_1622,N_1910);
xnor U2315 (N_2315,N_1505,N_1656);
or U2316 (N_2316,N_1806,N_1755);
or U2317 (N_2317,N_1677,N_1970);
and U2318 (N_2318,N_1573,N_1707);
nand U2319 (N_2319,N_1739,N_1639);
or U2320 (N_2320,N_1716,N_1983);
nor U2321 (N_2321,N_1721,N_1987);
and U2322 (N_2322,N_1907,N_1587);
or U2323 (N_2323,N_1902,N_1653);
or U2324 (N_2324,N_1805,N_1894);
or U2325 (N_2325,N_1913,N_1530);
nor U2326 (N_2326,N_1776,N_1943);
and U2327 (N_2327,N_1826,N_1571);
and U2328 (N_2328,N_1711,N_1977);
nand U2329 (N_2329,N_1566,N_1960);
xor U2330 (N_2330,N_1948,N_1727);
xnor U2331 (N_2331,N_1973,N_1711);
or U2332 (N_2332,N_1627,N_1923);
and U2333 (N_2333,N_1695,N_1590);
or U2334 (N_2334,N_1887,N_1929);
xnor U2335 (N_2335,N_1894,N_1763);
nor U2336 (N_2336,N_1678,N_1888);
and U2337 (N_2337,N_1737,N_1690);
nand U2338 (N_2338,N_1678,N_1902);
or U2339 (N_2339,N_1765,N_1565);
xnor U2340 (N_2340,N_1615,N_1835);
xnor U2341 (N_2341,N_1617,N_1832);
and U2342 (N_2342,N_1856,N_1879);
nor U2343 (N_2343,N_1666,N_1778);
nand U2344 (N_2344,N_1778,N_1553);
nand U2345 (N_2345,N_1768,N_1764);
nand U2346 (N_2346,N_1509,N_1856);
nand U2347 (N_2347,N_1970,N_1650);
or U2348 (N_2348,N_1566,N_1915);
and U2349 (N_2349,N_1874,N_1887);
xnor U2350 (N_2350,N_1906,N_1823);
xnor U2351 (N_2351,N_1863,N_1892);
nor U2352 (N_2352,N_1859,N_1961);
nor U2353 (N_2353,N_1981,N_1603);
nor U2354 (N_2354,N_1609,N_1671);
nor U2355 (N_2355,N_1809,N_1881);
nor U2356 (N_2356,N_1804,N_1576);
xor U2357 (N_2357,N_1510,N_1680);
xor U2358 (N_2358,N_1784,N_1575);
and U2359 (N_2359,N_1620,N_1688);
xor U2360 (N_2360,N_1852,N_1920);
or U2361 (N_2361,N_1561,N_1751);
nand U2362 (N_2362,N_1533,N_1557);
or U2363 (N_2363,N_1740,N_1582);
nand U2364 (N_2364,N_1793,N_1931);
nand U2365 (N_2365,N_1775,N_1641);
and U2366 (N_2366,N_1665,N_1503);
xor U2367 (N_2367,N_1612,N_1872);
or U2368 (N_2368,N_1861,N_1759);
and U2369 (N_2369,N_1592,N_1656);
and U2370 (N_2370,N_1939,N_1998);
xnor U2371 (N_2371,N_1711,N_1567);
or U2372 (N_2372,N_1951,N_1676);
and U2373 (N_2373,N_1565,N_1585);
and U2374 (N_2374,N_1530,N_1849);
xnor U2375 (N_2375,N_1901,N_1559);
and U2376 (N_2376,N_1809,N_1725);
xnor U2377 (N_2377,N_1964,N_1841);
or U2378 (N_2378,N_1661,N_1785);
nand U2379 (N_2379,N_1754,N_1927);
xor U2380 (N_2380,N_1798,N_1652);
or U2381 (N_2381,N_1578,N_1804);
nor U2382 (N_2382,N_1972,N_1668);
nand U2383 (N_2383,N_1541,N_1695);
and U2384 (N_2384,N_1594,N_1645);
or U2385 (N_2385,N_1658,N_1524);
xnor U2386 (N_2386,N_1894,N_1655);
or U2387 (N_2387,N_1551,N_1664);
nor U2388 (N_2388,N_1686,N_1931);
or U2389 (N_2389,N_1551,N_1834);
nand U2390 (N_2390,N_1536,N_1877);
and U2391 (N_2391,N_1949,N_1688);
and U2392 (N_2392,N_1868,N_1771);
or U2393 (N_2393,N_1938,N_1548);
and U2394 (N_2394,N_1960,N_1869);
xor U2395 (N_2395,N_1681,N_1537);
or U2396 (N_2396,N_1822,N_1634);
nor U2397 (N_2397,N_1575,N_1500);
nor U2398 (N_2398,N_1671,N_1694);
and U2399 (N_2399,N_1586,N_1549);
xor U2400 (N_2400,N_1967,N_1756);
xor U2401 (N_2401,N_1523,N_1831);
and U2402 (N_2402,N_1679,N_1821);
nor U2403 (N_2403,N_1930,N_1761);
or U2404 (N_2404,N_1949,N_1694);
and U2405 (N_2405,N_1608,N_1835);
and U2406 (N_2406,N_1602,N_1932);
xor U2407 (N_2407,N_1503,N_1719);
and U2408 (N_2408,N_1670,N_1991);
xor U2409 (N_2409,N_1796,N_1601);
xor U2410 (N_2410,N_1632,N_1527);
or U2411 (N_2411,N_1828,N_1845);
nor U2412 (N_2412,N_1986,N_1696);
or U2413 (N_2413,N_1521,N_1791);
nor U2414 (N_2414,N_1596,N_1716);
xnor U2415 (N_2415,N_1895,N_1829);
nand U2416 (N_2416,N_1571,N_1762);
and U2417 (N_2417,N_1926,N_1595);
and U2418 (N_2418,N_1695,N_1961);
nor U2419 (N_2419,N_1535,N_1539);
or U2420 (N_2420,N_1947,N_1917);
or U2421 (N_2421,N_1938,N_1885);
or U2422 (N_2422,N_1622,N_1737);
nand U2423 (N_2423,N_1684,N_1642);
and U2424 (N_2424,N_1505,N_1669);
or U2425 (N_2425,N_1862,N_1758);
and U2426 (N_2426,N_1763,N_1887);
xnor U2427 (N_2427,N_1747,N_1921);
xnor U2428 (N_2428,N_1713,N_1712);
or U2429 (N_2429,N_1556,N_1931);
nor U2430 (N_2430,N_1961,N_1715);
nand U2431 (N_2431,N_1870,N_1776);
nor U2432 (N_2432,N_1913,N_1849);
nor U2433 (N_2433,N_1921,N_1655);
or U2434 (N_2434,N_1614,N_1510);
xor U2435 (N_2435,N_1892,N_1793);
xnor U2436 (N_2436,N_1790,N_1862);
xnor U2437 (N_2437,N_1847,N_1986);
nand U2438 (N_2438,N_1844,N_1768);
and U2439 (N_2439,N_1612,N_1795);
or U2440 (N_2440,N_1702,N_1641);
nand U2441 (N_2441,N_1665,N_1596);
nor U2442 (N_2442,N_1736,N_1601);
or U2443 (N_2443,N_1555,N_1770);
and U2444 (N_2444,N_1785,N_1813);
or U2445 (N_2445,N_1502,N_1781);
nor U2446 (N_2446,N_1707,N_1909);
nor U2447 (N_2447,N_1822,N_1763);
and U2448 (N_2448,N_1662,N_1625);
or U2449 (N_2449,N_1810,N_1594);
xor U2450 (N_2450,N_1903,N_1515);
nor U2451 (N_2451,N_1573,N_1836);
nand U2452 (N_2452,N_1973,N_1854);
or U2453 (N_2453,N_1900,N_1600);
xor U2454 (N_2454,N_1863,N_1608);
xnor U2455 (N_2455,N_1950,N_1903);
and U2456 (N_2456,N_1809,N_1929);
xor U2457 (N_2457,N_1574,N_1895);
and U2458 (N_2458,N_1685,N_1819);
and U2459 (N_2459,N_1629,N_1788);
and U2460 (N_2460,N_1763,N_1945);
nand U2461 (N_2461,N_1705,N_1643);
nand U2462 (N_2462,N_1818,N_1659);
nor U2463 (N_2463,N_1819,N_1994);
nand U2464 (N_2464,N_1580,N_1574);
nand U2465 (N_2465,N_1854,N_1961);
and U2466 (N_2466,N_1750,N_1595);
and U2467 (N_2467,N_1775,N_1830);
and U2468 (N_2468,N_1959,N_1830);
and U2469 (N_2469,N_1573,N_1501);
nor U2470 (N_2470,N_1976,N_1701);
or U2471 (N_2471,N_1894,N_1970);
or U2472 (N_2472,N_1771,N_1913);
nand U2473 (N_2473,N_1867,N_1784);
nor U2474 (N_2474,N_1661,N_1630);
or U2475 (N_2475,N_1846,N_1635);
or U2476 (N_2476,N_1645,N_1504);
and U2477 (N_2477,N_1571,N_1946);
and U2478 (N_2478,N_1803,N_1727);
xnor U2479 (N_2479,N_1836,N_1765);
or U2480 (N_2480,N_1526,N_1868);
and U2481 (N_2481,N_1678,N_1681);
nor U2482 (N_2482,N_1986,N_1816);
and U2483 (N_2483,N_1512,N_1885);
and U2484 (N_2484,N_1559,N_1554);
or U2485 (N_2485,N_1794,N_1699);
or U2486 (N_2486,N_1583,N_1925);
and U2487 (N_2487,N_1784,N_1635);
nand U2488 (N_2488,N_1858,N_1981);
xnor U2489 (N_2489,N_1827,N_1813);
xor U2490 (N_2490,N_1890,N_1961);
and U2491 (N_2491,N_1503,N_1800);
and U2492 (N_2492,N_1920,N_1907);
xnor U2493 (N_2493,N_1907,N_1750);
nand U2494 (N_2494,N_1752,N_1510);
and U2495 (N_2495,N_1658,N_1930);
and U2496 (N_2496,N_1547,N_1712);
nand U2497 (N_2497,N_1880,N_1606);
or U2498 (N_2498,N_1640,N_1784);
and U2499 (N_2499,N_1896,N_1970);
or U2500 (N_2500,N_2372,N_2461);
xor U2501 (N_2501,N_2420,N_2245);
and U2502 (N_2502,N_2021,N_2264);
and U2503 (N_2503,N_2348,N_2206);
nor U2504 (N_2504,N_2107,N_2242);
xor U2505 (N_2505,N_2471,N_2033);
and U2506 (N_2506,N_2370,N_2199);
and U2507 (N_2507,N_2109,N_2266);
nand U2508 (N_2508,N_2086,N_2333);
xor U2509 (N_2509,N_2031,N_2295);
and U2510 (N_2510,N_2052,N_2490);
or U2511 (N_2511,N_2345,N_2185);
xnor U2512 (N_2512,N_2044,N_2045);
and U2513 (N_2513,N_2124,N_2169);
or U2514 (N_2514,N_2275,N_2284);
xor U2515 (N_2515,N_2120,N_2075);
xnor U2516 (N_2516,N_2176,N_2080);
xnor U2517 (N_2517,N_2493,N_2183);
xnor U2518 (N_2518,N_2391,N_2438);
nand U2519 (N_2519,N_2362,N_2177);
or U2520 (N_2520,N_2153,N_2323);
and U2521 (N_2521,N_2026,N_2322);
and U2522 (N_2522,N_2108,N_2152);
nor U2523 (N_2523,N_2316,N_2262);
nand U2524 (N_2524,N_2133,N_2016);
and U2525 (N_2525,N_2078,N_2378);
nor U2526 (N_2526,N_2306,N_2116);
and U2527 (N_2527,N_2427,N_2331);
xor U2528 (N_2528,N_2246,N_2201);
nor U2529 (N_2529,N_2138,N_2095);
nand U2530 (N_2530,N_2137,N_2130);
xnor U2531 (N_2531,N_2430,N_2288);
and U2532 (N_2532,N_2069,N_2175);
and U2533 (N_2533,N_2312,N_2478);
nand U2534 (N_2534,N_2117,N_2468);
nor U2535 (N_2535,N_2271,N_2261);
xor U2536 (N_2536,N_2101,N_2499);
or U2537 (N_2537,N_2233,N_2277);
and U2538 (N_2538,N_2325,N_2413);
or U2539 (N_2539,N_2278,N_2441);
nand U2540 (N_2540,N_2431,N_2005);
nor U2541 (N_2541,N_2327,N_2293);
nand U2542 (N_2542,N_2014,N_2215);
xor U2543 (N_2543,N_2047,N_2003);
and U2544 (N_2544,N_2172,N_2097);
nand U2545 (N_2545,N_2113,N_2477);
or U2546 (N_2546,N_2329,N_2416);
nor U2547 (N_2547,N_2415,N_2482);
nand U2548 (N_2548,N_2421,N_2213);
xor U2549 (N_2549,N_2168,N_2119);
and U2550 (N_2550,N_2292,N_2163);
nand U2551 (N_2551,N_2358,N_2207);
nor U2552 (N_2552,N_2324,N_2000);
xnor U2553 (N_2553,N_2311,N_2291);
nand U2554 (N_2554,N_2072,N_2286);
nor U2555 (N_2555,N_2382,N_2128);
and U2556 (N_2556,N_2229,N_2435);
and U2557 (N_2557,N_2191,N_2161);
xnor U2558 (N_2558,N_2463,N_2030);
nor U2559 (N_2559,N_2457,N_2068);
nor U2560 (N_2560,N_2301,N_2158);
and U2561 (N_2561,N_2450,N_2092);
nand U2562 (N_2562,N_2151,N_2453);
xnor U2563 (N_2563,N_2002,N_2056);
or U2564 (N_2564,N_2162,N_2355);
and U2565 (N_2565,N_2099,N_2218);
and U2566 (N_2566,N_2258,N_2313);
nor U2567 (N_2567,N_2340,N_2223);
nor U2568 (N_2568,N_2148,N_2051);
nor U2569 (N_2569,N_2352,N_2073);
or U2570 (N_2570,N_2318,N_2144);
xor U2571 (N_2571,N_2321,N_2209);
and U2572 (N_2572,N_2405,N_2257);
and U2573 (N_2573,N_2272,N_2127);
nor U2574 (N_2574,N_2254,N_2200);
and U2575 (N_2575,N_2319,N_2028);
xor U2576 (N_2576,N_2436,N_2303);
nand U2577 (N_2577,N_2354,N_2090);
nor U2578 (N_2578,N_2198,N_2432);
nor U2579 (N_2579,N_2429,N_2235);
nand U2580 (N_2580,N_2225,N_2081);
xor U2581 (N_2581,N_2433,N_2469);
nand U2582 (N_2582,N_2126,N_2193);
nor U2583 (N_2583,N_2243,N_2195);
nor U2584 (N_2584,N_2279,N_2424);
xnor U2585 (N_2585,N_2335,N_2473);
xnor U2586 (N_2586,N_2058,N_2377);
or U2587 (N_2587,N_2399,N_2167);
nor U2588 (N_2588,N_2308,N_2488);
xor U2589 (N_2589,N_2492,N_2139);
xor U2590 (N_2590,N_2070,N_2496);
and U2591 (N_2591,N_2360,N_2236);
nor U2592 (N_2592,N_2143,N_2350);
and U2593 (N_2593,N_2451,N_2012);
and U2594 (N_2594,N_2364,N_2210);
nand U2595 (N_2595,N_2001,N_2211);
nor U2596 (N_2596,N_2131,N_2023);
or U2597 (N_2597,N_2087,N_2226);
nor U2598 (N_2598,N_2224,N_2460);
nand U2599 (N_2599,N_2334,N_2443);
and U2600 (N_2600,N_2349,N_2196);
nor U2601 (N_2601,N_2479,N_2216);
nor U2602 (N_2602,N_2102,N_2204);
nor U2603 (N_2603,N_2297,N_2357);
or U2604 (N_2604,N_2423,N_2125);
nor U2605 (N_2605,N_2181,N_2486);
nor U2606 (N_2606,N_2466,N_2300);
xor U2607 (N_2607,N_2020,N_2426);
and U2608 (N_2608,N_2437,N_2076);
xnor U2609 (N_2609,N_2418,N_2228);
or U2610 (N_2610,N_2009,N_2449);
nor U2611 (N_2611,N_2179,N_2055);
xor U2612 (N_2612,N_2406,N_2011);
xnor U2613 (N_2613,N_2088,N_2013);
and U2614 (N_2614,N_2356,N_2403);
or U2615 (N_2615,N_2280,N_2192);
and U2616 (N_2616,N_2239,N_2342);
or U2617 (N_2617,N_2396,N_2018);
xnor U2618 (N_2618,N_2134,N_2386);
and U2619 (N_2619,N_2481,N_2458);
nor U2620 (N_2620,N_2497,N_2149);
nor U2621 (N_2621,N_2274,N_2412);
or U2622 (N_2622,N_2019,N_2351);
xnor U2623 (N_2623,N_2314,N_2285);
and U2624 (N_2624,N_2462,N_2170);
nand U2625 (N_2625,N_2470,N_2244);
nor U2626 (N_2626,N_2269,N_2414);
nor U2627 (N_2627,N_2428,N_2485);
nor U2628 (N_2628,N_2184,N_2039);
nand U2629 (N_2629,N_2214,N_2283);
xnor U2630 (N_2630,N_2157,N_2483);
or U2631 (N_2631,N_2132,N_2159);
or U2632 (N_2632,N_2096,N_2017);
nand U2633 (N_2633,N_2231,N_2273);
and U2634 (N_2634,N_2048,N_2221);
or U2635 (N_2635,N_2141,N_2155);
and U2636 (N_2636,N_2029,N_2118);
xnor U2637 (N_2637,N_2008,N_2383);
nor U2638 (N_2638,N_2142,N_2281);
nor U2639 (N_2639,N_2140,N_2232);
nor U2640 (N_2640,N_2103,N_2010);
nand U2641 (N_2641,N_2104,N_2135);
xor U2642 (N_2642,N_2267,N_2150);
nor U2643 (N_2643,N_2190,N_2004);
nor U2644 (N_2644,N_2160,N_2037);
and U2645 (N_2645,N_2397,N_2307);
nor U2646 (N_2646,N_2392,N_2344);
nand U2647 (N_2647,N_2455,N_2385);
nand U2648 (N_2648,N_2419,N_2240);
or U2649 (N_2649,N_2250,N_2178);
and U2650 (N_2650,N_2353,N_2027);
and U2651 (N_2651,N_2465,N_2110);
or U2652 (N_2652,N_2077,N_2064);
and U2653 (N_2653,N_2373,N_2467);
nor U2654 (N_2654,N_2060,N_2186);
nor U2655 (N_2655,N_2388,N_2253);
nand U2656 (N_2656,N_2252,N_2336);
xor U2657 (N_2657,N_2038,N_2374);
xnor U2658 (N_2658,N_2263,N_2040);
nand U2659 (N_2659,N_2442,N_2122);
or U2660 (N_2660,N_2480,N_2270);
or U2661 (N_2661,N_2251,N_2194);
nor U2662 (N_2662,N_2346,N_2491);
and U2663 (N_2663,N_2205,N_2282);
nor U2664 (N_2664,N_2091,N_2294);
nand U2665 (N_2665,N_2400,N_2067);
nor U2666 (N_2666,N_2456,N_2376);
and U2667 (N_2667,N_2022,N_2255);
and U2668 (N_2668,N_2381,N_2094);
and U2669 (N_2669,N_2290,N_2114);
nand U2670 (N_2670,N_2384,N_2380);
xnor U2671 (N_2671,N_2434,N_2136);
xnor U2672 (N_2672,N_2222,N_2289);
nand U2673 (N_2673,N_2057,N_2036);
xor U2674 (N_2674,N_2174,N_2459);
and U2675 (N_2675,N_2230,N_2024);
xor U2676 (N_2676,N_2444,N_2189);
nor U2677 (N_2677,N_2394,N_2310);
or U2678 (N_2678,N_2276,N_2407);
nand U2679 (N_2679,N_2476,N_2123);
or U2680 (N_2680,N_2452,N_2182);
xnor U2681 (N_2681,N_2085,N_2464);
nor U2682 (N_2682,N_2079,N_2105);
xor U2683 (N_2683,N_2154,N_2265);
and U2684 (N_2684,N_2445,N_2164);
or U2685 (N_2685,N_2417,N_2409);
xor U2686 (N_2686,N_2309,N_2089);
nand U2687 (N_2687,N_2146,N_2212);
nand U2688 (N_2688,N_2059,N_2389);
nor U2689 (N_2689,N_2098,N_2343);
or U2690 (N_2690,N_2165,N_2330);
nand U2691 (N_2691,N_2145,N_2446);
nand U2692 (N_2692,N_2234,N_2366);
xor U2693 (N_2693,N_2337,N_2112);
and U2694 (N_2694,N_2249,N_2341);
nand U2695 (N_2695,N_2043,N_2188);
or U2696 (N_2696,N_2365,N_2083);
or U2697 (N_2697,N_2296,N_2111);
nand U2698 (N_2698,N_2422,N_2025);
nor U2699 (N_2699,N_2129,N_2203);
nand U2700 (N_2700,N_2487,N_2454);
nor U2701 (N_2701,N_2338,N_2408);
nor U2702 (N_2702,N_2049,N_2006);
nand U2703 (N_2703,N_2371,N_2484);
xor U2704 (N_2704,N_2260,N_2171);
and U2705 (N_2705,N_2015,N_2495);
and U2706 (N_2706,N_2187,N_2066);
or U2707 (N_2707,N_2147,N_2106);
and U2708 (N_2708,N_2390,N_2363);
and U2709 (N_2709,N_2404,N_2268);
nor U2710 (N_2710,N_2401,N_2398);
and U2711 (N_2711,N_2448,N_2007);
or U2712 (N_2712,N_2042,N_2379);
nor U2713 (N_2713,N_2305,N_2359);
and U2714 (N_2714,N_2082,N_2220);
xor U2715 (N_2715,N_2202,N_2100);
and U2716 (N_2716,N_2304,N_2166);
nor U2717 (N_2717,N_2411,N_2440);
nand U2718 (N_2718,N_2368,N_2156);
and U2719 (N_2719,N_2410,N_2115);
or U2720 (N_2720,N_2326,N_2035);
nand U2721 (N_2721,N_2375,N_2474);
nand U2722 (N_2722,N_2393,N_2093);
and U2723 (N_2723,N_2367,N_2065);
xnor U2724 (N_2724,N_2062,N_2425);
nand U2725 (N_2725,N_2071,N_2032);
nand U2726 (N_2726,N_2317,N_2315);
and U2727 (N_2727,N_2387,N_2219);
or U2728 (N_2728,N_2238,N_2063);
and U2729 (N_2729,N_2061,N_2046);
or U2730 (N_2730,N_2320,N_2241);
and U2731 (N_2731,N_2054,N_2298);
or U2732 (N_2732,N_2361,N_2053);
and U2733 (N_2733,N_2041,N_2339);
nand U2734 (N_2734,N_2489,N_2227);
or U2735 (N_2735,N_2237,N_2299);
xnor U2736 (N_2736,N_2498,N_2074);
and U2737 (N_2737,N_2328,N_2197);
nand U2738 (N_2738,N_2439,N_2084);
or U2739 (N_2739,N_2256,N_2287);
and U2740 (N_2740,N_2472,N_2302);
nand U2741 (N_2741,N_2180,N_2347);
nor U2742 (N_2742,N_2034,N_2208);
nand U2743 (N_2743,N_2173,N_2494);
or U2744 (N_2744,N_2395,N_2050);
and U2745 (N_2745,N_2475,N_2247);
nand U2746 (N_2746,N_2332,N_2217);
nand U2747 (N_2747,N_2259,N_2121);
and U2748 (N_2748,N_2248,N_2369);
or U2749 (N_2749,N_2402,N_2447);
nand U2750 (N_2750,N_2040,N_2299);
nor U2751 (N_2751,N_2447,N_2310);
nor U2752 (N_2752,N_2337,N_2357);
and U2753 (N_2753,N_2086,N_2496);
and U2754 (N_2754,N_2211,N_2491);
nand U2755 (N_2755,N_2115,N_2021);
xnor U2756 (N_2756,N_2232,N_2142);
nor U2757 (N_2757,N_2195,N_2005);
nand U2758 (N_2758,N_2054,N_2173);
xor U2759 (N_2759,N_2233,N_2073);
and U2760 (N_2760,N_2296,N_2386);
xnor U2761 (N_2761,N_2487,N_2460);
and U2762 (N_2762,N_2468,N_2105);
nand U2763 (N_2763,N_2265,N_2255);
or U2764 (N_2764,N_2032,N_2054);
or U2765 (N_2765,N_2186,N_2472);
or U2766 (N_2766,N_2431,N_2448);
or U2767 (N_2767,N_2461,N_2137);
and U2768 (N_2768,N_2165,N_2278);
nor U2769 (N_2769,N_2222,N_2450);
and U2770 (N_2770,N_2484,N_2330);
and U2771 (N_2771,N_2071,N_2247);
nor U2772 (N_2772,N_2214,N_2139);
nand U2773 (N_2773,N_2068,N_2427);
nor U2774 (N_2774,N_2405,N_2086);
nand U2775 (N_2775,N_2486,N_2498);
and U2776 (N_2776,N_2138,N_2088);
or U2777 (N_2777,N_2007,N_2496);
nand U2778 (N_2778,N_2396,N_2317);
or U2779 (N_2779,N_2279,N_2398);
and U2780 (N_2780,N_2481,N_2317);
xnor U2781 (N_2781,N_2203,N_2366);
or U2782 (N_2782,N_2202,N_2052);
nand U2783 (N_2783,N_2298,N_2378);
nor U2784 (N_2784,N_2269,N_2381);
nand U2785 (N_2785,N_2141,N_2255);
and U2786 (N_2786,N_2024,N_2435);
nor U2787 (N_2787,N_2238,N_2103);
nor U2788 (N_2788,N_2315,N_2221);
xnor U2789 (N_2789,N_2462,N_2306);
or U2790 (N_2790,N_2338,N_2288);
and U2791 (N_2791,N_2173,N_2085);
and U2792 (N_2792,N_2180,N_2364);
or U2793 (N_2793,N_2206,N_2288);
or U2794 (N_2794,N_2304,N_2386);
xnor U2795 (N_2795,N_2101,N_2313);
xnor U2796 (N_2796,N_2178,N_2034);
nor U2797 (N_2797,N_2138,N_2411);
nand U2798 (N_2798,N_2035,N_2250);
and U2799 (N_2799,N_2016,N_2006);
and U2800 (N_2800,N_2175,N_2227);
xor U2801 (N_2801,N_2468,N_2092);
or U2802 (N_2802,N_2086,N_2353);
xnor U2803 (N_2803,N_2152,N_2160);
nand U2804 (N_2804,N_2004,N_2481);
nand U2805 (N_2805,N_2028,N_2181);
or U2806 (N_2806,N_2267,N_2087);
or U2807 (N_2807,N_2232,N_2459);
xnor U2808 (N_2808,N_2009,N_2003);
nand U2809 (N_2809,N_2120,N_2265);
or U2810 (N_2810,N_2141,N_2393);
and U2811 (N_2811,N_2149,N_2380);
xnor U2812 (N_2812,N_2373,N_2265);
nor U2813 (N_2813,N_2368,N_2417);
nor U2814 (N_2814,N_2424,N_2126);
xor U2815 (N_2815,N_2386,N_2178);
nand U2816 (N_2816,N_2419,N_2256);
xor U2817 (N_2817,N_2417,N_2365);
and U2818 (N_2818,N_2069,N_2237);
xnor U2819 (N_2819,N_2444,N_2306);
nand U2820 (N_2820,N_2369,N_2433);
nand U2821 (N_2821,N_2154,N_2212);
xnor U2822 (N_2822,N_2323,N_2055);
nand U2823 (N_2823,N_2407,N_2469);
nor U2824 (N_2824,N_2130,N_2334);
and U2825 (N_2825,N_2426,N_2383);
nand U2826 (N_2826,N_2253,N_2050);
xor U2827 (N_2827,N_2217,N_2471);
and U2828 (N_2828,N_2235,N_2440);
xnor U2829 (N_2829,N_2051,N_2267);
and U2830 (N_2830,N_2057,N_2281);
xnor U2831 (N_2831,N_2428,N_2275);
nand U2832 (N_2832,N_2250,N_2075);
xnor U2833 (N_2833,N_2066,N_2275);
xnor U2834 (N_2834,N_2087,N_2387);
nor U2835 (N_2835,N_2242,N_2272);
and U2836 (N_2836,N_2024,N_2347);
or U2837 (N_2837,N_2369,N_2452);
nor U2838 (N_2838,N_2249,N_2074);
nand U2839 (N_2839,N_2048,N_2479);
and U2840 (N_2840,N_2386,N_2030);
xnor U2841 (N_2841,N_2348,N_2372);
nor U2842 (N_2842,N_2282,N_2376);
nand U2843 (N_2843,N_2208,N_2114);
nor U2844 (N_2844,N_2326,N_2227);
xor U2845 (N_2845,N_2207,N_2115);
or U2846 (N_2846,N_2006,N_2355);
nand U2847 (N_2847,N_2496,N_2322);
or U2848 (N_2848,N_2160,N_2052);
xor U2849 (N_2849,N_2296,N_2283);
or U2850 (N_2850,N_2232,N_2393);
or U2851 (N_2851,N_2001,N_2108);
xor U2852 (N_2852,N_2161,N_2347);
nand U2853 (N_2853,N_2019,N_2200);
xnor U2854 (N_2854,N_2475,N_2201);
nand U2855 (N_2855,N_2327,N_2029);
and U2856 (N_2856,N_2430,N_2170);
xor U2857 (N_2857,N_2439,N_2278);
or U2858 (N_2858,N_2015,N_2423);
or U2859 (N_2859,N_2196,N_2416);
or U2860 (N_2860,N_2328,N_2324);
nor U2861 (N_2861,N_2338,N_2426);
xnor U2862 (N_2862,N_2402,N_2345);
or U2863 (N_2863,N_2356,N_2387);
or U2864 (N_2864,N_2495,N_2164);
or U2865 (N_2865,N_2300,N_2141);
or U2866 (N_2866,N_2170,N_2164);
xnor U2867 (N_2867,N_2136,N_2235);
xor U2868 (N_2868,N_2332,N_2128);
xor U2869 (N_2869,N_2271,N_2442);
and U2870 (N_2870,N_2308,N_2360);
xor U2871 (N_2871,N_2211,N_2230);
nor U2872 (N_2872,N_2052,N_2466);
and U2873 (N_2873,N_2036,N_2285);
or U2874 (N_2874,N_2010,N_2071);
or U2875 (N_2875,N_2274,N_2218);
and U2876 (N_2876,N_2473,N_2316);
nand U2877 (N_2877,N_2377,N_2485);
and U2878 (N_2878,N_2286,N_2458);
and U2879 (N_2879,N_2167,N_2164);
or U2880 (N_2880,N_2226,N_2057);
xnor U2881 (N_2881,N_2070,N_2218);
and U2882 (N_2882,N_2333,N_2309);
nand U2883 (N_2883,N_2376,N_2324);
nand U2884 (N_2884,N_2216,N_2401);
and U2885 (N_2885,N_2036,N_2463);
or U2886 (N_2886,N_2209,N_2039);
and U2887 (N_2887,N_2438,N_2167);
nand U2888 (N_2888,N_2004,N_2137);
nand U2889 (N_2889,N_2205,N_2174);
nor U2890 (N_2890,N_2207,N_2478);
and U2891 (N_2891,N_2323,N_2016);
nor U2892 (N_2892,N_2349,N_2122);
nand U2893 (N_2893,N_2337,N_2283);
xor U2894 (N_2894,N_2029,N_2143);
and U2895 (N_2895,N_2300,N_2399);
or U2896 (N_2896,N_2015,N_2209);
nand U2897 (N_2897,N_2028,N_2131);
xor U2898 (N_2898,N_2377,N_2436);
or U2899 (N_2899,N_2211,N_2452);
xor U2900 (N_2900,N_2424,N_2007);
nand U2901 (N_2901,N_2248,N_2276);
nor U2902 (N_2902,N_2182,N_2318);
or U2903 (N_2903,N_2283,N_2461);
or U2904 (N_2904,N_2269,N_2484);
or U2905 (N_2905,N_2140,N_2094);
or U2906 (N_2906,N_2090,N_2193);
and U2907 (N_2907,N_2289,N_2322);
or U2908 (N_2908,N_2005,N_2120);
or U2909 (N_2909,N_2263,N_2441);
nor U2910 (N_2910,N_2492,N_2373);
or U2911 (N_2911,N_2411,N_2005);
and U2912 (N_2912,N_2198,N_2250);
nand U2913 (N_2913,N_2177,N_2436);
or U2914 (N_2914,N_2043,N_2232);
or U2915 (N_2915,N_2344,N_2494);
nand U2916 (N_2916,N_2165,N_2482);
nand U2917 (N_2917,N_2195,N_2370);
or U2918 (N_2918,N_2337,N_2032);
xnor U2919 (N_2919,N_2115,N_2436);
xnor U2920 (N_2920,N_2139,N_2195);
nor U2921 (N_2921,N_2055,N_2409);
or U2922 (N_2922,N_2007,N_2368);
and U2923 (N_2923,N_2261,N_2301);
nor U2924 (N_2924,N_2269,N_2036);
or U2925 (N_2925,N_2350,N_2408);
xor U2926 (N_2926,N_2194,N_2127);
or U2927 (N_2927,N_2353,N_2154);
nor U2928 (N_2928,N_2189,N_2051);
or U2929 (N_2929,N_2255,N_2381);
or U2930 (N_2930,N_2394,N_2253);
or U2931 (N_2931,N_2293,N_2156);
nand U2932 (N_2932,N_2465,N_2442);
and U2933 (N_2933,N_2084,N_2283);
or U2934 (N_2934,N_2266,N_2352);
nor U2935 (N_2935,N_2194,N_2021);
xnor U2936 (N_2936,N_2215,N_2151);
nor U2937 (N_2937,N_2222,N_2362);
or U2938 (N_2938,N_2232,N_2084);
xnor U2939 (N_2939,N_2465,N_2137);
nor U2940 (N_2940,N_2023,N_2240);
nor U2941 (N_2941,N_2441,N_2039);
nor U2942 (N_2942,N_2120,N_2113);
and U2943 (N_2943,N_2015,N_2151);
nand U2944 (N_2944,N_2261,N_2485);
xnor U2945 (N_2945,N_2472,N_2486);
nand U2946 (N_2946,N_2459,N_2344);
nand U2947 (N_2947,N_2338,N_2343);
nor U2948 (N_2948,N_2419,N_2145);
or U2949 (N_2949,N_2281,N_2052);
xor U2950 (N_2950,N_2293,N_2175);
and U2951 (N_2951,N_2377,N_2387);
or U2952 (N_2952,N_2063,N_2464);
xor U2953 (N_2953,N_2318,N_2067);
nor U2954 (N_2954,N_2085,N_2001);
or U2955 (N_2955,N_2251,N_2429);
nor U2956 (N_2956,N_2172,N_2459);
and U2957 (N_2957,N_2203,N_2003);
nand U2958 (N_2958,N_2164,N_2466);
nand U2959 (N_2959,N_2314,N_2187);
or U2960 (N_2960,N_2142,N_2277);
xnor U2961 (N_2961,N_2471,N_2346);
nor U2962 (N_2962,N_2440,N_2343);
or U2963 (N_2963,N_2084,N_2188);
or U2964 (N_2964,N_2436,N_2428);
nand U2965 (N_2965,N_2096,N_2117);
nor U2966 (N_2966,N_2164,N_2387);
nand U2967 (N_2967,N_2188,N_2000);
nand U2968 (N_2968,N_2010,N_2171);
and U2969 (N_2969,N_2361,N_2304);
and U2970 (N_2970,N_2393,N_2358);
and U2971 (N_2971,N_2482,N_2166);
and U2972 (N_2972,N_2063,N_2399);
xor U2973 (N_2973,N_2498,N_2053);
nand U2974 (N_2974,N_2263,N_2457);
nor U2975 (N_2975,N_2148,N_2276);
xor U2976 (N_2976,N_2049,N_2203);
nand U2977 (N_2977,N_2093,N_2049);
and U2978 (N_2978,N_2290,N_2104);
nor U2979 (N_2979,N_2055,N_2205);
and U2980 (N_2980,N_2074,N_2400);
nor U2981 (N_2981,N_2279,N_2087);
nor U2982 (N_2982,N_2329,N_2130);
nand U2983 (N_2983,N_2163,N_2487);
and U2984 (N_2984,N_2151,N_2314);
nor U2985 (N_2985,N_2212,N_2148);
xor U2986 (N_2986,N_2259,N_2034);
nor U2987 (N_2987,N_2134,N_2276);
nor U2988 (N_2988,N_2468,N_2027);
and U2989 (N_2989,N_2030,N_2032);
xor U2990 (N_2990,N_2335,N_2082);
nand U2991 (N_2991,N_2027,N_2215);
and U2992 (N_2992,N_2049,N_2370);
and U2993 (N_2993,N_2019,N_2281);
xnor U2994 (N_2994,N_2364,N_2041);
or U2995 (N_2995,N_2117,N_2153);
xor U2996 (N_2996,N_2030,N_2105);
and U2997 (N_2997,N_2054,N_2095);
nand U2998 (N_2998,N_2105,N_2342);
nor U2999 (N_2999,N_2238,N_2279);
or U3000 (N_3000,N_2885,N_2594);
nor U3001 (N_3001,N_2558,N_2519);
or U3002 (N_3002,N_2824,N_2653);
or U3003 (N_3003,N_2698,N_2748);
nand U3004 (N_3004,N_2809,N_2630);
nor U3005 (N_3005,N_2680,N_2669);
or U3006 (N_3006,N_2566,N_2807);
nand U3007 (N_3007,N_2977,N_2887);
xnor U3008 (N_3008,N_2504,N_2736);
xor U3009 (N_3009,N_2837,N_2666);
xnor U3010 (N_3010,N_2581,N_2952);
or U3011 (N_3011,N_2593,N_2801);
and U3012 (N_3012,N_2909,N_2918);
nand U3013 (N_3013,N_2552,N_2522);
or U3014 (N_3014,N_2700,N_2777);
nand U3015 (N_3015,N_2521,N_2897);
xnor U3016 (N_3016,N_2720,N_2617);
nor U3017 (N_3017,N_2658,N_2815);
and U3018 (N_3018,N_2969,N_2834);
xnor U3019 (N_3019,N_2981,N_2990);
nor U3020 (N_3020,N_2673,N_2683);
nand U3021 (N_3021,N_2975,N_2710);
and U3022 (N_3022,N_2764,N_2670);
and U3023 (N_3023,N_2546,N_2964);
xnor U3024 (N_3024,N_2625,N_2967);
nor U3025 (N_3025,N_2852,N_2532);
and U3026 (N_3026,N_2999,N_2941);
nor U3027 (N_3027,N_2585,N_2946);
or U3028 (N_3028,N_2828,N_2765);
and U3029 (N_3029,N_2757,N_2712);
or U3030 (N_3030,N_2649,N_2867);
xnor U3031 (N_3031,N_2770,N_2760);
or U3032 (N_3032,N_2877,N_2746);
xnor U3033 (N_3033,N_2668,N_2699);
nor U3034 (N_3034,N_2703,N_2800);
and U3035 (N_3035,N_2995,N_2983);
nand U3036 (N_3036,N_2903,N_2963);
and U3037 (N_3037,N_2869,N_2934);
nand U3038 (N_3038,N_2604,N_2557);
or U3039 (N_3039,N_2634,N_2819);
xor U3040 (N_3040,N_2864,N_2664);
nand U3041 (N_3041,N_2541,N_2719);
xnor U3042 (N_3042,N_2539,N_2763);
and U3043 (N_3043,N_2635,N_2970);
and U3044 (N_3044,N_2985,N_2926);
and U3045 (N_3045,N_2832,N_2870);
xor U3046 (N_3046,N_2682,N_2709);
and U3047 (N_3047,N_2711,N_2958);
and U3048 (N_3048,N_2810,N_2553);
or U3049 (N_3049,N_2671,N_2904);
xnor U3050 (N_3050,N_2672,N_2761);
nand U3051 (N_3051,N_2913,N_2562);
nand U3052 (N_3052,N_2804,N_2560);
and U3053 (N_3053,N_2991,N_2880);
nand U3054 (N_3054,N_2621,N_2575);
nand U3055 (N_3055,N_2687,N_2846);
xor U3056 (N_3056,N_2895,N_2715);
and U3057 (N_3057,N_2652,N_2902);
nand U3058 (N_3058,N_2919,N_2729);
xnor U3059 (N_3059,N_2974,N_2749);
and U3060 (N_3060,N_2704,N_2578);
xor U3061 (N_3061,N_2582,N_2728);
nand U3062 (N_3062,N_2818,N_2708);
nand U3063 (N_3063,N_2656,N_2597);
and U3064 (N_3064,N_2953,N_2972);
or U3065 (N_3065,N_2697,N_2949);
xor U3066 (N_3066,N_2599,N_2986);
nor U3067 (N_3067,N_2962,N_2610);
and U3068 (N_3068,N_2858,N_2805);
nor U3069 (N_3069,N_2659,N_2802);
and U3070 (N_3070,N_2611,N_2798);
nand U3071 (N_3071,N_2542,N_2910);
nor U3072 (N_3072,N_2775,N_2608);
nand U3073 (N_3073,N_2745,N_2791);
and U3074 (N_3074,N_2780,N_2540);
or U3075 (N_3075,N_2734,N_2561);
or U3076 (N_3076,N_2943,N_2527);
nor U3077 (N_3077,N_2839,N_2718);
and U3078 (N_3078,N_2754,N_2901);
and U3079 (N_3079,N_2702,N_2848);
nand U3080 (N_3080,N_2771,N_2788);
nor U3081 (N_3081,N_2923,N_2998);
and U3082 (N_3082,N_2767,N_2722);
and U3083 (N_3083,N_2743,N_2549);
nand U3084 (N_3084,N_2694,N_2940);
or U3085 (N_3085,N_2841,N_2888);
or U3086 (N_3086,N_2654,N_2730);
and U3087 (N_3087,N_2871,N_2528);
xnor U3088 (N_3088,N_2808,N_2626);
nand U3089 (N_3089,N_2568,N_2931);
nand U3090 (N_3090,N_2739,N_2620);
and U3091 (N_3091,N_2782,N_2598);
xnor U3092 (N_3092,N_2847,N_2559);
nand U3093 (N_3093,N_2778,N_2922);
nor U3094 (N_3094,N_2851,N_2531);
nor U3095 (N_3095,N_2500,N_2735);
xor U3096 (N_3096,N_2883,N_2510);
xnor U3097 (N_3097,N_2744,N_2723);
xnor U3098 (N_3098,N_2667,N_2533);
or U3099 (N_3099,N_2688,N_2966);
and U3100 (N_3100,N_2979,N_2647);
nand U3101 (N_3101,N_2911,N_2956);
nor U3102 (N_3102,N_2890,N_2507);
or U3103 (N_3103,N_2517,N_2907);
nand U3104 (N_3104,N_2523,N_2811);
nor U3105 (N_3105,N_2564,N_2892);
nand U3106 (N_3106,N_2629,N_2938);
nor U3107 (N_3107,N_2752,N_2957);
or U3108 (N_3108,N_2679,N_2836);
nand U3109 (N_3109,N_2825,N_2845);
xor U3110 (N_3110,N_2886,N_2506);
xnor U3111 (N_3111,N_2982,N_2627);
xor U3112 (N_3112,N_2515,N_2917);
or U3113 (N_3113,N_2939,N_2584);
xor U3114 (N_3114,N_2950,N_2590);
or U3115 (N_3115,N_2795,N_2842);
or U3116 (N_3116,N_2865,N_2638);
and U3117 (N_3117,N_2936,N_2595);
and U3118 (N_3118,N_2548,N_2873);
and U3119 (N_3119,N_2550,N_2889);
and U3120 (N_3120,N_2721,N_2793);
and U3121 (N_3121,N_2534,N_2660);
nor U3122 (N_3122,N_2994,N_2577);
nand U3123 (N_3123,N_2965,N_2615);
nand U3124 (N_3124,N_2830,N_2993);
xor U3125 (N_3125,N_2861,N_2750);
nand U3126 (N_3126,N_2662,N_2769);
or U3127 (N_3127,N_2961,N_2536);
and U3128 (N_3128,N_2916,N_2947);
nand U3129 (N_3129,N_2573,N_2789);
and U3130 (N_3130,N_2505,N_2544);
xnor U3131 (N_3131,N_2929,N_2872);
and U3132 (N_3132,N_2650,N_2612);
nor U3133 (N_3133,N_2820,N_2605);
or U3134 (N_3134,N_2762,N_2792);
xnor U3135 (N_3135,N_2572,N_2645);
xor U3136 (N_3136,N_2874,N_2933);
nor U3137 (N_3137,N_2632,N_2678);
nor U3138 (N_3138,N_2740,N_2924);
nor U3139 (N_3139,N_2856,N_2690);
xor U3140 (N_3140,N_2755,N_2737);
and U3141 (N_3141,N_2591,N_2863);
xor U3142 (N_3142,N_2868,N_2583);
and U3143 (N_3143,N_2587,N_2600);
nand U3144 (N_3144,N_2618,N_2677);
xnor U3145 (N_3145,N_2607,N_2633);
and U3146 (N_3146,N_2648,N_2651);
and U3147 (N_3147,N_2827,N_2944);
nand U3148 (N_3148,N_2951,N_2565);
nor U3149 (N_3149,N_2996,N_2925);
or U3150 (N_3150,N_2772,N_2930);
xor U3151 (N_3151,N_2609,N_2823);
xnor U3152 (N_3152,N_2657,N_2602);
and U3153 (N_3153,N_2624,N_2636);
and U3154 (N_3154,N_2644,N_2731);
and U3155 (N_3155,N_2813,N_2696);
xor U3156 (N_3156,N_2787,N_2822);
or U3157 (N_3157,N_2525,N_2714);
nand U3158 (N_3158,N_2580,N_2753);
nand U3159 (N_3159,N_2705,N_2840);
and U3160 (N_3160,N_2516,N_2973);
nand U3161 (N_3161,N_2551,N_2716);
nand U3162 (N_3162,N_2642,N_2779);
xnor U3163 (N_3163,N_2826,N_2945);
nand U3164 (N_3164,N_2676,N_2843);
and U3165 (N_3165,N_2784,N_2799);
or U3166 (N_3166,N_2646,N_2742);
xnor U3167 (N_3167,N_2526,N_2751);
nor U3168 (N_3168,N_2535,N_2686);
nand U3169 (N_3169,N_2543,N_2968);
nor U3170 (N_3170,N_2576,N_2882);
or U3171 (N_3171,N_2537,N_2786);
nand U3172 (N_3172,N_2693,N_2850);
nor U3173 (N_3173,N_2921,N_2518);
xor U3174 (N_3174,N_2619,N_2655);
or U3175 (N_3175,N_2681,N_2741);
or U3176 (N_3176,N_2579,N_2601);
xnor U3177 (N_3177,N_2631,N_2643);
nor U3178 (N_3178,N_2684,N_2821);
nor U3179 (N_3179,N_2831,N_2733);
nor U3180 (N_3180,N_2773,N_2640);
or U3181 (N_3181,N_2976,N_2586);
xor U3182 (N_3182,N_2955,N_2768);
xnor U3183 (N_3183,N_2503,N_2978);
xnor U3184 (N_3184,N_2524,N_2724);
xnor U3185 (N_3185,N_2992,N_2674);
and U3186 (N_3186,N_2554,N_2606);
nand U3187 (N_3187,N_2876,N_2814);
and U3188 (N_3188,N_2896,N_2920);
nand U3189 (N_3189,N_2639,N_2988);
or U3190 (N_3190,N_2853,N_2812);
nor U3191 (N_3191,N_2783,N_2623);
xnor U3192 (N_3192,N_2908,N_2854);
xnor U3193 (N_3193,N_2756,N_2835);
nand U3194 (N_3194,N_2563,N_2637);
xnor U3195 (N_3195,N_2891,N_2695);
nor U3196 (N_3196,N_2614,N_2727);
or U3197 (N_3197,N_2790,N_2717);
nand U3198 (N_3198,N_2914,N_2588);
xnor U3199 (N_3199,N_2833,N_2747);
nand U3200 (N_3200,N_2529,N_2935);
or U3201 (N_3201,N_2857,N_2571);
xor U3202 (N_3202,N_2937,N_2927);
nand U3203 (N_3203,N_2774,N_2838);
nand U3204 (N_3204,N_2794,N_2898);
nor U3205 (N_3205,N_2884,N_2530);
and U3206 (N_3206,N_2641,N_2675);
and U3207 (N_3207,N_2661,N_2596);
nand U3208 (N_3208,N_2855,N_2685);
nand U3209 (N_3209,N_2567,N_2691);
and U3210 (N_3210,N_2603,N_2862);
or U3211 (N_3211,N_2980,N_2797);
xor U3212 (N_3212,N_2859,N_2502);
xnor U3213 (N_3213,N_2948,N_2829);
or U3214 (N_3214,N_2899,N_2893);
and U3215 (N_3215,N_2906,N_2665);
and U3216 (N_3216,N_2732,N_2912);
nor U3217 (N_3217,N_2781,N_2692);
and U3218 (N_3218,N_2860,N_2987);
and U3219 (N_3219,N_2513,N_2569);
and U3220 (N_3220,N_2905,N_2806);
or U3221 (N_3221,N_2707,N_2713);
xnor U3222 (N_3222,N_2538,N_2766);
and U3223 (N_3223,N_2706,N_2881);
or U3224 (N_3224,N_2997,N_2570);
and U3225 (N_3225,N_2628,N_2776);
nor U3226 (N_3226,N_2915,N_2622);
xnor U3227 (N_3227,N_2875,N_2785);
or U3228 (N_3228,N_2545,N_2520);
nand U3229 (N_3229,N_2817,N_2942);
xnor U3230 (N_3230,N_2514,N_2689);
nand U3231 (N_3231,N_2900,N_2879);
nand U3232 (N_3232,N_2984,N_2508);
xor U3233 (N_3233,N_2556,N_2928);
nor U3234 (N_3234,N_2894,N_2512);
and U3235 (N_3235,N_2701,N_2866);
or U3236 (N_3236,N_2589,N_2960);
xor U3237 (N_3237,N_2725,N_2959);
nor U3238 (N_3238,N_2932,N_2971);
xor U3239 (N_3239,N_2989,N_2758);
and U3240 (N_3240,N_2954,N_2803);
or U3241 (N_3241,N_2555,N_2592);
nand U3242 (N_3242,N_2511,N_2501);
nand U3243 (N_3243,N_2613,N_2547);
and U3244 (N_3244,N_2844,N_2738);
or U3245 (N_3245,N_2816,N_2616);
or U3246 (N_3246,N_2796,N_2509);
nor U3247 (N_3247,N_2574,N_2663);
or U3248 (N_3248,N_2759,N_2878);
xor U3249 (N_3249,N_2726,N_2849);
or U3250 (N_3250,N_2803,N_2549);
nor U3251 (N_3251,N_2986,N_2940);
and U3252 (N_3252,N_2846,N_2720);
nand U3253 (N_3253,N_2506,N_2759);
or U3254 (N_3254,N_2645,N_2686);
nand U3255 (N_3255,N_2943,N_2617);
nor U3256 (N_3256,N_2607,N_2697);
or U3257 (N_3257,N_2679,N_2635);
or U3258 (N_3258,N_2967,N_2966);
nor U3259 (N_3259,N_2831,N_2907);
or U3260 (N_3260,N_2591,N_2932);
or U3261 (N_3261,N_2868,N_2706);
and U3262 (N_3262,N_2682,N_2752);
xor U3263 (N_3263,N_2709,N_2940);
xnor U3264 (N_3264,N_2956,N_2617);
nor U3265 (N_3265,N_2736,N_2673);
nor U3266 (N_3266,N_2578,N_2856);
nor U3267 (N_3267,N_2765,N_2537);
or U3268 (N_3268,N_2844,N_2814);
nor U3269 (N_3269,N_2945,N_2880);
nor U3270 (N_3270,N_2947,N_2809);
nand U3271 (N_3271,N_2893,N_2915);
xnor U3272 (N_3272,N_2774,N_2888);
nand U3273 (N_3273,N_2970,N_2839);
or U3274 (N_3274,N_2648,N_2765);
nand U3275 (N_3275,N_2941,N_2860);
and U3276 (N_3276,N_2555,N_2977);
and U3277 (N_3277,N_2932,N_2943);
xor U3278 (N_3278,N_2902,N_2656);
nor U3279 (N_3279,N_2529,N_2527);
xnor U3280 (N_3280,N_2892,N_2660);
or U3281 (N_3281,N_2779,N_2684);
xor U3282 (N_3282,N_2859,N_2822);
nand U3283 (N_3283,N_2763,N_2737);
nand U3284 (N_3284,N_2978,N_2675);
nand U3285 (N_3285,N_2529,N_2813);
and U3286 (N_3286,N_2546,N_2999);
nand U3287 (N_3287,N_2817,N_2796);
nand U3288 (N_3288,N_2976,N_2729);
xor U3289 (N_3289,N_2865,N_2951);
nand U3290 (N_3290,N_2788,N_2511);
and U3291 (N_3291,N_2918,N_2873);
nand U3292 (N_3292,N_2955,N_2845);
and U3293 (N_3293,N_2982,N_2636);
nand U3294 (N_3294,N_2671,N_2538);
nand U3295 (N_3295,N_2860,N_2757);
xnor U3296 (N_3296,N_2639,N_2853);
or U3297 (N_3297,N_2757,N_2737);
nand U3298 (N_3298,N_2620,N_2996);
or U3299 (N_3299,N_2760,N_2699);
nor U3300 (N_3300,N_2561,N_2665);
nand U3301 (N_3301,N_2706,N_2790);
nand U3302 (N_3302,N_2744,N_2770);
nand U3303 (N_3303,N_2945,N_2562);
nor U3304 (N_3304,N_2616,N_2760);
or U3305 (N_3305,N_2994,N_2662);
nor U3306 (N_3306,N_2602,N_2754);
xnor U3307 (N_3307,N_2962,N_2870);
and U3308 (N_3308,N_2847,N_2963);
or U3309 (N_3309,N_2701,N_2751);
and U3310 (N_3310,N_2529,N_2723);
nor U3311 (N_3311,N_2778,N_2858);
or U3312 (N_3312,N_2856,N_2992);
xnor U3313 (N_3313,N_2991,N_2527);
or U3314 (N_3314,N_2837,N_2524);
nor U3315 (N_3315,N_2850,N_2538);
xnor U3316 (N_3316,N_2686,N_2597);
and U3317 (N_3317,N_2633,N_2603);
or U3318 (N_3318,N_2639,N_2937);
or U3319 (N_3319,N_2712,N_2638);
nor U3320 (N_3320,N_2598,N_2994);
xnor U3321 (N_3321,N_2703,N_2839);
xnor U3322 (N_3322,N_2940,N_2710);
or U3323 (N_3323,N_2527,N_2763);
or U3324 (N_3324,N_2865,N_2553);
or U3325 (N_3325,N_2966,N_2535);
xor U3326 (N_3326,N_2664,N_2761);
xor U3327 (N_3327,N_2803,N_2613);
nand U3328 (N_3328,N_2584,N_2503);
xor U3329 (N_3329,N_2525,N_2504);
xnor U3330 (N_3330,N_2725,N_2976);
nand U3331 (N_3331,N_2812,N_2953);
and U3332 (N_3332,N_2779,N_2529);
nand U3333 (N_3333,N_2742,N_2934);
nand U3334 (N_3334,N_2875,N_2836);
nand U3335 (N_3335,N_2662,N_2632);
or U3336 (N_3336,N_2620,N_2952);
and U3337 (N_3337,N_2693,N_2953);
nand U3338 (N_3338,N_2731,N_2533);
or U3339 (N_3339,N_2926,N_2678);
and U3340 (N_3340,N_2501,N_2522);
xnor U3341 (N_3341,N_2663,N_2581);
and U3342 (N_3342,N_2650,N_2995);
and U3343 (N_3343,N_2588,N_2570);
and U3344 (N_3344,N_2510,N_2710);
nand U3345 (N_3345,N_2714,N_2928);
nand U3346 (N_3346,N_2843,N_2761);
and U3347 (N_3347,N_2611,N_2785);
nor U3348 (N_3348,N_2925,N_2790);
nor U3349 (N_3349,N_2691,N_2679);
nand U3350 (N_3350,N_2677,N_2727);
nor U3351 (N_3351,N_2979,N_2847);
xnor U3352 (N_3352,N_2522,N_2938);
and U3353 (N_3353,N_2721,N_2930);
and U3354 (N_3354,N_2675,N_2802);
xnor U3355 (N_3355,N_2976,N_2985);
nand U3356 (N_3356,N_2998,N_2820);
xor U3357 (N_3357,N_2562,N_2706);
or U3358 (N_3358,N_2802,N_2857);
nor U3359 (N_3359,N_2520,N_2840);
and U3360 (N_3360,N_2784,N_2514);
xnor U3361 (N_3361,N_2988,N_2978);
xnor U3362 (N_3362,N_2633,N_2817);
xnor U3363 (N_3363,N_2664,N_2644);
xnor U3364 (N_3364,N_2971,N_2777);
or U3365 (N_3365,N_2660,N_2518);
and U3366 (N_3366,N_2711,N_2609);
nor U3367 (N_3367,N_2502,N_2869);
xor U3368 (N_3368,N_2888,N_2618);
nand U3369 (N_3369,N_2909,N_2771);
and U3370 (N_3370,N_2831,N_2900);
nand U3371 (N_3371,N_2562,N_2893);
nand U3372 (N_3372,N_2902,N_2508);
or U3373 (N_3373,N_2897,N_2586);
and U3374 (N_3374,N_2990,N_2976);
and U3375 (N_3375,N_2877,N_2984);
and U3376 (N_3376,N_2995,N_2793);
nor U3377 (N_3377,N_2975,N_2925);
xnor U3378 (N_3378,N_2953,N_2918);
or U3379 (N_3379,N_2653,N_2712);
nand U3380 (N_3380,N_2874,N_2591);
and U3381 (N_3381,N_2955,N_2602);
and U3382 (N_3382,N_2835,N_2540);
or U3383 (N_3383,N_2886,N_2902);
nor U3384 (N_3384,N_2504,N_2881);
or U3385 (N_3385,N_2614,N_2508);
xor U3386 (N_3386,N_2781,N_2601);
nor U3387 (N_3387,N_2677,N_2857);
nor U3388 (N_3388,N_2598,N_2858);
and U3389 (N_3389,N_2867,N_2541);
or U3390 (N_3390,N_2685,N_2604);
or U3391 (N_3391,N_2517,N_2618);
or U3392 (N_3392,N_2913,N_2901);
nand U3393 (N_3393,N_2766,N_2859);
or U3394 (N_3394,N_2537,N_2943);
or U3395 (N_3395,N_2738,N_2717);
or U3396 (N_3396,N_2599,N_2596);
or U3397 (N_3397,N_2657,N_2543);
nor U3398 (N_3398,N_2748,N_2596);
nand U3399 (N_3399,N_2997,N_2892);
xor U3400 (N_3400,N_2512,N_2590);
nor U3401 (N_3401,N_2784,N_2967);
nor U3402 (N_3402,N_2819,N_2720);
or U3403 (N_3403,N_2599,N_2547);
nor U3404 (N_3404,N_2502,N_2846);
nor U3405 (N_3405,N_2587,N_2619);
or U3406 (N_3406,N_2684,N_2833);
and U3407 (N_3407,N_2852,N_2521);
xor U3408 (N_3408,N_2883,N_2828);
nand U3409 (N_3409,N_2740,N_2575);
nor U3410 (N_3410,N_2900,N_2545);
nand U3411 (N_3411,N_2815,N_2699);
xnor U3412 (N_3412,N_2814,N_2761);
nor U3413 (N_3413,N_2609,N_2924);
nand U3414 (N_3414,N_2572,N_2670);
nand U3415 (N_3415,N_2836,N_2966);
xnor U3416 (N_3416,N_2838,N_2537);
xnor U3417 (N_3417,N_2578,N_2758);
xnor U3418 (N_3418,N_2768,N_2750);
or U3419 (N_3419,N_2517,N_2920);
xor U3420 (N_3420,N_2854,N_2833);
nor U3421 (N_3421,N_2868,N_2893);
nand U3422 (N_3422,N_2636,N_2521);
nand U3423 (N_3423,N_2894,N_2796);
xor U3424 (N_3424,N_2878,N_2588);
and U3425 (N_3425,N_2855,N_2592);
xor U3426 (N_3426,N_2941,N_2737);
nor U3427 (N_3427,N_2995,N_2842);
and U3428 (N_3428,N_2568,N_2536);
or U3429 (N_3429,N_2513,N_2577);
and U3430 (N_3430,N_2588,N_2773);
nor U3431 (N_3431,N_2673,N_2648);
and U3432 (N_3432,N_2928,N_2907);
or U3433 (N_3433,N_2965,N_2510);
and U3434 (N_3434,N_2691,N_2846);
or U3435 (N_3435,N_2956,N_2993);
nor U3436 (N_3436,N_2557,N_2666);
or U3437 (N_3437,N_2888,N_2793);
nor U3438 (N_3438,N_2792,N_2774);
nand U3439 (N_3439,N_2854,N_2531);
and U3440 (N_3440,N_2792,N_2683);
or U3441 (N_3441,N_2653,N_2916);
nor U3442 (N_3442,N_2803,N_2809);
xnor U3443 (N_3443,N_2843,N_2844);
xnor U3444 (N_3444,N_2772,N_2740);
or U3445 (N_3445,N_2565,N_2901);
nor U3446 (N_3446,N_2861,N_2672);
xnor U3447 (N_3447,N_2897,N_2650);
xnor U3448 (N_3448,N_2533,N_2857);
or U3449 (N_3449,N_2847,N_2865);
or U3450 (N_3450,N_2513,N_2732);
and U3451 (N_3451,N_2909,N_2738);
nor U3452 (N_3452,N_2545,N_2935);
xnor U3453 (N_3453,N_2693,N_2540);
nor U3454 (N_3454,N_2888,N_2839);
or U3455 (N_3455,N_2894,N_2592);
nand U3456 (N_3456,N_2532,N_2828);
xnor U3457 (N_3457,N_2711,N_2618);
xor U3458 (N_3458,N_2927,N_2901);
nor U3459 (N_3459,N_2808,N_2770);
nand U3460 (N_3460,N_2640,N_2950);
nand U3461 (N_3461,N_2778,N_2622);
and U3462 (N_3462,N_2949,N_2877);
xnor U3463 (N_3463,N_2796,N_2708);
nand U3464 (N_3464,N_2925,N_2720);
and U3465 (N_3465,N_2766,N_2556);
nor U3466 (N_3466,N_2509,N_2748);
and U3467 (N_3467,N_2824,N_2555);
nand U3468 (N_3468,N_2873,N_2647);
and U3469 (N_3469,N_2981,N_2873);
nor U3470 (N_3470,N_2993,N_2719);
xor U3471 (N_3471,N_2929,N_2691);
and U3472 (N_3472,N_2990,N_2969);
nor U3473 (N_3473,N_2797,N_2854);
nor U3474 (N_3474,N_2726,N_2872);
and U3475 (N_3475,N_2523,N_2872);
and U3476 (N_3476,N_2557,N_2633);
xor U3477 (N_3477,N_2905,N_2981);
nor U3478 (N_3478,N_2934,N_2640);
xor U3479 (N_3479,N_2549,N_2766);
or U3480 (N_3480,N_2845,N_2605);
or U3481 (N_3481,N_2968,N_2800);
and U3482 (N_3482,N_2770,N_2967);
xor U3483 (N_3483,N_2812,N_2995);
or U3484 (N_3484,N_2519,N_2959);
nand U3485 (N_3485,N_2711,N_2675);
nand U3486 (N_3486,N_2727,N_2649);
and U3487 (N_3487,N_2859,N_2746);
nor U3488 (N_3488,N_2582,N_2993);
xor U3489 (N_3489,N_2648,N_2806);
nand U3490 (N_3490,N_2555,N_2802);
nand U3491 (N_3491,N_2969,N_2503);
nand U3492 (N_3492,N_2835,N_2787);
nor U3493 (N_3493,N_2945,N_2637);
and U3494 (N_3494,N_2813,N_2612);
or U3495 (N_3495,N_2815,N_2736);
nand U3496 (N_3496,N_2553,N_2929);
nor U3497 (N_3497,N_2666,N_2667);
xor U3498 (N_3498,N_2711,N_2919);
nor U3499 (N_3499,N_2889,N_2622);
xnor U3500 (N_3500,N_3271,N_3190);
nand U3501 (N_3501,N_3444,N_3060);
or U3502 (N_3502,N_3235,N_3031);
or U3503 (N_3503,N_3193,N_3148);
and U3504 (N_3504,N_3278,N_3414);
xnor U3505 (N_3505,N_3055,N_3230);
and U3506 (N_3506,N_3110,N_3434);
xnor U3507 (N_3507,N_3012,N_3096);
or U3508 (N_3508,N_3013,N_3435);
xor U3509 (N_3509,N_3030,N_3391);
nand U3510 (N_3510,N_3138,N_3400);
nand U3511 (N_3511,N_3036,N_3395);
nor U3512 (N_3512,N_3404,N_3184);
nor U3513 (N_3513,N_3273,N_3181);
or U3514 (N_3514,N_3267,N_3356);
or U3515 (N_3515,N_3204,N_3474);
xnor U3516 (N_3516,N_3378,N_3092);
and U3517 (N_3517,N_3363,N_3179);
and U3518 (N_3518,N_3374,N_3019);
and U3519 (N_3519,N_3208,N_3468);
nand U3520 (N_3520,N_3089,N_3216);
xor U3521 (N_3521,N_3042,N_3280);
or U3522 (N_3522,N_3021,N_3413);
xnor U3523 (N_3523,N_3088,N_3073);
nand U3524 (N_3524,N_3274,N_3197);
nor U3525 (N_3525,N_3370,N_3126);
nor U3526 (N_3526,N_3229,N_3424);
nand U3527 (N_3527,N_3102,N_3282);
xnor U3528 (N_3528,N_3082,N_3106);
and U3529 (N_3529,N_3383,N_3086);
nor U3530 (N_3530,N_3319,N_3426);
nor U3531 (N_3531,N_3209,N_3408);
and U3532 (N_3532,N_3461,N_3220);
and U3533 (N_3533,N_3382,N_3063);
and U3534 (N_3534,N_3015,N_3497);
nand U3535 (N_3535,N_3000,N_3359);
nor U3536 (N_3536,N_3168,N_3486);
nor U3537 (N_3537,N_3398,N_3344);
xnor U3538 (N_3538,N_3299,N_3456);
nor U3539 (N_3539,N_3128,N_3460);
xor U3540 (N_3540,N_3249,N_3156);
nand U3541 (N_3541,N_3058,N_3315);
nor U3542 (N_3542,N_3471,N_3134);
xnor U3543 (N_3543,N_3150,N_3105);
nor U3544 (N_3544,N_3452,N_3392);
nor U3545 (N_3545,N_3300,N_3009);
and U3546 (N_3546,N_3125,N_3357);
nand U3547 (N_3547,N_3272,N_3368);
xnor U3548 (N_3548,N_3269,N_3258);
or U3549 (N_3549,N_3473,N_3187);
or U3550 (N_3550,N_3407,N_3048);
xor U3551 (N_3551,N_3289,N_3308);
and U3552 (N_3552,N_3399,N_3045);
xor U3553 (N_3553,N_3004,N_3483);
nor U3554 (N_3554,N_3306,N_3385);
xor U3555 (N_3555,N_3244,N_3242);
and U3556 (N_3556,N_3284,N_3183);
and U3557 (N_3557,N_3131,N_3265);
nand U3558 (N_3558,N_3389,N_3120);
nand U3559 (N_3559,N_3147,N_3263);
and U3560 (N_3560,N_3039,N_3298);
nand U3561 (N_3561,N_3079,N_3354);
nor U3562 (N_3562,N_3366,N_3369);
xnor U3563 (N_3563,N_3251,N_3453);
or U3564 (N_3564,N_3341,N_3254);
xor U3565 (N_3565,N_3129,N_3260);
xor U3566 (N_3566,N_3438,N_3075);
and U3567 (N_3567,N_3051,N_3288);
nor U3568 (N_3568,N_3202,N_3117);
xnor U3569 (N_3569,N_3169,N_3401);
nand U3570 (N_3570,N_3323,N_3330);
or U3571 (N_3571,N_3499,N_3432);
nor U3572 (N_3572,N_3339,N_3264);
xnor U3573 (N_3573,N_3135,N_3171);
and U3574 (N_3574,N_3490,N_3338);
and U3575 (N_3575,N_3433,N_3320);
nand U3576 (N_3576,N_3103,N_3302);
xor U3577 (N_3577,N_3084,N_3415);
nor U3578 (N_3578,N_3478,N_3108);
nor U3579 (N_3579,N_3384,N_3314);
xnor U3580 (N_3580,N_3346,N_3480);
or U3581 (N_3581,N_3481,N_3304);
xor U3582 (N_3582,N_3018,N_3005);
or U3583 (N_3583,N_3234,N_3351);
nor U3584 (N_3584,N_3059,N_3312);
or U3585 (N_3585,N_3322,N_3146);
nand U3586 (N_3586,N_3087,N_3310);
nor U3587 (N_3587,N_3140,N_3006);
and U3588 (N_3588,N_3430,N_3397);
xor U3589 (N_3589,N_3219,N_3008);
or U3590 (N_3590,N_3163,N_3491);
or U3591 (N_3591,N_3094,N_3062);
or U3592 (N_3592,N_3028,N_3143);
or U3593 (N_3593,N_3233,N_3136);
or U3594 (N_3594,N_3071,N_3349);
or U3595 (N_3595,N_3462,N_3137);
nand U3596 (N_3596,N_3429,N_3423);
and U3597 (N_3597,N_3340,N_3159);
xnor U3598 (N_3598,N_3227,N_3095);
nand U3599 (N_3599,N_3494,N_3056);
and U3600 (N_3600,N_3033,N_3498);
xnor U3601 (N_3601,N_3119,N_3180);
nand U3602 (N_3602,N_3248,N_3281);
xor U3603 (N_3603,N_3287,N_3333);
xnor U3604 (N_3604,N_3166,N_3017);
xnor U3605 (N_3605,N_3081,N_3161);
or U3606 (N_3606,N_3172,N_3296);
xnor U3607 (N_3607,N_3457,N_3224);
and U3608 (N_3608,N_3492,N_3182);
xor U3609 (N_3609,N_3077,N_3029);
nand U3610 (N_3610,N_3052,N_3201);
xor U3611 (N_3611,N_3164,N_3044);
or U3612 (N_3612,N_3297,N_3170);
xnor U3613 (N_3613,N_3205,N_3101);
xor U3614 (N_3614,N_3353,N_3294);
xnor U3615 (N_3615,N_3218,N_3212);
and U3616 (N_3616,N_3417,N_3347);
or U3617 (N_3617,N_3348,N_3065);
or U3618 (N_3618,N_3213,N_3496);
nor U3619 (N_3619,N_3231,N_3266);
or U3620 (N_3620,N_3074,N_3214);
xor U3621 (N_3621,N_3091,N_3387);
or U3622 (N_3622,N_3325,N_3343);
or U3623 (N_3623,N_3098,N_3449);
and U3624 (N_3624,N_3243,N_3240);
nor U3625 (N_3625,N_3291,N_3097);
nand U3626 (N_3626,N_3145,N_3355);
or U3627 (N_3627,N_3293,N_3425);
nand U3628 (N_3628,N_3286,N_3114);
or U3629 (N_3629,N_3035,N_3165);
xor U3630 (N_3630,N_3495,N_3024);
nand U3631 (N_3631,N_3133,N_3199);
and U3632 (N_3632,N_3144,N_3157);
xor U3633 (N_3633,N_3406,N_3459);
xor U3634 (N_3634,N_3023,N_3437);
nor U3635 (N_3635,N_3151,N_3041);
xor U3636 (N_3636,N_3203,N_3283);
nor U3637 (N_3637,N_3100,N_3107);
xnor U3638 (N_3638,N_3270,N_3371);
and U3639 (N_3639,N_3379,N_3447);
and U3640 (N_3640,N_3443,N_3390);
nor U3641 (N_3641,N_3068,N_3111);
xor U3642 (N_3642,N_3475,N_3345);
nand U3643 (N_3643,N_3334,N_3332);
and U3644 (N_3644,N_3466,N_3022);
xor U3645 (N_3645,N_3442,N_3259);
or U3646 (N_3646,N_3317,N_3295);
or U3647 (N_3647,N_3307,N_3255);
nand U3648 (N_3648,N_3275,N_3403);
nor U3649 (N_3649,N_3217,N_3245);
or U3650 (N_3650,N_3350,N_3421);
and U3651 (N_3651,N_3064,N_3153);
nand U3652 (N_3652,N_3050,N_3123);
xor U3653 (N_3653,N_3301,N_3313);
nand U3654 (N_3654,N_3493,N_3223);
nor U3655 (N_3655,N_3309,N_3207);
xor U3656 (N_3656,N_3477,N_3253);
xor U3657 (N_3657,N_3388,N_3487);
xnor U3658 (N_3658,N_3149,N_3215);
nor U3659 (N_3659,N_3049,N_3104);
or U3660 (N_3660,N_3246,N_3198);
xor U3661 (N_3661,N_3321,N_3154);
or U3662 (N_3662,N_3011,N_3311);
or U3663 (N_3663,N_3232,N_3364);
nand U3664 (N_3664,N_3465,N_3228);
or U3665 (N_3665,N_3003,N_3458);
nand U3666 (N_3666,N_3191,N_3372);
or U3667 (N_3667,N_3200,N_3099);
and U3668 (N_3668,N_3276,N_3410);
nand U3669 (N_3669,N_3416,N_3152);
nor U3670 (N_3670,N_3196,N_3360);
or U3671 (N_3671,N_3451,N_3377);
xor U3672 (N_3672,N_3115,N_3085);
or U3673 (N_3673,N_3327,N_3130);
and U3674 (N_3674,N_3122,N_3422);
and U3675 (N_3675,N_3155,N_3448);
xnor U3676 (N_3676,N_3427,N_3303);
and U3677 (N_3677,N_3194,N_3489);
or U3678 (N_3678,N_3070,N_3026);
nor U3679 (N_3679,N_3192,N_3261);
nand U3680 (N_3680,N_3305,N_3221);
or U3681 (N_3681,N_3066,N_3047);
or U3682 (N_3682,N_3210,N_3160);
and U3683 (N_3683,N_3464,N_3057);
xor U3684 (N_3684,N_3083,N_3211);
nand U3685 (N_3685,N_3257,N_3080);
xnor U3686 (N_3686,N_3316,N_3419);
nand U3687 (N_3687,N_3436,N_3185);
and U3688 (N_3688,N_3329,N_3420);
and U3689 (N_3689,N_3020,N_3124);
and U3690 (N_3690,N_3186,N_3001);
or U3691 (N_3691,N_3040,N_3409);
nor U3692 (N_3692,N_3237,N_3236);
xnor U3693 (N_3693,N_3162,N_3027);
nor U3694 (N_3694,N_3290,N_3174);
xor U3695 (N_3695,N_3337,N_3158);
and U3696 (N_3696,N_3470,N_3336);
nor U3697 (N_3697,N_3440,N_3324);
nor U3698 (N_3698,N_3238,N_3446);
nand U3699 (N_3699,N_3239,N_3484);
nand U3700 (N_3700,N_3431,N_3241);
nor U3701 (N_3701,N_3141,N_3279);
xnor U3702 (N_3702,N_3375,N_3488);
nand U3703 (N_3703,N_3247,N_3445);
xor U3704 (N_3704,N_3331,N_3454);
and U3705 (N_3705,N_3076,N_3121);
and U3706 (N_3706,N_3127,N_3176);
and U3707 (N_3707,N_3467,N_3318);
nand U3708 (N_3708,N_3376,N_3439);
and U3709 (N_3709,N_3002,N_3469);
nor U3710 (N_3710,N_3093,N_3195);
nor U3711 (N_3711,N_3472,N_3016);
nand U3712 (N_3712,N_3373,N_3078);
nand U3713 (N_3713,N_3067,N_3034);
and U3714 (N_3714,N_3173,N_3352);
xnor U3715 (N_3715,N_3367,N_3118);
nor U3716 (N_3716,N_3428,N_3268);
and U3717 (N_3717,N_3393,N_3010);
xnor U3718 (N_3718,N_3256,N_3225);
xor U3719 (N_3719,N_3476,N_3365);
and U3720 (N_3720,N_3116,N_3277);
xnor U3721 (N_3721,N_3032,N_3380);
or U3722 (N_3722,N_3188,N_3479);
and U3723 (N_3723,N_3342,N_3054);
xor U3724 (N_3724,N_3222,N_3412);
nor U3725 (N_3725,N_3038,N_3043);
and U3726 (N_3726,N_3167,N_3482);
or U3727 (N_3727,N_3069,N_3328);
or U3728 (N_3728,N_3046,N_3061);
and U3729 (N_3729,N_3485,N_3292);
or U3730 (N_3730,N_3007,N_3177);
or U3731 (N_3731,N_3139,N_3335);
nor U3732 (N_3732,N_3142,N_3025);
or U3733 (N_3733,N_3411,N_3014);
nor U3734 (N_3734,N_3381,N_3418);
xor U3735 (N_3735,N_3112,N_3441);
and U3736 (N_3736,N_3132,N_3386);
nor U3737 (N_3737,N_3405,N_3037);
xnor U3738 (N_3738,N_3175,N_3189);
xnor U3739 (N_3739,N_3455,N_3262);
or U3740 (N_3740,N_3285,N_3358);
nand U3741 (N_3741,N_3109,N_3463);
nor U3742 (N_3742,N_3252,N_3072);
and U3743 (N_3743,N_3053,N_3402);
xor U3744 (N_3744,N_3450,N_3394);
nor U3745 (N_3745,N_3206,N_3396);
nor U3746 (N_3746,N_3362,N_3226);
xor U3747 (N_3747,N_3326,N_3090);
or U3748 (N_3748,N_3178,N_3113);
nor U3749 (N_3749,N_3361,N_3250);
and U3750 (N_3750,N_3276,N_3387);
nand U3751 (N_3751,N_3067,N_3102);
nand U3752 (N_3752,N_3028,N_3415);
nand U3753 (N_3753,N_3006,N_3100);
and U3754 (N_3754,N_3454,N_3261);
or U3755 (N_3755,N_3458,N_3082);
xnor U3756 (N_3756,N_3114,N_3089);
nand U3757 (N_3757,N_3211,N_3119);
nand U3758 (N_3758,N_3005,N_3213);
or U3759 (N_3759,N_3033,N_3223);
and U3760 (N_3760,N_3016,N_3001);
nor U3761 (N_3761,N_3257,N_3110);
xnor U3762 (N_3762,N_3094,N_3135);
nor U3763 (N_3763,N_3471,N_3140);
nor U3764 (N_3764,N_3197,N_3118);
xor U3765 (N_3765,N_3038,N_3149);
and U3766 (N_3766,N_3418,N_3439);
or U3767 (N_3767,N_3043,N_3408);
or U3768 (N_3768,N_3410,N_3123);
nand U3769 (N_3769,N_3190,N_3399);
nor U3770 (N_3770,N_3454,N_3345);
nor U3771 (N_3771,N_3293,N_3383);
and U3772 (N_3772,N_3465,N_3377);
and U3773 (N_3773,N_3437,N_3331);
nor U3774 (N_3774,N_3163,N_3196);
and U3775 (N_3775,N_3010,N_3387);
and U3776 (N_3776,N_3286,N_3429);
xor U3777 (N_3777,N_3030,N_3157);
nand U3778 (N_3778,N_3183,N_3213);
xor U3779 (N_3779,N_3193,N_3000);
xor U3780 (N_3780,N_3427,N_3137);
xnor U3781 (N_3781,N_3337,N_3348);
nor U3782 (N_3782,N_3278,N_3319);
or U3783 (N_3783,N_3441,N_3156);
nand U3784 (N_3784,N_3245,N_3239);
and U3785 (N_3785,N_3001,N_3003);
nand U3786 (N_3786,N_3197,N_3237);
nand U3787 (N_3787,N_3266,N_3107);
nor U3788 (N_3788,N_3071,N_3348);
or U3789 (N_3789,N_3382,N_3053);
xnor U3790 (N_3790,N_3278,N_3498);
nand U3791 (N_3791,N_3067,N_3008);
or U3792 (N_3792,N_3034,N_3196);
xor U3793 (N_3793,N_3497,N_3259);
and U3794 (N_3794,N_3261,N_3249);
nor U3795 (N_3795,N_3277,N_3375);
and U3796 (N_3796,N_3262,N_3425);
nor U3797 (N_3797,N_3444,N_3080);
nor U3798 (N_3798,N_3454,N_3334);
nand U3799 (N_3799,N_3444,N_3045);
or U3800 (N_3800,N_3358,N_3224);
nor U3801 (N_3801,N_3232,N_3053);
and U3802 (N_3802,N_3111,N_3333);
or U3803 (N_3803,N_3292,N_3147);
xnor U3804 (N_3804,N_3105,N_3440);
or U3805 (N_3805,N_3387,N_3083);
xnor U3806 (N_3806,N_3264,N_3244);
nand U3807 (N_3807,N_3075,N_3123);
and U3808 (N_3808,N_3166,N_3425);
and U3809 (N_3809,N_3326,N_3022);
nand U3810 (N_3810,N_3189,N_3492);
or U3811 (N_3811,N_3121,N_3346);
nand U3812 (N_3812,N_3046,N_3098);
or U3813 (N_3813,N_3327,N_3474);
nor U3814 (N_3814,N_3179,N_3464);
and U3815 (N_3815,N_3479,N_3478);
xnor U3816 (N_3816,N_3176,N_3095);
or U3817 (N_3817,N_3250,N_3029);
xnor U3818 (N_3818,N_3456,N_3270);
or U3819 (N_3819,N_3186,N_3156);
nor U3820 (N_3820,N_3348,N_3216);
or U3821 (N_3821,N_3412,N_3391);
or U3822 (N_3822,N_3415,N_3150);
nor U3823 (N_3823,N_3140,N_3493);
or U3824 (N_3824,N_3127,N_3009);
xnor U3825 (N_3825,N_3095,N_3140);
nand U3826 (N_3826,N_3187,N_3324);
nor U3827 (N_3827,N_3091,N_3039);
nand U3828 (N_3828,N_3433,N_3212);
xor U3829 (N_3829,N_3254,N_3434);
nor U3830 (N_3830,N_3452,N_3256);
xnor U3831 (N_3831,N_3301,N_3062);
nand U3832 (N_3832,N_3448,N_3046);
or U3833 (N_3833,N_3072,N_3274);
nand U3834 (N_3834,N_3499,N_3293);
and U3835 (N_3835,N_3047,N_3439);
or U3836 (N_3836,N_3205,N_3111);
nor U3837 (N_3837,N_3002,N_3340);
xor U3838 (N_3838,N_3367,N_3026);
and U3839 (N_3839,N_3109,N_3188);
and U3840 (N_3840,N_3089,N_3146);
xor U3841 (N_3841,N_3114,N_3422);
xor U3842 (N_3842,N_3235,N_3187);
nand U3843 (N_3843,N_3068,N_3218);
xor U3844 (N_3844,N_3122,N_3366);
and U3845 (N_3845,N_3129,N_3474);
nand U3846 (N_3846,N_3391,N_3321);
nand U3847 (N_3847,N_3184,N_3096);
or U3848 (N_3848,N_3455,N_3458);
xnor U3849 (N_3849,N_3076,N_3216);
nor U3850 (N_3850,N_3211,N_3093);
or U3851 (N_3851,N_3431,N_3020);
nand U3852 (N_3852,N_3463,N_3023);
xor U3853 (N_3853,N_3176,N_3498);
xor U3854 (N_3854,N_3428,N_3277);
nand U3855 (N_3855,N_3253,N_3240);
nor U3856 (N_3856,N_3484,N_3123);
and U3857 (N_3857,N_3018,N_3141);
nand U3858 (N_3858,N_3037,N_3054);
xnor U3859 (N_3859,N_3157,N_3390);
nor U3860 (N_3860,N_3084,N_3073);
nand U3861 (N_3861,N_3044,N_3321);
xor U3862 (N_3862,N_3380,N_3464);
nor U3863 (N_3863,N_3273,N_3438);
or U3864 (N_3864,N_3293,N_3183);
nor U3865 (N_3865,N_3135,N_3357);
nand U3866 (N_3866,N_3331,N_3022);
xnor U3867 (N_3867,N_3129,N_3259);
and U3868 (N_3868,N_3469,N_3100);
nand U3869 (N_3869,N_3390,N_3136);
and U3870 (N_3870,N_3108,N_3176);
xor U3871 (N_3871,N_3015,N_3352);
nand U3872 (N_3872,N_3357,N_3496);
and U3873 (N_3873,N_3298,N_3018);
xor U3874 (N_3874,N_3381,N_3164);
and U3875 (N_3875,N_3144,N_3423);
nor U3876 (N_3876,N_3480,N_3461);
nand U3877 (N_3877,N_3061,N_3488);
nor U3878 (N_3878,N_3249,N_3263);
and U3879 (N_3879,N_3393,N_3170);
or U3880 (N_3880,N_3035,N_3300);
nand U3881 (N_3881,N_3226,N_3365);
and U3882 (N_3882,N_3083,N_3230);
or U3883 (N_3883,N_3468,N_3038);
and U3884 (N_3884,N_3451,N_3101);
and U3885 (N_3885,N_3048,N_3386);
and U3886 (N_3886,N_3083,N_3218);
or U3887 (N_3887,N_3385,N_3467);
or U3888 (N_3888,N_3395,N_3332);
nor U3889 (N_3889,N_3472,N_3400);
xor U3890 (N_3890,N_3165,N_3005);
nand U3891 (N_3891,N_3214,N_3324);
or U3892 (N_3892,N_3101,N_3029);
or U3893 (N_3893,N_3329,N_3470);
xor U3894 (N_3894,N_3398,N_3482);
nand U3895 (N_3895,N_3203,N_3141);
nand U3896 (N_3896,N_3178,N_3025);
nor U3897 (N_3897,N_3431,N_3098);
nor U3898 (N_3898,N_3318,N_3234);
or U3899 (N_3899,N_3036,N_3385);
or U3900 (N_3900,N_3102,N_3386);
xor U3901 (N_3901,N_3174,N_3381);
and U3902 (N_3902,N_3342,N_3011);
xor U3903 (N_3903,N_3344,N_3443);
nor U3904 (N_3904,N_3081,N_3349);
nor U3905 (N_3905,N_3230,N_3145);
nand U3906 (N_3906,N_3324,N_3276);
xor U3907 (N_3907,N_3492,N_3340);
and U3908 (N_3908,N_3206,N_3095);
xnor U3909 (N_3909,N_3249,N_3321);
xnor U3910 (N_3910,N_3167,N_3237);
and U3911 (N_3911,N_3260,N_3341);
nand U3912 (N_3912,N_3429,N_3344);
nand U3913 (N_3913,N_3026,N_3254);
and U3914 (N_3914,N_3495,N_3001);
and U3915 (N_3915,N_3408,N_3205);
or U3916 (N_3916,N_3364,N_3074);
or U3917 (N_3917,N_3331,N_3088);
nand U3918 (N_3918,N_3133,N_3282);
and U3919 (N_3919,N_3371,N_3257);
nand U3920 (N_3920,N_3140,N_3025);
nand U3921 (N_3921,N_3358,N_3448);
nor U3922 (N_3922,N_3382,N_3463);
xor U3923 (N_3923,N_3257,N_3165);
or U3924 (N_3924,N_3485,N_3070);
xnor U3925 (N_3925,N_3471,N_3234);
or U3926 (N_3926,N_3219,N_3235);
xnor U3927 (N_3927,N_3388,N_3054);
nand U3928 (N_3928,N_3327,N_3188);
and U3929 (N_3929,N_3328,N_3095);
nor U3930 (N_3930,N_3432,N_3421);
xnor U3931 (N_3931,N_3096,N_3273);
and U3932 (N_3932,N_3065,N_3372);
nor U3933 (N_3933,N_3123,N_3417);
nand U3934 (N_3934,N_3339,N_3185);
nor U3935 (N_3935,N_3421,N_3368);
or U3936 (N_3936,N_3020,N_3458);
and U3937 (N_3937,N_3159,N_3316);
or U3938 (N_3938,N_3141,N_3393);
nand U3939 (N_3939,N_3420,N_3255);
nand U3940 (N_3940,N_3449,N_3082);
nor U3941 (N_3941,N_3235,N_3314);
xnor U3942 (N_3942,N_3044,N_3066);
or U3943 (N_3943,N_3008,N_3337);
nand U3944 (N_3944,N_3325,N_3296);
xor U3945 (N_3945,N_3175,N_3239);
xor U3946 (N_3946,N_3370,N_3109);
nor U3947 (N_3947,N_3414,N_3444);
nand U3948 (N_3948,N_3447,N_3498);
xor U3949 (N_3949,N_3478,N_3080);
nand U3950 (N_3950,N_3341,N_3402);
or U3951 (N_3951,N_3249,N_3190);
or U3952 (N_3952,N_3489,N_3223);
or U3953 (N_3953,N_3111,N_3044);
or U3954 (N_3954,N_3235,N_3152);
or U3955 (N_3955,N_3199,N_3187);
nor U3956 (N_3956,N_3190,N_3356);
or U3957 (N_3957,N_3486,N_3050);
and U3958 (N_3958,N_3269,N_3457);
and U3959 (N_3959,N_3465,N_3411);
nor U3960 (N_3960,N_3382,N_3417);
nand U3961 (N_3961,N_3451,N_3415);
nand U3962 (N_3962,N_3120,N_3376);
nor U3963 (N_3963,N_3295,N_3090);
or U3964 (N_3964,N_3321,N_3470);
and U3965 (N_3965,N_3000,N_3170);
or U3966 (N_3966,N_3217,N_3134);
or U3967 (N_3967,N_3315,N_3020);
nor U3968 (N_3968,N_3388,N_3078);
and U3969 (N_3969,N_3314,N_3295);
xnor U3970 (N_3970,N_3212,N_3094);
xor U3971 (N_3971,N_3404,N_3185);
xnor U3972 (N_3972,N_3094,N_3140);
xor U3973 (N_3973,N_3130,N_3412);
or U3974 (N_3974,N_3126,N_3016);
and U3975 (N_3975,N_3438,N_3267);
xnor U3976 (N_3976,N_3333,N_3398);
nor U3977 (N_3977,N_3472,N_3219);
or U3978 (N_3978,N_3019,N_3216);
xor U3979 (N_3979,N_3000,N_3098);
and U3980 (N_3980,N_3420,N_3238);
or U3981 (N_3981,N_3413,N_3294);
nand U3982 (N_3982,N_3144,N_3465);
or U3983 (N_3983,N_3404,N_3498);
nand U3984 (N_3984,N_3115,N_3219);
nor U3985 (N_3985,N_3453,N_3142);
nand U3986 (N_3986,N_3296,N_3380);
xor U3987 (N_3987,N_3118,N_3434);
xor U3988 (N_3988,N_3360,N_3078);
nand U3989 (N_3989,N_3154,N_3211);
or U3990 (N_3990,N_3319,N_3122);
and U3991 (N_3991,N_3224,N_3363);
nand U3992 (N_3992,N_3271,N_3237);
and U3993 (N_3993,N_3382,N_3147);
or U3994 (N_3994,N_3270,N_3473);
or U3995 (N_3995,N_3242,N_3051);
and U3996 (N_3996,N_3386,N_3252);
nand U3997 (N_3997,N_3025,N_3400);
nand U3998 (N_3998,N_3053,N_3103);
nand U3999 (N_3999,N_3249,N_3027);
or U4000 (N_4000,N_3524,N_3838);
nand U4001 (N_4001,N_3741,N_3600);
and U4002 (N_4002,N_3509,N_3546);
and U4003 (N_4003,N_3749,N_3816);
and U4004 (N_4004,N_3672,N_3852);
nand U4005 (N_4005,N_3865,N_3963);
and U4006 (N_4006,N_3573,N_3925);
nor U4007 (N_4007,N_3800,N_3947);
nand U4008 (N_4008,N_3715,N_3647);
or U4009 (N_4009,N_3578,N_3878);
nand U4010 (N_4010,N_3751,N_3984);
xor U4011 (N_4011,N_3643,N_3784);
nor U4012 (N_4012,N_3683,N_3762);
nor U4013 (N_4013,N_3532,N_3894);
nor U4014 (N_4014,N_3540,N_3607);
or U4015 (N_4015,N_3661,N_3697);
nand U4016 (N_4016,N_3767,N_3864);
nor U4017 (N_4017,N_3732,N_3632);
xnor U4018 (N_4018,N_3770,N_3854);
nor U4019 (N_4019,N_3623,N_3620);
xor U4020 (N_4020,N_3863,N_3805);
xnor U4021 (N_4021,N_3610,N_3811);
and U4022 (N_4022,N_3669,N_3660);
nor U4023 (N_4023,N_3765,N_3750);
nand U4024 (N_4024,N_3889,N_3618);
xor U4025 (N_4025,N_3847,N_3659);
xnor U4026 (N_4026,N_3735,N_3710);
xnor U4027 (N_4027,N_3917,N_3849);
and U4028 (N_4028,N_3818,N_3827);
and U4029 (N_4029,N_3588,N_3909);
and U4030 (N_4030,N_3568,N_3712);
xor U4031 (N_4031,N_3996,N_3569);
and U4032 (N_4032,N_3918,N_3884);
xor U4033 (N_4033,N_3676,N_3929);
xnor U4034 (N_4034,N_3612,N_3558);
nor U4035 (N_4035,N_3948,N_3738);
nor U4036 (N_4036,N_3557,N_3763);
nand U4037 (N_4037,N_3862,N_3615);
and U4038 (N_4038,N_3571,N_3550);
nor U4039 (N_4039,N_3678,N_3512);
and U4040 (N_4040,N_3761,N_3914);
nor U4041 (N_4041,N_3686,N_3820);
and U4042 (N_4042,N_3562,N_3629);
nor U4043 (N_4043,N_3528,N_3788);
and U4044 (N_4044,N_3902,N_3961);
and U4045 (N_4045,N_3874,N_3802);
or U4046 (N_4046,N_3544,N_3664);
nand U4047 (N_4047,N_3783,N_3891);
nor U4048 (N_4048,N_3979,N_3570);
nand U4049 (N_4049,N_3527,N_3823);
and U4050 (N_4050,N_3752,N_3628);
nand U4051 (N_4051,N_3760,N_3791);
and U4052 (N_4052,N_3631,N_3911);
and U4053 (N_4053,N_3641,N_3966);
nor U4054 (N_4054,N_3590,N_3535);
and U4055 (N_4055,N_3598,N_3614);
nor U4056 (N_4056,N_3725,N_3837);
or U4057 (N_4057,N_3679,N_3775);
nand U4058 (N_4058,N_3815,N_3968);
xnor U4059 (N_4059,N_3936,N_3690);
or U4060 (N_4060,N_3939,N_3642);
nand U4061 (N_4061,N_3873,N_3807);
xor U4062 (N_4062,N_3887,N_3638);
nand U4063 (N_4063,N_3727,N_3764);
xnor U4064 (N_4064,N_3539,N_3603);
nand U4065 (N_4065,N_3988,N_3531);
xor U4066 (N_4066,N_3995,N_3594);
and U4067 (N_4067,N_3700,N_3699);
or U4068 (N_4068,N_3688,N_3771);
or U4069 (N_4069,N_3583,N_3604);
or U4070 (N_4070,N_3541,N_3739);
and U4071 (N_4071,N_3626,N_3759);
nand U4072 (N_4072,N_3658,N_3513);
or U4073 (N_4073,N_3844,N_3648);
nand U4074 (N_4074,N_3500,N_3876);
and U4075 (N_4075,N_3713,N_3855);
xnor U4076 (N_4076,N_3919,N_3987);
or U4077 (N_4077,N_3722,N_3799);
and U4078 (N_4078,N_3885,N_3935);
and U4079 (N_4079,N_3962,N_3662);
nor U4080 (N_4080,N_3960,N_3542);
nand U4081 (N_4081,N_3880,N_3976);
xor U4082 (N_4082,N_3729,N_3843);
nor U4083 (N_4083,N_3814,N_3942);
nand U4084 (N_4084,N_3768,N_3621);
nand U4085 (N_4085,N_3674,N_3602);
or U4086 (N_4086,N_3893,N_3908);
or U4087 (N_4087,N_3684,N_3521);
nor U4088 (N_4088,N_3834,N_3687);
and U4089 (N_4089,N_3515,N_3754);
nor U4090 (N_4090,N_3755,N_3666);
or U4091 (N_4091,N_3655,N_3582);
xor U4092 (N_4092,N_3986,N_3696);
and U4093 (N_4093,N_3653,N_3913);
nor U4094 (N_4094,N_3813,N_3910);
and U4095 (N_4095,N_3506,N_3974);
xor U4096 (N_4096,N_3777,N_3912);
and U4097 (N_4097,N_3786,N_3907);
nand U4098 (N_4098,N_3766,N_3959);
nor U4099 (N_4099,N_3932,N_3575);
and U4100 (N_4100,N_3999,N_3915);
or U4101 (N_4101,N_3740,N_3957);
nand U4102 (N_4102,N_3845,N_3654);
or U4103 (N_4103,N_3585,N_3599);
xnor U4104 (N_4104,N_3746,N_3776);
nand U4105 (N_4105,N_3572,N_3983);
nor U4106 (N_4106,N_3790,N_3523);
xnor U4107 (N_4107,N_3703,N_3903);
and U4108 (N_4108,N_3778,N_3870);
xor U4109 (N_4109,N_3529,N_3596);
nand U4110 (N_4110,N_3730,N_3501);
or U4111 (N_4111,N_3677,N_3720);
xnor U4112 (N_4112,N_3724,N_3559);
xor U4113 (N_4113,N_3923,N_3850);
or U4114 (N_4114,N_3973,N_3704);
nand U4115 (N_4115,N_3905,N_3906);
nand U4116 (N_4116,N_3519,N_3692);
nor U4117 (N_4117,N_3969,N_3920);
nand U4118 (N_4118,N_3639,N_3736);
or U4119 (N_4119,N_3924,N_3787);
nand U4120 (N_4120,N_3517,N_3990);
and U4121 (N_4121,N_3747,N_3993);
or U4122 (N_4122,N_3944,N_3680);
xnor U4123 (N_4123,N_3636,N_3848);
or U4124 (N_4124,N_3797,N_3556);
nand U4125 (N_4125,N_3756,N_3507);
and U4126 (N_4126,N_3856,N_3931);
xnor U4127 (N_4127,N_3955,N_3671);
xor U4128 (N_4128,N_3866,N_3812);
xnor U4129 (N_4129,N_3933,N_3789);
nor U4130 (N_4130,N_3564,N_3548);
and U4131 (N_4131,N_3792,N_3956);
and U4132 (N_4132,N_3657,N_3928);
nor U4133 (N_4133,N_3637,N_3951);
or U4134 (N_4134,N_3625,N_3875);
xnor U4135 (N_4135,N_3890,N_3744);
or U4136 (N_4136,N_3796,N_3613);
xor U4137 (N_4137,N_3971,N_3576);
or U4138 (N_4138,N_3719,N_3565);
and U4139 (N_4139,N_3581,N_3930);
nor U4140 (N_4140,N_3707,N_3616);
xor U4141 (N_4141,N_3773,N_3742);
xnor U4142 (N_4142,N_3520,N_3921);
and U4143 (N_4143,N_3701,N_3868);
nand U4144 (N_4144,N_3842,N_3651);
xor U4145 (N_4145,N_3593,N_3592);
or U4146 (N_4146,N_3859,N_3645);
xnor U4147 (N_4147,N_3977,N_3882);
and U4148 (N_4148,N_3927,N_3832);
or U4149 (N_4149,N_3934,N_3525);
xor U4150 (N_4150,N_3922,N_3808);
or U4151 (N_4151,N_3597,N_3897);
nor U4152 (N_4152,N_3649,N_3619);
xnor U4153 (N_4153,N_3846,N_3817);
nor U4154 (N_4154,N_3860,N_3691);
nand U4155 (N_4155,N_3985,N_3718);
and U4156 (N_4156,N_3839,N_3904);
or U4157 (N_4157,N_3980,N_3526);
or U4158 (N_4158,N_3705,N_3505);
nand U4159 (N_4159,N_3627,N_3693);
xnor U4160 (N_4160,N_3728,N_3634);
nand U4161 (N_4161,N_3853,N_3609);
nand U4162 (N_4162,N_3950,N_3745);
and U4163 (N_4163,N_3561,N_3534);
xnor U4164 (N_4164,N_3861,N_3895);
nor U4165 (N_4165,N_3538,N_3698);
nand U4166 (N_4166,N_3835,N_3685);
nand U4167 (N_4167,N_3668,N_3709);
nor U4168 (N_4168,N_3551,N_3958);
xor U4169 (N_4169,N_3833,N_3617);
xnor U4170 (N_4170,N_3731,N_3586);
xor U4171 (N_4171,N_3563,N_3896);
xnor U4172 (N_4172,N_3926,N_3809);
nand U4173 (N_4173,N_3667,N_3716);
and U4174 (N_4174,N_3821,N_3978);
nor U4175 (N_4175,N_3946,N_3721);
nor U4176 (N_4176,N_3587,N_3536);
or U4177 (N_4177,N_3781,N_3872);
and U4178 (N_4178,N_3970,N_3769);
nand U4179 (N_4179,N_3967,N_3656);
and U4180 (N_4180,N_3810,N_3595);
and U4181 (N_4181,N_3530,N_3577);
xnor U4182 (N_4182,N_3841,N_3591);
and U4183 (N_4183,N_3989,N_3819);
nor U4184 (N_4184,N_3916,N_3886);
nand U4185 (N_4185,N_3567,N_3549);
and U4186 (N_4186,N_3605,N_3840);
nand U4187 (N_4187,N_3574,N_3555);
and U4188 (N_4188,N_3682,N_3825);
nand U4189 (N_4189,N_3622,N_3652);
or U4190 (N_4190,N_3714,N_3734);
xor U4191 (N_4191,N_3793,N_3836);
nor U4192 (N_4192,N_3782,N_3611);
nor U4193 (N_4193,N_3824,N_3514);
nand U4194 (N_4194,N_3829,N_3552);
or U4195 (N_4195,N_3795,N_3547);
nor U4196 (N_4196,N_3780,N_3892);
nand U4197 (N_4197,N_3537,N_3624);
or U4198 (N_4198,N_3806,N_3723);
or U4199 (N_4199,N_3871,N_3994);
nand U4200 (N_4200,N_3997,N_3580);
xnor U4201 (N_4201,N_3516,N_3898);
nor U4202 (N_4202,N_3560,N_3681);
or U4203 (N_4203,N_3826,N_3689);
or U4204 (N_4204,N_3804,N_3635);
and U4205 (N_4205,N_3937,N_3608);
or U4206 (N_4206,N_3579,N_3758);
and U4207 (N_4207,N_3803,N_3901);
nor U4208 (N_4208,N_3858,N_3899);
nand U4209 (N_4209,N_3589,N_3828);
nor U4210 (N_4210,N_3522,N_3772);
nand U4211 (N_4211,N_3982,N_3774);
nor U4212 (N_4212,N_3566,N_3553);
xnor U4213 (N_4213,N_3708,N_3831);
and U4214 (N_4214,N_3867,N_3633);
and U4215 (N_4215,N_3801,N_3943);
or U4216 (N_4216,N_3508,N_3941);
nand U4217 (N_4217,N_3601,N_3952);
and U4218 (N_4218,N_3665,N_3881);
xor U4219 (N_4219,N_3964,N_3794);
nand U4220 (N_4220,N_3543,N_3733);
and U4221 (N_4221,N_3830,N_3822);
nor U4222 (N_4222,N_3981,N_3554);
nand U4223 (N_4223,N_3533,N_3972);
nand U4224 (N_4224,N_3851,N_3877);
nor U4225 (N_4225,N_3757,N_3644);
nor U4226 (N_4226,N_3646,N_3503);
and U4227 (N_4227,N_3753,N_3584);
nor U4228 (N_4228,N_3663,N_3900);
and U4229 (N_4229,N_3945,N_3949);
and U4230 (N_4230,N_3857,N_3938);
or U4231 (N_4231,N_3511,N_3726);
nand U4232 (N_4232,N_3695,N_3954);
xor U4233 (N_4233,N_3975,N_3883);
and U4234 (N_4234,N_3702,N_3953);
and U4235 (N_4235,N_3510,N_3706);
xnor U4236 (N_4236,N_3694,N_3998);
nor U4237 (N_4237,N_3545,N_3630);
nor U4238 (N_4238,N_3606,N_3717);
and U4239 (N_4239,N_3743,N_3879);
nor U4240 (N_4240,N_3504,N_3992);
xnor U4241 (N_4241,N_3798,N_3940);
xnor U4242 (N_4242,N_3650,N_3518);
nand U4243 (N_4243,N_3673,N_3748);
and U4244 (N_4244,N_3779,N_3869);
and U4245 (N_4245,N_3991,N_3888);
nand U4246 (N_4246,N_3640,N_3737);
and U4247 (N_4247,N_3711,N_3502);
and U4248 (N_4248,N_3965,N_3675);
or U4249 (N_4249,N_3785,N_3670);
nor U4250 (N_4250,N_3565,N_3540);
nor U4251 (N_4251,N_3806,N_3563);
or U4252 (N_4252,N_3707,N_3975);
xor U4253 (N_4253,N_3587,N_3588);
nor U4254 (N_4254,N_3868,N_3711);
and U4255 (N_4255,N_3872,N_3786);
nand U4256 (N_4256,N_3703,N_3879);
or U4257 (N_4257,N_3572,N_3513);
xor U4258 (N_4258,N_3610,N_3803);
nand U4259 (N_4259,N_3782,N_3883);
nand U4260 (N_4260,N_3897,N_3674);
or U4261 (N_4261,N_3628,N_3507);
or U4262 (N_4262,N_3515,N_3630);
and U4263 (N_4263,N_3853,N_3983);
nor U4264 (N_4264,N_3741,N_3595);
xor U4265 (N_4265,N_3895,N_3776);
nand U4266 (N_4266,N_3825,N_3803);
and U4267 (N_4267,N_3983,N_3596);
or U4268 (N_4268,N_3504,N_3580);
or U4269 (N_4269,N_3631,N_3967);
xnor U4270 (N_4270,N_3566,N_3942);
nand U4271 (N_4271,N_3627,N_3886);
and U4272 (N_4272,N_3586,N_3722);
and U4273 (N_4273,N_3659,N_3517);
and U4274 (N_4274,N_3943,N_3993);
xor U4275 (N_4275,N_3618,N_3884);
nand U4276 (N_4276,N_3538,N_3653);
xnor U4277 (N_4277,N_3767,N_3566);
xnor U4278 (N_4278,N_3934,N_3916);
nand U4279 (N_4279,N_3510,N_3665);
nand U4280 (N_4280,N_3677,N_3732);
or U4281 (N_4281,N_3711,N_3963);
and U4282 (N_4282,N_3836,N_3758);
nand U4283 (N_4283,N_3634,N_3963);
and U4284 (N_4284,N_3515,N_3770);
nand U4285 (N_4285,N_3743,N_3883);
xnor U4286 (N_4286,N_3645,N_3557);
nor U4287 (N_4287,N_3634,N_3537);
and U4288 (N_4288,N_3828,N_3807);
nand U4289 (N_4289,N_3882,N_3718);
xor U4290 (N_4290,N_3919,N_3851);
nor U4291 (N_4291,N_3727,N_3670);
xnor U4292 (N_4292,N_3802,N_3758);
or U4293 (N_4293,N_3542,N_3566);
xor U4294 (N_4294,N_3671,N_3877);
and U4295 (N_4295,N_3657,N_3855);
or U4296 (N_4296,N_3625,N_3784);
and U4297 (N_4297,N_3596,N_3950);
nor U4298 (N_4298,N_3782,N_3934);
xor U4299 (N_4299,N_3978,N_3955);
xnor U4300 (N_4300,N_3516,N_3853);
or U4301 (N_4301,N_3651,N_3873);
and U4302 (N_4302,N_3735,N_3512);
and U4303 (N_4303,N_3706,N_3828);
xor U4304 (N_4304,N_3745,N_3800);
nand U4305 (N_4305,N_3649,N_3695);
nor U4306 (N_4306,N_3538,N_3605);
or U4307 (N_4307,N_3954,N_3929);
or U4308 (N_4308,N_3838,N_3947);
nand U4309 (N_4309,N_3990,N_3826);
nand U4310 (N_4310,N_3742,N_3845);
nand U4311 (N_4311,N_3770,N_3603);
and U4312 (N_4312,N_3504,N_3834);
nand U4313 (N_4313,N_3878,N_3535);
and U4314 (N_4314,N_3851,N_3820);
and U4315 (N_4315,N_3912,N_3743);
or U4316 (N_4316,N_3673,N_3969);
and U4317 (N_4317,N_3691,N_3716);
or U4318 (N_4318,N_3880,N_3555);
nor U4319 (N_4319,N_3758,N_3664);
xor U4320 (N_4320,N_3671,N_3954);
nand U4321 (N_4321,N_3727,N_3822);
or U4322 (N_4322,N_3686,N_3751);
nand U4323 (N_4323,N_3941,N_3774);
xor U4324 (N_4324,N_3800,N_3532);
nor U4325 (N_4325,N_3935,N_3761);
nor U4326 (N_4326,N_3644,N_3901);
xor U4327 (N_4327,N_3787,N_3514);
and U4328 (N_4328,N_3849,N_3733);
and U4329 (N_4329,N_3991,N_3807);
nor U4330 (N_4330,N_3961,N_3599);
nand U4331 (N_4331,N_3625,N_3725);
or U4332 (N_4332,N_3518,N_3672);
or U4333 (N_4333,N_3568,N_3928);
or U4334 (N_4334,N_3679,N_3579);
or U4335 (N_4335,N_3854,N_3908);
or U4336 (N_4336,N_3847,N_3791);
and U4337 (N_4337,N_3830,N_3933);
nand U4338 (N_4338,N_3817,N_3759);
nor U4339 (N_4339,N_3514,N_3544);
xnor U4340 (N_4340,N_3880,N_3754);
xnor U4341 (N_4341,N_3758,N_3791);
nand U4342 (N_4342,N_3559,N_3907);
nor U4343 (N_4343,N_3629,N_3753);
nor U4344 (N_4344,N_3745,N_3628);
xor U4345 (N_4345,N_3763,N_3803);
and U4346 (N_4346,N_3946,N_3713);
and U4347 (N_4347,N_3770,N_3702);
and U4348 (N_4348,N_3896,N_3815);
nand U4349 (N_4349,N_3740,N_3762);
xnor U4350 (N_4350,N_3739,N_3807);
or U4351 (N_4351,N_3731,N_3612);
xnor U4352 (N_4352,N_3928,N_3919);
nand U4353 (N_4353,N_3687,N_3716);
xor U4354 (N_4354,N_3553,N_3853);
nand U4355 (N_4355,N_3739,N_3532);
xor U4356 (N_4356,N_3596,N_3645);
or U4357 (N_4357,N_3874,N_3533);
xnor U4358 (N_4358,N_3660,N_3899);
and U4359 (N_4359,N_3531,N_3545);
nor U4360 (N_4360,N_3971,N_3775);
nor U4361 (N_4361,N_3820,N_3843);
xnor U4362 (N_4362,N_3816,N_3633);
nand U4363 (N_4363,N_3839,N_3932);
xor U4364 (N_4364,N_3656,N_3811);
xnor U4365 (N_4365,N_3537,N_3535);
nor U4366 (N_4366,N_3742,N_3558);
xnor U4367 (N_4367,N_3736,N_3880);
nand U4368 (N_4368,N_3676,N_3764);
or U4369 (N_4369,N_3662,N_3707);
nand U4370 (N_4370,N_3755,N_3996);
nand U4371 (N_4371,N_3750,N_3629);
xor U4372 (N_4372,N_3525,N_3858);
xnor U4373 (N_4373,N_3707,N_3783);
or U4374 (N_4374,N_3754,N_3572);
nor U4375 (N_4375,N_3890,N_3687);
nand U4376 (N_4376,N_3571,N_3729);
nor U4377 (N_4377,N_3865,N_3538);
nand U4378 (N_4378,N_3906,N_3603);
or U4379 (N_4379,N_3827,N_3941);
nand U4380 (N_4380,N_3695,N_3910);
nand U4381 (N_4381,N_3804,N_3661);
nor U4382 (N_4382,N_3893,N_3787);
nand U4383 (N_4383,N_3995,N_3937);
or U4384 (N_4384,N_3519,N_3583);
and U4385 (N_4385,N_3525,N_3947);
and U4386 (N_4386,N_3949,N_3843);
and U4387 (N_4387,N_3819,N_3814);
nor U4388 (N_4388,N_3510,N_3538);
nor U4389 (N_4389,N_3646,N_3654);
and U4390 (N_4390,N_3959,N_3869);
nand U4391 (N_4391,N_3868,N_3819);
nand U4392 (N_4392,N_3527,N_3575);
and U4393 (N_4393,N_3735,N_3623);
and U4394 (N_4394,N_3870,N_3698);
nor U4395 (N_4395,N_3843,N_3557);
xor U4396 (N_4396,N_3953,N_3713);
nor U4397 (N_4397,N_3654,N_3589);
nand U4398 (N_4398,N_3998,N_3714);
or U4399 (N_4399,N_3824,N_3595);
nand U4400 (N_4400,N_3900,N_3806);
nor U4401 (N_4401,N_3868,N_3552);
xnor U4402 (N_4402,N_3713,N_3532);
nand U4403 (N_4403,N_3647,N_3516);
xnor U4404 (N_4404,N_3657,N_3588);
xnor U4405 (N_4405,N_3718,N_3587);
nand U4406 (N_4406,N_3794,N_3935);
nand U4407 (N_4407,N_3924,N_3728);
or U4408 (N_4408,N_3966,N_3580);
and U4409 (N_4409,N_3747,N_3604);
nor U4410 (N_4410,N_3623,N_3796);
and U4411 (N_4411,N_3678,N_3946);
nand U4412 (N_4412,N_3854,N_3978);
or U4413 (N_4413,N_3839,N_3840);
or U4414 (N_4414,N_3533,N_3777);
nor U4415 (N_4415,N_3910,N_3975);
xor U4416 (N_4416,N_3788,N_3621);
xnor U4417 (N_4417,N_3798,N_3569);
nand U4418 (N_4418,N_3577,N_3708);
nor U4419 (N_4419,N_3962,N_3553);
or U4420 (N_4420,N_3590,N_3735);
and U4421 (N_4421,N_3763,N_3862);
nand U4422 (N_4422,N_3619,N_3807);
and U4423 (N_4423,N_3725,N_3963);
and U4424 (N_4424,N_3582,N_3764);
nand U4425 (N_4425,N_3715,N_3544);
or U4426 (N_4426,N_3683,N_3544);
nand U4427 (N_4427,N_3836,N_3518);
or U4428 (N_4428,N_3518,N_3538);
xor U4429 (N_4429,N_3599,N_3745);
nand U4430 (N_4430,N_3852,N_3913);
xor U4431 (N_4431,N_3833,N_3969);
or U4432 (N_4432,N_3950,N_3789);
nor U4433 (N_4433,N_3942,N_3967);
and U4434 (N_4434,N_3605,N_3548);
or U4435 (N_4435,N_3760,N_3931);
nand U4436 (N_4436,N_3596,N_3993);
nand U4437 (N_4437,N_3509,N_3584);
xor U4438 (N_4438,N_3533,N_3505);
nor U4439 (N_4439,N_3573,N_3652);
nand U4440 (N_4440,N_3544,N_3786);
and U4441 (N_4441,N_3570,N_3925);
and U4442 (N_4442,N_3777,N_3672);
and U4443 (N_4443,N_3845,N_3622);
xnor U4444 (N_4444,N_3676,N_3680);
and U4445 (N_4445,N_3700,N_3767);
or U4446 (N_4446,N_3835,N_3743);
or U4447 (N_4447,N_3508,N_3616);
xnor U4448 (N_4448,N_3890,N_3957);
xor U4449 (N_4449,N_3649,N_3612);
xnor U4450 (N_4450,N_3672,N_3854);
nor U4451 (N_4451,N_3854,N_3565);
xor U4452 (N_4452,N_3518,N_3831);
or U4453 (N_4453,N_3538,N_3579);
nand U4454 (N_4454,N_3962,N_3853);
nor U4455 (N_4455,N_3662,N_3741);
xor U4456 (N_4456,N_3635,N_3924);
nor U4457 (N_4457,N_3618,N_3640);
and U4458 (N_4458,N_3983,N_3713);
nor U4459 (N_4459,N_3665,N_3976);
xor U4460 (N_4460,N_3533,N_3634);
nand U4461 (N_4461,N_3706,N_3634);
and U4462 (N_4462,N_3648,N_3682);
xnor U4463 (N_4463,N_3814,N_3950);
nand U4464 (N_4464,N_3836,N_3963);
xor U4465 (N_4465,N_3992,N_3719);
and U4466 (N_4466,N_3944,N_3603);
or U4467 (N_4467,N_3727,N_3622);
and U4468 (N_4468,N_3852,N_3721);
and U4469 (N_4469,N_3874,N_3708);
or U4470 (N_4470,N_3827,N_3970);
xnor U4471 (N_4471,N_3763,N_3697);
nor U4472 (N_4472,N_3798,N_3848);
nor U4473 (N_4473,N_3684,N_3936);
nand U4474 (N_4474,N_3760,N_3516);
nand U4475 (N_4475,N_3656,N_3638);
or U4476 (N_4476,N_3888,N_3928);
xnor U4477 (N_4477,N_3797,N_3840);
or U4478 (N_4478,N_3778,N_3555);
xnor U4479 (N_4479,N_3905,N_3519);
xor U4480 (N_4480,N_3546,N_3869);
and U4481 (N_4481,N_3656,N_3889);
or U4482 (N_4482,N_3657,N_3629);
nor U4483 (N_4483,N_3835,N_3643);
and U4484 (N_4484,N_3548,N_3958);
nand U4485 (N_4485,N_3672,N_3667);
and U4486 (N_4486,N_3646,N_3518);
nor U4487 (N_4487,N_3508,N_3700);
xnor U4488 (N_4488,N_3944,N_3656);
nor U4489 (N_4489,N_3777,N_3522);
nor U4490 (N_4490,N_3788,N_3799);
nor U4491 (N_4491,N_3870,N_3933);
nand U4492 (N_4492,N_3877,N_3978);
and U4493 (N_4493,N_3662,N_3876);
xnor U4494 (N_4494,N_3634,N_3862);
or U4495 (N_4495,N_3564,N_3605);
or U4496 (N_4496,N_3627,N_3611);
xnor U4497 (N_4497,N_3625,N_3946);
nand U4498 (N_4498,N_3879,N_3790);
or U4499 (N_4499,N_3881,N_3567);
or U4500 (N_4500,N_4002,N_4271);
and U4501 (N_4501,N_4243,N_4313);
nor U4502 (N_4502,N_4136,N_4408);
or U4503 (N_4503,N_4450,N_4381);
nor U4504 (N_4504,N_4253,N_4194);
nor U4505 (N_4505,N_4227,N_4319);
or U4506 (N_4506,N_4224,N_4162);
and U4507 (N_4507,N_4076,N_4184);
nor U4508 (N_4508,N_4081,N_4422);
nand U4509 (N_4509,N_4466,N_4402);
nand U4510 (N_4510,N_4373,N_4218);
and U4511 (N_4511,N_4153,N_4142);
nor U4512 (N_4512,N_4292,N_4093);
nor U4513 (N_4513,N_4445,N_4475);
xor U4514 (N_4514,N_4395,N_4433);
or U4515 (N_4515,N_4219,N_4095);
xnor U4516 (N_4516,N_4298,N_4116);
xnor U4517 (N_4517,N_4028,N_4336);
nor U4518 (N_4518,N_4177,N_4178);
nor U4519 (N_4519,N_4353,N_4003);
nand U4520 (N_4520,N_4469,N_4242);
nand U4521 (N_4521,N_4311,N_4419);
xnor U4522 (N_4522,N_4409,N_4148);
and U4523 (N_4523,N_4122,N_4046);
and U4524 (N_4524,N_4111,N_4055);
nand U4525 (N_4525,N_4364,N_4155);
or U4526 (N_4526,N_4251,N_4334);
nor U4527 (N_4527,N_4151,N_4415);
nand U4528 (N_4528,N_4316,N_4064);
nand U4529 (N_4529,N_4405,N_4492);
or U4530 (N_4530,N_4039,N_4132);
or U4531 (N_4531,N_4392,N_4185);
xnor U4532 (N_4532,N_4288,N_4362);
and U4533 (N_4533,N_4261,N_4421);
nand U4534 (N_4534,N_4009,N_4416);
xor U4535 (N_4535,N_4145,N_4379);
nor U4536 (N_4536,N_4380,N_4443);
nand U4537 (N_4537,N_4426,N_4041);
xor U4538 (N_4538,N_4065,N_4449);
or U4539 (N_4539,N_4268,N_4239);
or U4540 (N_4540,N_4296,N_4036);
or U4541 (N_4541,N_4393,N_4324);
nand U4542 (N_4542,N_4286,N_4451);
nand U4543 (N_4543,N_4091,N_4150);
and U4544 (N_4544,N_4420,N_4190);
nand U4545 (N_4545,N_4322,N_4038);
and U4546 (N_4546,N_4453,N_4283);
nor U4547 (N_4547,N_4225,N_4376);
xor U4548 (N_4548,N_4167,N_4183);
or U4549 (N_4549,N_4103,N_4086);
nor U4550 (N_4550,N_4310,N_4391);
xor U4551 (N_4551,N_4198,N_4293);
xnor U4552 (N_4552,N_4377,N_4303);
nand U4553 (N_4553,N_4208,N_4099);
or U4554 (N_4554,N_4390,N_4120);
or U4555 (N_4555,N_4314,N_4211);
and U4556 (N_4556,N_4474,N_4318);
nor U4557 (N_4557,N_4105,N_4497);
nor U4558 (N_4558,N_4335,N_4329);
nor U4559 (N_4559,N_4372,N_4192);
nand U4560 (N_4560,N_4473,N_4438);
nor U4561 (N_4561,N_4189,N_4214);
and U4562 (N_4562,N_4212,N_4355);
and U4563 (N_4563,N_4435,N_4312);
or U4564 (N_4564,N_4258,N_4053);
and U4565 (N_4565,N_4174,N_4423);
xor U4566 (N_4566,N_4282,N_4035);
nand U4567 (N_4567,N_4315,N_4273);
or U4568 (N_4568,N_4398,N_4401);
xor U4569 (N_4569,N_4204,N_4487);
nand U4570 (N_4570,N_4112,N_4403);
or U4571 (N_4571,N_4436,N_4343);
and U4572 (N_4572,N_4179,N_4368);
nand U4573 (N_4573,N_4005,N_4220);
or U4574 (N_4574,N_4187,N_4340);
xor U4575 (N_4575,N_4356,N_4068);
xnor U4576 (N_4576,N_4460,N_4387);
nor U4577 (N_4577,N_4096,N_4094);
or U4578 (N_4578,N_4191,N_4452);
nor U4579 (N_4579,N_4305,N_4083);
nand U4580 (N_4580,N_4321,N_4197);
nor U4581 (N_4581,N_4146,N_4428);
nand U4582 (N_4582,N_4044,N_4418);
xor U4583 (N_4583,N_4207,N_4066);
xnor U4584 (N_4584,N_4172,N_4490);
xnor U4585 (N_4585,N_4455,N_4202);
xnor U4586 (N_4586,N_4470,N_4232);
nor U4587 (N_4587,N_4071,N_4245);
or U4588 (N_4588,N_4020,N_4131);
xor U4589 (N_4589,N_4431,N_4017);
or U4590 (N_4590,N_4217,N_4287);
or U4591 (N_4591,N_4240,N_4429);
or U4592 (N_4592,N_4238,N_4498);
or U4593 (N_4593,N_4259,N_4388);
nand U4594 (N_4594,N_4216,N_4168);
and U4595 (N_4595,N_4375,N_4047);
and U4596 (N_4596,N_4295,N_4163);
xor U4597 (N_4597,N_4366,N_4249);
nand U4598 (N_4598,N_4333,N_4165);
or U4599 (N_4599,N_4080,N_4430);
xnor U4600 (N_4600,N_4458,N_4459);
xor U4601 (N_4601,N_4326,N_4135);
nor U4602 (N_4602,N_4223,N_4203);
and U4603 (N_4603,N_4141,N_4247);
nor U4604 (N_4604,N_4444,N_4468);
xor U4605 (N_4605,N_4365,N_4457);
nor U4606 (N_4606,N_4033,N_4193);
and U4607 (N_4607,N_4357,N_4025);
nor U4608 (N_4608,N_4210,N_4482);
nand U4609 (N_4609,N_4317,N_4158);
nand U4610 (N_4610,N_4010,N_4118);
nand U4611 (N_4611,N_4186,N_4260);
and U4612 (N_4612,N_4462,N_4031);
and U4613 (N_4613,N_4327,N_4137);
nor U4614 (N_4614,N_4058,N_4359);
and U4615 (N_4615,N_4417,N_4256);
or U4616 (N_4616,N_4264,N_4048);
nor U4617 (N_4617,N_4117,N_4109);
and U4618 (N_4618,N_4289,N_4008);
xnor U4619 (N_4619,N_4266,N_4037);
xor U4620 (N_4620,N_4199,N_4342);
nor U4621 (N_4621,N_4016,N_4139);
xor U4622 (N_4622,N_4060,N_4156);
and U4623 (N_4623,N_4125,N_4015);
nand U4624 (N_4624,N_4309,N_4472);
nor U4625 (N_4625,N_4351,N_4078);
nor U4626 (N_4626,N_4115,N_4486);
or U4627 (N_4627,N_4241,N_4491);
or U4628 (N_4628,N_4488,N_4007);
or U4629 (N_4629,N_4425,N_4050);
and U4630 (N_4630,N_4481,N_4485);
nand U4631 (N_4631,N_4332,N_4045);
or U4632 (N_4632,N_4084,N_4348);
and U4633 (N_4633,N_4383,N_4069);
and U4634 (N_4634,N_4478,N_4265);
nor U4635 (N_4635,N_4371,N_4284);
nor U4636 (N_4636,N_4280,N_4344);
xnor U4637 (N_4637,N_4244,N_4275);
nor U4638 (N_4638,N_4171,N_4367);
xor U4639 (N_4639,N_4442,N_4213);
nor U4640 (N_4640,N_4014,N_4480);
or U4641 (N_4641,N_4072,N_4175);
nor U4642 (N_4642,N_4032,N_4206);
xnor U4643 (N_4643,N_4440,N_4149);
xnor U4644 (N_4644,N_4030,N_4108);
xnor U4645 (N_4645,N_4427,N_4496);
or U4646 (N_4646,N_4300,N_4128);
or U4647 (N_4647,N_4350,N_4325);
nor U4648 (N_4648,N_4098,N_4154);
or U4649 (N_4649,N_4101,N_4196);
and U4650 (N_4650,N_4307,N_4339);
nor U4651 (N_4651,N_4360,N_4346);
nor U4652 (N_4652,N_4308,N_4006);
and U4653 (N_4653,N_4042,N_4236);
or U4654 (N_4654,N_4411,N_4463);
nand U4655 (N_4655,N_4121,N_4018);
and U4656 (N_4656,N_4447,N_4089);
xnor U4657 (N_4657,N_4262,N_4205);
xnor U4658 (N_4658,N_4338,N_4056);
and U4659 (N_4659,N_4011,N_4267);
or U4660 (N_4660,N_4229,N_4161);
or U4661 (N_4661,N_4057,N_4147);
nor U4662 (N_4662,N_4277,N_4024);
and U4663 (N_4663,N_4022,N_4026);
nor U4664 (N_4664,N_4363,N_4144);
and U4665 (N_4665,N_4441,N_4230);
or U4666 (N_4666,N_4023,N_4345);
and U4667 (N_4667,N_4157,N_4233);
and U4668 (N_4668,N_4434,N_4181);
and U4669 (N_4669,N_4126,N_4323);
nor U4670 (N_4670,N_4404,N_4255);
nor U4671 (N_4671,N_4467,N_4097);
nand U4672 (N_4672,N_4087,N_4476);
nor U4673 (N_4673,N_4130,N_4274);
or U4674 (N_4674,N_4437,N_4133);
nor U4675 (N_4675,N_4297,N_4299);
or U4676 (N_4676,N_4234,N_4104);
xor U4677 (N_4677,N_4027,N_4140);
nor U4678 (N_4678,N_4389,N_4301);
and U4679 (N_4679,N_4396,N_4019);
nand U4680 (N_4680,N_4201,N_4079);
nand U4681 (N_4681,N_4034,N_4354);
nand U4682 (N_4682,N_4063,N_4013);
and U4683 (N_4683,N_4250,N_4159);
or U4684 (N_4684,N_4290,N_4209);
nor U4685 (N_4685,N_4123,N_4285);
and U4686 (N_4686,N_4100,N_4110);
nor U4687 (N_4687,N_4059,N_4143);
or U4688 (N_4688,N_4246,N_4374);
xnor U4689 (N_4689,N_4021,N_4235);
or U4690 (N_4690,N_4328,N_4067);
nand U4691 (N_4691,N_4370,N_4252);
or U4692 (N_4692,N_4341,N_4294);
nand U4693 (N_4693,N_4493,N_4477);
nor U4694 (N_4694,N_4465,N_4439);
or U4695 (N_4695,N_4051,N_4400);
or U4696 (N_4696,N_4062,N_4170);
nor U4697 (N_4697,N_4479,N_4291);
nor U4698 (N_4698,N_4306,N_4043);
nor U4699 (N_4699,N_4361,N_4129);
or U4700 (N_4700,N_4052,N_4231);
nand U4701 (N_4701,N_4082,N_4254);
nand U4702 (N_4702,N_4070,N_4413);
nor U4703 (N_4703,N_4378,N_4173);
or U4704 (N_4704,N_4138,N_4074);
or U4705 (N_4705,N_4088,N_4269);
and U4706 (N_4706,N_4085,N_4358);
nor U4707 (N_4707,N_4263,N_4215);
and U4708 (N_4708,N_4029,N_4407);
or U4709 (N_4709,N_4432,N_4397);
xor U4710 (N_4710,N_4221,N_4385);
and U4711 (N_4711,N_4134,N_4276);
nand U4712 (N_4712,N_4337,N_4279);
and U4713 (N_4713,N_4107,N_4499);
nor U4714 (N_4714,N_4483,N_4160);
and U4715 (N_4715,N_4237,N_4257);
nand U4716 (N_4716,N_4456,N_4406);
xor U4717 (N_4717,N_4272,N_4320);
nor U4718 (N_4718,N_4352,N_4330);
and U4719 (N_4719,N_4114,N_4448);
and U4720 (N_4720,N_4226,N_4195);
or U4721 (N_4721,N_4424,N_4494);
xor U4722 (N_4722,N_4061,N_4049);
or U4723 (N_4723,N_4169,N_4278);
nor U4724 (N_4724,N_4484,N_4248);
nor U4725 (N_4725,N_4075,N_4302);
xnor U4726 (N_4726,N_4012,N_4077);
nor U4727 (N_4727,N_4412,N_4410);
nand U4728 (N_4728,N_4106,N_4414);
xor U4729 (N_4729,N_4394,N_4040);
or U4730 (N_4730,N_4281,N_4166);
xor U4731 (N_4731,N_4495,N_4004);
and U4732 (N_4732,N_4127,N_4331);
nor U4733 (N_4733,N_4054,N_4188);
xor U4734 (N_4734,N_4347,N_4270);
and U4735 (N_4735,N_4119,N_4464);
or U4736 (N_4736,N_4000,N_4102);
and U4737 (N_4737,N_4349,N_4113);
or U4738 (N_4738,N_4152,N_4461);
and U4739 (N_4739,N_4124,N_4092);
xnor U4740 (N_4740,N_4369,N_4073);
nand U4741 (N_4741,N_4228,N_4454);
nand U4742 (N_4742,N_4446,N_4489);
nor U4743 (N_4743,N_4471,N_4399);
xor U4744 (N_4744,N_4180,N_4176);
or U4745 (N_4745,N_4001,N_4182);
and U4746 (N_4746,N_4222,N_4090);
nand U4747 (N_4747,N_4164,N_4200);
xor U4748 (N_4748,N_4384,N_4304);
and U4749 (N_4749,N_4382,N_4386);
nor U4750 (N_4750,N_4225,N_4475);
xor U4751 (N_4751,N_4099,N_4137);
nor U4752 (N_4752,N_4138,N_4422);
nor U4753 (N_4753,N_4425,N_4308);
nand U4754 (N_4754,N_4467,N_4450);
xor U4755 (N_4755,N_4220,N_4460);
xor U4756 (N_4756,N_4136,N_4089);
nand U4757 (N_4757,N_4458,N_4103);
and U4758 (N_4758,N_4448,N_4340);
nor U4759 (N_4759,N_4474,N_4388);
and U4760 (N_4760,N_4005,N_4440);
nor U4761 (N_4761,N_4112,N_4120);
and U4762 (N_4762,N_4167,N_4419);
nand U4763 (N_4763,N_4094,N_4028);
nand U4764 (N_4764,N_4310,N_4297);
nor U4765 (N_4765,N_4354,N_4041);
and U4766 (N_4766,N_4007,N_4081);
or U4767 (N_4767,N_4232,N_4072);
and U4768 (N_4768,N_4338,N_4095);
nand U4769 (N_4769,N_4352,N_4400);
or U4770 (N_4770,N_4006,N_4088);
or U4771 (N_4771,N_4437,N_4135);
xor U4772 (N_4772,N_4203,N_4499);
or U4773 (N_4773,N_4235,N_4249);
nand U4774 (N_4774,N_4432,N_4241);
and U4775 (N_4775,N_4356,N_4476);
and U4776 (N_4776,N_4239,N_4404);
or U4777 (N_4777,N_4038,N_4181);
or U4778 (N_4778,N_4297,N_4250);
xor U4779 (N_4779,N_4254,N_4196);
xnor U4780 (N_4780,N_4043,N_4247);
xor U4781 (N_4781,N_4418,N_4142);
xor U4782 (N_4782,N_4478,N_4284);
or U4783 (N_4783,N_4492,N_4218);
and U4784 (N_4784,N_4385,N_4177);
nand U4785 (N_4785,N_4362,N_4281);
and U4786 (N_4786,N_4458,N_4403);
and U4787 (N_4787,N_4257,N_4419);
nand U4788 (N_4788,N_4112,N_4080);
nor U4789 (N_4789,N_4371,N_4389);
or U4790 (N_4790,N_4004,N_4334);
and U4791 (N_4791,N_4186,N_4213);
nand U4792 (N_4792,N_4074,N_4481);
nor U4793 (N_4793,N_4484,N_4492);
xnor U4794 (N_4794,N_4019,N_4308);
xor U4795 (N_4795,N_4448,N_4208);
nand U4796 (N_4796,N_4225,N_4023);
or U4797 (N_4797,N_4089,N_4151);
nor U4798 (N_4798,N_4186,N_4226);
nand U4799 (N_4799,N_4394,N_4168);
nor U4800 (N_4800,N_4354,N_4158);
and U4801 (N_4801,N_4173,N_4470);
xor U4802 (N_4802,N_4394,N_4046);
xnor U4803 (N_4803,N_4017,N_4261);
nor U4804 (N_4804,N_4109,N_4248);
or U4805 (N_4805,N_4020,N_4280);
nor U4806 (N_4806,N_4167,N_4281);
or U4807 (N_4807,N_4353,N_4107);
xor U4808 (N_4808,N_4233,N_4439);
nand U4809 (N_4809,N_4135,N_4032);
xor U4810 (N_4810,N_4029,N_4046);
and U4811 (N_4811,N_4258,N_4143);
or U4812 (N_4812,N_4157,N_4301);
nand U4813 (N_4813,N_4101,N_4095);
and U4814 (N_4814,N_4042,N_4321);
nor U4815 (N_4815,N_4347,N_4492);
nor U4816 (N_4816,N_4333,N_4292);
nand U4817 (N_4817,N_4085,N_4181);
nand U4818 (N_4818,N_4260,N_4184);
and U4819 (N_4819,N_4330,N_4148);
nand U4820 (N_4820,N_4232,N_4331);
and U4821 (N_4821,N_4298,N_4037);
and U4822 (N_4822,N_4168,N_4103);
nor U4823 (N_4823,N_4476,N_4272);
nand U4824 (N_4824,N_4237,N_4132);
nor U4825 (N_4825,N_4277,N_4053);
nand U4826 (N_4826,N_4020,N_4302);
xor U4827 (N_4827,N_4200,N_4013);
and U4828 (N_4828,N_4224,N_4337);
xor U4829 (N_4829,N_4046,N_4188);
and U4830 (N_4830,N_4049,N_4439);
or U4831 (N_4831,N_4431,N_4254);
nand U4832 (N_4832,N_4057,N_4297);
and U4833 (N_4833,N_4251,N_4302);
nor U4834 (N_4834,N_4181,N_4243);
nor U4835 (N_4835,N_4218,N_4480);
nor U4836 (N_4836,N_4171,N_4349);
xnor U4837 (N_4837,N_4344,N_4364);
nand U4838 (N_4838,N_4093,N_4425);
and U4839 (N_4839,N_4196,N_4455);
nor U4840 (N_4840,N_4479,N_4029);
and U4841 (N_4841,N_4473,N_4143);
or U4842 (N_4842,N_4404,N_4048);
xor U4843 (N_4843,N_4187,N_4219);
or U4844 (N_4844,N_4317,N_4426);
or U4845 (N_4845,N_4370,N_4220);
or U4846 (N_4846,N_4124,N_4462);
and U4847 (N_4847,N_4166,N_4016);
xor U4848 (N_4848,N_4475,N_4281);
nand U4849 (N_4849,N_4218,N_4423);
and U4850 (N_4850,N_4344,N_4146);
or U4851 (N_4851,N_4400,N_4338);
xor U4852 (N_4852,N_4250,N_4141);
nor U4853 (N_4853,N_4491,N_4237);
nand U4854 (N_4854,N_4122,N_4238);
nor U4855 (N_4855,N_4384,N_4216);
xor U4856 (N_4856,N_4022,N_4418);
nor U4857 (N_4857,N_4340,N_4174);
nor U4858 (N_4858,N_4241,N_4457);
xnor U4859 (N_4859,N_4267,N_4051);
nor U4860 (N_4860,N_4222,N_4427);
and U4861 (N_4861,N_4203,N_4492);
nand U4862 (N_4862,N_4280,N_4389);
nand U4863 (N_4863,N_4172,N_4463);
xnor U4864 (N_4864,N_4428,N_4041);
and U4865 (N_4865,N_4040,N_4217);
nand U4866 (N_4866,N_4104,N_4198);
and U4867 (N_4867,N_4438,N_4011);
or U4868 (N_4868,N_4428,N_4163);
and U4869 (N_4869,N_4468,N_4240);
xor U4870 (N_4870,N_4365,N_4089);
nand U4871 (N_4871,N_4068,N_4346);
and U4872 (N_4872,N_4015,N_4390);
nand U4873 (N_4873,N_4206,N_4130);
xor U4874 (N_4874,N_4137,N_4215);
nor U4875 (N_4875,N_4484,N_4489);
nand U4876 (N_4876,N_4475,N_4451);
nand U4877 (N_4877,N_4432,N_4072);
nand U4878 (N_4878,N_4081,N_4360);
nand U4879 (N_4879,N_4219,N_4145);
and U4880 (N_4880,N_4176,N_4406);
or U4881 (N_4881,N_4161,N_4146);
nand U4882 (N_4882,N_4170,N_4362);
and U4883 (N_4883,N_4260,N_4116);
and U4884 (N_4884,N_4156,N_4140);
xnor U4885 (N_4885,N_4204,N_4394);
xor U4886 (N_4886,N_4233,N_4295);
xor U4887 (N_4887,N_4205,N_4475);
xor U4888 (N_4888,N_4073,N_4377);
or U4889 (N_4889,N_4085,N_4397);
or U4890 (N_4890,N_4119,N_4301);
and U4891 (N_4891,N_4404,N_4044);
nor U4892 (N_4892,N_4434,N_4210);
xor U4893 (N_4893,N_4372,N_4132);
nand U4894 (N_4894,N_4181,N_4314);
or U4895 (N_4895,N_4197,N_4139);
nand U4896 (N_4896,N_4155,N_4466);
nor U4897 (N_4897,N_4420,N_4021);
and U4898 (N_4898,N_4248,N_4399);
and U4899 (N_4899,N_4268,N_4164);
nor U4900 (N_4900,N_4090,N_4419);
or U4901 (N_4901,N_4178,N_4163);
or U4902 (N_4902,N_4491,N_4065);
and U4903 (N_4903,N_4400,N_4010);
xor U4904 (N_4904,N_4054,N_4313);
nor U4905 (N_4905,N_4198,N_4319);
and U4906 (N_4906,N_4012,N_4486);
nor U4907 (N_4907,N_4327,N_4008);
or U4908 (N_4908,N_4162,N_4159);
xnor U4909 (N_4909,N_4220,N_4381);
or U4910 (N_4910,N_4020,N_4413);
or U4911 (N_4911,N_4248,N_4498);
xor U4912 (N_4912,N_4296,N_4406);
nand U4913 (N_4913,N_4349,N_4418);
nor U4914 (N_4914,N_4320,N_4174);
or U4915 (N_4915,N_4084,N_4424);
xor U4916 (N_4916,N_4450,N_4246);
nand U4917 (N_4917,N_4346,N_4103);
nand U4918 (N_4918,N_4270,N_4455);
xor U4919 (N_4919,N_4151,N_4093);
nand U4920 (N_4920,N_4341,N_4087);
and U4921 (N_4921,N_4271,N_4048);
or U4922 (N_4922,N_4266,N_4419);
and U4923 (N_4923,N_4367,N_4229);
or U4924 (N_4924,N_4425,N_4268);
or U4925 (N_4925,N_4274,N_4049);
and U4926 (N_4926,N_4029,N_4307);
or U4927 (N_4927,N_4068,N_4396);
or U4928 (N_4928,N_4216,N_4022);
and U4929 (N_4929,N_4237,N_4445);
xnor U4930 (N_4930,N_4285,N_4114);
and U4931 (N_4931,N_4260,N_4339);
nor U4932 (N_4932,N_4456,N_4458);
and U4933 (N_4933,N_4219,N_4004);
nor U4934 (N_4934,N_4461,N_4391);
nand U4935 (N_4935,N_4024,N_4473);
xor U4936 (N_4936,N_4194,N_4215);
nand U4937 (N_4937,N_4308,N_4367);
nand U4938 (N_4938,N_4072,N_4091);
xor U4939 (N_4939,N_4155,N_4454);
or U4940 (N_4940,N_4025,N_4079);
nand U4941 (N_4941,N_4411,N_4067);
nand U4942 (N_4942,N_4145,N_4193);
nand U4943 (N_4943,N_4071,N_4214);
or U4944 (N_4944,N_4368,N_4424);
nand U4945 (N_4945,N_4233,N_4264);
or U4946 (N_4946,N_4439,N_4282);
nand U4947 (N_4947,N_4377,N_4029);
nor U4948 (N_4948,N_4165,N_4016);
xnor U4949 (N_4949,N_4186,N_4136);
nor U4950 (N_4950,N_4206,N_4489);
or U4951 (N_4951,N_4449,N_4292);
nand U4952 (N_4952,N_4094,N_4343);
or U4953 (N_4953,N_4470,N_4013);
and U4954 (N_4954,N_4481,N_4198);
xor U4955 (N_4955,N_4021,N_4166);
or U4956 (N_4956,N_4211,N_4137);
nor U4957 (N_4957,N_4182,N_4297);
or U4958 (N_4958,N_4437,N_4041);
xnor U4959 (N_4959,N_4376,N_4016);
nor U4960 (N_4960,N_4412,N_4082);
and U4961 (N_4961,N_4213,N_4495);
or U4962 (N_4962,N_4114,N_4060);
xor U4963 (N_4963,N_4475,N_4194);
nor U4964 (N_4964,N_4427,N_4050);
nor U4965 (N_4965,N_4426,N_4445);
nor U4966 (N_4966,N_4412,N_4070);
nor U4967 (N_4967,N_4490,N_4041);
or U4968 (N_4968,N_4246,N_4345);
nor U4969 (N_4969,N_4339,N_4372);
and U4970 (N_4970,N_4447,N_4058);
xnor U4971 (N_4971,N_4281,N_4390);
nand U4972 (N_4972,N_4064,N_4219);
nor U4973 (N_4973,N_4479,N_4412);
nand U4974 (N_4974,N_4080,N_4261);
nor U4975 (N_4975,N_4243,N_4341);
nor U4976 (N_4976,N_4274,N_4248);
and U4977 (N_4977,N_4081,N_4119);
or U4978 (N_4978,N_4338,N_4297);
and U4979 (N_4979,N_4401,N_4350);
and U4980 (N_4980,N_4437,N_4218);
xnor U4981 (N_4981,N_4448,N_4473);
or U4982 (N_4982,N_4232,N_4057);
nor U4983 (N_4983,N_4238,N_4378);
nor U4984 (N_4984,N_4380,N_4261);
and U4985 (N_4985,N_4272,N_4151);
nand U4986 (N_4986,N_4168,N_4386);
nand U4987 (N_4987,N_4295,N_4171);
nand U4988 (N_4988,N_4336,N_4457);
or U4989 (N_4989,N_4137,N_4360);
nor U4990 (N_4990,N_4228,N_4356);
and U4991 (N_4991,N_4403,N_4225);
nand U4992 (N_4992,N_4471,N_4146);
nor U4993 (N_4993,N_4167,N_4350);
nand U4994 (N_4994,N_4156,N_4080);
nand U4995 (N_4995,N_4083,N_4304);
xor U4996 (N_4996,N_4417,N_4476);
nand U4997 (N_4997,N_4383,N_4025);
nand U4998 (N_4998,N_4111,N_4452);
or U4999 (N_4999,N_4096,N_4097);
or U5000 (N_5000,N_4700,N_4882);
and U5001 (N_5001,N_4999,N_4802);
xor U5002 (N_5002,N_4838,N_4710);
or U5003 (N_5003,N_4753,N_4867);
nand U5004 (N_5004,N_4889,N_4827);
xor U5005 (N_5005,N_4797,N_4879);
nand U5006 (N_5006,N_4915,N_4973);
nor U5007 (N_5007,N_4637,N_4796);
or U5008 (N_5008,N_4703,N_4876);
nor U5009 (N_5009,N_4986,N_4606);
nor U5010 (N_5010,N_4854,N_4596);
or U5011 (N_5011,N_4800,N_4823);
and U5012 (N_5012,N_4971,N_4729);
nand U5013 (N_5013,N_4885,N_4545);
xnor U5014 (N_5014,N_4759,N_4899);
and U5015 (N_5015,N_4922,N_4506);
and U5016 (N_5016,N_4589,N_4904);
or U5017 (N_5017,N_4511,N_4745);
xor U5018 (N_5018,N_4592,N_4584);
and U5019 (N_5019,N_4547,N_4909);
xnor U5020 (N_5020,N_4788,N_4868);
or U5021 (N_5021,N_4508,N_4649);
nand U5022 (N_5022,N_4888,N_4910);
or U5023 (N_5023,N_4911,N_4805);
nand U5024 (N_5024,N_4801,N_4689);
nand U5025 (N_5025,N_4569,N_4956);
xnor U5026 (N_5026,N_4976,N_4990);
and U5027 (N_5027,N_4857,N_4526);
or U5028 (N_5028,N_4559,N_4556);
nand U5029 (N_5029,N_4713,N_4845);
xor U5030 (N_5030,N_4836,N_4578);
nor U5031 (N_5031,N_4648,N_4757);
and U5032 (N_5032,N_4894,N_4718);
or U5033 (N_5033,N_4624,N_4880);
xnor U5034 (N_5034,N_4977,N_4568);
and U5035 (N_5035,N_4622,N_4647);
nand U5036 (N_5036,N_4929,N_4519);
nor U5037 (N_5037,N_4708,N_4617);
nand U5038 (N_5038,N_4528,N_4505);
nand U5039 (N_5039,N_4810,N_4539);
nor U5040 (N_5040,N_4983,N_4724);
and U5041 (N_5041,N_4570,N_4590);
and U5042 (N_5042,N_4735,N_4982);
nor U5043 (N_5043,N_4787,N_4856);
or U5044 (N_5044,N_4962,N_4618);
xnor U5045 (N_5045,N_4761,N_4791);
and U5046 (N_5046,N_4935,N_4604);
or U5047 (N_5047,N_4641,N_4985);
xor U5048 (N_5048,N_4987,N_4830);
nand U5049 (N_5049,N_4679,N_4793);
nand U5050 (N_5050,N_4936,N_4813);
and U5051 (N_5051,N_4931,N_4835);
or U5052 (N_5052,N_4615,N_4642);
nor U5053 (N_5053,N_4549,N_4771);
or U5054 (N_5054,N_4979,N_4851);
nand U5055 (N_5055,N_4565,N_4881);
nor U5056 (N_5056,N_4825,N_4755);
or U5057 (N_5057,N_4864,N_4638);
nand U5058 (N_5058,N_4968,N_4597);
or U5059 (N_5059,N_4583,N_4668);
nand U5060 (N_5060,N_4947,N_4540);
nor U5061 (N_5061,N_4733,N_4917);
nor U5062 (N_5062,N_4548,N_4863);
or U5063 (N_5063,N_4581,N_4934);
xnor U5064 (N_5064,N_4869,N_4628);
xnor U5065 (N_5065,N_4953,N_4819);
nand U5066 (N_5066,N_4930,N_4727);
nor U5067 (N_5067,N_4636,N_4538);
and U5068 (N_5068,N_4646,N_4704);
nand U5069 (N_5069,N_4698,N_4705);
nor U5070 (N_5070,N_4969,N_4814);
nor U5071 (N_5071,N_4966,N_4503);
and U5072 (N_5072,N_4780,N_4643);
nand U5073 (N_5073,N_4877,N_4655);
nand U5074 (N_5074,N_4893,N_4776);
or U5075 (N_5075,N_4716,N_4551);
nand U5076 (N_5076,N_4507,N_4599);
or U5077 (N_5077,N_4984,N_4870);
nor U5078 (N_5078,N_4672,N_4840);
or U5079 (N_5079,N_4883,N_4758);
nand U5080 (N_5080,N_4842,N_4747);
xnor U5081 (N_5081,N_4919,N_4937);
xnor U5082 (N_5082,N_4886,N_4730);
nand U5083 (N_5083,N_4783,N_4573);
nor U5084 (N_5084,N_4946,N_4921);
and U5085 (N_5085,N_4812,N_4572);
nand U5086 (N_5086,N_4752,N_4964);
and U5087 (N_5087,N_4501,N_4785);
xor U5088 (N_5088,N_4737,N_4678);
nand U5089 (N_5089,N_4995,N_4792);
nor U5090 (N_5090,N_4804,N_4690);
xor U5091 (N_5091,N_4715,N_4920);
xor U5092 (N_5092,N_4858,N_4865);
nand U5093 (N_5093,N_4616,N_4900);
or U5094 (N_5094,N_4952,N_4558);
and U5095 (N_5095,N_4607,N_4586);
xor U5096 (N_5096,N_4587,N_4773);
and U5097 (N_5097,N_4996,N_4843);
or U5098 (N_5098,N_4872,N_4890);
nor U5099 (N_5099,N_4702,N_4520);
nand U5100 (N_5100,N_4645,N_4906);
nor U5101 (N_5101,N_4699,N_4714);
and U5102 (N_5102,N_4871,N_4631);
xnor U5103 (N_5103,N_4633,N_4512);
xor U5104 (N_5104,N_4666,N_4799);
and U5105 (N_5105,N_4701,N_4566);
and U5106 (N_5106,N_4510,N_4564);
and U5107 (N_5107,N_4772,N_4670);
and U5108 (N_5108,N_4938,N_4960);
nor U5109 (N_5109,N_4933,N_4907);
nor U5110 (N_5110,N_4691,N_4654);
xor U5111 (N_5111,N_4504,N_4866);
xor U5112 (N_5112,N_4914,N_4859);
nand U5113 (N_5113,N_4562,N_4826);
nand U5114 (N_5114,N_4707,N_4750);
or U5115 (N_5115,N_4774,N_4652);
xnor U5116 (N_5116,N_4958,N_4571);
and U5117 (N_5117,N_4903,N_4591);
xor U5118 (N_5118,N_4536,N_4623);
and U5119 (N_5119,N_4582,N_4898);
xnor U5120 (N_5120,N_4576,N_4656);
or U5121 (N_5121,N_4822,N_4594);
nand U5122 (N_5122,N_4719,N_4602);
and U5123 (N_5123,N_4908,N_4664);
nor U5124 (N_5124,N_4731,N_4709);
xnor U5125 (N_5125,N_4575,N_4782);
or U5126 (N_5126,N_4673,N_4809);
xor U5127 (N_5127,N_4789,N_4660);
xor U5128 (N_5128,N_4831,N_4820);
xor U5129 (N_5129,N_4878,N_4963);
nand U5130 (N_5130,N_4884,N_4683);
nand U5131 (N_5131,N_4850,N_4502);
xnor U5132 (N_5132,N_4777,N_4613);
nand U5133 (N_5133,N_4693,N_4741);
nor U5134 (N_5134,N_4650,N_4957);
xnor U5135 (N_5135,N_4897,N_4769);
and U5136 (N_5136,N_4967,N_4663);
xor U5137 (N_5137,N_4756,N_4852);
nor U5138 (N_5138,N_4529,N_4738);
or U5139 (N_5139,N_4754,N_4644);
or U5140 (N_5140,N_4561,N_4726);
nor U5141 (N_5141,N_4674,N_4524);
or U5142 (N_5142,N_4684,N_4912);
nor U5143 (N_5143,N_4994,N_4516);
nand U5144 (N_5144,N_4837,N_4530);
nand U5145 (N_5145,N_4535,N_4627);
xnor U5146 (N_5146,N_4546,N_4790);
or U5147 (N_5147,N_4686,N_4762);
xnor U5148 (N_5148,N_4665,N_4742);
xnor U5149 (N_5149,N_4766,N_4775);
xnor U5150 (N_5150,N_4577,N_4598);
and U5151 (N_5151,N_4661,N_4640);
and U5152 (N_5152,N_4696,N_4860);
nand U5153 (N_5153,N_4926,N_4816);
xor U5154 (N_5154,N_4717,N_4891);
and U5155 (N_5155,N_4605,N_4728);
nand U5156 (N_5156,N_4841,N_4625);
xor U5157 (N_5157,N_4736,N_4676);
and U5158 (N_5158,N_4657,N_4658);
or U5159 (N_5159,N_4853,N_4629);
or U5160 (N_5160,N_4687,N_4961);
and U5161 (N_5161,N_4849,N_4828);
xor U5162 (N_5162,N_4531,N_4744);
nand U5163 (N_5163,N_4610,N_4944);
or U5164 (N_5164,N_4579,N_4550);
xor U5165 (N_5165,N_4950,N_4651);
xnor U5166 (N_5166,N_4720,N_4895);
or U5167 (N_5167,N_4552,N_4974);
or U5168 (N_5168,N_4740,N_4778);
nand U5169 (N_5169,N_4611,N_4659);
nand U5170 (N_5170,N_4913,N_4544);
and U5171 (N_5171,N_4989,N_4517);
or U5172 (N_5172,N_4669,N_4749);
or U5173 (N_5173,N_4940,N_4580);
or U5174 (N_5174,N_4833,N_4692);
or U5175 (N_5175,N_4553,N_4887);
and U5176 (N_5176,N_4991,N_4721);
nor U5177 (N_5177,N_4513,N_4824);
nor U5178 (N_5178,N_4939,N_4518);
and U5179 (N_5179,N_4815,N_4560);
and U5180 (N_5180,N_4639,N_4975);
nor U5181 (N_5181,N_4525,N_4734);
nor U5182 (N_5182,N_4998,N_4839);
nor U5183 (N_5183,N_4896,N_4786);
nand U5184 (N_5184,N_4563,N_4765);
nand U5185 (N_5185,N_4806,N_4509);
or U5186 (N_5186,N_4965,N_4732);
and U5187 (N_5187,N_4993,N_4588);
nand U5188 (N_5188,N_4981,N_4954);
and U5189 (N_5189,N_4794,N_4601);
and U5190 (N_5190,N_4927,N_4768);
and U5191 (N_5191,N_4861,N_4847);
nor U5192 (N_5192,N_4523,N_4600);
nor U5193 (N_5193,N_4542,N_4992);
xnor U5194 (N_5194,N_4630,N_4534);
and U5195 (N_5195,N_4557,N_4862);
nor U5196 (N_5196,N_4697,N_4751);
nand U5197 (N_5197,N_4807,N_4817);
nand U5198 (N_5198,N_4892,N_4667);
nor U5199 (N_5199,N_4725,N_4902);
nor U5200 (N_5200,N_4739,N_4500);
xnor U5201 (N_5201,N_4923,N_4695);
nor U5202 (N_5202,N_4541,N_4634);
or U5203 (N_5203,N_4988,N_4608);
xnor U5204 (N_5204,N_4593,N_4671);
xor U5205 (N_5205,N_4875,N_4711);
nor U5206 (N_5206,N_4978,N_4743);
xnor U5207 (N_5207,N_4945,N_4626);
or U5208 (N_5208,N_4653,N_4533);
and U5209 (N_5209,N_4972,N_4585);
or U5210 (N_5210,N_4970,N_4924);
or U5211 (N_5211,N_4574,N_4941);
nand U5212 (N_5212,N_4619,N_4808);
and U5213 (N_5213,N_4722,N_4948);
nor U5214 (N_5214,N_4677,N_4829);
or U5215 (N_5215,N_4521,N_4763);
and U5216 (N_5216,N_4942,N_4621);
nor U5217 (N_5217,N_4918,N_4925);
nand U5218 (N_5218,N_4818,N_4834);
nor U5219 (N_5219,N_4955,N_4770);
xor U5220 (N_5220,N_4905,N_4848);
or U5221 (N_5221,N_4675,N_4980);
nand U5222 (N_5222,N_4688,N_4784);
or U5223 (N_5223,N_4959,N_4662);
nor U5224 (N_5224,N_4712,N_4832);
nor U5225 (N_5225,N_4928,N_4767);
or U5226 (N_5226,N_4803,N_4949);
and U5227 (N_5227,N_4694,N_4603);
and U5228 (N_5228,N_4681,N_4873);
nand U5229 (N_5229,N_4522,N_4620);
nor U5230 (N_5230,N_4567,N_4682);
nor U5231 (N_5231,N_4685,N_4795);
nand U5232 (N_5232,N_4532,N_4781);
and U5233 (N_5233,N_4943,N_4764);
nand U5234 (N_5234,N_4746,N_4614);
nand U5235 (N_5235,N_4997,N_4932);
and U5236 (N_5236,N_4901,N_4537);
or U5237 (N_5237,N_4609,N_4515);
or U5238 (N_5238,N_4543,N_4723);
nor U5239 (N_5239,N_4811,N_4612);
and U5240 (N_5240,N_4748,N_4760);
xnor U5241 (N_5241,N_4779,N_4555);
nor U5242 (N_5242,N_4846,N_4855);
nor U5243 (N_5243,N_4632,N_4635);
xnor U5244 (N_5244,N_4951,N_4844);
nand U5245 (N_5245,N_4554,N_4680);
nor U5246 (N_5246,N_4798,N_4821);
xor U5247 (N_5247,N_4706,N_4514);
nor U5248 (N_5248,N_4527,N_4916);
nor U5249 (N_5249,N_4595,N_4874);
nor U5250 (N_5250,N_4895,N_4746);
nand U5251 (N_5251,N_4843,N_4610);
or U5252 (N_5252,N_4949,N_4990);
or U5253 (N_5253,N_4703,N_4670);
xor U5254 (N_5254,N_4662,N_4705);
xor U5255 (N_5255,N_4747,N_4762);
nand U5256 (N_5256,N_4513,N_4911);
and U5257 (N_5257,N_4823,N_4992);
and U5258 (N_5258,N_4937,N_4662);
xor U5259 (N_5259,N_4642,N_4692);
nand U5260 (N_5260,N_4529,N_4538);
nor U5261 (N_5261,N_4945,N_4813);
and U5262 (N_5262,N_4532,N_4576);
or U5263 (N_5263,N_4607,N_4954);
nand U5264 (N_5264,N_4801,N_4503);
nand U5265 (N_5265,N_4886,N_4833);
nor U5266 (N_5266,N_4584,N_4808);
nand U5267 (N_5267,N_4599,N_4683);
nor U5268 (N_5268,N_4728,N_4949);
or U5269 (N_5269,N_4841,N_4557);
nor U5270 (N_5270,N_4836,N_4642);
nor U5271 (N_5271,N_4931,N_4691);
nor U5272 (N_5272,N_4662,N_4801);
and U5273 (N_5273,N_4761,N_4641);
or U5274 (N_5274,N_4983,N_4936);
and U5275 (N_5275,N_4532,N_4605);
or U5276 (N_5276,N_4978,N_4562);
nor U5277 (N_5277,N_4616,N_4680);
or U5278 (N_5278,N_4911,N_4752);
and U5279 (N_5279,N_4935,N_4907);
nand U5280 (N_5280,N_4785,N_4695);
or U5281 (N_5281,N_4971,N_4941);
nor U5282 (N_5282,N_4561,N_4924);
or U5283 (N_5283,N_4572,N_4600);
nor U5284 (N_5284,N_4736,N_4818);
or U5285 (N_5285,N_4750,N_4757);
or U5286 (N_5286,N_4666,N_4787);
or U5287 (N_5287,N_4606,N_4824);
and U5288 (N_5288,N_4700,N_4840);
xnor U5289 (N_5289,N_4898,N_4542);
nand U5290 (N_5290,N_4645,N_4747);
or U5291 (N_5291,N_4631,N_4984);
and U5292 (N_5292,N_4734,N_4533);
nor U5293 (N_5293,N_4893,N_4637);
and U5294 (N_5294,N_4834,N_4757);
nor U5295 (N_5295,N_4607,N_4890);
nand U5296 (N_5296,N_4867,N_4831);
and U5297 (N_5297,N_4656,N_4685);
or U5298 (N_5298,N_4563,N_4725);
nor U5299 (N_5299,N_4862,N_4589);
xor U5300 (N_5300,N_4580,N_4505);
nor U5301 (N_5301,N_4509,N_4501);
nand U5302 (N_5302,N_4604,N_4934);
xnor U5303 (N_5303,N_4969,N_4753);
and U5304 (N_5304,N_4954,N_4980);
nand U5305 (N_5305,N_4880,N_4732);
nor U5306 (N_5306,N_4747,N_4992);
or U5307 (N_5307,N_4817,N_4686);
or U5308 (N_5308,N_4940,N_4539);
xor U5309 (N_5309,N_4689,N_4569);
xnor U5310 (N_5310,N_4524,N_4558);
nand U5311 (N_5311,N_4994,N_4815);
nand U5312 (N_5312,N_4939,N_4628);
and U5313 (N_5313,N_4816,N_4801);
nor U5314 (N_5314,N_4600,N_4566);
or U5315 (N_5315,N_4693,N_4914);
or U5316 (N_5316,N_4593,N_4860);
xnor U5317 (N_5317,N_4511,N_4613);
or U5318 (N_5318,N_4534,N_4516);
nand U5319 (N_5319,N_4549,N_4768);
or U5320 (N_5320,N_4741,N_4665);
and U5321 (N_5321,N_4894,N_4857);
xnor U5322 (N_5322,N_4954,N_4973);
nand U5323 (N_5323,N_4816,N_4711);
nand U5324 (N_5324,N_4716,N_4791);
nor U5325 (N_5325,N_4788,N_4753);
and U5326 (N_5326,N_4598,N_4863);
or U5327 (N_5327,N_4684,N_4730);
nand U5328 (N_5328,N_4510,N_4897);
or U5329 (N_5329,N_4955,N_4894);
nand U5330 (N_5330,N_4779,N_4879);
nand U5331 (N_5331,N_4898,N_4900);
nor U5332 (N_5332,N_4522,N_4664);
or U5333 (N_5333,N_4504,N_4974);
or U5334 (N_5334,N_4859,N_4831);
nand U5335 (N_5335,N_4569,N_4809);
and U5336 (N_5336,N_4934,N_4720);
nand U5337 (N_5337,N_4726,N_4662);
nor U5338 (N_5338,N_4746,N_4695);
nor U5339 (N_5339,N_4669,N_4883);
nand U5340 (N_5340,N_4827,N_4513);
nor U5341 (N_5341,N_4575,N_4700);
nand U5342 (N_5342,N_4852,N_4613);
xnor U5343 (N_5343,N_4549,N_4816);
nand U5344 (N_5344,N_4710,N_4955);
nand U5345 (N_5345,N_4945,N_4867);
nand U5346 (N_5346,N_4808,N_4972);
nand U5347 (N_5347,N_4754,N_4668);
xnor U5348 (N_5348,N_4959,N_4806);
nor U5349 (N_5349,N_4624,N_4668);
nor U5350 (N_5350,N_4718,N_4553);
or U5351 (N_5351,N_4830,N_4667);
nand U5352 (N_5352,N_4926,N_4990);
or U5353 (N_5353,N_4984,N_4832);
xor U5354 (N_5354,N_4589,N_4541);
or U5355 (N_5355,N_4718,N_4575);
or U5356 (N_5356,N_4988,N_4698);
nand U5357 (N_5357,N_4913,N_4723);
nand U5358 (N_5358,N_4838,N_4939);
nand U5359 (N_5359,N_4597,N_4993);
nor U5360 (N_5360,N_4662,N_4905);
xnor U5361 (N_5361,N_4978,N_4928);
nor U5362 (N_5362,N_4834,N_4549);
nor U5363 (N_5363,N_4770,N_4771);
nand U5364 (N_5364,N_4927,N_4697);
xor U5365 (N_5365,N_4548,N_4502);
nand U5366 (N_5366,N_4976,N_4766);
xor U5367 (N_5367,N_4615,N_4881);
or U5368 (N_5368,N_4960,N_4735);
nand U5369 (N_5369,N_4694,N_4572);
nand U5370 (N_5370,N_4693,N_4947);
xnor U5371 (N_5371,N_4863,N_4728);
or U5372 (N_5372,N_4801,N_4532);
nor U5373 (N_5373,N_4849,N_4567);
or U5374 (N_5374,N_4646,N_4635);
nand U5375 (N_5375,N_4956,N_4996);
nand U5376 (N_5376,N_4505,N_4502);
xnor U5377 (N_5377,N_4994,N_4798);
nand U5378 (N_5378,N_4534,N_4775);
nor U5379 (N_5379,N_4575,N_4539);
nor U5380 (N_5380,N_4573,N_4526);
nand U5381 (N_5381,N_4694,N_4766);
nand U5382 (N_5382,N_4621,N_4654);
and U5383 (N_5383,N_4978,N_4932);
and U5384 (N_5384,N_4567,N_4596);
nor U5385 (N_5385,N_4803,N_4805);
or U5386 (N_5386,N_4517,N_4556);
or U5387 (N_5387,N_4871,N_4832);
xnor U5388 (N_5388,N_4709,N_4792);
and U5389 (N_5389,N_4990,N_4968);
or U5390 (N_5390,N_4950,N_4648);
xor U5391 (N_5391,N_4904,N_4794);
nand U5392 (N_5392,N_4705,N_4771);
and U5393 (N_5393,N_4551,N_4585);
or U5394 (N_5394,N_4684,N_4872);
xor U5395 (N_5395,N_4917,N_4591);
and U5396 (N_5396,N_4774,N_4839);
nor U5397 (N_5397,N_4724,N_4897);
or U5398 (N_5398,N_4560,N_4524);
nand U5399 (N_5399,N_4584,N_4654);
xnor U5400 (N_5400,N_4613,N_4505);
nor U5401 (N_5401,N_4871,N_4736);
nand U5402 (N_5402,N_4980,N_4521);
nor U5403 (N_5403,N_4629,N_4778);
nand U5404 (N_5404,N_4618,N_4926);
and U5405 (N_5405,N_4834,N_4795);
xor U5406 (N_5406,N_4767,N_4821);
xnor U5407 (N_5407,N_4977,N_4748);
nand U5408 (N_5408,N_4772,N_4633);
nand U5409 (N_5409,N_4534,N_4784);
nand U5410 (N_5410,N_4892,N_4698);
and U5411 (N_5411,N_4568,N_4849);
xnor U5412 (N_5412,N_4799,N_4865);
nand U5413 (N_5413,N_4905,N_4619);
or U5414 (N_5414,N_4846,N_4539);
or U5415 (N_5415,N_4837,N_4656);
and U5416 (N_5416,N_4976,N_4724);
and U5417 (N_5417,N_4603,N_4609);
nor U5418 (N_5418,N_4583,N_4717);
nand U5419 (N_5419,N_4718,N_4753);
nand U5420 (N_5420,N_4922,N_4540);
xnor U5421 (N_5421,N_4537,N_4714);
nand U5422 (N_5422,N_4864,N_4521);
nand U5423 (N_5423,N_4518,N_4686);
nor U5424 (N_5424,N_4709,N_4956);
and U5425 (N_5425,N_4950,N_4760);
nor U5426 (N_5426,N_4747,N_4812);
or U5427 (N_5427,N_4800,N_4853);
nand U5428 (N_5428,N_4609,N_4528);
or U5429 (N_5429,N_4896,N_4966);
or U5430 (N_5430,N_4708,N_4522);
and U5431 (N_5431,N_4889,N_4909);
xor U5432 (N_5432,N_4589,N_4544);
xnor U5433 (N_5433,N_4678,N_4511);
nor U5434 (N_5434,N_4663,N_4821);
and U5435 (N_5435,N_4893,N_4922);
nand U5436 (N_5436,N_4882,N_4824);
xnor U5437 (N_5437,N_4676,N_4822);
nand U5438 (N_5438,N_4505,N_4787);
nand U5439 (N_5439,N_4931,N_4941);
or U5440 (N_5440,N_4575,N_4511);
and U5441 (N_5441,N_4564,N_4899);
nor U5442 (N_5442,N_4600,N_4796);
or U5443 (N_5443,N_4512,N_4926);
nand U5444 (N_5444,N_4863,N_4788);
nor U5445 (N_5445,N_4548,N_4736);
xor U5446 (N_5446,N_4797,N_4929);
nand U5447 (N_5447,N_4745,N_4670);
or U5448 (N_5448,N_4742,N_4934);
or U5449 (N_5449,N_4949,N_4593);
or U5450 (N_5450,N_4725,N_4691);
or U5451 (N_5451,N_4806,N_4565);
and U5452 (N_5452,N_4964,N_4791);
and U5453 (N_5453,N_4622,N_4950);
xor U5454 (N_5454,N_4579,N_4540);
and U5455 (N_5455,N_4508,N_4868);
nor U5456 (N_5456,N_4784,N_4553);
nand U5457 (N_5457,N_4790,N_4899);
nor U5458 (N_5458,N_4848,N_4913);
xnor U5459 (N_5459,N_4508,N_4686);
nor U5460 (N_5460,N_4653,N_4775);
or U5461 (N_5461,N_4571,N_4624);
or U5462 (N_5462,N_4913,N_4875);
xnor U5463 (N_5463,N_4848,N_4583);
xnor U5464 (N_5464,N_4644,N_4989);
and U5465 (N_5465,N_4623,N_4692);
nor U5466 (N_5466,N_4830,N_4802);
nor U5467 (N_5467,N_4598,N_4997);
and U5468 (N_5468,N_4954,N_4795);
or U5469 (N_5469,N_4843,N_4511);
and U5470 (N_5470,N_4889,N_4516);
xor U5471 (N_5471,N_4836,N_4933);
xor U5472 (N_5472,N_4997,N_4635);
nand U5473 (N_5473,N_4565,N_4696);
xnor U5474 (N_5474,N_4705,N_4857);
or U5475 (N_5475,N_4932,N_4603);
and U5476 (N_5476,N_4966,N_4849);
nor U5477 (N_5477,N_4945,N_4589);
nand U5478 (N_5478,N_4714,N_4973);
nand U5479 (N_5479,N_4748,N_4682);
nor U5480 (N_5480,N_4510,N_4644);
and U5481 (N_5481,N_4741,N_4938);
or U5482 (N_5482,N_4704,N_4936);
or U5483 (N_5483,N_4608,N_4977);
and U5484 (N_5484,N_4585,N_4986);
nor U5485 (N_5485,N_4725,N_4724);
and U5486 (N_5486,N_4685,N_4868);
xor U5487 (N_5487,N_4541,N_4854);
xnor U5488 (N_5488,N_4561,N_4553);
nor U5489 (N_5489,N_4894,N_4699);
xnor U5490 (N_5490,N_4585,N_4859);
and U5491 (N_5491,N_4895,N_4676);
nor U5492 (N_5492,N_4805,N_4534);
nor U5493 (N_5493,N_4650,N_4967);
xnor U5494 (N_5494,N_4603,N_4987);
and U5495 (N_5495,N_4742,N_4913);
and U5496 (N_5496,N_4765,N_4759);
xor U5497 (N_5497,N_4519,N_4868);
and U5498 (N_5498,N_4982,N_4839);
or U5499 (N_5499,N_4848,N_4566);
nor U5500 (N_5500,N_5092,N_5440);
xor U5501 (N_5501,N_5168,N_5485);
or U5502 (N_5502,N_5378,N_5363);
nor U5503 (N_5503,N_5045,N_5468);
and U5504 (N_5504,N_5303,N_5035);
xor U5505 (N_5505,N_5419,N_5191);
nand U5506 (N_5506,N_5308,N_5342);
xor U5507 (N_5507,N_5403,N_5186);
nand U5508 (N_5508,N_5269,N_5421);
and U5509 (N_5509,N_5277,N_5345);
and U5510 (N_5510,N_5249,N_5404);
xnor U5511 (N_5511,N_5085,N_5260);
xnor U5512 (N_5512,N_5270,N_5413);
nand U5513 (N_5513,N_5040,N_5450);
nand U5514 (N_5514,N_5401,N_5020);
nor U5515 (N_5515,N_5391,N_5087);
or U5516 (N_5516,N_5012,N_5102);
nand U5517 (N_5517,N_5252,N_5321);
xnor U5518 (N_5518,N_5365,N_5228);
and U5519 (N_5519,N_5212,N_5390);
nor U5520 (N_5520,N_5197,N_5209);
nor U5521 (N_5521,N_5352,N_5013);
nor U5522 (N_5522,N_5354,N_5145);
xnor U5523 (N_5523,N_5036,N_5077);
or U5524 (N_5524,N_5106,N_5198);
xor U5525 (N_5525,N_5499,N_5446);
nor U5526 (N_5526,N_5187,N_5067);
xnor U5527 (N_5527,N_5193,N_5332);
and U5528 (N_5528,N_5152,N_5215);
or U5529 (N_5529,N_5165,N_5283);
xnor U5530 (N_5530,N_5163,N_5090);
nor U5531 (N_5531,N_5483,N_5177);
nand U5532 (N_5532,N_5052,N_5002);
or U5533 (N_5533,N_5431,N_5096);
and U5534 (N_5534,N_5107,N_5079);
xnor U5535 (N_5535,N_5100,N_5451);
and U5536 (N_5536,N_5465,N_5392);
and U5537 (N_5537,N_5007,N_5267);
nand U5538 (N_5538,N_5299,N_5147);
or U5539 (N_5539,N_5072,N_5495);
nand U5540 (N_5540,N_5005,N_5449);
or U5541 (N_5541,N_5098,N_5211);
nor U5542 (N_5542,N_5222,N_5441);
and U5543 (N_5543,N_5349,N_5265);
and U5544 (N_5544,N_5157,N_5080);
nor U5545 (N_5545,N_5289,N_5395);
nand U5546 (N_5546,N_5280,N_5353);
nor U5547 (N_5547,N_5261,N_5083);
xnor U5548 (N_5548,N_5455,N_5396);
and U5549 (N_5549,N_5358,N_5425);
or U5550 (N_5550,N_5438,N_5161);
nand U5551 (N_5551,N_5134,N_5302);
nor U5552 (N_5552,N_5316,N_5082);
nor U5553 (N_5553,N_5307,N_5015);
nand U5554 (N_5554,N_5498,N_5330);
nor U5555 (N_5555,N_5482,N_5114);
xor U5556 (N_5556,N_5324,N_5304);
or U5557 (N_5557,N_5070,N_5429);
xor U5558 (N_5558,N_5164,N_5377);
nor U5559 (N_5559,N_5169,N_5227);
nor U5560 (N_5560,N_5028,N_5056);
xor U5561 (N_5561,N_5050,N_5296);
or U5562 (N_5562,N_5472,N_5051);
and U5563 (N_5563,N_5207,N_5481);
and U5564 (N_5564,N_5104,N_5266);
and U5565 (N_5565,N_5009,N_5117);
and U5566 (N_5566,N_5412,N_5210);
nand U5567 (N_5567,N_5016,N_5146);
nand U5568 (N_5568,N_5244,N_5325);
or U5569 (N_5569,N_5124,N_5359);
and U5570 (N_5570,N_5469,N_5194);
xnor U5571 (N_5571,N_5411,N_5370);
xnor U5572 (N_5572,N_5199,N_5356);
xnor U5573 (N_5573,N_5291,N_5360);
nand U5574 (N_5574,N_5043,N_5433);
and U5575 (N_5575,N_5427,N_5057);
xor U5576 (N_5576,N_5301,N_5258);
nand U5577 (N_5577,N_5017,N_5357);
or U5578 (N_5578,N_5306,N_5093);
nor U5579 (N_5579,N_5122,N_5158);
nand U5580 (N_5580,N_5263,N_5133);
or U5581 (N_5581,N_5150,N_5381);
and U5582 (N_5582,N_5407,N_5179);
xnor U5583 (N_5583,N_5091,N_5064);
nand U5584 (N_5584,N_5128,N_5167);
nand U5585 (N_5585,N_5213,N_5275);
xor U5586 (N_5586,N_5251,N_5497);
nor U5587 (N_5587,N_5366,N_5166);
or U5588 (N_5588,N_5019,N_5350);
or U5589 (N_5589,N_5333,N_5162);
nor U5590 (N_5590,N_5334,N_5273);
nor U5591 (N_5591,N_5470,N_5143);
nand U5592 (N_5592,N_5063,N_5241);
xor U5593 (N_5593,N_5111,N_5027);
or U5594 (N_5594,N_5118,N_5250);
xnor U5595 (N_5595,N_5402,N_5417);
nor U5596 (N_5596,N_5119,N_5081);
xor U5597 (N_5597,N_5322,N_5214);
or U5598 (N_5598,N_5101,N_5320);
xor U5599 (N_5599,N_5371,N_5400);
nor U5600 (N_5600,N_5201,N_5113);
nand U5601 (N_5601,N_5397,N_5340);
xnor U5602 (N_5602,N_5039,N_5327);
xnor U5603 (N_5603,N_5399,N_5439);
and U5604 (N_5604,N_5243,N_5484);
xnor U5605 (N_5605,N_5406,N_5149);
xnor U5606 (N_5606,N_5038,N_5226);
nand U5607 (N_5607,N_5463,N_5132);
and U5608 (N_5608,N_5315,N_5493);
nand U5609 (N_5609,N_5135,N_5492);
and U5610 (N_5610,N_5346,N_5264);
xnor U5611 (N_5611,N_5021,N_5123);
nand U5612 (N_5612,N_5206,N_5058);
nor U5613 (N_5613,N_5000,N_5130);
and U5614 (N_5614,N_5443,N_5127);
xor U5615 (N_5615,N_5178,N_5294);
xor U5616 (N_5616,N_5071,N_5225);
and U5617 (N_5617,N_5240,N_5276);
or U5618 (N_5618,N_5285,N_5192);
xnor U5619 (N_5619,N_5182,N_5245);
and U5620 (N_5620,N_5231,N_5023);
nor U5621 (N_5621,N_5125,N_5311);
nand U5622 (N_5622,N_5060,N_5305);
xor U5623 (N_5623,N_5108,N_5183);
nand U5624 (N_5624,N_5233,N_5151);
or U5625 (N_5625,N_5076,N_5061);
nor U5626 (N_5626,N_5338,N_5208);
and U5627 (N_5627,N_5084,N_5385);
and U5628 (N_5628,N_5105,N_5398);
nor U5629 (N_5629,N_5202,N_5310);
xor U5630 (N_5630,N_5328,N_5094);
or U5631 (N_5631,N_5144,N_5042);
or U5632 (N_5632,N_5180,N_5435);
nand U5633 (N_5633,N_5314,N_5116);
and U5634 (N_5634,N_5355,N_5216);
or U5635 (N_5635,N_5424,N_5386);
or U5636 (N_5636,N_5099,N_5459);
and U5637 (N_5637,N_5029,N_5297);
nor U5638 (N_5638,N_5078,N_5480);
nor U5639 (N_5639,N_5159,N_5437);
and U5640 (N_5640,N_5255,N_5362);
nand U5641 (N_5641,N_5382,N_5171);
nand U5642 (N_5642,N_5282,N_5287);
nand U5643 (N_5643,N_5474,N_5298);
xnor U5644 (N_5644,N_5136,N_5293);
and U5645 (N_5645,N_5220,N_5218);
xnor U5646 (N_5646,N_5479,N_5008);
xor U5647 (N_5647,N_5237,N_5138);
and U5648 (N_5648,N_5317,N_5010);
or U5649 (N_5649,N_5488,N_5312);
nor U5650 (N_5650,N_5313,N_5453);
or U5651 (N_5651,N_5066,N_5248);
and U5652 (N_5652,N_5466,N_5054);
nor U5653 (N_5653,N_5257,N_5430);
nand U5654 (N_5654,N_5367,N_5131);
and U5655 (N_5655,N_5478,N_5309);
nand U5656 (N_5656,N_5335,N_5239);
xnor U5657 (N_5657,N_5494,N_5154);
and U5658 (N_5658,N_5268,N_5242);
xnor U5659 (N_5659,N_5256,N_5047);
or U5660 (N_5660,N_5288,N_5300);
nor U5661 (N_5661,N_5048,N_5203);
nor U5662 (N_5662,N_5383,N_5292);
xnor U5663 (N_5663,N_5236,N_5121);
nor U5664 (N_5664,N_5318,N_5423);
and U5665 (N_5665,N_5075,N_5348);
nor U5666 (N_5666,N_5148,N_5062);
nor U5667 (N_5667,N_5232,N_5223);
nor U5668 (N_5668,N_5323,N_5073);
and U5669 (N_5669,N_5436,N_5184);
nor U5670 (N_5670,N_5103,N_5126);
nor U5671 (N_5671,N_5409,N_5139);
and U5672 (N_5672,N_5095,N_5112);
or U5673 (N_5673,N_5279,N_5156);
nor U5674 (N_5674,N_5022,N_5490);
nand U5675 (N_5675,N_5331,N_5496);
or U5676 (N_5676,N_5031,N_5388);
or U5677 (N_5677,N_5410,N_5069);
nor U5678 (N_5678,N_5175,N_5337);
or U5679 (N_5679,N_5253,N_5055);
nor U5680 (N_5680,N_5476,N_5375);
xor U5681 (N_5681,N_5384,N_5246);
nor U5682 (N_5682,N_5428,N_5447);
or U5683 (N_5683,N_5467,N_5120);
and U5684 (N_5684,N_5172,N_5046);
or U5685 (N_5685,N_5109,N_5452);
xor U5686 (N_5686,N_5088,N_5217);
or U5687 (N_5687,N_5189,N_5434);
xor U5688 (N_5688,N_5387,N_5489);
nand U5689 (N_5689,N_5457,N_5341);
nand U5690 (N_5690,N_5238,N_5456);
and U5691 (N_5691,N_5374,N_5160);
nor U5692 (N_5692,N_5471,N_5284);
nor U5693 (N_5693,N_5053,N_5364);
xor U5694 (N_5694,N_5074,N_5174);
nor U5695 (N_5695,N_5477,N_5181);
and U5696 (N_5696,N_5030,N_5196);
nor U5697 (N_5697,N_5281,N_5110);
nand U5698 (N_5698,N_5219,N_5004);
and U5699 (N_5699,N_5408,N_5204);
nand U5700 (N_5700,N_5014,N_5034);
nor U5701 (N_5701,N_5229,N_5272);
nand U5702 (N_5702,N_5176,N_5205);
xnor U5703 (N_5703,N_5380,N_5278);
or U5704 (N_5704,N_5343,N_5271);
nand U5705 (N_5705,N_5361,N_5234);
xnor U5706 (N_5706,N_5011,N_5037);
nand U5707 (N_5707,N_5086,N_5140);
nor U5708 (N_5708,N_5418,N_5460);
and U5709 (N_5709,N_5221,N_5141);
nand U5710 (N_5710,N_5373,N_5049);
and U5711 (N_5711,N_5394,N_5155);
and U5712 (N_5712,N_5097,N_5442);
xnor U5713 (N_5713,N_5487,N_5129);
xnor U5714 (N_5714,N_5259,N_5041);
nor U5715 (N_5715,N_5432,N_5372);
or U5716 (N_5716,N_5329,N_5368);
and U5717 (N_5717,N_5445,N_5415);
xnor U5718 (N_5718,N_5065,N_5068);
nand U5719 (N_5719,N_5461,N_5190);
nand U5720 (N_5720,N_5224,N_5024);
and U5721 (N_5721,N_5185,N_5448);
or U5722 (N_5722,N_5414,N_5274);
nor U5723 (N_5723,N_5351,N_5444);
and U5724 (N_5724,N_5369,N_5464);
nand U5725 (N_5725,N_5170,N_5336);
nand U5726 (N_5726,N_5295,N_5235);
xor U5727 (N_5727,N_5290,N_5344);
nor U5728 (N_5728,N_5018,N_5230);
xnor U5729 (N_5729,N_5405,N_5059);
xnor U5730 (N_5730,N_5142,N_5188);
or U5731 (N_5731,N_5393,N_5173);
or U5732 (N_5732,N_5254,N_5486);
or U5733 (N_5733,N_5379,N_5003);
nand U5734 (N_5734,N_5001,N_5347);
nand U5735 (N_5735,N_5475,N_5006);
nand U5736 (N_5736,N_5454,N_5153);
xor U5737 (N_5737,N_5339,N_5286);
nand U5738 (N_5738,N_5458,N_5462);
nand U5739 (N_5739,N_5089,N_5420);
nand U5740 (N_5740,N_5473,N_5416);
nand U5741 (N_5741,N_5376,N_5195);
nand U5742 (N_5742,N_5491,N_5426);
nand U5743 (N_5743,N_5025,N_5033);
or U5744 (N_5744,N_5115,N_5026);
nor U5745 (N_5745,N_5200,N_5137);
xor U5746 (N_5746,N_5422,N_5326);
and U5747 (N_5747,N_5262,N_5247);
nand U5748 (N_5748,N_5389,N_5319);
or U5749 (N_5749,N_5044,N_5032);
nor U5750 (N_5750,N_5123,N_5091);
nor U5751 (N_5751,N_5158,N_5496);
or U5752 (N_5752,N_5295,N_5232);
and U5753 (N_5753,N_5250,N_5115);
or U5754 (N_5754,N_5186,N_5266);
nor U5755 (N_5755,N_5058,N_5063);
nor U5756 (N_5756,N_5451,N_5042);
nor U5757 (N_5757,N_5288,N_5472);
and U5758 (N_5758,N_5135,N_5279);
xnor U5759 (N_5759,N_5249,N_5071);
xor U5760 (N_5760,N_5260,N_5188);
and U5761 (N_5761,N_5025,N_5073);
or U5762 (N_5762,N_5371,N_5318);
xor U5763 (N_5763,N_5108,N_5218);
xor U5764 (N_5764,N_5375,N_5118);
nand U5765 (N_5765,N_5269,N_5205);
or U5766 (N_5766,N_5448,N_5492);
nand U5767 (N_5767,N_5377,N_5425);
nand U5768 (N_5768,N_5280,N_5432);
or U5769 (N_5769,N_5023,N_5377);
nand U5770 (N_5770,N_5386,N_5041);
nand U5771 (N_5771,N_5349,N_5263);
nor U5772 (N_5772,N_5425,N_5114);
and U5773 (N_5773,N_5383,N_5180);
and U5774 (N_5774,N_5158,N_5218);
xor U5775 (N_5775,N_5346,N_5427);
or U5776 (N_5776,N_5032,N_5448);
xor U5777 (N_5777,N_5485,N_5483);
nand U5778 (N_5778,N_5002,N_5495);
and U5779 (N_5779,N_5342,N_5068);
nor U5780 (N_5780,N_5345,N_5284);
or U5781 (N_5781,N_5071,N_5345);
or U5782 (N_5782,N_5393,N_5325);
xor U5783 (N_5783,N_5153,N_5437);
or U5784 (N_5784,N_5083,N_5144);
and U5785 (N_5785,N_5022,N_5491);
or U5786 (N_5786,N_5240,N_5263);
xor U5787 (N_5787,N_5040,N_5007);
nand U5788 (N_5788,N_5329,N_5371);
nand U5789 (N_5789,N_5250,N_5441);
nand U5790 (N_5790,N_5377,N_5182);
or U5791 (N_5791,N_5402,N_5259);
or U5792 (N_5792,N_5229,N_5110);
nor U5793 (N_5793,N_5199,N_5475);
and U5794 (N_5794,N_5245,N_5341);
nor U5795 (N_5795,N_5326,N_5318);
nor U5796 (N_5796,N_5040,N_5394);
nand U5797 (N_5797,N_5246,N_5144);
and U5798 (N_5798,N_5315,N_5326);
or U5799 (N_5799,N_5423,N_5030);
nand U5800 (N_5800,N_5196,N_5229);
nand U5801 (N_5801,N_5187,N_5071);
nand U5802 (N_5802,N_5013,N_5387);
nand U5803 (N_5803,N_5214,N_5274);
and U5804 (N_5804,N_5126,N_5211);
nand U5805 (N_5805,N_5323,N_5091);
xnor U5806 (N_5806,N_5078,N_5477);
or U5807 (N_5807,N_5440,N_5033);
nand U5808 (N_5808,N_5424,N_5179);
xnor U5809 (N_5809,N_5089,N_5367);
nor U5810 (N_5810,N_5388,N_5016);
and U5811 (N_5811,N_5412,N_5422);
or U5812 (N_5812,N_5120,N_5300);
and U5813 (N_5813,N_5299,N_5460);
xnor U5814 (N_5814,N_5045,N_5025);
xor U5815 (N_5815,N_5360,N_5430);
or U5816 (N_5816,N_5293,N_5241);
nor U5817 (N_5817,N_5068,N_5476);
and U5818 (N_5818,N_5327,N_5110);
xor U5819 (N_5819,N_5101,N_5300);
and U5820 (N_5820,N_5396,N_5334);
nand U5821 (N_5821,N_5122,N_5164);
nor U5822 (N_5822,N_5395,N_5193);
nand U5823 (N_5823,N_5083,N_5443);
nand U5824 (N_5824,N_5395,N_5272);
and U5825 (N_5825,N_5032,N_5420);
nand U5826 (N_5826,N_5105,N_5298);
and U5827 (N_5827,N_5280,N_5169);
or U5828 (N_5828,N_5446,N_5164);
xnor U5829 (N_5829,N_5006,N_5396);
or U5830 (N_5830,N_5318,N_5224);
nand U5831 (N_5831,N_5219,N_5260);
xor U5832 (N_5832,N_5306,N_5257);
or U5833 (N_5833,N_5365,N_5485);
nor U5834 (N_5834,N_5069,N_5417);
xor U5835 (N_5835,N_5391,N_5116);
or U5836 (N_5836,N_5200,N_5392);
or U5837 (N_5837,N_5484,N_5038);
or U5838 (N_5838,N_5312,N_5378);
nor U5839 (N_5839,N_5305,N_5027);
nand U5840 (N_5840,N_5017,N_5346);
and U5841 (N_5841,N_5322,N_5179);
nand U5842 (N_5842,N_5279,N_5382);
nand U5843 (N_5843,N_5212,N_5260);
xnor U5844 (N_5844,N_5241,N_5384);
nand U5845 (N_5845,N_5284,N_5292);
or U5846 (N_5846,N_5296,N_5279);
xnor U5847 (N_5847,N_5371,N_5495);
or U5848 (N_5848,N_5071,N_5295);
nand U5849 (N_5849,N_5485,N_5122);
nand U5850 (N_5850,N_5253,N_5422);
and U5851 (N_5851,N_5462,N_5450);
nor U5852 (N_5852,N_5127,N_5425);
or U5853 (N_5853,N_5144,N_5159);
nand U5854 (N_5854,N_5230,N_5330);
or U5855 (N_5855,N_5069,N_5346);
nor U5856 (N_5856,N_5101,N_5109);
and U5857 (N_5857,N_5065,N_5349);
xnor U5858 (N_5858,N_5204,N_5396);
xnor U5859 (N_5859,N_5464,N_5057);
or U5860 (N_5860,N_5055,N_5039);
nand U5861 (N_5861,N_5442,N_5035);
xor U5862 (N_5862,N_5004,N_5234);
nand U5863 (N_5863,N_5376,N_5409);
nor U5864 (N_5864,N_5226,N_5243);
and U5865 (N_5865,N_5076,N_5353);
or U5866 (N_5866,N_5423,N_5350);
and U5867 (N_5867,N_5455,N_5324);
xor U5868 (N_5868,N_5131,N_5446);
or U5869 (N_5869,N_5211,N_5355);
and U5870 (N_5870,N_5013,N_5128);
xnor U5871 (N_5871,N_5415,N_5131);
or U5872 (N_5872,N_5331,N_5111);
nand U5873 (N_5873,N_5460,N_5470);
nand U5874 (N_5874,N_5324,N_5033);
or U5875 (N_5875,N_5055,N_5273);
nor U5876 (N_5876,N_5157,N_5088);
xnor U5877 (N_5877,N_5424,N_5365);
nor U5878 (N_5878,N_5052,N_5464);
xor U5879 (N_5879,N_5234,N_5257);
xor U5880 (N_5880,N_5400,N_5071);
nand U5881 (N_5881,N_5124,N_5463);
nor U5882 (N_5882,N_5096,N_5015);
xnor U5883 (N_5883,N_5459,N_5162);
nand U5884 (N_5884,N_5476,N_5249);
or U5885 (N_5885,N_5167,N_5432);
xor U5886 (N_5886,N_5233,N_5351);
or U5887 (N_5887,N_5289,N_5397);
nand U5888 (N_5888,N_5487,N_5495);
or U5889 (N_5889,N_5105,N_5236);
or U5890 (N_5890,N_5037,N_5056);
nor U5891 (N_5891,N_5371,N_5203);
nor U5892 (N_5892,N_5047,N_5117);
nand U5893 (N_5893,N_5006,N_5057);
or U5894 (N_5894,N_5124,N_5233);
xnor U5895 (N_5895,N_5116,N_5241);
nor U5896 (N_5896,N_5085,N_5223);
nor U5897 (N_5897,N_5373,N_5311);
and U5898 (N_5898,N_5406,N_5068);
nand U5899 (N_5899,N_5345,N_5495);
nor U5900 (N_5900,N_5086,N_5189);
or U5901 (N_5901,N_5286,N_5280);
or U5902 (N_5902,N_5449,N_5401);
and U5903 (N_5903,N_5446,N_5056);
and U5904 (N_5904,N_5491,N_5414);
nor U5905 (N_5905,N_5435,N_5339);
nand U5906 (N_5906,N_5089,N_5345);
or U5907 (N_5907,N_5122,N_5416);
or U5908 (N_5908,N_5086,N_5412);
or U5909 (N_5909,N_5393,N_5075);
or U5910 (N_5910,N_5418,N_5060);
or U5911 (N_5911,N_5495,N_5037);
and U5912 (N_5912,N_5318,N_5352);
or U5913 (N_5913,N_5381,N_5310);
and U5914 (N_5914,N_5373,N_5112);
and U5915 (N_5915,N_5285,N_5281);
xnor U5916 (N_5916,N_5219,N_5454);
xor U5917 (N_5917,N_5029,N_5334);
nand U5918 (N_5918,N_5075,N_5338);
xnor U5919 (N_5919,N_5010,N_5064);
nand U5920 (N_5920,N_5193,N_5094);
and U5921 (N_5921,N_5014,N_5141);
or U5922 (N_5922,N_5488,N_5307);
nor U5923 (N_5923,N_5310,N_5496);
or U5924 (N_5924,N_5203,N_5370);
nand U5925 (N_5925,N_5149,N_5274);
or U5926 (N_5926,N_5151,N_5253);
xor U5927 (N_5927,N_5410,N_5240);
nor U5928 (N_5928,N_5272,N_5183);
and U5929 (N_5929,N_5361,N_5055);
or U5930 (N_5930,N_5291,N_5418);
or U5931 (N_5931,N_5492,N_5342);
nor U5932 (N_5932,N_5059,N_5280);
nor U5933 (N_5933,N_5216,N_5280);
nor U5934 (N_5934,N_5039,N_5324);
nand U5935 (N_5935,N_5386,N_5089);
nor U5936 (N_5936,N_5327,N_5428);
nand U5937 (N_5937,N_5032,N_5464);
xnor U5938 (N_5938,N_5289,N_5245);
nor U5939 (N_5939,N_5191,N_5245);
xnor U5940 (N_5940,N_5076,N_5082);
and U5941 (N_5941,N_5366,N_5338);
nand U5942 (N_5942,N_5362,N_5167);
and U5943 (N_5943,N_5143,N_5320);
nand U5944 (N_5944,N_5087,N_5321);
and U5945 (N_5945,N_5420,N_5065);
nor U5946 (N_5946,N_5444,N_5415);
nand U5947 (N_5947,N_5267,N_5074);
nand U5948 (N_5948,N_5357,N_5484);
xnor U5949 (N_5949,N_5178,N_5074);
xnor U5950 (N_5950,N_5187,N_5364);
nor U5951 (N_5951,N_5402,N_5229);
or U5952 (N_5952,N_5239,N_5319);
xor U5953 (N_5953,N_5413,N_5309);
or U5954 (N_5954,N_5282,N_5013);
and U5955 (N_5955,N_5487,N_5464);
or U5956 (N_5956,N_5443,N_5498);
and U5957 (N_5957,N_5360,N_5200);
nand U5958 (N_5958,N_5112,N_5483);
and U5959 (N_5959,N_5188,N_5144);
nand U5960 (N_5960,N_5457,N_5232);
or U5961 (N_5961,N_5351,N_5473);
or U5962 (N_5962,N_5032,N_5415);
nand U5963 (N_5963,N_5277,N_5223);
nand U5964 (N_5964,N_5304,N_5442);
or U5965 (N_5965,N_5099,N_5420);
xor U5966 (N_5966,N_5285,N_5465);
and U5967 (N_5967,N_5108,N_5289);
or U5968 (N_5968,N_5075,N_5418);
xor U5969 (N_5969,N_5209,N_5340);
nor U5970 (N_5970,N_5060,N_5372);
nor U5971 (N_5971,N_5236,N_5487);
nand U5972 (N_5972,N_5274,N_5346);
or U5973 (N_5973,N_5326,N_5022);
or U5974 (N_5974,N_5233,N_5044);
nand U5975 (N_5975,N_5273,N_5194);
or U5976 (N_5976,N_5402,N_5294);
or U5977 (N_5977,N_5468,N_5106);
or U5978 (N_5978,N_5272,N_5039);
and U5979 (N_5979,N_5455,N_5306);
xnor U5980 (N_5980,N_5062,N_5006);
or U5981 (N_5981,N_5248,N_5291);
and U5982 (N_5982,N_5485,N_5172);
or U5983 (N_5983,N_5410,N_5436);
and U5984 (N_5984,N_5246,N_5256);
xor U5985 (N_5985,N_5301,N_5416);
xor U5986 (N_5986,N_5241,N_5287);
nor U5987 (N_5987,N_5251,N_5210);
and U5988 (N_5988,N_5436,N_5062);
nand U5989 (N_5989,N_5467,N_5043);
xnor U5990 (N_5990,N_5222,N_5145);
or U5991 (N_5991,N_5216,N_5253);
xnor U5992 (N_5992,N_5343,N_5121);
nand U5993 (N_5993,N_5336,N_5094);
nor U5994 (N_5994,N_5443,N_5447);
and U5995 (N_5995,N_5367,N_5352);
and U5996 (N_5996,N_5129,N_5185);
nor U5997 (N_5997,N_5239,N_5158);
and U5998 (N_5998,N_5056,N_5411);
nand U5999 (N_5999,N_5388,N_5334);
nor U6000 (N_6000,N_5802,N_5819);
or U6001 (N_6001,N_5542,N_5950);
nor U6002 (N_6002,N_5522,N_5554);
and U6003 (N_6003,N_5866,N_5698);
nor U6004 (N_6004,N_5711,N_5713);
and U6005 (N_6005,N_5971,N_5995);
nor U6006 (N_6006,N_5692,N_5694);
nor U6007 (N_6007,N_5619,N_5920);
nand U6008 (N_6008,N_5651,N_5500);
nor U6009 (N_6009,N_5839,N_5818);
nand U6010 (N_6010,N_5639,N_5567);
nor U6011 (N_6011,N_5641,N_5759);
nor U6012 (N_6012,N_5533,N_5530);
or U6013 (N_6013,N_5836,N_5782);
nand U6014 (N_6014,N_5784,N_5805);
or U6015 (N_6015,N_5521,N_5709);
and U6016 (N_6016,N_5792,N_5969);
nand U6017 (N_6017,N_5664,N_5745);
nor U6018 (N_6018,N_5677,N_5555);
nor U6019 (N_6019,N_5510,N_5863);
and U6020 (N_6020,N_5850,N_5826);
or U6021 (N_6021,N_5642,N_5848);
or U6022 (N_6022,N_5882,N_5993);
nand U6023 (N_6023,N_5874,N_5879);
xnor U6024 (N_6024,N_5520,N_5858);
or U6025 (N_6025,N_5734,N_5925);
xor U6026 (N_6026,N_5987,N_5777);
nor U6027 (N_6027,N_5684,N_5944);
nand U6028 (N_6028,N_5834,N_5615);
and U6029 (N_6029,N_5962,N_5600);
nor U6030 (N_6030,N_5970,N_5561);
nand U6031 (N_6031,N_5785,N_5643);
nand U6032 (N_6032,N_5742,N_5838);
xor U6033 (N_6033,N_5895,N_5655);
and U6034 (N_6034,N_5562,N_5748);
nor U6035 (N_6035,N_5652,N_5846);
or U6036 (N_6036,N_5775,N_5699);
and U6037 (N_6037,N_5519,N_5945);
nand U6038 (N_6038,N_5978,N_5931);
and U6039 (N_6039,N_5956,N_5597);
xor U6040 (N_6040,N_5587,N_5695);
and U6041 (N_6041,N_5772,N_5531);
or U6042 (N_6042,N_5508,N_5766);
or U6043 (N_6043,N_5549,N_5696);
or U6044 (N_6044,N_5509,N_5608);
and U6045 (N_6045,N_5660,N_5718);
and U6046 (N_6046,N_5973,N_5813);
or U6047 (N_6047,N_5963,N_5682);
and U6048 (N_6048,N_5663,N_5983);
nand U6049 (N_6049,N_5765,N_5602);
or U6050 (N_6050,N_5793,N_5937);
nor U6051 (N_6051,N_5653,N_5590);
xor U6052 (N_6052,N_5690,N_5881);
nor U6053 (N_6053,N_5708,N_5853);
nor U6054 (N_6054,N_5706,N_5659);
nor U6055 (N_6055,N_5800,N_5909);
or U6056 (N_6056,N_5668,N_5592);
and U6057 (N_6057,N_5816,N_5598);
nand U6058 (N_6058,N_5893,N_5605);
xnor U6059 (N_6059,N_5683,N_5886);
nand U6060 (N_6060,N_5612,N_5907);
nor U6061 (N_6061,N_5649,N_5671);
and U6062 (N_6062,N_5992,N_5676);
nand U6063 (N_6063,N_5725,N_5941);
xnor U6064 (N_6064,N_5908,N_5697);
nor U6065 (N_6065,N_5568,N_5905);
nor U6066 (N_6066,N_5638,N_5832);
and U6067 (N_6067,N_5722,N_5923);
and U6068 (N_6068,N_5753,N_5936);
xor U6069 (N_6069,N_5583,N_5679);
and U6070 (N_6070,N_5998,N_5825);
xor U6071 (N_6071,N_5943,N_5735);
or U6072 (N_6072,N_5762,N_5738);
and U6073 (N_6073,N_5505,N_5861);
nand U6074 (N_6074,N_5835,N_5894);
nand U6075 (N_6075,N_5644,N_5565);
nor U6076 (N_6076,N_5873,N_5952);
nor U6077 (N_6077,N_5661,N_5974);
nor U6078 (N_6078,N_5593,N_5501);
or U6079 (N_6079,N_5575,N_5731);
or U6080 (N_6080,N_5740,N_5650);
or U6081 (N_6081,N_5871,N_5657);
xor U6082 (N_6082,N_5914,N_5552);
nand U6083 (N_6083,N_5700,N_5573);
nand U6084 (N_6084,N_5902,N_5537);
nor U6085 (N_6085,N_5877,N_5566);
and U6086 (N_6086,N_5553,N_5633);
nand U6087 (N_6087,N_5511,N_5716);
nand U6088 (N_6088,N_5609,N_5704);
nand U6089 (N_6089,N_5724,N_5623);
nand U6090 (N_6090,N_5751,N_5559);
xor U6091 (N_6091,N_5527,N_5997);
nor U6092 (N_6092,N_5647,N_5930);
and U6093 (N_6093,N_5535,N_5670);
xor U6094 (N_6094,N_5747,N_5551);
or U6095 (N_6095,N_5662,N_5958);
nand U6096 (N_6096,N_5582,N_5658);
nor U6097 (N_6097,N_5611,N_5667);
nand U6098 (N_6098,N_5924,N_5955);
nand U6099 (N_6099,N_5548,N_5788);
and U6100 (N_6100,N_5584,N_5812);
or U6101 (N_6101,N_5875,N_5932);
nand U6102 (N_6102,N_5991,N_5778);
xnor U6103 (N_6103,N_5984,N_5547);
nand U6104 (N_6104,N_5503,N_5860);
or U6105 (N_6105,N_5940,N_5712);
nor U6106 (N_6106,N_5870,N_5769);
nor U6107 (N_6107,N_5733,N_5786);
nor U6108 (N_6108,N_5539,N_5701);
nand U6109 (N_6109,N_5814,N_5915);
or U6110 (N_6110,N_5571,N_5981);
and U6111 (N_6111,N_5545,N_5514);
nor U6112 (N_6112,N_5746,N_5689);
and U6113 (N_6113,N_5960,N_5631);
xor U6114 (N_6114,N_5703,N_5666);
nand U6115 (N_6115,N_5804,N_5726);
or U6116 (N_6116,N_5938,N_5911);
or U6117 (N_6117,N_5616,N_5841);
nand U6118 (N_6118,N_5538,N_5946);
nor U6119 (N_6119,N_5771,N_5904);
and U6120 (N_6120,N_5688,N_5933);
xnor U6121 (N_6121,N_5576,N_5687);
nand U6122 (N_6122,N_5577,N_5790);
xnor U6123 (N_6123,N_5743,N_5961);
or U6124 (N_6124,N_5516,N_5648);
nand U6125 (N_6125,N_5868,N_5621);
or U6126 (N_6126,N_5730,N_5614);
xnor U6127 (N_6127,N_5986,N_5756);
nand U6128 (N_6128,N_5764,N_5957);
xor U6129 (N_6129,N_5721,N_5729);
xor U6130 (N_6130,N_5705,N_5919);
nand U6131 (N_6131,N_5796,N_5680);
or U6132 (N_6132,N_5646,N_5912);
and U6133 (N_6133,N_5770,N_5776);
nor U6134 (N_6134,N_5601,N_5989);
or U6135 (N_6135,N_5557,N_5768);
or U6136 (N_6136,N_5578,N_5710);
nand U6137 (N_6137,N_5686,N_5821);
or U6138 (N_6138,N_5791,N_5885);
xor U6139 (N_6139,N_5951,N_5596);
and U6140 (N_6140,N_5723,N_5669);
nor U6141 (N_6141,N_5574,N_5580);
and U6142 (N_6142,N_5595,N_5857);
nor U6143 (N_6143,N_5529,N_5840);
or U6144 (N_6144,N_5627,N_5604);
xor U6145 (N_6145,N_5843,N_5675);
nor U6146 (N_6146,N_5720,N_5833);
nand U6147 (N_6147,N_5900,N_5532);
nand U6148 (N_6148,N_5588,N_5524);
nor U6149 (N_6149,N_5618,N_5523);
nand U6150 (N_6150,N_5851,N_5589);
xnor U6151 (N_6151,N_5996,N_5854);
nand U6152 (N_6152,N_5613,N_5632);
nor U6153 (N_6153,N_5579,N_5635);
nor U6154 (N_6154,N_5672,N_5717);
or U6155 (N_6155,N_5967,N_5829);
nand U6156 (N_6156,N_5954,N_5727);
nand U6157 (N_6157,N_5855,N_5830);
xor U6158 (N_6158,N_5892,N_5599);
xor U6159 (N_6159,N_5630,N_5528);
and U6160 (N_6160,N_5922,N_5849);
nand U6161 (N_6161,N_5787,N_5773);
and U6162 (N_6162,N_5808,N_5707);
or U6163 (N_6163,N_5517,N_5719);
nor U6164 (N_6164,N_5678,N_5525);
nor U6165 (N_6165,N_5585,N_5736);
nor U6166 (N_6166,N_5750,N_5896);
and U6167 (N_6167,N_5754,N_5815);
xor U6168 (N_6168,N_5901,N_5506);
and U6169 (N_6169,N_5691,N_5757);
or U6170 (N_6170,N_5888,N_5864);
xor U6171 (N_6171,N_5890,N_5982);
or U6172 (N_6172,N_5801,N_5610);
and U6173 (N_6173,N_5968,N_5674);
xor U6174 (N_6174,N_5789,N_5856);
xnor U6175 (N_6175,N_5564,N_5994);
xor U6176 (N_6176,N_5640,N_5887);
nor U6177 (N_6177,N_5504,N_5617);
xor U6178 (N_6178,N_5779,N_5763);
or U6179 (N_6179,N_5507,N_5570);
or U6180 (N_6180,N_5884,N_5999);
and U6181 (N_6181,N_5947,N_5737);
xnor U6182 (N_6182,N_5809,N_5827);
xnor U6183 (N_6183,N_5546,N_5822);
or U6184 (N_6184,N_5867,N_5990);
xnor U6185 (N_6185,N_5797,N_5685);
nand U6186 (N_6186,N_5603,N_5847);
nor U6187 (N_6187,N_5558,N_5556);
or U6188 (N_6188,N_5512,N_5714);
nand U6189 (N_6189,N_5965,N_5979);
or U6190 (N_6190,N_5903,N_5752);
and U6191 (N_6191,N_5628,N_5810);
or U6192 (N_6192,N_5749,N_5693);
xnor U6193 (N_6193,N_5935,N_5803);
nand U6194 (N_6194,N_5844,N_5928);
and U6195 (N_6195,N_5852,N_5744);
nand U6196 (N_6196,N_5629,N_5767);
or U6197 (N_6197,N_5980,N_5591);
nand U6198 (N_6198,N_5972,N_5761);
nand U6199 (N_6199,N_5625,N_5891);
xnor U6200 (N_6200,N_5518,N_5702);
xnor U6201 (N_6201,N_5794,N_5654);
nand U6202 (N_6202,N_5883,N_5799);
and U6203 (N_6203,N_5926,N_5502);
nand U6204 (N_6204,N_5878,N_5939);
nand U6205 (N_6205,N_5637,N_5934);
and U6206 (N_6206,N_5634,N_5820);
and U6207 (N_6207,N_5550,N_5910);
nor U6208 (N_6208,N_5774,N_5927);
and U6209 (N_6209,N_5942,N_5948);
xor U6210 (N_6210,N_5798,N_5917);
nor U6211 (N_6211,N_5918,N_5544);
xor U6212 (N_6212,N_5869,N_5606);
nand U6213 (N_6213,N_5607,N_5966);
nor U6214 (N_6214,N_5572,N_5586);
and U6215 (N_6215,N_5828,N_5862);
nand U6216 (N_6216,N_5536,N_5673);
nor U6217 (N_6217,N_5758,N_5859);
xor U6218 (N_6218,N_5715,N_5656);
nor U6219 (N_6219,N_5817,N_5949);
or U6220 (N_6220,N_5824,N_5732);
or U6221 (N_6221,N_5897,N_5959);
nand U6222 (N_6222,N_5515,N_5977);
nand U6223 (N_6223,N_5889,N_5921);
and U6224 (N_6224,N_5837,N_5880);
and U6225 (N_6225,N_5563,N_5755);
or U6226 (N_6226,N_5540,N_5872);
and U6227 (N_6227,N_5842,N_5728);
nand U6228 (N_6228,N_5645,N_5665);
nand U6229 (N_6229,N_5526,N_5964);
or U6230 (N_6230,N_5845,N_5541);
xor U6231 (N_6231,N_5622,N_5899);
xnor U6232 (N_6232,N_5906,N_5985);
and U6233 (N_6233,N_5534,N_5953);
or U6234 (N_6234,N_5913,N_5624);
or U6235 (N_6235,N_5975,N_5560);
and U6236 (N_6236,N_5543,N_5636);
xnor U6237 (N_6237,N_5916,N_5806);
xnor U6238 (N_6238,N_5739,N_5831);
xnor U6239 (N_6239,N_5795,N_5594);
nand U6240 (N_6240,N_5898,N_5988);
or U6241 (N_6241,N_5626,N_5929);
or U6242 (N_6242,N_5569,N_5741);
or U6243 (N_6243,N_5807,N_5581);
xnor U6244 (N_6244,N_5780,N_5513);
or U6245 (N_6245,N_5681,N_5620);
xor U6246 (N_6246,N_5876,N_5823);
nor U6247 (N_6247,N_5811,N_5865);
nand U6248 (N_6248,N_5783,N_5781);
or U6249 (N_6249,N_5976,N_5760);
nand U6250 (N_6250,N_5826,N_5761);
or U6251 (N_6251,N_5664,N_5958);
xnor U6252 (N_6252,N_5765,N_5844);
or U6253 (N_6253,N_5885,N_5588);
xor U6254 (N_6254,N_5750,N_5909);
nand U6255 (N_6255,N_5623,N_5954);
nor U6256 (N_6256,N_5754,N_5712);
and U6257 (N_6257,N_5841,N_5630);
nand U6258 (N_6258,N_5836,N_5678);
nand U6259 (N_6259,N_5515,N_5662);
xor U6260 (N_6260,N_5512,N_5603);
nand U6261 (N_6261,N_5876,N_5564);
or U6262 (N_6262,N_5817,N_5769);
nand U6263 (N_6263,N_5925,N_5638);
nand U6264 (N_6264,N_5968,N_5671);
nor U6265 (N_6265,N_5931,N_5526);
and U6266 (N_6266,N_5815,N_5723);
nand U6267 (N_6267,N_5958,N_5887);
xnor U6268 (N_6268,N_5804,N_5838);
nor U6269 (N_6269,N_5931,N_5878);
and U6270 (N_6270,N_5563,N_5680);
nor U6271 (N_6271,N_5736,N_5802);
or U6272 (N_6272,N_5685,N_5714);
xnor U6273 (N_6273,N_5541,N_5825);
xor U6274 (N_6274,N_5699,N_5658);
nor U6275 (N_6275,N_5858,N_5564);
nand U6276 (N_6276,N_5691,N_5551);
or U6277 (N_6277,N_5922,N_5776);
and U6278 (N_6278,N_5940,N_5655);
xor U6279 (N_6279,N_5787,N_5930);
or U6280 (N_6280,N_5872,N_5706);
or U6281 (N_6281,N_5557,N_5838);
nor U6282 (N_6282,N_5966,N_5928);
xor U6283 (N_6283,N_5646,N_5527);
nor U6284 (N_6284,N_5713,N_5520);
or U6285 (N_6285,N_5794,N_5692);
xor U6286 (N_6286,N_5810,N_5867);
nand U6287 (N_6287,N_5566,N_5831);
nand U6288 (N_6288,N_5537,N_5758);
or U6289 (N_6289,N_5683,N_5578);
and U6290 (N_6290,N_5738,N_5655);
xor U6291 (N_6291,N_5526,N_5703);
or U6292 (N_6292,N_5842,N_5585);
or U6293 (N_6293,N_5723,N_5747);
nor U6294 (N_6294,N_5904,N_5611);
nor U6295 (N_6295,N_5868,N_5672);
or U6296 (N_6296,N_5549,N_5686);
nor U6297 (N_6297,N_5895,N_5750);
xor U6298 (N_6298,N_5536,N_5868);
and U6299 (N_6299,N_5625,N_5610);
or U6300 (N_6300,N_5776,N_5915);
nor U6301 (N_6301,N_5936,N_5752);
nand U6302 (N_6302,N_5575,N_5689);
nand U6303 (N_6303,N_5787,N_5786);
xnor U6304 (N_6304,N_5853,N_5866);
or U6305 (N_6305,N_5724,N_5505);
xnor U6306 (N_6306,N_5890,N_5529);
nor U6307 (N_6307,N_5692,N_5503);
xor U6308 (N_6308,N_5617,N_5786);
nand U6309 (N_6309,N_5747,N_5629);
or U6310 (N_6310,N_5553,N_5897);
xnor U6311 (N_6311,N_5963,N_5814);
nor U6312 (N_6312,N_5861,N_5916);
or U6313 (N_6313,N_5561,N_5827);
or U6314 (N_6314,N_5961,N_5987);
nand U6315 (N_6315,N_5991,N_5841);
nor U6316 (N_6316,N_5558,N_5598);
xnor U6317 (N_6317,N_5708,N_5549);
nand U6318 (N_6318,N_5507,N_5654);
or U6319 (N_6319,N_5751,N_5511);
nor U6320 (N_6320,N_5773,N_5918);
xor U6321 (N_6321,N_5704,N_5504);
nand U6322 (N_6322,N_5795,N_5742);
nand U6323 (N_6323,N_5727,N_5601);
or U6324 (N_6324,N_5797,N_5922);
nor U6325 (N_6325,N_5560,N_5509);
or U6326 (N_6326,N_5942,N_5542);
xor U6327 (N_6327,N_5929,N_5551);
and U6328 (N_6328,N_5710,N_5745);
and U6329 (N_6329,N_5596,N_5781);
or U6330 (N_6330,N_5671,N_5638);
nor U6331 (N_6331,N_5755,N_5988);
xnor U6332 (N_6332,N_5614,N_5735);
or U6333 (N_6333,N_5821,N_5588);
and U6334 (N_6334,N_5953,N_5533);
xor U6335 (N_6335,N_5845,N_5607);
xnor U6336 (N_6336,N_5863,N_5827);
xor U6337 (N_6337,N_5629,N_5773);
nor U6338 (N_6338,N_5714,N_5883);
nor U6339 (N_6339,N_5809,N_5636);
nor U6340 (N_6340,N_5571,N_5848);
nand U6341 (N_6341,N_5846,N_5539);
or U6342 (N_6342,N_5929,N_5710);
and U6343 (N_6343,N_5802,N_5848);
or U6344 (N_6344,N_5679,N_5775);
and U6345 (N_6345,N_5863,N_5902);
xor U6346 (N_6346,N_5896,N_5752);
nand U6347 (N_6347,N_5539,N_5838);
and U6348 (N_6348,N_5861,N_5730);
nand U6349 (N_6349,N_5774,N_5904);
xnor U6350 (N_6350,N_5593,N_5964);
nand U6351 (N_6351,N_5986,N_5873);
or U6352 (N_6352,N_5849,N_5956);
nor U6353 (N_6353,N_5516,N_5999);
or U6354 (N_6354,N_5726,N_5612);
xor U6355 (N_6355,N_5929,N_5849);
and U6356 (N_6356,N_5989,N_5552);
nand U6357 (N_6357,N_5506,N_5508);
nor U6358 (N_6358,N_5843,N_5880);
or U6359 (N_6359,N_5826,N_5824);
nand U6360 (N_6360,N_5849,N_5825);
nand U6361 (N_6361,N_5583,N_5714);
xnor U6362 (N_6362,N_5698,N_5770);
or U6363 (N_6363,N_5588,N_5928);
and U6364 (N_6364,N_5701,N_5599);
nand U6365 (N_6365,N_5605,N_5519);
xor U6366 (N_6366,N_5540,N_5664);
nand U6367 (N_6367,N_5975,N_5806);
or U6368 (N_6368,N_5794,N_5729);
xnor U6369 (N_6369,N_5754,N_5613);
and U6370 (N_6370,N_5921,N_5688);
nand U6371 (N_6371,N_5948,N_5665);
xor U6372 (N_6372,N_5744,N_5842);
xor U6373 (N_6373,N_5604,N_5713);
or U6374 (N_6374,N_5830,N_5510);
and U6375 (N_6375,N_5780,N_5800);
xnor U6376 (N_6376,N_5616,N_5851);
or U6377 (N_6377,N_5618,N_5824);
and U6378 (N_6378,N_5781,N_5541);
nand U6379 (N_6379,N_5630,N_5552);
nor U6380 (N_6380,N_5884,N_5891);
nor U6381 (N_6381,N_5809,N_5869);
or U6382 (N_6382,N_5758,N_5617);
nor U6383 (N_6383,N_5735,N_5698);
nand U6384 (N_6384,N_5886,N_5725);
nor U6385 (N_6385,N_5907,N_5908);
xor U6386 (N_6386,N_5628,N_5721);
xor U6387 (N_6387,N_5848,N_5540);
nand U6388 (N_6388,N_5861,N_5918);
xor U6389 (N_6389,N_5874,N_5542);
xnor U6390 (N_6390,N_5833,N_5614);
nor U6391 (N_6391,N_5901,N_5840);
and U6392 (N_6392,N_5857,N_5764);
or U6393 (N_6393,N_5503,N_5897);
xor U6394 (N_6394,N_5762,N_5584);
xor U6395 (N_6395,N_5916,N_5802);
nand U6396 (N_6396,N_5780,N_5649);
xnor U6397 (N_6397,N_5766,N_5687);
nand U6398 (N_6398,N_5940,N_5509);
and U6399 (N_6399,N_5885,N_5615);
nor U6400 (N_6400,N_5596,N_5835);
nor U6401 (N_6401,N_5648,N_5869);
xor U6402 (N_6402,N_5895,N_5555);
nand U6403 (N_6403,N_5779,N_5654);
xor U6404 (N_6404,N_5611,N_5728);
nand U6405 (N_6405,N_5725,N_5514);
xor U6406 (N_6406,N_5627,N_5702);
nor U6407 (N_6407,N_5709,N_5971);
and U6408 (N_6408,N_5656,N_5685);
xor U6409 (N_6409,N_5935,N_5575);
nor U6410 (N_6410,N_5854,N_5589);
or U6411 (N_6411,N_5817,N_5501);
or U6412 (N_6412,N_5913,N_5934);
nor U6413 (N_6413,N_5706,N_5735);
and U6414 (N_6414,N_5698,N_5612);
nand U6415 (N_6415,N_5515,N_5608);
nor U6416 (N_6416,N_5505,N_5837);
or U6417 (N_6417,N_5811,N_5950);
nor U6418 (N_6418,N_5743,N_5507);
and U6419 (N_6419,N_5533,N_5723);
xor U6420 (N_6420,N_5616,N_5900);
nor U6421 (N_6421,N_5717,N_5531);
and U6422 (N_6422,N_5526,N_5822);
nand U6423 (N_6423,N_5766,N_5545);
or U6424 (N_6424,N_5849,N_5902);
nor U6425 (N_6425,N_5640,N_5509);
nor U6426 (N_6426,N_5612,N_5959);
or U6427 (N_6427,N_5743,N_5691);
nand U6428 (N_6428,N_5928,N_5579);
nor U6429 (N_6429,N_5608,N_5577);
nor U6430 (N_6430,N_5913,N_5747);
or U6431 (N_6431,N_5619,N_5929);
and U6432 (N_6432,N_5592,N_5744);
and U6433 (N_6433,N_5854,N_5670);
nand U6434 (N_6434,N_5704,N_5732);
nand U6435 (N_6435,N_5978,N_5969);
xnor U6436 (N_6436,N_5789,N_5550);
xnor U6437 (N_6437,N_5718,N_5735);
and U6438 (N_6438,N_5847,N_5984);
and U6439 (N_6439,N_5803,N_5839);
or U6440 (N_6440,N_5835,N_5569);
xnor U6441 (N_6441,N_5765,N_5570);
or U6442 (N_6442,N_5964,N_5903);
or U6443 (N_6443,N_5642,N_5983);
nand U6444 (N_6444,N_5935,N_5595);
and U6445 (N_6445,N_5538,N_5713);
nand U6446 (N_6446,N_5527,N_5666);
and U6447 (N_6447,N_5604,N_5772);
or U6448 (N_6448,N_5630,N_5948);
nand U6449 (N_6449,N_5507,N_5873);
and U6450 (N_6450,N_5625,N_5565);
and U6451 (N_6451,N_5573,N_5836);
or U6452 (N_6452,N_5932,N_5798);
xnor U6453 (N_6453,N_5740,N_5856);
nor U6454 (N_6454,N_5724,N_5918);
xnor U6455 (N_6455,N_5787,N_5956);
nand U6456 (N_6456,N_5922,N_5514);
or U6457 (N_6457,N_5874,N_5791);
nor U6458 (N_6458,N_5815,N_5803);
nor U6459 (N_6459,N_5880,N_5739);
xor U6460 (N_6460,N_5950,N_5782);
xnor U6461 (N_6461,N_5963,N_5832);
xnor U6462 (N_6462,N_5902,N_5801);
and U6463 (N_6463,N_5765,N_5948);
and U6464 (N_6464,N_5683,N_5630);
nand U6465 (N_6465,N_5585,N_5918);
and U6466 (N_6466,N_5817,N_5674);
nand U6467 (N_6467,N_5823,N_5741);
nor U6468 (N_6468,N_5586,N_5981);
and U6469 (N_6469,N_5943,N_5586);
or U6470 (N_6470,N_5608,N_5847);
nor U6471 (N_6471,N_5884,N_5753);
nor U6472 (N_6472,N_5986,N_5726);
nor U6473 (N_6473,N_5662,N_5685);
or U6474 (N_6474,N_5560,N_5505);
nand U6475 (N_6475,N_5958,N_5860);
nand U6476 (N_6476,N_5565,N_5882);
or U6477 (N_6477,N_5879,N_5922);
nor U6478 (N_6478,N_5606,N_5640);
or U6479 (N_6479,N_5746,N_5930);
nor U6480 (N_6480,N_5726,N_5885);
xor U6481 (N_6481,N_5636,N_5746);
nand U6482 (N_6482,N_5972,N_5949);
xnor U6483 (N_6483,N_5836,N_5803);
and U6484 (N_6484,N_5561,N_5862);
or U6485 (N_6485,N_5949,N_5776);
or U6486 (N_6486,N_5602,N_5745);
and U6487 (N_6487,N_5614,N_5742);
or U6488 (N_6488,N_5938,N_5925);
nand U6489 (N_6489,N_5519,N_5713);
or U6490 (N_6490,N_5564,N_5568);
nor U6491 (N_6491,N_5543,N_5701);
nand U6492 (N_6492,N_5983,N_5736);
and U6493 (N_6493,N_5980,N_5535);
or U6494 (N_6494,N_5576,N_5641);
nor U6495 (N_6495,N_5863,N_5875);
nand U6496 (N_6496,N_5506,N_5752);
or U6497 (N_6497,N_5532,N_5796);
nand U6498 (N_6498,N_5809,N_5617);
nand U6499 (N_6499,N_5668,N_5643);
nand U6500 (N_6500,N_6404,N_6240);
nand U6501 (N_6501,N_6082,N_6360);
nor U6502 (N_6502,N_6416,N_6341);
and U6503 (N_6503,N_6207,N_6287);
nand U6504 (N_6504,N_6153,N_6024);
nor U6505 (N_6505,N_6047,N_6149);
nand U6506 (N_6506,N_6262,N_6395);
xor U6507 (N_6507,N_6011,N_6461);
nor U6508 (N_6508,N_6107,N_6193);
nor U6509 (N_6509,N_6392,N_6484);
and U6510 (N_6510,N_6489,N_6407);
xor U6511 (N_6511,N_6179,N_6085);
nand U6512 (N_6512,N_6091,N_6454);
or U6513 (N_6513,N_6006,N_6173);
and U6514 (N_6514,N_6297,N_6337);
nand U6515 (N_6515,N_6046,N_6374);
nand U6516 (N_6516,N_6311,N_6352);
and U6517 (N_6517,N_6401,N_6027);
or U6518 (N_6518,N_6217,N_6384);
and U6519 (N_6519,N_6100,N_6129);
nor U6520 (N_6520,N_6292,N_6277);
xnor U6521 (N_6521,N_6417,N_6368);
nand U6522 (N_6522,N_6089,N_6381);
and U6523 (N_6523,N_6005,N_6326);
or U6524 (N_6524,N_6393,N_6450);
and U6525 (N_6525,N_6069,N_6252);
nand U6526 (N_6526,N_6142,N_6034);
nor U6527 (N_6527,N_6185,N_6195);
or U6528 (N_6528,N_6075,N_6105);
nor U6529 (N_6529,N_6296,N_6446);
xor U6530 (N_6530,N_6014,N_6436);
xnor U6531 (N_6531,N_6108,N_6203);
nand U6532 (N_6532,N_6270,N_6167);
xor U6533 (N_6533,N_6044,N_6357);
and U6534 (N_6534,N_6307,N_6369);
xor U6535 (N_6535,N_6045,N_6244);
or U6536 (N_6536,N_6176,N_6397);
or U6537 (N_6537,N_6471,N_6439);
xor U6538 (N_6538,N_6229,N_6093);
nand U6539 (N_6539,N_6221,N_6135);
nor U6540 (N_6540,N_6134,N_6039);
nand U6541 (N_6541,N_6486,N_6218);
or U6542 (N_6542,N_6467,N_6268);
and U6543 (N_6543,N_6037,N_6259);
nand U6544 (N_6544,N_6377,N_6096);
nand U6545 (N_6545,N_6216,N_6498);
or U6546 (N_6546,N_6449,N_6370);
nor U6547 (N_6547,N_6480,N_6007);
nand U6548 (N_6548,N_6354,N_6121);
and U6549 (N_6549,N_6265,N_6496);
nand U6550 (N_6550,N_6049,N_6399);
or U6551 (N_6551,N_6191,N_6116);
and U6552 (N_6552,N_6257,N_6494);
or U6553 (N_6553,N_6119,N_6400);
nor U6554 (N_6554,N_6367,N_6373);
or U6555 (N_6555,N_6260,N_6474);
xor U6556 (N_6556,N_6133,N_6380);
nand U6557 (N_6557,N_6396,N_6224);
and U6558 (N_6558,N_6281,N_6302);
or U6559 (N_6559,N_6227,N_6347);
and U6560 (N_6560,N_6363,N_6452);
nand U6561 (N_6561,N_6258,N_6250);
nand U6562 (N_6562,N_6422,N_6201);
xnor U6563 (N_6563,N_6271,N_6205);
nand U6564 (N_6564,N_6033,N_6478);
xor U6565 (N_6565,N_6177,N_6414);
nand U6566 (N_6566,N_6123,N_6077);
nor U6567 (N_6567,N_6267,N_6314);
and U6568 (N_6568,N_6350,N_6237);
and U6569 (N_6569,N_6163,N_6066);
nand U6570 (N_6570,N_6055,N_6375);
and U6571 (N_6571,N_6432,N_6394);
nand U6572 (N_6572,N_6318,N_6102);
nor U6573 (N_6573,N_6194,N_6018);
nand U6574 (N_6574,N_6332,N_6025);
nand U6575 (N_6575,N_6309,N_6303);
nand U6576 (N_6576,N_6483,N_6095);
xor U6577 (N_6577,N_6162,N_6204);
and U6578 (N_6578,N_6086,N_6349);
nand U6579 (N_6579,N_6181,N_6435);
xor U6580 (N_6580,N_6264,N_6101);
and U6581 (N_6581,N_6188,N_6061);
nand U6582 (N_6582,N_6159,N_6234);
nand U6583 (N_6583,N_6021,N_6189);
or U6584 (N_6584,N_6468,N_6458);
nor U6585 (N_6585,N_6490,N_6183);
xor U6586 (N_6586,N_6273,N_6226);
nor U6587 (N_6587,N_6065,N_6158);
and U6588 (N_6588,N_6492,N_6346);
xor U6589 (N_6589,N_6012,N_6230);
or U6590 (N_6590,N_6092,N_6058);
and U6591 (N_6591,N_6481,N_6285);
and U6592 (N_6592,N_6168,N_6111);
or U6593 (N_6593,N_6245,N_6340);
and U6594 (N_6594,N_6081,N_6088);
nand U6595 (N_6595,N_6462,N_6141);
nor U6596 (N_6596,N_6317,N_6356);
and U6597 (N_6597,N_6236,N_6079);
or U6598 (N_6598,N_6109,N_6198);
nand U6599 (N_6599,N_6146,N_6387);
nor U6600 (N_6600,N_6488,N_6442);
nor U6601 (N_6601,N_6154,N_6219);
xnor U6602 (N_6602,N_6148,N_6444);
or U6603 (N_6603,N_6335,N_6054);
nand U6604 (N_6604,N_6313,N_6473);
nor U6605 (N_6605,N_6321,N_6269);
nand U6606 (N_6606,N_6115,N_6379);
nor U6607 (N_6607,N_6125,N_6160);
and U6608 (N_6608,N_6098,N_6345);
nand U6609 (N_6609,N_6113,N_6056);
and U6610 (N_6610,N_6074,N_6348);
nand U6611 (N_6611,N_6304,N_6301);
xor U6612 (N_6612,N_6080,N_6294);
xnor U6613 (N_6613,N_6283,N_6222);
or U6614 (N_6614,N_6437,N_6402);
xnor U6615 (N_6615,N_6043,N_6291);
xor U6616 (N_6616,N_6305,N_6165);
nor U6617 (N_6617,N_6094,N_6084);
nor U6618 (N_6618,N_6112,N_6275);
nor U6619 (N_6619,N_6248,N_6306);
nand U6620 (N_6620,N_6428,N_6353);
nand U6621 (N_6621,N_6124,N_6147);
and U6622 (N_6622,N_6329,N_6060);
and U6623 (N_6623,N_6213,N_6364);
xnor U6624 (N_6624,N_6434,N_6362);
nand U6625 (N_6625,N_6420,N_6122);
or U6626 (N_6626,N_6343,N_6278);
or U6627 (N_6627,N_6320,N_6310);
nor U6628 (N_6628,N_6151,N_6386);
or U6629 (N_6629,N_6425,N_6184);
and U6630 (N_6630,N_6254,N_6495);
xor U6631 (N_6631,N_6050,N_6447);
nand U6632 (N_6632,N_6186,N_6272);
xnor U6633 (N_6633,N_6336,N_6324);
or U6634 (N_6634,N_6118,N_6202);
nor U6635 (N_6635,N_6323,N_6175);
nand U6636 (N_6636,N_6015,N_6316);
nand U6637 (N_6637,N_6366,N_6456);
or U6638 (N_6638,N_6466,N_6412);
and U6639 (N_6639,N_6448,N_6126);
and U6640 (N_6640,N_6327,N_6322);
nand U6641 (N_6641,N_6064,N_6427);
or U6642 (N_6642,N_6460,N_6187);
or U6643 (N_6643,N_6090,N_6182);
or U6644 (N_6644,N_6127,N_6411);
or U6645 (N_6645,N_6274,N_6013);
and U6646 (N_6646,N_6199,N_6312);
nor U6647 (N_6647,N_6212,N_6215);
and U6648 (N_6648,N_6300,N_6433);
nand U6649 (N_6649,N_6280,N_6128);
nand U6650 (N_6650,N_6156,N_6256);
xnor U6651 (N_6651,N_6382,N_6378);
xor U6652 (N_6652,N_6443,N_6003);
xnor U6653 (N_6653,N_6228,N_6023);
and U6654 (N_6654,N_6223,N_6130);
nor U6655 (N_6655,N_6288,N_6339);
xnor U6656 (N_6656,N_6431,N_6371);
nand U6657 (N_6657,N_6491,N_6166);
nand U6658 (N_6658,N_6499,N_6405);
and U6659 (N_6659,N_6365,N_6457);
nand U6660 (N_6660,N_6197,N_6026);
xor U6661 (N_6661,N_6103,N_6251);
and U6662 (N_6662,N_6419,N_6057);
nand U6663 (N_6663,N_6106,N_6004);
nor U6664 (N_6664,N_6036,N_6476);
nor U6665 (N_6665,N_6029,N_6152);
or U6666 (N_6666,N_6235,N_6220);
xnor U6667 (N_6667,N_6247,N_6391);
or U6668 (N_6668,N_6465,N_6415);
and U6669 (N_6669,N_6242,N_6214);
or U6670 (N_6670,N_6019,N_6000);
or U6671 (N_6671,N_6208,N_6067);
nor U6672 (N_6672,N_6063,N_6286);
or U6673 (N_6673,N_6426,N_6233);
or U6674 (N_6674,N_6172,N_6136);
nor U6675 (N_6675,N_6031,N_6319);
nand U6676 (N_6676,N_6232,N_6358);
or U6677 (N_6677,N_6359,N_6464);
nand U6678 (N_6678,N_6161,N_6174);
or U6679 (N_6679,N_6487,N_6010);
xnor U6680 (N_6680,N_6351,N_6389);
or U6681 (N_6681,N_6110,N_6279);
nor U6682 (N_6682,N_6048,N_6298);
xnor U6683 (N_6683,N_6038,N_6403);
or U6684 (N_6684,N_6469,N_6209);
nor U6685 (N_6685,N_6139,N_6413);
and U6686 (N_6686,N_6051,N_6295);
or U6687 (N_6687,N_6097,N_6440);
nor U6688 (N_6688,N_6083,N_6338);
nand U6689 (N_6689,N_6143,N_6290);
nor U6690 (N_6690,N_6120,N_6241);
and U6691 (N_6691,N_6052,N_6438);
nand U6692 (N_6692,N_6087,N_6239);
and U6693 (N_6693,N_6001,N_6225);
nand U6694 (N_6694,N_6453,N_6017);
nor U6695 (N_6695,N_6164,N_6114);
xor U6696 (N_6696,N_6211,N_6390);
nor U6697 (N_6697,N_6073,N_6190);
nand U6698 (N_6698,N_6068,N_6150);
nor U6699 (N_6699,N_6497,N_6040);
nor U6700 (N_6700,N_6104,N_6059);
nand U6701 (N_6701,N_6028,N_6171);
nor U6702 (N_6702,N_6138,N_6385);
and U6703 (N_6703,N_6117,N_6410);
nor U6704 (N_6704,N_6376,N_6459);
nor U6705 (N_6705,N_6263,N_6409);
nor U6706 (N_6706,N_6016,N_6170);
or U6707 (N_6707,N_6493,N_6408);
xnor U6708 (N_6708,N_6289,N_6282);
nand U6709 (N_6709,N_6388,N_6042);
nand U6710 (N_6710,N_6423,N_6331);
and U6711 (N_6711,N_6062,N_6200);
nor U6712 (N_6712,N_6424,N_6253);
xor U6713 (N_6713,N_6406,N_6255);
or U6714 (N_6714,N_6009,N_6137);
xor U6715 (N_6715,N_6455,N_6441);
or U6716 (N_6716,N_6330,N_6210);
and U6717 (N_6717,N_6315,N_6261);
and U6718 (N_6718,N_6477,N_6002);
nor U6719 (N_6719,N_6470,N_6131);
nand U6720 (N_6720,N_6342,N_6022);
or U6721 (N_6721,N_6398,N_6430);
nand U6722 (N_6722,N_6284,N_6293);
and U6723 (N_6723,N_6020,N_6479);
xor U6724 (N_6724,N_6231,N_6078);
and U6725 (N_6725,N_6355,N_6008);
or U6726 (N_6726,N_6144,N_6032);
nor U6727 (N_6727,N_6238,N_6071);
or U6728 (N_6728,N_6145,N_6475);
nand U6729 (N_6729,N_6485,N_6372);
or U6730 (N_6730,N_6418,N_6180);
nand U6731 (N_6731,N_6482,N_6308);
and U6732 (N_6732,N_6325,N_6072);
or U6733 (N_6733,N_6196,N_6132);
and U6734 (N_6734,N_6076,N_6035);
nand U6735 (N_6735,N_6192,N_6472);
xor U6736 (N_6736,N_6429,N_6344);
xnor U6737 (N_6737,N_6041,N_6169);
or U6738 (N_6738,N_6155,N_6451);
xnor U6739 (N_6739,N_6334,N_6333);
xor U6740 (N_6740,N_6299,N_6445);
nor U6741 (N_6741,N_6206,N_6246);
or U6742 (N_6742,N_6053,N_6243);
and U6743 (N_6743,N_6140,N_6361);
or U6744 (N_6744,N_6266,N_6157);
nor U6745 (N_6745,N_6383,N_6328);
nor U6746 (N_6746,N_6070,N_6421);
xnor U6747 (N_6747,N_6030,N_6178);
xnor U6748 (N_6748,N_6099,N_6463);
xnor U6749 (N_6749,N_6276,N_6249);
xnor U6750 (N_6750,N_6124,N_6152);
xnor U6751 (N_6751,N_6173,N_6432);
xnor U6752 (N_6752,N_6338,N_6067);
nor U6753 (N_6753,N_6227,N_6388);
nand U6754 (N_6754,N_6216,N_6300);
xor U6755 (N_6755,N_6276,N_6061);
nand U6756 (N_6756,N_6086,N_6096);
nor U6757 (N_6757,N_6336,N_6062);
nor U6758 (N_6758,N_6093,N_6037);
or U6759 (N_6759,N_6282,N_6468);
nand U6760 (N_6760,N_6288,N_6250);
or U6761 (N_6761,N_6224,N_6200);
nor U6762 (N_6762,N_6313,N_6250);
nor U6763 (N_6763,N_6307,N_6267);
or U6764 (N_6764,N_6131,N_6059);
nor U6765 (N_6765,N_6201,N_6031);
nor U6766 (N_6766,N_6436,N_6238);
nor U6767 (N_6767,N_6148,N_6154);
nor U6768 (N_6768,N_6129,N_6154);
nor U6769 (N_6769,N_6388,N_6328);
nor U6770 (N_6770,N_6459,N_6479);
nand U6771 (N_6771,N_6085,N_6094);
and U6772 (N_6772,N_6168,N_6243);
nor U6773 (N_6773,N_6446,N_6162);
nor U6774 (N_6774,N_6204,N_6317);
nand U6775 (N_6775,N_6015,N_6017);
or U6776 (N_6776,N_6081,N_6328);
xor U6777 (N_6777,N_6238,N_6392);
and U6778 (N_6778,N_6298,N_6158);
nand U6779 (N_6779,N_6160,N_6203);
nand U6780 (N_6780,N_6292,N_6178);
or U6781 (N_6781,N_6200,N_6491);
or U6782 (N_6782,N_6496,N_6203);
or U6783 (N_6783,N_6335,N_6090);
and U6784 (N_6784,N_6251,N_6294);
and U6785 (N_6785,N_6198,N_6496);
xnor U6786 (N_6786,N_6472,N_6259);
and U6787 (N_6787,N_6487,N_6337);
and U6788 (N_6788,N_6384,N_6441);
or U6789 (N_6789,N_6400,N_6408);
or U6790 (N_6790,N_6093,N_6077);
or U6791 (N_6791,N_6100,N_6269);
nand U6792 (N_6792,N_6258,N_6143);
nor U6793 (N_6793,N_6196,N_6311);
nand U6794 (N_6794,N_6162,N_6411);
and U6795 (N_6795,N_6044,N_6414);
or U6796 (N_6796,N_6364,N_6357);
xor U6797 (N_6797,N_6231,N_6042);
xnor U6798 (N_6798,N_6037,N_6474);
or U6799 (N_6799,N_6073,N_6347);
nand U6800 (N_6800,N_6498,N_6151);
xnor U6801 (N_6801,N_6367,N_6461);
xor U6802 (N_6802,N_6382,N_6331);
and U6803 (N_6803,N_6497,N_6135);
or U6804 (N_6804,N_6421,N_6367);
or U6805 (N_6805,N_6276,N_6442);
and U6806 (N_6806,N_6194,N_6477);
nor U6807 (N_6807,N_6091,N_6456);
nand U6808 (N_6808,N_6004,N_6192);
nand U6809 (N_6809,N_6389,N_6446);
and U6810 (N_6810,N_6324,N_6217);
nand U6811 (N_6811,N_6126,N_6092);
xor U6812 (N_6812,N_6023,N_6018);
nand U6813 (N_6813,N_6440,N_6015);
xor U6814 (N_6814,N_6434,N_6460);
and U6815 (N_6815,N_6473,N_6179);
nand U6816 (N_6816,N_6312,N_6401);
or U6817 (N_6817,N_6196,N_6384);
or U6818 (N_6818,N_6040,N_6134);
and U6819 (N_6819,N_6435,N_6332);
xnor U6820 (N_6820,N_6300,N_6499);
nand U6821 (N_6821,N_6054,N_6465);
and U6822 (N_6822,N_6237,N_6076);
nand U6823 (N_6823,N_6094,N_6268);
or U6824 (N_6824,N_6499,N_6138);
nor U6825 (N_6825,N_6302,N_6040);
or U6826 (N_6826,N_6335,N_6263);
nand U6827 (N_6827,N_6087,N_6424);
and U6828 (N_6828,N_6017,N_6169);
nand U6829 (N_6829,N_6222,N_6255);
nand U6830 (N_6830,N_6174,N_6411);
xnor U6831 (N_6831,N_6315,N_6099);
nand U6832 (N_6832,N_6345,N_6385);
nand U6833 (N_6833,N_6447,N_6275);
xor U6834 (N_6834,N_6080,N_6499);
and U6835 (N_6835,N_6330,N_6110);
or U6836 (N_6836,N_6238,N_6177);
nand U6837 (N_6837,N_6117,N_6084);
nor U6838 (N_6838,N_6116,N_6054);
xor U6839 (N_6839,N_6290,N_6241);
xor U6840 (N_6840,N_6495,N_6384);
and U6841 (N_6841,N_6108,N_6419);
nor U6842 (N_6842,N_6075,N_6440);
xnor U6843 (N_6843,N_6348,N_6098);
nand U6844 (N_6844,N_6381,N_6232);
nor U6845 (N_6845,N_6028,N_6169);
and U6846 (N_6846,N_6275,N_6267);
nand U6847 (N_6847,N_6418,N_6298);
xor U6848 (N_6848,N_6040,N_6436);
nor U6849 (N_6849,N_6416,N_6061);
or U6850 (N_6850,N_6396,N_6262);
xor U6851 (N_6851,N_6229,N_6231);
nand U6852 (N_6852,N_6357,N_6379);
xor U6853 (N_6853,N_6098,N_6343);
xnor U6854 (N_6854,N_6061,N_6008);
xor U6855 (N_6855,N_6397,N_6323);
xor U6856 (N_6856,N_6206,N_6012);
or U6857 (N_6857,N_6154,N_6464);
nor U6858 (N_6858,N_6377,N_6294);
or U6859 (N_6859,N_6413,N_6291);
nand U6860 (N_6860,N_6348,N_6367);
nand U6861 (N_6861,N_6171,N_6293);
nand U6862 (N_6862,N_6205,N_6027);
nor U6863 (N_6863,N_6046,N_6316);
nand U6864 (N_6864,N_6117,N_6415);
xnor U6865 (N_6865,N_6172,N_6309);
nand U6866 (N_6866,N_6354,N_6372);
nand U6867 (N_6867,N_6366,N_6448);
xor U6868 (N_6868,N_6127,N_6379);
and U6869 (N_6869,N_6004,N_6273);
and U6870 (N_6870,N_6468,N_6362);
and U6871 (N_6871,N_6367,N_6213);
nand U6872 (N_6872,N_6493,N_6364);
nand U6873 (N_6873,N_6037,N_6086);
and U6874 (N_6874,N_6372,N_6155);
nand U6875 (N_6875,N_6273,N_6218);
nand U6876 (N_6876,N_6258,N_6153);
xnor U6877 (N_6877,N_6099,N_6207);
nand U6878 (N_6878,N_6454,N_6404);
nand U6879 (N_6879,N_6282,N_6218);
nor U6880 (N_6880,N_6319,N_6176);
and U6881 (N_6881,N_6297,N_6259);
or U6882 (N_6882,N_6414,N_6411);
nand U6883 (N_6883,N_6077,N_6103);
nor U6884 (N_6884,N_6324,N_6195);
xnor U6885 (N_6885,N_6407,N_6121);
and U6886 (N_6886,N_6229,N_6094);
xor U6887 (N_6887,N_6332,N_6007);
nor U6888 (N_6888,N_6357,N_6354);
nor U6889 (N_6889,N_6456,N_6241);
nor U6890 (N_6890,N_6411,N_6320);
nor U6891 (N_6891,N_6474,N_6133);
xnor U6892 (N_6892,N_6067,N_6305);
nor U6893 (N_6893,N_6335,N_6252);
xor U6894 (N_6894,N_6077,N_6069);
nand U6895 (N_6895,N_6355,N_6219);
or U6896 (N_6896,N_6096,N_6058);
or U6897 (N_6897,N_6172,N_6083);
nand U6898 (N_6898,N_6340,N_6298);
and U6899 (N_6899,N_6424,N_6223);
nand U6900 (N_6900,N_6083,N_6176);
xnor U6901 (N_6901,N_6097,N_6175);
or U6902 (N_6902,N_6117,N_6317);
xnor U6903 (N_6903,N_6073,N_6295);
and U6904 (N_6904,N_6449,N_6120);
nand U6905 (N_6905,N_6049,N_6482);
xor U6906 (N_6906,N_6464,N_6086);
and U6907 (N_6907,N_6117,N_6092);
xnor U6908 (N_6908,N_6151,N_6207);
or U6909 (N_6909,N_6410,N_6206);
nor U6910 (N_6910,N_6137,N_6100);
and U6911 (N_6911,N_6139,N_6407);
or U6912 (N_6912,N_6058,N_6083);
or U6913 (N_6913,N_6460,N_6422);
and U6914 (N_6914,N_6475,N_6157);
nor U6915 (N_6915,N_6261,N_6229);
nor U6916 (N_6916,N_6219,N_6229);
or U6917 (N_6917,N_6373,N_6369);
nor U6918 (N_6918,N_6358,N_6380);
nand U6919 (N_6919,N_6254,N_6011);
nand U6920 (N_6920,N_6390,N_6226);
xor U6921 (N_6921,N_6492,N_6450);
xor U6922 (N_6922,N_6458,N_6211);
nand U6923 (N_6923,N_6339,N_6401);
xor U6924 (N_6924,N_6161,N_6164);
and U6925 (N_6925,N_6261,N_6214);
nor U6926 (N_6926,N_6229,N_6283);
and U6927 (N_6927,N_6171,N_6464);
and U6928 (N_6928,N_6299,N_6262);
and U6929 (N_6929,N_6341,N_6176);
and U6930 (N_6930,N_6177,N_6127);
xor U6931 (N_6931,N_6110,N_6396);
and U6932 (N_6932,N_6140,N_6228);
and U6933 (N_6933,N_6177,N_6170);
or U6934 (N_6934,N_6045,N_6189);
nand U6935 (N_6935,N_6245,N_6440);
nor U6936 (N_6936,N_6125,N_6275);
xor U6937 (N_6937,N_6254,N_6055);
and U6938 (N_6938,N_6184,N_6395);
or U6939 (N_6939,N_6251,N_6454);
nor U6940 (N_6940,N_6032,N_6460);
or U6941 (N_6941,N_6173,N_6158);
or U6942 (N_6942,N_6498,N_6302);
or U6943 (N_6943,N_6340,N_6263);
nand U6944 (N_6944,N_6412,N_6329);
and U6945 (N_6945,N_6316,N_6214);
xnor U6946 (N_6946,N_6360,N_6035);
and U6947 (N_6947,N_6465,N_6306);
or U6948 (N_6948,N_6360,N_6157);
xor U6949 (N_6949,N_6177,N_6187);
or U6950 (N_6950,N_6160,N_6271);
nand U6951 (N_6951,N_6073,N_6044);
nand U6952 (N_6952,N_6366,N_6141);
and U6953 (N_6953,N_6222,N_6344);
and U6954 (N_6954,N_6031,N_6116);
and U6955 (N_6955,N_6295,N_6095);
nand U6956 (N_6956,N_6057,N_6357);
nor U6957 (N_6957,N_6341,N_6152);
and U6958 (N_6958,N_6350,N_6139);
nor U6959 (N_6959,N_6258,N_6168);
nor U6960 (N_6960,N_6267,N_6211);
xnor U6961 (N_6961,N_6306,N_6385);
nand U6962 (N_6962,N_6083,N_6349);
xor U6963 (N_6963,N_6189,N_6459);
nor U6964 (N_6964,N_6479,N_6322);
nor U6965 (N_6965,N_6302,N_6288);
nor U6966 (N_6966,N_6409,N_6432);
or U6967 (N_6967,N_6238,N_6379);
xor U6968 (N_6968,N_6092,N_6373);
xor U6969 (N_6969,N_6494,N_6228);
xor U6970 (N_6970,N_6069,N_6255);
nand U6971 (N_6971,N_6034,N_6317);
and U6972 (N_6972,N_6347,N_6138);
xor U6973 (N_6973,N_6402,N_6435);
and U6974 (N_6974,N_6449,N_6483);
nor U6975 (N_6975,N_6145,N_6065);
xnor U6976 (N_6976,N_6203,N_6023);
xor U6977 (N_6977,N_6313,N_6097);
and U6978 (N_6978,N_6005,N_6243);
xor U6979 (N_6979,N_6189,N_6271);
or U6980 (N_6980,N_6208,N_6132);
and U6981 (N_6981,N_6164,N_6465);
nor U6982 (N_6982,N_6057,N_6127);
xor U6983 (N_6983,N_6150,N_6180);
nand U6984 (N_6984,N_6486,N_6148);
and U6985 (N_6985,N_6354,N_6196);
and U6986 (N_6986,N_6139,N_6447);
or U6987 (N_6987,N_6080,N_6257);
nor U6988 (N_6988,N_6265,N_6218);
and U6989 (N_6989,N_6419,N_6079);
nand U6990 (N_6990,N_6471,N_6402);
nand U6991 (N_6991,N_6363,N_6265);
xnor U6992 (N_6992,N_6168,N_6431);
nor U6993 (N_6993,N_6194,N_6124);
or U6994 (N_6994,N_6220,N_6420);
xnor U6995 (N_6995,N_6287,N_6022);
and U6996 (N_6996,N_6436,N_6187);
or U6997 (N_6997,N_6436,N_6046);
nor U6998 (N_6998,N_6449,N_6416);
or U6999 (N_6999,N_6043,N_6388);
nor U7000 (N_7000,N_6642,N_6963);
nand U7001 (N_7001,N_6676,N_6536);
nand U7002 (N_7002,N_6543,N_6955);
nand U7003 (N_7003,N_6881,N_6643);
and U7004 (N_7004,N_6695,N_6786);
nor U7005 (N_7005,N_6895,N_6887);
or U7006 (N_7006,N_6933,N_6912);
xnor U7007 (N_7007,N_6573,N_6645);
and U7008 (N_7008,N_6575,N_6908);
or U7009 (N_7009,N_6918,N_6858);
nor U7010 (N_7010,N_6799,N_6501);
nand U7011 (N_7011,N_6586,N_6898);
and U7012 (N_7012,N_6552,N_6820);
and U7013 (N_7013,N_6865,N_6979);
nor U7014 (N_7014,N_6869,N_6606);
and U7015 (N_7015,N_6698,N_6768);
nor U7016 (N_7016,N_6960,N_6894);
nand U7017 (N_7017,N_6787,N_6623);
nand U7018 (N_7018,N_6861,N_6655);
and U7019 (N_7019,N_6677,N_6774);
xnor U7020 (N_7020,N_6944,N_6562);
and U7021 (N_7021,N_6977,N_6760);
or U7022 (N_7022,N_6605,N_6783);
nor U7023 (N_7023,N_6802,N_6968);
nor U7024 (N_7024,N_6672,N_6974);
xnor U7025 (N_7025,N_6807,N_6632);
nand U7026 (N_7026,N_6539,N_6791);
nand U7027 (N_7027,N_6519,N_6524);
xor U7028 (N_7028,N_6665,N_6907);
nor U7029 (N_7029,N_6884,N_6548);
or U7030 (N_7030,N_6617,N_6981);
or U7031 (N_7031,N_6763,N_6663);
xor U7032 (N_7032,N_6812,N_6965);
xor U7033 (N_7033,N_6806,N_6794);
xnor U7034 (N_7034,N_6888,N_6889);
nor U7035 (N_7035,N_6972,N_6624);
nor U7036 (N_7036,N_6615,N_6694);
nor U7037 (N_7037,N_6725,N_6506);
or U7038 (N_7038,N_6594,N_6722);
nor U7039 (N_7039,N_6830,N_6915);
nor U7040 (N_7040,N_6599,N_6510);
and U7041 (N_7041,N_6701,N_6565);
nand U7042 (N_7042,N_6998,N_6772);
nand U7043 (N_7043,N_6815,N_6983);
nor U7044 (N_7044,N_6756,N_6658);
xnor U7045 (N_7045,N_6638,N_6595);
and U7046 (N_7046,N_6618,N_6603);
xnor U7047 (N_7047,N_6890,N_6538);
nand U7048 (N_7048,N_6800,N_6704);
nand U7049 (N_7049,N_6596,N_6578);
nor U7050 (N_7050,N_6532,N_6954);
and U7051 (N_7051,N_6639,N_6921);
nor U7052 (N_7052,N_6669,N_6734);
and U7053 (N_7053,N_6999,N_6518);
or U7054 (N_7054,N_6987,N_6932);
and U7055 (N_7055,N_6721,N_6724);
xor U7056 (N_7056,N_6937,N_6857);
or U7057 (N_7057,N_6516,N_6929);
or U7058 (N_7058,N_6529,N_6927);
nand U7059 (N_7059,N_6530,N_6626);
and U7060 (N_7060,N_6534,N_6710);
and U7061 (N_7061,N_6950,N_6556);
nand U7062 (N_7062,N_6732,N_6686);
or U7063 (N_7063,N_6607,N_6742);
xor U7064 (N_7064,N_6610,N_6572);
xor U7065 (N_7065,N_6917,N_6608);
nor U7066 (N_7066,N_6664,N_6943);
nand U7067 (N_7067,N_6614,N_6719);
and U7068 (N_7068,N_6587,N_6600);
xor U7069 (N_7069,N_6997,N_6823);
and U7070 (N_7070,N_6592,N_6796);
xor U7071 (N_7071,N_6916,N_6566);
and U7072 (N_7072,N_6754,N_6844);
or U7073 (N_7073,N_6993,N_6941);
nor U7074 (N_7074,N_6708,N_6805);
xnor U7075 (N_7075,N_6711,N_6528);
nor U7076 (N_7076,N_6714,N_6847);
nor U7077 (N_7077,N_6854,N_6577);
xor U7078 (N_7078,N_6690,N_6641);
or U7079 (N_7079,N_6507,N_6718);
and U7080 (N_7080,N_6561,N_6604);
nor U7081 (N_7081,N_6931,N_6938);
xnor U7082 (N_7082,N_6728,N_6836);
nand U7083 (N_7083,N_6588,N_6553);
and U7084 (N_7084,N_6652,N_6750);
nand U7085 (N_7085,N_6852,N_6782);
nand U7086 (N_7086,N_6925,N_6923);
nand U7087 (N_7087,N_6991,N_6970);
nand U7088 (N_7088,N_6909,N_6576);
or U7089 (N_7089,N_6531,N_6511);
nand U7090 (N_7090,N_6737,N_6567);
and U7091 (N_7091,N_6810,N_6976);
nand U7092 (N_7092,N_6648,N_6619);
and U7093 (N_7093,N_6650,N_6770);
or U7094 (N_7094,N_6825,N_6706);
and U7095 (N_7095,N_6814,N_6700);
nand U7096 (N_7096,N_6744,N_6526);
or U7097 (N_7097,N_6570,N_6735);
nor U7098 (N_7098,N_6591,N_6827);
and U7099 (N_7099,N_6637,N_6930);
nor U7100 (N_7100,N_6952,N_6776);
nand U7101 (N_7101,N_6837,N_6855);
nor U7102 (N_7102,N_6731,N_6883);
nand U7103 (N_7103,N_6873,N_6579);
or U7104 (N_7104,N_6853,N_6967);
nand U7105 (N_7105,N_6559,N_6597);
or U7106 (N_7106,N_6792,N_6699);
nand U7107 (N_7107,N_6634,N_6761);
nand U7108 (N_7108,N_6824,N_6514);
nor U7109 (N_7109,N_6947,N_6697);
xor U7110 (N_7110,N_6777,N_6613);
nand U7111 (N_7111,N_6990,N_6903);
nand U7112 (N_7112,N_6753,N_6590);
and U7113 (N_7113,N_6891,N_6920);
nor U7114 (N_7114,N_6752,N_6911);
nor U7115 (N_7115,N_6520,N_6733);
nand U7116 (N_7116,N_6503,N_6517);
or U7117 (N_7117,N_6871,N_6816);
nor U7118 (N_7118,N_6966,N_6549);
nand U7119 (N_7119,N_6957,N_6961);
nand U7120 (N_7120,N_6747,N_6537);
xnor U7121 (N_7121,N_6727,N_6662);
nand U7122 (N_7122,N_6533,N_6877);
nand U7123 (N_7123,N_6829,N_6545);
nor U7124 (N_7124,N_6502,N_6885);
or U7125 (N_7125,N_6771,N_6571);
nor U7126 (N_7126,N_6896,N_6901);
nor U7127 (N_7127,N_6583,N_6715);
and U7128 (N_7128,N_6942,N_6859);
and U7129 (N_7129,N_6584,N_6696);
and U7130 (N_7130,N_6996,N_6525);
or U7131 (N_7131,N_6679,N_6730);
or U7132 (N_7132,N_6654,N_6984);
and U7133 (N_7133,N_6601,N_6843);
and U7134 (N_7134,N_6512,N_6860);
xor U7135 (N_7135,N_6628,N_6897);
nand U7136 (N_7136,N_6946,N_6554);
nand U7137 (N_7137,N_6804,N_6779);
nor U7138 (N_7138,N_6832,N_6817);
nor U7139 (N_7139,N_6759,N_6822);
nand U7140 (N_7140,N_6969,N_6793);
or U7141 (N_7141,N_6555,N_6846);
xnor U7142 (N_7142,N_6707,N_6971);
xor U7143 (N_7143,N_6646,N_6717);
xnor U7144 (N_7144,N_6521,N_6716);
nand U7145 (N_7145,N_6821,N_6673);
and U7146 (N_7146,N_6535,N_6922);
nor U7147 (N_7147,N_6746,N_6789);
xnor U7148 (N_7148,N_6546,N_6809);
or U7149 (N_7149,N_6928,N_6801);
nor U7150 (N_7150,N_6851,N_6982);
xnor U7151 (N_7151,N_6712,N_6948);
and U7152 (N_7152,N_6994,N_6540);
xnor U7153 (N_7153,N_6839,N_6705);
nor U7154 (N_7154,N_6835,N_6616);
and U7155 (N_7155,N_6647,N_6765);
nand U7156 (N_7156,N_6818,N_6940);
and U7157 (N_7157,N_6803,N_6755);
and U7158 (N_7158,N_6563,N_6685);
nand U7159 (N_7159,N_6527,N_6985);
xnor U7160 (N_7160,N_6653,N_6568);
nor U7161 (N_7161,N_6879,N_6790);
xor U7162 (N_7162,N_6681,N_6515);
nand U7163 (N_7163,N_6692,N_6689);
nand U7164 (N_7164,N_6934,N_6989);
nor U7165 (N_7165,N_6778,N_6609);
nor U7166 (N_7166,N_6602,N_6866);
and U7167 (N_7167,N_6541,N_6936);
nand U7168 (N_7168,N_6935,N_6867);
xnor U7169 (N_7169,N_6878,N_6951);
xor U7170 (N_7170,N_6956,N_6767);
or U7171 (N_7171,N_6644,N_6551);
nand U7172 (N_7172,N_6547,N_6995);
nand U7173 (N_7173,N_6621,N_6876);
or U7174 (N_7174,N_6964,N_6649);
xor U7175 (N_7175,N_6508,N_6899);
nor U7176 (N_7176,N_6880,N_6550);
nor U7177 (N_7177,N_6975,N_6682);
nand U7178 (N_7178,N_6666,N_6739);
or U7179 (N_7179,N_6622,N_6640);
nand U7180 (N_7180,N_6688,N_6900);
xnor U7181 (N_7181,N_6625,N_6862);
xor U7182 (N_7182,N_6986,N_6741);
and U7183 (N_7183,N_6906,N_6726);
and U7184 (N_7184,N_6992,N_6833);
nand U7185 (N_7185,N_6939,N_6838);
or U7186 (N_7186,N_6914,N_6775);
nor U7187 (N_7187,N_6749,N_6523);
or U7188 (N_7188,N_6978,N_6636);
or U7189 (N_7189,N_6740,N_6840);
nand U7190 (N_7190,N_6560,N_6808);
and U7191 (N_7191,N_6945,N_6748);
nand U7192 (N_7192,N_6635,N_6798);
nor U7193 (N_7193,N_6558,N_6850);
nor U7194 (N_7194,N_6893,N_6574);
nand U7195 (N_7195,N_6667,N_6769);
nor U7196 (N_7196,N_6743,N_6926);
nor U7197 (N_7197,N_6611,N_6720);
xnor U7198 (N_7198,N_6904,N_6848);
or U7199 (N_7199,N_6842,N_6905);
or U7200 (N_7200,N_6589,N_6882);
nand U7201 (N_7201,N_6845,N_6849);
nand U7202 (N_7202,N_6819,N_6738);
nand U7203 (N_7203,N_6693,N_6831);
and U7204 (N_7204,N_6736,N_6766);
nand U7205 (N_7205,N_6509,N_6569);
or U7206 (N_7206,N_6962,N_6863);
xor U7207 (N_7207,N_6745,N_6627);
nor U7208 (N_7208,N_6780,N_6902);
nand U7209 (N_7209,N_6886,N_6557);
and U7210 (N_7210,N_6670,N_6811);
nor U7211 (N_7211,N_6703,N_6834);
nor U7212 (N_7212,N_6729,N_6683);
xnor U7213 (N_7213,N_6651,N_6702);
xnor U7214 (N_7214,N_6762,N_6633);
xor U7215 (N_7215,N_6875,N_6630);
xor U7216 (N_7216,N_6504,N_6631);
xnor U7217 (N_7217,N_6910,N_6675);
and U7218 (N_7218,N_6542,N_6585);
xor U7219 (N_7219,N_6564,N_6856);
xnor U7220 (N_7220,N_6713,N_6892);
xor U7221 (N_7221,N_6656,N_6620);
or U7222 (N_7222,N_6687,N_6788);
xor U7223 (N_7223,N_6784,N_6659);
or U7224 (N_7224,N_6513,N_6522);
nor U7225 (N_7225,N_6924,N_6773);
nand U7226 (N_7226,N_6913,N_6500);
nand U7227 (N_7227,N_6751,N_6668);
and U7228 (N_7228,N_6505,N_6764);
and U7229 (N_7229,N_6797,N_6758);
or U7230 (N_7230,N_6973,N_6868);
nor U7231 (N_7231,N_6581,N_6629);
and U7232 (N_7232,N_6795,N_6612);
and U7233 (N_7233,N_6691,N_6813);
nand U7234 (N_7234,N_6680,N_6580);
nand U7235 (N_7235,N_6872,N_6674);
nand U7236 (N_7236,N_6671,N_6781);
or U7237 (N_7237,N_6723,N_6919);
or U7238 (N_7238,N_6864,N_6988);
xor U7239 (N_7239,N_6661,N_6757);
or U7240 (N_7240,N_6657,N_6709);
or U7241 (N_7241,N_6582,N_6874);
and U7242 (N_7242,N_6593,N_6841);
nand U7243 (N_7243,N_6959,N_6684);
xor U7244 (N_7244,N_6870,N_6678);
nor U7245 (N_7245,N_6828,N_6598);
nor U7246 (N_7246,N_6544,N_6826);
and U7247 (N_7247,N_6958,N_6980);
and U7248 (N_7248,N_6660,N_6785);
xor U7249 (N_7249,N_6949,N_6953);
nand U7250 (N_7250,N_6950,N_6614);
or U7251 (N_7251,N_6884,N_6711);
and U7252 (N_7252,N_6920,N_6710);
nand U7253 (N_7253,N_6765,N_6930);
nand U7254 (N_7254,N_6603,N_6799);
xor U7255 (N_7255,N_6837,N_6832);
or U7256 (N_7256,N_6899,N_6777);
xor U7257 (N_7257,N_6622,N_6892);
nor U7258 (N_7258,N_6701,N_6530);
or U7259 (N_7259,N_6998,N_6901);
and U7260 (N_7260,N_6892,N_6608);
and U7261 (N_7261,N_6700,N_6639);
nand U7262 (N_7262,N_6922,N_6948);
or U7263 (N_7263,N_6600,N_6510);
nor U7264 (N_7264,N_6637,N_6647);
or U7265 (N_7265,N_6938,N_6876);
xor U7266 (N_7266,N_6977,N_6711);
xnor U7267 (N_7267,N_6765,N_6881);
nor U7268 (N_7268,N_6526,N_6603);
xnor U7269 (N_7269,N_6620,N_6985);
nand U7270 (N_7270,N_6923,N_6580);
or U7271 (N_7271,N_6733,N_6701);
or U7272 (N_7272,N_6597,N_6576);
xor U7273 (N_7273,N_6939,N_6850);
xnor U7274 (N_7274,N_6642,N_6566);
nor U7275 (N_7275,N_6513,N_6674);
and U7276 (N_7276,N_6906,N_6510);
xor U7277 (N_7277,N_6670,N_6776);
nand U7278 (N_7278,N_6864,N_6807);
xnor U7279 (N_7279,N_6773,N_6596);
or U7280 (N_7280,N_6903,N_6563);
and U7281 (N_7281,N_6646,N_6749);
or U7282 (N_7282,N_6923,N_6871);
xor U7283 (N_7283,N_6506,N_6717);
nor U7284 (N_7284,N_6883,N_6667);
nor U7285 (N_7285,N_6878,N_6502);
or U7286 (N_7286,N_6639,N_6575);
or U7287 (N_7287,N_6683,N_6959);
nand U7288 (N_7288,N_6778,N_6526);
and U7289 (N_7289,N_6528,N_6613);
and U7290 (N_7290,N_6519,N_6538);
xor U7291 (N_7291,N_6968,N_6550);
xnor U7292 (N_7292,N_6948,N_6805);
and U7293 (N_7293,N_6747,N_6772);
nand U7294 (N_7294,N_6869,N_6754);
or U7295 (N_7295,N_6518,N_6923);
xor U7296 (N_7296,N_6915,N_6552);
nand U7297 (N_7297,N_6887,N_6530);
xor U7298 (N_7298,N_6604,N_6567);
nor U7299 (N_7299,N_6747,N_6722);
and U7300 (N_7300,N_6731,N_6913);
xnor U7301 (N_7301,N_6586,N_6529);
or U7302 (N_7302,N_6874,N_6588);
nand U7303 (N_7303,N_6695,N_6906);
nor U7304 (N_7304,N_6834,N_6511);
nor U7305 (N_7305,N_6749,N_6803);
nor U7306 (N_7306,N_6801,N_6635);
nand U7307 (N_7307,N_6956,N_6715);
nand U7308 (N_7308,N_6773,N_6981);
nand U7309 (N_7309,N_6991,N_6605);
and U7310 (N_7310,N_6691,N_6736);
nor U7311 (N_7311,N_6542,N_6620);
and U7312 (N_7312,N_6505,N_6512);
and U7313 (N_7313,N_6739,N_6935);
nand U7314 (N_7314,N_6702,N_6992);
nand U7315 (N_7315,N_6587,N_6772);
or U7316 (N_7316,N_6558,N_6537);
and U7317 (N_7317,N_6552,N_6804);
nor U7318 (N_7318,N_6869,N_6749);
nor U7319 (N_7319,N_6763,N_6931);
nand U7320 (N_7320,N_6859,N_6722);
nor U7321 (N_7321,N_6530,N_6801);
nor U7322 (N_7322,N_6615,N_6786);
or U7323 (N_7323,N_6586,N_6583);
and U7324 (N_7324,N_6817,N_6968);
xor U7325 (N_7325,N_6624,N_6507);
xor U7326 (N_7326,N_6602,N_6865);
and U7327 (N_7327,N_6584,N_6564);
nor U7328 (N_7328,N_6694,N_6865);
nor U7329 (N_7329,N_6868,N_6863);
nand U7330 (N_7330,N_6566,N_6896);
xor U7331 (N_7331,N_6742,N_6612);
nor U7332 (N_7332,N_6534,N_6700);
and U7333 (N_7333,N_6654,N_6678);
and U7334 (N_7334,N_6579,N_6810);
nand U7335 (N_7335,N_6595,N_6960);
or U7336 (N_7336,N_6615,N_6749);
xnor U7337 (N_7337,N_6568,N_6947);
nor U7338 (N_7338,N_6613,N_6641);
or U7339 (N_7339,N_6894,N_6964);
nand U7340 (N_7340,N_6648,N_6843);
xnor U7341 (N_7341,N_6996,N_6772);
xnor U7342 (N_7342,N_6896,N_6613);
nand U7343 (N_7343,N_6643,N_6552);
xor U7344 (N_7344,N_6727,N_6887);
nand U7345 (N_7345,N_6948,N_6834);
xor U7346 (N_7346,N_6654,N_6627);
nand U7347 (N_7347,N_6798,N_6547);
nand U7348 (N_7348,N_6723,N_6543);
and U7349 (N_7349,N_6574,N_6712);
and U7350 (N_7350,N_6522,N_6781);
nand U7351 (N_7351,N_6793,N_6594);
or U7352 (N_7352,N_6710,N_6654);
nand U7353 (N_7353,N_6880,N_6545);
nand U7354 (N_7354,N_6659,N_6755);
nand U7355 (N_7355,N_6866,N_6667);
and U7356 (N_7356,N_6756,N_6719);
and U7357 (N_7357,N_6982,N_6899);
or U7358 (N_7358,N_6744,N_6912);
nor U7359 (N_7359,N_6892,N_6912);
and U7360 (N_7360,N_6705,N_6639);
nor U7361 (N_7361,N_6832,N_6733);
or U7362 (N_7362,N_6639,N_6685);
nor U7363 (N_7363,N_6790,N_6777);
nor U7364 (N_7364,N_6886,N_6574);
or U7365 (N_7365,N_6969,N_6771);
nand U7366 (N_7366,N_6891,N_6807);
and U7367 (N_7367,N_6925,N_6788);
nor U7368 (N_7368,N_6706,N_6816);
nand U7369 (N_7369,N_6568,N_6869);
xnor U7370 (N_7370,N_6760,N_6840);
nand U7371 (N_7371,N_6703,N_6747);
nand U7372 (N_7372,N_6539,N_6841);
or U7373 (N_7373,N_6514,N_6685);
and U7374 (N_7374,N_6709,N_6690);
and U7375 (N_7375,N_6980,N_6969);
nand U7376 (N_7376,N_6718,N_6853);
and U7377 (N_7377,N_6740,N_6694);
xnor U7378 (N_7378,N_6794,N_6721);
nor U7379 (N_7379,N_6601,N_6930);
and U7380 (N_7380,N_6592,N_6702);
xnor U7381 (N_7381,N_6876,N_6886);
nor U7382 (N_7382,N_6589,N_6971);
and U7383 (N_7383,N_6829,N_6524);
xnor U7384 (N_7384,N_6596,N_6763);
nor U7385 (N_7385,N_6818,N_6857);
nor U7386 (N_7386,N_6812,N_6646);
or U7387 (N_7387,N_6893,N_6817);
and U7388 (N_7388,N_6767,N_6515);
nor U7389 (N_7389,N_6529,N_6870);
and U7390 (N_7390,N_6564,N_6828);
nor U7391 (N_7391,N_6784,N_6948);
or U7392 (N_7392,N_6830,N_6709);
nand U7393 (N_7393,N_6592,N_6525);
nand U7394 (N_7394,N_6708,N_6589);
xnor U7395 (N_7395,N_6637,N_6737);
xor U7396 (N_7396,N_6860,N_6671);
or U7397 (N_7397,N_6550,N_6879);
or U7398 (N_7398,N_6993,N_6860);
or U7399 (N_7399,N_6863,N_6589);
nand U7400 (N_7400,N_6522,N_6983);
or U7401 (N_7401,N_6534,N_6589);
nor U7402 (N_7402,N_6649,N_6944);
and U7403 (N_7403,N_6632,N_6847);
and U7404 (N_7404,N_6730,N_6966);
nand U7405 (N_7405,N_6776,N_6947);
or U7406 (N_7406,N_6689,N_6788);
nand U7407 (N_7407,N_6518,N_6714);
and U7408 (N_7408,N_6779,N_6902);
nor U7409 (N_7409,N_6831,N_6858);
nor U7410 (N_7410,N_6565,N_6537);
and U7411 (N_7411,N_6805,N_6651);
nand U7412 (N_7412,N_6893,N_6538);
and U7413 (N_7413,N_6896,N_6858);
or U7414 (N_7414,N_6973,N_6943);
and U7415 (N_7415,N_6590,N_6796);
or U7416 (N_7416,N_6675,N_6920);
and U7417 (N_7417,N_6670,N_6707);
nand U7418 (N_7418,N_6767,N_6660);
or U7419 (N_7419,N_6800,N_6735);
and U7420 (N_7420,N_6506,N_6513);
xor U7421 (N_7421,N_6762,N_6944);
or U7422 (N_7422,N_6932,N_6539);
and U7423 (N_7423,N_6696,N_6659);
xnor U7424 (N_7424,N_6926,N_6763);
or U7425 (N_7425,N_6672,N_6548);
nor U7426 (N_7426,N_6557,N_6813);
nand U7427 (N_7427,N_6696,N_6902);
nor U7428 (N_7428,N_6554,N_6976);
or U7429 (N_7429,N_6900,N_6701);
or U7430 (N_7430,N_6826,N_6768);
or U7431 (N_7431,N_6553,N_6570);
nor U7432 (N_7432,N_6925,N_6779);
and U7433 (N_7433,N_6693,N_6943);
xnor U7434 (N_7434,N_6764,N_6551);
or U7435 (N_7435,N_6734,N_6717);
nor U7436 (N_7436,N_6700,N_6659);
nor U7437 (N_7437,N_6800,N_6597);
xor U7438 (N_7438,N_6966,N_6604);
xnor U7439 (N_7439,N_6985,N_6927);
nand U7440 (N_7440,N_6940,N_6547);
nand U7441 (N_7441,N_6631,N_6621);
xnor U7442 (N_7442,N_6950,N_6540);
and U7443 (N_7443,N_6702,N_6718);
xnor U7444 (N_7444,N_6852,N_6611);
and U7445 (N_7445,N_6717,N_6568);
nand U7446 (N_7446,N_6599,N_6855);
nand U7447 (N_7447,N_6829,N_6701);
nand U7448 (N_7448,N_6945,N_6759);
and U7449 (N_7449,N_6871,N_6578);
nor U7450 (N_7450,N_6605,N_6643);
nor U7451 (N_7451,N_6501,N_6990);
nand U7452 (N_7452,N_6705,N_6514);
nand U7453 (N_7453,N_6999,N_6730);
xnor U7454 (N_7454,N_6853,N_6893);
or U7455 (N_7455,N_6792,N_6530);
nand U7456 (N_7456,N_6702,N_6893);
nand U7457 (N_7457,N_6996,N_6800);
xor U7458 (N_7458,N_6979,N_6688);
nor U7459 (N_7459,N_6716,N_6909);
or U7460 (N_7460,N_6669,N_6832);
nor U7461 (N_7461,N_6602,N_6605);
xor U7462 (N_7462,N_6661,N_6977);
nand U7463 (N_7463,N_6919,N_6957);
or U7464 (N_7464,N_6563,N_6949);
nand U7465 (N_7465,N_6888,N_6565);
nand U7466 (N_7466,N_6557,N_6795);
xor U7467 (N_7467,N_6969,N_6924);
and U7468 (N_7468,N_6766,N_6792);
nor U7469 (N_7469,N_6593,N_6601);
or U7470 (N_7470,N_6740,N_6950);
nand U7471 (N_7471,N_6591,N_6718);
nand U7472 (N_7472,N_6945,N_6951);
nor U7473 (N_7473,N_6686,N_6929);
and U7474 (N_7474,N_6707,N_6571);
xor U7475 (N_7475,N_6865,N_6930);
xnor U7476 (N_7476,N_6691,N_6793);
or U7477 (N_7477,N_6801,N_6720);
and U7478 (N_7478,N_6518,N_6848);
nand U7479 (N_7479,N_6929,N_6527);
nor U7480 (N_7480,N_6741,N_6629);
and U7481 (N_7481,N_6591,N_6866);
xnor U7482 (N_7482,N_6602,N_6523);
nand U7483 (N_7483,N_6704,N_6606);
nor U7484 (N_7484,N_6642,N_6735);
nor U7485 (N_7485,N_6750,N_6850);
xnor U7486 (N_7486,N_6896,N_6925);
nor U7487 (N_7487,N_6687,N_6703);
nand U7488 (N_7488,N_6824,N_6532);
and U7489 (N_7489,N_6677,N_6686);
nand U7490 (N_7490,N_6650,N_6708);
nand U7491 (N_7491,N_6618,N_6826);
xor U7492 (N_7492,N_6621,N_6808);
and U7493 (N_7493,N_6698,N_6759);
nor U7494 (N_7494,N_6530,N_6503);
or U7495 (N_7495,N_6945,N_6632);
xnor U7496 (N_7496,N_6983,N_6596);
nand U7497 (N_7497,N_6584,N_6828);
nand U7498 (N_7498,N_6669,N_6600);
xor U7499 (N_7499,N_6882,N_6673);
or U7500 (N_7500,N_7288,N_7001);
xnor U7501 (N_7501,N_7172,N_7460);
and U7502 (N_7502,N_7209,N_7355);
nand U7503 (N_7503,N_7370,N_7032);
xor U7504 (N_7504,N_7093,N_7264);
nand U7505 (N_7505,N_7280,N_7246);
and U7506 (N_7506,N_7396,N_7429);
xnor U7507 (N_7507,N_7114,N_7217);
and U7508 (N_7508,N_7241,N_7420);
nor U7509 (N_7509,N_7210,N_7405);
or U7510 (N_7510,N_7021,N_7358);
xor U7511 (N_7511,N_7281,N_7235);
and U7512 (N_7512,N_7224,N_7380);
xor U7513 (N_7513,N_7256,N_7274);
and U7514 (N_7514,N_7293,N_7208);
nor U7515 (N_7515,N_7439,N_7020);
nor U7516 (N_7516,N_7386,N_7453);
nand U7517 (N_7517,N_7059,N_7259);
and U7518 (N_7518,N_7363,N_7492);
nand U7519 (N_7519,N_7286,N_7427);
xnor U7520 (N_7520,N_7227,N_7393);
or U7521 (N_7521,N_7130,N_7174);
nand U7522 (N_7522,N_7195,N_7468);
nor U7523 (N_7523,N_7131,N_7069);
and U7524 (N_7524,N_7212,N_7335);
xnor U7525 (N_7525,N_7449,N_7013);
and U7526 (N_7526,N_7411,N_7399);
nand U7527 (N_7527,N_7015,N_7373);
nor U7528 (N_7528,N_7138,N_7162);
and U7529 (N_7529,N_7478,N_7082);
nor U7530 (N_7530,N_7310,N_7118);
nand U7531 (N_7531,N_7400,N_7487);
or U7532 (N_7532,N_7051,N_7379);
or U7533 (N_7533,N_7446,N_7056);
and U7534 (N_7534,N_7495,N_7490);
or U7535 (N_7535,N_7254,N_7315);
or U7536 (N_7536,N_7119,N_7002);
xnor U7537 (N_7537,N_7035,N_7479);
nand U7538 (N_7538,N_7070,N_7282);
nand U7539 (N_7539,N_7270,N_7340);
xor U7540 (N_7540,N_7458,N_7301);
or U7541 (N_7541,N_7213,N_7475);
nor U7542 (N_7542,N_7110,N_7216);
nand U7543 (N_7543,N_7333,N_7247);
xnor U7544 (N_7544,N_7237,N_7409);
nand U7545 (N_7545,N_7451,N_7322);
or U7546 (N_7546,N_7108,N_7101);
or U7547 (N_7547,N_7024,N_7023);
and U7548 (N_7548,N_7145,N_7090);
xnor U7549 (N_7549,N_7161,N_7248);
or U7550 (N_7550,N_7218,N_7179);
nor U7551 (N_7551,N_7499,N_7206);
and U7552 (N_7552,N_7245,N_7250);
and U7553 (N_7553,N_7125,N_7403);
or U7554 (N_7554,N_7025,N_7154);
xnor U7555 (N_7555,N_7215,N_7252);
and U7556 (N_7556,N_7463,N_7151);
nand U7557 (N_7557,N_7238,N_7207);
and U7558 (N_7558,N_7229,N_7220);
xor U7559 (N_7559,N_7311,N_7223);
xnor U7560 (N_7560,N_7075,N_7387);
or U7561 (N_7561,N_7324,N_7257);
or U7562 (N_7562,N_7494,N_7077);
or U7563 (N_7563,N_7361,N_7074);
and U7564 (N_7564,N_7291,N_7294);
and U7565 (N_7565,N_7395,N_7197);
or U7566 (N_7566,N_7042,N_7159);
nand U7567 (N_7567,N_7203,N_7349);
nor U7568 (N_7568,N_7033,N_7292);
or U7569 (N_7569,N_7312,N_7022);
nand U7570 (N_7570,N_7255,N_7419);
nor U7571 (N_7571,N_7234,N_7461);
or U7572 (N_7572,N_7413,N_7457);
or U7573 (N_7573,N_7408,N_7342);
nor U7574 (N_7574,N_7450,N_7103);
and U7575 (N_7575,N_7092,N_7422);
or U7576 (N_7576,N_7120,N_7474);
xnor U7577 (N_7577,N_7417,N_7144);
or U7578 (N_7578,N_7117,N_7231);
xnor U7579 (N_7579,N_7378,N_7276);
nand U7580 (N_7580,N_7006,N_7049);
or U7581 (N_7581,N_7389,N_7230);
or U7582 (N_7582,N_7438,N_7171);
or U7583 (N_7583,N_7320,N_7236);
or U7584 (N_7584,N_7390,N_7347);
nor U7585 (N_7585,N_7076,N_7260);
and U7586 (N_7586,N_7432,N_7484);
xor U7587 (N_7587,N_7155,N_7316);
nor U7588 (N_7588,N_7477,N_7476);
nand U7589 (N_7589,N_7410,N_7081);
nor U7590 (N_7590,N_7200,N_7201);
nand U7591 (N_7591,N_7214,N_7331);
and U7592 (N_7592,N_7242,N_7462);
and U7593 (N_7593,N_7455,N_7191);
xnor U7594 (N_7594,N_7375,N_7034);
and U7595 (N_7595,N_7123,N_7030);
and U7596 (N_7596,N_7038,N_7431);
nor U7597 (N_7597,N_7019,N_7481);
or U7598 (N_7598,N_7482,N_7228);
nand U7599 (N_7599,N_7163,N_7416);
nor U7600 (N_7600,N_7415,N_7087);
or U7601 (N_7601,N_7485,N_7078);
nand U7602 (N_7602,N_7444,N_7364);
nand U7603 (N_7603,N_7440,N_7266);
nor U7604 (N_7604,N_7135,N_7047);
nand U7605 (N_7605,N_7066,N_7426);
and U7606 (N_7606,N_7044,N_7425);
and U7607 (N_7607,N_7423,N_7263);
or U7608 (N_7608,N_7096,N_7351);
or U7609 (N_7609,N_7299,N_7164);
and U7610 (N_7610,N_7048,N_7326);
and U7611 (N_7611,N_7243,N_7459);
nand U7612 (N_7612,N_7268,N_7063);
xor U7613 (N_7613,N_7313,N_7343);
nand U7614 (N_7614,N_7057,N_7088);
and U7615 (N_7615,N_7008,N_7412);
or U7616 (N_7616,N_7177,N_7065);
xnor U7617 (N_7617,N_7337,N_7004);
nand U7618 (N_7618,N_7339,N_7404);
or U7619 (N_7619,N_7128,N_7445);
nor U7620 (N_7620,N_7436,N_7061);
xor U7621 (N_7621,N_7398,N_7045);
nand U7622 (N_7622,N_7287,N_7308);
xor U7623 (N_7623,N_7132,N_7198);
nand U7624 (N_7624,N_7165,N_7356);
or U7625 (N_7625,N_7369,N_7433);
nor U7626 (N_7626,N_7041,N_7367);
or U7627 (N_7627,N_7107,N_7284);
xor U7628 (N_7628,N_7084,N_7302);
or U7629 (N_7629,N_7491,N_7289);
and U7630 (N_7630,N_7493,N_7202);
nor U7631 (N_7631,N_7384,N_7007);
nor U7632 (N_7632,N_7300,N_7376);
xnor U7633 (N_7633,N_7095,N_7028);
or U7634 (N_7634,N_7105,N_7112);
nand U7635 (N_7635,N_7014,N_7297);
nand U7636 (N_7636,N_7321,N_7486);
nand U7637 (N_7637,N_7498,N_7170);
or U7638 (N_7638,N_7072,N_7193);
xnor U7639 (N_7639,N_7158,N_7497);
xor U7640 (N_7640,N_7178,N_7157);
and U7641 (N_7641,N_7345,N_7346);
xnor U7642 (N_7642,N_7186,N_7012);
xor U7643 (N_7643,N_7183,N_7290);
and U7644 (N_7644,N_7083,N_7388);
or U7645 (N_7645,N_7421,N_7106);
or U7646 (N_7646,N_7122,N_7225);
or U7647 (N_7647,N_7189,N_7332);
and U7648 (N_7648,N_7141,N_7139);
or U7649 (N_7649,N_7382,N_7187);
and U7650 (N_7650,N_7113,N_7050);
or U7651 (N_7651,N_7115,N_7488);
or U7652 (N_7652,N_7273,N_7173);
and U7653 (N_7653,N_7317,N_7226);
nand U7654 (N_7654,N_7116,N_7053);
xnor U7655 (N_7655,N_7272,N_7153);
nor U7656 (N_7656,N_7418,N_7064);
nand U7657 (N_7657,N_7442,N_7329);
or U7658 (N_7658,N_7239,N_7129);
or U7659 (N_7659,N_7039,N_7185);
xor U7660 (N_7660,N_7085,N_7447);
or U7661 (N_7661,N_7244,N_7043);
nand U7662 (N_7662,N_7037,N_7307);
xor U7663 (N_7663,N_7348,N_7296);
nor U7664 (N_7664,N_7192,N_7441);
or U7665 (N_7665,N_7430,N_7111);
xor U7666 (N_7666,N_7464,N_7146);
or U7667 (N_7667,N_7143,N_7222);
xor U7668 (N_7668,N_7211,N_7062);
or U7669 (N_7669,N_7334,N_7055);
and U7670 (N_7670,N_7327,N_7283);
or U7671 (N_7671,N_7149,N_7167);
nand U7672 (N_7672,N_7052,N_7277);
xor U7673 (N_7673,N_7469,N_7434);
and U7674 (N_7674,N_7309,N_7018);
nand U7675 (N_7675,N_7303,N_7233);
or U7676 (N_7676,N_7219,N_7199);
and U7677 (N_7677,N_7029,N_7104);
xor U7678 (N_7678,N_7134,N_7181);
or U7679 (N_7679,N_7323,N_7188);
xor U7680 (N_7680,N_7168,N_7190);
xor U7681 (N_7681,N_7344,N_7318);
xor U7682 (N_7682,N_7005,N_7150);
nor U7683 (N_7683,N_7182,N_7091);
or U7684 (N_7684,N_7362,N_7046);
and U7685 (N_7685,N_7269,N_7319);
and U7686 (N_7686,N_7133,N_7080);
xor U7687 (N_7687,N_7397,N_7454);
or U7688 (N_7688,N_7278,N_7184);
and U7689 (N_7689,N_7466,N_7295);
nand U7690 (N_7690,N_7058,N_7251);
or U7691 (N_7691,N_7341,N_7194);
nand U7692 (N_7692,N_7160,N_7054);
and U7693 (N_7693,N_7325,N_7240);
or U7694 (N_7694,N_7169,N_7456);
nor U7695 (N_7695,N_7094,N_7371);
xor U7696 (N_7696,N_7465,N_7428);
nor U7697 (N_7697,N_7489,N_7031);
xor U7698 (N_7698,N_7306,N_7142);
nand U7699 (N_7699,N_7424,N_7435);
and U7700 (N_7700,N_7180,N_7067);
xor U7701 (N_7701,N_7480,N_7279);
and U7702 (N_7702,N_7406,N_7175);
or U7703 (N_7703,N_7330,N_7102);
nand U7704 (N_7704,N_7009,N_7097);
xnor U7705 (N_7705,N_7147,N_7353);
and U7706 (N_7706,N_7261,N_7467);
nand U7707 (N_7707,N_7140,N_7121);
or U7708 (N_7708,N_7402,N_7026);
and U7709 (N_7709,N_7359,N_7285);
and U7710 (N_7710,N_7368,N_7099);
or U7711 (N_7711,N_7068,N_7338);
and U7712 (N_7712,N_7221,N_7360);
and U7713 (N_7713,N_7124,N_7016);
nor U7714 (N_7714,N_7437,N_7414);
or U7715 (N_7715,N_7071,N_7152);
xor U7716 (N_7716,N_7253,N_7471);
or U7717 (N_7717,N_7452,N_7298);
and U7718 (N_7718,N_7328,N_7472);
nor U7719 (N_7719,N_7401,N_7470);
nand U7720 (N_7720,N_7496,N_7365);
or U7721 (N_7721,N_7377,N_7205);
and U7722 (N_7722,N_7448,N_7100);
xor U7723 (N_7723,N_7204,N_7109);
or U7724 (N_7724,N_7262,N_7258);
xor U7725 (N_7725,N_7267,N_7086);
nor U7726 (N_7726,N_7148,N_7060);
nor U7727 (N_7727,N_7372,N_7089);
nand U7728 (N_7728,N_7232,N_7079);
or U7729 (N_7729,N_7304,N_7381);
and U7730 (N_7730,N_7443,N_7483);
xor U7731 (N_7731,N_7036,N_7196);
xnor U7732 (N_7732,N_7383,N_7350);
and U7733 (N_7733,N_7000,N_7040);
nor U7734 (N_7734,N_7366,N_7003);
xor U7735 (N_7735,N_7473,N_7126);
and U7736 (N_7736,N_7305,N_7166);
nand U7737 (N_7737,N_7336,N_7073);
xor U7738 (N_7738,N_7394,N_7275);
or U7739 (N_7739,N_7249,N_7385);
and U7740 (N_7740,N_7314,N_7017);
nor U7741 (N_7741,N_7010,N_7407);
or U7742 (N_7742,N_7357,N_7176);
and U7743 (N_7743,N_7352,N_7127);
nor U7744 (N_7744,N_7011,N_7391);
nand U7745 (N_7745,N_7271,N_7374);
nor U7746 (N_7746,N_7156,N_7136);
nand U7747 (N_7747,N_7137,N_7265);
nor U7748 (N_7748,N_7392,N_7354);
nand U7749 (N_7749,N_7098,N_7027);
xnor U7750 (N_7750,N_7239,N_7177);
nand U7751 (N_7751,N_7480,N_7010);
xnor U7752 (N_7752,N_7393,N_7275);
nor U7753 (N_7753,N_7414,N_7446);
nand U7754 (N_7754,N_7236,N_7080);
nand U7755 (N_7755,N_7369,N_7177);
or U7756 (N_7756,N_7395,N_7250);
and U7757 (N_7757,N_7414,N_7040);
or U7758 (N_7758,N_7097,N_7347);
nand U7759 (N_7759,N_7374,N_7413);
nand U7760 (N_7760,N_7220,N_7005);
xnor U7761 (N_7761,N_7333,N_7487);
xor U7762 (N_7762,N_7394,N_7187);
nand U7763 (N_7763,N_7350,N_7492);
and U7764 (N_7764,N_7388,N_7046);
nand U7765 (N_7765,N_7355,N_7429);
nand U7766 (N_7766,N_7335,N_7246);
nor U7767 (N_7767,N_7369,N_7001);
nor U7768 (N_7768,N_7065,N_7075);
xnor U7769 (N_7769,N_7343,N_7009);
xor U7770 (N_7770,N_7407,N_7276);
nor U7771 (N_7771,N_7034,N_7383);
or U7772 (N_7772,N_7277,N_7348);
nor U7773 (N_7773,N_7135,N_7046);
or U7774 (N_7774,N_7392,N_7118);
nand U7775 (N_7775,N_7174,N_7222);
or U7776 (N_7776,N_7182,N_7469);
and U7777 (N_7777,N_7294,N_7071);
and U7778 (N_7778,N_7117,N_7241);
or U7779 (N_7779,N_7162,N_7282);
nor U7780 (N_7780,N_7204,N_7224);
xnor U7781 (N_7781,N_7387,N_7008);
or U7782 (N_7782,N_7068,N_7257);
and U7783 (N_7783,N_7091,N_7122);
nor U7784 (N_7784,N_7228,N_7119);
nor U7785 (N_7785,N_7085,N_7419);
or U7786 (N_7786,N_7380,N_7373);
xor U7787 (N_7787,N_7041,N_7115);
xnor U7788 (N_7788,N_7063,N_7291);
xnor U7789 (N_7789,N_7375,N_7363);
nand U7790 (N_7790,N_7313,N_7036);
or U7791 (N_7791,N_7390,N_7283);
and U7792 (N_7792,N_7171,N_7126);
xor U7793 (N_7793,N_7260,N_7360);
nor U7794 (N_7794,N_7227,N_7065);
or U7795 (N_7795,N_7258,N_7478);
and U7796 (N_7796,N_7252,N_7396);
xnor U7797 (N_7797,N_7234,N_7332);
xnor U7798 (N_7798,N_7337,N_7287);
and U7799 (N_7799,N_7041,N_7338);
or U7800 (N_7800,N_7444,N_7313);
or U7801 (N_7801,N_7244,N_7474);
xnor U7802 (N_7802,N_7344,N_7314);
and U7803 (N_7803,N_7159,N_7403);
nand U7804 (N_7804,N_7091,N_7068);
nor U7805 (N_7805,N_7217,N_7141);
xnor U7806 (N_7806,N_7233,N_7159);
or U7807 (N_7807,N_7072,N_7460);
nand U7808 (N_7808,N_7294,N_7293);
or U7809 (N_7809,N_7055,N_7488);
or U7810 (N_7810,N_7256,N_7271);
xnor U7811 (N_7811,N_7459,N_7338);
nand U7812 (N_7812,N_7003,N_7247);
or U7813 (N_7813,N_7248,N_7166);
xor U7814 (N_7814,N_7144,N_7148);
and U7815 (N_7815,N_7461,N_7121);
or U7816 (N_7816,N_7053,N_7150);
and U7817 (N_7817,N_7182,N_7256);
nor U7818 (N_7818,N_7068,N_7130);
or U7819 (N_7819,N_7206,N_7272);
and U7820 (N_7820,N_7497,N_7293);
nor U7821 (N_7821,N_7261,N_7459);
nor U7822 (N_7822,N_7174,N_7301);
and U7823 (N_7823,N_7312,N_7368);
or U7824 (N_7824,N_7062,N_7240);
or U7825 (N_7825,N_7233,N_7136);
or U7826 (N_7826,N_7293,N_7283);
nand U7827 (N_7827,N_7294,N_7156);
and U7828 (N_7828,N_7472,N_7027);
nand U7829 (N_7829,N_7419,N_7070);
nor U7830 (N_7830,N_7194,N_7044);
or U7831 (N_7831,N_7245,N_7184);
nand U7832 (N_7832,N_7331,N_7187);
or U7833 (N_7833,N_7307,N_7405);
and U7834 (N_7834,N_7341,N_7237);
nand U7835 (N_7835,N_7370,N_7314);
and U7836 (N_7836,N_7217,N_7109);
and U7837 (N_7837,N_7471,N_7464);
xnor U7838 (N_7838,N_7465,N_7146);
nor U7839 (N_7839,N_7334,N_7185);
and U7840 (N_7840,N_7353,N_7405);
or U7841 (N_7841,N_7227,N_7079);
nor U7842 (N_7842,N_7107,N_7199);
nand U7843 (N_7843,N_7020,N_7413);
xor U7844 (N_7844,N_7205,N_7197);
nand U7845 (N_7845,N_7079,N_7013);
and U7846 (N_7846,N_7237,N_7022);
xnor U7847 (N_7847,N_7436,N_7025);
or U7848 (N_7848,N_7186,N_7129);
and U7849 (N_7849,N_7145,N_7125);
nor U7850 (N_7850,N_7319,N_7366);
nor U7851 (N_7851,N_7430,N_7273);
nor U7852 (N_7852,N_7287,N_7487);
or U7853 (N_7853,N_7197,N_7090);
nand U7854 (N_7854,N_7221,N_7418);
and U7855 (N_7855,N_7023,N_7232);
nand U7856 (N_7856,N_7400,N_7319);
nand U7857 (N_7857,N_7004,N_7072);
xor U7858 (N_7858,N_7109,N_7463);
xor U7859 (N_7859,N_7239,N_7418);
or U7860 (N_7860,N_7081,N_7050);
nor U7861 (N_7861,N_7034,N_7045);
or U7862 (N_7862,N_7268,N_7029);
nand U7863 (N_7863,N_7348,N_7206);
nand U7864 (N_7864,N_7313,N_7212);
or U7865 (N_7865,N_7291,N_7482);
nor U7866 (N_7866,N_7073,N_7149);
xnor U7867 (N_7867,N_7089,N_7387);
nor U7868 (N_7868,N_7423,N_7243);
nor U7869 (N_7869,N_7046,N_7121);
nor U7870 (N_7870,N_7452,N_7286);
and U7871 (N_7871,N_7261,N_7333);
nor U7872 (N_7872,N_7019,N_7395);
nor U7873 (N_7873,N_7009,N_7288);
and U7874 (N_7874,N_7029,N_7216);
or U7875 (N_7875,N_7285,N_7166);
and U7876 (N_7876,N_7343,N_7344);
xor U7877 (N_7877,N_7423,N_7155);
or U7878 (N_7878,N_7318,N_7065);
nor U7879 (N_7879,N_7211,N_7342);
or U7880 (N_7880,N_7079,N_7358);
xnor U7881 (N_7881,N_7217,N_7132);
nor U7882 (N_7882,N_7406,N_7482);
xor U7883 (N_7883,N_7255,N_7192);
nand U7884 (N_7884,N_7332,N_7208);
nor U7885 (N_7885,N_7122,N_7498);
nand U7886 (N_7886,N_7415,N_7028);
and U7887 (N_7887,N_7291,N_7149);
nor U7888 (N_7888,N_7445,N_7293);
and U7889 (N_7889,N_7134,N_7404);
nor U7890 (N_7890,N_7239,N_7220);
and U7891 (N_7891,N_7075,N_7323);
and U7892 (N_7892,N_7366,N_7251);
nand U7893 (N_7893,N_7158,N_7301);
and U7894 (N_7894,N_7259,N_7455);
and U7895 (N_7895,N_7428,N_7238);
nor U7896 (N_7896,N_7062,N_7290);
nand U7897 (N_7897,N_7151,N_7180);
xor U7898 (N_7898,N_7413,N_7052);
xnor U7899 (N_7899,N_7068,N_7112);
or U7900 (N_7900,N_7288,N_7294);
and U7901 (N_7901,N_7242,N_7426);
nand U7902 (N_7902,N_7312,N_7015);
nand U7903 (N_7903,N_7405,N_7114);
and U7904 (N_7904,N_7287,N_7053);
and U7905 (N_7905,N_7314,N_7256);
or U7906 (N_7906,N_7167,N_7127);
xor U7907 (N_7907,N_7081,N_7250);
or U7908 (N_7908,N_7424,N_7032);
xor U7909 (N_7909,N_7155,N_7137);
xnor U7910 (N_7910,N_7419,N_7034);
xor U7911 (N_7911,N_7158,N_7393);
nor U7912 (N_7912,N_7215,N_7032);
xnor U7913 (N_7913,N_7277,N_7140);
and U7914 (N_7914,N_7087,N_7341);
xnor U7915 (N_7915,N_7487,N_7232);
nor U7916 (N_7916,N_7289,N_7209);
nand U7917 (N_7917,N_7187,N_7291);
and U7918 (N_7918,N_7237,N_7440);
or U7919 (N_7919,N_7009,N_7346);
nor U7920 (N_7920,N_7008,N_7118);
or U7921 (N_7921,N_7325,N_7024);
and U7922 (N_7922,N_7335,N_7251);
xor U7923 (N_7923,N_7400,N_7144);
nand U7924 (N_7924,N_7372,N_7454);
nand U7925 (N_7925,N_7288,N_7273);
nand U7926 (N_7926,N_7477,N_7295);
or U7927 (N_7927,N_7422,N_7103);
or U7928 (N_7928,N_7368,N_7189);
nor U7929 (N_7929,N_7268,N_7428);
nor U7930 (N_7930,N_7029,N_7132);
or U7931 (N_7931,N_7123,N_7214);
xnor U7932 (N_7932,N_7292,N_7294);
nor U7933 (N_7933,N_7299,N_7460);
nor U7934 (N_7934,N_7371,N_7158);
nand U7935 (N_7935,N_7067,N_7301);
and U7936 (N_7936,N_7467,N_7432);
nor U7937 (N_7937,N_7195,N_7197);
nand U7938 (N_7938,N_7144,N_7102);
or U7939 (N_7939,N_7067,N_7292);
or U7940 (N_7940,N_7010,N_7089);
nand U7941 (N_7941,N_7065,N_7074);
xnor U7942 (N_7942,N_7426,N_7194);
and U7943 (N_7943,N_7140,N_7148);
xor U7944 (N_7944,N_7004,N_7193);
nor U7945 (N_7945,N_7078,N_7291);
or U7946 (N_7946,N_7349,N_7227);
xor U7947 (N_7947,N_7158,N_7182);
and U7948 (N_7948,N_7001,N_7210);
nor U7949 (N_7949,N_7445,N_7303);
xor U7950 (N_7950,N_7097,N_7243);
xnor U7951 (N_7951,N_7116,N_7304);
nor U7952 (N_7952,N_7443,N_7234);
xnor U7953 (N_7953,N_7343,N_7462);
and U7954 (N_7954,N_7038,N_7324);
or U7955 (N_7955,N_7259,N_7075);
and U7956 (N_7956,N_7453,N_7263);
xor U7957 (N_7957,N_7099,N_7422);
nor U7958 (N_7958,N_7431,N_7382);
or U7959 (N_7959,N_7167,N_7256);
nor U7960 (N_7960,N_7226,N_7274);
or U7961 (N_7961,N_7437,N_7212);
nor U7962 (N_7962,N_7301,N_7101);
nor U7963 (N_7963,N_7461,N_7262);
or U7964 (N_7964,N_7108,N_7130);
or U7965 (N_7965,N_7464,N_7402);
or U7966 (N_7966,N_7373,N_7158);
nor U7967 (N_7967,N_7414,N_7130);
nor U7968 (N_7968,N_7441,N_7055);
or U7969 (N_7969,N_7014,N_7124);
nor U7970 (N_7970,N_7486,N_7480);
and U7971 (N_7971,N_7247,N_7290);
and U7972 (N_7972,N_7201,N_7465);
nor U7973 (N_7973,N_7007,N_7245);
xor U7974 (N_7974,N_7015,N_7256);
nand U7975 (N_7975,N_7157,N_7185);
nand U7976 (N_7976,N_7162,N_7259);
xor U7977 (N_7977,N_7304,N_7362);
nand U7978 (N_7978,N_7234,N_7051);
nand U7979 (N_7979,N_7490,N_7131);
and U7980 (N_7980,N_7103,N_7495);
nand U7981 (N_7981,N_7229,N_7273);
nor U7982 (N_7982,N_7337,N_7495);
xnor U7983 (N_7983,N_7011,N_7223);
or U7984 (N_7984,N_7116,N_7069);
nor U7985 (N_7985,N_7322,N_7275);
and U7986 (N_7986,N_7228,N_7173);
or U7987 (N_7987,N_7323,N_7080);
nand U7988 (N_7988,N_7233,N_7427);
nor U7989 (N_7989,N_7199,N_7257);
and U7990 (N_7990,N_7474,N_7450);
nand U7991 (N_7991,N_7467,N_7095);
nor U7992 (N_7992,N_7361,N_7481);
or U7993 (N_7993,N_7160,N_7494);
or U7994 (N_7994,N_7163,N_7094);
xnor U7995 (N_7995,N_7201,N_7469);
nor U7996 (N_7996,N_7229,N_7499);
nor U7997 (N_7997,N_7218,N_7027);
xnor U7998 (N_7998,N_7283,N_7234);
or U7999 (N_7999,N_7071,N_7355);
nand U8000 (N_8000,N_7995,N_7643);
nand U8001 (N_8001,N_7659,N_7953);
or U8002 (N_8002,N_7554,N_7522);
or U8003 (N_8003,N_7834,N_7913);
and U8004 (N_8004,N_7757,N_7610);
and U8005 (N_8005,N_7745,N_7993);
nand U8006 (N_8006,N_7883,N_7588);
nor U8007 (N_8007,N_7678,N_7507);
and U8008 (N_8008,N_7889,N_7662);
or U8009 (N_8009,N_7839,N_7682);
and U8010 (N_8010,N_7797,N_7840);
and U8011 (N_8011,N_7697,N_7653);
nor U8012 (N_8012,N_7894,N_7852);
and U8013 (N_8013,N_7543,N_7742);
xor U8014 (N_8014,N_7957,N_7578);
xor U8015 (N_8015,N_7676,N_7885);
nand U8016 (N_8016,N_7509,N_7517);
and U8017 (N_8017,N_7639,N_7626);
nand U8018 (N_8018,N_7560,N_7825);
or U8019 (N_8019,N_7919,N_7935);
nand U8020 (N_8020,N_7506,N_7743);
and U8021 (N_8021,N_7673,N_7977);
and U8022 (N_8022,N_7669,N_7955);
or U8023 (N_8023,N_7721,N_7739);
nand U8024 (N_8024,N_7633,N_7573);
nand U8025 (N_8025,N_7539,N_7727);
nand U8026 (N_8026,N_7777,N_7966);
xor U8027 (N_8027,N_7814,N_7500);
and U8028 (N_8028,N_7803,N_7950);
nor U8029 (N_8029,N_7940,N_7774);
and U8030 (N_8030,N_7606,N_7783);
xor U8031 (N_8031,N_7901,N_7635);
and U8032 (N_8032,N_7607,N_7971);
and U8033 (N_8033,N_7645,N_7609);
or U8034 (N_8034,N_7579,N_7587);
xor U8035 (N_8035,N_7747,N_7824);
nand U8036 (N_8036,N_7755,N_7740);
and U8037 (N_8037,N_7851,N_7605);
and U8038 (N_8038,N_7594,N_7680);
and U8039 (N_8039,N_7695,N_7799);
and U8040 (N_8040,N_7722,N_7880);
nand U8041 (N_8041,N_7692,N_7984);
xnor U8042 (N_8042,N_7709,N_7693);
nor U8043 (N_8043,N_7846,N_7884);
and U8044 (N_8044,N_7881,N_7780);
or U8045 (N_8045,N_7925,N_7705);
or U8046 (N_8046,N_7903,N_7862);
and U8047 (N_8047,N_7703,N_7915);
nor U8048 (N_8048,N_7823,N_7948);
or U8049 (N_8049,N_7752,N_7636);
nand U8050 (N_8050,N_7656,N_7949);
and U8051 (N_8051,N_7535,N_7622);
nor U8052 (N_8052,N_7991,N_7658);
or U8053 (N_8053,N_7572,N_7976);
xor U8054 (N_8054,N_7891,N_7576);
xor U8055 (N_8055,N_7688,N_7627);
or U8056 (N_8056,N_7530,N_7537);
or U8057 (N_8057,N_7741,N_7564);
nand U8058 (N_8058,N_7638,N_7833);
xnor U8059 (N_8059,N_7596,N_7683);
or U8060 (N_8060,N_7524,N_7865);
or U8061 (N_8061,N_7598,N_7951);
nor U8062 (N_8062,N_7921,N_7972);
nand U8063 (N_8063,N_7569,N_7781);
nand U8064 (N_8064,N_7749,N_7544);
xor U8065 (N_8065,N_7527,N_7860);
or U8066 (N_8066,N_7603,N_7973);
nor U8067 (N_8067,N_7748,N_7580);
or U8068 (N_8068,N_7581,N_7806);
xnor U8069 (N_8069,N_7735,N_7649);
nor U8070 (N_8070,N_7821,N_7808);
and U8071 (N_8071,N_7967,N_7734);
nand U8072 (N_8072,N_7952,N_7687);
and U8073 (N_8073,N_7796,N_7556);
xor U8074 (N_8074,N_7947,N_7970);
and U8075 (N_8075,N_7988,N_7866);
or U8076 (N_8076,N_7856,N_7829);
xnor U8077 (N_8077,N_7779,N_7983);
xnor U8078 (N_8078,N_7784,N_7864);
nand U8079 (N_8079,N_7545,N_7912);
nor U8080 (N_8080,N_7667,N_7763);
nor U8081 (N_8081,N_7718,N_7514);
and U8082 (N_8082,N_7920,N_7845);
and U8083 (N_8083,N_7512,N_7548);
xor U8084 (N_8084,N_7801,N_7657);
xnor U8085 (N_8085,N_7532,N_7867);
xor U8086 (N_8086,N_7922,N_7505);
xnor U8087 (N_8087,N_7761,N_7561);
nand U8088 (N_8088,N_7965,N_7568);
nor U8089 (N_8089,N_7769,N_7508);
or U8090 (N_8090,N_7802,N_7835);
or U8091 (N_8091,N_7621,N_7759);
nor U8092 (N_8092,N_7652,N_7790);
xor U8093 (N_8093,N_7736,N_7661);
nor U8094 (N_8094,N_7617,N_7985);
nor U8095 (N_8095,N_7744,N_7758);
nand U8096 (N_8096,N_7869,N_7832);
xnor U8097 (N_8097,N_7665,N_7997);
and U8098 (N_8098,N_7941,N_7675);
nor U8099 (N_8099,N_7521,N_7904);
nand U8100 (N_8100,N_7936,N_7751);
nor U8101 (N_8101,N_7716,N_7592);
nor U8102 (N_8102,N_7956,N_7926);
or U8103 (N_8103,N_7786,N_7504);
or U8104 (N_8104,N_7859,N_7690);
and U8105 (N_8105,N_7794,N_7525);
or U8106 (N_8106,N_7644,N_7989);
or U8107 (N_8107,N_7932,N_7830);
or U8108 (N_8108,N_7681,N_7520);
or U8109 (N_8109,N_7529,N_7927);
nor U8110 (N_8110,N_7563,N_7874);
xor U8111 (N_8111,N_7717,N_7879);
or U8112 (N_8112,N_7651,N_7708);
nor U8113 (N_8113,N_7551,N_7642);
or U8114 (N_8114,N_7836,N_7728);
nand U8115 (N_8115,N_7768,N_7618);
xnor U8116 (N_8116,N_7906,N_7677);
and U8117 (N_8117,N_7704,N_7929);
xor U8118 (N_8118,N_7961,N_7730);
and U8119 (N_8119,N_7600,N_7624);
xor U8120 (N_8120,N_7898,N_7994);
nand U8121 (N_8121,N_7637,N_7646);
or U8122 (N_8122,N_7868,N_7798);
or U8123 (N_8123,N_7541,N_7733);
nor U8124 (N_8124,N_7540,N_7987);
xor U8125 (N_8125,N_7619,N_7582);
and U8126 (N_8126,N_7907,N_7756);
or U8127 (N_8127,N_7788,N_7583);
or U8128 (N_8128,N_7914,N_7818);
nand U8129 (N_8129,N_7902,N_7844);
or U8130 (N_8130,N_7899,N_7555);
and U8131 (N_8131,N_7848,N_7738);
nand U8132 (N_8132,N_7916,N_7893);
nor U8133 (N_8133,N_7599,N_7820);
and U8134 (N_8134,N_7723,N_7699);
xnor U8135 (N_8135,N_7562,N_7849);
nor U8136 (N_8136,N_7910,N_7791);
xor U8137 (N_8137,N_7767,N_7625);
and U8138 (N_8138,N_7511,N_7623);
nand U8139 (N_8139,N_7574,N_7945);
nand U8140 (N_8140,N_7978,N_7855);
nor U8141 (N_8141,N_7776,N_7773);
xnor U8142 (N_8142,N_7770,N_7990);
or U8143 (N_8143,N_7700,N_7655);
nor U8144 (N_8144,N_7558,N_7611);
xor U8145 (N_8145,N_7577,N_7602);
nand U8146 (N_8146,N_7533,N_7567);
and U8147 (N_8147,N_7595,N_7672);
and U8148 (N_8148,N_7895,N_7519);
or U8149 (N_8149,N_7584,N_7805);
or U8150 (N_8150,N_7996,N_7954);
or U8151 (N_8151,N_7754,N_7559);
nor U8152 (N_8152,N_7842,N_7850);
xor U8153 (N_8153,N_7597,N_7931);
xor U8154 (N_8154,N_7946,N_7992);
and U8155 (N_8155,N_7974,N_7923);
and U8156 (N_8156,N_7890,N_7590);
or U8157 (N_8157,N_7979,N_7710);
or U8158 (N_8158,N_7612,N_7811);
nor U8159 (N_8159,N_7944,N_7817);
nor U8160 (N_8160,N_7601,N_7650);
xor U8161 (N_8161,N_7882,N_7765);
or U8162 (N_8162,N_7552,N_7518);
or U8163 (N_8163,N_7795,N_7875);
or U8164 (N_8164,N_7760,N_7831);
nand U8165 (N_8165,N_7613,N_7571);
and U8166 (N_8166,N_7968,N_7629);
nor U8167 (N_8167,N_7871,N_7711);
xnor U8168 (N_8168,N_7648,N_7822);
nor U8169 (N_8169,N_7538,N_7837);
nor U8170 (N_8170,N_7557,N_7876);
xnor U8171 (N_8171,N_7698,N_7707);
xnor U8172 (N_8172,N_7685,N_7816);
nor U8173 (N_8173,N_7838,N_7604);
or U8174 (N_8174,N_7887,N_7691);
xor U8175 (N_8175,N_7523,N_7515);
xnor U8176 (N_8176,N_7980,N_7666);
or U8177 (N_8177,N_7960,N_7858);
or U8178 (N_8178,N_7812,N_7775);
and U8179 (N_8179,N_7719,N_7958);
xnor U8180 (N_8180,N_7975,N_7510);
nand U8181 (N_8181,N_7826,N_7789);
and U8182 (N_8182,N_7905,N_7632);
xor U8183 (N_8183,N_7917,N_7939);
nand U8184 (N_8184,N_7702,N_7663);
xnor U8185 (N_8185,N_7896,N_7766);
nor U8186 (N_8186,N_7872,N_7550);
or U8187 (N_8187,N_7679,N_7696);
or U8188 (N_8188,N_7892,N_7746);
and U8189 (N_8189,N_7634,N_7998);
nor U8190 (N_8190,N_7918,N_7706);
xor U8191 (N_8191,N_7565,N_7531);
nand U8192 (N_8192,N_7630,N_7999);
and U8193 (N_8193,N_7566,N_7782);
nand U8194 (N_8194,N_7647,N_7857);
or U8195 (N_8195,N_7615,N_7620);
nand U8196 (N_8196,N_7962,N_7528);
nand U8197 (N_8197,N_7593,N_7928);
nor U8198 (N_8198,N_7726,N_7686);
and U8199 (N_8199,N_7668,N_7516);
and U8200 (N_8200,N_7715,N_7841);
and U8201 (N_8201,N_7526,N_7942);
nor U8202 (N_8202,N_7843,N_7877);
and U8203 (N_8203,N_7720,N_7713);
xnor U8204 (N_8204,N_7809,N_7753);
nand U8205 (N_8205,N_7986,N_7724);
nor U8206 (N_8206,N_7654,N_7810);
nand U8207 (N_8207,N_7847,N_7542);
or U8208 (N_8208,N_7959,N_7828);
and U8209 (N_8209,N_7502,N_7701);
nor U8210 (N_8210,N_7764,N_7964);
xor U8211 (N_8211,N_7900,N_7793);
nand U8212 (N_8212,N_7750,N_7553);
nor U8213 (N_8213,N_7897,N_7870);
nand U8214 (N_8214,N_7631,N_7501);
nand U8215 (N_8215,N_7863,N_7924);
nor U8216 (N_8216,N_7819,N_7725);
or U8217 (N_8217,N_7547,N_7772);
and U8218 (N_8218,N_7640,N_7908);
or U8219 (N_8219,N_7614,N_7660);
nor U8220 (N_8220,N_7591,N_7787);
or U8221 (N_8221,N_7714,N_7981);
or U8222 (N_8222,N_7549,N_7873);
xnor U8223 (N_8223,N_7616,N_7513);
nor U8224 (N_8224,N_7503,N_7813);
xnor U8225 (N_8225,N_7674,N_7628);
nand U8226 (N_8226,N_7778,N_7854);
xor U8227 (N_8227,N_7943,N_7732);
xnor U8228 (N_8228,N_7888,N_7608);
and U8229 (N_8229,N_7963,N_7815);
nor U8230 (N_8230,N_7546,N_7689);
and U8231 (N_8231,N_7712,N_7586);
nor U8232 (N_8232,N_7878,N_7771);
xor U8233 (N_8233,N_7737,N_7969);
nor U8234 (N_8234,N_7534,N_7575);
or U8235 (N_8235,N_7807,N_7585);
nor U8236 (N_8236,N_7827,N_7536);
or U8237 (N_8237,N_7886,N_7729);
and U8238 (N_8238,N_7933,N_7909);
nor U8239 (N_8239,N_7731,N_7861);
nand U8240 (N_8240,N_7670,N_7937);
and U8241 (N_8241,N_7938,N_7664);
nor U8242 (N_8242,N_7589,N_7804);
nand U8243 (N_8243,N_7694,N_7930);
nand U8244 (N_8244,N_7982,N_7853);
or U8245 (N_8245,N_7934,N_7762);
or U8246 (N_8246,N_7911,N_7684);
xnor U8247 (N_8247,N_7570,N_7785);
xnor U8248 (N_8248,N_7792,N_7800);
nor U8249 (N_8249,N_7641,N_7671);
nor U8250 (N_8250,N_7846,N_7943);
or U8251 (N_8251,N_7697,N_7836);
or U8252 (N_8252,N_7937,N_7839);
nand U8253 (N_8253,N_7504,N_7867);
and U8254 (N_8254,N_7996,N_7515);
or U8255 (N_8255,N_7987,N_7582);
and U8256 (N_8256,N_7765,N_7687);
or U8257 (N_8257,N_7580,N_7612);
or U8258 (N_8258,N_7518,N_7594);
or U8259 (N_8259,N_7613,N_7780);
xor U8260 (N_8260,N_7717,N_7516);
xor U8261 (N_8261,N_7796,N_7755);
and U8262 (N_8262,N_7907,N_7776);
and U8263 (N_8263,N_7727,N_7933);
nand U8264 (N_8264,N_7731,N_7711);
and U8265 (N_8265,N_7777,N_7828);
xor U8266 (N_8266,N_7686,N_7953);
nor U8267 (N_8267,N_7640,N_7874);
xnor U8268 (N_8268,N_7945,N_7587);
and U8269 (N_8269,N_7526,N_7551);
and U8270 (N_8270,N_7636,N_7889);
and U8271 (N_8271,N_7660,N_7781);
nand U8272 (N_8272,N_7542,N_7851);
xor U8273 (N_8273,N_7794,N_7745);
nand U8274 (N_8274,N_7884,N_7879);
nand U8275 (N_8275,N_7994,N_7939);
nor U8276 (N_8276,N_7698,N_7846);
xor U8277 (N_8277,N_7651,N_7559);
and U8278 (N_8278,N_7983,N_7961);
and U8279 (N_8279,N_7767,N_7782);
nand U8280 (N_8280,N_7814,N_7755);
nor U8281 (N_8281,N_7671,N_7882);
or U8282 (N_8282,N_7518,N_7805);
xor U8283 (N_8283,N_7692,N_7968);
or U8284 (N_8284,N_7961,N_7713);
or U8285 (N_8285,N_7630,N_7628);
and U8286 (N_8286,N_7745,N_7817);
and U8287 (N_8287,N_7809,N_7745);
or U8288 (N_8288,N_7869,N_7839);
and U8289 (N_8289,N_7837,N_7938);
xor U8290 (N_8290,N_7851,N_7639);
nor U8291 (N_8291,N_7986,N_7722);
or U8292 (N_8292,N_7979,N_7928);
and U8293 (N_8293,N_7665,N_7699);
xor U8294 (N_8294,N_7790,N_7716);
or U8295 (N_8295,N_7515,N_7992);
nand U8296 (N_8296,N_7791,N_7847);
and U8297 (N_8297,N_7733,N_7572);
xnor U8298 (N_8298,N_7882,N_7605);
xnor U8299 (N_8299,N_7672,N_7737);
xor U8300 (N_8300,N_7722,N_7634);
nand U8301 (N_8301,N_7628,N_7963);
nor U8302 (N_8302,N_7637,N_7556);
nor U8303 (N_8303,N_7988,N_7763);
and U8304 (N_8304,N_7507,N_7660);
or U8305 (N_8305,N_7922,N_7959);
xor U8306 (N_8306,N_7900,N_7657);
nand U8307 (N_8307,N_7960,N_7967);
and U8308 (N_8308,N_7958,N_7517);
nor U8309 (N_8309,N_7920,N_7559);
and U8310 (N_8310,N_7544,N_7715);
or U8311 (N_8311,N_7725,N_7661);
nor U8312 (N_8312,N_7504,N_7559);
nand U8313 (N_8313,N_7714,N_7938);
xor U8314 (N_8314,N_7765,N_7908);
or U8315 (N_8315,N_7884,N_7908);
nor U8316 (N_8316,N_7983,N_7967);
or U8317 (N_8317,N_7988,N_7679);
and U8318 (N_8318,N_7663,N_7970);
nand U8319 (N_8319,N_7938,N_7585);
nand U8320 (N_8320,N_7839,N_7509);
xor U8321 (N_8321,N_7849,N_7764);
xor U8322 (N_8322,N_7821,N_7905);
nor U8323 (N_8323,N_7615,N_7770);
xnor U8324 (N_8324,N_7923,N_7838);
nor U8325 (N_8325,N_7753,N_7607);
xnor U8326 (N_8326,N_7850,N_7906);
and U8327 (N_8327,N_7843,N_7610);
nor U8328 (N_8328,N_7868,N_7570);
and U8329 (N_8329,N_7928,N_7701);
or U8330 (N_8330,N_7841,N_7599);
xor U8331 (N_8331,N_7767,N_7535);
and U8332 (N_8332,N_7916,N_7621);
or U8333 (N_8333,N_7891,N_7995);
and U8334 (N_8334,N_7813,N_7839);
nor U8335 (N_8335,N_7850,N_7641);
or U8336 (N_8336,N_7641,N_7992);
or U8337 (N_8337,N_7662,N_7634);
xnor U8338 (N_8338,N_7786,N_7587);
or U8339 (N_8339,N_7621,N_7567);
and U8340 (N_8340,N_7910,N_7635);
and U8341 (N_8341,N_7702,N_7533);
xnor U8342 (N_8342,N_7761,N_7900);
xor U8343 (N_8343,N_7568,N_7867);
or U8344 (N_8344,N_7705,N_7749);
nand U8345 (N_8345,N_7975,N_7922);
nor U8346 (N_8346,N_7782,N_7944);
nor U8347 (N_8347,N_7925,N_7554);
and U8348 (N_8348,N_7789,N_7816);
xor U8349 (N_8349,N_7882,N_7536);
or U8350 (N_8350,N_7962,N_7710);
nor U8351 (N_8351,N_7885,N_7863);
or U8352 (N_8352,N_7959,N_7606);
and U8353 (N_8353,N_7817,N_7599);
and U8354 (N_8354,N_7624,N_7581);
nor U8355 (N_8355,N_7783,N_7805);
and U8356 (N_8356,N_7511,N_7728);
and U8357 (N_8357,N_7857,N_7629);
nor U8358 (N_8358,N_7639,N_7861);
nor U8359 (N_8359,N_7651,N_7874);
xor U8360 (N_8360,N_7583,N_7963);
and U8361 (N_8361,N_7966,N_7590);
and U8362 (N_8362,N_7625,N_7520);
nor U8363 (N_8363,N_7648,N_7915);
or U8364 (N_8364,N_7651,N_7524);
xor U8365 (N_8365,N_7972,N_7577);
nor U8366 (N_8366,N_7521,N_7687);
or U8367 (N_8367,N_7895,N_7543);
or U8368 (N_8368,N_7924,N_7622);
xor U8369 (N_8369,N_7957,N_7735);
nand U8370 (N_8370,N_7850,N_7690);
xnor U8371 (N_8371,N_7889,N_7677);
or U8372 (N_8372,N_7995,N_7740);
and U8373 (N_8373,N_7962,N_7818);
xor U8374 (N_8374,N_7829,N_7925);
or U8375 (N_8375,N_7574,N_7751);
or U8376 (N_8376,N_7668,N_7959);
nor U8377 (N_8377,N_7903,N_7778);
nor U8378 (N_8378,N_7719,N_7527);
or U8379 (N_8379,N_7837,N_7887);
xor U8380 (N_8380,N_7911,N_7663);
and U8381 (N_8381,N_7855,N_7940);
xnor U8382 (N_8382,N_7909,N_7641);
nor U8383 (N_8383,N_7748,N_7581);
nor U8384 (N_8384,N_7732,N_7635);
nand U8385 (N_8385,N_7645,N_7594);
nand U8386 (N_8386,N_7707,N_7972);
or U8387 (N_8387,N_7718,N_7842);
or U8388 (N_8388,N_7888,N_7675);
nor U8389 (N_8389,N_7562,N_7558);
nand U8390 (N_8390,N_7970,N_7526);
or U8391 (N_8391,N_7978,N_7868);
and U8392 (N_8392,N_7577,N_7631);
xor U8393 (N_8393,N_7821,N_7840);
and U8394 (N_8394,N_7584,N_7524);
xor U8395 (N_8395,N_7531,N_7580);
xnor U8396 (N_8396,N_7524,N_7867);
or U8397 (N_8397,N_7783,N_7878);
and U8398 (N_8398,N_7890,N_7858);
nor U8399 (N_8399,N_7768,N_7587);
nand U8400 (N_8400,N_7998,N_7960);
nor U8401 (N_8401,N_7639,N_7808);
xnor U8402 (N_8402,N_7771,N_7990);
or U8403 (N_8403,N_7763,N_7932);
and U8404 (N_8404,N_7903,N_7766);
or U8405 (N_8405,N_7898,N_7869);
xor U8406 (N_8406,N_7651,N_7564);
nor U8407 (N_8407,N_7661,N_7595);
or U8408 (N_8408,N_7506,N_7976);
xnor U8409 (N_8409,N_7615,N_7678);
nor U8410 (N_8410,N_7822,N_7918);
and U8411 (N_8411,N_7825,N_7717);
or U8412 (N_8412,N_7988,N_7655);
or U8413 (N_8413,N_7810,N_7989);
or U8414 (N_8414,N_7684,N_7561);
xnor U8415 (N_8415,N_7514,N_7576);
or U8416 (N_8416,N_7750,N_7952);
xnor U8417 (N_8417,N_7848,N_7913);
or U8418 (N_8418,N_7879,N_7719);
or U8419 (N_8419,N_7906,N_7817);
or U8420 (N_8420,N_7810,N_7628);
xor U8421 (N_8421,N_7784,N_7530);
nand U8422 (N_8422,N_7734,N_7671);
or U8423 (N_8423,N_7619,N_7819);
or U8424 (N_8424,N_7660,N_7983);
and U8425 (N_8425,N_7503,N_7753);
and U8426 (N_8426,N_7773,N_7702);
or U8427 (N_8427,N_7880,N_7937);
or U8428 (N_8428,N_7829,N_7815);
nor U8429 (N_8429,N_7995,N_7523);
nand U8430 (N_8430,N_7926,N_7611);
xnor U8431 (N_8431,N_7549,N_7705);
nand U8432 (N_8432,N_7766,N_7724);
or U8433 (N_8433,N_7651,N_7671);
nand U8434 (N_8434,N_7658,N_7906);
and U8435 (N_8435,N_7521,N_7715);
and U8436 (N_8436,N_7559,N_7916);
or U8437 (N_8437,N_7790,N_7810);
nor U8438 (N_8438,N_7914,N_7525);
nor U8439 (N_8439,N_7845,N_7755);
nand U8440 (N_8440,N_7696,N_7996);
nor U8441 (N_8441,N_7728,N_7733);
nand U8442 (N_8442,N_7570,N_7979);
xnor U8443 (N_8443,N_7858,N_7525);
xnor U8444 (N_8444,N_7875,N_7557);
nand U8445 (N_8445,N_7917,N_7586);
nand U8446 (N_8446,N_7599,N_7584);
nand U8447 (N_8447,N_7519,N_7626);
nand U8448 (N_8448,N_7967,N_7543);
xnor U8449 (N_8449,N_7807,N_7752);
and U8450 (N_8450,N_7945,N_7511);
nand U8451 (N_8451,N_7587,N_7852);
or U8452 (N_8452,N_7579,N_7527);
or U8453 (N_8453,N_7690,N_7726);
and U8454 (N_8454,N_7575,N_7666);
or U8455 (N_8455,N_7562,N_7584);
and U8456 (N_8456,N_7638,N_7856);
nand U8457 (N_8457,N_7607,N_7519);
xnor U8458 (N_8458,N_7562,N_7888);
xor U8459 (N_8459,N_7670,N_7909);
xor U8460 (N_8460,N_7993,N_7623);
xnor U8461 (N_8461,N_7848,N_7824);
nand U8462 (N_8462,N_7858,N_7568);
or U8463 (N_8463,N_7805,N_7593);
and U8464 (N_8464,N_7881,N_7684);
nand U8465 (N_8465,N_7952,N_7937);
or U8466 (N_8466,N_7706,N_7584);
xor U8467 (N_8467,N_7645,N_7600);
nand U8468 (N_8468,N_7785,N_7762);
nor U8469 (N_8469,N_7866,N_7929);
nand U8470 (N_8470,N_7710,N_7741);
nand U8471 (N_8471,N_7589,N_7963);
or U8472 (N_8472,N_7787,N_7576);
nor U8473 (N_8473,N_7636,N_7527);
and U8474 (N_8474,N_7834,N_7534);
xor U8475 (N_8475,N_7762,N_7944);
or U8476 (N_8476,N_7855,N_7595);
xnor U8477 (N_8477,N_7962,N_7888);
nand U8478 (N_8478,N_7537,N_7861);
and U8479 (N_8479,N_7729,N_7766);
and U8480 (N_8480,N_7921,N_7548);
and U8481 (N_8481,N_7985,N_7735);
or U8482 (N_8482,N_7987,N_7979);
nor U8483 (N_8483,N_7920,N_7910);
xor U8484 (N_8484,N_7579,N_7551);
nand U8485 (N_8485,N_7535,N_7634);
or U8486 (N_8486,N_7985,N_7791);
nand U8487 (N_8487,N_7654,N_7601);
nand U8488 (N_8488,N_7830,N_7653);
or U8489 (N_8489,N_7975,N_7999);
or U8490 (N_8490,N_7609,N_7779);
xor U8491 (N_8491,N_7926,N_7512);
or U8492 (N_8492,N_7824,N_7920);
xnor U8493 (N_8493,N_7544,N_7556);
and U8494 (N_8494,N_7676,N_7917);
nor U8495 (N_8495,N_7922,N_7794);
nand U8496 (N_8496,N_7949,N_7748);
or U8497 (N_8497,N_7566,N_7570);
and U8498 (N_8498,N_7542,N_7890);
nor U8499 (N_8499,N_7811,N_7710);
or U8500 (N_8500,N_8314,N_8300);
or U8501 (N_8501,N_8195,N_8013);
and U8502 (N_8502,N_8169,N_8163);
nand U8503 (N_8503,N_8157,N_8331);
and U8504 (N_8504,N_8346,N_8342);
xor U8505 (N_8505,N_8375,N_8414);
xor U8506 (N_8506,N_8036,N_8381);
nand U8507 (N_8507,N_8485,N_8246);
or U8508 (N_8508,N_8389,N_8451);
and U8509 (N_8509,N_8085,N_8274);
nand U8510 (N_8510,N_8227,N_8339);
or U8511 (N_8511,N_8432,N_8341);
xor U8512 (N_8512,N_8348,N_8373);
nand U8513 (N_8513,N_8042,N_8398);
and U8514 (N_8514,N_8426,N_8210);
and U8515 (N_8515,N_8333,N_8197);
nor U8516 (N_8516,N_8135,N_8316);
nor U8517 (N_8517,N_8001,N_8264);
and U8518 (N_8518,N_8468,N_8477);
xnor U8519 (N_8519,N_8248,N_8196);
nand U8520 (N_8520,N_8482,N_8077);
xor U8521 (N_8521,N_8450,N_8464);
nand U8522 (N_8522,N_8129,N_8265);
xor U8523 (N_8523,N_8325,N_8453);
or U8524 (N_8524,N_8288,N_8067);
or U8525 (N_8525,N_8437,N_8235);
nor U8526 (N_8526,N_8494,N_8447);
nor U8527 (N_8527,N_8054,N_8062);
nor U8528 (N_8528,N_8297,N_8489);
nor U8529 (N_8529,N_8440,N_8005);
xnor U8530 (N_8530,N_8417,N_8155);
or U8531 (N_8531,N_8383,N_8142);
xor U8532 (N_8532,N_8154,N_8206);
or U8533 (N_8533,N_8324,N_8237);
xnor U8534 (N_8534,N_8467,N_8170);
or U8535 (N_8535,N_8216,N_8117);
nand U8536 (N_8536,N_8349,N_8213);
and U8537 (N_8537,N_8362,N_8483);
and U8538 (N_8538,N_8038,N_8111);
and U8539 (N_8539,N_8037,N_8205);
or U8540 (N_8540,N_8277,N_8069);
nand U8541 (N_8541,N_8397,N_8379);
nand U8542 (N_8542,N_8409,N_8366);
or U8543 (N_8543,N_8025,N_8020);
xnor U8544 (N_8544,N_8484,N_8360);
nand U8545 (N_8545,N_8445,N_8204);
nor U8546 (N_8546,N_8175,N_8420);
and U8547 (N_8547,N_8439,N_8189);
nor U8548 (N_8548,N_8328,N_8030);
nor U8549 (N_8549,N_8088,N_8291);
or U8550 (N_8550,N_8322,N_8177);
xnor U8551 (N_8551,N_8463,N_8161);
or U8552 (N_8552,N_8008,N_8113);
nand U8553 (N_8553,N_8148,N_8416);
xnor U8554 (N_8554,N_8159,N_8101);
nor U8555 (N_8555,N_8065,N_8167);
xor U8556 (N_8556,N_8469,N_8402);
nor U8557 (N_8557,N_8207,N_8405);
or U8558 (N_8558,N_8119,N_8406);
nand U8559 (N_8559,N_8185,N_8344);
xor U8560 (N_8560,N_8260,N_8089);
nor U8561 (N_8561,N_8374,N_8240);
or U8562 (N_8562,N_8456,N_8474);
nand U8563 (N_8563,N_8052,N_8149);
or U8564 (N_8564,N_8329,N_8449);
nand U8565 (N_8565,N_8178,N_8302);
nor U8566 (N_8566,N_8239,N_8462);
xnor U8567 (N_8567,N_8198,N_8433);
and U8568 (N_8568,N_8306,N_8303);
or U8569 (N_8569,N_8243,N_8128);
xor U8570 (N_8570,N_8337,N_8040);
or U8571 (N_8571,N_8047,N_8269);
and U8572 (N_8572,N_8011,N_8233);
and U8573 (N_8573,N_8238,N_8224);
or U8574 (N_8574,N_8024,N_8347);
xor U8575 (N_8575,N_8022,N_8123);
and U8576 (N_8576,N_8340,N_8285);
and U8577 (N_8577,N_8095,N_8415);
and U8578 (N_8578,N_8311,N_8404);
and U8579 (N_8579,N_8292,N_8221);
nor U8580 (N_8580,N_8232,N_8275);
or U8581 (N_8581,N_8493,N_8035);
nand U8582 (N_8582,N_8384,N_8122);
nor U8583 (N_8583,N_8390,N_8293);
xor U8584 (N_8584,N_8106,N_8215);
or U8585 (N_8585,N_8307,N_8225);
xnor U8586 (N_8586,N_8199,N_8470);
or U8587 (N_8587,N_8434,N_8133);
nor U8588 (N_8588,N_8218,N_8211);
nand U8589 (N_8589,N_8317,N_8168);
nand U8590 (N_8590,N_8066,N_8353);
and U8591 (N_8591,N_8299,N_8338);
or U8592 (N_8592,N_8029,N_8446);
or U8593 (N_8593,N_8308,N_8372);
xnor U8594 (N_8594,N_8388,N_8202);
or U8595 (N_8595,N_8112,N_8244);
xnor U8596 (N_8596,N_8130,N_8352);
nand U8597 (N_8597,N_8043,N_8438);
nand U8598 (N_8598,N_8153,N_8137);
nor U8599 (N_8599,N_8368,N_8051);
nor U8600 (N_8600,N_8027,N_8002);
or U8601 (N_8601,N_8249,N_8105);
nor U8602 (N_8602,N_8487,N_8096);
nor U8603 (N_8603,N_8162,N_8378);
or U8604 (N_8604,N_8430,N_8336);
and U8605 (N_8605,N_8026,N_8071);
or U8606 (N_8606,N_8080,N_8012);
nand U8607 (N_8607,N_8212,N_8055);
and U8608 (N_8608,N_8230,N_8284);
nand U8609 (N_8609,N_8323,N_8152);
and U8610 (N_8610,N_8241,N_8190);
nor U8611 (N_8611,N_8072,N_8127);
xor U8612 (N_8612,N_8173,N_8121);
xnor U8613 (N_8613,N_8003,N_8156);
or U8614 (N_8614,N_8073,N_8321);
nand U8615 (N_8615,N_8472,N_8318);
or U8616 (N_8616,N_8257,N_8326);
nand U8617 (N_8617,N_8425,N_8018);
xor U8618 (N_8618,N_8354,N_8496);
or U8619 (N_8619,N_8017,N_8343);
and U8620 (N_8620,N_8074,N_8120);
nor U8621 (N_8621,N_8259,N_8041);
nor U8622 (N_8622,N_8330,N_8138);
and U8623 (N_8623,N_8165,N_8186);
and U8624 (N_8624,N_8465,N_8092);
xnor U8625 (N_8625,N_8403,N_8361);
and U8626 (N_8626,N_8242,N_8283);
and U8627 (N_8627,N_8455,N_8049);
xor U8628 (N_8628,N_8282,N_8102);
nor U8629 (N_8629,N_8201,N_8247);
nand U8630 (N_8630,N_8411,N_8234);
nor U8631 (N_8631,N_8441,N_8401);
nand U8632 (N_8632,N_8287,N_8399);
xnor U8633 (N_8633,N_8050,N_8236);
and U8634 (N_8634,N_8393,N_8457);
nand U8635 (N_8635,N_8126,N_8454);
xnor U8636 (N_8636,N_8083,N_8193);
nor U8637 (N_8637,N_8486,N_8222);
nand U8638 (N_8638,N_8476,N_8315);
or U8639 (N_8639,N_8164,N_8082);
nand U8640 (N_8640,N_8116,N_8488);
or U8641 (N_8641,N_8394,N_8104);
or U8642 (N_8642,N_8034,N_8160);
xnor U8643 (N_8643,N_8363,N_8079);
nand U8644 (N_8644,N_8498,N_8256);
and U8645 (N_8645,N_8320,N_8053);
or U8646 (N_8646,N_8107,N_8253);
nand U8647 (N_8647,N_8281,N_8332);
or U8648 (N_8648,N_8408,N_8109);
nand U8649 (N_8649,N_8499,N_8098);
or U8650 (N_8650,N_8100,N_8427);
nand U8651 (N_8651,N_8407,N_8396);
nor U8652 (N_8652,N_8436,N_8214);
xnor U8653 (N_8653,N_8471,N_8171);
nor U8654 (N_8654,N_8431,N_8444);
and U8655 (N_8655,N_8473,N_8060);
or U8656 (N_8656,N_8174,N_8021);
and U8657 (N_8657,N_8391,N_8219);
nand U8658 (N_8658,N_8369,N_8423);
xnor U8659 (N_8659,N_8028,N_8377);
xor U8660 (N_8660,N_8004,N_8191);
and U8661 (N_8661,N_8097,N_8443);
xor U8662 (N_8662,N_8007,N_8015);
xor U8663 (N_8663,N_8327,N_8309);
or U8664 (N_8664,N_8422,N_8263);
xnor U8665 (N_8665,N_8412,N_8166);
nor U8666 (N_8666,N_8298,N_8048);
or U8667 (N_8667,N_8084,N_8192);
or U8668 (N_8668,N_8478,N_8200);
nand U8669 (N_8669,N_8355,N_8245);
and U8670 (N_8670,N_8495,N_8187);
xnor U8671 (N_8671,N_8124,N_8305);
xnor U8672 (N_8672,N_8480,N_8076);
or U8673 (N_8673,N_8086,N_8270);
and U8674 (N_8674,N_8118,N_8176);
nor U8675 (N_8675,N_8180,N_8370);
or U8676 (N_8676,N_8458,N_8087);
or U8677 (N_8677,N_8250,N_8057);
nand U8678 (N_8678,N_8358,N_8497);
nor U8679 (N_8679,N_8364,N_8271);
nor U8680 (N_8680,N_8070,N_8386);
and U8681 (N_8681,N_8385,N_8461);
nand U8682 (N_8682,N_8146,N_8217);
or U8683 (N_8683,N_8075,N_8081);
xnor U8684 (N_8684,N_8115,N_8421);
xnor U8685 (N_8685,N_8045,N_8276);
or U8686 (N_8686,N_8139,N_8475);
xnor U8687 (N_8687,N_8382,N_8261);
or U8688 (N_8688,N_8194,N_8428);
and U8689 (N_8689,N_8481,N_8351);
and U8690 (N_8690,N_8273,N_8345);
nand U8691 (N_8691,N_8365,N_8304);
nor U8692 (N_8692,N_8290,N_8172);
and U8693 (N_8693,N_8278,N_8289);
nor U8694 (N_8694,N_8229,N_8424);
nand U8695 (N_8695,N_8387,N_8078);
nand U8696 (N_8696,N_8151,N_8359);
or U8697 (N_8697,N_8479,N_8108);
or U8698 (N_8698,N_8091,N_8254);
and U8699 (N_8699,N_8286,N_8114);
nand U8700 (N_8700,N_8145,N_8371);
nor U8701 (N_8701,N_8182,N_8367);
nand U8702 (N_8702,N_8031,N_8132);
xor U8703 (N_8703,N_8255,N_8136);
nand U8704 (N_8704,N_8295,N_8090);
xor U8705 (N_8705,N_8357,N_8103);
nand U8706 (N_8706,N_8044,N_8296);
and U8707 (N_8707,N_8228,N_8014);
nand U8708 (N_8708,N_8064,N_8183);
nor U8709 (N_8709,N_8310,N_8376);
and U8710 (N_8710,N_8061,N_8140);
and U8711 (N_8711,N_8039,N_8063);
xnor U8712 (N_8712,N_8429,N_8334);
nor U8713 (N_8713,N_8350,N_8262);
xor U8714 (N_8714,N_8059,N_8279);
nor U8715 (N_8715,N_8460,N_8413);
and U8716 (N_8716,N_8144,N_8125);
xor U8717 (N_8717,N_8058,N_8010);
xor U8718 (N_8718,N_8395,N_8000);
or U8719 (N_8719,N_8150,N_8442);
nand U8720 (N_8720,N_8452,N_8032);
or U8721 (N_8721,N_8312,N_8143);
or U8722 (N_8722,N_8068,N_8046);
nor U8723 (N_8723,N_8223,N_8006);
nor U8724 (N_8724,N_8147,N_8459);
xnor U8725 (N_8725,N_8466,N_8094);
or U8726 (N_8726,N_8184,N_8272);
nor U8727 (N_8727,N_8016,N_8179);
nor U8728 (N_8728,N_8220,N_8418);
nand U8729 (N_8729,N_8410,N_8188);
nand U8730 (N_8730,N_8280,N_8301);
nand U8731 (N_8731,N_8099,N_8181);
nand U8732 (N_8732,N_8268,N_8258);
or U8733 (N_8733,N_8266,N_8251);
and U8734 (N_8734,N_8208,N_8492);
nand U8735 (N_8735,N_8267,N_8380);
nand U8736 (N_8736,N_8033,N_8356);
nand U8737 (N_8737,N_8203,N_8056);
nand U8738 (N_8738,N_8294,N_8448);
nand U8739 (N_8739,N_8313,N_8110);
nor U8740 (N_8740,N_8491,N_8335);
nand U8741 (N_8741,N_8252,N_8023);
or U8742 (N_8742,N_8400,N_8134);
xnor U8743 (N_8743,N_8392,N_8009);
nand U8744 (N_8744,N_8419,N_8019);
xnor U8745 (N_8745,N_8093,N_8231);
xnor U8746 (N_8746,N_8490,N_8131);
or U8747 (N_8747,N_8158,N_8435);
nand U8748 (N_8748,N_8209,N_8319);
and U8749 (N_8749,N_8141,N_8226);
and U8750 (N_8750,N_8192,N_8287);
nor U8751 (N_8751,N_8103,N_8011);
xnor U8752 (N_8752,N_8393,N_8231);
and U8753 (N_8753,N_8210,N_8419);
nand U8754 (N_8754,N_8469,N_8239);
nor U8755 (N_8755,N_8111,N_8150);
or U8756 (N_8756,N_8469,N_8062);
and U8757 (N_8757,N_8243,N_8388);
or U8758 (N_8758,N_8164,N_8166);
or U8759 (N_8759,N_8333,N_8150);
xor U8760 (N_8760,N_8464,N_8180);
nor U8761 (N_8761,N_8466,N_8005);
xnor U8762 (N_8762,N_8185,N_8017);
xnor U8763 (N_8763,N_8307,N_8051);
nor U8764 (N_8764,N_8496,N_8072);
or U8765 (N_8765,N_8453,N_8044);
nand U8766 (N_8766,N_8199,N_8442);
nand U8767 (N_8767,N_8245,N_8207);
or U8768 (N_8768,N_8427,N_8226);
and U8769 (N_8769,N_8343,N_8487);
or U8770 (N_8770,N_8279,N_8321);
and U8771 (N_8771,N_8189,N_8495);
nor U8772 (N_8772,N_8293,N_8258);
nand U8773 (N_8773,N_8208,N_8064);
or U8774 (N_8774,N_8085,N_8124);
or U8775 (N_8775,N_8305,N_8443);
or U8776 (N_8776,N_8022,N_8291);
nor U8777 (N_8777,N_8044,N_8157);
nand U8778 (N_8778,N_8047,N_8456);
xnor U8779 (N_8779,N_8392,N_8414);
nand U8780 (N_8780,N_8112,N_8289);
and U8781 (N_8781,N_8194,N_8449);
and U8782 (N_8782,N_8453,N_8329);
or U8783 (N_8783,N_8492,N_8326);
and U8784 (N_8784,N_8333,N_8196);
or U8785 (N_8785,N_8041,N_8388);
or U8786 (N_8786,N_8404,N_8433);
nor U8787 (N_8787,N_8057,N_8120);
and U8788 (N_8788,N_8282,N_8499);
nor U8789 (N_8789,N_8385,N_8404);
and U8790 (N_8790,N_8192,N_8289);
xor U8791 (N_8791,N_8040,N_8113);
or U8792 (N_8792,N_8302,N_8060);
or U8793 (N_8793,N_8108,N_8071);
and U8794 (N_8794,N_8044,N_8330);
and U8795 (N_8795,N_8113,N_8166);
nand U8796 (N_8796,N_8157,N_8489);
and U8797 (N_8797,N_8492,N_8413);
nor U8798 (N_8798,N_8376,N_8319);
nor U8799 (N_8799,N_8488,N_8212);
xor U8800 (N_8800,N_8475,N_8101);
nand U8801 (N_8801,N_8038,N_8153);
xnor U8802 (N_8802,N_8178,N_8117);
and U8803 (N_8803,N_8489,N_8482);
or U8804 (N_8804,N_8245,N_8292);
nor U8805 (N_8805,N_8092,N_8217);
nand U8806 (N_8806,N_8430,N_8272);
nand U8807 (N_8807,N_8014,N_8241);
and U8808 (N_8808,N_8231,N_8038);
xnor U8809 (N_8809,N_8296,N_8299);
and U8810 (N_8810,N_8323,N_8026);
nand U8811 (N_8811,N_8295,N_8321);
or U8812 (N_8812,N_8440,N_8468);
or U8813 (N_8813,N_8176,N_8438);
nor U8814 (N_8814,N_8167,N_8222);
nor U8815 (N_8815,N_8434,N_8455);
xor U8816 (N_8816,N_8253,N_8090);
and U8817 (N_8817,N_8091,N_8224);
and U8818 (N_8818,N_8230,N_8334);
nor U8819 (N_8819,N_8479,N_8125);
xnor U8820 (N_8820,N_8161,N_8132);
or U8821 (N_8821,N_8290,N_8392);
or U8822 (N_8822,N_8427,N_8135);
and U8823 (N_8823,N_8047,N_8249);
or U8824 (N_8824,N_8064,N_8457);
xor U8825 (N_8825,N_8175,N_8053);
and U8826 (N_8826,N_8439,N_8096);
xnor U8827 (N_8827,N_8174,N_8414);
nor U8828 (N_8828,N_8240,N_8030);
and U8829 (N_8829,N_8255,N_8015);
nand U8830 (N_8830,N_8405,N_8408);
and U8831 (N_8831,N_8367,N_8217);
or U8832 (N_8832,N_8323,N_8264);
nor U8833 (N_8833,N_8173,N_8105);
and U8834 (N_8834,N_8132,N_8055);
xor U8835 (N_8835,N_8107,N_8045);
nor U8836 (N_8836,N_8315,N_8267);
xnor U8837 (N_8837,N_8132,N_8374);
nor U8838 (N_8838,N_8401,N_8367);
xnor U8839 (N_8839,N_8376,N_8201);
or U8840 (N_8840,N_8246,N_8461);
nor U8841 (N_8841,N_8303,N_8360);
nor U8842 (N_8842,N_8390,N_8275);
or U8843 (N_8843,N_8024,N_8232);
xor U8844 (N_8844,N_8471,N_8415);
and U8845 (N_8845,N_8222,N_8133);
and U8846 (N_8846,N_8362,N_8053);
xor U8847 (N_8847,N_8347,N_8137);
xor U8848 (N_8848,N_8299,N_8231);
nor U8849 (N_8849,N_8384,N_8113);
nand U8850 (N_8850,N_8025,N_8340);
and U8851 (N_8851,N_8072,N_8134);
nor U8852 (N_8852,N_8170,N_8261);
nor U8853 (N_8853,N_8252,N_8334);
nor U8854 (N_8854,N_8009,N_8122);
xor U8855 (N_8855,N_8349,N_8325);
nand U8856 (N_8856,N_8053,N_8182);
or U8857 (N_8857,N_8219,N_8093);
xor U8858 (N_8858,N_8152,N_8087);
nand U8859 (N_8859,N_8320,N_8262);
xnor U8860 (N_8860,N_8042,N_8406);
xor U8861 (N_8861,N_8137,N_8239);
or U8862 (N_8862,N_8294,N_8434);
nor U8863 (N_8863,N_8224,N_8024);
or U8864 (N_8864,N_8188,N_8379);
and U8865 (N_8865,N_8301,N_8303);
or U8866 (N_8866,N_8471,N_8244);
or U8867 (N_8867,N_8433,N_8446);
or U8868 (N_8868,N_8174,N_8237);
xor U8869 (N_8869,N_8058,N_8282);
nand U8870 (N_8870,N_8338,N_8189);
nand U8871 (N_8871,N_8495,N_8358);
or U8872 (N_8872,N_8251,N_8029);
xnor U8873 (N_8873,N_8294,N_8499);
nand U8874 (N_8874,N_8311,N_8460);
nor U8875 (N_8875,N_8437,N_8430);
nand U8876 (N_8876,N_8184,N_8136);
nor U8877 (N_8877,N_8366,N_8092);
xnor U8878 (N_8878,N_8194,N_8148);
or U8879 (N_8879,N_8186,N_8085);
or U8880 (N_8880,N_8022,N_8130);
nand U8881 (N_8881,N_8344,N_8376);
xnor U8882 (N_8882,N_8344,N_8115);
and U8883 (N_8883,N_8241,N_8016);
and U8884 (N_8884,N_8044,N_8328);
xor U8885 (N_8885,N_8486,N_8255);
nor U8886 (N_8886,N_8431,N_8364);
xor U8887 (N_8887,N_8133,N_8459);
nor U8888 (N_8888,N_8178,N_8327);
xnor U8889 (N_8889,N_8314,N_8329);
xor U8890 (N_8890,N_8247,N_8280);
and U8891 (N_8891,N_8406,N_8005);
and U8892 (N_8892,N_8280,N_8184);
nor U8893 (N_8893,N_8073,N_8288);
xor U8894 (N_8894,N_8497,N_8333);
nand U8895 (N_8895,N_8350,N_8144);
nor U8896 (N_8896,N_8468,N_8365);
xor U8897 (N_8897,N_8169,N_8486);
nor U8898 (N_8898,N_8143,N_8247);
or U8899 (N_8899,N_8470,N_8473);
nor U8900 (N_8900,N_8338,N_8302);
xnor U8901 (N_8901,N_8174,N_8477);
xor U8902 (N_8902,N_8285,N_8332);
and U8903 (N_8903,N_8311,N_8456);
nand U8904 (N_8904,N_8375,N_8336);
nor U8905 (N_8905,N_8142,N_8153);
or U8906 (N_8906,N_8449,N_8285);
or U8907 (N_8907,N_8488,N_8494);
xor U8908 (N_8908,N_8416,N_8288);
or U8909 (N_8909,N_8251,N_8307);
and U8910 (N_8910,N_8342,N_8010);
and U8911 (N_8911,N_8177,N_8411);
or U8912 (N_8912,N_8327,N_8460);
or U8913 (N_8913,N_8405,N_8158);
or U8914 (N_8914,N_8113,N_8457);
and U8915 (N_8915,N_8239,N_8455);
and U8916 (N_8916,N_8167,N_8385);
xor U8917 (N_8917,N_8381,N_8249);
and U8918 (N_8918,N_8355,N_8332);
xor U8919 (N_8919,N_8478,N_8203);
or U8920 (N_8920,N_8112,N_8203);
xnor U8921 (N_8921,N_8301,N_8358);
xnor U8922 (N_8922,N_8091,N_8188);
xor U8923 (N_8923,N_8277,N_8007);
or U8924 (N_8924,N_8460,N_8477);
nand U8925 (N_8925,N_8463,N_8024);
xor U8926 (N_8926,N_8081,N_8208);
and U8927 (N_8927,N_8202,N_8095);
and U8928 (N_8928,N_8024,N_8276);
nand U8929 (N_8929,N_8175,N_8059);
or U8930 (N_8930,N_8021,N_8468);
and U8931 (N_8931,N_8382,N_8226);
nor U8932 (N_8932,N_8304,N_8164);
and U8933 (N_8933,N_8087,N_8310);
or U8934 (N_8934,N_8416,N_8449);
nand U8935 (N_8935,N_8433,N_8201);
and U8936 (N_8936,N_8193,N_8353);
nor U8937 (N_8937,N_8316,N_8020);
nand U8938 (N_8938,N_8317,N_8276);
xor U8939 (N_8939,N_8296,N_8100);
nor U8940 (N_8940,N_8184,N_8247);
xnor U8941 (N_8941,N_8382,N_8105);
nor U8942 (N_8942,N_8132,N_8231);
xnor U8943 (N_8943,N_8285,N_8036);
xnor U8944 (N_8944,N_8434,N_8112);
nor U8945 (N_8945,N_8448,N_8059);
nor U8946 (N_8946,N_8133,N_8053);
nor U8947 (N_8947,N_8036,N_8373);
or U8948 (N_8948,N_8343,N_8080);
and U8949 (N_8949,N_8495,N_8394);
or U8950 (N_8950,N_8112,N_8387);
xnor U8951 (N_8951,N_8083,N_8478);
or U8952 (N_8952,N_8204,N_8294);
xnor U8953 (N_8953,N_8402,N_8336);
xnor U8954 (N_8954,N_8426,N_8051);
nor U8955 (N_8955,N_8348,N_8269);
nand U8956 (N_8956,N_8427,N_8073);
and U8957 (N_8957,N_8051,N_8241);
xnor U8958 (N_8958,N_8452,N_8172);
xor U8959 (N_8959,N_8301,N_8282);
xor U8960 (N_8960,N_8099,N_8325);
nand U8961 (N_8961,N_8339,N_8183);
nor U8962 (N_8962,N_8248,N_8318);
and U8963 (N_8963,N_8234,N_8139);
nand U8964 (N_8964,N_8123,N_8145);
or U8965 (N_8965,N_8090,N_8126);
xnor U8966 (N_8966,N_8120,N_8109);
or U8967 (N_8967,N_8447,N_8428);
nand U8968 (N_8968,N_8063,N_8021);
and U8969 (N_8969,N_8222,N_8090);
xnor U8970 (N_8970,N_8029,N_8161);
xor U8971 (N_8971,N_8332,N_8258);
nand U8972 (N_8972,N_8002,N_8315);
nor U8973 (N_8973,N_8437,N_8294);
or U8974 (N_8974,N_8193,N_8477);
xnor U8975 (N_8975,N_8041,N_8223);
nand U8976 (N_8976,N_8104,N_8123);
nor U8977 (N_8977,N_8425,N_8058);
and U8978 (N_8978,N_8296,N_8095);
or U8979 (N_8979,N_8384,N_8255);
nand U8980 (N_8980,N_8413,N_8392);
nand U8981 (N_8981,N_8192,N_8204);
or U8982 (N_8982,N_8272,N_8361);
nand U8983 (N_8983,N_8397,N_8443);
or U8984 (N_8984,N_8196,N_8171);
nor U8985 (N_8985,N_8145,N_8143);
and U8986 (N_8986,N_8457,N_8126);
or U8987 (N_8987,N_8028,N_8424);
or U8988 (N_8988,N_8404,N_8346);
or U8989 (N_8989,N_8042,N_8495);
xor U8990 (N_8990,N_8152,N_8021);
xor U8991 (N_8991,N_8482,N_8384);
or U8992 (N_8992,N_8032,N_8218);
nand U8993 (N_8993,N_8494,N_8091);
or U8994 (N_8994,N_8168,N_8098);
nor U8995 (N_8995,N_8149,N_8326);
nand U8996 (N_8996,N_8334,N_8326);
nand U8997 (N_8997,N_8431,N_8343);
nor U8998 (N_8998,N_8244,N_8175);
xnor U8999 (N_8999,N_8057,N_8413);
nand U9000 (N_9000,N_8808,N_8801);
and U9001 (N_9001,N_8932,N_8735);
nand U9002 (N_9002,N_8928,N_8580);
nand U9003 (N_9003,N_8714,N_8552);
xor U9004 (N_9004,N_8763,N_8931);
nand U9005 (N_9005,N_8718,N_8600);
xnor U9006 (N_9006,N_8601,N_8972);
xnor U9007 (N_9007,N_8994,N_8539);
or U9008 (N_9008,N_8775,N_8665);
nand U9009 (N_9009,N_8686,N_8560);
xor U9010 (N_9010,N_8661,N_8833);
nand U9011 (N_9011,N_8620,N_8897);
and U9012 (N_9012,N_8992,N_8966);
nor U9013 (N_9013,N_8645,N_8762);
nand U9014 (N_9014,N_8811,N_8975);
nand U9015 (N_9015,N_8904,N_8985);
xor U9016 (N_9016,N_8802,N_8732);
nand U9017 (N_9017,N_8852,N_8671);
xor U9018 (N_9018,N_8835,N_8970);
xor U9019 (N_9019,N_8887,N_8940);
nor U9020 (N_9020,N_8923,N_8517);
nor U9021 (N_9021,N_8642,N_8984);
and U9022 (N_9022,N_8544,N_8838);
and U9023 (N_9023,N_8949,N_8871);
or U9024 (N_9024,N_8702,N_8860);
or U9025 (N_9025,N_8510,N_8537);
and U9026 (N_9026,N_8689,N_8706);
and U9027 (N_9027,N_8895,N_8562);
nand U9028 (N_9028,N_8595,N_8640);
and U9029 (N_9029,N_8857,N_8783);
nor U9030 (N_9030,N_8503,N_8694);
or U9031 (N_9031,N_8758,N_8893);
xnor U9032 (N_9032,N_8549,N_8800);
nand U9033 (N_9033,N_8813,N_8791);
xor U9034 (N_9034,N_8619,N_8742);
nand U9035 (N_9035,N_8959,N_8873);
and U9036 (N_9036,N_8778,N_8740);
nor U9037 (N_9037,N_8729,N_8824);
or U9038 (N_9038,N_8683,N_8961);
xor U9039 (N_9039,N_8710,N_8776);
nand U9040 (N_9040,N_8656,N_8715);
and U9041 (N_9041,N_8990,N_8607);
xor U9042 (N_9042,N_8896,N_8638);
nand U9043 (N_9043,N_8599,N_8588);
xnor U9044 (N_9044,N_8861,N_8789);
xnor U9045 (N_9045,N_8500,N_8854);
or U9046 (N_9046,N_8643,N_8713);
xnor U9047 (N_9047,N_8839,N_8846);
or U9048 (N_9048,N_8698,N_8799);
nand U9049 (N_9049,N_8945,N_8546);
or U9050 (N_9050,N_8681,N_8901);
nor U9051 (N_9051,N_8894,N_8612);
or U9052 (N_9052,N_8953,N_8613);
xnor U9053 (N_9053,N_8981,N_8616);
nand U9054 (N_9054,N_8830,N_8797);
nor U9055 (N_9055,N_8739,N_8991);
xor U9056 (N_9056,N_8687,N_8724);
and U9057 (N_9057,N_8964,N_8826);
nand U9058 (N_9058,N_8764,N_8850);
nand U9059 (N_9059,N_8529,N_8829);
nor U9060 (N_9060,N_8907,N_8520);
nand U9061 (N_9061,N_8809,N_8976);
or U9062 (N_9062,N_8633,N_8569);
nor U9063 (N_9063,N_8900,N_8880);
or U9064 (N_9064,N_8886,N_8551);
nand U9065 (N_9065,N_8627,N_8986);
nand U9066 (N_9066,N_8704,N_8963);
xnor U9067 (N_9067,N_8807,N_8818);
xnor U9068 (N_9068,N_8837,N_8636);
or U9069 (N_9069,N_8793,N_8559);
and U9070 (N_9070,N_8697,N_8618);
nand U9071 (N_9071,N_8617,N_8574);
or U9072 (N_9072,N_8507,N_8635);
nor U9073 (N_9073,N_8858,N_8744);
nand U9074 (N_9074,N_8676,N_8815);
nand U9075 (N_9075,N_8920,N_8624);
xnor U9076 (N_9076,N_8957,N_8805);
nand U9077 (N_9077,N_8667,N_8670);
xnor U9078 (N_9078,N_8557,N_8575);
nand U9079 (N_9079,N_8745,N_8980);
nand U9080 (N_9080,N_8699,N_8653);
nand U9081 (N_9081,N_8501,N_8812);
xor U9082 (N_9082,N_8918,N_8564);
or U9083 (N_9083,N_8622,N_8743);
or U9084 (N_9084,N_8626,N_8581);
xnor U9085 (N_9085,N_8936,N_8777);
nor U9086 (N_9086,N_8711,N_8673);
nand U9087 (N_9087,N_8505,N_8577);
nand U9088 (N_9088,N_8817,N_8662);
or U9089 (N_9089,N_8703,N_8696);
or U9090 (N_9090,N_8716,N_8870);
or U9091 (N_9091,N_8736,N_8658);
xnor U9092 (N_9092,N_8726,N_8543);
nand U9093 (N_9093,N_8891,N_8663);
or U9094 (N_9094,N_8593,N_8722);
nand U9095 (N_9095,N_8561,N_8610);
nor U9096 (N_9096,N_8605,N_8779);
or U9097 (N_9097,N_8965,N_8614);
nor U9098 (N_9098,N_8760,N_8885);
or U9099 (N_9099,N_8631,N_8921);
nor U9100 (N_9100,N_8769,N_8946);
xnor U9101 (N_9101,N_8563,N_8834);
xor U9102 (N_9102,N_8952,N_8590);
xnor U9103 (N_9103,N_8844,N_8608);
xor U9104 (N_9104,N_8664,N_8987);
and U9105 (N_9105,N_8705,N_8855);
nand U9106 (N_9106,N_8875,N_8524);
xnor U9107 (N_9107,N_8602,N_8848);
xor U9108 (N_9108,N_8866,N_8514);
and U9109 (N_9109,N_8814,N_8788);
nand U9110 (N_9110,N_8504,N_8721);
xnor U9111 (N_9111,N_8556,N_8910);
xor U9112 (N_9112,N_8578,N_8916);
nand U9113 (N_9113,N_8816,N_8655);
nor U9114 (N_9114,N_8755,N_8948);
and U9115 (N_9115,N_8541,N_8565);
xor U9116 (N_9116,N_8795,N_8958);
xor U9117 (N_9117,N_8765,N_8822);
or U9118 (N_9118,N_8749,N_8516);
nand U9119 (N_9119,N_8538,N_8908);
or U9120 (N_9120,N_8934,N_8584);
nand U9121 (N_9121,N_8840,N_8652);
nand U9122 (N_9122,N_8892,N_8654);
nand U9123 (N_9123,N_8634,N_8604);
or U9124 (N_9124,N_8796,N_8862);
and U9125 (N_9125,N_8935,N_8585);
xnor U9126 (N_9126,N_8929,N_8682);
and U9127 (N_9127,N_8913,N_8508);
nand U9128 (N_9128,N_8869,N_8956);
or U9129 (N_9129,N_8821,N_8511);
nand U9130 (N_9130,N_8919,N_8877);
nor U9131 (N_9131,N_8629,N_8810);
and U9132 (N_9132,N_8917,N_8962);
or U9133 (N_9133,N_8679,N_8864);
or U9134 (N_9134,N_8554,N_8926);
nor U9135 (N_9135,N_8521,N_8576);
nor U9136 (N_9136,N_8725,N_8641);
nor U9137 (N_9137,N_8836,N_8573);
nand U9138 (N_9138,N_8941,N_8659);
nor U9139 (N_9139,N_8657,N_8847);
xor U9140 (N_9140,N_8566,N_8727);
nor U9141 (N_9141,N_8644,N_8666);
and U9142 (N_9142,N_8794,N_8933);
nor U9143 (N_9143,N_8693,N_8533);
nand U9144 (N_9144,N_8648,N_8567);
or U9145 (N_9145,N_8609,N_8526);
nand U9146 (N_9146,N_8519,N_8823);
or U9147 (N_9147,N_8555,N_8773);
nor U9148 (N_9148,N_8688,N_8939);
or U9149 (N_9149,N_8995,N_8603);
xnor U9150 (N_9150,N_8832,N_8872);
or U9151 (N_9151,N_8954,N_8781);
xnor U9152 (N_9152,N_8540,N_8571);
xor U9153 (N_9153,N_8730,N_8632);
nand U9154 (N_9154,N_8979,N_8591);
and U9155 (N_9155,N_8927,N_8884);
and U9156 (N_9156,N_8532,N_8771);
nor U9157 (N_9157,N_8868,N_8733);
xor U9158 (N_9158,N_8903,N_8579);
xor U9159 (N_9159,N_8530,N_8598);
nor U9160 (N_9160,N_8851,N_8525);
nand U9161 (N_9161,N_8534,N_8512);
and U9162 (N_9162,N_8768,N_8915);
nor U9163 (N_9163,N_8867,N_8660);
or U9164 (N_9164,N_8942,N_8842);
nand U9165 (N_9165,N_8523,N_8787);
nand U9166 (N_9166,N_8951,N_8649);
nor U9167 (N_9167,N_8905,N_8938);
nand U9168 (N_9168,N_8675,N_8708);
xor U9169 (N_9169,N_8820,N_8754);
nor U9170 (N_9170,N_8527,N_8888);
nor U9171 (N_9171,N_8582,N_8535);
or U9172 (N_9172,N_8761,N_8882);
or U9173 (N_9173,N_8784,N_8678);
nand U9174 (N_9174,N_8700,N_8912);
nor U9175 (N_9175,N_8930,N_8684);
or U9176 (N_9176,N_8606,N_8651);
nand U9177 (N_9177,N_8752,N_8690);
xnor U9178 (N_9178,N_8922,N_8738);
nor U9179 (N_9179,N_8548,N_8828);
and U9180 (N_9180,N_8717,N_8757);
or U9181 (N_9181,N_8843,N_8906);
or U9182 (N_9182,N_8669,N_8550);
nor U9183 (N_9183,N_8782,N_8513);
and U9184 (N_9184,N_8630,N_8691);
and U9185 (N_9185,N_8914,N_8943);
xnor U9186 (N_9186,N_8547,N_8774);
xor U9187 (N_9187,N_8672,N_8583);
or U9188 (N_9188,N_8748,N_8746);
nor U9189 (N_9189,N_8586,N_8879);
or U9190 (N_9190,N_8753,N_8646);
xor U9191 (N_9191,N_8845,N_8647);
and U9192 (N_9192,N_8621,N_8924);
nor U9193 (N_9193,N_8998,N_8719);
nand U9194 (N_9194,N_8874,N_8841);
or U9195 (N_9195,N_8728,N_8996);
nand U9196 (N_9196,N_8925,N_8751);
nand U9197 (N_9197,N_8780,N_8883);
and U9198 (N_9198,N_8955,N_8960);
and U9199 (N_9199,N_8518,N_8989);
nor U9200 (N_9200,N_8701,N_8737);
and U9201 (N_9201,N_8685,N_8709);
nor U9202 (N_9202,N_8937,N_8568);
xnor U9203 (N_9203,N_8853,N_8950);
xor U9204 (N_9204,N_8531,N_8899);
or U9205 (N_9205,N_8878,N_8712);
and U9206 (N_9206,N_8628,N_8509);
xnor U9207 (N_9207,N_8973,N_8756);
and U9208 (N_9208,N_8637,N_8790);
and U9209 (N_9209,N_8890,N_8993);
nand U9210 (N_9210,N_8997,N_8515);
nand U9211 (N_9211,N_8785,N_8589);
and U9212 (N_9212,N_8572,N_8819);
xor U9213 (N_9213,N_8977,N_8898);
nand U9214 (N_9214,N_8881,N_8982);
or U9215 (N_9215,N_8969,N_8902);
nor U9216 (N_9216,N_8831,N_8741);
nor U9217 (N_9217,N_8911,N_8570);
nand U9218 (N_9218,N_8798,N_8720);
xor U9219 (N_9219,N_8806,N_8971);
nand U9220 (N_9220,N_8772,N_8974);
and U9221 (N_9221,N_8506,N_8978);
or U9222 (N_9222,N_8792,N_8623);
nand U9223 (N_9223,N_8587,N_8750);
or U9224 (N_9224,N_8849,N_8594);
xnor U9225 (N_9225,N_8804,N_8889);
xor U9226 (N_9226,N_8786,N_8766);
nor U9227 (N_9227,N_8639,N_8502);
nor U9228 (N_9228,N_8692,N_8947);
nor U9229 (N_9229,N_8859,N_8650);
xnor U9230 (N_9230,N_8967,N_8677);
or U9231 (N_9231,N_8759,N_8983);
and U9232 (N_9232,N_8856,N_8770);
nor U9233 (N_9233,N_8536,N_8825);
and U9234 (N_9234,N_8597,N_8734);
nand U9235 (N_9235,N_8988,N_8723);
nand U9236 (N_9236,N_8625,N_8747);
or U9237 (N_9237,N_8522,N_8528);
nor U9238 (N_9238,N_8999,N_8592);
xnor U9239 (N_9239,N_8545,N_8767);
and U9240 (N_9240,N_8596,N_8707);
nor U9241 (N_9241,N_8909,N_8863);
nand U9242 (N_9242,N_8558,N_8542);
nor U9243 (N_9243,N_8668,N_8553);
xnor U9244 (N_9244,N_8944,N_8803);
nand U9245 (N_9245,N_8968,N_8876);
and U9246 (N_9246,N_8827,N_8865);
and U9247 (N_9247,N_8695,N_8611);
nand U9248 (N_9248,N_8731,N_8680);
and U9249 (N_9249,N_8615,N_8674);
nand U9250 (N_9250,N_8971,N_8532);
or U9251 (N_9251,N_8847,N_8908);
xor U9252 (N_9252,N_8847,N_8606);
nand U9253 (N_9253,N_8922,N_8747);
nor U9254 (N_9254,N_8729,N_8664);
nand U9255 (N_9255,N_8758,N_8768);
or U9256 (N_9256,N_8996,N_8670);
or U9257 (N_9257,N_8990,N_8796);
nor U9258 (N_9258,N_8727,N_8638);
and U9259 (N_9259,N_8668,N_8771);
xor U9260 (N_9260,N_8645,N_8952);
or U9261 (N_9261,N_8700,N_8863);
nor U9262 (N_9262,N_8735,N_8617);
or U9263 (N_9263,N_8962,N_8843);
or U9264 (N_9264,N_8694,N_8650);
and U9265 (N_9265,N_8528,N_8962);
nand U9266 (N_9266,N_8841,N_8772);
xor U9267 (N_9267,N_8972,N_8610);
and U9268 (N_9268,N_8537,N_8793);
or U9269 (N_9269,N_8833,N_8518);
xor U9270 (N_9270,N_8780,N_8629);
nand U9271 (N_9271,N_8644,N_8770);
and U9272 (N_9272,N_8760,N_8944);
nor U9273 (N_9273,N_8648,N_8957);
nand U9274 (N_9274,N_8834,N_8523);
xor U9275 (N_9275,N_8677,N_8769);
nor U9276 (N_9276,N_8549,N_8668);
nand U9277 (N_9277,N_8714,N_8776);
and U9278 (N_9278,N_8968,N_8879);
or U9279 (N_9279,N_8867,N_8577);
nor U9280 (N_9280,N_8864,N_8759);
xor U9281 (N_9281,N_8925,N_8953);
or U9282 (N_9282,N_8684,N_8562);
or U9283 (N_9283,N_8822,N_8635);
or U9284 (N_9284,N_8911,N_8669);
and U9285 (N_9285,N_8807,N_8946);
or U9286 (N_9286,N_8973,N_8552);
or U9287 (N_9287,N_8730,N_8706);
and U9288 (N_9288,N_8755,N_8903);
nand U9289 (N_9289,N_8562,N_8510);
nor U9290 (N_9290,N_8957,N_8636);
nor U9291 (N_9291,N_8731,N_8833);
xnor U9292 (N_9292,N_8622,N_8529);
or U9293 (N_9293,N_8630,N_8509);
xnor U9294 (N_9294,N_8575,N_8888);
xnor U9295 (N_9295,N_8505,N_8581);
or U9296 (N_9296,N_8935,N_8793);
nand U9297 (N_9297,N_8606,N_8560);
nand U9298 (N_9298,N_8709,N_8699);
nor U9299 (N_9299,N_8567,N_8800);
nor U9300 (N_9300,N_8821,N_8561);
or U9301 (N_9301,N_8964,N_8665);
and U9302 (N_9302,N_8834,N_8733);
xnor U9303 (N_9303,N_8719,N_8665);
xnor U9304 (N_9304,N_8821,N_8749);
or U9305 (N_9305,N_8589,N_8845);
or U9306 (N_9306,N_8662,N_8549);
and U9307 (N_9307,N_8594,N_8855);
and U9308 (N_9308,N_8761,N_8583);
nor U9309 (N_9309,N_8843,N_8733);
or U9310 (N_9310,N_8993,N_8514);
or U9311 (N_9311,N_8692,N_8962);
nand U9312 (N_9312,N_8738,N_8657);
nor U9313 (N_9313,N_8765,N_8850);
and U9314 (N_9314,N_8673,N_8585);
xor U9315 (N_9315,N_8935,N_8577);
nand U9316 (N_9316,N_8817,N_8807);
nand U9317 (N_9317,N_8727,N_8740);
xor U9318 (N_9318,N_8928,N_8617);
and U9319 (N_9319,N_8845,N_8548);
or U9320 (N_9320,N_8916,N_8855);
and U9321 (N_9321,N_8991,N_8607);
and U9322 (N_9322,N_8864,N_8676);
xnor U9323 (N_9323,N_8727,N_8524);
xnor U9324 (N_9324,N_8965,N_8774);
xnor U9325 (N_9325,N_8983,N_8801);
and U9326 (N_9326,N_8641,N_8813);
xor U9327 (N_9327,N_8712,N_8834);
xnor U9328 (N_9328,N_8967,N_8674);
and U9329 (N_9329,N_8639,N_8525);
nand U9330 (N_9330,N_8861,N_8988);
nor U9331 (N_9331,N_8887,N_8892);
and U9332 (N_9332,N_8566,N_8759);
nor U9333 (N_9333,N_8888,N_8639);
nand U9334 (N_9334,N_8898,N_8895);
and U9335 (N_9335,N_8924,N_8906);
and U9336 (N_9336,N_8809,N_8871);
or U9337 (N_9337,N_8645,N_8854);
or U9338 (N_9338,N_8686,N_8715);
xnor U9339 (N_9339,N_8966,N_8749);
nand U9340 (N_9340,N_8849,N_8651);
xor U9341 (N_9341,N_8673,N_8565);
and U9342 (N_9342,N_8519,N_8597);
xnor U9343 (N_9343,N_8767,N_8607);
or U9344 (N_9344,N_8915,N_8606);
nand U9345 (N_9345,N_8627,N_8837);
nor U9346 (N_9346,N_8759,N_8672);
or U9347 (N_9347,N_8977,N_8891);
nor U9348 (N_9348,N_8981,N_8958);
or U9349 (N_9349,N_8795,N_8618);
nand U9350 (N_9350,N_8917,N_8870);
nand U9351 (N_9351,N_8809,N_8995);
nor U9352 (N_9352,N_8712,N_8793);
or U9353 (N_9353,N_8718,N_8842);
nor U9354 (N_9354,N_8997,N_8791);
and U9355 (N_9355,N_8755,N_8797);
and U9356 (N_9356,N_8709,N_8842);
nor U9357 (N_9357,N_8667,N_8801);
or U9358 (N_9358,N_8730,N_8997);
nand U9359 (N_9359,N_8924,N_8758);
and U9360 (N_9360,N_8512,N_8786);
xor U9361 (N_9361,N_8896,N_8888);
and U9362 (N_9362,N_8929,N_8983);
xnor U9363 (N_9363,N_8502,N_8771);
xnor U9364 (N_9364,N_8889,N_8657);
xor U9365 (N_9365,N_8794,N_8584);
nand U9366 (N_9366,N_8541,N_8967);
and U9367 (N_9367,N_8652,N_8555);
xnor U9368 (N_9368,N_8539,N_8721);
nand U9369 (N_9369,N_8584,N_8883);
or U9370 (N_9370,N_8863,N_8666);
xor U9371 (N_9371,N_8964,N_8644);
or U9372 (N_9372,N_8782,N_8718);
nor U9373 (N_9373,N_8526,N_8814);
xor U9374 (N_9374,N_8627,N_8848);
and U9375 (N_9375,N_8764,N_8959);
or U9376 (N_9376,N_8616,N_8697);
xor U9377 (N_9377,N_8609,N_8568);
nand U9378 (N_9378,N_8637,N_8676);
or U9379 (N_9379,N_8890,N_8635);
nand U9380 (N_9380,N_8550,N_8956);
or U9381 (N_9381,N_8651,N_8856);
or U9382 (N_9382,N_8529,N_8715);
nand U9383 (N_9383,N_8816,N_8715);
xor U9384 (N_9384,N_8845,N_8524);
and U9385 (N_9385,N_8653,N_8792);
or U9386 (N_9386,N_8711,N_8597);
and U9387 (N_9387,N_8726,N_8988);
and U9388 (N_9388,N_8946,N_8697);
and U9389 (N_9389,N_8695,N_8712);
and U9390 (N_9390,N_8760,N_8656);
nand U9391 (N_9391,N_8883,N_8857);
nor U9392 (N_9392,N_8740,N_8738);
nand U9393 (N_9393,N_8697,N_8832);
or U9394 (N_9394,N_8915,N_8842);
xnor U9395 (N_9395,N_8514,N_8688);
nand U9396 (N_9396,N_8936,N_8952);
nor U9397 (N_9397,N_8665,N_8836);
xnor U9398 (N_9398,N_8966,N_8714);
and U9399 (N_9399,N_8627,N_8637);
and U9400 (N_9400,N_8678,N_8570);
xor U9401 (N_9401,N_8962,N_8564);
xor U9402 (N_9402,N_8834,N_8852);
and U9403 (N_9403,N_8898,N_8999);
xnor U9404 (N_9404,N_8966,N_8623);
xnor U9405 (N_9405,N_8612,N_8760);
or U9406 (N_9406,N_8619,N_8671);
xnor U9407 (N_9407,N_8924,N_8978);
xor U9408 (N_9408,N_8547,N_8708);
nor U9409 (N_9409,N_8535,N_8521);
nand U9410 (N_9410,N_8811,N_8531);
and U9411 (N_9411,N_8946,N_8688);
and U9412 (N_9412,N_8740,N_8969);
nor U9413 (N_9413,N_8840,N_8667);
xnor U9414 (N_9414,N_8891,N_8658);
xnor U9415 (N_9415,N_8827,N_8999);
and U9416 (N_9416,N_8538,N_8854);
nor U9417 (N_9417,N_8650,N_8524);
or U9418 (N_9418,N_8595,N_8920);
nor U9419 (N_9419,N_8534,N_8674);
and U9420 (N_9420,N_8913,N_8673);
nand U9421 (N_9421,N_8780,N_8753);
and U9422 (N_9422,N_8964,N_8806);
xor U9423 (N_9423,N_8914,N_8696);
and U9424 (N_9424,N_8672,N_8529);
nor U9425 (N_9425,N_8863,N_8735);
xor U9426 (N_9426,N_8565,N_8944);
or U9427 (N_9427,N_8741,N_8819);
or U9428 (N_9428,N_8827,N_8725);
xor U9429 (N_9429,N_8708,N_8743);
xor U9430 (N_9430,N_8792,N_8764);
nand U9431 (N_9431,N_8582,N_8506);
xor U9432 (N_9432,N_8806,N_8976);
and U9433 (N_9433,N_8600,N_8865);
or U9434 (N_9434,N_8533,N_8819);
xor U9435 (N_9435,N_8816,N_8569);
nor U9436 (N_9436,N_8799,N_8873);
and U9437 (N_9437,N_8812,N_8598);
and U9438 (N_9438,N_8874,N_8677);
and U9439 (N_9439,N_8881,N_8560);
xnor U9440 (N_9440,N_8588,N_8795);
or U9441 (N_9441,N_8537,N_8844);
and U9442 (N_9442,N_8765,N_8702);
nand U9443 (N_9443,N_8932,N_8784);
nor U9444 (N_9444,N_8823,N_8761);
and U9445 (N_9445,N_8661,N_8950);
or U9446 (N_9446,N_8651,N_8590);
or U9447 (N_9447,N_8947,N_8772);
nor U9448 (N_9448,N_8819,N_8573);
xor U9449 (N_9449,N_8702,N_8970);
nor U9450 (N_9450,N_8980,N_8964);
nor U9451 (N_9451,N_8516,N_8813);
nand U9452 (N_9452,N_8552,N_8528);
xor U9453 (N_9453,N_8938,N_8917);
nand U9454 (N_9454,N_8786,N_8993);
or U9455 (N_9455,N_8921,N_8748);
nor U9456 (N_9456,N_8594,N_8683);
xnor U9457 (N_9457,N_8762,N_8787);
xor U9458 (N_9458,N_8718,N_8964);
or U9459 (N_9459,N_8895,N_8877);
xor U9460 (N_9460,N_8538,N_8824);
or U9461 (N_9461,N_8626,N_8906);
and U9462 (N_9462,N_8929,N_8579);
or U9463 (N_9463,N_8934,N_8731);
and U9464 (N_9464,N_8930,N_8960);
xor U9465 (N_9465,N_8652,N_8660);
nor U9466 (N_9466,N_8617,N_8892);
xnor U9467 (N_9467,N_8855,N_8558);
or U9468 (N_9468,N_8566,N_8588);
or U9469 (N_9469,N_8600,N_8572);
or U9470 (N_9470,N_8569,N_8972);
nand U9471 (N_9471,N_8753,N_8741);
xnor U9472 (N_9472,N_8823,N_8624);
nor U9473 (N_9473,N_8539,N_8821);
and U9474 (N_9474,N_8767,N_8952);
nor U9475 (N_9475,N_8921,N_8718);
and U9476 (N_9476,N_8548,N_8730);
nand U9477 (N_9477,N_8546,N_8703);
nand U9478 (N_9478,N_8737,N_8789);
xor U9479 (N_9479,N_8578,N_8624);
xor U9480 (N_9480,N_8720,N_8690);
and U9481 (N_9481,N_8782,N_8857);
and U9482 (N_9482,N_8865,N_8832);
nor U9483 (N_9483,N_8930,N_8500);
or U9484 (N_9484,N_8644,N_8534);
and U9485 (N_9485,N_8960,N_8904);
nand U9486 (N_9486,N_8555,N_8780);
nand U9487 (N_9487,N_8664,N_8931);
and U9488 (N_9488,N_8689,N_8672);
or U9489 (N_9489,N_8567,N_8883);
xnor U9490 (N_9490,N_8922,N_8915);
or U9491 (N_9491,N_8795,N_8938);
nor U9492 (N_9492,N_8575,N_8518);
and U9493 (N_9493,N_8686,N_8776);
nand U9494 (N_9494,N_8939,N_8787);
nand U9495 (N_9495,N_8557,N_8953);
or U9496 (N_9496,N_8941,N_8917);
xor U9497 (N_9497,N_8569,N_8564);
or U9498 (N_9498,N_8831,N_8573);
or U9499 (N_9499,N_8868,N_8580);
xor U9500 (N_9500,N_9361,N_9385);
nor U9501 (N_9501,N_9312,N_9037);
nor U9502 (N_9502,N_9131,N_9046);
nor U9503 (N_9503,N_9396,N_9486);
or U9504 (N_9504,N_9042,N_9337);
nor U9505 (N_9505,N_9184,N_9422);
xor U9506 (N_9506,N_9241,N_9217);
nand U9507 (N_9507,N_9034,N_9243);
or U9508 (N_9508,N_9237,N_9466);
nor U9509 (N_9509,N_9317,N_9149);
nand U9510 (N_9510,N_9225,N_9138);
nor U9511 (N_9511,N_9137,N_9366);
or U9512 (N_9512,N_9354,N_9006);
nor U9513 (N_9513,N_9259,N_9304);
nor U9514 (N_9514,N_9438,N_9244);
or U9515 (N_9515,N_9093,N_9356);
nand U9516 (N_9516,N_9120,N_9004);
nand U9517 (N_9517,N_9443,N_9347);
and U9518 (N_9518,N_9122,N_9095);
and U9519 (N_9519,N_9033,N_9088);
or U9520 (N_9520,N_9160,N_9276);
nand U9521 (N_9521,N_9079,N_9104);
nor U9522 (N_9522,N_9399,N_9091);
and U9523 (N_9523,N_9447,N_9235);
and U9524 (N_9524,N_9305,N_9099);
or U9525 (N_9525,N_9424,N_9287);
nand U9526 (N_9526,N_9472,N_9448);
or U9527 (N_9527,N_9142,N_9014);
nand U9528 (N_9528,N_9064,N_9412);
nor U9529 (N_9529,N_9446,N_9417);
xnor U9530 (N_9530,N_9487,N_9303);
nand U9531 (N_9531,N_9152,N_9496);
and U9532 (N_9532,N_9299,N_9389);
and U9533 (N_9533,N_9023,N_9169);
xor U9534 (N_9534,N_9136,N_9199);
xor U9535 (N_9535,N_9035,N_9163);
nand U9536 (N_9536,N_9094,N_9031);
nor U9537 (N_9537,N_9390,N_9344);
xor U9538 (N_9538,N_9076,N_9371);
xnor U9539 (N_9539,N_9269,N_9148);
and U9540 (N_9540,N_9436,N_9231);
xor U9541 (N_9541,N_9271,N_9154);
xor U9542 (N_9542,N_9408,N_9039);
or U9543 (N_9543,N_9192,N_9497);
and U9544 (N_9544,N_9156,N_9189);
nand U9545 (N_9545,N_9464,N_9194);
nand U9546 (N_9546,N_9100,N_9202);
xor U9547 (N_9547,N_9043,N_9196);
nor U9548 (N_9548,N_9092,N_9162);
and U9549 (N_9549,N_9207,N_9261);
or U9550 (N_9550,N_9198,N_9461);
xnor U9551 (N_9551,N_9368,N_9178);
or U9552 (N_9552,N_9116,N_9168);
nor U9553 (N_9553,N_9020,N_9059);
nor U9554 (N_9554,N_9286,N_9260);
and U9555 (N_9555,N_9313,N_9330);
and U9556 (N_9556,N_9378,N_9019);
nor U9557 (N_9557,N_9326,N_9352);
and U9558 (N_9558,N_9074,N_9265);
and U9559 (N_9559,N_9255,N_9355);
xor U9560 (N_9560,N_9161,N_9423);
xnor U9561 (N_9561,N_9258,N_9082);
nand U9562 (N_9562,N_9405,N_9103);
nor U9563 (N_9563,N_9011,N_9348);
nor U9564 (N_9564,N_9343,N_9444);
and U9565 (N_9565,N_9476,N_9054);
nand U9566 (N_9566,N_9346,N_9084);
or U9567 (N_9567,N_9146,N_9197);
nand U9568 (N_9568,N_9324,N_9377);
nor U9569 (N_9569,N_9065,N_9195);
and U9570 (N_9570,N_9188,N_9167);
nor U9571 (N_9571,N_9185,N_9016);
and U9572 (N_9572,N_9278,N_9058);
and U9573 (N_9573,N_9205,N_9239);
or U9574 (N_9574,N_9393,N_9481);
xnor U9575 (N_9575,N_9489,N_9052);
or U9576 (N_9576,N_9395,N_9310);
xor U9577 (N_9577,N_9294,N_9402);
or U9578 (N_9578,N_9426,N_9248);
and U9579 (N_9579,N_9308,N_9249);
nand U9580 (N_9580,N_9290,N_9097);
and U9581 (N_9581,N_9349,N_9441);
nand U9582 (N_9582,N_9381,N_9157);
and U9583 (N_9583,N_9080,N_9172);
and U9584 (N_9584,N_9204,N_9328);
or U9585 (N_9585,N_9108,N_9460);
nand U9586 (N_9586,N_9158,N_9485);
nand U9587 (N_9587,N_9075,N_9141);
xor U9588 (N_9588,N_9338,N_9070);
and U9589 (N_9589,N_9191,N_9367);
or U9590 (N_9590,N_9474,N_9021);
xor U9591 (N_9591,N_9109,N_9482);
xor U9592 (N_9592,N_9250,N_9270);
nand U9593 (N_9593,N_9127,N_9289);
nor U9594 (N_9594,N_9442,N_9106);
or U9595 (N_9595,N_9041,N_9434);
or U9596 (N_9596,N_9087,N_9362);
nor U9597 (N_9597,N_9220,N_9471);
or U9598 (N_9598,N_9394,N_9325);
and U9599 (N_9599,N_9242,N_9200);
and U9600 (N_9600,N_9067,N_9047);
or U9601 (N_9601,N_9245,N_9266);
nor U9602 (N_9602,N_9277,N_9000);
xor U9603 (N_9603,N_9114,N_9430);
nor U9604 (N_9604,N_9263,N_9421);
nor U9605 (N_9605,N_9085,N_9128);
nand U9606 (N_9606,N_9425,N_9469);
nand U9607 (N_9607,N_9036,N_9003);
or U9608 (N_9608,N_9063,N_9272);
nand U9609 (N_9609,N_9057,N_9468);
and U9610 (N_9610,N_9360,N_9044);
xor U9611 (N_9611,N_9240,N_9340);
or U9612 (N_9612,N_9323,N_9224);
or U9613 (N_9613,N_9236,N_9397);
or U9614 (N_9614,N_9038,N_9073);
nand U9615 (N_9615,N_9401,N_9359);
nor U9616 (N_9616,N_9384,N_9267);
and U9617 (N_9617,N_9252,N_9314);
xor U9618 (N_9618,N_9414,N_9339);
nor U9619 (N_9619,N_9130,N_9180);
or U9620 (N_9620,N_9433,N_9013);
nor U9621 (N_9621,N_9211,N_9322);
or U9622 (N_9622,N_9400,N_9246);
xnor U9623 (N_9623,N_9222,N_9372);
and U9624 (N_9624,N_9418,N_9380);
xor U9625 (N_9625,N_9420,N_9451);
and U9626 (N_9626,N_9379,N_9210);
xnor U9627 (N_9627,N_9253,N_9432);
nor U9628 (N_9628,N_9415,N_9370);
nand U9629 (N_9629,N_9427,N_9483);
nand U9630 (N_9630,N_9488,N_9435);
and U9631 (N_9631,N_9090,N_9437);
nand U9632 (N_9632,N_9297,N_9111);
and U9633 (N_9633,N_9445,N_9293);
or U9634 (N_9634,N_9376,N_9140);
and U9635 (N_9635,N_9144,N_9134);
nor U9636 (N_9636,N_9077,N_9386);
nand U9637 (N_9637,N_9457,N_9369);
or U9638 (N_9638,N_9030,N_9186);
nand U9639 (N_9639,N_9493,N_9391);
nand U9640 (N_9640,N_9072,N_9238);
or U9641 (N_9641,N_9285,N_9176);
nor U9642 (N_9642,N_9406,N_9086);
nand U9643 (N_9643,N_9153,N_9350);
or U9644 (N_9644,N_9398,N_9212);
or U9645 (N_9645,N_9478,N_9459);
xnor U9646 (N_9646,N_9281,N_9101);
nand U9647 (N_9647,N_9491,N_9334);
or U9648 (N_9648,N_9123,N_9280);
nor U9649 (N_9649,N_9268,N_9319);
xor U9650 (N_9650,N_9327,N_9190);
and U9651 (N_9651,N_9066,N_9440);
xnor U9652 (N_9652,N_9477,N_9419);
or U9653 (N_9653,N_9320,N_9494);
or U9654 (N_9654,N_9193,N_9115);
nand U9655 (N_9655,N_9335,N_9392);
nor U9656 (N_9656,N_9133,N_9129);
xnor U9657 (N_9657,N_9264,N_9139);
nand U9658 (N_9658,N_9135,N_9365);
nand U9659 (N_9659,N_9221,N_9292);
xnor U9660 (N_9660,N_9300,N_9452);
or U9661 (N_9661,N_9179,N_9201);
nand U9662 (N_9662,N_9456,N_9404);
nand U9663 (N_9663,N_9007,N_9208);
xnor U9664 (N_9664,N_9490,N_9216);
nand U9665 (N_9665,N_9467,N_9032);
nand U9666 (N_9666,N_9040,N_9357);
and U9667 (N_9667,N_9470,N_9229);
nor U9668 (N_9668,N_9341,N_9022);
xor U9669 (N_9669,N_9219,N_9045);
or U9670 (N_9670,N_9410,N_9015);
xor U9671 (N_9671,N_9175,N_9251);
and U9672 (N_9672,N_9449,N_9454);
nand U9673 (N_9673,N_9089,N_9453);
xor U9674 (N_9674,N_9413,N_9049);
nand U9675 (N_9675,N_9177,N_9403);
nor U9676 (N_9676,N_9318,N_9098);
and U9677 (N_9677,N_9048,N_9256);
or U9678 (N_9678,N_9060,N_9078);
or U9679 (N_9679,N_9288,N_9273);
nor U9680 (N_9680,N_9055,N_9455);
or U9681 (N_9681,N_9374,N_9150);
or U9682 (N_9682,N_9302,N_9105);
nor U9683 (N_9683,N_9363,N_9121);
or U9684 (N_9684,N_9387,N_9068);
and U9685 (N_9685,N_9017,N_9375);
xnor U9686 (N_9686,N_9247,N_9409);
nand U9687 (N_9687,N_9351,N_9462);
xnor U9688 (N_9688,N_9155,N_9183);
nor U9689 (N_9689,N_9234,N_9069);
xnor U9690 (N_9690,N_9126,N_9062);
nor U9691 (N_9691,N_9203,N_9254);
xor U9692 (N_9692,N_9336,N_9102);
or U9693 (N_9693,N_9206,N_9001);
nand U9694 (N_9694,N_9479,N_9275);
and U9695 (N_9695,N_9024,N_9051);
nor U9696 (N_9696,N_9232,N_9315);
nor U9697 (N_9697,N_9182,N_9473);
xor U9698 (N_9698,N_9495,N_9307);
nor U9699 (N_9699,N_9475,N_9373);
nor U9700 (N_9700,N_9429,N_9165);
nand U9701 (N_9701,N_9009,N_9223);
and U9702 (N_9702,N_9113,N_9056);
and U9703 (N_9703,N_9416,N_9284);
xor U9704 (N_9704,N_9081,N_9333);
xnor U9705 (N_9705,N_9342,N_9458);
xor U9706 (N_9706,N_9439,N_9383);
xnor U9707 (N_9707,N_9226,N_9110);
nand U9708 (N_9708,N_9181,N_9257);
nand U9709 (N_9709,N_9029,N_9159);
or U9710 (N_9710,N_9164,N_9061);
nand U9711 (N_9711,N_9331,N_9227);
nor U9712 (N_9712,N_9311,N_9214);
and U9713 (N_9713,N_9262,N_9296);
nand U9714 (N_9714,N_9018,N_9301);
and U9715 (N_9715,N_9010,N_9005);
and U9716 (N_9716,N_9118,N_9213);
xnor U9717 (N_9717,N_9450,N_9145);
nand U9718 (N_9718,N_9283,N_9364);
or U9719 (N_9719,N_9124,N_9465);
or U9720 (N_9720,N_9050,N_9187);
nor U9721 (N_9721,N_9492,N_9431);
and U9722 (N_9722,N_9008,N_9166);
nand U9723 (N_9723,N_9174,N_9096);
nor U9724 (N_9724,N_9358,N_9480);
nor U9725 (N_9725,N_9332,N_9295);
xor U9726 (N_9726,N_9002,N_9025);
nand U9727 (N_9727,N_9228,N_9012);
and U9728 (N_9728,N_9298,N_9053);
or U9729 (N_9729,N_9388,N_9027);
xnor U9730 (N_9730,N_9143,N_9306);
or U9731 (N_9731,N_9071,N_9215);
or U9732 (N_9732,N_9499,N_9233);
xor U9733 (N_9733,N_9484,N_9321);
nand U9734 (N_9734,N_9498,N_9026);
or U9735 (N_9735,N_9463,N_9083);
and U9736 (N_9736,N_9147,N_9230);
xor U9737 (N_9737,N_9353,N_9382);
nor U9738 (N_9738,N_9170,N_9282);
and U9739 (N_9739,N_9428,N_9107);
and U9740 (N_9740,N_9291,N_9125);
or U9741 (N_9741,N_9279,N_9171);
xor U9742 (N_9742,N_9132,N_9274);
nand U9743 (N_9743,N_9407,N_9209);
and U9744 (N_9744,N_9119,N_9151);
and U9745 (N_9745,N_9218,N_9411);
or U9746 (N_9746,N_9316,N_9309);
xnor U9747 (N_9747,N_9173,N_9112);
xnor U9748 (N_9748,N_9117,N_9329);
nand U9749 (N_9749,N_9028,N_9345);
nand U9750 (N_9750,N_9090,N_9343);
nand U9751 (N_9751,N_9394,N_9310);
xnor U9752 (N_9752,N_9078,N_9279);
or U9753 (N_9753,N_9154,N_9058);
xor U9754 (N_9754,N_9146,N_9177);
and U9755 (N_9755,N_9030,N_9157);
and U9756 (N_9756,N_9156,N_9336);
and U9757 (N_9757,N_9468,N_9269);
nand U9758 (N_9758,N_9478,N_9237);
and U9759 (N_9759,N_9480,N_9426);
or U9760 (N_9760,N_9026,N_9188);
or U9761 (N_9761,N_9135,N_9486);
or U9762 (N_9762,N_9050,N_9192);
or U9763 (N_9763,N_9170,N_9476);
nand U9764 (N_9764,N_9124,N_9417);
nor U9765 (N_9765,N_9005,N_9375);
xor U9766 (N_9766,N_9427,N_9133);
nand U9767 (N_9767,N_9316,N_9116);
xor U9768 (N_9768,N_9229,N_9461);
and U9769 (N_9769,N_9074,N_9229);
nor U9770 (N_9770,N_9465,N_9279);
nand U9771 (N_9771,N_9238,N_9197);
xnor U9772 (N_9772,N_9429,N_9066);
and U9773 (N_9773,N_9154,N_9351);
or U9774 (N_9774,N_9398,N_9347);
xnor U9775 (N_9775,N_9099,N_9254);
and U9776 (N_9776,N_9322,N_9161);
and U9777 (N_9777,N_9253,N_9468);
xor U9778 (N_9778,N_9305,N_9484);
and U9779 (N_9779,N_9193,N_9222);
and U9780 (N_9780,N_9252,N_9485);
xnor U9781 (N_9781,N_9274,N_9165);
or U9782 (N_9782,N_9049,N_9246);
and U9783 (N_9783,N_9080,N_9432);
nor U9784 (N_9784,N_9207,N_9231);
and U9785 (N_9785,N_9447,N_9057);
xor U9786 (N_9786,N_9417,N_9308);
nor U9787 (N_9787,N_9074,N_9200);
or U9788 (N_9788,N_9393,N_9020);
xor U9789 (N_9789,N_9113,N_9428);
or U9790 (N_9790,N_9153,N_9156);
or U9791 (N_9791,N_9312,N_9172);
or U9792 (N_9792,N_9153,N_9047);
or U9793 (N_9793,N_9225,N_9131);
nor U9794 (N_9794,N_9078,N_9480);
nand U9795 (N_9795,N_9406,N_9428);
nand U9796 (N_9796,N_9467,N_9012);
or U9797 (N_9797,N_9421,N_9163);
or U9798 (N_9798,N_9358,N_9139);
and U9799 (N_9799,N_9117,N_9148);
nor U9800 (N_9800,N_9453,N_9157);
nand U9801 (N_9801,N_9026,N_9048);
or U9802 (N_9802,N_9160,N_9439);
xnor U9803 (N_9803,N_9490,N_9396);
nand U9804 (N_9804,N_9144,N_9019);
nand U9805 (N_9805,N_9060,N_9384);
nand U9806 (N_9806,N_9310,N_9481);
nand U9807 (N_9807,N_9477,N_9136);
or U9808 (N_9808,N_9068,N_9123);
and U9809 (N_9809,N_9360,N_9400);
and U9810 (N_9810,N_9442,N_9457);
xnor U9811 (N_9811,N_9215,N_9157);
or U9812 (N_9812,N_9029,N_9226);
xnor U9813 (N_9813,N_9216,N_9055);
or U9814 (N_9814,N_9392,N_9226);
xor U9815 (N_9815,N_9272,N_9229);
and U9816 (N_9816,N_9385,N_9202);
nor U9817 (N_9817,N_9405,N_9413);
nand U9818 (N_9818,N_9218,N_9109);
nand U9819 (N_9819,N_9222,N_9289);
xor U9820 (N_9820,N_9107,N_9195);
or U9821 (N_9821,N_9091,N_9403);
and U9822 (N_9822,N_9381,N_9055);
xor U9823 (N_9823,N_9332,N_9172);
nor U9824 (N_9824,N_9359,N_9377);
nand U9825 (N_9825,N_9333,N_9061);
nand U9826 (N_9826,N_9123,N_9278);
or U9827 (N_9827,N_9018,N_9422);
nor U9828 (N_9828,N_9451,N_9358);
xnor U9829 (N_9829,N_9033,N_9485);
xor U9830 (N_9830,N_9094,N_9039);
nor U9831 (N_9831,N_9029,N_9260);
or U9832 (N_9832,N_9136,N_9195);
or U9833 (N_9833,N_9203,N_9214);
or U9834 (N_9834,N_9486,N_9450);
and U9835 (N_9835,N_9191,N_9218);
xor U9836 (N_9836,N_9439,N_9144);
xor U9837 (N_9837,N_9455,N_9172);
xor U9838 (N_9838,N_9288,N_9283);
and U9839 (N_9839,N_9402,N_9330);
xor U9840 (N_9840,N_9475,N_9103);
xor U9841 (N_9841,N_9255,N_9291);
and U9842 (N_9842,N_9346,N_9433);
nand U9843 (N_9843,N_9096,N_9315);
nand U9844 (N_9844,N_9160,N_9034);
or U9845 (N_9845,N_9070,N_9499);
nor U9846 (N_9846,N_9196,N_9379);
and U9847 (N_9847,N_9202,N_9463);
xor U9848 (N_9848,N_9196,N_9218);
or U9849 (N_9849,N_9103,N_9421);
nand U9850 (N_9850,N_9200,N_9376);
nand U9851 (N_9851,N_9351,N_9099);
xnor U9852 (N_9852,N_9433,N_9312);
nor U9853 (N_9853,N_9350,N_9483);
xor U9854 (N_9854,N_9106,N_9195);
nor U9855 (N_9855,N_9184,N_9071);
or U9856 (N_9856,N_9015,N_9121);
or U9857 (N_9857,N_9397,N_9460);
nand U9858 (N_9858,N_9455,N_9277);
nor U9859 (N_9859,N_9241,N_9374);
and U9860 (N_9860,N_9162,N_9493);
or U9861 (N_9861,N_9204,N_9322);
nand U9862 (N_9862,N_9418,N_9127);
nor U9863 (N_9863,N_9470,N_9424);
and U9864 (N_9864,N_9462,N_9213);
or U9865 (N_9865,N_9146,N_9189);
or U9866 (N_9866,N_9376,N_9164);
and U9867 (N_9867,N_9187,N_9114);
or U9868 (N_9868,N_9167,N_9215);
xor U9869 (N_9869,N_9280,N_9082);
nand U9870 (N_9870,N_9201,N_9069);
nor U9871 (N_9871,N_9153,N_9396);
or U9872 (N_9872,N_9192,N_9242);
nor U9873 (N_9873,N_9169,N_9399);
nor U9874 (N_9874,N_9294,N_9302);
nand U9875 (N_9875,N_9471,N_9183);
and U9876 (N_9876,N_9117,N_9400);
nand U9877 (N_9877,N_9297,N_9344);
xor U9878 (N_9878,N_9216,N_9373);
xor U9879 (N_9879,N_9076,N_9254);
or U9880 (N_9880,N_9368,N_9390);
xor U9881 (N_9881,N_9457,N_9176);
nand U9882 (N_9882,N_9420,N_9263);
nor U9883 (N_9883,N_9365,N_9229);
or U9884 (N_9884,N_9484,N_9101);
or U9885 (N_9885,N_9426,N_9015);
xor U9886 (N_9886,N_9453,N_9485);
nand U9887 (N_9887,N_9422,N_9173);
nand U9888 (N_9888,N_9317,N_9487);
nand U9889 (N_9889,N_9133,N_9149);
nand U9890 (N_9890,N_9450,N_9423);
or U9891 (N_9891,N_9122,N_9400);
nor U9892 (N_9892,N_9244,N_9187);
nand U9893 (N_9893,N_9371,N_9326);
or U9894 (N_9894,N_9399,N_9031);
nand U9895 (N_9895,N_9309,N_9307);
xnor U9896 (N_9896,N_9284,N_9372);
and U9897 (N_9897,N_9488,N_9311);
xnor U9898 (N_9898,N_9023,N_9377);
xnor U9899 (N_9899,N_9464,N_9483);
and U9900 (N_9900,N_9367,N_9306);
or U9901 (N_9901,N_9169,N_9054);
or U9902 (N_9902,N_9233,N_9306);
and U9903 (N_9903,N_9184,N_9081);
xor U9904 (N_9904,N_9386,N_9411);
xor U9905 (N_9905,N_9122,N_9331);
xor U9906 (N_9906,N_9361,N_9029);
xnor U9907 (N_9907,N_9423,N_9113);
xnor U9908 (N_9908,N_9041,N_9126);
and U9909 (N_9909,N_9070,N_9127);
xnor U9910 (N_9910,N_9132,N_9431);
nand U9911 (N_9911,N_9499,N_9465);
and U9912 (N_9912,N_9236,N_9340);
and U9913 (N_9913,N_9083,N_9198);
nor U9914 (N_9914,N_9156,N_9070);
nor U9915 (N_9915,N_9458,N_9265);
and U9916 (N_9916,N_9166,N_9069);
and U9917 (N_9917,N_9246,N_9293);
nor U9918 (N_9918,N_9230,N_9337);
and U9919 (N_9919,N_9499,N_9431);
or U9920 (N_9920,N_9223,N_9283);
or U9921 (N_9921,N_9396,N_9275);
nand U9922 (N_9922,N_9274,N_9414);
xor U9923 (N_9923,N_9306,N_9041);
xnor U9924 (N_9924,N_9321,N_9151);
nand U9925 (N_9925,N_9491,N_9103);
or U9926 (N_9926,N_9460,N_9496);
or U9927 (N_9927,N_9346,N_9466);
or U9928 (N_9928,N_9466,N_9325);
or U9929 (N_9929,N_9439,N_9068);
and U9930 (N_9930,N_9496,N_9401);
xor U9931 (N_9931,N_9154,N_9196);
nand U9932 (N_9932,N_9443,N_9017);
or U9933 (N_9933,N_9016,N_9320);
xor U9934 (N_9934,N_9140,N_9260);
and U9935 (N_9935,N_9252,N_9341);
nor U9936 (N_9936,N_9015,N_9235);
xor U9937 (N_9937,N_9438,N_9279);
nor U9938 (N_9938,N_9423,N_9044);
nand U9939 (N_9939,N_9385,N_9238);
or U9940 (N_9940,N_9027,N_9342);
xor U9941 (N_9941,N_9054,N_9057);
xnor U9942 (N_9942,N_9096,N_9306);
nor U9943 (N_9943,N_9185,N_9023);
or U9944 (N_9944,N_9447,N_9380);
nand U9945 (N_9945,N_9344,N_9109);
or U9946 (N_9946,N_9101,N_9431);
nor U9947 (N_9947,N_9085,N_9110);
nand U9948 (N_9948,N_9282,N_9256);
nand U9949 (N_9949,N_9037,N_9319);
xnor U9950 (N_9950,N_9446,N_9110);
nand U9951 (N_9951,N_9363,N_9442);
nor U9952 (N_9952,N_9231,N_9118);
nor U9953 (N_9953,N_9419,N_9011);
nor U9954 (N_9954,N_9430,N_9479);
nor U9955 (N_9955,N_9281,N_9006);
xor U9956 (N_9956,N_9312,N_9365);
nor U9957 (N_9957,N_9217,N_9005);
nand U9958 (N_9958,N_9028,N_9243);
nor U9959 (N_9959,N_9106,N_9125);
and U9960 (N_9960,N_9212,N_9145);
nor U9961 (N_9961,N_9124,N_9171);
xor U9962 (N_9962,N_9497,N_9409);
nor U9963 (N_9963,N_9387,N_9297);
or U9964 (N_9964,N_9204,N_9231);
nand U9965 (N_9965,N_9298,N_9117);
and U9966 (N_9966,N_9400,N_9080);
nor U9967 (N_9967,N_9462,N_9467);
or U9968 (N_9968,N_9370,N_9409);
or U9969 (N_9969,N_9119,N_9129);
and U9970 (N_9970,N_9256,N_9233);
xor U9971 (N_9971,N_9344,N_9336);
or U9972 (N_9972,N_9439,N_9467);
nor U9973 (N_9973,N_9184,N_9383);
xor U9974 (N_9974,N_9412,N_9264);
xor U9975 (N_9975,N_9187,N_9031);
and U9976 (N_9976,N_9406,N_9378);
nand U9977 (N_9977,N_9241,N_9455);
and U9978 (N_9978,N_9043,N_9371);
or U9979 (N_9979,N_9014,N_9404);
nor U9980 (N_9980,N_9164,N_9495);
xor U9981 (N_9981,N_9042,N_9454);
nand U9982 (N_9982,N_9368,N_9074);
nand U9983 (N_9983,N_9381,N_9435);
xor U9984 (N_9984,N_9046,N_9241);
nand U9985 (N_9985,N_9443,N_9240);
nand U9986 (N_9986,N_9166,N_9199);
or U9987 (N_9987,N_9441,N_9365);
nor U9988 (N_9988,N_9345,N_9088);
or U9989 (N_9989,N_9495,N_9016);
or U9990 (N_9990,N_9475,N_9357);
nand U9991 (N_9991,N_9121,N_9430);
and U9992 (N_9992,N_9230,N_9399);
nand U9993 (N_9993,N_9235,N_9416);
and U9994 (N_9994,N_9176,N_9189);
xnor U9995 (N_9995,N_9261,N_9336);
or U9996 (N_9996,N_9127,N_9002);
xor U9997 (N_9997,N_9198,N_9025);
xnor U9998 (N_9998,N_9297,N_9394);
and U9999 (N_9999,N_9121,N_9242);
xor UO_0 (O_0,N_9788,N_9822);
or UO_1 (O_1,N_9624,N_9856);
nor UO_2 (O_2,N_9500,N_9738);
xor UO_3 (O_3,N_9714,N_9945);
or UO_4 (O_4,N_9579,N_9506);
and UO_5 (O_5,N_9516,N_9511);
nand UO_6 (O_6,N_9768,N_9935);
nor UO_7 (O_7,N_9853,N_9510);
xnor UO_8 (O_8,N_9791,N_9849);
xnor UO_9 (O_9,N_9669,N_9797);
xor UO_10 (O_10,N_9867,N_9507);
and UO_11 (O_11,N_9586,N_9731);
nor UO_12 (O_12,N_9801,N_9934);
or UO_13 (O_13,N_9686,N_9843);
xor UO_14 (O_14,N_9895,N_9874);
nor UO_15 (O_15,N_9705,N_9562);
and UO_16 (O_16,N_9529,N_9855);
xnor UO_17 (O_17,N_9694,N_9829);
and UO_18 (O_18,N_9555,N_9543);
nor UO_19 (O_19,N_9621,N_9539);
or UO_20 (O_20,N_9972,N_9818);
nand UO_21 (O_21,N_9959,N_9885);
xor UO_22 (O_22,N_9827,N_9927);
nor UO_23 (O_23,N_9613,N_9983);
nand UO_24 (O_24,N_9701,N_9527);
nand UO_25 (O_25,N_9643,N_9965);
and UO_26 (O_26,N_9990,N_9651);
and UO_27 (O_27,N_9854,N_9661);
and UO_28 (O_28,N_9821,N_9743);
and UO_29 (O_29,N_9864,N_9870);
nand UO_30 (O_30,N_9876,N_9541);
nand UO_31 (O_31,N_9559,N_9536);
nor UO_32 (O_32,N_9671,N_9750);
nor UO_33 (O_33,N_9588,N_9781);
nand UO_34 (O_34,N_9515,N_9745);
and UO_35 (O_35,N_9626,N_9761);
and UO_36 (O_36,N_9863,N_9615);
or UO_37 (O_37,N_9834,N_9937);
or UO_38 (O_38,N_9968,N_9755);
or UO_39 (O_39,N_9703,N_9711);
and UO_40 (O_40,N_9544,N_9609);
xnor UO_41 (O_41,N_9660,N_9760);
xor UO_42 (O_42,N_9597,N_9540);
nand UO_43 (O_43,N_9950,N_9587);
nand UO_44 (O_44,N_9599,N_9675);
or UO_45 (O_45,N_9975,N_9938);
and UO_46 (O_46,N_9779,N_9986);
or UO_47 (O_47,N_9592,N_9717);
xor UO_48 (O_48,N_9948,N_9535);
xor UO_49 (O_49,N_9908,N_9673);
nand UO_50 (O_50,N_9891,N_9851);
or UO_51 (O_51,N_9570,N_9632);
and UO_52 (O_52,N_9958,N_9780);
and UO_53 (O_53,N_9978,N_9769);
nand UO_54 (O_54,N_9848,N_9756);
or UO_55 (O_55,N_9922,N_9709);
nor UO_56 (O_56,N_9973,N_9608);
nand UO_57 (O_57,N_9702,N_9551);
and UO_58 (O_58,N_9641,N_9678);
and UO_59 (O_59,N_9954,N_9682);
nor UO_60 (O_60,N_9502,N_9590);
and UO_61 (O_61,N_9635,N_9850);
nor UO_62 (O_62,N_9857,N_9905);
xnor UO_63 (O_63,N_9815,N_9886);
or UO_64 (O_64,N_9787,N_9839);
xnor UO_65 (O_65,N_9554,N_9795);
nand UO_66 (O_66,N_9931,N_9556);
or UO_67 (O_67,N_9698,N_9774);
or UO_68 (O_68,N_9837,N_9676);
nand UO_69 (O_69,N_9976,N_9593);
nand UO_70 (O_70,N_9674,N_9580);
or UO_71 (O_71,N_9881,N_9812);
and UO_72 (O_72,N_9523,N_9913);
xnor UO_73 (O_73,N_9636,N_9748);
and UO_74 (O_74,N_9899,N_9569);
or UO_75 (O_75,N_9557,N_9566);
xor UO_76 (O_76,N_9670,N_9893);
and UO_77 (O_77,N_9681,N_9877);
nor UO_78 (O_78,N_9658,N_9627);
or UO_79 (O_79,N_9879,N_9806);
or UO_80 (O_80,N_9503,N_9604);
xnor UO_81 (O_81,N_9776,N_9645);
or UO_82 (O_82,N_9939,N_9524);
nand UO_83 (O_83,N_9929,N_9716);
or UO_84 (O_84,N_9966,N_9949);
or UO_85 (O_85,N_9573,N_9517);
or UO_86 (O_86,N_9718,N_9900);
or UO_87 (O_87,N_9648,N_9552);
nor UO_88 (O_88,N_9647,N_9871);
and UO_89 (O_89,N_9794,N_9969);
nor UO_90 (O_90,N_9538,N_9697);
and UO_91 (O_91,N_9724,N_9928);
xor UO_92 (O_92,N_9962,N_9987);
and UO_93 (O_93,N_9630,N_9649);
nor UO_94 (O_94,N_9810,N_9764);
nor UO_95 (O_95,N_9833,N_9578);
and UO_96 (O_96,N_9904,N_9875);
and UO_97 (O_97,N_9943,N_9998);
nand UO_98 (O_98,N_9662,N_9903);
nor UO_99 (O_99,N_9751,N_9816);
and UO_100 (O_100,N_9501,N_9991);
and UO_101 (O_101,N_9811,N_9634);
and UO_102 (O_102,N_9898,N_9677);
nand UO_103 (O_103,N_9633,N_9988);
or UO_104 (O_104,N_9808,N_9901);
nand UO_105 (O_105,N_9719,N_9666);
xor UO_106 (O_106,N_9690,N_9866);
nand UO_107 (O_107,N_9800,N_9721);
and UO_108 (O_108,N_9894,N_9663);
or UO_109 (O_109,N_9548,N_9957);
nor UO_110 (O_110,N_9777,N_9610);
xnor UO_111 (O_111,N_9942,N_9672);
xnor UO_112 (O_112,N_9622,N_9880);
and UO_113 (O_113,N_9730,N_9519);
nor UO_114 (O_114,N_9915,N_9656);
xnor UO_115 (O_115,N_9897,N_9955);
and UO_116 (O_116,N_9842,N_9838);
or UO_117 (O_117,N_9923,N_9553);
or UO_118 (O_118,N_9979,N_9531);
and UO_119 (O_119,N_9728,N_9653);
and UO_120 (O_120,N_9936,N_9512);
or UO_121 (O_121,N_9947,N_9888);
nor UO_122 (O_122,N_9932,N_9530);
nor UO_123 (O_123,N_9605,N_9504);
and UO_124 (O_124,N_9558,N_9873);
or UO_125 (O_125,N_9642,N_9933);
nand UO_126 (O_126,N_9679,N_9723);
nor UO_127 (O_127,N_9970,N_9542);
and UO_128 (O_128,N_9712,N_9537);
or UO_129 (O_129,N_9865,N_9757);
nor UO_130 (O_130,N_9737,N_9759);
nand UO_131 (O_131,N_9884,N_9992);
nand UO_132 (O_132,N_9889,N_9509);
nand UO_133 (O_133,N_9665,N_9868);
nand UO_134 (O_134,N_9963,N_9692);
xnor UO_135 (O_135,N_9583,N_9550);
nand UO_136 (O_136,N_9980,N_9704);
and UO_137 (O_137,N_9646,N_9726);
xnor UO_138 (O_138,N_9786,N_9734);
xnor UO_139 (O_139,N_9652,N_9591);
nand UO_140 (O_140,N_9926,N_9564);
nor UO_141 (O_141,N_9775,N_9532);
and UO_142 (O_142,N_9982,N_9999);
xor UO_143 (O_143,N_9577,N_9766);
nor UO_144 (O_144,N_9773,N_9740);
or UO_145 (O_145,N_9802,N_9925);
or UO_146 (O_146,N_9930,N_9872);
nor UO_147 (O_147,N_9572,N_9568);
and UO_148 (O_148,N_9585,N_9984);
or UO_149 (O_149,N_9520,N_9807);
or UO_150 (O_150,N_9598,N_9616);
or UO_151 (O_151,N_9817,N_9911);
and UO_152 (O_152,N_9747,N_9637);
nor UO_153 (O_153,N_9944,N_9770);
or UO_154 (O_154,N_9765,N_9639);
nor UO_155 (O_155,N_9561,N_9789);
and UO_156 (O_156,N_9892,N_9575);
and UO_157 (O_157,N_9623,N_9790);
nor UO_158 (O_158,N_9887,N_9890);
and UO_159 (O_159,N_9582,N_9846);
or UO_160 (O_160,N_9912,N_9819);
nand UO_161 (O_161,N_9852,N_9534);
or UO_162 (O_162,N_9741,N_9700);
xor UO_163 (O_163,N_9798,N_9725);
and UO_164 (O_164,N_9640,N_9657);
nand UO_165 (O_165,N_9840,N_9828);
or UO_166 (O_166,N_9859,N_9513);
xnor UO_167 (O_167,N_9971,N_9735);
or UO_168 (O_168,N_9707,N_9563);
nor UO_169 (O_169,N_9514,N_9906);
or UO_170 (O_170,N_9878,N_9584);
nand UO_171 (O_171,N_9691,N_9917);
and UO_172 (O_172,N_9739,N_9771);
nor UO_173 (O_173,N_9589,N_9919);
or UO_174 (O_174,N_9618,N_9758);
xor UO_175 (O_175,N_9985,N_9754);
or UO_176 (O_176,N_9744,N_9638);
xnor UO_177 (O_177,N_9547,N_9767);
nand UO_178 (O_178,N_9628,N_9956);
nand UO_179 (O_179,N_9614,N_9727);
nand UO_180 (O_180,N_9625,N_9720);
nand UO_181 (O_181,N_9823,N_9820);
nand UO_182 (O_182,N_9782,N_9909);
nor UO_183 (O_183,N_9752,N_9805);
xor UO_184 (O_184,N_9668,N_9687);
xor UO_185 (O_185,N_9841,N_9545);
xor UO_186 (O_186,N_9736,N_9994);
xnor UO_187 (O_187,N_9862,N_9804);
or UO_188 (O_188,N_9964,N_9960);
or UO_189 (O_189,N_9629,N_9785);
and UO_190 (O_190,N_9961,N_9784);
and UO_191 (O_191,N_9710,N_9600);
nand UO_192 (O_192,N_9549,N_9611);
nand UO_193 (O_193,N_9977,N_9920);
and UO_194 (O_194,N_9596,N_9924);
nor UO_195 (O_195,N_9921,N_9683);
nor UO_196 (O_196,N_9619,N_9722);
nand UO_197 (O_197,N_9941,N_9825);
xnor UO_198 (O_198,N_9940,N_9799);
or UO_199 (O_199,N_9729,N_9644);
nand UO_200 (O_200,N_9595,N_9996);
nand UO_201 (O_201,N_9581,N_9847);
xor UO_202 (O_202,N_9508,N_9831);
xor UO_203 (O_203,N_9792,N_9505);
nor UO_204 (O_204,N_9688,N_9796);
nand UO_205 (O_205,N_9574,N_9813);
and UO_206 (O_206,N_9860,N_9601);
nand UO_207 (O_207,N_9902,N_9606);
and UO_208 (O_208,N_9525,N_9607);
nor UO_209 (O_209,N_9809,N_9650);
and UO_210 (O_210,N_9953,N_9708);
nand UO_211 (O_211,N_9617,N_9783);
nor UO_212 (O_212,N_9685,N_9762);
and UO_213 (O_213,N_9946,N_9793);
xor UO_214 (O_214,N_9689,N_9655);
nor UO_215 (O_215,N_9715,N_9612);
and UO_216 (O_216,N_9733,N_9989);
xor UO_217 (O_217,N_9995,N_9916);
nor UO_218 (O_218,N_9526,N_9654);
nand UO_219 (O_219,N_9993,N_9835);
xnor UO_220 (O_220,N_9845,N_9603);
xor UO_221 (O_221,N_9861,N_9753);
xor UO_222 (O_222,N_9858,N_9997);
nand UO_223 (O_223,N_9824,N_9567);
xnor UO_224 (O_224,N_9882,N_9560);
nor UO_225 (O_225,N_9533,N_9620);
nor UO_226 (O_226,N_9844,N_9830);
nor UO_227 (O_227,N_9576,N_9742);
nand UO_228 (O_228,N_9695,N_9680);
or UO_229 (O_229,N_9565,N_9706);
nor UO_230 (O_230,N_9518,N_9746);
and UO_231 (O_231,N_9952,N_9664);
xor UO_232 (O_232,N_9749,N_9910);
nand UO_233 (O_233,N_9699,N_9522);
or UO_234 (O_234,N_9732,N_9826);
xnor UO_235 (O_235,N_9814,N_9832);
xor UO_236 (O_236,N_9907,N_9974);
and UO_237 (O_237,N_9981,N_9836);
nor UO_238 (O_238,N_9896,N_9763);
xor UO_239 (O_239,N_9528,N_9667);
xnor UO_240 (O_240,N_9693,N_9869);
xnor UO_241 (O_241,N_9772,N_9696);
and UO_242 (O_242,N_9951,N_9778);
xnor UO_243 (O_243,N_9684,N_9631);
xnor UO_244 (O_244,N_9883,N_9803);
xor UO_245 (O_245,N_9713,N_9521);
nand UO_246 (O_246,N_9594,N_9602);
or UO_247 (O_247,N_9918,N_9571);
nand UO_248 (O_248,N_9659,N_9546);
nor UO_249 (O_249,N_9914,N_9967);
xnor UO_250 (O_250,N_9639,N_9881);
nand UO_251 (O_251,N_9990,N_9995);
nor UO_252 (O_252,N_9701,N_9925);
or UO_253 (O_253,N_9860,N_9576);
and UO_254 (O_254,N_9849,N_9989);
nand UO_255 (O_255,N_9626,N_9979);
or UO_256 (O_256,N_9556,N_9640);
xnor UO_257 (O_257,N_9921,N_9729);
or UO_258 (O_258,N_9888,N_9670);
or UO_259 (O_259,N_9664,N_9614);
and UO_260 (O_260,N_9862,N_9731);
and UO_261 (O_261,N_9647,N_9600);
nor UO_262 (O_262,N_9903,N_9842);
nand UO_263 (O_263,N_9657,N_9617);
xnor UO_264 (O_264,N_9920,N_9536);
or UO_265 (O_265,N_9958,N_9762);
nor UO_266 (O_266,N_9507,N_9569);
nand UO_267 (O_267,N_9890,N_9737);
nand UO_268 (O_268,N_9873,N_9767);
and UO_269 (O_269,N_9747,N_9804);
xor UO_270 (O_270,N_9527,N_9671);
nand UO_271 (O_271,N_9659,N_9592);
or UO_272 (O_272,N_9958,N_9550);
nand UO_273 (O_273,N_9867,N_9727);
xor UO_274 (O_274,N_9988,N_9615);
or UO_275 (O_275,N_9571,N_9816);
and UO_276 (O_276,N_9626,N_9709);
xor UO_277 (O_277,N_9905,N_9968);
and UO_278 (O_278,N_9575,N_9986);
and UO_279 (O_279,N_9957,N_9507);
nand UO_280 (O_280,N_9747,N_9534);
nor UO_281 (O_281,N_9855,N_9956);
nor UO_282 (O_282,N_9936,N_9978);
nor UO_283 (O_283,N_9704,N_9720);
and UO_284 (O_284,N_9973,N_9686);
xor UO_285 (O_285,N_9632,N_9989);
nor UO_286 (O_286,N_9706,N_9666);
or UO_287 (O_287,N_9838,N_9971);
nor UO_288 (O_288,N_9778,N_9687);
and UO_289 (O_289,N_9557,N_9976);
nor UO_290 (O_290,N_9954,N_9880);
nand UO_291 (O_291,N_9500,N_9769);
and UO_292 (O_292,N_9551,N_9989);
nor UO_293 (O_293,N_9844,N_9877);
xnor UO_294 (O_294,N_9986,N_9946);
xnor UO_295 (O_295,N_9929,N_9676);
or UO_296 (O_296,N_9710,N_9828);
xor UO_297 (O_297,N_9871,N_9614);
nand UO_298 (O_298,N_9569,N_9908);
xnor UO_299 (O_299,N_9898,N_9700);
xnor UO_300 (O_300,N_9570,N_9608);
or UO_301 (O_301,N_9741,N_9703);
and UO_302 (O_302,N_9517,N_9825);
or UO_303 (O_303,N_9917,N_9880);
xnor UO_304 (O_304,N_9720,N_9933);
xor UO_305 (O_305,N_9586,N_9988);
and UO_306 (O_306,N_9526,N_9821);
and UO_307 (O_307,N_9587,N_9934);
nand UO_308 (O_308,N_9539,N_9533);
xnor UO_309 (O_309,N_9612,N_9889);
nor UO_310 (O_310,N_9726,N_9705);
nor UO_311 (O_311,N_9777,N_9825);
or UO_312 (O_312,N_9914,N_9506);
nor UO_313 (O_313,N_9761,N_9983);
and UO_314 (O_314,N_9685,N_9898);
nor UO_315 (O_315,N_9963,N_9956);
xor UO_316 (O_316,N_9779,N_9953);
nand UO_317 (O_317,N_9522,N_9614);
nor UO_318 (O_318,N_9575,N_9599);
xnor UO_319 (O_319,N_9764,N_9903);
and UO_320 (O_320,N_9984,N_9724);
nand UO_321 (O_321,N_9671,N_9634);
nand UO_322 (O_322,N_9516,N_9847);
and UO_323 (O_323,N_9868,N_9644);
and UO_324 (O_324,N_9646,N_9711);
xnor UO_325 (O_325,N_9892,N_9577);
nor UO_326 (O_326,N_9541,N_9865);
nand UO_327 (O_327,N_9753,N_9549);
nor UO_328 (O_328,N_9962,N_9509);
or UO_329 (O_329,N_9938,N_9533);
nor UO_330 (O_330,N_9658,N_9851);
or UO_331 (O_331,N_9678,N_9662);
nor UO_332 (O_332,N_9924,N_9631);
xor UO_333 (O_333,N_9723,N_9749);
nor UO_334 (O_334,N_9685,N_9967);
or UO_335 (O_335,N_9696,N_9537);
nor UO_336 (O_336,N_9624,N_9601);
nand UO_337 (O_337,N_9772,N_9940);
nand UO_338 (O_338,N_9633,N_9667);
nor UO_339 (O_339,N_9673,N_9644);
nor UO_340 (O_340,N_9718,N_9996);
nor UO_341 (O_341,N_9664,N_9773);
or UO_342 (O_342,N_9608,N_9631);
nor UO_343 (O_343,N_9952,N_9832);
nand UO_344 (O_344,N_9814,N_9753);
nor UO_345 (O_345,N_9909,N_9613);
nand UO_346 (O_346,N_9842,N_9607);
nand UO_347 (O_347,N_9995,N_9948);
or UO_348 (O_348,N_9856,N_9977);
nand UO_349 (O_349,N_9796,N_9542);
and UO_350 (O_350,N_9578,N_9519);
or UO_351 (O_351,N_9877,N_9946);
xor UO_352 (O_352,N_9742,N_9838);
or UO_353 (O_353,N_9761,N_9876);
nor UO_354 (O_354,N_9561,N_9606);
or UO_355 (O_355,N_9764,N_9908);
and UO_356 (O_356,N_9613,N_9670);
and UO_357 (O_357,N_9852,N_9975);
and UO_358 (O_358,N_9773,N_9548);
nor UO_359 (O_359,N_9586,N_9625);
nand UO_360 (O_360,N_9838,N_9586);
xnor UO_361 (O_361,N_9574,N_9723);
and UO_362 (O_362,N_9694,N_9628);
xor UO_363 (O_363,N_9653,N_9950);
or UO_364 (O_364,N_9833,N_9503);
nor UO_365 (O_365,N_9757,N_9898);
nor UO_366 (O_366,N_9836,N_9681);
nor UO_367 (O_367,N_9679,N_9500);
xor UO_368 (O_368,N_9526,N_9912);
nor UO_369 (O_369,N_9797,N_9707);
nand UO_370 (O_370,N_9868,N_9825);
and UO_371 (O_371,N_9557,N_9834);
nor UO_372 (O_372,N_9901,N_9512);
nand UO_373 (O_373,N_9625,N_9615);
nand UO_374 (O_374,N_9905,N_9524);
and UO_375 (O_375,N_9835,N_9916);
and UO_376 (O_376,N_9588,N_9969);
nand UO_377 (O_377,N_9843,N_9571);
nor UO_378 (O_378,N_9764,N_9841);
xor UO_379 (O_379,N_9589,N_9876);
nor UO_380 (O_380,N_9512,N_9865);
nor UO_381 (O_381,N_9651,N_9548);
nor UO_382 (O_382,N_9768,N_9547);
nor UO_383 (O_383,N_9576,N_9962);
xnor UO_384 (O_384,N_9878,N_9856);
nor UO_385 (O_385,N_9879,N_9673);
nand UO_386 (O_386,N_9556,N_9665);
nand UO_387 (O_387,N_9669,N_9788);
nor UO_388 (O_388,N_9865,N_9597);
xor UO_389 (O_389,N_9965,N_9552);
nand UO_390 (O_390,N_9736,N_9505);
nor UO_391 (O_391,N_9611,N_9507);
nand UO_392 (O_392,N_9540,N_9927);
nor UO_393 (O_393,N_9942,N_9822);
and UO_394 (O_394,N_9513,N_9922);
nor UO_395 (O_395,N_9621,N_9685);
xnor UO_396 (O_396,N_9552,N_9949);
xor UO_397 (O_397,N_9599,N_9688);
nand UO_398 (O_398,N_9753,N_9658);
or UO_399 (O_399,N_9552,N_9508);
nand UO_400 (O_400,N_9771,N_9629);
and UO_401 (O_401,N_9525,N_9813);
nand UO_402 (O_402,N_9784,N_9986);
and UO_403 (O_403,N_9932,N_9858);
and UO_404 (O_404,N_9943,N_9871);
or UO_405 (O_405,N_9902,N_9723);
xnor UO_406 (O_406,N_9876,N_9894);
nand UO_407 (O_407,N_9842,N_9869);
xor UO_408 (O_408,N_9965,N_9765);
and UO_409 (O_409,N_9857,N_9686);
nand UO_410 (O_410,N_9963,N_9839);
and UO_411 (O_411,N_9541,N_9966);
xor UO_412 (O_412,N_9529,N_9839);
or UO_413 (O_413,N_9655,N_9853);
xor UO_414 (O_414,N_9917,N_9764);
nor UO_415 (O_415,N_9615,N_9633);
xor UO_416 (O_416,N_9881,N_9979);
and UO_417 (O_417,N_9569,N_9939);
nor UO_418 (O_418,N_9864,N_9933);
and UO_419 (O_419,N_9500,N_9602);
and UO_420 (O_420,N_9886,N_9586);
nand UO_421 (O_421,N_9754,N_9724);
and UO_422 (O_422,N_9794,N_9876);
nand UO_423 (O_423,N_9594,N_9593);
xnor UO_424 (O_424,N_9713,N_9958);
or UO_425 (O_425,N_9579,N_9655);
xor UO_426 (O_426,N_9786,N_9961);
xnor UO_427 (O_427,N_9825,N_9758);
xnor UO_428 (O_428,N_9902,N_9957);
nor UO_429 (O_429,N_9680,N_9538);
xnor UO_430 (O_430,N_9964,N_9755);
and UO_431 (O_431,N_9591,N_9668);
or UO_432 (O_432,N_9535,N_9516);
and UO_433 (O_433,N_9527,N_9669);
and UO_434 (O_434,N_9709,N_9577);
xnor UO_435 (O_435,N_9591,N_9831);
or UO_436 (O_436,N_9612,N_9734);
and UO_437 (O_437,N_9525,N_9928);
or UO_438 (O_438,N_9779,N_9512);
xor UO_439 (O_439,N_9912,N_9913);
nand UO_440 (O_440,N_9973,N_9674);
and UO_441 (O_441,N_9772,N_9503);
nand UO_442 (O_442,N_9999,N_9882);
or UO_443 (O_443,N_9726,N_9676);
or UO_444 (O_444,N_9598,N_9857);
and UO_445 (O_445,N_9751,N_9797);
nor UO_446 (O_446,N_9776,N_9921);
nand UO_447 (O_447,N_9951,N_9589);
nand UO_448 (O_448,N_9932,N_9787);
xnor UO_449 (O_449,N_9787,N_9766);
and UO_450 (O_450,N_9849,N_9619);
or UO_451 (O_451,N_9707,N_9679);
or UO_452 (O_452,N_9591,N_9709);
nor UO_453 (O_453,N_9592,N_9732);
xnor UO_454 (O_454,N_9738,N_9992);
nand UO_455 (O_455,N_9634,N_9704);
xnor UO_456 (O_456,N_9968,N_9892);
nand UO_457 (O_457,N_9892,N_9570);
and UO_458 (O_458,N_9812,N_9525);
or UO_459 (O_459,N_9567,N_9825);
and UO_460 (O_460,N_9770,N_9943);
xor UO_461 (O_461,N_9680,N_9602);
xor UO_462 (O_462,N_9869,N_9748);
nor UO_463 (O_463,N_9816,N_9696);
and UO_464 (O_464,N_9725,N_9940);
xor UO_465 (O_465,N_9982,N_9996);
nand UO_466 (O_466,N_9609,N_9590);
and UO_467 (O_467,N_9640,N_9630);
xnor UO_468 (O_468,N_9866,N_9522);
nand UO_469 (O_469,N_9795,N_9544);
and UO_470 (O_470,N_9880,N_9712);
and UO_471 (O_471,N_9739,N_9902);
nand UO_472 (O_472,N_9936,N_9805);
nor UO_473 (O_473,N_9992,N_9608);
xor UO_474 (O_474,N_9637,N_9740);
xnor UO_475 (O_475,N_9725,N_9996);
or UO_476 (O_476,N_9795,N_9986);
xor UO_477 (O_477,N_9531,N_9923);
xor UO_478 (O_478,N_9841,N_9713);
xnor UO_479 (O_479,N_9978,N_9717);
nor UO_480 (O_480,N_9732,N_9903);
and UO_481 (O_481,N_9827,N_9600);
xor UO_482 (O_482,N_9670,N_9976);
nor UO_483 (O_483,N_9868,N_9582);
or UO_484 (O_484,N_9783,N_9847);
and UO_485 (O_485,N_9834,N_9859);
nand UO_486 (O_486,N_9725,N_9571);
xnor UO_487 (O_487,N_9904,N_9522);
or UO_488 (O_488,N_9578,N_9778);
nand UO_489 (O_489,N_9949,N_9718);
xor UO_490 (O_490,N_9882,N_9626);
and UO_491 (O_491,N_9608,N_9683);
nand UO_492 (O_492,N_9832,N_9818);
nand UO_493 (O_493,N_9885,N_9824);
and UO_494 (O_494,N_9847,N_9757);
nand UO_495 (O_495,N_9980,N_9629);
and UO_496 (O_496,N_9809,N_9589);
nand UO_497 (O_497,N_9769,N_9667);
nand UO_498 (O_498,N_9579,N_9685);
xor UO_499 (O_499,N_9740,N_9512);
nand UO_500 (O_500,N_9878,N_9907);
nor UO_501 (O_501,N_9844,N_9620);
xnor UO_502 (O_502,N_9779,N_9526);
nor UO_503 (O_503,N_9997,N_9947);
nor UO_504 (O_504,N_9513,N_9589);
or UO_505 (O_505,N_9512,N_9868);
and UO_506 (O_506,N_9785,N_9536);
or UO_507 (O_507,N_9638,N_9862);
nor UO_508 (O_508,N_9690,N_9942);
nor UO_509 (O_509,N_9643,N_9765);
and UO_510 (O_510,N_9869,N_9611);
xor UO_511 (O_511,N_9997,N_9853);
and UO_512 (O_512,N_9657,N_9660);
nand UO_513 (O_513,N_9990,N_9818);
and UO_514 (O_514,N_9740,N_9619);
or UO_515 (O_515,N_9681,N_9872);
and UO_516 (O_516,N_9711,N_9595);
or UO_517 (O_517,N_9733,N_9808);
nand UO_518 (O_518,N_9559,N_9856);
nand UO_519 (O_519,N_9579,N_9661);
and UO_520 (O_520,N_9971,N_9562);
nor UO_521 (O_521,N_9988,N_9845);
nor UO_522 (O_522,N_9611,N_9932);
or UO_523 (O_523,N_9554,N_9870);
nand UO_524 (O_524,N_9819,N_9539);
nor UO_525 (O_525,N_9613,N_9505);
nor UO_526 (O_526,N_9969,N_9852);
nand UO_527 (O_527,N_9821,N_9610);
and UO_528 (O_528,N_9527,N_9649);
nand UO_529 (O_529,N_9667,N_9705);
xnor UO_530 (O_530,N_9524,N_9549);
xnor UO_531 (O_531,N_9985,N_9505);
xor UO_532 (O_532,N_9682,N_9508);
and UO_533 (O_533,N_9669,N_9991);
or UO_534 (O_534,N_9675,N_9820);
nand UO_535 (O_535,N_9868,N_9782);
or UO_536 (O_536,N_9910,N_9616);
or UO_537 (O_537,N_9602,N_9566);
and UO_538 (O_538,N_9935,N_9763);
or UO_539 (O_539,N_9595,N_9789);
and UO_540 (O_540,N_9736,N_9923);
nand UO_541 (O_541,N_9825,N_9830);
xor UO_542 (O_542,N_9751,N_9719);
xor UO_543 (O_543,N_9991,N_9516);
nor UO_544 (O_544,N_9849,N_9905);
nor UO_545 (O_545,N_9538,N_9565);
and UO_546 (O_546,N_9697,N_9592);
xor UO_547 (O_547,N_9556,N_9534);
or UO_548 (O_548,N_9561,N_9757);
nand UO_549 (O_549,N_9803,N_9794);
or UO_550 (O_550,N_9906,N_9535);
nor UO_551 (O_551,N_9739,N_9664);
and UO_552 (O_552,N_9530,N_9905);
nor UO_553 (O_553,N_9788,N_9514);
or UO_554 (O_554,N_9603,N_9831);
or UO_555 (O_555,N_9547,N_9927);
nor UO_556 (O_556,N_9755,N_9732);
xor UO_557 (O_557,N_9573,N_9508);
nor UO_558 (O_558,N_9640,N_9699);
xor UO_559 (O_559,N_9988,N_9732);
nor UO_560 (O_560,N_9625,N_9767);
and UO_561 (O_561,N_9779,N_9566);
xor UO_562 (O_562,N_9558,N_9638);
and UO_563 (O_563,N_9814,N_9732);
nor UO_564 (O_564,N_9759,N_9613);
xor UO_565 (O_565,N_9757,N_9746);
or UO_566 (O_566,N_9794,N_9920);
nand UO_567 (O_567,N_9831,N_9947);
nand UO_568 (O_568,N_9636,N_9912);
or UO_569 (O_569,N_9848,N_9944);
and UO_570 (O_570,N_9776,N_9946);
or UO_571 (O_571,N_9629,N_9669);
nand UO_572 (O_572,N_9896,N_9550);
nor UO_573 (O_573,N_9979,N_9627);
nor UO_574 (O_574,N_9918,N_9537);
nand UO_575 (O_575,N_9876,N_9679);
and UO_576 (O_576,N_9885,N_9802);
nor UO_577 (O_577,N_9861,N_9990);
xor UO_578 (O_578,N_9631,N_9612);
nor UO_579 (O_579,N_9587,N_9993);
xor UO_580 (O_580,N_9784,N_9555);
and UO_581 (O_581,N_9962,N_9526);
and UO_582 (O_582,N_9891,N_9669);
xnor UO_583 (O_583,N_9772,N_9677);
nor UO_584 (O_584,N_9624,N_9807);
xnor UO_585 (O_585,N_9568,N_9862);
or UO_586 (O_586,N_9540,N_9890);
and UO_587 (O_587,N_9953,N_9601);
and UO_588 (O_588,N_9953,N_9618);
or UO_589 (O_589,N_9794,N_9641);
xor UO_590 (O_590,N_9576,N_9562);
nor UO_591 (O_591,N_9668,N_9872);
or UO_592 (O_592,N_9978,N_9602);
nand UO_593 (O_593,N_9955,N_9566);
xnor UO_594 (O_594,N_9626,N_9694);
xor UO_595 (O_595,N_9804,N_9600);
and UO_596 (O_596,N_9595,N_9719);
nand UO_597 (O_597,N_9609,N_9555);
nor UO_598 (O_598,N_9655,N_9696);
or UO_599 (O_599,N_9923,N_9850);
or UO_600 (O_600,N_9664,N_9799);
nand UO_601 (O_601,N_9581,N_9981);
nand UO_602 (O_602,N_9979,N_9997);
or UO_603 (O_603,N_9690,N_9773);
and UO_604 (O_604,N_9840,N_9505);
nand UO_605 (O_605,N_9543,N_9623);
nand UO_606 (O_606,N_9770,N_9849);
xor UO_607 (O_607,N_9953,N_9530);
xor UO_608 (O_608,N_9730,N_9952);
and UO_609 (O_609,N_9922,N_9618);
or UO_610 (O_610,N_9820,N_9836);
nand UO_611 (O_611,N_9835,N_9990);
xor UO_612 (O_612,N_9591,N_9716);
xor UO_613 (O_613,N_9955,N_9764);
and UO_614 (O_614,N_9933,N_9836);
nand UO_615 (O_615,N_9667,N_9548);
or UO_616 (O_616,N_9548,N_9879);
nor UO_617 (O_617,N_9843,N_9624);
xor UO_618 (O_618,N_9951,N_9806);
nor UO_619 (O_619,N_9587,N_9779);
xor UO_620 (O_620,N_9875,N_9922);
nor UO_621 (O_621,N_9572,N_9649);
nor UO_622 (O_622,N_9628,N_9861);
or UO_623 (O_623,N_9830,N_9718);
xnor UO_624 (O_624,N_9714,N_9677);
nand UO_625 (O_625,N_9960,N_9759);
nor UO_626 (O_626,N_9619,N_9538);
and UO_627 (O_627,N_9610,N_9802);
xnor UO_628 (O_628,N_9712,N_9860);
and UO_629 (O_629,N_9712,N_9600);
or UO_630 (O_630,N_9522,N_9902);
nor UO_631 (O_631,N_9537,N_9870);
or UO_632 (O_632,N_9928,N_9504);
nand UO_633 (O_633,N_9640,N_9781);
nor UO_634 (O_634,N_9627,N_9686);
nor UO_635 (O_635,N_9933,N_9983);
nand UO_636 (O_636,N_9713,N_9949);
or UO_637 (O_637,N_9818,N_9902);
and UO_638 (O_638,N_9600,N_9791);
xnor UO_639 (O_639,N_9638,N_9612);
nor UO_640 (O_640,N_9838,N_9849);
or UO_641 (O_641,N_9647,N_9635);
xor UO_642 (O_642,N_9983,N_9779);
and UO_643 (O_643,N_9983,N_9957);
nand UO_644 (O_644,N_9994,N_9556);
or UO_645 (O_645,N_9559,N_9916);
or UO_646 (O_646,N_9979,N_9684);
or UO_647 (O_647,N_9921,N_9568);
or UO_648 (O_648,N_9848,N_9502);
nor UO_649 (O_649,N_9586,N_9851);
nor UO_650 (O_650,N_9873,N_9579);
xor UO_651 (O_651,N_9903,N_9793);
nor UO_652 (O_652,N_9641,N_9851);
nor UO_653 (O_653,N_9626,N_9544);
or UO_654 (O_654,N_9581,N_9811);
or UO_655 (O_655,N_9779,N_9699);
xor UO_656 (O_656,N_9645,N_9563);
or UO_657 (O_657,N_9803,N_9762);
nor UO_658 (O_658,N_9549,N_9764);
nand UO_659 (O_659,N_9731,N_9529);
nor UO_660 (O_660,N_9940,N_9956);
xnor UO_661 (O_661,N_9581,N_9534);
or UO_662 (O_662,N_9741,N_9607);
and UO_663 (O_663,N_9754,N_9877);
and UO_664 (O_664,N_9992,N_9928);
nor UO_665 (O_665,N_9944,N_9958);
and UO_666 (O_666,N_9574,N_9556);
xor UO_667 (O_667,N_9778,N_9777);
nand UO_668 (O_668,N_9946,N_9545);
nand UO_669 (O_669,N_9708,N_9750);
nor UO_670 (O_670,N_9645,N_9961);
nor UO_671 (O_671,N_9696,N_9822);
or UO_672 (O_672,N_9570,N_9784);
xor UO_673 (O_673,N_9872,N_9914);
xnor UO_674 (O_674,N_9754,N_9750);
and UO_675 (O_675,N_9574,N_9687);
nand UO_676 (O_676,N_9830,N_9779);
xnor UO_677 (O_677,N_9551,N_9765);
and UO_678 (O_678,N_9959,N_9549);
nand UO_679 (O_679,N_9922,N_9531);
nand UO_680 (O_680,N_9784,N_9669);
nor UO_681 (O_681,N_9664,N_9561);
xnor UO_682 (O_682,N_9885,N_9676);
nor UO_683 (O_683,N_9558,N_9799);
and UO_684 (O_684,N_9964,N_9931);
xor UO_685 (O_685,N_9818,N_9982);
xor UO_686 (O_686,N_9753,N_9567);
nand UO_687 (O_687,N_9656,N_9899);
nor UO_688 (O_688,N_9558,N_9877);
or UO_689 (O_689,N_9636,N_9930);
and UO_690 (O_690,N_9851,N_9994);
or UO_691 (O_691,N_9902,N_9969);
xnor UO_692 (O_692,N_9656,N_9582);
or UO_693 (O_693,N_9874,N_9561);
and UO_694 (O_694,N_9852,N_9811);
nand UO_695 (O_695,N_9957,N_9569);
and UO_696 (O_696,N_9860,N_9657);
nand UO_697 (O_697,N_9861,N_9958);
or UO_698 (O_698,N_9865,N_9912);
and UO_699 (O_699,N_9833,N_9968);
or UO_700 (O_700,N_9538,N_9862);
nand UO_701 (O_701,N_9979,N_9864);
or UO_702 (O_702,N_9771,N_9878);
nor UO_703 (O_703,N_9803,N_9959);
nand UO_704 (O_704,N_9951,N_9874);
nor UO_705 (O_705,N_9750,N_9904);
xor UO_706 (O_706,N_9713,N_9672);
or UO_707 (O_707,N_9711,N_9577);
or UO_708 (O_708,N_9606,N_9978);
or UO_709 (O_709,N_9879,N_9788);
nor UO_710 (O_710,N_9943,N_9819);
nand UO_711 (O_711,N_9651,N_9589);
xnor UO_712 (O_712,N_9782,N_9815);
xnor UO_713 (O_713,N_9817,N_9976);
nand UO_714 (O_714,N_9943,N_9799);
nor UO_715 (O_715,N_9502,N_9918);
nand UO_716 (O_716,N_9601,N_9535);
xor UO_717 (O_717,N_9735,N_9853);
xnor UO_718 (O_718,N_9606,N_9549);
or UO_719 (O_719,N_9969,N_9505);
nor UO_720 (O_720,N_9880,N_9719);
xor UO_721 (O_721,N_9630,N_9587);
xnor UO_722 (O_722,N_9532,N_9721);
nor UO_723 (O_723,N_9522,N_9591);
and UO_724 (O_724,N_9824,N_9798);
or UO_725 (O_725,N_9691,N_9883);
nand UO_726 (O_726,N_9661,N_9796);
xnor UO_727 (O_727,N_9768,N_9650);
and UO_728 (O_728,N_9794,N_9629);
xnor UO_729 (O_729,N_9709,N_9589);
nor UO_730 (O_730,N_9998,N_9530);
xnor UO_731 (O_731,N_9690,N_9889);
or UO_732 (O_732,N_9780,N_9715);
nand UO_733 (O_733,N_9850,N_9959);
and UO_734 (O_734,N_9702,N_9815);
xnor UO_735 (O_735,N_9680,N_9653);
or UO_736 (O_736,N_9939,N_9620);
xnor UO_737 (O_737,N_9987,N_9895);
or UO_738 (O_738,N_9925,N_9691);
xor UO_739 (O_739,N_9841,N_9516);
nand UO_740 (O_740,N_9741,N_9819);
and UO_741 (O_741,N_9755,N_9670);
xor UO_742 (O_742,N_9593,N_9533);
or UO_743 (O_743,N_9714,N_9964);
nand UO_744 (O_744,N_9910,N_9842);
and UO_745 (O_745,N_9749,N_9921);
and UO_746 (O_746,N_9795,N_9635);
nand UO_747 (O_747,N_9550,N_9798);
xor UO_748 (O_748,N_9627,N_9704);
and UO_749 (O_749,N_9638,N_9585);
and UO_750 (O_750,N_9742,N_9658);
nand UO_751 (O_751,N_9712,N_9804);
or UO_752 (O_752,N_9701,N_9599);
and UO_753 (O_753,N_9654,N_9649);
xor UO_754 (O_754,N_9524,N_9902);
nand UO_755 (O_755,N_9849,N_9723);
nor UO_756 (O_756,N_9614,N_9685);
and UO_757 (O_757,N_9669,N_9801);
nand UO_758 (O_758,N_9817,N_9807);
and UO_759 (O_759,N_9539,N_9669);
nand UO_760 (O_760,N_9935,N_9893);
or UO_761 (O_761,N_9761,N_9914);
nor UO_762 (O_762,N_9697,N_9649);
xor UO_763 (O_763,N_9847,N_9852);
nand UO_764 (O_764,N_9838,N_9516);
nand UO_765 (O_765,N_9840,N_9598);
nor UO_766 (O_766,N_9610,N_9551);
xor UO_767 (O_767,N_9809,N_9770);
nand UO_768 (O_768,N_9746,N_9592);
and UO_769 (O_769,N_9764,N_9819);
nor UO_770 (O_770,N_9745,N_9680);
and UO_771 (O_771,N_9679,N_9702);
or UO_772 (O_772,N_9650,N_9558);
and UO_773 (O_773,N_9568,N_9773);
nor UO_774 (O_774,N_9914,N_9871);
or UO_775 (O_775,N_9665,N_9848);
nand UO_776 (O_776,N_9637,N_9713);
nor UO_777 (O_777,N_9687,N_9801);
xnor UO_778 (O_778,N_9506,N_9764);
nand UO_779 (O_779,N_9777,N_9947);
nand UO_780 (O_780,N_9731,N_9859);
nand UO_781 (O_781,N_9518,N_9816);
nand UO_782 (O_782,N_9546,N_9886);
xnor UO_783 (O_783,N_9603,N_9540);
nand UO_784 (O_784,N_9989,N_9673);
and UO_785 (O_785,N_9507,N_9953);
or UO_786 (O_786,N_9835,N_9856);
and UO_787 (O_787,N_9610,N_9634);
and UO_788 (O_788,N_9926,N_9977);
nor UO_789 (O_789,N_9626,N_9911);
and UO_790 (O_790,N_9812,N_9575);
xor UO_791 (O_791,N_9956,N_9646);
nand UO_792 (O_792,N_9747,N_9650);
xor UO_793 (O_793,N_9809,N_9747);
nor UO_794 (O_794,N_9845,N_9643);
xnor UO_795 (O_795,N_9608,N_9532);
nor UO_796 (O_796,N_9853,N_9905);
nor UO_797 (O_797,N_9906,N_9788);
nand UO_798 (O_798,N_9793,N_9852);
and UO_799 (O_799,N_9966,N_9830);
xor UO_800 (O_800,N_9865,N_9733);
and UO_801 (O_801,N_9884,N_9937);
nand UO_802 (O_802,N_9827,N_9529);
nor UO_803 (O_803,N_9778,N_9519);
nand UO_804 (O_804,N_9605,N_9681);
or UO_805 (O_805,N_9839,N_9507);
or UO_806 (O_806,N_9771,N_9647);
and UO_807 (O_807,N_9668,N_9672);
nor UO_808 (O_808,N_9627,N_9673);
and UO_809 (O_809,N_9863,N_9830);
xor UO_810 (O_810,N_9852,N_9598);
nand UO_811 (O_811,N_9860,N_9767);
xnor UO_812 (O_812,N_9934,N_9992);
nand UO_813 (O_813,N_9540,N_9532);
and UO_814 (O_814,N_9757,N_9530);
xnor UO_815 (O_815,N_9831,N_9910);
nor UO_816 (O_816,N_9892,N_9713);
nand UO_817 (O_817,N_9844,N_9685);
nand UO_818 (O_818,N_9858,N_9915);
and UO_819 (O_819,N_9869,N_9553);
or UO_820 (O_820,N_9967,N_9792);
or UO_821 (O_821,N_9675,N_9855);
and UO_822 (O_822,N_9818,N_9648);
xor UO_823 (O_823,N_9707,N_9875);
nor UO_824 (O_824,N_9731,N_9799);
xnor UO_825 (O_825,N_9558,N_9608);
and UO_826 (O_826,N_9549,N_9819);
nor UO_827 (O_827,N_9855,N_9987);
and UO_828 (O_828,N_9956,N_9950);
nor UO_829 (O_829,N_9728,N_9813);
xor UO_830 (O_830,N_9886,N_9701);
and UO_831 (O_831,N_9920,N_9778);
or UO_832 (O_832,N_9574,N_9815);
or UO_833 (O_833,N_9639,N_9951);
and UO_834 (O_834,N_9536,N_9760);
or UO_835 (O_835,N_9630,N_9766);
nor UO_836 (O_836,N_9871,N_9689);
and UO_837 (O_837,N_9796,N_9715);
nand UO_838 (O_838,N_9760,N_9963);
xnor UO_839 (O_839,N_9618,N_9791);
nand UO_840 (O_840,N_9557,N_9567);
xnor UO_841 (O_841,N_9743,N_9892);
or UO_842 (O_842,N_9808,N_9987);
nand UO_843 (O_843,N_9609,N_9671);
and UO_844 (O_844,N_9683,N_9997);
or UO_845 (O_845,N_9521,N_9806);
and UO_846 (O_846,N_9872,N_9818);
nand UO_847 (O_847,N_9621,N_9627);
nor UO_848 (O_848,N_9919,N_9823);
xor UO_849 (O_849,N_9796,N_9548);
or UO_850 (O_850,N_9701,N_9754);
nor UO_851 (O_851,N_9585,N_9820);
nand UO_852 (O_852,N_9577,N_9516);
or UO_853 (O_853,N_9605,N_9592);
xnor UO_854 (O_854,N_9653,N_9883);
nand UO_855 (O_855,N_9557,N_9921);
nand UO_856 (O_856,N_9564,N_9539);
nand UO_857 (O_857,N_9607,N_9599);
xnor UO_858 (O_858,N_9843,N_9944);
nor UO_859 (O_859,N_9963,N_9922);
or UO_860 (O_860,N_9934,N_9819);
nor UO_861 (O_861,N_9644,N_9601);
or UO_862 (O_862,N_9531,N_9723);
nor UO_863 (O_863,N_9577,N_9977);
or UO_864 (O_864,N_9592,N_9789);
and UO_865 (O_865,N_9603,N_9579);
nand UO_866 (O_866,N_9966,N_9840);
or UO_867 (O_867,N_9608,N_9825);
nand UO_868 (O_868,N_9625,N_9618);
nor UO_869 (O_869,N_9567,N_9726);
nor UO_870 (O_870,N_9990,N_9934);
or UO_871 (O_871,N_9852,N_9740);
nand UO_872 (O_872,N_9717,N_9643);
and UO_873 (O_873,N_9507,N_9598);
nor UO_874 (O_874,N_9605,N_9557);
or UO_875 (O_875,N_9562,N_9745);
nor UO_876 (O_876,N_9652,N_9557);
and UO_877 (O_877,N_9996,N_9878);
xor UO_878 (O_878,N_9671,N_9743);
and UO_879 (O_879,N_9993,N_9599);
xnor UO_880 (O_880,N_9796,N_9968);
nand UO_881 (O_881,N_9571,N_9752);
nor UO_882 (O_882,N_9558,N_9579);
xnor UO_883 (O_883,N_9979,N_9588);
nand UO_884 (O_884,N_9877,N_9521);
or UO_885 (O_885,N_9898,N_9679);
xor UO_886 (O_886,N_9917,N_9947);
or UO_887 (O_887,N_9503,N_9995);
xor UO_888 (O_888,N_9791,N_9653);
xor UO_889 (O_889,N_9745,N_9937);
nand UO_890 (O_890,N_9999,N_9640);
nand UO_891 (O_891,N_9949,N_9924);
nor UO_892 (O_892,N_9915,N_9727);
nand UO_893 (O_893,N_9744,N_9946);
nor UO_894 (O_894,N_9905,N_9765);
nand UO_895 (O_895,N_9683,N_9955);
nand UO_896 (O_896,N_9663,N_9512);
or UO_897 (O_897,N_9978,N_9683);
xnor UO_898 (O_898,N_9755,N_9596);
and UO_899 (O_899,N_9754,N_9987);
and UO_900 (O_900,N_9980,N_9925);
xor UO_901 (O_901,N_9697,N_9528);
nor UO_902 (O_902,N_9938,N_9595);
nor UO_903 (O_903,N_9792,N_9698);
nor UO_904 (O_904,N_9906,N_9750);
xnor UO_905 (O_905,N_9903,N_9972);
nor UO_906 (O_906,N_9844,N_9703);
xnor UO_907 (O_907,N_9577,N_9505);
and UO_908 (O_908,N_9896,N_9696);
nand UO_909 (O_909,N_9741,N_9598);
and UO_910 (O_910,N_9531,N_9753);
nand UO_911 (O_911,N_9706,N_9967);
nand UO_912 (O_912,N_9738,N_9935);
and UO_913 (O_913,N_9727,N_9589);
nand UO_914 (O_914,N_9503,N_9886);
xor UO_915 (O_915,N_9550,N_9658);
and UO_916 (O_916,N_9845,N_9674);
nand UO_917 (O_917,N_9995,N_9518);
or UO_918 (O_918,N_9817,N_9647);
xnor UO_919 (O_919,N_9897,N_9635);
nand UO_920 (O_920,N_9502,N_9516);
and UO_921 (O_921,N_9704,N_9719);
nor UO_922 (O_922,N_9818,N_9745);
nor UO_923 (O_923,N_9851,N_9812);
nor UO_924 (O_924,N_9580,N_9666);
nand UO_925 (O_925,N_9992,N_9529);
nor UO_926 (O_926,N_9652,N_9822);
and UO_927 (O_927,N_9740,N_9991);
nor UO_928 (O_928,N_9938,N_9721);
and UO_929 (O_929,N_9864,N_9653);
and UO_930 (O_930,N_9787,N_9645);
nor UO_931 (O_931,N_9614,N_9687);
or UO_932 (O_932,N_9630,N_9891);
nand UO_933 (O_933,N_9971,N_9584);
or UO_934 (O_934,N_9784,N_9694);
nor UO_935 (O_935,N_9509,N_9878);
or UO_936 (O_936,N_9512,N_9808);
or UO_937 (O_937,N_9650,N_9884);
xor UO_938 (O_938,N_9997,N_9776);
nor UO_939 (O_939,N_9799,N_9721);
or UO_940 (O_940,N_9632,N_9943);
nand UO_941 (O_941,N_9820,N_9914);
nand UO_942 (O_942,N_9547,N_9573);
nand UO_943 (O_943,N_9680,N_9658);
xnor UO_944 (O_944,N_9627,N_9708);
or UO_945 (O_945,N_9651,N_9742);
xnor UO_946 (O_946,N_9928,N_9954);
nor UO_947 (O_947,N_9760,N_9789);
xnor UO_948 (O_948,N_9529,N_9678);
xor UO_949 (O_949,N_9755,N_9677);
xnor UO_950 (O_950,N_9970,N_9548);
or UO_951 (O_951,N_9756,N_9581);
xor UO_952 (O_952,N_9793,N_9785);
or UO_953 (O_953,N_9710,N_9816);
and UO_954 (O_954,N_9552,N_9733);
xor UO_955 (O_955,N_9657,N_9559);
and UO_956 (O_956,N_9713,N_9852);
xor UO_957 (O_957,N_9990,N_9952);
or UO_958 (O_958,N_9939,N_9663);
xor UO_959 (O_959,N_9968,N_9950);
nor UO_960 (O_960,N_9527,N_9542);
and UO_961 (O_961,N_9622,N_9500);
nand UO_962 (O_962,N_9659,N_9981);
nor UO_963 (O_963,N_9835,N_9942);
nor UO_964 (O_964,N_9704,N_9692);
nand UO_965 (O_965,N_9718,N_9796);
nand UO_966 (O_966,N_9893,N_9559);
nand UO_967 (O_967,N_9829,N_9524);
nor UO_968 (O_968,N_9876,N_9554);
and UO_969 (O_969,N_9961,N_9601);
nand UO_970 (O_970,N_9908,N_9763);
nand UO_971 (O_971,N_9813,N_9616);
nand UO_972 (O_972,N_9681,N_9632);
nor UO_973 (O_973,N_9694,N_9529);
xor UO_974 (O_974,N_9943,N_9995);
or UO_975 (O_975,N_9531,N_9517);
nand UO_976 (O_976,N_9808,N_9762);
nor UO_977 (O_977,N_9778,N_9703);
nand UO_978 (O_978,N_9824,N_9812);
nor UO_979 (O_979,N_9908,N_9806);
or UO_980 (O_980,N_9796,N_9549);
nand UO_981 (O_981,N_9769,N_9717);
xnor UO_982 (O_982,N_9739,N_9856);
nand UO_983 (O_983,N_9595,N_9624);
and UO_984 (O_984,N_9712,N_9997);
nor UO_985 (O_985,N_9952,N_9764);
or UO_986 (O_986,N_9584,N_9703);
or UO_987 (O_987,N_9591,N_9997);
xor UO_988 (O_988,N_9606,N_9965);
or UO_989 (O_989,N_9706,N_9778);
or UO_990 (O_990,N_9970,N_9629);
xnor UO_991 (O_991,N_9566,N_9897);
or UO_992 (O_992,N_9645,N_9636);
nand UO_993 (O_993,N_9621,N_9523);
or UO_994 (O_994,N_9885,N_9590);
or UO_995 (O_995,N_9596,N_9900);
xor UO_996 (O_996,N_9604,N_9749);
nor UO_997 (O_997,N_9508,N_9766);
nand UO_998 (O_998,N_9850,N_9509);
and UO_999 (O_999,N_9877,N_9537);
or UO_1000 (O_1000,N_9967,N_9763);
nand UO_1001 (O_1001,N_9805,N_9767);
xor UO_1002 (O_1002,N_9776,N_9957);
and UO_1003 (O_1003,N_9930,N_9969);
and UO_1004 (O_1004,N_9984,N_9791);
nand UO_1005 (O_1005,N_9891,N_9965);
nand UO_1006 (O_1006,N_9686,N_9616);
nor UO_1007 (O_1007,N_9622,N_9810);
or UO_1008 (O_1008,N_9772,N_9790);
nand UO_1009 (O_1009,N_9797,N_9631);
xor UO_1010 (O_1010,N_9793,N_9963);
and UO_1011 (O_1011,N_9561,N_9978);
nand UO_1012 (O_1012,N_9665,N_9666);
or UO_1013 (O_1013,N_9706,N_9760);
nor UO_1014 (O_1014,N_9855,N_9919);
nand UO_1015 (O_1015,N_9500,N_9703);
and UO_1016 (O_1016,N_9716,N_9605);
nand UO_1017 (O_1017,N_9942,N_9528);
or UO_1018 (O_1018,N_9895,N_9691);
nand UO_1019 (O_1019,N_9979,N_9653);
xor UO_1020 (O_1020,N_9994,N_9996);
or UO_1021 (O_1021,N_9856,N_9858);
nand UO_1022 (O_1022,N_9508,N_9759);
nor UO_1023 (O_1023,N_9570,N_9638);
nand UO_1024 (O_1024,N_9594,N_9878);
xor UO_1025 (O_1025,N_9654,N_9811);
nand UO_1026 (O_1026,N_9787,N_9743);
nor UO_1027 (O_1027,N_9672,N_9767);
nor UO_1028 (O_1028,N_9760,N_9754);
or UO_1029 (O_1029,N_9892,N_9644);
and UO_1030 (O_1030,N_9656,N_9620);
or UO_1031 (O_1031,N_9825,N_9722);
nand UO_1032 (O_1032,N_9750,N_9694);
nand UO_1033 (O_1033,N_9584,N_9937);
or UO_1034 (O_1034,N_9663,N_9839);
nor UO_1035 (O_1035,N_9552,N_9745);
nor UO_1036 (O_1036,N_9998,N_9673);
xor UO_1037 (O_1037,N_9544,N_9573);
and UO_1038 (O_1038,N_9811,N_9781);
nand UO_1039 (O_1039,N_9540,N_9905);
nand UO_1040 (O_1040,N_9852,N_9944);
and UO_1041 (O_1041,N_9978,N_9856);
and UO_1042 (O_1042,N_9797,N_9723);
nand UO_1043 (O_1043,N_9507,N_9557);
nor UO_1044 (O_1044,N_9634,N_9665);
xnor UO_1045 (O_1045,N_9949,N_9700);
nor UO_1046 (O_1046,N_9718,N_9995);
nand UO_1047 (O_1047,N_9578,N_9968);
and UO_1048 (O_1048,N_9851,N_9840);
and UO_1049 (O_1049,N_9955,N_9550);
or UO_1050 (O_1050,N_9502,N_9537);
xnor UO_1051 (O_1051,N_9706,N_9757);
and UO_1052 (O_1052,N_9564,N_9579);
nand UO_1053 (O_1053,N_9632,N_9904);
xnor UO_1054 (O_1054,N_9660,N_9531);
xnor UO_1055 (O_1055,N_9535,N_9816);
xor UO_1056 (O_1056,N_9885,N_9778);
or UO_1057 (O_1057,N_9948,N_9904);
nand UO_1058 (O_1058,N_9870,N_9560);
and UO_1059 (O_1059,N_9526,N_9648);
nor UO_1060 (O_1060,N_9763,N_9716);
xor UO_1061 (O_1061,N_9564,N_9807);
nor UO_1062 (O_1062,N_9616,N_9858);
nand UO_1063 (O_1063,N_9757,N_9868);
nand UO_1064 (O_1064,N_9756,N_9604);
and UO_1065 (O_1065,N_9990,N_9994);
nor UO_1066 (O_1066,N_9566,N_9799);
nand UO_1067 (O_1067,N_9848,N_9620);
or UO_1068 (O_1068,N_9851,N_9583);
or UO_1069 (O_1069,N_9613,N_9835);
nand UO_1070 (O_1070,N_9902,N_9787);
nand UO_1071 (O_1071,N_9695,N_9575);
or UO_1072 (O_1072,N_9902,N_9736);
or UO_1073 (O_1073,N_9788,N_9661);
nand UO_1074 (O_1074,N_9788,N_9777);
nand UO_1075 (O_1075,N_9715,N_9869);
nand UO_1076 (O_1076,N_9714,N_9955);
nand UO_1077 (O_1077,N_9807,N_9814);
nor UO_1078 (O_1078,N_9728,N_9600);
nor UO_1079 (O_1079,N_9771,N_9535);
and UO_1080 (O_1080,N_9895,N_9907);
and UO_1081 (O_1081,N_9750,N_9861);
xnor UO_1082 (O_1082,N_9731,N_9526);
nand UO_1083 (O_1083,N_9687,N_9842);
or UO_1084 (O_1084,N_9589,N_9821);
xor UO_1085 (O_1085,N_9578,N_9956);
or UO_1086 (O_1086,N_9927,N_9601);
xor UO_1087 (O_1087,N_9575,N_9760);
xnor UO_1088 (O_1088,N_9665,N_9798);
and UO_1089 (O_1089,N_9775,N_9988);
or UO_1090 (O_1090,N_9889,N_9569);
and UO_1091 (O_1091,N_9622,N_9909);
xnor UO_1092 (O_1092,N_9894,N_9722);
nor UO_1093 (O_1093,N_9719,N_9607);
or UO_1094 (O_1094,N_9822,N_9955);
nand UO_1095 (O_1095,N_9882,N_9737);
nor UO_1096 (O_1096,N_9997,N_9973);
nor UO_1097 (O_1097,N_9714,N_9720);
and UO_1098 (O_1098,N_9867,N_9500);
or UO_1099 (O_1099,N_9545,N_9748);
nor UO_1100 (O_1100,N_9598,N_9590);
and UO_1101 (O_1101,N_9648,N_9536);
xor UO_1102 (O_1102,N_9836,N_9713);
nor UO_1103 (O_1103,N_9979,N_9944);
nor UO_1104 (O_1104,N_9897,N_9615);
and UO_1105 (O_1105,N_9846,N_9638);
or UO_1106 (O_1106,N_9718,N_9755);
nand UO_1107 (O_1107,N_9670,N_9868);
or UO_1108 (O_1108,N_9922,N_9882);
nand UO_1109 (O_1109,N_9785,N_9922);
or UO_1110 (O_1110,N_9579,N_9662);
and UO_1111 (O_1111,N_9663,N_9708);
xnor UO_1112 (O_1112,N_9627,N_9535);
and UO_1113 (O_1113,N_9757,N_9562);
xor UO_1114 (O_1114,N_9921,N_9808);
or UO_1115 (O_1115,N_9560,N_9537);
and UO_1116 (O_1116,N_9999,N_9601);
or UO_1117 (O_1117,N_9854,N_9508);
nor UO_1118 (O_1118,N_9852,N_9734);
and UO_1119 (O_1119,N_9702,N_9598);
or UO_1120 (O_1120,N_9915,N_9792);
and UO_1121 (O_1121,N_9939,N_9863);
and UO_1122 (O_1122,N_9996,N_9884);
nor UO_1123 (O_1123,N_9862,N_9519);
nand UO_1124 (O_1124,N_9711,N_9777);
nand UO_1125 (O_1125,N_9641,N_9951);
xnor UO_1126 (O_1126,N_9656,N_9995);
or UO_1127 (O_1127,N_9976,N_9659);
nand UO_1128 (O_1128,N_9536,N_9606);
nand UO_1129 (O_1129,N_9600,N_9577);
nand UO_1130 (O_1130,N_9625,N_9656);
or UO_1131 (O_1131,N_9733,N_9797);
nand UO_1132 (O_1132,N_9696,N_9762);
or UO_1133 (O_1133,N_9817,N_9853);
xor UO_1134 (O_1134,N_9680,N_9616);
xor UO_1135 (O_1135,N_9682,N_9918);
nand UO_1136 (O_1136,N_9661,N_9889);
or UO_1137 (O_1137,N_9760,N_9731);
or UO_1138 (O_1138,N_9576,N_9931);
xnor UO_1139 (O_1139,N_9561,N_9932);
nand UO_1140 (O_1140,N_9872,N_9888);
nand UO_1141 (O_1141,N_9624,N_9946);
or UO_1142 (O_1142,N_9930,N_9977);
nor UO_1143 (O_1143,N_9523,N_9628);
xnor UO_1144 (O_1144,N_9762,N_9787);
and UO_1145 (O_1145,N_9548,N_9735);
nand UO_1146 (O_1146,N_9611,N_9757);
and UO_1147 (O_1147,N_9551,N_9746);
xor UO_1148 (O_1148,N_9634,N_9550);
or UO_1149 (O_1149,N_9536,N_9793);
nand UO_1150 (O_1150,N_9658,N_9970);
and UO_1151 (O_1151,N_9839,N_9906);
xor UO_1152 (O_1152,N_9572,N_9819);
nand UO_1153 (O_1153,N_9927,N_9872);
nor UO_1154 (O_1154,N_9932,N_9590);
nor UO_1155 (O_1155,N_9910,N_9939);
xnor UO_1156 (O_1156,N_9554,N_9615);
and UO_1157 (O_1157,N_9690,N_9742);
xor UO_1158 (O_1158,N_9868,N_9584);
and UO_1159 (O_1159,N_9640,N_9950);
nand UO_1160 (O_1160,N_9668,N_9650);
xor UO_1161 (O_1161,N_9513,N_9955);
xnor UO_1162 (O_1162,N_9978,N_9593);
xnor UO_1163 (O_1163,N_9600,N_9860);
nand UO_1164 (O_1164,N_9931,N_9749);
or UO_1165 (O_1165,N_9840,N_9913);
and UO_1166 (O_1166,N_9541,N_9630);
nand UO_1167 (O_1167,N_9516,N_9661);
nand UO_1168 (O_1168,N_9999,N_9576);
xnor UO_1169 (O_1169,N_9703,N_9950);
nor UO_1170 (O_1170,N_9724,N_9695);
or UO_1171 (O_1171,N_9955,N_9993);
nor UO_1172 (O_1172,N_9540,N_9815);
or UO_1173 (O_1173,N_9937,N_9587);
xor UO_1174 (O_1174,N_9585,N_9915);
nand UO_1175 (O_1175,N_9784,N_9976);
or UO_1176 (O_1176,N_9756,N_9889);
and UO_1177 (O_1177,N_9823,N_9909);
and UO_1178 (O_1178,N_9962,N_9979);
or UO_1179 (O_1179,N_9532,N_9916);
nand UO_1180 (O_1180,N_9648,N_9701);
nor UO_1181 (O_1181,N_9830,N_9908);
nand UO_1182 (O_1182,N_9582,N_9949);
nor UO_1183 (O_1183,N_9861,N_9819);
and UO_1184 (O_1184,N_9766,N_9538);
or UO_1185 (O_1185,N_9750,N_9836);
nor UO_1186 (O_1186,N_9936,N_9727);
xor UO_1187 (O_1187,N_9520,N_9962);
nand UO_1188 (O_1188,N_9800,N_9585);
nand UO_1189 (O_1189,N_9626,N_9746);
or UO_1190 (O_1190,N_9546,N_9836);
or UO_1191 (O_1191,N_9905,N_9628);
nand UO_1192 (O_1192,N_9774,N_9693);
nand UO_1193 (O_1193,N_9739,N_9727);
and UO_1194 (O_1194,N_9849,N_9985);
nand UO_1195 (O_1195,N_9504,N_9719);
or UO_1196 (O_1196,N_9592,N_9808);
nor UO_1197 (O_1197,N_9975,N_9837);
nor UO_1198 (O_1198,N_9772,N_9541);
nand UO_1199 (O_1199,N_9642,N_9987);
nand UO_1200 (O_1200,N_9988,N_9939);
and UO_1201 (O_1201,N_9691,N_9884);
xor UO_1202 (O_1202,N_9567,N_9747);
xor UO_1203 (O_1203,N_9737,N_9730);
nor UO_1204 (O_1204,N_9937,N_9783);
xor UO_1205 (O_1205,N_9612,N_9935);
nor UO_1206 (O_1206,N_9849,N_9994);
nand UO_1207 (O_1207,N_9841,N_9709);
or UO_1208 (O_1208,N_9976,N_9909);
xnor UO_1209 (O_1209,N_9682,N_9555);
nor UO_1210 (O_1210,N_9851,N_9732);
nand UO_1211 (O_1211,N_9820,N_9907);
or UO_1212 (O_1212,N_9826,N_9752);
nand UO_1213 (O_1213,N_9801,N_9862);
xnor UO_1214 (O_1214,N_9655,N_9940);
and UO_1215 (O_1215,N_9603,N_9900);
or UO_1216 (O_1216,N_9990,N_9855);
and UO_1217 (O_1217,N_9637,N_9917);
nand UO_1218 (O_1218,N_9509,N_9778);
or UO_1219 (O_1219,N_9784,N_9682);
nor UO_1220 (O_1220,N_9805,N_9983);
and UO_1221 (O_1221,N_9810,N_9984);
nand UO_1222 (O_1222,N_9730,N_9771);
nand UO_1223 (O_1223,N_9542,N_9780);
and UO_1224 (O_1224,N_9538,N_9947);
nand UO_1225 (O_1225,N_9889,N_9790);
nor UO_1226 (O_1226,N_9756,N_9800);
xor UO_1227 (O_1227,N_9965,N_9569);
nor UO_1228 (O_1228,N_9916,N_9828);
nor UO_1229 (O_1229,N_9653,N_9591);
or UO_1230 (O_1230,N_9622,N_9736);
and UO_1231 (O_1231,N_9724,N_9638);
or UO_1232 (O_1232,N_9565,N_9881);
and UO_1233 (O_1233,N_9767,N_9512);
xnor UO_1234 (O_1234,N_9949,N_9937);
xor UO_1235 (O_1235,N_9711,N_9762);
and UO_1236 (O_1236,N_9629,N_9898);
nor UO_1237 (O_1237,N_9821,N_9614);
and UO_1238 (O_1238,N_9557,N_9851);
xor UO_1239 (O_1239,N_9870,N_9744);
nor UO_1240 (O_1240,N_9559,N_9508);
and UO_1241 (O_1241,N_9590,N_9747);
nand UO_1242 (O_1242,N_9611,N_9867);
or UO_1243 (O_1243,N_9662,N_9924);
and UO_1244 (O_1244,N_9809,N_9921);
nand UO_1245 (O_1245,N_9642,N_9604);
xnor UO_1246 (O_1246,N_9562,N_9841);
xor UO_1247 (O_1247,N_9833,N_9961);
and UO_1248 (O_1248,N_9818,N_9678);
and UO_1249 (O_1249,N_9753,N_9569);
xor UO_1250 (O_1250,N_9507,N_9636);
nor UO_1251 (O_1251,N_9622,N_9595);
nor UO_1252 (O_1252,N_9895,N_9696);
xnor UO_1253 (O_1253,N_9996,N_9557);
and UO_1254 (O_1254,N_9617,N_9879);
or UO_1255 (O_1255,N_9826,N_9936);
and UO_1256 (O_1256,N_9764,N_9721);
or UO_1257 (O_1257,N_9602,N_9940);
or UO_1258 (O_1258,N_9522,N_9957);
and UO_1259 (O_1259,N_9544,N_9557);
and UO_1260 (O_1260,N_9550,N_9829);
and UO_1261 (O_1261,N_9738,N_9852);
or UO_1262 (O_1262,N_9874,N_9615);
xor UO_1263 (O_1263,N_9709,N_9521);
nor UO_1264 (O_1264,N_9903,N_9545);
nand UO_1265 (O_1265,N_9500,N_9524);
nor UO_1266 (O_1266,N_9863,N_9682);
nor UO_1267 (O_1267,N_9617,N_9687);
or UO_1268 (O_1268,N_9594,N_9810);
or UO_1269 (O_1269,N_9899,N_9588);
nor UO_1270 (O_1270,N_9588,N_9587);
and UO_1271 (O_1271,N_9991,N_9639);
xnor UO_1272 (O_1272,N_9838,N_9529);
nand UO_1273 (O_1273,N_9551,N_9873);
nor UO_1274 (O_1274,N_9504,N_9743);
xnor UO_1275 (O_1275,N_9668,N_9530);
or UO_1276 (O_1276,N_9557,N_9684);
or UO_1277 (O_1277,N_9651,N_9758);
and UO_1278 (O_1278,N_9526,N_9607);
or UO_1279 (O_1279,N_9513,N_9998);
or UO_1280 (O_1280,N_9713,N_9691);
nand UO_1281 (O_1281,N_9844,N_9764);
nand UO_1282 (O_1282,N_9774,N_9736);
or UO_1283 (O_1283,N_9948,N_9699);
nor UO_1284 (O_1284,N_9623,N_9885);
xnor UO_1285 (O_1285,N_9583,N_9624);
nor UO_1286 (O_1286,N_9980,N_9770);
or UO_1287 (O_1287,N_9905,N_9800);
nand UO_1288 (O_1288,N_9811,N_9925);
nor UO_1289 (O_1289,N_9583,N_9891);
and UO_1290 (O_1290,N_9905,N_9908);
and UO_1291 (O_1291,N_9971,N_9707);
nor UO_1292 (O_1292,N_9674,N_9984);
or UO_1293 (O_1293,N_9696,N_9685);
nor UO_1294 (O_1294,N_9961,N_9581);
nand UO_1295 (O_1295,N_9627,N_9720);
and UO_1296 (O_1296,N_9945,N_9938);
nand UO_1297 (O_1297,N_9633,N_9521);
and UO_1298 (O_1298,N_9510,N_9655);
xnor UO_1299 (O_1299,N_9660,N_9778);
and UO_1300 (O_1300,N_9690,N_9555);
or UO_1301 (O_1301,N_9904,N_9839);
and UO_1302 (O_1302,N_9646,N_9555);
xnor UO_1303 (O_1303,N_9630,N_9574);
nand UO_1304 (O_1304,N_9784,N_9581);
nand UO_1305 (O_1305,N_9789,N_9752);
and UO_1306 (O_1306,N_9962,N_9600);
or UO_1307 (O_1307,N_9680,N_9896);
xnor UO_1308 (O_1308,N_9586,N_9952);
nor UO_1309 (O_1309,N_9754,N_9621);
and UO_1310 (O_1310,N_9625,N_9878);
nor UO_1311 (O_1311,N_9902,N_9603);
and UO_1312 (O_1312,N_9511,N_9600);
xor UO_1313 (O_1313,N_9989,N_9535);
or UO_1314 (O_1314,N_9712,N_9677);
xor UO_1315 (O_1315,N_9783,N_9543);
nand UO_1316 (O_1316,N_9924,N_9910);
and UO_1317 (O_1317,N_9637,N_9569);
nor UO_1318 (O_1318,N_9776,N_9991);
and UO_1319 (O_1319,N_9795,N_9926);
nor UO_1320 (O_1320,N_9814,N_9981);
and UO_1321 (O_1321,N_9877,N_9551);
nor UO_1322 (O_1322,N_9734,N_9575);
nor UO_1323 (O_1323,N_9625,N_9580);
nand UO_1324 (O_1324,N_9605,N_9607);
nand UO_1325 (O_1325,N_9682,N_9525);
nor UO_1326 (O_1326,N_9698,N_9641);
and UO_1327 (O_1327,N_9961,N_9927);
nand UO_1328 (O_1328,N_9557,N_9580);
and UO_1329 (O_1329,N_9808,N_9711);
or UO_1330 (O_1330,N_9888,N_9696);
xnor UO_1331 (O_1331,N_9927,N_9587);
xor UO_1332 (O_1332,N_9992,N_9826);
xor UO_1333 (O_1333,N_9502,N_9829);
or UO_1334 (O_1334,N_9701,N_9523);
nand UO_1335 (O_1335,N_9831,N_9722);
nor UO_1336 (O_1336,N_9826,N_9528);
or UO_1337 (O_1337,N_9826,N_9817);
or UO_1338 (O_1338,N_9948,N_9885);
nand UO_1339 (O_1339,N_9939,N_9802);
xnor UO_1340 (O_1340,N_9856,N_9832);
nor UO_1341 (O_1341,N_9655,N_9959);
and UO_1342 (O_1342,N_9617,N_9950);
and UO_1343 (O_1343,N_9922,N_9660);
and UO_1344 (O_1344,N_9794,N_9806);
and UO_1345 (O_1345,N_9689,N_9515);
nand UO_1346 (O_1346,N_9523,N_9648);
or UO_1347 (O_1347,N_9698,N_9853);
and UO_1348 (O_1348,N_9925,N_9739);
nor UO_1349 (O_1349,N_9909,N_9693);
nand UO_1350 (O_1350,N_9848,N_9833);
nand UO_1351 (O_1351,N_9500,N_9774);
xor UO_1352 (O_1352,N_9793,N_9838);
nand UO_1353 (O_1353,N_9888,N_9752);
xor UO_1354 (O_1354,N_9711,N_9820);
or UO_1355 (O_1355,N_9950,N_9974);
xnor UO_1356 (O_1356,N_9626,N_9856);
xor UO_1357 (O_1357,N_9627,N_9501);
and UO_1358 (O_1358,N_9602,N_9734);
xnor UO_1359 (O_1359,N_9780,N_9859);
or UO_1360 (O_1360,N_9934,N_9531);
nor UO_1361 (O_1361,N_9757,N_9977);
nor UO_1362 (O_1362,N_9950,N_9537);
or UO_1363 (O_1363,N_9645,N_9809);
and UO_1364 (O_1364,N_9576,N_9605);
and UO_1365 (O_1365,N_9637,N_9861);
nor UO_1366 (O_1366,N_9595,N_9726);
nor UO_1367 (O_1367,N_9657,N_9947);
nand UO_1368 (O_1368,N_9713,N_9529);
nor UO_1369 (O_1369,N_9696,N_9869);
and UO_1370 (O_1370,N_9765,N_9522);
nor UO_1371 (O_1371,N_9761,N_9716);
xnor UO_1372 (O_1372,N_9646,N_9717);
nand UO_1373 (O_1373,N_9954,N_9912);
or UO_1374 (O_1374,N_9862,N_9717);
nor UO_1375 (O_1375,N_9777,N_9735);
and UO_1376 (O_1376,N_9515,N_9990);
or UO_1377 (O_1377,N_9744,N_9869);
nor UO_1378 (O_1378,N_9726,N_9851);
nand UO_1379 (O_1379,N_9556,N_9812);
and UO_1380 (O_1380,N_9975,N_9945);
or UO_1381 (O_1381,N_9552,N_9926);
xor UO_1382 (O_1382,N_9961,N_9955);
or UO_1383 (O_1383,N_9963,N_9737);
and UO_1384 (O_1384,N_9940,N_9540);
nor UO_1385 (O_1385,N_9923,N_9667);
and UO_1386 (O_1386,N_9613,N_9569);
or UO_1387 (O_1387,N_9505,N_9971);
and UO_1388 (O_1388,N_9500,N_9866);
nand UO_1389 (O_1389,N_9536,N_9823);
nor UO_1390 (O_1390,N_9762,N_9880);
and UO_1391 (O_1391,N_9746,N_9842);
and UO_1392 (O_1392,N_9641,N_9950);
xor UO_1393 (O_1393,N_9525,N_9500);
and UO_1394 (O_1394,N_9644,N_9593);
nand UO_1395 (O_1395,N_9709,N_9970);
nand UO_1396 (O_1396,N_9736,N_9670);
xor UO_1397 (O_1397,N_9516,N_9753);
xnor UO_1398 (O_1398,N_9833,N_9958);
nor UO_1399 (O_1399,N_9762,N_9959);
nor UO_1400 (O_1400,N_9714,N_9724);
or UO_1401 (O_1401,N_9853,N_9957);
nor UO_1402 (O_1402,N_9600,N_9652);
xor UO_1403 (O_1403,N_9781,N_9662);
or UO_1404 (O_1404,N_9873,N_9977);
nand UO_1405 (O_1405,N_9676,N_9660);
and UO_1406 (O_1406,N_9995,N_9852);
nand UO_1407 (O_1407,N_9793,N_9951);
nor UO_1408 (O_1408,N_9875,N_9538);
nand UO_1409 (O_1409,N_9945,N_9790);
xor UO_1410 (O_1410,N_9603,N_9878);
xor UO_1411 (O_1411,N_9758,N_9851);
xnor UO_1412 (O_1412,N_9864,N_9993);
nand UO_1413 (O_1413,N_9662,N_9925);
xnor UO_1414 (O_1414,N_9996,N_9759);
nand UO_1415 (O_1415,N_9930,N_9542);
xnor UO_1416 (O_1416,N_9812,N_9543);
xor UO_1417 (O_1417,N_9675,N_9821);
xor UO_1418 (O_1418,N_9772,N_9788);
or UO_1419 (O_1419,N_9755,N_9662);
xor UO_1420 (O_1420,N_9529,N_9729);
xor UO_1421 (O_1421,N_9815,N_9820);
nor UO_1422 (O_1422,N_9813,N_9605);
and UO_1423 (O_1423,N_9711,N_9978);
nor UO_1424 (O_1424,N_9609,N_9694);
xnor UO_1425 (O_1425,N_9908,N_9616);
nor UO_1426 (O_1426,N_9620,N_9592);
and UO_1427 (O_1427,N_9745,N_9623);
nor UO_1428 (O_1428,N_9904,N_9574);
or UO_1429 (O_1429,N_9969,N_9725);
nand UO_1430 (O_1430,N_9991,N_9758);
nor UO_1431 (O_1431,N_9583,N_9885);
or UO_1432 (O_1432,N_9680,N_9977);
nand UO_1433 (O_1433,N_9843,N_9998);
nand UO_1434 (O_1434,N_9684,N_9538);
or UO_1435 (O_1435,N_9806,N_9867);
nand UO_1436 (O_1436,N_9657,N_9638);
nand UO_1437 (O_1437,N_9630,N_9838);
xnor UO_1438 (O_1438,N_9967,N_9749);
nand UO_1439 (O_1439,N_9655,N_9981);
nand UO_1440 (O_1440,N_9510,N_9832);
xor UO_1441 (O_1441,N_9815,N_9761);
or UO_1442 (O_1442,N_9772,N_9959);
nor UO_1443 (O_1443,N_9540,N_9968);
and UO_1444 (O_1444,N_9993,N_9555);
nor UO_1445 (O_1445,N_9846,N_9630);
xnor UO_1446 (O_1446,N_9927,N_9713);
and UO_1447 (O_1447,N_9605,N_9622);
or UO_1448 (O_1448,N_9768,N_9699);
and UO_1449 (O_1449,N_9937,N_9672);
and UO_1450 (O_1450,N_9999,N_9504);
or UO_1451 (O_1451,N_9915,N_9572);
xnor UO_1452 (O_1452,N_9993,N_9753);
nor UO_1453 (O_1453,N_9523,N_9849);
nor UO_1454 (O_1454,N_9988,N_9681);
xor UO_1455 (O_1455,N_9807,N_9593);
xor UO_1456 (O_1456,N_9636,N_9740);
and UO_1457 (O_1457,N_9807,N_9871);
nand UO_1458 (O_1458,N_9842,N_9666);
or UO_1459 (O_1459,N_9994,N_9654);
and UO_1460 (O_1460,N_9927,N_9522);
and UO_1461 (O_1461,N_9913,N_9615);
nor UO_1462 (O_1462,N_9950,N_9685);
nor UO_1463 (O_1463,N_9932,N_9929);
nand UO_1464 (O_1464,N_9844,N_9853);
xnor UO_1465 (O_1465,N_9736,N_9867);
xor UO_1466 (O_1466,N_9531,N_9727);
nor UO_1467 (O_1467,N_9574,N_9739);
and UO_1468 (O_1468,N_9887,N_9773);
or UO_1469 (O_1469,N_9932,N_9909);
xnor UO_1470 (O_1470,N_9615,N_9761);
and UO_1471 (O_1471,N_9509,N_9738);
xnor UO_1472 (O_1472,N_9711,N_9581);
xor UO_1473 (O_1473,N_9681,N_9664);
or UO_1474 (O_1474,N_9852,N_9854);
nand UO_1475 (O_1475,N_9526,N_9846);
nand UO_1476 (O_1476,N_9980,N_9777);
nor UO_1477 (O_1477,N_9922,N_9952);
nor UO_1478 (O_1478,N_9729,N_9860);
and UO_1479 (O_1479,N_9806,N_9518);
xor UO_1480 (O_1480,N_9667,N_9797);
or UO_1481 (O_1481,N_9742,N_9574);
nor UO_1482 (O_1482,N_9535,N_9662);
nor UO_1483 (O_1483,N_9631,N_9534);
nand UO_1484 (O_1484,N_9959,N_9797);
or UO_1485 (O_1485,N_9518,N_9911);
nor UO_1486 (O_1486,N_9898,N_9550);
and UO_1487 (O_1487,N_9823,N_9753);
nor UO_1488 (O_1488,N_9849,N_9508);
nor UO_1489 (O_1489,N_9872,N_9765);
and UO_1490 (O_1490,N_9964,N_9712);
nor UO_1491 (O_1491,N_9842,N_9515);
or UO_1492 (O_1492,N_9536,N_9910);
xnor UO_1493 (O_1493,N_9815,N_9778);
or UO_1494 (O_1494,N_9981,N_9951);
xor UO_1495 (O_1495,N_9917,N_9791);
nand UO_1496 (O_1496,N_9529,N_9940);
nand UO_1497 (O_1497,N_9574,N_9977);
xor UO_1498 (O_1498,N_9798,N_9618);
and UO_1499 (O_1499,N_9536,N_9828);
endmodule