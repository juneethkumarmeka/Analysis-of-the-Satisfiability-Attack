module basic_1500_15000_2000_3_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10035,N_10038,N_10039,N_10040,N_10041,N_10043,N_10044,N_10046,N_10047,N_10048,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10057,N_10058,N_10060,N_10061,N_10062,N_10064,N_10066,N_10067,N_10068,N_10071,N_10072,N_10074,N_10075,N_10076,N_10077,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10093,N_10094,N_10096,N_10097,N_10098,N_10099,N_10100,N_10103,N_10105,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10114,N_10115,N_10118,N_10119,N_10120,N_10121,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10145,N_10146,N_10148,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10167,N_10169,N_10170,N_10172,N_10174,N_10176,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10188,N_10189,N_10190,N_10192,N_10193,N_10194,N_10195,N_10196,N_10198,N_10199,N_10201,N_10202,N_10203,N_10204,N_10205,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10257,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10269,N_10270,N_10274,N_10275,N_10276,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10292,N_10293,N_10294,N_10296,N_10297,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10308,N_10309,N_10310,N_10311,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10324,N_10325,N_10327,N_10328,N_10329,N_10330,N_10332,N_10333,N_10334,N_10335,N_10336,N_10338,N_10339,N_10340,N_10341,N_10342,N_10344,N_10345,N_10346,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10358,N_10359,N_10360,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10374,N_10375,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10387,N_10389,N_10390,N_10391,N_10392,N_10393,N_10395,N_10397,N_10398,N_10399,N_10401,N_10402,N_10404,N_10406,N_10407,N_10408,N_10409,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10418,N_10419,N_10421,N_10422,N_10424,N_10425,N_10426,N_10428,N_10430,N_10431,N_10432,N_10434,N_10435,N_10436,N_10438,N_10440,N_10441,N_10442,N_10443,N_10445,N_10446,N_10447,N_10448,N_10449,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10466,N_10467,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10493,N_10494,N_10495,N_10498,N_10499,N_10501,N_10502,N_10504,N_10505,N_10506,N_10507,N_10508,N_10510,N_10512,N_10513,N_10514,N_10515,N_10516,N_10519,N_10520,N_10521,N_10522,N_10524,N_10527,N_10529,N_10532,N_10533,N_10534,N_10535,N_10536,N_10538,N_10539,N_10540,N_10541,N_10546,N_10547,N_10548,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10564,N_10565,N_10566,N_10567,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10577,N_10578,N_10579,N_10580,N_10581,N_10583,N_10584,N_10587,N_10588,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10617,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10627,N_10628,N_10630,N_10631,N_10632,N_10634,N_10636,N_10639,N_10641,N_10642,N_10643,N_10644,N_10646,N_10647,N_10648,N_10649,N_10653,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10664,N_10665,N_10667,N_10669,N_10670,N_10671,N_10672,N_10674,N_10676,N_10678,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10697,N_10699,N_10700,N_10701,N_10703,N_10704,N_10706,N_10708,N_10709,N_10710,N_10711,N_10713,N_10714,N_10716,N_10717,N_10718,N_10719,N_10720,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10740,N_10741,N_10742,N_10745,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10759,N_10760,N_10761,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10770,N_10771,N_10772,N_10773,N_10777,N_10778,N_10781,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10791,N_10792,N_10793,N_10795,N_10796,N_10797,N_10798,N_10800,N_10801,N_10802,N_10803,N_10805,N_10807,N_10808,N_10809,N_10810,N_10811,N_10813,N_10814,N_10817,N_10818,N_10821,N_10822,N_10823,N_10825,N_10826,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10841,N_10843,N_10844,N_10845,N_10850,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10861,N_10862,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10874,N_10876,N_10878,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10890,N_10892,N_10893,N_10895,N_10896,N_10897,N_10900,N_10901,N_10903,N_10904,N_10905,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10922,N_10923,N_10924,N_10925,N_10928,N_10929,N_10930,N_10931,N_10934,N_10935,N_10936,N_10938,N_10939,N_10940,N_10941,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10961,N_10962,N_10963,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10991,N_10992,N_10993,N_10994,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11009,N_11010,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11030,N_11031,N_11032,N_11036,N_11038,N_11040,N_11041,N_11042,N_11043,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11053,N_11054,N_11055,N_11056,N_11058,N_11059,N_11060,N_11061,N_11062,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11085,N_11087,N_11088,N_11089,N_11092,N_11093,N_11094,N_11095,N_11097,N_11098,N_11099,N_11100,N_11101,N_11103,N_11104,N_11105,N_11106,N_11107,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11137,N_11138,N_11139,N_11140,N_11141,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11153,N_11154,N_11156,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11181,N_11183,N_11184,N_11185,N_11186,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11225,N_11226,N_11227,N_11228,N_11230,N_11231,N_11233,N_11235,N_11236,N_11237,N_11238,N_11240,N_11242,N_11243,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11272,N_11274,N_11275,N_11276,N_11279,N_11280,N_11281,N_11282,N_11284,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11294,N_11295,N_11296,N_11297,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11330,N_11331,N_11332,N_11333,N_11334,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11378,N_11379,N_11380,N_11381,N_11382,N_11384,N_11385,N_11386,N_11387,N_11388,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11400,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11411,N_11412,N_11413,N_11414,N_11417,N_11419,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11437,N_11438,N_11439,N_11441,N_11443,N_11444,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11474,N_11475,N_11476,N_11478,N_11480,N_11481,N_11483,N_11484,N_11485,N_11486,N_11487,N_11489,N_11490,N_11491,N_11493,N_11494,N_11497,N_11498,N_11499,N_11500,N_11503,N_11504,N_11505,N_11506,N_11507,N_11509,N_11510,N_11511,N_11512,N_11514,N_11515,N_11518,N_11519,N_11520,N_11521,N_11522,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11548,N_11549,N_11550,N_11551,N_11552,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11561,N_11562,N_11563,N_11564,N_11566,N_11567,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11577,N_11578,N_11579,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11626,N_11627,N_11628,N_11631,N_11632,N_11633,N_11635,N_11636,N_11637,N_11638,N_11640,N_11641,N_11642,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11653,N_11654,N_11655,N_11656,N_11659,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11677,N_11678,N_11680,N_11681,N_11682,N_11683,N_11685,N_11687,N_11688,N_11689,N_11690,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11713,N_11714,N_11715,N_11717,N_11718,N_11719,N_11720,N_11722,N_11724,N_11725,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11742,N_11744,N_11745,N_11746,N_11750,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11763,N_11764,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11790,N_11791,N_11793,N_11794,N_11795,N_11797,N_11799,N_11800,N_11801,N_11803,N_11804,N_11806,N_11807,N_11808,N_11809,N_11810,N_11812,N_11813,N_11814,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11824,N_11825,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11839,N_11841,N_11842,N_11843,N_11844,N_11846,N_11847,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11865,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11892,N_11893,N_11894,N_11895,N_11896,N_11898,N_11899,N_11900,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11921,N_11922,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11932,N_11933,N_11934,N_11935,N_11936,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11948,N_11949,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11969,N_11970,N_11972,N_11973,N_11974,N_11976,N_11977,N_11978,N_11979,N_11980,N_11982,N_11983,N_11984,N_11985,N_11987,N_11988,N_11989,N_11990,N_11991,N_11993,N_11994,N_11995,N_11998,N_11999,N_12000,N_12001,N_12003,N_12004,N_12005,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12018,N_12019,N_12020,N_12021,N_12022,N_12025,N_12026,N_12027,N_12028,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12038,N_12039,N_12041,N_12042,N_12043,N_12044,N_12045,N_12047,N_12048,N_12049,N_12050,N_12051,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12065,N_12066,N_12067,N_12068,N_12069,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12098,N_12100,N_12101,N_12102,N_12104,N_12105,N_12106,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12116,N_12117,N_12119,N_12120,N_12121,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12158,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12182,N_12183,N_12184,N_12186,N_12187,N_12188,N_12189,N_12190,N_12193,N_12194,N_12195,N_12196,N_12198,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12217,N_12218,N_12219,N_12220,N_12221,N_12224,N_12225,N_12227,N_12228,N_12230,N_12231,N_12233,N_12234,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12244,N_12246,N_12247,N_12249,N_12250,N_12251,N_12252,N_12254,N_12255,N_12258,N_12260,N_12262,N_12263,N_12264,N_12265,N_12267,N_12268,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12285,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12325,N_12326,N_12327,N_12329,N_12331,N_12332,N_12333,N_12337,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12364,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12376,N_12377,N_12378,N_12379,N_12380,N_12383,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12395,N_12396,N_12398,N_12399,N_12400,N_12401,N_12402,N_12404,N_12406,N_12407,N_12408,N_12409,N_12411,N_12412,N_12413,N_12414,N_12415,N_12417,N_12418,N_12419,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12433,N_12435,N_12436,N_12437,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12455,N_12457,N_12458,N_12462,N_12464,N_12465,N_12466,N_12468,N_12469,N_12470,N_12471,N_12472,N_12476,N_12477,N_12478,N_12479,N_12480,N_12482,N_12483,N_12484,N_12487,N_12488,N_12490,N_12491,N_12492,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12531,N_12532,N_12533,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12555,N_12556,N_12557,N_12558,N_12560,N_12561,N_12562,N_12564,N_12565,N_12566,N_12567,N_12568,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12582,N_12583,N_12584,N_12585,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12594,N_12595,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12605,N_12606,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12616,N_12617,N_12618,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12641,N_12644,N_12645,N_12646,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12686,N_12688,N_12690,N_12693,N_12694,N_12695,N_12696,N_12698,N_12699,N_12700,N_12703,N_12704,N_12705,N_12707,N_12708,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12721,N_12723,N_12725,N_12726,N_12727,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12742,N_12743,N_12745,N_12746,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12767,N_12768,N_12769,N_12770,N_12771,N_12773,N_12774,N_12775,N_12776,N_12777,N_12779,N_12780,N_12781,N_12782,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12793,N_12795,N_12796,N_12797,N_12798,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12818,N_12819,N_12820,N_12821,N_12823,N_12824,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12835,N_12836,N_12837,N_12838,N_12839,N_12842,N_12843,N_12844,N_12845,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12860,N_12861,N_12862,N_12863,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12875,N_12876,N_12879,N_12880,N_12881,N_12883,N_12884,N_12886,N_12887,N_12888,N_12889,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12913,N_12915,N_12916,N_12917,N_12918,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12979,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12999,N_13000,N_13001,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13014,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13025,N_13027,N_13028,N_13030,N_13031,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13054,N_13055,N_13056,N_13059,N_13060,N_13061,N_13063,N_13064,N_13065,N_13066,N_13068,N_13069,N_13070,N_13072,N_13073,N_13074,N_13075,N_13077,N_13079,N_13080,N_13081,N_13082,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13093,N_13094,N_13097,N_13099,N_13101,N_13102,N_13103,N_13105,N_13106,N_13107,N_13108,N_13109,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13125,N_13126,N_13127,N_13128,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13167,N_13168,N_13170,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13189,N_13190,N_13191,N_13192,N_13194,N_13195,N_13198,N_13200,N_13201,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13224,N_13225,N_13226,N_13228,N_13229,N_13230,N_13231,N_13234,N_13235,N_13236,N_13238,N_13239,N_13240,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13250,N_13251,N_13252,N_13254,N_13256,N_13258,N_13259,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13272,N_13276,N_13277,N_13278,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13290,N_13291,N_13292,N_13293,N_13294,N_13296,N_13297,N_13298,N_13299,N_13301,N_13302,N_13304,N_13305,N_13306,N_13307,N_13308,N_13310,N_13311,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13360,N_13363,N_13364,N_13365,N_13367,N_13368,N_13369,N_13371,N_13372,N_13373,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13387,N_13388,N_13389,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13400,N_13401,N_13402,N_13403,N_13405,N_13406,N_13407,N_13408,N_13410,N_13411,N_13413,N_13414,N_13416,N_13417,N_13419,N_13420,N_13421,N_13422,N_13423,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13435,N_13436,N_13437,N_13439,N_13440,N_13441,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13450,N_13454,N_13455,N_13456,N_13457,N_13458,N_13460,N_13462,N_13463,N_13464,N_13466,N_13467,N_13468,N_13469,N_13470,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13494,N_13495,N_13496,N_13497,N_13499,N_13501,N_13502,N_13503,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13514,N_13515,N_13516,N_13517,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13526,N_13528,N_13530,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13539,N_13540,N_13541,N_13544,N_13545,N_13546,N_13547,N_13549,N_13550,N_13551,N_13553,N_13555,N_13557,N_13558,N_13559,N_13560,N_13561,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13600,N_13601,N_13603,N_13604,N_13605,N_13607,N_13608,N_13609,N_13612,N_13613,N_13615,N_13616,N_13617,N_13618,N_13622,N_13623,N_13624,N_13626,N_13627,N_13628,N_13629,N_13630,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13639,N_13640,N_13641,N_13643,N_13645,N_13646,N_13647,N_13648,N_13649,N_13651,N_13652,N_13653,N_13654,N_13656,N_13657,N_13658,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13684,N_13685,N_13688,N_13689,N_13690,N_13692,N_13693,N_13694,N_13697,N_13698,N_13699,N_13700,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13724,N_13725,N_13726,N_13727,N_13729,N_13730,N_13731,N_13732,N_13733,N_13735,N_13736,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13754,N_13756,N_13758,N_13760,N_13761,N_13762,N_13763,N_13765,N_13766,N_13767,N_13769,N_13770,N_13771,N_13773,N_13774,N_13775,N_13776,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13793,N_13794,N_13797,N_13798,N_13802,N_13804,N_13805,N_13806,N_13807,N_13809,N_13811,N_13812,N_13814,N_13815,N_13816,N_13817,N_13818,N_13820,N_13821,N_13822,N_13823,N_13825,N_13826,N_13827,N_13828,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13840,N_13841,N_13843,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13854,N_13855,N_13857,N_13859,N_13860,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13874,N_13875,N_13876,N_13877,N_13879,N_13880,N_13881,N_13882,N_13884,N_13886,N_13887,N_13888,N_13891,N_13893,N_13894,N_13896,N_13897,N_13898,N_13900,N_13901,N_13902,N_13903,N_13904,N_13906,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13924,N_13925,N_13926,N_13928,N_13930,N_13931,N_13932,N_13933,N_13935,N_13936,N_13937,N_13938,N_13939,N_13942,N_13943,N_13944,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13955,N_13958,N_13959,N_13960,N_13961,N_13962,N_13964,N_13965,N_13966,N_13967,N_13969,N_13971,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13983,N_13984,N_13985,N_13988,N_13992,N_13993,N_13994,N_13996,N_13997,N_13998,N_14001,N_14002,N_14003,N_14004,N_14006,N_14007,N_14008,N_14010,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14022,N_14023,N_14024,N_14025,N_14028,N_14029,N_14030,N_14031,N_14032,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14061,N_14062,N_14064,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14076,N_14077,N_14078,N_14079,N_14081,N_14082,N_14083,N_14084,N_14085,N_14087,N_14089,N_14093,N_14095,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14105,N_14106,N_14108,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14119,N_14120,N_14121,N_14122,N_14123,N_14126,N_14127,N_14128,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14168,N_14171,N_14173,N_14174,N_14176,N_14177,N_14178,N_14179,N_14180,N_14182,N_14183,N_14184,N_14185,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14200,N_14201,N_14202,N_14204,N_14205,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14222,N_14223,N_14224,N_14225,N_14226,N_14228,N_14229,N_14230,N_14231,N_14234,N_14236,N_14238,N_14239,N_14240,N_14241,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14258,N_14259,N_14260,N_14261,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14302,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14316,N_14320,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14330,N_14334,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14343,N_14344,N_14345,N_14347,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14364,N_14366,N_14368,N_14370,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14383,N_14384,N_14385,N_14386,N_14388,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14398,N_14399,N_14400,N_14401,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14428,N_14429,N_14431,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14448,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14463,N_14464,N_14465,N_14466,N_14469,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14500,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14540,N_14541,N_14542,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14562,N_14563,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14578,N_14579,N_14580,N_14581,N_14583,N_14584,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14606,N_14607,N_14608,N_14610,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14656,N_14658,N_14659,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14668,N_14669,N_14670,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14681,N_14682,N_14683,N_14684,N_14685,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14714,N_14715,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14746,N_14748,N_14750,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14768,N_14769,N_14770,N_14771,N_14773,N_14775,N_14776,N_14777,N_14778,N_14779,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14788,N_14789,N_14790,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14817,N_14824,N_14826,N_14827,N_14828,N_14829,N_14830,N_14832,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14849,N_14851,N_14852,N_14854,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14864,N_14865,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14875,N_14876,N_14877,N_14879,N_14880,N_14882,N_14883,N_14884,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14899,N_14900,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14915,N_14916,N_14917,N_14920,N_14922,N_14923,N_14927,N_14928,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14940,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_61,In_1229);
and U1 (N_1,In_343,In_984);
and U2 (N_2,In_1366,In_852);
or U3 (N_3,In_938,In_176);
or U4 (N_4,In_1056,In_111);
nor U5 (N_5,In_1011,In_1419);
and U6 (N_6,In_225,In_1096);
or U7 (N_7,In_1160,In_1023);
and U8 (N_8,In_528,In_368);
nand U9 (N_9,In_1027,In_1061);
nor U10 (N_10,In_575,In_499);
xor U11 (N_11,In_1481,In_865);
xor U12 (N_12,In_1048,In_1000);
nor U13 (N_13,In_996,In_412);
xnor U14 (N_14,In_502,In_1070);
nor U15 (N_15,In_526,In_1051);
and U16 (N_16,In_681,In_604);
xnor U17 (N_17,In_1141,In_1112);
and U18 (N_18,In_71,In_1242);
xnor U19 (N_19,In_193,In_86);
and U20 (N_20,In_900,In_829);
nor U21 (N_21,In_1327,In_1068);
nor U22 (N_22,In_919,In_710);
and U23 (N_23,In_565,In_1081);
nand U24 (N_24,In_406,In_1474);
nand U25 (N_25,In_1405,In_1188);
xor U26 (N_26,In_123,In_701);
nor U27 (N_27,In_1363,In_339);
nor U28 (N_28,In_391,In_448);
nor U29 (N_29,In_1337,In_597);
nand U30 (N_30,In_1085,In_127);
or U31 (N_31,In_402,In_130);
nor U32 (N_32,In_779,In_312);
nand U33 (N_33,In_1269,In_1256);
or U34 (N_34,In_1468,In_52);
or U35 (N_35,In_188,In_138);
xor U36 (N_36,In_1288,In_767);
nor U37 (N_37,In_1454,In_1305);
xor U38 (N_38,In_1278,In_1470);
nand U39 (N_39,In_1120,In_1039);
xnor U40 (N_40,In_727,In_667);
xor U41 (N_41,In_758,In_1429);
or U42 (N_42,In_508,In_640);
nand U43 (N_43,In_847,In_1099);
xnor U44 (N_44,In_743,In_1187);
xor U45 (N_45,In_1064,In_781);
xor U46 (N_46,In_1456,In_103);
or U47 (N_47,In_398,In_706);
xnor U48 (N_48,In_432,In_8);
xnor U49 (N_49,In_1346,In_95);
xnor U50 (N_50,In_860,In_1371);
and U51 (N_51,In_1424,In_601);
and U52 (N_52,In_322,In_1493);
or U53 (N_53,In_1435,In_978);
nor U54 (N_54,In_821,In_1072);
or U55 (N_55,In_1417,In_458);
nor U56 (N_56,In_328,In_114);
and U57 (N_57,In_39,In_913);
nand U58 (N_58,In_1237,In_884);
nor U59 (N_59,In_660,In_538);
nand U60 (N_60,In_1486,In_1257);
or U61 (N_61,In_107,In_467);
nor U62 (N_62,In_636,In_119);
xor U63 (N_63,In_1028,In_1035);
nor U64 (N_64,In_255,In_1388);
nand U65 (N_65,In_126,In_461);
or U66 (N_66,In_995,In_1054);
nand U67 (N_67,In_1398,In_1220);
nor U68 (N_68,In_644,In_213);
xnor U69 (N_69,In_911,In_836);
and U70 (N_70,In_1149,In_778);
and U71 (N_71,In_456,In_13);
nand U72 (N_72,In_68,In_493);
and U73 (N_73,In_902,In_1375);
and U74 (N_74,In_963,In_1351);
nor U75 (N_75,In_650,In_1155);
nand U76 (N_76,In_1031,In_329);
and U77 (N_77,In_292,In_1377);
and U78 (N_78,In_480,In_285);
and U79 (N_79,In_626,In_1408);
or U80 (N_80,In_72,In_1128);
nor U81 (N_81,In_1362,In_845);
nand U82 (N_82,In_171,In_338);
or U83 (N_83,In_1394,In_905);
xor U84 (N_84,In_1249,In_1342);
nor U85 (N_85,In_484,In_278);
nor U86 (N_86,In_1244,In_1368);
xnor U87 (N_87,In_959,In_1040);
nand U88 (N_88,In_1207,In_998);
nand U89 (N_89,In_823,In_1029);
nor U90 (N_90,In_53,In_1421);
or U91 (N_91,In_3,In_359);
nand U92 (N_92,In_291,In_1194);
and U93 (N_93,In_179,In_896);
xor U94 (N_94,In_1320,In_868);
nand U95 (N_95,In_997,In_65);
nor U96 (N_96,In_449,In_788);
xnor U97 (N_97,In_986,In_629);
nand U98 (N_98,In_1492,In_124);
nand U99 (N_99,In_624,In_979);
and U100 (N_100,In_614,In_704);
and U101 (N_101,In_1147,In_300);
and U102 (N_102,In_909,In_337);
and U103 (N_103,In_1344,In_232);
nor U104 (N_104,In_642,In_268);
and U105 (N_105,In_4,In_699);
nand U106 (N_106,In_128,In_944);
or U107 (N_107,In_1222,In_1045);
nor U108 (N_108,In_417,In_739);
nor U109 (N_109,In_90,In_464);
nor U110 (N_110,In_1459,In_513);
nand U111 (N_111,In_286,In_748);
xnor U112 (N_112,In_655,In_1240);
xnor U113 (N_113,In_1125,In_587);
or U114 (N_114,In_1418,In_506);
nand U115 (N_115,In_1361,In_488);
and U116 (N_116,In_332,In_1004);
nand U117 (N_117,In_915,In_1267);
nor U118 (N_118,In_1176,In_732);
xnor U119 (N_119,In_738,In_664);
xnor U120 (N_120,In_1005,In_1428);
or U121 (N_121,In_1034,In_532);
nand U122 (N_122,In_1338,In_723);
and U123 (N_123,In_81,In_351);
and U124 (N_124,In_26,In_1271);
nor U125 (N_125,In_204,In_1432);
nor U126 (N_126,In_888,In_1233);
nor U127 (N_127,In_298,In_874);
nand U128 (N_128,In_1183,In_570);
and U129 (N_129,In_1313,In_440);
nand U130 (N_130,In_152,In_638);
xnor U131 (N_131,In_29,In_651);
or U132 (N_132,In_1379,In_828);
nor U133 (N_133,In_215,In_1392);
nand U134 (N_134,In_811,In_36);
or U135 (N_135,In_1019,In_1339);
nand U136 (N_136,In_290,In_192);
or U137 (N_137,In_381,In_364);
nand U138 (N_138,In_142,In_725);
nand U139 (N_139,In_798,In_1251);
nor U140 (N_140,In_573,In_542);
or U141 (N_141,In_91,In_610);
or U142 (N_142,In_830,In_1100);
nand U143 (N_143,In_594,In_46);
xnor U144 (N_144,In_964,In_1227);
nand U145 (N_145,In_953,In_853);
or U146 (N_146,In_1404,In_140);
nor U147 (N_147,In_856,In_691);
or U148 (N_148,In_410,In_507);
and U149 (N_149,In_304,In_1438);
nor U150 (N_150,In_267,In_1219);
or U151 (N_151,In_409,In_205);
xnor U152 (N_152,In_315,In_1234);
nand U153 (N_153,In_1014,In_1108);
nand U154 (N_154,In_447,In_1228);
or U155 (N_155,In_397,In_1300);
nand U156 (N_156,In_492,In_362);
xnor U157 (N_157,In_420,In_980);
nand U158 (N_158,In_1494,In_363);
or U159 (N_159,In_1445,In_1186);
nor U160 (N_160,In_721,In_209);
or U161 (N_161,In_280,In_987);
and U162 (N_162,In_1292,In_1103);
nor U163 (N_163,In_937,In_975);
xnor U164 (N_164,In_32,In_730);
and U165 (N_165,In_1043,In_731);
and U166 (N_166,In_317,In_797);
or U167 (N_167,In_117,In_372);
and U168 (N_168,In_314,In_607);
nand U169 (N_169,In_559,In_195);
and U170 (N_170,In_1197,In_620);
xnor U171 (N_171,In_952,In_189);
nor U172 (N_172,In_876,In_705);
nor U173 (N_173,In_139,In_84);
nor U174 (N_174,In_679,In_490);
nor U175 (N_175,In_1097,In_161);
or U176 (N_176,In_1347,In_1358);
nor U177 (N_177,In_104,In_1464);
nand U178 (N_178,In_1010,In_530);
nand U179 (N_179,In_170,In_234);
and U180 (N_180,In_541,In_1426);
nor U181 (N_181,In_1472,In_50);
nand U182 (N_182,In_603,In_407);
xnor U183 (N_183,In_524,In_23);
or U184 (N_184,In_791,In_360);
nand U185 (N_185,In_833,In_1441);
nor U186 (N_186,In_825,In_297);
or U187 (N_187,In_1461,In_951);
nor U188 (N_188,In_954,In_1403);
or U189 (N_189,In_672,In_1166);
nor U190 (N_190,In_1025,In_1198);
and U191 (N_191,In_1077,In_970);
or U192 (N_192,In_385,In_776);
xnor U193 (N_193,In_253,In_1480);
or U194 (N_194,In_912,In_948);
xnor U195 (N_195,In_934,In_1431);
nor U196 (N_196,In_678,In_1210);
nand U197 (N_197,In_231,In_415);
and U198 (N_198,In_454,In_137);
xnor U199 (N_199,In_1190,In_94);
nor U200 (N_200,In_931,In_848);
nor U201 (N_201,In_54,In_533);
xor U202 (N_202,In_635,In_1387);
xor U203 (N_203,In_1323,In_849);
and U204 (N_204,In_668,In_1469);
nand U205 (N_205,In_422,In_974);
and U206 (N_206,In_752,In_403);
xnor U207 (N_207,In_521,In_822);
and U208 (N_208,In_76,In_973);
nor U209 (N_209,In_1478,In_486);
or U210 (N_210,In_1032,In_74);
nand U211 (N_211,In_707,In_1400);
nor U212 (N_212,In_1317,In_843);
xnor U213 (N_213,In_1127,In_303);
nand U214 (N_214,In_875,In_387);
or U215 (N_215,In_914,In_375);
and U216 (N_216,In_321,In_237);
xnor U217 (N_217,In_211,In_308);
xnor U218 (N_218,In_181,In_643);
or U219 (N_219,In_1049,In_1255);
nor U220 (N_220,In_971,In_165);
xor U221 (N_221,In_718,In_1129);
xor U222 (N_222,In_1450,In_1236);
or U223 (N_223,In_516,In_51);
nor U224 (N_224,In_1243,In_1226);
or U225 (N_225,In_1266,In_946);
xor U226 (N_226,In_457,In_945);
nand U227 (N_227,In_450,In_1248);
nor U228 (N_228,In_613,In_1283);
or U229 (N_229,In_235,In_881);
and U230 (N_230,In_1307,In_77);
or U231 (N_231,In_983,In_851);
nand U232 (N_232,In_1,In_100);
nand U233 (N_233,In_595,In_56);
nor U234 (N_234,In_1277,In_720);
nand U235 (N_235,In_1433,In_306);
nand U236 (N_236,In_1448,In_10);
and U237 (N_237,In_1336,In_1425);
xnor U238 (N_238,In_413,In_1225);
and U239 (N_239,In_1066,In_1109);
nand U240 (N_240,In_481,In_968);
or U241 (N_241,In_641,In_1416);
xor U242 (N_242,In_1293,In_159);
and U243 (N_243,In_1084,In_862);
or U244 (N_244,In_742,In_1137);
nor U245 (N_245,In_1017,In_47);
xor U246 (N_246,In_148,In_14);
nand U247 (N_247,In_1439,In_112);
nor U248 (N_248,In_302,In_1488);
nand U249 (N_249,In_1178,In_977);
and U250 (N_250,In_248,In_769);
xnor U251 (N_251,In_229,In_196);
and U252 (N_252,In_878,In_0);
or U253 (N_253,In_1091,In_583);
or U254 (N_254,In_1465,In_110);
nand U255 (N_255,In_44,In_1089);
and U256 (N_256,In_872,In_1062);
nand U257 (N_257,In_1216,In_1374);
and U258 (N_258,In_150,In_358);
and U259 (N_259,In_677,In_272);
or U260 (N_260,In_344,In_514);
nor U261 (N_261,In_435,In_438);
and U262 (N_262,In_729,In_579);
xnor U263 (N_263,In_352,In_459);
nor U264 (N_264,In_645,In_1013);
and U265 (N_265,In_1087,In_1304);
nand U266 (N_266,In_961,In_1422);
nand U267 (N_267,In_346,In_652);
or U268 (N_268,In_156,In_1158);
xor U269 (N_269,In_763,In_1151);
xnor U270 (N_270,In_759,In_890);
xnor U271 (N_271,In_365,In_1086);
and U272 (N_272,In_616,In_1314);
or U273 (N_273,In_1383,In_442);
xnor U274 (N_274,In_325,In_745);
xor U275 (N_275,In_348,In_1442);
or U276 (N_276,In_1487,In_1261);
nor U277 (N_277,In_200,In_907);
or U278 (N_278,In_108,In_1075);
xnor U279 (N_279,In_82,In_261);
xnor U280 (N_280,In_675,In_1495);
or U281 (N_281,In_1270,In_460);
or U282 (N_282,In_1065,In_585);
nand U283 (N_283,In_79,In_904);
nand U284 (N_284,In_198,In_494);
xnor U285 (N_285,In_1399,In_177);
nand U286 (N_286,In_1407,In_772);
or U287 (N_287,In_728,In_969);
or U288 (N_288,In_1462,In_1202);
nor U289 (N_289,In_734,In_175);
xnor U290 (N_290,In_482,In_157);
or U291 (N_291,In_1209,In_1095);
nor U292 (N_292,In_544,In_1322);
nand U293 (N_293,In_1440,In_1106);
xnor U294 (N_294,In_1378,In_589);
xnor U295 (N_295,In_281,In_1059);
nor U296 (N_296,In_639,In_498);
and U297 (N_297,In_208,In_649);
and U298 (N_298,In_840,In_994);
nor U299 (N_299,In_1284,In_41);
nor U300 (N_300,In_578,In_1038);
and U301 (N_301,In_1258,In_174);
xor U302 (N_302,In_653,In_96);
xor U303 (N_303,In_1491,In_331);
nor U304 (N_304,In_1093,In_495);
nor U305 (N_305,In_894,In_816);
and U306 (N_306,In_503,In_279);
xnor U307 (N_307,In_527,In_12);
xor U308 (N_308,In_657,In_892);
nand U309 (N_309,In_433,In_1148);
or U310 (N_310,In_891,In_378);
nand U311 (N_311,In_569,In_1179);
or U312 (N_312,In_1069,In_665);
or U313 (N_313,In_1200,In_1175);
nand U314 (N_314,In_556,In_618);
nand U315 (N_315,In_453,In_1296);
or U316 (N_316,In_563,In_125);
and U317 (N_317,In_399,In_491);
xor U318 (N_318,In_269,In_698);
nand U319 (N_319,In_648,In_382);
nor U320 (N_320,In_859,In_1163);
xor U321 (N_321,In_501,In_1335);
or U322 (N_322,In_1185,In_1490);
and U323 (N_323,In_925,In_773);
nand U324 (N_324,In_414,In_1352);
and U325 (N_325,In_275,In_680);
nand U326 (N_326,In_584,In_88);
nand U327 (N_327,In_49,In_801);
nand U328 (N_328,In_592,In_832);
or U329 (N_329,In_887,In_11);
nand U330 (N_330,In_250,In_1246);
nor U331 (N_331,In_371,In_591);
and U332 (N_332,In_958,In_558);
nor U333 (N_333,In_478,In_416);
nor U334 (N_334,In_1451,In_560);
nand U335 (N_335,In_1309,In_855);
xor U336 (N_336,In_666,In_1180);
xnor U337 (N_337,In_850,In_245);
and U338 (N_338,In_430,In_1310);
or U339 (N_339,In_73,In_886);
xnor U340 (N_340,In_361,In_608);
nand U341 (N_341,In_1389,In_1218);
nand U342 (N_342,In_1250,In_120);
and U343 (N_343,In_804,In_345);
or U344 (N_344,In_550,In_1437);
nor U345 (N_345,In_101,In_927);
or U346 (N_346,In_1232,In_1355);
and U347 (N_347,In_153,In_1140);
nand U348 (N_348,In_87,In_1205);
and U349 (N_349,In_113,In_355);
xnor U350 (N_350,In_1098,In_1326);
xnor U351 (N_351,In_1396,In_571);
and U352 (N_352,In_1423,In_238);
nor U353 (N_353,In_247,In_1333);
nand U354 (N_354,In_1015,In_1489);
xor U355 (N_355,In_287,In_342);
xor U356 (N_356,In_19,In_222);
nor U357 (N_357,In_260,In_795);
and U358 (N_358,In_697,In_525);
xnor U359 (N_359,In_426,In_155);
nor U360 (N_360,In_1189,In_28);
or U361 (N_361,In_1156,In_1348);
xnor U362 (N_362,In_185,In_1321);
xor U363 (N_363,In_1130,In_988);
nor U364 (N_364,In_418,In_1033);
and U365 (N_365,In_168,In_939);
and U366 (N_366,In_755,In_370);
xor U367 (N_367,In_842,In_441);
and U368 (N_368,In_1238,In_324);
and U369 (N_369,In_1275,In_682);
or U370 (N_370,In_1057,In_813);
nor U371 (N_371,In_831,In_805);
xor U372 (N_372,In_1359,In_479);
nor U373 (N_373,In_863,In_580);
xnor U374 (N_374,In_452,In_1286);
and U375 (N_375,In_227,In_932);
nor U376 (N_376,In_374,In_992);
nor U377 (N_377,In_1146,In_146);
xor U378 (N_378,In_1074,In_1058);
nand U379 (N_379,In_340,In_1133);
nor U380 (N_380,In_1298,In_468);
nand U381 (N_381,In_1131,In_1050);
nor U382 (N_382,In_561,In_1341);
nand U383 (N_383,In_7,In_5);
and U384 (N_384,In_1410,In_1297);
xnor U385 (N_385,In_443,In_1088);
nor U386 (N_386,In_737,In_1123);
or U387 (N_387,In_803,In_239);
or U388 (N_388,In_1191,In_326);
nor U389 (N_389,In_588,In_700);
xnor U390 (N_390,In_1311,In_218);
and U391 (N_391,In_197,In_48);
and U392 (N_392,In_34,In_1026);
nor U393 (N_393,In_1079,In_1415);
nor U394 (N_394,In_145,In_309);
or U395 (N_395,In_955,In_1102);
xor U396 (N_396,In_765,In_709);
or U397 (N_397,In_899,In_754);
and U398 (N_398,In_1214,In_257);
xnor U399 (N_399,In_431,In_796);
or U400 (N_400,In_895,In_1107);
nor U401 (N_401,In_350,In_619);
and U402 (N_402,In_217,In_673);
xor U403 (N_403,In_80,In_1482);
or U404 (N_404,In_622,In_1245);
and U405 (N_405,In_1002,In_207);
nor U406 (N_406,In_1414,In_330);
or U407 (N_407,In_598,In_132);
or U408 (N_408,In_462,In_815);
and U409 (N_409,In_1150,In_568);
or U410 (N_410,In_202,In_1285);
xor U411 (N_411,In_879,In_473);
nand U412 (N_412,In_1262,In_711);
or U413 (N_413,In_252,In_985);
or U414 (N_414,In_131,In_392);
nor U415 (N_415,In_719,In_935);
or U416 (N_416,In_747,In_910);
or U417 (N_417,In_548,In_136);
nor U418 (N_418,In_1036,In_838);
nor U419 (N_419,In_31,In_857);
nand U420 (N_420,In_621,In_962);
and U421 (N_421,In_1308,In_1299);
nor U422 (N_422,In_522,In_802);
or U423 (N_423,In_45,In_357);
nand U424 (N_424,In_694,In_66);
or U425 (N_425,In_898,In_472);
xor U426 (N_426,In_485,In_611);
or U427 (N_427,In_824,In_266);
and U428 (N_428,In_576,In_1276);
nand U429 (N_429,In_670,In_947);
nor U430 (N_430,In_349,In_606);
nand U431 (N_431,In_518,In_1092);
or U432 (N_432,In_134,In_790);
nor U433 (N_433,In_510,In_158);
or U434 (N_434,In_1367,In_1372);
or U435 (N_435,In_477,In_24);
nand U436 (N_436,In_921,In_474);
nor U437 (N_437,In_817,In_662);
xor U438 (N_438,In_1124,In_893);
and U439 (N_439,In_722,In_249);
and U440 (N_440,In_1047,In_1090);
xor U441 (N_441,In_336,In_335);
nor U442 (N_442,In_265,In_808);
and U443 (N_443,In_323,In_1364);
and U444 (N_444,In_783,In_1302);
xor U445 (N_445,In_692,In_933);
and U446 (N_446,In_950,In_685);
and U447 (N_447,In_820,In_1473);
and U448 (N_448,In_633,In_178);
and U449 (N_449,In_436,In_121);
nor U450 (N_450,In_557,In_419);
nand U451 (N_451,In_751,In_1443);
nor U452 (N_452,In_889,In_993);
xor U453 (N_453,In_1485,In_22);
nand U454 (N_454,In_1263,In_1330);
xnor U455 (N_455,In_1199,In_1119);
and U456 (N_456,In_63,In_386);
nor U457 (N_457,In_630,In_703);
nor U458 (N_458,In_943,In_301);
or U459 (N_459,In_1152,In_105);
nand U460 (N_460,In_809,In_1390);
nand U461 (N_461,In_1252,In_184);
xnor U462 (N_462,In_172,In_182);
and U463 (N_463,In_839,In_552);
nand U464 (N_464,In_1386,In_540);
nand U465 (N_465,In_296,In_674);
xnor U466 (N_466,In_1496,In_30);
xnor U467 (N_467,In_547,In_870);
xnor U468 (N_468,In_744,In_259);
nor U469 (N_469,In_60,In_497);
nor U470 (N_470,In_1221,In_390);
and U471 (N_471,In_989,In_310);
and U472 (N_472,In_982,In_966);
nand U473 (N_473,In_885,In_1067);
or U474 (N_474,In_1325,In_487);
nand U475 (N_475,In_122,In_379);
xor U476 (N_476,In_1181,In_1007);
and U477 (N_477,In_1280,In_1174);
and U478 (N_478,In_930,In_276);
nor U479 (N_479,In_936,In_1212);
xnor U480 (N_480,In_318,In_1447);
nand U481 (N_481,In_354,In_1409);
nor U482 (N_482,In_186,In_1094);
xor U483 (N_483,In_1260,In_1016);
or U484 (N_484,In_1213,In_226);
or U485 (N_485,In_835,In_221);
nand U486 (N_486,In_313,In_1171);
or U487 (N_487,In_389,In_273);
or U488 (N_488,In_129,In_733);
xnor U489 (N_489,In_741,In_1060);
xnor U490 (N_490,In_299,In_717);
nor U491 (N_491,In_6,In_810);
or U492 (N_492,In_427,In_512);
and U493 (N_493,In_240,In_1020);
nand U494 (N_494,In_496,In_1273);
nor U495 (N_495,In_846,In_17);
xor U496 (N_496,In_1012,In_543);
nand U497 (N_497,In_320,In_531);
xor U498 (N_498,In_940,In_1476);
or U499 (N_499,In_1008,In_1172);
or U500 (N_500,In_70,In_1145);
and U501 (N_501,In_877,In_1170);
xnor U502 (N_502,In_1078,In_646);
or U503 (N_503,In_1498,In_37);
xnor U504 (N_504,In_423,In_564);
nor U505 (N_505,In_246,In_1165);
or U506 (N_506,In_827,In_401);
nor U507 (N_507,In_369,In_787);
or U508 (N_508,In_18,In_883);
and U509 (N_509,In_1101,In_289);
nor U510 (N_510,In_1201,In_256);
and U511 (N_511,In_58,In_469);
nor U512 (N_512,In_736,In_294);
and U513 (N_513,In_714,In_546);
or U514 (N_514,In_1042,In_444);
or U515 (N_515,In_1265,In_806);
nor U516 (N_516,In_434,In_917);
or U517 (N_517,In_1206,In_762);
nand U518 (N_518,In_1370,In_164);
nand U519 (N_519,In_251,In_991);
nand U520 (N_520,In_1453,In_1115);
xnor U521 (N_521,In_1455,In_702);
nor U522 (N_522,In_1239,In_819);
or U523 (N_523,In_380,In_1231);
xnor U524 (N_524,In_466,In_115);
nand U525 (N_525,In_782,In_1173);
or U526 (N_526,In_1161,In_768);
or U527 (N_527,In_1452,In_1458);
and U528 (N_528,In_149,In_689);
nor U529 (N_529,In_1471,In_393);
nor U530 (N_530,In_194,In_1446);
or U531 (N_531,In_596,In_577);
nand U532 (N_532,In_1009,In_1215);
or U533 (N_533,In_210,In_1082);
and U534 (N_534,In_567,In_928);
or U535 (N_535,In_429,In_637);
or U536 (N_536,In_224,In_428);
nor U537 (N_537,In_116,In_244);
or U538 (N_538,In_1162,In_715);
and U539 (N_539,In_228,In_534);
and U540 (N_540,In_284,In_135);
nand U541 (N_541,In_214,In_1457);
nor U542 (N_542,In_1143,In_180);
xor U543 (N_543,In_612,In_471);
and U544 (N_544,In_599,In_1055);
or U545 (N_545,In_421,In_212);
nand U546 (N_546,In_750,In_529);
xor U547 (N_547,In_1353,In_236);
nor U548 (N_548,In_1073,In_923);
nor U549 (N_549,In_1167,In_1272);
nor U550 (N_550,In_1349,In_437);
and U551 (N_551,In_305,In_271);
and U552 (N_552,In_404,In_967);
nand U553 (N_553,In_373,In_789);
or U554 (N_554,In_696,In_1329);
nand U555 (N_555,In_470,In_341);
nor U556 (N_556,In_411,In_1479);
and U557 (N_557,In_574,In_1463);
xor U558 (N_558,In_242,In_133);
xnor U559 (N_559,In_1105,In_27);
or U560 (N_560,In_1037,In_1195);
or U561 (N_561,In_42,In_1204);
and U562 (N_562,In_799,In_1328);
nor U563 (N_563,In_1434,In_523);
or U564 (N_564,In_1315,In_99);
or U565 (N_565,In_519,In_1306);
nand U566 (N_566,In_511,In_716);
nand U567 (N_567,In_647,In_794);
nor U568 (N_568,In_949,In_295);
xor U569 (N_569,In_1196,In_1113);
and U570 (N_570,In_555,In_483);
nor U571 (N_571,In_1076,In_1357);
nand U572 (N_572,In_687,In_377);
and U573 (N_573,In_187,In_1044);
nand U574 (N_574,In_858,In_1235);
xor U575 (N_575,In_141,In_683);
xnor U576 (N_576,In_1281,In_169);
xor U577 (N_577,In_190,In_627);
nand U578 (N_578,In_1324,In_764);
xor U579 (N_579,In_1318,In_770);
and U580 (N_580,In_871,In_85);
nor U581 (N_581,In_97,In_713);
nand U582 (N_582,In_760,In_1203);
nand U583 (N_583,In_600,In_143);
or U584 (N_584,In_1169,In_43);
xnor U585 (N_585,In_283,In_463);
nand U586 (N_586,In_632,In_981);
and U587 (N_587,In_1142,In_792);
nor U588 (N_588,In_1052,In_1153);
xnor U589 (N_589,In_241,In_21);
and U590 (N_590,In_1376,In_976);
nand U591 (N_591,In_1312,In_671);
xor U592 (N_592,In_445,In_771);
xor U593 (N_593,In_1154,In_656);
nor U594 (N_594,In_465,In_658);
and U595 (N_595,In_554,In_903);
or U596 (N_596,In_774,In_897);
nor U597 (N_597,In_118,In_535);
nor U598 (N_598,In_924,In_439);
nand U599 (N_599,In_793,In_311);
xnor U600 (N_600,In_258,In_366);
or U601 (N_601,In_16,In_1022);
nand U602 (N_602,In_1483,In_1182);
or U603 (N_603,In_1230,In_1006);
and U604 (N_604,In_356,In_775);
nand U605 (N_605,In_784,In_1126);
and U606 (N_606,In_777,In_686);
or U607 (N_607,In_1177,In_1294);
and U608 (N_608,In_307,In_1287);
xnor U609 (N_609,In_394,In_1030);
nor U610 (N_610,In_220,In_1334);
xor U611 (N_611,In_766,In_628);
nor U612 (N_612,In_749,In_882);
and U613 (N_613,In_1118,In_277);
nor U614 (N_614,In_586,In_1393);
or U615 (N_615,In_1289,In_35);
and U616 (N_616,In_1268,In_1373);
xor U617 (N_617,In_785,In_695);
nand U618 (N_618,In_92,In_1467);
nand U619 (N_619,In_475,In_1083);
nor U620 (N_620,In_965,In_33);
nor U621 (N_621,In_219,In_1411);
nor U622 (N_622,In_941,In_75);
nor U623 (N_623,In_353,In_384);
nor U624 (N_624,In_388,In_1134);
or U625 (N_625,In_1144,In_93);
xor U626 (N_626,In_1475,In_167);
or U627 (N_627,In_1224,In_1135);
and U628 (N_628,In_396,In_1382);
nand U629 (N_629,In_376,In_807);
xor U630 (N_630,In_1136,In_590);
xnor U631 (N_631,In_83,In_1259);
nand U632 (N_632,In_1279,In_999);
and U633 (N_633,In_263,In_800);
nand U634 (N_634,In_1018,In_262);
nand U635 (N_635,In_243,In_1241);
or U636 (N_636,In_1021,In_1164);
xor U637 (N_637,In_1122,In_254);
xnor U638 (N_638,In_451,In_1274);
nor U639 (N_639,In_203,In_408);
nand U640 (N_640,In_690,In_1071);
nor U641 (N_641,In_1168,In_106);
nor U642 (N_642,In_55,In_395);
xor U643 (N_643,In_282,In_582);
and U644 (N_644,In_1365,In_1121);
nor U645 (N_645,In_1484,In_867);
xnor U646 (N_646,In_593,In_724);
nor U647 (N_647,In_424,In_676);
and U648 (N_648,In_1412,In_1138);
xnor U649 (N_649,In_1436,In_89);
nand U650 (N_650,In_183,In_1444);
xor U651 (N_651,In_623,In_753);
and U652 (N_652,In_956,In_1449);
and U653 (N_653,In_509,In_160);
and U654 (N_654,In_1356,In_756);
or U655 (N_655,In_367,In_163);
nor U656 (N_656,In_1157,In_1295);
nor U657 (N_657,In_144,In_1117);
xnor U658 (N_658,In_918,In_1046);
nand U659 (N_659,In_1354,In_78);
nor U660 (N_660,In_1104,In_708);
nand U661 (N_661,In_274,In_230);
or U662 (N_662,In_1208,In_780);
nor U663 (N_663,In_1499,In_786);
xnor U664 (N_664,In_57,In_38);
and U665 (N_665,In_500,In_1413);
nand U666 (N_666,In_504,In_539);
or U667 (N_667,In_1497,In_1385);
nor U668 (N_668,In_562,In_1331);
xor U669 (N_669,In_69,In_1466);
and U670 (N_670,In_1381,In_960);
and U671 (N_671,In_669,In_2);
and U672 (N_672,In_873,In_553);
xnor U673 (N_673,In_319,In_1110);
xor U674 (N_674,In_489,In_551);
xor U675 (N_675,In_1063,In_40);
or U676 (N_676,In_1319,In_537);
and U677 (N_677,In_1003,In_631);
xor U678 (N_678,In_1401,In_1116);
nand U679 (N_679,In_663,In_929);
nor U680 (N_680,In_844,In_216);
nor U681 (N_681,In_1420,In_549);
nand U682 (N_682,In_659,In_837);
xor U683 (N_683,In_625,In_834);
nand U684 (N_684,In_1041,In_1395);
xnor U685 (N_685,In_383,In_288);
nor U686 (N_686,In_615,In_405);
nor U687 (N_687,In_520,In_1114);
and U688 (N_688,In_901,In_264);
and U689 (N_689,In_293,In_926);
or U690 (N_690,In_166,In_206);
xnor U691 (N_691,In_581,In_1159);
xor U692 (N_692,In_201,In_233);
or U693 (N_693,In_757,In_1430);
or U694 (N_694,In_1406,In_1192);
and U695 (N_695,In_1264,In_654);
nor U696 (N_696,In_866,In_62);
nand U697 (N_697,In_446,In_1111);
or U698 (N_698,In_64,In_1053);
and U699 (N_699,In_942,In_861);
nand U700 (N_700,In_572,In_223);
xor U701 (N_701,In_1282,In_814);
xor U702 (N_702,In_400,In_1340);
and U703 (N_703,In_712,In_605);
xnor U704 (N_704,In_515,In_1303);
and U705 (N_705,In_688,In_1024);
and U706 (N_706,In_864,In_191);
nand U707 (N_707,In_347,In_455);
nor U708 (N_708,In_922,In_726);
and U709 (N_709,In_162,In_818);
nand U710 (N_710,In_1343,In_1254);
nor U711 (N_711,In_536,In_1460);
nor U712 (N_712,In_1350,In_1384);
nor U713 (N_713,In_102,In_1345);
nand U714 (N_714,In_20,In_1402);
or U715 (N_715,In_1427,In_9);
and U716 (N_716,In_517,In_1253);
and U717 (N_717,In_609,In_1080);
xnor U718 (N_718,In_1380,In_1391);
nand U719 (N_719,In_746,In_1223);
xnor U720 (N_720,In_916,In_920);
and U721 (N_721,In_1001,In_1184);
nand U722 (N_722,In_761,In_1139);
nor U723 (N_723,In_505,In_740);
or U724 (N_724,In_476,In_333);
nor U725 (N_725,In_826,In_1477);
xnor U726 (N_726,In_869,In_1290);
and U727 (N_727,In_59,In_1193);
or U728 (N_728,In_98,In_735);
or U729 (N_729,In_908,In_602);
nor U730 (N_730,In_1132,In_854);
and U731 (N_731,In_957,In_1247);
and U732 (N_732,In_1301,In_1397);
xnor U733 (N_733,In_67,In_327);
nor U734 (N_734,In_880,In_812);
nand U735 (N_735,In_1217,In_15);
or U736 (N_736,In_990,In_634);
or U737 (N_737,In_154,In_1332);
nand U738 (N_738,In_566,In_661);
xor U739 (N_739,In_25,In_906);
xnor U740 (N_740,In_109,In_425);
nor U741 (N_741,In_334,In_147);
or U742 (N_742,In_617,In_684);
nand U743 (N_743,In_316,In_1360);
xnor U744 (N_744,In_1291,In_151);
or U745 (N_745,In_972,In_1316);
nor U746 (N_746,In_1369,In_545);
nor U747 (N_747,In_173,In_1211);
xnor U748 (N_748,In_841,In_199);
xor U749 (N_749,In_693,In_270);
nor U750 (N_750,In_337,In_186);
nor U751 (N_751,In_793,In_919);
nor U752 (N_752,In_579,In_1318);
and U753 (N_753,In_1249,In_885);
and U754 (N_754,In_523,In_406);
and U755 (N_755,In_613,In_650);
or U756 (N_756,In_1427,In_52);
nand U757 (N_757,In_1467,In_866);
xor U758 (N_758,In_747,In_441);
and U759 (N_759,In_140,In_79);
and U760 (N_760,In_893,In_407);
nor U761 (N_761,In_694,In_316);
nand U762 (N_762,In_1090,In_1113);
nand U763 (N_763,In_1367,In_79);
nor U764 (N_764,In_432,In_27);
or U765 (N_765,In_523,In_1452);
nand U766 (N_766,In_62,In_221);
and U767 (N_767,In_1188,In_1105);
and U768 (N_768,In_736,In_699);
xnor U769 (N_769,In_90,In_750);
and U770 (N_770,In_51,In_986);
nand U771 (N_771,In_37,In_131);
and U772 (N_772,In_1385,In_503);
nor U773 (N_773,In_1273,In_63);
nor U774 (N_774,In_1437,In_665);
nand U775 (N_775,In_943,In_987);
or U776 (N_776,In_6,In_597);
nor U777 (N_777,In_697,In_1377);
xor U778 (N_778,In_84,In_602);
nand U779 (N_779,In_649,In_588);
nor U780 (N_780,In_1083,In_3);
nand U781 (N_781,In_268,In_539);
and U782 (N_782,In_519,In_505);
nand U783 (N_783,In_1006,In_23);
nor U784 (N_784,In_1474,In_571);
nand U785 (N_785,In_640,In_1190);
nand U786 (N_786,In_848,In_144);
nand U787 (N_787,In_657,In_885);
nand U788 (N_788,In_1485,In_1001);
xnor U789 (N_789,In_1498,In_832);
nor U790 (N_790,In_1016,In_1445);
or U791 (N_791,In_233,In_227);
nor U792 (N_792,In_989,In_859);
xor U793 (N_793,In_103,In_1177);
or U794 (N_794,In_559,In_140);
xor U795 (N_795,In_645,In_1229);
nor U796 (N_796,In_585,In_1332);
xor U797 (N_797,In_41,In_268);
nand U798 (N_798,In_1360,In_809);
nor U799 (N_799,In_593,In_693);
or U800 (N_800,In_0,In_1330);
nand U801 (N_801,In_161,In_408);
and U802 (N_802,In_14,In_1456);
and U803 (N_803,In_436,In_1016);
or U804 (N_804,In_912,In_848);
and U805 (N_805,In_409,In_508);
nand U806 (N_806,In_1300,In_242);
and U807 (N_807,In_326,In_241);
nand U808 (N_808,In_1036,In_592);
or U809 (N_809,In_1309,In_337);
or U810 (N_810,In_734,In_651);
xnor U811 (N_811,In_317,In_1246);
xnor U812 (N_812,In_287,In_670);
and U813 (N_813,In_1437,In_1025);
or U814 (N_814,In_772,In_1355);
nor U815 (N_815,In_119,In_560);
nor U816 (N_816,In_1016,In_1171);
nor U817 (N_817,In_851,In_225);
and U818 (N_818,In_185,In_49);
and U819 (N_819,In_236,In_57);
and U820 (N_820,In_913,In_362);
or U821 (N_821,In_290,In_1356);
or U822 (N_822,In_782,In_680);
or U823 (N_823,In_1244,In_272);
or U824 (N_824,In_12,In_1182);
or U825 (N_825,In_571,In_799);
nand U826 (N_826,In_92,In_413);
nor U827 (N_827,In_1188,In_1497);
nand U828 (N_828,In_1444,In_680);
nand U829 (N_829,In_1184,In_655);
xnor U830 (N_830,In_701,In_288);
and U831 (N_831,In_284,In_574);
and U832 (N_832,In_1283,In_1126);
nand U833 (N_833,In_1423,In_346);
xnor U834 (N_834,In_941,In_1058);
nand U835 (N_835,In_1030,In_753);
and U836 (N_836,In_1015,In_1026);
nor U837 (N_837,In_1417,In_1036);
or U838 (N_838,In_771,In_160);
nand U839 (N_839,In_536,In_664);
or U840 (N_840,In_49,In_994);
xor U841 (N_841,In_297,In_333);
xor U842 (N_842,In_276,In_1094);
and U843 (N_843,In_57,In_49);
nand U844 (N_844,In_355,In_1466);
xnor U845 (N_845,In_971,In_204);
or U846 (N_846,In_905,In_315);
and U847 (N_847,In_1115,In_1021);
or U848 (N_848,In_814,In_617);
or U849 (N_849,In_732,In_462);
and U850 (N_850,In_151,In_1008);
xor U851 (N_851,In_102,In_227);
nand U852 (N_852,In_1156,In_728);
and U853 (N_853,In_648,In_951);
and U854 (N_854,In_927,In_1203);
and U855 (N_855,In_1279,In_1213);
xnor U856 (N_856,In_558,In_752);
nor U857 (N_857,In_1076,In_253);
nor U858 (N_858,In_918,In_1055);
xor U859 (N_859,In_128,In_485);
nand U860 (N_860,In_597,In_897);
and U861 (N_861,In_1260,In_546);
nand U862 (N_862,In_1324,In_94);
nor U863 (N_863,In_920,In_822);
nand U864 (N_864,In_93,In_1485);
nor U865 (N_865,In_1241,In_768);
or U866 (N_866,In_826,In_23);
nand U867 (N_867,In_628,In_334);
nand U868 (N_868,In_1337,In_948);
nor U869 (N_869,In_559,In_1041);
and U870 (N_870,In_1373,In_236);
nand U871 (N_871,In_229,In_684);
nor U872 (N_872,In_682,In_1263);
and U873 (N_873,In_665,In_726);
or U874 (N_874,In_911,In_592);
xor U875 (N_875,In_1376,In_327);
and U876 (N_876,In_1053,In_434);
nor U877 (N_877,In_899,In_473);
and U878 (N_878,In_1033,In_696);
and U879 (N_879,In_341,In_1317);
nand U880 (N_880,In_526,In_1368);
or U881 (N_881,In_1432,In_988);
nor U882 (N_882,In_1251,In_245);
nand U883 (N_883,In_198,In_712);
and U884 (N_884,In_424,In_753);
and U885 (N_885,In_1102,In_1351);
nand U886 (N_886,In_695,In_349);
nor U887 (N_887,In_1140,In_637);
nor U888 (N_888,In_195,In_523);
xnor U889 (N_889,In_1470,In_1017);
nor U890 (N_890,In_634,In_81);
xnor U891 (N_891,In_187,In_991);
or U892 (N_892,In_19,In_975);
xnor U893 (N_893,In_268,In_1301);
and U894 (N_894,In_1173,In_1254);
nor U895 (N_895,In_193,In_1250);
xnor U896 (N_896,In_200,In_1045);
and U897 (N_897,In_614,In_140);
or U898 (N_898,In_679,In_905);
xnor U899 (N_899,In_1250,In_279);
nand U900 (N_900,In_1461,In_608);
nor U901 (N_901,In_906,In_518);
and U902 (N_902,In_17,In_512);
xor U903 (N_903,In_721,In_1397);
and U904 (N_904,In_213,In_116);
nor U905 (N_905,In_388,In_859);
nand U906 (N_906,In_475,In_1230);
or U907 (N_907,In_36,In_810);
nand U908 (N_908,In_435,In_285);
nand U909 (N_909,In_1144,In_137);
or U910 (N_910,In_90,In_1327);
xnor U911 (N_911,In_1345,In_1490);
xor U912 (N_912,In_829,In_1169);
xor U913 (N_913,In_899,In_428);
or U914 (N_914,In_1122,In_133);
or U915 (N_915,In_48,In_154);
or U916 (N_916,In_324,In_1352);
and U917 (N_917,In_1408,In_354);
nor U918 (N_918,In_1250,In_134);
or U919 (N_919,In_30,In_172);
and U920 (N_920,In_581,In_752);
xor U921 (N_921,In_229,In_877);
xnor U922 (N_922,In_1360,In_690);
and U923 (N_923,In_1267,In_1492);
nand U924 (N_924,In_291,In_443);
nor U925 (N_925,In_817,In_1327);
or U926 (N_926,In_1452,In_816);
or U927 (N_927,In_1046,In_705);
xor U928 (N_928,In_1376,In_853);
and U929 (N_929,In_776,In_1062);
and U930 (N_930,In_1409,In_196);
and U931 (N_931,In_650,In_506);
nor U932 (N_932,In_979,In_607);
nor U933 (N_933,In_1056,In_259);
and U934 (N_934,In_664,In_1393);
nand U935 (N_935,In_1135,In_1383);
xnor U936 (N_936,In_926,In_34);
and U937 (N_937,In_258,In_195);
nor U938 (N_938,In_110,In_1357);
nor U939 (N_939,In_652,In_1363);
and U940 (N_940,In_49,In_209);
nor U941 (N_941,In_129,In_346);
nand U942 (N_942,In_1068,In_408);
or U943 (N_943,In_646,In_722);
and U944 (N_944,In_391,In_539);
or U945 (N_945,In_1473,In_468);
nor U946 (N_946,In_1462,In_79);
nor U947 (N_947,In_291,In_372);
xor U948 (N_948,In_1035,In_619);
nor U949 (N_949,In_601,In_1495);
or U950 (N_950,In_553,In_453);
or U951 (N_951,In_1370,In_997);
and U952 (N_952,In_478,In_155);
nor U953 (N_953,In_923,In_423);
xnor U954 (N_954,In_1310,In_1126);
xor U955 (N_955,In_1363,In_1061);
nand U956 (N_956,In_197,In_382);
xnor U957 (N_957,In_1041,In_1446);
or U958 (N_958,In_1036,In_531);
nand U959 (N_959,In_195,In_370);
or U960 (N_960,In_285,In_701);
nor U961 (N_961,In_1235,In_999);
nand U962 (N_962,In_891,In_658);
or U963 (N_963,In_955,In_53);
xnor U964 (N_964,In_975,In_1026);
nand U965 (N_965,In_1420,In_1446);
and U966 (N_966,In_564,In_200);
and U967 (N_967,In_225,In_971);
and U968 (N_968,In_643,In_794);
nor U969 (N_969,In_1474,In_1362);
nor U970 (N_970,In_1000,In_323);
nand U971 (N_971,In_723,In_145);
nor U972 (N_972,In_440,In_750);
nand U973 (N_973,In_1103,In_1138);
or U974 (N_974,In_1437,In_782);
nor U975 (N_975,In_108,In_198);
nand U976 (N_976,In_630,In_942);
nor U977 (N_977,In_1413,In_1143);
nor U978 (N_978,In_112,In_315);
or U979 (N_979,In_813,In_51);
nand U980 (N_980,In_712,In_290);
nor U981 (N_981,In_846,In_1150);
and U982 (N_982,In_286,In_272);
nand U983 (N_983,In_909,In_283);
nor U984 (N_984,In_128,In_908);
and U985 (N_985,In_1046,In_879);
nor U986 (N_986,In_160,In_494);
and U987 (N_987,In_229,In_174);
and U988 (N_988,In_143,In_1368);
and U989 (N_989,In_254,In_308);
xor U990 (N_990,In_697,In_987);
or U991 (N_991,In_545,In_1237);
nand U992 (N_992,In_855,In_1039);
or U993 (N_993,In_1160,In_1219);
nor U994 (N_994,In_1401,In_913);
and U995 (N_995,In_950,In_1188);
and U996 (N_996,In_488,In_572);
and U997 (N_997,In_1448,In_343);
nor U998 (N_998,In_535,In_1377);
and U999 (N_999,In_750,In_50);
nand U1000 (N_1000,In_315,In_1271);
xnor U1001 (N_1001,In_1140,In_485);
or U1002 (N_1002,In_1437,In_781);
nor U1003 (N_1003,In_1357,In_549);
nor U1004 (N_1004,In_1232,In_1007);
nor U1005 (N_1005,In_908,In_992);
and U1006 (N_1006,In_1393,In_997);
and U1007 (N_1007,In_713,In_611);
nor U1008 (N_1008,In_824,In_1215);
nand U1009 (N_1009,In_437,In_971);
nand U1010 (N_1010,In_144,In_526);
or U1011 (N_1011,In_163,In_545);
nand U1012 (N_1012,In_132,In_817);
nand U1013 (N_1013,In_1042,In_486);
or U1014 (N_1014,In_303,In_798);
nor U1015 (N_1015,In_1146,In_401);
and U1016 (N_1016,In_150,In_1022);
or U1017 (N_1017,In_224,In_83);
nor U1018 (N_1018,In_1327,In_94);
or U1019 (N_1019,In_266,In_504);
or U1020 (N_1020,In_500,In_318);
or U1021 (N_1021,In_1411,In_732);
or U1022 (N_1022,In_791,In_1229);
and U1023 (N_1023,In_772,In_79);
and U1024 (N_1024,In_35,In_451);
nor U1025 (N_1025,In_516,In_1033);
or U1026 (N_1026,In_190,In_669);
or U1027 (N_1027,In_206,In_313);
nand U1028 (N_1028,In_69,In_149);
and U1029 (N_1029,In_326,In_1113);
xnor U1030 (N_1030,In_1009,In_1100);
and U1031 (N_1031,In_1127,In_1418);
nand U1032 (N_1032,In_257,In_1224);
nor U1033 (N_1033,In_946,In_606);
and U1034 (N_1034,In_1408,In_143);
and U1035 (N_1035,In_41,In_971);
nand U1036 (N_1036,In_1195,In_1440);
and U1037 (N_1037,In_311,In_551);
nor U1038 (N_1038,In_1137,In_406);
nor U1039 (N_1039,In_1477,In_125);
xnor U1040 (N_1040,In_929,In_626);
or U1041 (N_1041,In_809,In_633);
nand U1042 (N_1042,In_372,In_1136);
or U1043 (N_1043,In_316,In_131);
nand U1044 (N_1044,In_1425,In_738);
and U1045 (N_1045,In_888,In_1158);
xor U1046 (N_1046,In_1043,In_1069);
and U1047 (N_1047,In_598,In_0);
or U1048 (N_1048,In_529,In_773);
or U1049 (N_1049,In_1178,In_493);
nand U1050 (N_1050,In_548,In_739);
or U1051 (N_1051,In_16,In_1363);
and U1052 (N_1052,In_922,In_1169);
or U1053 (N_1053,In_1077,In_456);
nor U1054 (N_1054,In_1468,In_1345);
xnor U1055 (N_1055,In_667,In_1334);
xnor U1056 (N_1056,In_1158,In_1277);
xor U1057 (N_1057,In_1174,In_831);
nand U1058 (N_1058,In_611,In_551);
nor U1059 (N_1059,In_839,In_596);
nor U1060 (N_1060,In_1348,In_514);
and U1061 (N_1061,In_501,In_752);
or U1062 (N_1062,In_816,In_1398);
nand U1063 (N_1063,In_278,In_1392);
xnor U1064 (N_1064,In_720,In_674);
and U1065 (N_1065,In_1419,In_342);
nor U1066 (N_1066,In_542,In_434);
or U1067 (N_1067,In_75,In_118);
nor U1068 (N_1068,In_106,In_1218);
nand U1069 (N_1069,In_894,In_1342);
and U1070 (N_1070,In_667,In_639);
or U1071 (N_1071,In_1060,In_615);
or U1072 (N_1072,In_399,In_790);
nand U1073 (N_1073,In_1336,In_92);
xor U1074 (N_1074,In_594,In_829);
and U1075 (N_1075,In_160,In_1490);
and U1076 (N_1076,In_443,In_841);
xnor U1077 (N_1077,In_412,In_1153);
xor U1078 (N_1078,In_397,In_456);
nand U1079 (N_1079,In_502,In_1235);
nor U1080 (N_1080,In_1064,In_1190);
and U1081 (N_1081,In_887,In_294);
and U1082 (N_1082,In_686,In_1000);
and U1083 (N_1083,In_278,In_68);
nand U1084 (N_1084,In_1439,In_554);
nor U1085 (N_1085,In_1238,In_302);
nor U1086 (N_1086,In_662,In_1443);
nor U1087 (N_1087,In_55,In_799);
nand U1088 (N_1088,In_1172,In_680);
or U1089 (N_1089,In_632,In_1238);
or U1090 (N_1090,In_240,In_537);
nor U1091 (N_1091,In_605,In_1427);
or U1092 (N_1092,In_452,In_1455);
xnor U1093 (N_1093,In_1149,In_334);
or U1094 (N_1094,In_176,In_933);
or U1095 (N_1095,In_107,In_1301);
or U1096 (N_1096,In_502,In_1394);
or U1097 (N_1097,In_1147,In_972);
xor U1098 (N_1098,In_511,In_1412);
nand U1099 (N_1099,In_911,In_636);
nor U1100 (N_1100,In_860,In_276);
and U1101 (N_1101,In_709,In_639);
and U1102 (N_1102,In_795,In_1185);
nand U1103 (N_1103,In_531,In_470);
xor U1104 (N_1104,In_189,In_611);
xnor U1105 (N_1105,In_796,In_1072);
and U1106 (N_1106,In_913,In_571);
xnor U1107 (N_1107,In_195,In_602);
and U1108 (N_1108,In_51,In_837);
and U1109 (N_1109,In_1259,In_153);
nor U1110 (N_1110,In_993,In_1104);
nor U1111 (N_1111,In_1130,In_1415);
nand U1112 (N_1112,In_820,In_1209);
or U1113 (N_1113,In_336,In_1172);
nand U1114 (N_1114,In_1332,In_183);
nor U1115 (N_1115,In_249,In_1211);
nor U1116 (N_1116,In_76,In_511);
nand U1117 (N_1117,In_69,In_295);
and U1118 (N_1118,In_201,In_1010);
or U1119 (N_1119,In_478,In_1084);
or U1120 (N_1120,In_778,In_1026);
nand U1121 (N_1121,In_344,In_629);
xnor U1122 (N_1122,In_1034,In_40);
nand U1123 (N_1123,In_160,In_561);
and U1124 (N_1124,In_66,In_1275);
or U1125 (N_1125,In_550,In_1216);
nand U1126 (N_1126,In_55,In_121);
or U1127 (N_1127,In_377,In_1323);
xnor U1128 (N_1128,In_1091,In_703);
nand U1129 (N_1129,In_776,In_20);
and U1130 (N_1130,In_1366,In_720);
and U1131 (N_1131,In_1439,In_985);
xnor U1132 (N_1132,In_1491,In_1115);
and U1133 (N_1133,In_1491,In_613);
or U1134 (N_1134,In_828,In_192);
and U1135 (N_1135,In_1182,In_94);
nand U1136 (N_1136,In_931,In_1082);
or U1137 (N_1137,In_963,In_429);
xnor U1138 (N_1138,In_381,In_1329);
or U1139 (N_1139,In_82,In_1007);
nor U1140 (N_1140,In_1273,In_332);
or U1141 (N_1141,In_1498,In_601);
nor U1142 (N_1142,In_1019,In_463);
xor U1143 (N_1143,In_105,In_1361);
nor U1144 (N_1144,In_1289,In_847);
or U1145 (N_1145,In_1431,In_132);
or U1146 (N_1146,In_473,In_715);
or U1147 (N_1147,In_734,In_768);
and U1148 (N_1148,In_700,In_923);
xnor U1149 (N_1149,In_790,In_158);
nand U1150 (N_1150,In_687,In_128);
and U1151 (N_1151,In_794,In_509);
or U1152 (N_1152,In_1230,In_1198);
and U1153 (N_1153,In_810,In_368);
or U1154 (N_1154,In_1267,In_676);
nor U1155 (N_1155,In_802,In_58);
and U1156 (N_1156,In_1127,In_698);
nand U1157 (N_1157,In_314,In_372);
xor U1158 (N_1158,In_1396,In_1171);
or U1159 (N_1159,In_1364,In_218);
nand U1160 (N_1160,In_949,In_271);
or U1161 (N_1161,In_1267,In_943);
and U1162 (N_1162,In_907,In_1373);
xnor U1163 (N_1163,In_767,In_1293);
and U1164 (N_1164,In_726,In_620);
xnor U1165 (N_1165,In_1347,In_615);
xnor U1166 (N_1166,In_1170,In_1338);
and U1167 (N_1167,In_247,In_69);
and U1168 (N_1168,In_969,In_1078);
xnor U1169 (N_1169,In_1217,In_1078);
and U1170 (N_1170,In_890,In_73);
or U1171 (N_1171,In_810,In_1373);
and U1172 (N_1172,In_1036,In_646);
nand U1173 (N_1173,In_716,In_442);
or U1174 (N_1174,In_685,In_237);
or U1175 (N_1175,In_1310,In_145);
and U1176 (N_1176,In_917,In_808);
xor U1177 (N_1177,In_992,In_1239);
or U1178 (N_1178,In_1067,In_124);
or U1179 (N_1179,In_135,In_1373);
or U1180 (N_1180,In_440,In_446);
xor U1181 (N_1181,In_253,In_1288);
and U1182 (N_1182,In_847,In_988);
xor U1183 (N_1183,In_285,In_244);
or U1184 (N_1184,In_1261,In_639);
xnor U1185 (N_1185,In_100,In_1063);
xor U1186 (N_1186,In_329,In_514);
nand U1187 (N_1187,In_1234,In_1294);
or U1188 (N_1188,In_1236,In_1484);
nor U1189 (N_1189,In_1097,In_1208);
nor U1190 (N_1190,In_1202,In_881);
or U1191 (N_1191,In_33,In_1107);
and U1192 (N_1192,In_125,In_1214);
and U1193 (N_1193,In_312,In_761);
or U1194 (N_1194,In_541,In_909);
nor U1195 (N_1195,In_953,In_158);
and U1196 (N_1196,In_1490,In_1151);
nand U1197 (N_1197,In_797,In_343);
nor U1198 (N_1198,In_1356,In_936);
xor U1199 (N_1199,In_795,In_548);
nand U1200 (N_1200,In_116,In_668);
and U1201 (N_1201,In_421,In_140);
xor U1202 (N_1202,In_432,In_1144);
or U1203 (N_1203,In_279,In_1058);
xnor U1204 (N_1204,In_1275,In_1466);
nand U1205 (N_1205,In_1278,In_232);
xnor U1206 (N_1206,In_759,In_558);
nor U1207 (N_1207,In_1020,In_812);
and U1208 (N_1208,In_1131,In_32);
nor U1209 (N_1209,In_137,In_611);
xor U1210 (N_1210,In_550,In_456);
xor U1211 (N_1211,In_438,In_212);
and U1212 (N_1212,In_1279,In_36);
and U1213 (N_1213,In_996,In_722);
xnor U1214 (N_1214,In_696,In_1114);
nor U1215 (N_1215,In_1134,In_327);
nor U1216 (N_1216,In_285,In_1182);
or U1217 (N_1217,In_1382,In_409);
nor U1218 (N_1218,In_1043,In_555);
nand U1219 (N_1219,In_898,In_1016);
and U1220 (N_1220,In_549,In_1406);
nor U1221 (N_1221,In_887,In_1302);
xor U1222 (N_1222,In_1277,In_971);
or U1223 (N_1223,In_1355,In_1264);
and U1224 (N_1224,In_224,In_221);
xnor U1225 (N_1225,In_540,In_626);
nor U1226 (N_1226,In_1491,In_95);
xnor U1227 (N_1227,In_971,In_487);
nand U1228 (N_1228,In_371,In_112);
nand U1229 (N_1229,In_1221,In_139);
or U1230 (N_1230,In_531,In_1226);
nor U1231 (N_1231,In_853,In_566);
and U1232 (N_1232,In_1073,In_171);
xor U1233 (N_1233,In_821,In_382);
or U1234 (N_1234,In_645,In_1280);
nand U1235 (N_1235,In_1052,In_926);
nand U1236 (N_1236,In_404,In_301);
and U1237 (N_1237,In_391,In_1186);
nand U1238 (N_1238,In_1208,In_1419);
nor U1239 (N_1239,In_551,In_293);
or U1240 (N_1240,In_464,In_1398);
xnor U1241 (N_1241,In_499,In_100);
nor U1242 (N_1242,In_1103,In_1493);
nor U1243 (N_1243,In_1362,In_1022);
or U1244 (N_1244,In_363,In_5);
nor U1245 (N_1245,In_142,In_553);
nor U1246 (N_1246,In_446,In_913);
nor U1247 (N_1247,In_356,In_1416);
and U1248 (N_1248,In_667,In_464);
nor U1249 (N_1249,In_887,In_1429);
and U1250 (N_1250,In_419,In_1244);
xnor U1251 (N_1251,In_514,In_190);
xor U1252 (N_1252,In_1382,In_1434);
or U1253 (N_1253,In_118,In_1450);
xor U1254 (N_1254,In_1190,In_643);
xnor U1255 (N_1255,In_1011,In_998);
xor U1256 (N_1256,In_580,In_489);
xor U1257 (N_1257,In_687,In_65);
or U1258 (N_1258,In_846,In_161);
nand U1259 (N_1259,In_1466,In_262);
and U1260 (N_1260,In_1071,In_1178);
nor U1261 (N_1261,In_452,In_523);
or U1262 (N_1262,In_958,In_1245);
nand U1263 (N_1263,In_9,In_427);
and U1264 (N_1264,In_1237,In_1441);
or U1265 (N_1265,In_667,In_1290);
xor U1266 (N_1266,In_792,In_853);
xor U1267 (N_1267,In_1202,In_12);
or U1268 (N_1268,In_962,In_1497);
or U1269 (N_1269,In_473,In_381);
nand U1270 (N_1270,In_542,In_523);
nand U1271 (N_1271,In_1351,In_106);
and U1272 (N_1272,In_1326,In_710);
and U1273 (N_1273,In_1215,In_263);
xnor U1274 (N_1274,In_1095,In_1199);
xor U1275 (N_1275,In_761,In_604);
xnor U1276 (N_1276,In_833,In_23);
and U1277 (N_1277,In_288,In_1498);
and U1278 (N_1278,In_696,In_1336);
and U1279 (N_1279,In_1470,In_574);
xor U1280 (N_1280,In_585,In_828);
or U1281 (N_1281,In_438,In_1233);
and U1282 (N_1282,In_1113,In_1190);
and U1283 (N_1283,In_1159,In_755);
and U1284 (N_1284,In_302,In_1060);
and U1285 (N_1285,In_44,In_152);
nand U1286 (N_1286,In_140,In_1444);
xnor U1287 (N_1287,In_562,In_1453);
xnor U1288 (N_1288,In_1171,In_65);
or U1289 (N_1289,In_14,In_877);
nand U1290 (N_1290,In_112,In_1469);
and U1291 (N_1291,In_943,In_1045);
or U1292 (N_1292,In_809,In_289);
xnor U1293 (N_1293,In_1036,In_1411);
and U1294 (N_1294,In_80,In_302);
and U1295 (N_1295,In_1465,In_474);
xor U1296 (N_1296,In_837,In_1079);
xor U1297 (N_1297,In_344,In_371);
and U1298 (N_1298,In_182,In_1255);
nand U1299 (N_1299,In_1048,In_303);
xnor U1300 (N_1300,In_930,In_1271);
and U1301 (N_1301,In_1460,In_1337);
nand U1302 (N_1302,In_601,In_596);
or U1303 (N_1303,In_814,In_1006);
nor U1304 (N_1304,In_140,In_921);
nor U1305 (N_1305,In_845,In_1401);
and U1306 (N_1306,In_868,In_1277);
xor U1307 (N_1307,In_932,In_154);
xnor U1308 (N_1308,In_686,In_928);
xnor U1309 (N_1309,In_845,In_476);
nand U1310 (N_1310,In_1082,In_1442);
nor U1311 (N_1311,In_689,In_1388);
nand U1312 (N_1312,In_975,In_299);
nor U1313 (N_1313,In_1018,In_1494);
xor U1314 (N_1314,In_1409,In_1357);
xnor U1315 (N_1315,In_1073,In_886);
nor U1316 (N_1316,In_779,In_675);
and U1317 (N_1317,In_777,In_1142);
nand U1318 (N_1318,In_349,In_387);
or U1319 (N_1319,In_1424,In_472);
nor U1320 (N_1320,In_1112,In_735);
or U1321 (N_1321,In_833,In_1088);
and U1322 (N_1322,In_576,In_893);
nor U1323 (N_1323,In_1468,In_1040);
or U1324 (N_1324,In_1251,In_1449);
or U1325 (N_1325,In_930,In_325);
nor U1326 (N_1326,In_1489,In_647);
nor U1327 (N_1327,In_1446,In_1215);
xnor U1328 (N_1328,In_959,In_550);
nor U1329 (N_1329,In_257,In_951);
nand U1330 (N_1330,In_130,In_374);
and U1331 (N_1331,In_722,In_448);
and U1332 (N_1332,In_1494,In_1372);
or U1333 (N_1333,In_126,In_718);
nor U1334 (N_1334,In_1046,In_1031);
xor U1335 (N_1335,In_793,In_1430);
nor U1336 (N_1336,In_625,In_984);
or U1337 (N_1337,In_1080,In_430);
nor U1338 (N_1338,In_691,In_1164);
and U1339 (N_1339,In_7,In_1280);
nand U1340 (N_1340,In_384,In_112);
nand U1341 (N_1341,In_976,In_66);
nor U1342 (N_1342,In_517,In_208);
nor U1343 (N_1343,In_720,In_203);
nand U1344 (N_1344,In_850,In_726);
nor U1345 (N_1345,In_64,In_916);
or U1346 (N_1346,In_1344,In_355);
and U1347 (N_1347,In_685,In_980);
xnor U1348 (N_1348,In_236,In_879);
nor U1349 (N_1349,In_10,In_410);
or U1350 (N_1350,In_1230,In_1407);
nor U1351 (N_1351,In_146,In_964);
and U1352 (N_1352,In_1052,In_1393);
xnor U1353 (N_1353,In_201,In_272);
nor U1354 (N_1354,In_1197,In_773);
xnor U1355 (N_1355,In_834,In_1322);
and U1356 (N_1356,In_157,In_523);
and U1357 (N_1357,In_708,In_1049);
and U1358 (N_1358,In_1236,In_14);
nand U1359 (N_1359,In_1193,In_886);
xor U1360 (N_1360,In_899,In_1412);
xnor U1361 (N_1361,In_1300,In_456);
and U1362 (N_1362,In_623,In_1355);
or U1363 (N_1363,In_1235,In_1444);
nand U1364 (N_1364,In_1466,In_641);
xnor U1365 (N_1365,In_1049,In_403);
nand U1366 (N_1366,In_60,In_1389);
or U1367 (N_1367,In_365,In_1025);
and U1368 (N_1368,In_187,In_1224);
nand U1369 (N_1369,In_154,In_689);
or U1370 (N_1370,In_528,In_1217);
and U1371 (N_1371,In_1425,In_564);
nand U1372 (N_1372,In_835,In_239);
and U1373 (N_1373,In_1386,In_929);
xor U1374 (N_1374,In_651,In_1350);
xor U1375 (N_1375,In_1477,In_63);
and U1376 (N_1376,In_143,In_1410);
nand U1377 (N_1377,In_873,In_37);
xor U1378 (N_1378,In_917,In_318);
nor U1379 (N_1379,In_1167,In_1361);
xor U1380 (N_1380,In_1402,In_1396);
and U1381 (N_1381,In_112,In_901);
xnor U1382 (N_1382,In_1418,In_915);
nand U1383 (N_1383,In_981,In_32);
nand U1384 (N_1384,In_183,In_1337);
and U1385 (N_1385,In_645,In_60);
or U1386 (N_1386,In_774,In_34);
and U1387 (N_1387,In_830,In_1110);
nor U1388 (N_1388,In_1358,In_771);
xor U1389 (N_1389,In_1030,In_223);
nor U1390 (N_1390,In_1102,In_1189);
or U1391 (N_1391,In_171,In_596);
nand U1392 (N_1392,In_380,In_239);
xnor U1393 (N_1393,In_1150,In_348);
nor U1394 (N_1394,In_143,In_64);
nand U1395 (N_1395,In_778,In_995);
nor U1396 (N_1396,In_391,In_1054);
and U1397 (N_1397,In_0,In_1404);
or U1398 (N_1398,In_127,In_1112);
nor U1399 (N_1399,In_446,In_1238);
nor U1400 (N_1400,In_275,In_73);
and U1401 (N_1401,In_334,In_489);
nand U1402 (N_1402,In_208,In_609);
and U1403 (N_1403,In_1387,In_26);
nor U1404 (N_1404,In_76,In_314);
xnor U1405 (N_1405,In_350,In_537);
or U1406 (N_1406,In_1361,In_969);
or U1407 (N_1407,In_231,In_1059);
xnor U1408 (N_1408,In_1308,In_1159);
or U1409 (N_1409,In_1482,In_1400);
or U1410 (N_1410,In_780,In_1273);
nor U1411 (N_1411,In_157,In_145);
nor U1412 (N_1412,In_127,In_998);
nor U1413 (N_1413,In_281,In_1340);
nand U1414 (N_1414,In_636,In_1116);
and U1415 (N_1415,In_1237,In_620);
or U1416 (N_1416,In_1239,In_18);
nor U1417 (N_1417,In_48,In_1209);
nor U1418 (N_1418,In_611,In_394);
or U1419 (N_1419,In_1477,In_664);
and U1420 (N_1420,In_40,In_1474);
and U1421 (N_1421,In_1203,In_424);
and U1422 (N_1422,In_113,In_1484);
or U1423 (N_1423,In_1374,In_60);
xor U1424 (N_1424,In_680,In_1009);
nand U1425 (N_1425,In_90,In_1396);
and U1426 (N_1426,In_447,In_1330);
and U1427 (N_1427,In_911,In_176);
xor U1428 (N_1428,In_962,In_1360);
xor U1429 (N_1429,In_1311,In_607);
xor U1430 (N_1430,In_742,In_1143);
and U1431 (N_1431,In_1096,In_893);
xnor U1432 (N_1432,In_402,In_580);
or U1433 (N_1433,In_1226,In_303);
or U1434 (N_1434,In_716,In_1003);
or U1435 (N_1435,In_987,In_692);
nor U1436 (N_1436,In_1329,In_636);
and U1437 (N_1437,In_0,In_726);
xnor U1438 (N_1438,In_324,In_1130);
xor U1439 (N_1439,In_1144,In_1457);
or U1440 (N_1440,In_698,In_976);
nand U1441 (N_1441,In_330,In_1069);
nor U1442 (N_1442,In_947,In_1393);
or U1443 (N_1443,In_1124,In_1015);
nor U1444 (N_1444,In_320,In_1134);
nor U1445 (N_1445,In_1024,In_1097);
xnor U1446 (N_1446,In_1121,In_785);
nand U1447 (N_1447,In_1168,In_662);
and U1448 (N_1448,In_1365,In_503);
nor U1449 (N_1449,In_1212,In_257);
or U1450 (N_1450,In_639,In_443);
nand U1451 (N_1451,In_1459,In_835);
nand U1452 (N_1452,In_186,In_1346);
nand U1453 (N_1453,In_716,In_1031);
and U1454 (N_1454,In_354,In_1244);
nand U1455 (N_1455,In_252,In_1289);
nand U1456 (N_1456,In_1447,In_1271);
nor U1457 (N_1457,In_394,In_837);
or U1458 (N_1458,In_413,In_1187);
or U1459 (N_1459,In_92,In_549);
xnor U1460 (N_1460,In_325,In_1457);
nand U1461 (N_1461,In_745,In_1317);
nand U1462 (N_1462,In_1271,In_990);
nor U1463 (N_1463,In_1421,In_628);
nor U1464 (N_1464,In_431,In_320);
and U1465 (N_1465,In_52,In_106);
xor U1466 (N_1466,In_1366,In_969);
nor U1467 (N_1467,In_207,In_1070);
xor U1468 (N_1468,In_1295,In_836);
nor U1469 (N_1469,In_252,In_13);
or U1470 (N_1470,In_301,In_1420);
xor U1471 (N_1471,In_609,In_28);
nand U1472 (N_1472,In_216,In_1447);
nor U1473 (N_1473,In_1039,In_222);
nand U1474 (N_1474,In_189,In_503);
or U1475 (N_1475,In_644,In_146);
nor U1476 (N_1476,In_1273,In_1439);
or U1477 (N_1477,In_556,In_690);
nand U1478 (N_1478,In_91,In_194);
or U1479 (N_1479,In_1231,In_21);
xor U1480 (N_1480,In_1311,In_275);
and U1481 (N_1481,In_895,In_65);
nor U1482 (N_1482,In_469,In_672);
or U1483 (N_1483,In_326,In_1263);
and U1484 (N_1484,In_437,In_1247);
and U1485 (N_1485,In_1239,In_1264);
xnor U1486 (N_1486,In_1126,In_499);
xnor U1487 (N_1487,In_118,In_1329);
xor U1488 (N_1488,In_556,In_1303);
or U1489 (N_1489,In_294,In_477);
nor U1490 (N_1490,In_802,In_533);
or U1491 (N_1491,In_834,In_612);
xor U1492 (N_1492,In_400,In_1245);
or U1493 (N_1493,In_1319,In_98);
and U1494 (N_1494,In_1297,In_411);
nor U1495 (N_1495,In_286,In_64);
nor U1496 (N_1496,In_814,In_811);
and U1497 (N_1497,In_665,In_735);
and U1498 (N_1498,In_45,In_679);
or U1499 (N_1499,In_939,In_1437);
nand U1500 (N_1500,In_719,In_767);
nand U1501 (N_1501,In_584,In_1100);
xnor U1502 (N_1502,In_1277,In_670);
nand U1503 (N_1503,In_166,In_1213);
and U1504 (N_1504,In_384,In_331);
or U1505 (N_1505,In_602,In_330);
xnor U1506 (N_1506,In_347,In_1292);
xor U1507 (N_1507,In_823,In_1168);
nor U1508 (N_1508,In_937,In_840);
xnor U1509 (N_1509,In_1439,In_698);
or U1510 (N_1510,In_634,In_1249);
xor U1511 (N_1511,In_356,In_729);
nand U1512 (N_1512,In_1157,In_37);
nor U1513 (N_1513,In_927,In_1270);
nand U1514 (N_1514,In_1462,In_989);
nor U1515 (N_1515,In_1331,In_690);
and U1516 (N_1516,In_364,In_1247);
xnor U1517 (N_1517,In_829,In_690);
xnor U1518 (N_1518,In_1212,In_593);
nand U1519 (N_1519,In_182,In_559);
nor U1520 (N_1520,In_1363,In_68);
nand U1521 (N_1521,In_1304,In_805);
nand U1522 (N_1522,In_205,In_655);
nor U1523 (N_1523,In_300,In_978);
nor U1524 (N_1524,In_100,In_791);
nor U1525 (N_1525,In_1019,In_564);
nor U1526 (N_1526,In_574,In_872);
and U1527 (N_1527,In_19,In_1466);
nand U1528 (N_1528,In_785,In_175);
nor U1529 (N_1529,In_1313,In_1124);
nor U1530 (N_1530,In_978,In_997);
nor U1531 (N_1531,In_476,In_219);
nand U1532 (N_1532,In_794,In_274);
or U1533 (N_1533,In_377,In_1368);
or U1534 (N_1534,In_433,In_1481);
or U1535 (N_1535,In_482,In_798);
and U1536 (N_1536,In_375,In_626);
xor U1537 (N_1537,In_312,In_7);
or U1538 (N_1538,In_524,In_400);
nor U1539 (N_1539,In_534,In_1344);
or U1540 (N_1540,In_769,In_132);
and U1541 (N_1541,In_145,In_279);
or U1542 (N_1542,In_1081,In_1494);
nand U1543 (N_1543,In_1261,In_121);
nor U1544 (N_1544,In_498,In_1416);
nor U1545 (N_1545,In_355,In_232);
nand U1546 (N_1546,In_201,In_717);
and U1547 (N_1547,In_592,In_976);
xnor U1548 (N_1548,In_678,In_1188);
and U1549 (N_1549,In_603,In_944);
nor U1550 (N_1550,In_285,In_221);
xnor U1551 (N_1551,In_628,In_78);
nor U1552 (N_1552,In_145,In_1044);
or U1553 (N_1553,In_654,In_1255);
and U1554 (N_1554,In_944,In_921);
and U1555 (N_1555,In_1140,In_963);
nand U1556 (N_1556,In_128,In_782);
nor U1557 (N_1557,In_527,In_229);
xnor U1558 (N_1558,In_1245,In_1125);
nor U1559 (N_1559,In_1059,In_455);
nor U1560 (N_1560,In_278,In_770);
nor U1561 (N_1561,In_657,In_950);
or U1562 (N_1562,In_671,In_197);
nand U1563 (N_1563,In_1344,In_48);
nand U1564 (N_1564,In_394,In_557);
nor U1565 (N_1565,In_815,In_468);
or U1566 (N_1566,In_1115,In_1405);
xor U1567 (N_1567,In_209,In_1062);
nor U1568 (N_1568,In_206,In_157);
nor U1569 (N_1569,In_1342,In_846);
nor U1570 (N_1570,In_1226,In_895);
nor U1571 (N_1571,In_1121,In_720);
nand U1572 (N_1572,In_390,In_1101);
nor U1573 (N_1573,In_1231,In_476);
nor U1574 (N_1574,In_1031,In_256);
nor U1575 (N_1575,In_1087,In_289);
or U1576 (N_1576,In_253,In_322);
and U1577 (N_1577,In_774,In_334);
nor U1578 (N_1578,In_140,In_624);
xnor U1579 (N_1579,In_1138,In_422);
or U1580 (N_1580,In_65,In_51);
xor U1581 (N_1581,In_1142,In_102);
or U1582 (N_1582,In_1247,In_1388);
nand U1583 (N_1583,In_57,In_1331);
nor U1584 (N_1584,In_22,In_485);
and U1585 (N_1585,In_1442,In_153);
or U1586 (N_1586,In_358,In_1114);
and U1587 (N_1587,In_40,In_876);
and U1588 (N_1588,In_393,In_569);
nor U1589 (N_1589,In_179,In_1430);
and U1590 (N_1590,In_1264,In_1307);
or U1591 (N_1591,In_941,In_78);
and U1592 (N_1592,In_972,In_941);
and U1593 (N_1593,In_1298,In_313);
xnor U1594 (N_1594,In_495,In_331);
nor U1595 (N_1595,In_341,In_1419);
nand U1596 (N_1596,In_1301,In_332);
and U1597 (N_1597,In_1224,In_981);
nand U1598 (N_1598,In_685,In_1474);
or U1599 (N_1599,In_902,In_456);
xor U1600 (N_1600,In_596,In_1369);
or U1601 (N_1601,In_1444,In_456);
nor U1602 (N_1602,In_780,In_462);
or U1603 (N_1603,In_1481,In_612);
or U1604 (N_1604,In_119,In_342);
xnor U1605 (N_1605,In_1243,In_1194);
or U1606 (N_1606,In_1443,In_1025);
xor U1607 (N_1607,In_77,In_909);
and U1608 (N_1608,In_359,In_427);
xor U1609 (N_1609,In_982,In_1347);
nand U1610 (N_1610,In_726,In_1384);
and U1611 (N_1611,In_1152,In_611);
xor U1612 (N_1612,In_713,In_95);
xnor U1613 (N_1613,In_825,In_897);
or U1614 (N_1614,In_1038,In_1122);
nand U1615 (N_1615,In_1421,In_944);
nor U1616 (N_1616,In_862,In_534);
and U1617 (N_1617,In_506,In_949);
xnor U1618 (N_1618,In_287,In_1340);
xor U1619 (N_1619,In_660,In_120);
nor U1620 (N_1620,In_224,In_796);
or U1621 (N_1621,In_885,In_789);
nor U1622 (N_1622,In_811,In_242);
nand U1623 (N_1623,In_69,In_134);
nor U1624 (N_1624,In_141,In_482);
nor U1625 (N_1625,In_916,In_677);
nand U1626 (N_1626,In_240,In_402);
nand U1627 (N_1627,In_762,In_1396);
nand U1628 (N_1628,In_840,In_145);
xnor U1629 (N_1629,In_1115,In_904);
or U1630 (N_1630,In_254,In_452);
and U1631 (N_1631,In_359,In_97);
xnor U1632 (N_1632,In_240,In_1286);
nor U1633 (N_1633,In_405,In_723);
nand U1634 (N_1634,In_710,In_489);
nor U1635 (N_1635,In_1138,In_378);
nor U1636 (N_1636,In_1083,In_955);
xor U1637 (N_1637,In_361,In_615);
nor U1638 (N_1638,In_422,In_10);
or U1639 (N_1639,In_425,In_1429);
and U1640 (N_1640,In_803,In_1373);
or U1641 (N_1641,In_208,In_1415);
nand U1642 (N_1642,In_174,In_383);
nand U1643 (N_1643,In_956,In_230);
and U1644 (N_1644,In_169,In_332);
xnor U1645 (N_1645,In_970,In_1029);
nand U1646 (N_1646,In_291,In_949);
or U1647 (N_1647,In_415,In_669);
xnor U1648 (N_1648,In_338,In_819);
and U1649 (N_1649,In_96,In_200);
or U1650 (N_1650,In_470,In_589);
and U1651 (N_1651,In_96,In_1173);
or U1652 (N_1652,In_443,In_440);
nor U1653 (N_1653,In_1302,In_1213);
nor U1654 (N_1654,In_792,In_599);
and U1655 (N_1655,In_1079,In_274);
xor U1656 (N_1656,In_468,In_146);
and U1657 (N_1657,In_876,In_82);
xor U1658 (N_1658,In_19,In_9);
and U1659 (N_1659,In_34,In_975);
nand U1660 (N_1660,In_766,In_448);
and U1661 (N_1661,In_161,In_950);
xnor U1662 (N_1662,In_437,In_467);
or U1663 (N_1663,In_1084,In_330);
and U1664 (N_1664,In_925,In_199);
xor U1665 (N_1665,In_1430,In_925);
or U1666 (N_1666,In_584,In_1432);
or U1667 (N_1667,In_331,In_71);
nor U1668 (N_1668,In_1407,In_1186);
or U1669 (N_1669,In_919,In_1461);
xor U1670 (N_1670,In_653,In_469);
nand U1671 (N_1671,In_920,In_664);
or U1672 (N_1672,In_454,In_303);
or U1673 (N_1673,In_1213,In_292);
and U1674 (N_1674,In_609,In_421);
and U1675 (N_1675,In_1267,In_722);
nor U1676 (N_1676,In_888,In_32);
nand U1677 (N_1677,In_1180,In_369);
and U1678 (N_1678,In_763,In_949);
or U1679 (N_1679,In_983,In_1335);
nand U1680 (N_1680,In_492,In_1156);
xnor U1681 (N_1681,In_123,In_1007);
nand U1682 (N_1682,In_891,In_10);
and U1683 (N_1683,In_516,In_500);
nand U1684 (N_1684,In_1129,In_985);
or U1685 (N_1685,In_223,In_613);
or U1686 (N_1686,In_1480,In_520);
nand U1687 (N_1687,In_1048,In_448);
or U1688 (N_1688,In_1424,In_47);
or U1689 (N_1689,In_259,In_637);
nor U1690 (N_1690,In_521,In_13);
and U1691 (N_1691,In_1260,In_804);
and U1692 (N_1692,In_973,In_860);
xor U1693 (N_1693,In_1265,In_1277);
xnor U1694 (N_1694,In_1394,In_1438);
nand U1695 (N_1695,In_1340,In_780);
nor U1696 (N_1696,In_953,In_1168);
and U1697 (N_1697,In_9,In_1010);
nand U1698 (N_1698,In_686,In_1233);
nor U1699 (N_1699,In_320,In_877);
nand U1700 (N_1700,In_318,In_894);
nor U1701 (N_1701,In_578,In_400);
or U1702 (N_1702,In_570,In_433);
or U1703 (N_1703,In_522,In_683);
nand U1704 (N_1704,In_997,In_1135);
and U1705 (N_1705,In_167,In_1234);
nand U1706 (N_1706,In_760,In_721);
xnor U1707 (N_1707,In_463,In_553);
xnor U1708 (N_1708,In_1258,In_122);
and U1709 (N_1709,In_482,In_264);
and U1710 (N_1710,In_250,In_734);
xnor U1711 (N_1711,In_1241,In_1323);
xnor U1712 (N_1712,In_1312,In_626);
nor U1713 (N_1713,In_383,In_714);
nand U1714 (N_1714,In_1493,In_663);
xor U1715 (N_1715,In_1344,In_807);
nand U1716 (N_1716,In_1473,In_1499);
and U1717 (N_1717,In_27,In_532);
and U1718 (N_1718,In_1055,In_1000);
or U1719 (N_1719,In_5,In_927);
or U1720 (N_1720,In_257,In_461);
xor U1721 (N_1721,In_880,In_667);
or U1722 (N_1722,In_1227,In_602);
nand U1723 (N_1723,In_1273,In_347);
nor U1724 (N_1724,In_996,In_1001);
or U1725 (N_1725,In_929,In_388);
nand U1726 (N_1726,In_338,In_1440);
nand U1727 (N_1727,In_1417,In_1327);
nand U1728 (N_1728,In_408,In_4);
or U1729 (N_1729,In_221,In_1407);
xor U1730 (N_1730,In_774,In_537);
or U1731 (N_1731,In_72,In_759);
and U1732 (N_1732,In_758,In_603);
nand U1733 (N_1733,In_978,In_1074);
nor U1734 (N_1734,In_549,In_863);
and U1735 (N_1735,In_376,In_962);
nand U1736 (N_1736,In_1304,In_146);
nor U1737 (N_1737,In_1163,In_904);
and U1738 (N_1738,In_1351,In_135);
and U1739 (N_1739,In_141,In_316);
or U1740 (N_1740,In_1111,In_994);
xor U1741 (N_1741,In_974,In_1098);
nor U1742 (N_1742,In_1390,In_286);
nor U1743 (N_1743,In_881,In_1144);
xor U1744 (N_1744,In_494,In_815);
xor U1745 (N_1745,In_1073,In_110);
nand U1746 (N_1746,In_255,In_608);
nor U1747 (N_1747,In_747,In_528);
xnor U1748 (N_1748,In_1262,In_726);
xor U1749 (N_1749,In_644,In_1011);
and U1750 (N_1750,In_622,In_1087);
and U1751 (N_1751,In_1370,In_152);
and U1752 (N_1752,In_52,In_1099);
nor U1753 (N_1753,In_353,In_348);
nand U1754 (N_1754,In_1278,In_35);
and U1755 (N_1755,In_301,In_585);
nor U1756 (N_1756,In_574,In_134);
or U1757 (N_1757,In_539,In_297);
nor U1758 (N_1758,In_327,In_147);
nand U1759 (N_1759,In_856,In_264);
and U1760 (N_1760,In_740,In_1135);
nand U1761 (N_1761,In_1369,In_798);
nand U1762 (N_1762,In_854,In_449);
xnor U1763 (N_1763,In_339,In_611);
nand U1764 (N_1764,In_167,In_1221);
nand U1765 (N_1765,In_1098,In_351);
or U1766 (N_1766,In_1295,In_572);
nor U1767 (N_1767,In_141,In_843);
xnor U1768 (N_1768,In_132,In_1234);
nand U1769 (N_1769,In_445,In_883);
and U1770 (N_1770,In_505,In_899);
and U1771 (N_1771,In_288,In_1411);
and U1772 (N_1772,In_650,In_1323);
nor U1773 (N_1773,In_1191,In_718);
or U1774 (N_1774,In_418,In_1430);
xor U1775 (N_1775,In_1196,In_810);
xor U1776 (N_1776,In_1421,In_1086);
or U1777 (N_1777,In_216,In_1080);
nand U1778 (N_1778,In_321,In_1381);
nand U1779 (N_1779,In_1239,In_213);
and U1780 (N_1780,In_275,In_338);
nand U1781 (N_1781,In_937,In_90);
and U1782 (N_1782,In_1212,In_847);
nor U1783 (N_1783,In_955,In_1124);
nor U1784 (N_1784,In_202,In_1038);
or U1785 (N_1785,In_1083,In_871);
nand U1786 (N_1786,In_1167,In_1232);
nand U1787 (N_1787,In_708,In_1266);
nor U1788 (N_1788,In_418,In_1227);
xnor U1789 (N_1789,In_638,In_1265);
and U1790 (N_1790,In_1238,In_1014);
nand U1791 (N_1791,In_21,In_1293);
xor U1792 (N_1792,In_1038,In_432);
and U1793 (N_1793,In_1415,In_861);
nor U1794 (N_1794,In_1011,In_155);
nand U1795 (N_1795,In_260,In_430);
nand U1796 (N_1796,In_1331,In_1252);
xnor U1797 (N_1797,In_463,In_1048);
or U1798 (N_1798,In_835,In_1028);
nand U1799 (N_1799,In_1132,In_98);
xnor U1800 (N_1800,In_769,In_642);
nand U1801 (N_1801,In_1015,In_535);
xnor U1802 (N_1802,In_59,In_487);
or U1803 (N_1803,In_121,In_891);
and U1804 (N_1804,In_1114,In_815);
and U1805 (N_1805,In_454,In_1384);
xor U1806 (N_1806,In_1334,In_112);
nand U1807 (N_1807,In_286,In_1163);
xnor U1808 (N_1808,In_323,In_883);
or U1809 (N_1809,In_980,In_1487);
or U1810 (N_1810,In_1396,In_814);
xor U1811 (N_1811,In_1291,In_842);
xnor U1812 (N_1812,In_121,In_954);
xnor U1813 (N_1813,In_2,In_1052);
xnor U1814 (N_1814,In_1176,In_485);
and U1815 (N_1815,In_1014,In_221);
and U1816 (N_1816,In_791,In_44);
or U1817 (N_1817,In_1073,In_180);
xnor U1818 (N_1818,In_886,In_632);
xor U1819 (N_1819,In_320,In_100);
or U1820 (N_1820,In_592,In_1119);
nor U1821 (N_1821,In_616,In_1017);
or U1822 (N_1822,In_44,In_1488);
nor U1823 (N_1823,In_542,In_707);
xor U1824 (N_1824,In_208,In_1021);
and U1825 (N_1825,In_1102,In_488);
nand U1826 (N_1826,In_101,In_1061);
nor U1827 (N_1827,In_1328,In_1352);
and U1828 (N_1828,In_964,In_9);
nand U1829 (N_1829,In_858,In_1426);
xnor U1830 (N_1830,In_919,In_85);
and U1831 (N_1831,In_1081,In_764);
xnor U1832 (N_1832,In_646,In_680);
or U1833 (N_1833,In_1444,In_1340);
xnor U1834 (N_1834,In_154,In_877);
nand U1835 (N_1835,In_591,In_1064);
and U1836 (N_1836,In_578,In_1030);
nand U1837 (N_1837,In_29,In_907);
or U1838 (N_1838,In_916,In_1268);
or U1839 (N_1839,In_381,In_851);
xnor U1840 (N_1840,In_794,In_139);
nand U1841 (N_1841,In_698,In_1265);
and U1842 (N_1842,In_414,In_1313);
or U1843 (N_1843,In_934,In_1363);
nand U1844 (N_1844,In_1392,In_128);
or U1845 (N_1845,In_536,In_687);
or U1846 (N_1846,In_1431,In_1128);
and U1847 (N_1847,In_501,In_1251);
nor U1848 (N_1848,In_892,In_203);
nand U1849 (N_1849,In_167,In_470);
or U1850 (N_1850,In_1046,In_1305);
xor U1851 (N_1851,In_265,In_432);
or U1852 (N_1852,In_303,In_1181);
and U1853 (N_1853,In_263,In_1393);
or U1854 (N_1854,In_1328,In_671);
or U1855 (N_1855,In_556,In_601);
nor U1856 (N_1856,In_207,In_578);
and U1857 (N_1857,In_95,In_1025);
and U1858 (N_1858,In_798,In_1392);
and U1859 (N_1859,In_482,In_715);
or U1860 (N_1860,In_39,In_650);
xnor U1861 (N_1861,In_101,In_478);
xnor U1862 (N_1862,In_1202,In_213);
xnor U1863 (N_1863,In_32,In_1043);
and U1864 (N_1864,In_704,In_8);
nand U1865 (N_1865,In_781,In_3);
nand U1866 (N_1866,In_377,In_1031);
and U1867 (N_1867,In_1152,In_481);
xor U1868 (N_1868,In_1374,In_1398);
xor U1869 (N_1869,In_833,In_1079);
or U1870 (N_1870,In_297,In_1102);
nor U1871 (N_1871,In_1423,In_244);
and U1872 (N_1872,In_1047,In_1499);
nor U1873 (N_1873,In_686,In_632);
or U1874 (N_1874,In_857,In_1453);
xnor U1875 (N_1875,In_785,In_488);
and U1876 (N_1876,In_880,In_1244);
nor U1877 (N_1877,In_1115,In_1116);
or U1878 (N_1878,In_1130,In_316);
and U1879 (N_1879,In_1479,In_1156);
or U1880 (N_1880,In_40,In_135);
xnor U1881 (N_1881,In_370,In_57);
and U1882 (N_1882,In_561,In_479);
and U1883 (N_1883,In_44,In_852);
or U1884 (N_1884,In_508,In_991);
xor U1885 (N_1885,In_1326,In_1318);
or U1886 (N_1886,In_1036,In_441);
or U1887 (N_1887,In_1091,In_663);
nor U1888 (N_1888,In_849,In_268);
or U1889 (N_1889,In_1215,In_1059);
or U1890 (N_1890,In_42,In_1128);
and U1891 (N_1891,In_323,In_1256);
nor U1892 (N_1892,In_1252,In_1022);
or U1893 (N_1893,In_969,In_1397);
xor U1894 (N_1894,In_1413,In_1308);
xnor U1895 (N_1895,In_839,In_769);
nor U1896 (N_1896,In_38,In_1187);
and U1897 (N_1897,In_371,In_14);
and U1898 (N_1898,In_1461,In_1284);
or U1899 (N_1899,In_113,In_1149);
nand U1900 (N_1900,In_1377,In_771);
or U1901 (N_1901,In_322,In_237);
or U1902 (N_1902,In_444,In_756);
nor U1903 (N_1903,In_1419,In_433);
or U1904 (N_1904,In_710,In_1334);
nand U1905 (N_1905,In_1474,In_918);
and U1906 (N_1906,In_300,In_1202);
nor U1907 (N_1907,In_921,In_36);
and U1908 (N_1908,In_178,In_892);
nor U1909 (N_1909,In_85,In_837);
nor U1910 (N_1910,In_1494,In_992);
xnor U1911 (N_1911,In_1110,In_131);
or U1912 (N_1912,In_206,In_537);
or U1913 (N_1913,In_855,In_1363);
or U1914 (N_1914,In_1229,In_541);
xor U1915 (N_1915,In_453,In_244);
nor U1916 (N_1916,In_77,In_545);
xnor U1917 (N_1917,In_768,In_636);
nor U1918 (N_1918,In_1457,In_858);
or U1919 (N_1919,In_199,In_646);
nor U1920 (N_1920,In_70,In_286);
and U1921 (N_1921,In_1026,In_852);
or U1922 (N_1922,In_747,In_433);
nand U1923 (N_1923,In_771,In_706);
nor U1924 (N_1924,In_948,In_635);
nand U1925 (N_1925,In_1297,In_1408);
nor U1926 (N_1926,In_1172,In_669);
or U1927 (N_1927,In_421,In_1013);
xnor U1928 (N_1928,In_483,In_865);
xor U1929 (N_1929,In_724,In_1258);
xnor U1930 (N_1930,In_371,In_763);
nand U1931 (N_1931,In_724,In_1496);
and U1932 (N_1932,In_714,In_1272);
and U1933 (N_1933,In_484,In_1404);
and U1934 (N_1934,In_1495,In_902);
nor U1935 (N_1935,In_355,In_884);
or U1936 (N_1936,In_985,In_731);
nand U1937 (N_1937,In_590,In_737);
and U1938 (N_1938,In_332,In_605);
nand U1939 (N_1939,In_1476,In_200);
and U1940 (N_1940,In_487,In_800);
nand U1941 (N_1941,In_603,In_650);
and U1942 (N_1942,In_837,In_860);
nor U1943 (N_1943,In_1177,In_818);
or U1944 (N_1944,In_1211,In_1048);
or U1945 (N_1945,In_799,In_1189);
xor U1946 (N_1946,In_1078,In_616);
and U1947 (N_1947,In_1375,In_140);
nand U1948 (N_1948,In_446,In_1026);
nand U1949 (N_1949,In_475,In_1393);
nor U1950 (N_1950,In_212,In_678);
xor U1951 (N_1951,In_1054,In_829);
nand U1952 (N_1952,In_158,In_1368);
xor U1953 (N_1953,In_198,In_1492);
nand U1954 (N_1954,In_993,In_935);
and U1955 (N_1955,In_963,In_374);
and U1956 (N_1956,In_1187,In_385);
and U1957 (N_1957,In_922,In_1088);
and U1958 (N_1958,In_325,In_680);
nand U1959 (N_1959,In_193,In_248);
xor U1960 (N_1960,In_321,In_943);
nor U1961 (N_1961,In_1237,In_10);
and U1962 (N_1962,In_1106,In_554);
nor U1963 (N_1963,In_1110,In_1137);
nand U1964 (N_1964,In_688,In_1039);
xnor U1965 (N_1965,In_904,In_1100);
nor U1966 (N_1966,In_698,In_1118);
and U1967 (N_1967,In_1163,In_778);
xor U1968 (N_1968,In_1178,In_41);
nor U1969 (N_1969,In_1113,In_744);
nor U1970 (N_1970,In_1004,In_612);
nand U1971 (N_1971,In_582,In_1108);
or U1972 (N_1972,In_511,In_1203);
xnor U1973 (N_1973,In_144,In_515);
and U1974 (N_1974,In_540,In_291);
xor U1975 (N_1975,In_1431,In_1021);
nand U1976 (N_1976,In_923,In_757);
and U1977 (N_1977,In_159,In_887);
or U1978 (N_1978,In_1270,In_620);
nand U1979 (N_1979,In_731,In_1311);
nand U1980 (N_1980,In_1434,In_145);
nand U1981 (N_1981,In_549,In_834);
nand U1982 (N_1982,In_983,In_1177);
and U1983 (N_1983,In_603,In_942);
xnor U1984 (N_1984,In_914,In_1103);
nand U1985 (N_1985,In_420,In_92);
and U1986 (N_1986,In_1115,In_357);
xnor U1987 (N_1987,In_552,In_401);
nand U1988 (N_1988,In_1334,In_210);
xor U1989 (N_1989,In_479,In_372);
nand U1990 (N_1990,In_300,In_1390);
nand U1991 (N_1991,In_566,In_1062);
and U1992 (N_1992,In_747,In_1110);
nand U1993 (N_1993,In_1153,In_1199);
nand U1994 (N_1994,In_1467,In_372);
or U1995 (N_1995,In_642,In_1199);
or U1996 (N_1996,In_482,In_1439);
and U1997 (N_1997,In_550,In_490);
nor U1998 (N_1998,In_267,In_1375);
or U1999 (N_1999,In_89,In_744);
nor U2000 (N_2000,In_1081,In_1130);
and U2001 (N_2001,In_56,In_952);
and U2002 (N_2002,In_26,In_953);
or U2003 (N_2003,In_6,In_1469);
nor U2004 (N_2004,In_899,In_1121);
xor U2005 (N_2005,In_544,In_957);
nor U2006 (N_2006,In_1095,In_1158);
or U2007 (N_2007,In_392,In_688);
xor U2008 (N_2008,In_1065,In_916);
xnor U2009 (N_2009,In_367,In_1201);
nor U2010 (N_2010,In_1303,In_658);
nand U2011 (N_2011,In_936,In_1083);
xnor U2012 (N_2012,In_647,In_1418);
xnor U2013 (N_2013,In_1194,In_837);
and U2014 (N_2014,In_330,In_247);
nor U2015 (N_2015,In_792,In_1162);
nor U2016 (N_2016,In_1246,In_759);
nor U2017 (N_2017,In_285,In_606);
nor U2018 (N_2018,In_395,In_648);
or U2019 (N_2019,In_904,In_1277);
and U2020 (N_2020,In_861,In_1052);
nand U2021 (N_2021,In_1302,In_1327);
or U2022 (N_2022,In_170,In_467);
nor U2023 (N_2023,In_1013,In_2);
nor U2024 (N_2024,In_97,In_273);
nand U2025 (N_2025,In_108,In_186);
nor U2026 (N_2026,In_237,In_518);
nand U2027 (N_2027,In_286,In_1287);
or U2028 (N_2028,In_1272,In_373);
xor U2029 (N_2029,In_427,In_1076);
nor U2030 (N_2030,In_1309,In_384);
nand U2031 (N_2031,In_134,In_96);
nor U2032 (N_2032,In_1451,In_417);
or U2033 (N_2033,In_213,In_473);
xor U2034 (N_2034,In_1350,In_310);
or U2035 (N_2035,In_1434,In_625);
nand U2036 (N_2036,In_1195,In_645);
and U2037 (N_2037,In_704,In_846);
nand U2038 (N_2038,In_67,In_1336);
or U2039 (N_2039,In_222,In_1255);
xor U2040 (N_2040,In_1077,In_7);
or U2041 (N_2041,In_372,In_748);
and U2042 (N_2042,In_1412,In_836);
and U2043 (N_2043,In_430,In_868);
nor U2044 (N_2044,In_429,In_904);
and U2045 (N_2045,In_397,In_851);
nand U2046 (N_2046,In_701,In_1396);
nand U2047 (N_2047,In_862,In_105);
nor U2048 (N_2048,In_616,In_719);
nand U2049 (N_2049,In_1079,In_700);
nor U2050 (N_2050,In_780,In_987);
nand U2051 (N_2051,In_682,In_918);
xnor U2052 (N_2052,In_1237,In_265);
nor U2053 (N_2053,In_289,In_649);
nor U2054 (N_2054,In_1348,In_29);
nand U2055 (N_2055,In_1294,In_254);
xnor U2056 (N_2056,In_577,In_1183);
and U2057 (N_2057,In_313,In_294);
nor U2058 (N_2058,In_828,In_661);
nand U2059 (N_2059,In_677,In_726);
or U2060 (N_2060,In_585,In_1190);
nor U2061 (N_2061,In_107,In_4);
and U2062 (N_2062,In_1366,In_303);
or U2063 (N_2063,In_1127,In_456);
xnor U2064 (N_2064,In_1237,In_921);
and U2065 (N_2065,In_516,In_803);
xnor U2066 (N_2066,In_972,In_424);
nor U2067 (N_2067,In_984,In_511);
nand U2068 (N_2068,In_266,In_1434);
or U2069 (N_2069,In_699,In_1365);
xor U2070 (N_2070,In_993,In_81);
xnor U2071 (N_2071,In_326,In_877);
and U2072 (N_2072,In_439,In_1358);
or U2073 (N_2073,In_1262,In_1352);
or U2074 (N_2074,In_262,In_1393);
or U2075 (N_2075,In_453,In_903);
nand U2076 (N_2076,In_648,In_1274);
nand U2077 (N_2077,In_310,In_34);
nor U2078 (N_2078,In_1203,In_439);
nor U2079 (N_2079,In_508,In_751);
nand U2080 (N_2080,In_366,In_996);
or U2081 (N_2081,In_1141,In_346);
or U2082 (N_2082,In_95,In_1371);
or U2083 (N_2083,In_851,In_433);
or U2084 (N_2084,In_749,In_501);
nor U2085 (N_2085,In_1266,In_304);
or U2086 (N_2086,In_344,In_581);
nor U2087 (N_2087,In_1041,In_1483);
or U2088 (N_2088,In_1456,In_136);
nor U2089 (N_2089,In_59,In_263);
or U2090 (N_2090,In_1270,In_1483);
nor U2091 (N_2091,In_781,In_473);
or U2092 (N_2092,In_87,In_246);
or U2093 (N_2093,In_740,In_723);
xor U2094 (N_2094,In_580,In_1008);
nor U2095 (N_2095,In_36,In_467);
nand U2096 (N_2096,In_208,In_837);
nor U2097 (N_2097,In_676,In_998);
nor U2098 (N_2098,In_362,In_1413);
nor U2099 (N_2099,In_368,In_1069);
xor U2100 (N_2100,In_160,In_395);
nor U2101 (N_2101,In_886,In_309);
nand U2102 (N_2102,In_433,In_641);
and U2103 (N_2103,In_769,In_1415);
nand U2104 (N_2104,In_1214,In_1002);
and U2105 (N_2105,In_1427,In_1405);
or U2106 (N_2106,In_875,In_1110);
nand U2107 (N_2107,In_785,In_866);
nand U2108 (N_2108,In_690,In_332);
xor U2109 (N_2109,In_1046,In_347);
nor U2110 (N_2110,In_285,In_969);
nand U2111 (N_2111,In_909,In_1351);
nand U2112 (N_2112,In_663,In_38);
nand U2113 (N_2113,In_646,In_564);
nand U2114 (N_2114,In_1458,In_696);
or U2115 (N_2115,In_928,In_974);
nor U2116 (N_2116,In_448,In_1029);
and U2117 (N_2117,In_1112,In_842);
xor U2118 (N_2118,In_994,In_1214);
nor U2119 (N_2119,In_49,In_134);
and U2120 (N_2120,In_505,In_982);
and U2121 (N_2121,In_1101,In_316);
nor U2122 (N_2122,In_1154,In_1336);
and U2123 (N_2123,In_546,In_804);
and U2124 (N_2124,In_901,In_529);
nor U2125 (N_2125,In_362,In_334);
or U2126 (N_2126,In_940,In_1432);
or U2127 (N_2127,In_1089,In_835);
and U2128 (N_2128,In_1439,In_58);
or U2129 (N_2129,In_163,In_106);
xor U2130 (N_2130,In_838,In_494);
nor U2131 (N_2131,In_1243,In_714);
and U2132 (N_2132,In_1206,In_459);
or U2133 (N_2133,In_344,In_7);
and U2134 (N_2134,In_438,In_729);
nor U2135 (N_2135,In_176,In_20);
nand U2136 (N_2136,In_161,In_86);
or U2137 (N_2137,In_32,In_855);
and U2138 (N_2138,In_724,In_284);
and U2139 (N_2139,In_526,In_744);
xnor U2140 (N_2140,In_283,In_1346);
or U2141 (N_2141,In_610,In_703);
nand U2142 (N_2142,In_1123,In_689);
xnor U2143 (N_2143,In_43,In_380);
nand U2144 (N_2144,In_1139,In_852);
or U2145 (N_2145,In_21,In_1307);
and U2146 (N_2146,In_1294,In_800);
and U2147 (N_2147,In_1117,In_1216);
nand U2148 (N_2148,In_483,In_263);
or U2149 (N_2149,In_640,In_7);
nand U2150 (N_2150,In_273,In_749);
xnor U2151 (N_2151,In_815,In_885);
nor U2152 (N_2152,In_1211,In_950);
or U2153 (N_2153,In_1045,In_340);
nor U2154 (N_2154,In_1217,In_957);
nor U2155 (N_2155,In_1101,In_1080);
xor U2156 (N_2156,In_1038,In_1496);
and U2157 (N_2157,In_841,In_1449);
nand U2158 (N_2158,In_748,In_1301);
nor U2159 (N_2159,In_596,In_1210);
nor U2160 (N_2160,In_447,In_1137);
or U2161 (N_2161,In_551,In_782);
xor U2162 (N_2162,In_254,In_915);
and U2163 (N_2163,In_747,In_1213);
or U2164 (N_2164,In_704,In_75);
nand U2165 (N_2165,In_1370,In_842);
nor U2166 (N_2166,In_91,In_1123);
and U2167 (N_2167,In_610,In_328);
nand U2168 (N_2168,In_214,In_1354);
nor U2169 (N_2169,In_44,In_474);
nor U2170 (N_2170,In_291,In_1212);
or U2171 (N_2171,In_1196,In_30);
and U2172 (N_2172,In_343,In_1393);
nand U2173 (N_2173,In_651,In_885);
xnor U2174 (N_2174,In_416,In_1313);
nor U2175 (N_2175,In_946,In_367);
xor U2176 (N_2176,In_1022,In_758);
and U2177 (N_2177,In_121,In_1196);
xor U2178 (N_2178,In_601,In_112);
and U2179 (N_2179,In_111,In_558);
nor U2180 (N_2180,In_632,In_712);
nand U2181 (N_2181,In_120,In_938);
or U2182 (N_2182,In_1150,In_494);
xor U2183 (N_2183,In_822,In_279);
nor U2184 (N_2184,In_103,In_1090);
or U2185 (N_2185,In_1276,In_929);
or U2186 (N_2186,In_556,In_1094);
xor U2187 (N_2187,In_654,In_665);
or U2188 (N_2188,In_56,In_716);
and U2189 (N_2189,In_1186,In_269);
nor U2190 (N_2190,In_1330,In_567);
or U2191 (N_2191,In_1146,In_739);
or U2192 (N_2192,In_202,In_1129);
and U2193 (N_2193,In_1295,In_472);
nor U2194 (N_2194,In_1440,In_1133);
and U2195 (N_2195,In_17,In_1062);
xnor U2196 (N_2196,In_1222,In_613);
nand U2197 (N_2197,In_363,In_335);
and U2198 (N_2198,In_1452,In_1265);
or U2199 (N_2199,In_253,In_515);
or U2200 (N_2200,In_1461,In_402);
or U2201 (N_2201,In_613,In_936);
or U2202 (N_2202,In_42,In_845);
or U2203 (N_2203,In_1107,In_1001);
xnor U2204 (N_2204,In_32,In_836);
xnor U2205 (N_2205,In_561,In_601);
nand U2206 (N_2206,In_252,In_396);
or U2207 (N_2207,In_861,In_452);
xor U2208 (N_2208,In_1299,In_540);
and U2209 (N_2209,In_1410,In_478);
nor U2210 (N_2210,In_1131,In_1312);
nand U2211 (N_2211,In_1193,In_99);
nor U2212 (N_2212,In_870,In_1384);
nor U2213 (N_2213,In_605,In_923);
nor U2214 (N_2214,In_61,In_899);
xor U2215 (N_2215,In_823,In_1052);
nor U2216 (N_2216,In_281,In_90);
nor U2217 (N_2217,In_201,In_693);
and U2218 (N_2218,In_974,In_1449);
xnor U2219 (N_2219,In_1242,In_994);
nor U2220 (N_2220,In_105,In_530);
nor U2221 (N_2221,In_722,In_885);
xor U2222 (N_2222,In_595,In_709);
xor U2223 (N_2223,In_1013,In_450);
or U2224 (N_2224,In_119,In_575);
nor U2225 (N_2225,In_373,In_1372);
nand U2226 (N_2226,In_181,In_469);
xnor U2227 (N_2227,In_447,In_244);
nor U2228 (N_2228,In_204,In_481);
and U2229 (N_2229,In_378,In_1237);
and U2230 (N_2230,In_956,In_1112);
or U2231 (N_2231,In_495,In_366);
nand U2232 (N_2232,In_51,In_1221);
or U2233 (N_2233,In_1042,In_1021);
or U2234 (N_2234,In_589,In_29);
nor U2235 (N_2235,In_216,In_1129);
or U2236 (N_2236,In_781,In_1222);
xnor U2237 (N_2237,In_519,In_1430);
xnor U2238 (N_2238,In_374,In_651);
nand U2239 (N_2239,In_215,In_898);
or U2240 (N_2240,In_792,In_848);
nor U2241 (N_2241,In_763,In_1247);
or U2242 (N_2242,In_1089,In_1072);
xor U2243 (N_2243,In_44,In_1206);
nand U2244 (N_2244,In_762,In_185);
xnor U2245 (N_2245,In_1400,In_1421);
xnor U2246 (N_2246,In_922,In_1355);
nor U2247 (N_2247,In_48,In_484);
nand U2248 (N_2248,In_1283,In_526);
nand U2249 (N_2249,In_118,In_454);
and U2250 (N_2250,In_1433,In_131);
and U2251 (N_2251,In_11,In_217);
xor U2252 (N_2252,In_1246,In_861);
nand U2253 (N_2253,In_1413,In_820);
nand U2254 (N_2254,In_403,In_894);
nand U2255 (N_2255,In_67,In_129);
nand U2256 (N_2256,In_253,In_543);
xor U2257 (N_2257,In_537,In_868);
or U2258 (N_2258,In_299,In_1213);
nand U2259 (N_2259,In_570,In_1325);
xnor U2260 (N_2260,In_233,In_1071);
or U2261 (N_2261,In_308,In_667);
or U2262 (N_2262,In_346,In_515);
and U2263 (N_2263,In_99,In_119);
nor U2264 (N_2264,In_422,In_988);
nor U2265 (N_2265,In_129,In_370);
nand U2266 (N_2266,In_1146,In_1389);
or U2267 (N_2267,In_932,In_403);
nor U2268 (N_2268,In_991,In_364);
or U2269 (N_2269,In_1283,In_439);
nor U2270 (N_2270,In_95,In_1495);
xor U2271 (N_2271,In_876,In_388);
and U2272 (N_2272,In_377,In_1098);
and U2273 (N_2273,In_426,In_859);
and U2274 (N_2274,In_580,In_1216);
or U2275 (N_2275,In_488,In_123);
xnor U2276 (N_2276,In_666,In_3);
nor U2277 (N_2277,In_1165,In_189);
nor U2278 (N_2278,In_1056,In_967);
nand U2279 (N_2279,In_166,In_1387);
nand U2280 (N_2280,In_668,In_1441);
nor U2281 (N_2281,In_290,In_43);
nor U2282 (N_2282,In_3,In_1389);
and U2283 (N_2283,In_1433,In_575);
and U2284 (N_2284,In_1079,In_386);
xor U2285 (N_2285,In_1226,In_1258);
and U2286 (N_2286,In_1294,In_284);
xor U2287 (N_2287,In_1426,In_268);
or U2288 (N_2288,In_18,In_964);
or U2289 (N_2289,In_778,In_1389);
nand U2290 (N_2290,In_203,In_217);
or U2291 (N_2291,In_79,In_1440);
or U2292 (N_2292,In_1102,In_1481);
or U2293 (N_2293,In_1025,In_536);
xor U2294 (N_2294,In_1230,In_486);
or U2295 (N_2295,In_812,In_1327);
nand U2296 (N_2296,In_504,In_11);
or U2297 (N_2297,In_1457,In_1029);
nor U2298 (N_2298,In_776,In_177);
nor U2299 (N_2299,In_235,In_1225);
or U2300 (N_2300,In_281,In_796);
xor U2301 (N_2301,In_1128,In_104);
or U2302 (N_2302,In_443,In_1085);
nor U2303 (N_2303,In_905,In_962);
xnor U2304 (N_2304,In_198,In_297);
nand U2305 (N_2305,In_1319,In_395);
or U2306 (N_2306,In_9,In_431);
xor U2307 (N_2307,In_239,In_637);
and U2308 (N_2308,In_543,In_452);
nand U2309 (N_2309,In_618,In_100);
or U2310 (N_2310,In_86,In_1007);
xor U2311 (N_2311,In_849,In_40);
nor U2312 (N_2312,In_16,In_262);
and U2313 (N_2313,In_649,In_82);
or U2314 (N_2314,In_1142,In_988);
and U2315 (N_2315,In_651,In_875);
and U2316 (N_2316,In_651,In_392);
nand U2317 (N_2317,In_1054,In_1297);
and U2318 (N_2318,In_1129,In_209);
and U2319 (N_2319,In_761,In_831);
nand U2320 (N_2320,In_735,In_152);
nand U2321 (N_2321,In_553,In_766);
or U2322 (N_2322,In_941,In_136);
nand U2323 (N_2323,In_492,In_767);
or U2324 (N_2324,In_867,In_32);
and U2325 (N_2325,In_517,In_969);
nor U2326 (N_2326,In_1236,In_825);
nand U2327 (N_2327,In_440,In_1295);
xnor U2328 (N_2328,In_1065,In_74);
xor U2329 (N_2329,In_272,In_491);
and U2330 (N_2330,In_998,In_275);
xnor U2331 (N_2331,In_26,In_208);
and U2332 (N_2332,In_529,In_908);
or U2333 (N_2333,In_1319,In_864);
nor U2334 (N_2334,In_917,In_430);
nand U2335 (N_2335,In_294,In_187);
or U2336 (N_2336,In_1179,In_335);
nor U2337 (N_2337,In_380,In_188);
or U2338 (N_2338,In_1333,In_1427);
xor U2339 (N_2339,In_769,In_351);
nor U2340 (N_2340,In_426,In_887);
and U2341 (N_2341,In_1324,In_471);
nor U2342 (N_2342,In_42,In_279);
xnor U2343 (N_2343,In_612,In_1301);
or U2344 (N_2344,In_1041,In_996);
nor U2345 (N_2345,In_1102,In_463);
or U2346 (N_2346,In_1239,In_1490);
nor U2347 (N_2347,In_870,In_205);
and U2348 (N_2348,In_1262,In_1379);
nand U2349 (N_2349,In_467,In_141);
nor U2350 (N_2350,In_75,In_1484);
or U2351 (N_2351,In_1178,In_472);
and U2352 (N_2352,In_423,In_1209);
or U2353 (N_2353,In_1334,In_450);
xnor U2354 (N_2354,In_888,In_1038);
xnor U2355 (N_2355,In_206,In_1049);
xor U2356 (N_2356,In_81,In_203);
nor U2357 (N_2357,In_53,In_546);
nand U2358 (N_2358,In_565,In_1156);
or U2359 (N_2359,In_649,In_891);
and U2360 (N_2360,In_1199,In_1286);
nand U2361 (N_2361,In_1092,In_1227);
or U2362 (N_2362,In_801,In_610);
xor U2363 (N_2363,In_79,In_1113);
xor U2364 (N_2364,In_1093,In_628);
xnor U2365 (N_2365,In_93,In_1132);
xor U2366 (N_2366,In_434,In_275);
or U2367 (N_2367,In_652,In_268);
and U2368 (N_2368,In_268,In_888);
nand U2369 (N_2369,In_1238,In_1423);
nand U2370 (N_2370,In_473,In_1176);
and U2371 (N_2371,In_389,In_799);
and U2372 (N_2372,In_749,In_783);
xnor U2373 (N_2373,In_760,In_913);
and U2374 (N_2374,In_878,In_1248);
nor U2375 (N_2375,In_581,In_671);
xnor U2376 (N_2376,In_603,In_1245);
or U2377 (N_2377,In_476,In_1181);
xnor U2378 (N_2378,In_968,In_449);
or U2379 (N_2379,In_1045,In_380);
nand U2380 (N_2380,In_861,In_569);
nor U2381 (N_2381,In_329,In_1221);
xnor U2382 (N_2382,In_1206,In_1385);
or U2383 (N_2383,In_1149,In_1484);
xnor U2384 (N_2384,In_256,In_328);
and U2385 (N_2385,In_770,In_744);
nor U2386 (N_2386,In_661,In_788);
and U2387 (N_2387,In_279,In_330);
nand U2388 (N_2388,In_351,In_462);
and U2389 (N_2389,In_846,In_440);
and U2390 (N_2390,In_842,In_1135);
nor U2391 (N_2391,In_1302,In_1041);
nor U2392 (N_2392,In_81,In_852);
nand U2393 (N_2393,In_906,In_281);
or U2394 (N_2394,In_1061,In_375);
xnor U2395 (N_2395,In_1055,In_772);
nand U2396 (N_2396,In_1446,In_46);
nor U2397 (N_2397,In_1248,In_1276);
xnor U2398 (N_2398,In_1494,In_970);
or U2399 (N_2399,In_971,In_496);
nand U2400 (N_2400,In_1378,In_1198);
nand U2401 (N_2401,In_445,In_969);
and U2402 (N_2402,In_1299,In_1340);
or U2403 (N_2403,In_914,In_949);
or U2404 (N_2404,In_1166,In_433);
or U2405 (N_2405,In_1339,In_608);
or U2406 (N_2406,In_265,In_245);
and U2407 (N_2407,In_792,In_172);
nand U2408 (N_2408,In_1341,In_325);
nand U2409 (N_2409,In_766,In_1327);
and U2410 (N_2410,In_446,In_1307);
and U2411 (N_2411,In_194,In_897);
nand U2412 (N_2412,In_340,In_1476);
and U2413 (N_2413,In_1309,In_429);
nor U2414 (N_2414,In_925,In_1379);
xnor U2415 (N_2415,In_698,In_262);
and U2416 (N_2416,In_764,In_367);
or U2417 (N_2417,In_1499,In_396);
nor U2418 (N_2418,In_921,In_241);
or U2419 (N_2419,In_1400,In_124);
and U2420 (N_2420,In_832,In_1131);
or U2421 (N_2421,In_910,In_709);
nand U2422 (N_2422,In_236,In_316);
or U2423 (N_2423,In_992,In_106);
nand U2424 (N_2424,In_480,In_835);
nand U2425 (N_2425,In_689,In_982);
or U2426 (N_2426,In_52,In_898);
nand U2427 (N_2427,In_36,In_945);
nor U2428 (N_2428,In_1234,In_268);
nor U2429 (N_2429,In_1187,In_1150);
or U2430 (N_2430,In_667,In_930);
or U2431 (N_2431,In_704,In_32);
and U2432 (N_2432,In_492,In_791);
nor U2433 (N_2433,In_1439,In_1103);
xnor U2434 (N_2434,In_268,In_904);
nand U2435 (N_2435,In_188,In_1344);
and U2436 (N_2436,In_912,In_1363);
nor U2437 (N_2437,In_1412,In_420);
nand U2438 (N_2438,In_1476,In_253);
xnor U2439 (N_2439,In_1486,In_22);
nor U2440 (N_2440,In_1202,In_922);
and U2441 (N_2441,In_146,In_119);
xnor U2442 (N_2442,In_1463,In_1399);
nand U2443 (N_2443,In_799,In_107);
nor U2444 (N_2444,In_1007,In_1201);
nand U2445 (N_2445,In_130,In_952);
xnor U2446 (N_2446,In_1319,In_1424);
nand U2447 (N_2447,In_1090,In_571);
nor U2448 (N_2448,In_1466,In_554);
or U2449 (N_2449,In_1342,In_656);
nand U2450 (N_2450,In_363,In_820);
nor U2451 (N_2451,In_1226,In_1036);
xnor U2452 (N_2452,In_346,In_1373);
xnor U2453 (N_2453,In_1136,In_798);
xor U2454 (N_2454,In_741,In_594);
xor U2455 (N_2455,In_386,In_1298);
nor U2456 (N_2456,In_853,In_740);
and U2457 (N_2457,In_1,In_502);
nand U2458 (N_2458,In_336,In_434);
or U2459 (N_2459,In_522,In_60);
or U2460 (N_2460,In_930,In_1421);
and U2461 (N_2461,In_515,In_466);
nor U2462 (N_2462,In_157,In_1126);
xor U2463 (N_2463,In_1487,In_714);
nor U2464 (N_2464,In_527,In_141);
xnor U2465 (N_2465,In_1449,In_1264);
nand U2466 (N_2466,In_172,In_1321);
nand U2467 (N_2467,In_52,In_1428);
and U2468 (N_2468,In_107,In_754);
or U2469 (N_2469,In_248,In_991);
xor U2470 (N_2470,In_1235,In_584);
and U2471 (N_2471,In_1279,In_436);
and U2472 (N_2472,In_382,In_290);
nor U2473 (N_2473,In_415,In_1118);
and U2474 (N_2474,In_1038,In_1473);
or U2475 (N_2475,In_347,In_1422);
xnor U2476 (N_2476,In_812,In_1412);
and U2477 (N_2477,In_735,In_523);
or U2478 (N_2478,In_676,In_1268);
nor U2479 (N_2479,In_1129,In_827);
nor U2480 (N_2480,In_1251,In_1474);
nor U2481 (N_2481,In_486,In_60);
or U2482 (N_2482,In_236,In_1211);
or U2483 (N_2483,In_1197,In_1273);
nand U2484 (N_2484,In_773,In_1004);
nand U2485 (N_2485,In_942,In_1001);
nor U2486 (N_2486,In_1029,In_960);
nor U2487 (N_2487,In_96,In_136);
nand U2488 (N_2488,In_352,In_805);
or U2489 (N_2489,In_1006,In_450);
xor U2490 (N_2490,In_638,In_569);
nand U2491 (N_2491,In_602,In_97);
xnor U2492 (N_2492,In_731,In_179);
nand U2493 (N_2493,In_1421,In_1295);
xor U2494 (N_2494,In_1271,In_965);
nor U2495 (N_2495,In_634,In_1283);
nand U2496 (N_2496,In_825,In_243);
and U2497 (N_2497,In_1333,In_548);
xor U2498 (N_2498,In_861,In_302);
nor U2499 (N_2499,In_884,In_1401);
nand U2500 (N_2500,In_277,In_275);
or U2501 (N_2501,In_403,In_1189);
or U2502 (N_2502,In_844,In_532);
and U2503 (N_2503,In_1168,In_915);
nand U2504 (N_2504,In_392,In_186);
and U2505 (N_2505,In_207,In_1353);
nand U2506 (N_2506,In_879,In_835);
nand U2507 (N_2507,In_52,In_1333);
nand U2508 (N_2508,In_0,In_631);
and U2509 (N_2509,In_1344,In_638);
nand U2510 (N_2510,In_611,In_190);
or U2511 (N_2511,In_350,In_1087);
or U2512 (N_2512,In_30,In_1249);
nor U2513 (N_2513,In_461,In_388);
xor U2514 (N_2514,In_938,In_769);
nor U2515 (N_2515,In_804,In_1157);
nand U2516 (N_2516,In_1403,In_906);
and U2517 (N_2517,In_418,In_99);
nand U2518 (N_2518,In_703,In_1481);
or U2519 (N_2519,In_591,In_344);
or U2520 (N_2520,In_1178,In_1078);
or U2521 (N_2521,In_1352,In_163);
nor U2522 (N_2522,In_126,In_790);
nand U2523 (N_2523,In_484,In_448);
nand U2524 (N_2524,In_370,In_388);
xor U2525 (N_2525,In_614,In_167);
xnor U2526 (N_2526,In_1154,In_323);
or U2527 (N_2527,In_990,In_404);
and U2528 (N_2528,In_820,In_1237);
or U2529 (N_2529,In_72,In_135);
or U2530 (N_2530,In_316,In_1246);
nor U2531 (N_2531,In_498,In_160);
xnor U2532 (N_2532,In_1069,In_486);
or U2533 (N_2533,In_440,In_426);
and U2534 (N_2534,In_940,In_337);
or U2535 (N_2535,In_1379,In_1343);
nor U2536 (N_2536,In_1346,In_484);
or U2537 (N_2537,In_24,In_1027);
xnor U2538 (N_2538,In_390,In_259);
xor U2539 (N_2539,In_245,In_286);
and U2540 (N_2540,In_644,In_2);
xnor U2541 (N_2541,In_1137,In_807);
and U2542 (N_2542,In_345,In_442);
nor U2543 (N_2543,In_1133,In_478);
or U2544 (N_2544,In_912,In_1085);
nor U2545 (N_2545,In_1492,In_1341);
nand U2546 (N_2546,In_36,In_1377);
nand U2547 (N_2547,In_247,In_1366);
nand U2548 (N_2548,In_70,In_478);
xor U2549 (N_2549,In_676,In_1489);
and U2550 (N_2550,In_1164,In_266);
nor U2551 (N_2551,In_855,In_492);
or U2552 (N_2552,In_107,In_452);
and U2553 (N_2553,In_987,In_1252);
or U2554 (N_2554,In_1172,In_281);
xor U2555 (N_2555,In_1175,In_1085);
nor U2556 (N_2556,In_1351,In_661);
xnor U2557 (N_2557,In_402,In_139);
nand U2558 (N_2558,In_443,In_632);
or U2559 (N_2559,In_354,In_1213);
xnor U2560 (N_2560,In_1255,In_1018);
and U2561 (N_2561,In_120,In_1492);
nand U2562 (N_2562,In_73,In_958);
nor U2563 (N_2563,In_1036,In_579);
or U2564 (N_2564,In_1158,In_220);
nand U2565 (N_2565,In_1032,In_1254);
nand U2566 (N_2566,In_1487,In_1472);
xor U2567 (N_2567,In_948,In_379);
xnor U2568 (N_2568,In_267,In_776);
and U2569 (N_2569,In_61,In_408);
and U2570 (N_2570,In_816,In_469);
or U2571 (N_2571,In_1051,In_1116);
and U2572 (N_2572,In_1493,In_1391);
and U2573 (N_2573,In_229,In_83);
or U2574 (N_2574,In_620,In_313);
and U2575 (N_2575,In_690,In_740);
xnor U2576 (N_2576,In_291,In_1499);
and U2577 (N_2577,In_76,In_1162);
or U2578 (N_2578,In_696,In_17);
or U2579 (N_2579,In_183,In_434);
or U2580 (N_2580,In_105,In_1168);
xor U2581 (N_2581,In_1132,In_200);
nand U2582 (N_2582,In_1378,In_122);
or U2583 (N_2583,In_1440,In_836);
nor U2584 (N_2584,In_1228,In_494);
nor U2585 (N_2585,In_1004,In_1084);
or U2586 (N_2586,In_678,In_1496);
xor U2587 (N_2587,In_959,In_149);
nand U2588 (N_2588,In_314,In_616);
or U2589 (N_2589,In_1076,In_765);
nand U2590 (N_2590,In_132,In_760);
and U2591 (N_2591,In_442,In_1264);
nand U2592 (N_2592,In_961,In_1472);
nand U2593 (N_2593,In_1224,In_1082);
xnor U2594 (N_2594,In_699,In_471);
and U2595 (N_2595,In_88,In_406);
xnor U2596 (N_2596,In_460,In_373);
nand U2597 (N_2597,In_878,In_1059);
xnor U2598 (N_2598,In_1139,In_775);
or U2599 (N_2599,In_182,In_604);
or U2600 (N_2600,In_527,In_70);
nor U2601 (N_2601,In_1229,In_863);
and U2602 (N_2602,In_788,In_765);
xor U2603 (N_2603,In_76,In_1042);
nor U2604 (N_2604,In_1473,In_552);
nor U2605 (N_2605,In_691,In_8);
nor U2606 (N_2606,In_992,In_1490);
nand U2607 (N_2607,In_209,In_141);
nand U2608 (N_2608,In_105,In_1242);
xnor U2609 (N_2609,In_969,In_823);
nand U2610 (N_2610,In_1367,In_1002);
and U2611 (N_2611,In_60,In_1117);
or U2612 (N_2612,In_293,In_953);
nand U2613 (N_2613,In_609,In_1279);
nor U2614 (N_2614,In_1379,In_306);
nand U2615 (N_2615,In_374,In_393);
or U2616 (N_2616,In_667,In_522);
nor U2617 (N_2617,In_1347,In_1473);
nand U2618 (N_2618,In_123,In_226);
or U2619 (N_2619,In_1373,In_600);
nand U2620 (N_2620,In_899,In_1418);
nor U2621 (N_2621,In_1481,In_1295);
or U2622 (N_2622,In_558,In_979);
or U2623 (N_2623,In_1359,In_750);
nand U2624 (N_2624,In_997,In_1285);
xnor U2625 (N_2625,In_92,In_1006);
xor U2626 (N_2626,In_672,In_332);
nand U2627 (N_2627,In_571,In_1388);
and U2628 (N_2628,In_806,In_958);
xor U2629 (N_2629,In_564,In_1471);
nor U2630 (N_2630,In_956,In_805);
nor U2631 (N_2631,In_783,In_1462);
nand U2632 (N_2632,In_854,In_1232);
or U2633 (N_2633,In_270,In_698);
nand U2634 (N_2634,In_262,In_705);
nor U2635 (N_2635,In_101,In_1039);
and U2636 (N_2636,In_9,In_1271);
or U2637 (N_2637,In_524,In_937);
or U2638 (N_2638,In_866,In_1214);
xnor U2639 (N_2639,In_16,In_87);
or U2640 (N_2640,In_1279,In_603);
nor U2641 (N_2641,In_650,In_844);
xor U2642 (N_2642,In_1368,In_398);
nand U2643 (N_2643,In_1131,In_1110);
nor U2644 (N_2644,In_1222,In_299);
or U2645 (N_2645,In_1182,In_540);
or U2646 (N_2646,In_1039,In_568);
xnor U2647 (N_2647,In_1273,In_375);
xnor U2648 (N_2648,In_262,In_1340);
nor U2649 (N_2649,In_8,In_272);
and U2650 (N_2650,In_1398,In_858);
or U2651 (N_2651,In_315,In_761);
xnor U2652 (N_2652,In_1253,In_1020);
and U2653 (N_2653,In_765,In_258);
or U2654 (N_2654,In_677,In_532);
and U2655 (N_2655,In_1362,In_1023);
xnor U2656 (N_2656,In_492,In_202);
nor U2657 (N_2657,In_1110,In_780);
nand U2658 (N_2658,In_858,In_937);
xnor U2659 (N_2659,In_992,In_77);
nand U2660 (N_2660,In_517,In_427);
nand U2661 (N_2661,In_790,In_1060);
nor U2662 (N_2662,In_480,In_1398);
and U2663 (N_2663,In_713,In_1001);
and U2664 (N_2664,In_780,In_246);
or U2665 (N_2665,In_703,In_1422);
and U2666 (N_2666,In_1231,In_1342);
xor U2667 (N_2667,In_1370,In_808);
and U2668 (N_2668,In_975,In_705);
xnor U2669 (N_2669,In_166,In_184);
or U2670 (N_2670,In_94,In_842);
nand U2671 (N_2671,In_166,In_811);
xnor U2672 (N_2672,In_735,In_680);
and U2673 (N_2673,In_596,In_1461);
xnor U2674 (N_2674,In_51,In_848);
or U2675 (N_2675,In_598,In_657);
nand U2676 (N_2676,In_131,In_1331);
nand U2677 (N_2677,In_840,In_71);
and U2678 (N_2678,In_724,In_1349);
xor U2679 (N_2679,In_781,In_751);
xnor U2680 (N_2680,In_1388,In_347);
nor U2681 (N_2681,In_504,In_1179);
xor U2682 (N_2682,In_575,In_1484);
nand U2683 (N_2683,In_77,In_99);
nand U2684 (N_2684,In_663,In_270);
nand U2685 (N_2685,In_373,In_497);
and U2686 (N_2686,In_269,In_254);
xnor U2687 (N_2687,In_1125,In_581);
nand U2688 (N_2688,In_453,In_920);
xnor U2689 (N_2689,In_1026,In_324);
and U2690 (N_2690,In_1254,In_970);
nand U2691 (N_2691,In_180,In_1351);
and U2692 (N_2692,In_357,In_284);
nand U2693 (N_2693,In_1268,In_781);
nor U2694 (N_2694,In_1389,In_1438);
nor U2695 (N_2695,In_1,In_748);
xor U2696 (N_2696,In_1071,In_278);
nor U2697 (N_2697,In_222,In_633);
or U2698 (N_2698,In_1216,In_834);
nand U2699 (N_2699,In_252,In_712);
and U2700 (N_2700,In_704,In_346);
or U2701 (N_2701,In_939,In_88);
nor U2702 (N_2702,In_1176,In_623);
xor U2703 (N_2703,In_1365,In_887);
or U2704 (N_2704,In_838,In_1438);
or U2705 (N_2705,In_513,In_901);
or U2706 (N_2706,In_1442,In_710);
or U2707 (N_2707,In_167,In_358);
nand U2708 (N_2708,In_1364,In_1169);
nand U2709 (N_2709,In_884,In_1426);
xnor U2710 (N_2710,In_819,In_931);
and U2711 (N_2711,In_747,In_447);
nand U2712 (N_2712,In_634,In_249);
nand U2713 (N_2713,In_1116,In_252);
or U2714 (N_2714,In_961,In_887);
nor U2715 (N_2715,In_97,In_408);
nand U2716 (N_2716,In_843,In_1174);
nand U2717 (N_2717,In_75,In_147);
nand U2718 (N_2718,In_454,In_769);
nand U2719 (N_2719,In_858,In_1205);
xnor U2720 (N_2720,In_1369,In_430);
nand U2721 (N_2721,In_612,In_1056);
or U2722 (N_2722,In_1085,In_1485);
nand U2723 (N_2723,In_1384,In_1245);
nor U2724 (N_2724,In_684,In_155);
and U2725 (N_2725,In_1048,In_1443);
and U2726 (N_2726,In_797,In_976);
xor U2727 (N_2727,In_920,In_1236);
and U2728 (N_2728,In_819,In_590);
or U2729 (N_2729,In_731,In_368);
xnor U2730 (N_2730,In_721,In_1391);
xor U2731 (N_2731,In_326,In_189);
xnor U2732 (N_2732,In_555,In_532);
nand U2733 (N_2733,In_1326,In_272);
nand U2734 (N_2734,In_480,In_1108);
or U2735 (N_2735,In_63,In_1251);
or U2736 (N_2736,In_191,In_583);
and U2737 (N_2737,In_858,In_743);
nand U2738 (N_2738,In_1438,In_596);
nand U2739 (N_2739,In_656,In_756);
and U2740 (N_2740,In_1156,In_1221);
or U2741 (N_2741,In_753,In_999);
nor U2742 (N_2742,In_1171,In_386);
nor U2743 (N_2743,In_755,In_615);
nand U2744 (N_2744,In_1313,In_1059);
nand U2745 (N_2745,In_364,In_352);
and U2746 (N_2746,In_332,In_69);
nor U2747 (N_2747,In_1010,In_1034);
nor U2748 (N_2748,In_968,In_527);
nand U2749 (N_2749,In_788,In_1144);
and U2750 (N_2750,In_1342,In_711);
or U2751 (N_2751,In_906,In_1076);
or U2752 (N_2752,In_77,In_54);
and U2753 (N_2753,In_347,In_752);
nor U2754 (N_2754,In_1354,In_93);
nor U2755 (N_2755,In_429,In_1461);
xnor U2756 (N_2756,In_246,In_1092);
and U2757 (N_2757,In_683,In_317);
and U2758 (N_2758,In_1027,In_160);
or U2759 (N_2759,In_321,In_1022);
and U2760 (N_2760,In_1244,In_660);
xnor U2761 (N_2761,In_1073,In_1223);
nor U2762 (N_2762,In_1338,In_1302);
xnor U2763 (N_2763,In_1177,In_1091);
or U2764 (N_2764,In_493,In_631);
or U2765 (N_2765,In_450,In_93);
xor U2766 (N_2766,In_710,In_719);
or U2767 (N_2767,In_955,In_209);
nand U2768 (N_2768,In_1312,In_411);
and U2769 (N_2769,In_1408,In_525);
xor U2770 (N_2770,In_153,In_1471);
and U2771 (N_2771,In_1261,In_667);
nand U2772 (N_2772,In_425,In_1416);
and U2773 (N_2773,In_449,In_872);
and U2774 (N_2774,In_278,In_1162);
or U2775 (N_2775,In_815,In_691);
nand U2776 (N_2776,In_415,In_871);
nand U2777 (N_2777,In_811,In_1478);
xor U2778 (N_2778,In_923,In_1067);
or U2779 (N_2779,In_401,In_469);
nand U2780 (N_2780,In_854,In_639);
or U2781 (N_2781,In_615,In_1054);
or U2782 (N_2782,In_1035,In_863);
and U2783 (N_2783,In_286,In_1485);
and U2784 (N_2784,In_477,In_1151);
nand U2785 (N_2785,In_297,In_745);
nand U2786 (N_2786,In_549,In_266);
xor U2787 (N_2787,In_1142,In_1213);
and U2788 (N_2788,In_879,In_130);
or U2789 (N_2789,In_891,In_1263);
nand U2790 (N_2790,In_433,In_911);
or U2791 (N_2791,In_1206,In_867);
xor U2792 (N_2792,In_543,In_1327);
or U2793 (N_2793,In_826,In_966);
nor U2794 (N_2794,In_1327,In_532);
nand U2795 (N_2795,In_1242,In_452);
and U2796 (N_2796,In_134,In_777);
or U2797 (N_2797,In_803,In_1021);
xor U2798 (N_2798,In_151,In_1412);
nand U2799 (N_2799,In_239,In_889);
nand U2800 (N_2800,In_219,In_274);
and U2801 (N_2801,In_1465,In_15);
xnor U2802 (N_2802,In_1319,In_1365);
or U2803 (N_2803,In_255,In_775);
xnor U2804 (N_2804,In_1429,In_97);
xor U2805 (N_2805,In_632,In_296);
or U2806 (N_2806,In_1460,In_597);
xor U2807 (N_2807,In_1002,In_273);
or U2808 (N_2808,In_19,In_716);
xnor U2809 (N_2809,In_219,In_1178);
and U2810 (N_2810,In_1320,In_1209);
xor U2811 (N_2811,In_181,In_30);
and U2812 (N_2812,In_1371,In_704);
xor U2813 (N_2813,In_1202,In_1456);
nor U2814 (N_2814,In_1206,In_504);
and U2815 (N_2815,In_1478,In_136);
and U2816 (N_2816,In_1242,In_816);
or U2817 (N_2817,In_1206,In_591);
xor U2818 (N_2818,In_879,In_561);
or U2819 (N_2819,In_733,In_697);
and U2820 (N_2820,In_1131,In_370);
nor U2821 (N_2821,In_531,In_122);
nand U2822 (N_2822,In_238,In_730);
nand U2823 (N_2823,In_214,In_1233);
and U2824 (N_2824,In_963,In_353);
or U2825 (N_2825,In_723,In_1184);
xor U2826 (N_2826,In_81,In_807);
nand U2827 (N_2827,In_1004,In_1450);
or U2828 (N_2828,In_525,In_167);
nand U2829 (N_2829,In_933,In_682);
nor U2830 (N_2830,In_1151,In_1410);
and U2831 (N_2831,In_312,In_1078);
or U2832 (N_2832,In_398,In_1347);
nand U2833 (N_2833,In_1356,In_883);
xnor U2834 (N_2834,In_627,In_1460);
nor U2835 (N_2835,In_1278,In_152);
nand U2836 (N_2836,In_1188,In_108);
nand U2837 (N_2837,In_1275,In_1046);
xor U2838 (N_2838,In_516,In_1345);
and U2839 (N_2839,In_283,In_627);
nor U2840 (N_2840,In_384,In_1166);
and U2841 (N_2841,In_870,In_206);
and U2842 (N_2842,In_128,In_320);
nand U2843 (N_2843,In_450,In_104);
nand U2844 (N_2844,In_567,In_101);
nor U2845 (N_2845,In_832,In_1149);
nand U2846 (N_2846,In_540,In_1141);
or U2847 (N_2847,In_419,In_1000);
and U2848 (N_2848,In_747,In_1157);
or U2849 (N_2849,In_671,In_1081);
nor U2850 (N_2850,In_946,In_1259);
and U2851 (N_2851,In_1367,In_1098);
xnor U2852 (N_2852,In_504,In_1378);
nor U2853 (N_2853,In_1065,In_771);
or U2854 (N_2854,In_552,In_1489);
nand U2855 (N_2855,In_40,In_74);
and U2856 (N_2856,In_700,In_780);
nor U2857 (N_2857,In_1433,In_178);
and U2858 (N_2858,In_823,In_639);
nor U2859 (N_2859,In_782,In_1412);
or U2860 (N_2860,In_373,In_34);
and U2861 (N_2861,In_1179,In_597);
xnor U2862 (N_2862,In_154,In_1394);
and U2863 (N_2863,In_165,In_258);
nand U2864 (N_2864,In_1286,In_362);
or U2865 (N_2865,In_1024,In_743);
and U2866 (N_2866,In_673,In_1383);
or U2867 (N_2867,In_1129,In_465);
xnor U2868 (N_2868,In_1063,In_1220);
or U2869 (N_2869,In_325,In_392);
and U2870 (N_2870,In_1158,In_875);
and U2871 (N_2871,In_879,In_476);
or U2872 (N_2872,In_1446,In_436);
nor U2873 (N_2873,In_653,In_390);
or U2874 (N_2874,In_794,In_1249);
nand U2875 (N_2875,In_1366,In_1034);
or U2876 (N_2876,In_1053,In_205);
nor U2877 (N_2877,In_391,In_393);
or U2878 (N_2878,In_1464,In_1051);
nand U2879 (N_2879,In_724,In_1352);
or U2880 (N_2880,In_949,In_129);
or U2881 (N_2881,In_955,In_1440);
nand U2882 (N_2882,In_1071,In_1182);
xor U2883 (N_2883,In_630,In_1028);
and U2884 (N_2884,In_734,In_880);
and U2885 (N_2885,In_1269,In_367);
and U2886 (N_2886,In_930,In_1405);
xnor U2887 (N_2887,In_1328,In_1428);
and U2888 (N_2888,In_1066,In_1127);
nand U2889 (N_2889,In_1224,In_297);
or U2890 (N_2890,In_429,In_160);
xor U2891 (N_2891,In_924,In_677);
nor U2892 (N_2892,In_364,In_964);
or U2893 (N_2893,In_941,In_1203);
nand U2894 (N_2894,In_817,In_1079);
nand U2895 (N_2895,In_208,In_266);
xnor U2896 (N_2896,In_567,In_307);
nand U2897 (N_2897,In_51,In_625);
nand U2898 (N_2898,In_183,In_910);
and U2899 (N_2899,In_1045,In_215);
nand U2900 (N_2900,In_46,In_1164);
nand U2901 (N_2901,In_829,In_1192);
xor U2902 (N_2902,In_243,In_487);
and U2903 (N_2903,In_1205,In_778);
nor U2904 (N_2904,In_276,In_1102);
or U2905 (N_2905,In_1293,In_324);
nand U2906 (N_2906,In_1219,In_1484);
nor U2907 (N_2907,In_190,In_164);
xnor U2908 (N_2908,In_819,In_1449);
nor U2909 (N_2909,In_577,In_224);
or U2910 (N_2910,In_1004,In_208);
and U2911 (N_2911,In_1050,In_1058);
nand U2912 (N_2912,In_242,In_808);
or U2913 (N_2913,In_185,In_1154);
or U2914 (N_2914,In_509,In_1003);
xor U2915 (N_2915,In_328,In_1093);
xor U2916 (N_2916,In_1426,In_1027);
xnor U2917 (N_2917,In_1339,In_366);
nand U2918 (N_2918,In_1180,In_1086);
xnor U2919 (N_2919,In_1225,In_433);
nor U2920 (N_2920,In_378,In_293);
xor U2921 (N_2921,In_401,In_268);
or U2922 (N_2922,In_404,In_912);
nor U2923 (N_2923,In_428,In_778);
or U2924 (N_2924,In_954,In_16);
nand U2925 (N_2925,In_941,In_631);
or U2926 (N_2926,In_502,In_472);
nor U2927 (N_2927,In_1147,In_835);
nor U2928 (N_2928,In_772,In_724);
nor U2929 (N_2929,In_994,In_970);
and U2930 (N_2930,In_289,In_1180);
xor U2931 (N_2931,In_466,In_1348);
nand U2932 (N_2932,In_906,In_718);
nor U2933 (N_2933,In_371,In_1430);
and U2934 (N_2934,In_689,In_364);
and U2935 (N_2935,In_293,In_959);
xor U2936 (N_2936,In_1432,In_315);
nor U2937 (N_2937,In_575,In_794);
and U2938 (N_2938,In_1066,In_921);
nor U2939 (N_2939,In_1140,In_1448);
and U2940 (N_2940,In_682,In_291);
xor U2941 (N_2941,In_478,In_717);
or U2942 (N_2942,In_173,In_1045);
xnor U2943 (N_2943,In_833,In_896);
nor U2944 (N_2944,In_611,In_985);
nand U2945 (N_2945,In_947,In_1476);
nor U2946 (N_2946,In_669,In_1137);
nand U2947 (N_2947,In_802,In_952);
nand U2948 (N_2948,In_684,In_138);
xnor U2949 (N_2949,In_1471,In_953);
or U2950 (N_2950,In_190,In_361);
or U2951 (N_2951,In_945,In_701);
and U2952 (N_2952,In_83,In_556);
xor U2953 (N_2953,In_1490,In_1325);
nand U2954 (N_2954,In_1370,In_1132);
or U2955 (N_2955,In_585,In_329);
and U2956 (N_2956,In_1255,In_55);
and U2957 (N_2957,In_1165,In_799);
or U2958 (N_2958,In_845,In_282);
and U2959 (N_2959,In_1254,In_1324);
and U2960 (N_2960,In_1187,In_762);
xor U2961 (N_2961,In_121,In_790);
and U2962 (N_2962,In_975,In_934);
nor U2963 (N_2963,In_1048,In_441);
nand U2964 (N_2964,In_510,In_1258);
or U2965 (N_2965,In_761,In_841);
and U2966 (N_2966,In_967,In_1349);
xor U2967 (N_2967,In_318,In_857);
and U2968 (N_2968,In_1074,In_808);
nor U2969 (N_2969,In_1298,In_554);
nor U2970 (N_2970,In_816,In_1404);
nor U2971 (N_2971,In_695,In_148);
xor U2972 (N_2972,In_750,In_129);
nor U2973 (N_2973,In_667,In_626);
xnor U2974 (N_2974,In_253,In_1452);
or U2975 (N_2975,In_1317,In_1231);
nand U2976 (N_2976,In_210,In_948);
or U2977 (N_2977,In_547,In_249);
or U2978 (N_2978,In_120,In_767);
or U2979 (N_2979,In_796,In_1365);
and U2980 (N_2980,In_1403,In_997);
nor U2981 (N_2981,In_1394,In_1436);
or U2982 (N_2982,In_1213,In_1286);
xnor U2983 (N_2983,In_424,In_790);
nand U2984 (N_2984,In_807,In_1266);
and U2985 (N_2985,In_1187,In_859);
nand U2986 (N_2986,In_1358,In_878);
nor U2987 (N_2987,In_912,In_1469);
and U2988 (N_2988,In_1092,In_730);
and U2989 (N_2989,In_1177,In_1466);
nor U2990 (N_2990,In_256,In_1108);
xor U2991 (N_2991,In_758,In_178);
nand U2992 (N_2992,In_564,In_766);
nand U2993 (N_2993,In_492,In_1043);
or U2994 (N_2994,In_1329,In_325);
or U2995 (N_2995,In_54,In_1246);
or U2996 (N_2996,In_1116,In_1373);
or U2997 (N_2997,In_61,In_1050);
nand U2998 (N_2998,In_359,In_393);
and U2999 (N_2999,In_448,In_1241);
nor U3000 (N_3000,In_139,In_625);
nor U3001 (N_3001,In_1227,In_1000);
and U3002 (N_3002,In_534,In_1232);
or U3003 (N_3003,In_1154,In_42);
nor U3004 (N_3004,In_321,In_404);
xor U3005 (N_3005,In_714,In_52);
xnor U3006 (N_3006,In_513,In_1010);
nand U3007 (N_3007,In_702,In_493);
nand U3008 (N_3008,In_507,In_849);
or U3009 (N_3009,In_692,In_877);
and U3010 (N_3010,In_1123,In_627);
nand U3011 (N_3011,In_1421,In_710);
or U3012 (N_3012,In_28,In_178);
xor U3013 (N_3013,In_1183,In_658);
nand U3014 (N_3014,In_75,In_800);
or U3015 (N_3015,In_1358,In_57);
nand U3016 (N_3016,In_16,In_575);
nand U3017 (N_3017,In_1333,In_884);
nand U3018 (N_3018,In_809,In_981);
or U3019 (N_3019,In_676,In_1319);
nor U3020 (N_3020,In_1266,In_819);
nand U3021 (N_3021,In_1438,In_530);
or U3022 (N_3022,In_345,In_227);
nor U3023 (N_3023,In_1015,In_1394);
xor U3024 (N_3024,In_1188,In_309);
nand U3025 (N_3025,In_129,In_18);
and U3026 (N_3026,In_164,In_535);
nand U3027 (N_3027,In_1243,In_927);
or U3028 (N_3028,In_553,In_1289);
xor U3029 (N_3029,In_1326,In_516);
xnor U3030 (N_3030,In_1025,In_624);
nand U3031 (N_3031,In_1306,In_454);
or U3032 (N_3032,In_1217,In_1040);
xnor U3033 (N_3033,In_1103,In_1419);
or U3034 (N_3034,In_393,In_721);
nand U3035 (N_3035,In_768,In_821);
xnor U3036 (N_3036,In_312,In_679);
nand U3037 (N_3037,In_364,In_930);
nand U3038 (N_3038,In_559,In_693);
and U3039 (N_3039,In_345,In_280);
nand U3040 (N_3040,In_490,In_594);
nor U3041 (N_3041,In_1283,In_1469);
nor U3042 (N_3042,In_4,In_907);
xnor U3043 (N_3043,In_252,In_1499);
nand U3044 (N_3044,In_474,In_1253);
xor U3045 (N_3045,In_485,In_882);
nor U3046 (N_3046,In_1434,In_880);
xnor U3047 (N_3047,In_581,In_1481);
and U3048 (N_3048,In_1354,In_932);
and U3049 (N_3049,In_268,In_977);
or U3050 (N_3050,In_1385,In_838);
and U3051 (N_3051,In_1438,In_439);
nor U3052 (N_3052,In_894,In_548);
nand U3053 (N_3053,In_915,In_348);
xnor U3054 (N_3054,In_1154,In_815);
and U3055 (N_3055,In_1395,In_161);
xor U3056 (N_3056,In_1307,In_858);
nand U3057 (N_3057,In_1171,In_1139);
xor U3058 (N_3058,In_99,In_363);
xnor U3059 (N_3059,In_1270,In_168);
or U3060 (N_3060,In_1286,In_833);
xor U3061 (N_3061,In_572,In_1442);
and U3062 (N_3062,In_963,In_996);
xnor U3063 (N_3063,In_488,In_650);
and U3064 (N_3064,In_793,In_213);
or U3065 (N_3065,In_896,In_753);
nor U3066 (N_3066,In_81,In_1080);
or U3067 (N_3067,In_1269,In_339);
or U3068 (N_3068,In_390,In_1159);
xnor U3069 (N_3069,In_716,In_1235);
or U3070 (N_3070,In_1483,In_981);
or U3071 (N_3071,In_950,In_1352);
and U3072 (N_3072,In_156,In_653);
and U3073 (N_3073,In_704,In_486);
nor U3074 (N_3074,In_842,In_379);
and U3075 (N_3075,In_857,In_955);
and U3076 (N_3076,In_466,In_1216);
and U3077 (N_3077,In_623,In_103);
nor U3078 (N_3078,In_506,In_967);
and U3079 (N_3079,In_504,In_1034);
nor U3080 (N_3080,In_604,In_1300);
xnor U3081 (N_3081,In_204,In_677);
xnor U3082 (N_3082,In_650,In_1104);
and U3083 (N_3083,In_509,In_995);
nor U3084 (N_3084,In_421,In_676);
nand U3085 (N_3085,In_1125,In_1201);
nor U3086 (N_3086,In_792,In_674);
and U3087 (N_3087,In_1194,In_1090);
nand U3088 (N_3088,In_556,In_826);
nor U3089 (N_3089,In_268,In_200);
xor U3090 (N_3090,In_1252,In_1467);
nand U3091 (N_3091,In_5,In_399);
and U3092 (N_3092,In_712,In_320);
nand U3093 (N_3093,In_724,In_594);
nand U3094 (N_3094,In_778,In_1032);
and U3095 (N_3095,In_576,In_442);
xnor U3096 (N_3096,In_220,In_348);
and U3097 (N_3097,In_763,In_308);
xnor U3098 (N_3098,In_666,In_1096);
nor U3099 (N_3099,In_1357,In_580);
xnor U3100 (N_3100,In_449,In_483);
or U3101 (N_3101,In_765,In_1247);
and U3102 (N_3102,In_767,In_321);
xnor U3103 (N_3103,In_542,In_4);
nand U3104 (N_3104,In_1283,In_1393);
xnor U3105 (N_3105,In_5,In_1257);
nor U3106 (N_3106,In_264,In_122);
xor U3107 (N_3107,In_747,In_250);
or U3108 (N_3108,In_1491,In_431);
xor U3109 (N_3109,In_308,In_1490);
nor U3110 (N_3110,In_916,In_965);
nand U3111 (N_3111,In_1438,In_55);
or U3112 (N_3112,In_1164,In_35);
and U3113 (N_3113,In_235,In_1354);
and U3114 (N_3114,In_893,In_476);
xnor U3115 (N_3115,In_644,In_235);
nor U3116 (N_3116,In_878,In_1328);
or U3117 (N_3117,In_1237,In_440);
or U3118 (N_3118,In_181,In_1321);
nand U3119 (N_3119,In_27,In_591);
nand U3120 (N_3120,In_534,In_264);
xnor U3121 (N_3121,In_823,In_419);
or U3122 (N_3122,In_642,In_120);
nand U3123 (N_3123,In_998,In_34);
and U3124 (N_3124,In_1037,In_512);
or U3125 (N_3125,In_195,In_1157);
nand U3126 (N_3126,In_1393,In_774);
and U3127 (N_3127,In_297,In_199);
nor U3128 (N_3128,In_22,In_464);
xnor U3129 (N_3129,In_774,In_1240);
nand U3130 (N_3130,In_1132,In_923);
nor U3131 (N_3131,In_710,In_667);
and U3132 (N_3132,In_797,In_69);
xnor U3133 (N_3133,In_1366,In_170);
nand U3134 (N_3134,In_960,In_580);
and U3135 (N_3135,In_821,In_556);
nor U3136 (N_3136,In_1293,In_1016);
nor U3137 (N_3137,In_965,In_1255);
nor U3138 (N_3138,In_730,In_303);
nand U3139 (N_3139,In_1230,In_663);
or U3140 (N_3140,In_278,In_619);
and U3141 (N_3141,In_105,In_518);
or U3142 (N_3142,In_800,In_671);
nor U3143 (N_3143,In_500,In_135);
nand U3144 (N_3144,In_158,In_993);
nor U3145 (N_3145,In_1456,In_1130);
nor U3146 (N_3146,In_175,In_553);
xor U3147 (N_3147,In_1222,In_202);
and U3148 (N_3148,In_1084,In_261);
xnor U3149 (N_3149,In_1203,In_202);
xnor U3150 (N_3150,In_802,In_470);
or U3151 (N_3151,In_1483,In_498);
nand U3152 (N_3152,In_1167,In_633);
or U3153 (N_3153,In_1428,In_1169);
xor U3154 (N_3154,In_15,In_902);
xor U3155 (N_3155,In_1091,In_256);
or U3156 (N_3156,In_877,In_1375);
and U3157 (N_3157,In_277,In_974);
xnor U3158 (N_3158,In_1014,In_842);
and U3159 (N_3159,In_262,In_1051);
and U3160 (N_3160,In_809,In_1170);
or U3161 (N_3161,In_1397,In_531);
or U3162 (N_3162,In_825,In_1334);
nand U3163 (N_3163,In_1060,In_829);
nor U3164 (N_3164,In_27,In_1137);
nand U3165 (N_3165,In_482,In_1490);
nand U3166 (N_3166,In_928,In_995);
xnor U3167 (N_3167,In_852,In_937);
or U3168 (N_3168,In_392,In_1227);
nand U3169 (N_3169,In_146,In_638);
nand U3170 (N_3170,In_871,In_587);
xnor U3171 (N_3171,In_318,In_1115);
and U3172 (N_3172,In_575,In_533);
or U3173 (N_3173,In_1133,In_1360);
nand U3174 (N_3174,In_359,In_86);
nor U3175 (N_3175,In_659,In_172);
nor U3176 (N_3176,In_878,In_1273);
and U3177 (N_3177,In_904,In_410);
and U3178 (N_3178,In_967,In_748);
and U3179 (N_3179,In_1357,In_1410);
xnor U3180 (N_3180,In_805,In_63);
xnor U3181 (N_3181,In_263,In_757);
nand U3182 (N_3182,In_305,In_170);
xor U3183 (N_3183,In_705,In_1244);
and U3184 (N_3184,In_1200,In_944);
and U3185 (N_3185,In_869,In_1197);
xnor U3186 (N_3186,In_498,In_1492);
and U3187 (N_3187,In_1260,In_1207);
or U3188 (N_3188,In_939,In_561);
nor U3189 (N_3189,In_853,In_383);
or U3190 (N_3190,In_927,In_1041);
nor U3191 (N_3191,In_569,In_654);
and U3192 (N_3192,In_675,In_1260);
and U3193 (N_3193,In_987,In_1130);
nor U3194 (N_3194,In_1467,In_131);
nand U3195 (N_3195,In_509,In_8);
or U3196 (N_3196,In_450,In_781);
or U3197 (N_3197,In_490,In_1217);
and U3198 (N_3198,In_77,In_1211);
xor U3199 (N_3199,In_1189,In_284);
xnor U3200 (N_3200,In_1372,In_1055);
or U3201 (N_3201,In_431,In_463);
and U3202 (N_3202,In_975,In_1393);
xnor U3203 (N_3203,In_646,In_327);
xor U3204 (N_3204,In_1219,In_324);
xor U3205 (N_3205,In_962,In_86);
or U3206 (N_3206,In_341,In_698);
nor U3207 (N_3207,In_1388,In_373);
or U3208 (N_3208,In_1307,In_861);
and U3209 (N_3209,In_766,In_1223);
nand U3210 (N_3210,In_330,In_49);
xor U3211 (N_3211,In_540,In_514);
and U3212 (N_3212,In_1077,In_169);
nand U3213 (N_3213,In_467,In_39);
xnor U3214 (N_3214,In_1252,In_510);
xor U3215 (N_3215,In_278,In_857);
xor U3216 (N_3216,In_707,In_842);
xor U3217 (N_3217,In_331,In_635);
or U3218 (N_3218,In_1221,In_823);
xnor U3219 (N_3219,In_1002,In_782);
nand U3220 (N_3220,In_714,In_1120);
xor U3221 (N_3221,In_1076,In_1146);
nand U3222 (N_3222,In_1165,In_1233);
xnor U3223 (N_3223,In_319,In_192);
nor U3224 (N_3224,In_863,In_179);
nand U3225 (N_3225,In_444,In_1268);
nor U3226 (N_3226,In_278,In_1379);
nand U3227 (N_3227,In_1272,In_1346);
xor U3228 (N_3228,In_1480,In_849);
xor U3229 (N_3229,In_773,In_530);
or U3230 (N_3230,In_686,In_1254);
xor U3231 (N_3231,In_477,In_865);
xor U3232 (N_3232,In_715,In_1140);
xor U3233 (N_3233,In_539,In_549);
xnor U3234 (N_3234,In_945,In_1467);
nand U3235 (N_3235,In_651,In_825);
xnor U3236 (N_3236,In_978,In_170);
and U3237 (N_3237,In_160,In_550);
and U3238 (N_3238,In_61,In_1371);
nand U3239 (N_3239,In_438,In_661);
nor U3240 (N_3240,In_456,In_1400);
and U3241 (N_3241,In_1405,In_113);
xor U3242 (N_3242,In_578,In_184);
nor U3243 (N_3243,In_1018,In_296);
and U3244 (N_3244,In_1248,In_797);
nand U3245 (N_3245,In_368,In_865);
xnor U3246 (N_3246,In_404,In_1023);
xnor U3247 (N_3247,In_445,In_269);
and U3248 (N_3248,In_664,In_928);
or U3249 (N_3249,In_928,In_481);
or U3250 (N_3250,In_508,In_889);
nand U3251 (N_3251,In_420,In_1019);
xor U3252 (N_3252,In_1463,In_506);
or U3253 (N_3253,In_334,In_872);
nor U3254 (N_3254,In_1164,In_1109);
nor U3255 (N_3255,In_1436,In_111);
and U3256 (N_3256,In_983,In_999);
nand U3257 (N_3257,In_785,In_892);
nand U3258 (N_3258,In_111,In_1313);
and U3259 (N_3259,In_1387,In_1311);
nand U3260 (N_3260,In_276,In_1143);
or U3261 (N_3261,In_1113,In_1421);
or U3262 (N_3262,In_746,In_342);
or U3263 (N_3263,In_705,In_1140);
or U3264 (N_3264,In_652,In_218);
or U3265 (N_3265,In_353,In_377);
nand U3266 (N_3266,In_1407,In_974);
and U3267 (N_3267,In_198,In_902);
nor U3268 (N_3268,In_1062,In_475);
nor U3269 (N_3269,In_1132,In_1272);
or U3270 (N_3270,In_563,In_1087);
xor U3271 (N_3271,In_668,In_1110);
nor U3272 (N_3272,In_512,In_1115);
nor U3273 (N_3273,In_495,In_549);
nor U3274 (N_3274,In_31,In_1103);
or U3275 (N_3275,In_1389,In_179);
xnor U3276 (N_3276,In_563,In_1248);
xor U3277 (N_3277,In_156,In_1224);
nand U3278 (N_3278,In_633,In_514);
nand U3279 (N_3279,In_366,In_193);
xor U3280 (N_3280,In_957,In_661);
or U3281 (N_3281,In_1456,In_828);
nor U3282 (N_3282,In_1334,In_1113);
nor U3283 (N_3283,In_1209,In_158);
xor U3284 (N_3284,In_847,In_1373);
and U3285 (N_3285,In_338,In_53);
nand U3286 (N_3286,In_1401,In_206);
nor U3287 (N_3287,In_1290,In_1446);
nor U3288 (N_3288,In_565,In_460);
nor U3289 (N_3289,In_606,In_188);
nor U3290 (N_3290,In_1234,In_306);
xnor U3291 (N_3291,In_1313,In_1146);
nand U3292 (N_3292,In_804,In_104);
nor U3293 (N_3293,In_386,In_700);
and U3294 (N_3294,In_138,In_532);
xnor U3295 (N_3295,In_1444,In_1085);
or U3296 (N_3296,In_1191,In_1102);
or U3297 (N_3297,In_498,In_1274);
xnor U3298 (N_3298,In_639,In_62);
and U3299 (N_3299,In_1103,In_223);
nor U3300 (N_3300,In_619,In_1048);
nand U3301 (N_3301,In_24,In_987);
nand U3302 (N_3302,In_1262,In_954);
or U3303 (N_3303,In_799,In_1299);
xor U3304 (N_3304,In_26,In_1481);
and U3305 (N_3305,In_1205,In_71);
nand U3306 (N_3306,In_695,In_189);
or U3307 (N_3307,In_643,In_24);
or U3308 (N_3308,In_1251,In_1433);
nor U3309 (N_3309,In_166,In_1463);
nor U3310 (N_3310,In_796,In_1136);
nand U3311 (N_3311,In_1487,In_460);
and U3312 (N_3312,In_709,In_376);
xnor U3313 (N_3313,In_883,In_35);
or U3314 (N_3314,In_639,In_755);
xnor U3315 (N_3315,In_724,In_1384);
nor U3316 (N_3316,In_1470,In_986);
nor U3317 (N_3317,In_1309,In_1315);
nor U3318 (N_3318,In_928,In_145);
and U3319 (N_3319,In_694,In_61);
nor U3320 (N_3320,In_304,In_465);
xor U3321 (N_3321,In_566,In_1004);
xor U3322 (N_3322,In_371,In_1373);
and U3323 (N_3323,In_1379,In_418);
or U3324 (N_3324,In_875,In_236);
xor U3325 (N_3325,In_284,In_830);
or U3326 (N_3326,In_841,In_970);
nand U3327 (N_3327,In_1402,In_51);
and U3328 (N_3328,In_877,In_144);
nand U3329 (N_3329,In_1081,In_839);
nor U3330 (N_3330,In_822,In_1186);
nand U3331 (N_3331,In_269,In_708);
nor U3332 (N_3332,In_1427,In_684);
or U3333 (N_3333,In_449,In_305);
nor U3334 (N_3334,In_82,In_502);
or U3335 (N_3335,In_981,In_764);
or U3336 (N_3336,In_1377,In_549);
xnor U3337 (N_3337,In_726,In_528);
and U3338 (N_3338,In_414,In_816);
or U3339 (N_3339,In_1231,In_1306);
or U3340 (N_3340,In_1303,In_935);
nand U3341 (N_3341,In_52,In_366);
nor U3342 (N_3342,In_533,In_845);
or U3343 (N_3343,In_0,In_1451);
and U3344 (N_3344,In_502,In_302);
nor U3345 (N_3345,In_351,In_544);
and U3346 (N_3346,In_741,In_538);
and U3347 (N_3347,In_824,In_1175);
nand U3348 (N_3348,In_1476,In_542);
or U3349 (N_3349,In_814,In_919);
or U3350 (N_3350,In_648,In_892);
and U3351 (N_3351,In_511,In_1020);
xor U3352 (N_3352,In_539,In_1145);
nor U3353 (N_3353,In_521,In_675);
and U3354 (N_3354,In_965,In_1023);
or U3355 (N_3355,In_695,In_331);
and U3356 (N_3356,In_317,In_398);
or U3357 (N_3357,In_200,In_66);
or U3358 (N_3358,In_609,In_1178);
nor U3359 (N_3359,In_1023,In_394);
or U3360 (N_3360,In_223,In_1170);
xnor U3361 (N_3361,In_307,In_157);
nand U3362 (N_3362,In_934,In_670);
xnor U3363 (N_3363,In_1087,In_990);
and U3364 (N_3364,In_1037,In_1494);
or U3365 (N_3365,In_549,In_349);
or U3366 (N_3366,In_1099,In_883);
or U3367 (N_3367,In_94,In_1157);
or U3368 (N_3368,In_157,In_840);
xor U3369 (N_3369,In_1142,In_633);
and U3370 (N_3370,In_1432,In_428);
nand U3371 (N_3371,In_220,In_1080);
xor U3372 (N_3372,In_1301,In_1481);
or U3373 (N_3373,In_83,In_904);
and U3374 (N_3374,In_581,In_1049);
and U3375 (N_3375,In_42,In_516);
xnor U3376 (N_3376,In_1433,In_353);
or U3377 (N_3377,In_1144,In_1364);
and U3378 (N_3378,In_362,In_617);
xor U3379 (N_3379,In_674,In_488);
nand U3380 (N_3380,In_1244,In_605);
nor U3381 (N_3381,In_218,In_269);
nand U3382 (N_3382,In_1271,In_730);
and U3383 (N_3383,In_786,In_242);
and U3384 (N_3384,In_1281,In_849);
or U3385 (N_3385,In_1209,In_403);
and U3386 (N_3386,In_1223,In_879);
xor U3387 (N_3387,In_867,In_273);
and U3388 (N_3388,In_817,In_412);
nand U3389 (N_3389,In_664,In_670);
nor U3390 (N_3390,In_1331,In_164);
nand U3391 (N_3391,In_741,In_1218);
nand U3392 (N_3392,In_502,In_344);
or U3393 (N_3393,In_224,In_407);
xor U3394 (N_3394,In_586,In_623);
xnor U3395 (N_3395,In_874,In_1132);
and U3396 (N_3396,In_333,In_1167);
nor U3397 (N_3397,In_896,In_1425);
and U3398 (N_3398,In_379,In_687);
and U3399 (N_3399,In_1103,In_225);
xnor U3400 (N_3400,In_1245,In_371);
xnor U3401 (N_3401,In_1042,In_1187);
xor U3402 (N_3402,In_484,In_1073);
nand U3403 (N_3403,In_89,In_768);
nor U3404 (N_3404,In_1469,In_111);
or U3405 (N_3405,In_14,In_334);
nor U3406 (N_3406,In_692,In_631);
nand U3407 (N_3407,In_1172,In_274);
nor U3408 (N_3408,In_958,In_1369);
and U3409 (N_3409,In_10,In_556);
and U3410 (N_3410,In_96,In_1161);
nand U3411 (N_3411,In_4,In_587);
nor U3412 (N_3412,In_522,In_639);
nand U3413 (N_3413,In_71,In_1235);
and U3414 (N_3414,In_816,In_1002);
nor U3415 (N_3415,In_592,In_252);
nor U3416 (N_3416,In_634,In_1323);
and U3417 (N_3417,In_1039,In_1063);
or U3418 (N_3418,In_163,In_804);
and U3419 (N_3419,In_905,In_165);
xnor U3420 (N_3420,In_265,In_173);
or U3421 (N_3421,In_405,In_869);
nor U3422 (N_3422,In_1421,In_1464);
and U3423 (N_3423,In_772,In_491);
or U3424 (N_3424,In_307,In_699);
or U3425 (N_3425,In_205,In_1079);
nand U3426 (N_3426,In_1227,In_782);
nor U3427 (N_3427,In_771,In_280);
xor U3428 (N_3428,In_815,In_162);
nand U3429 (N_3429,In_1198,In_550);
and U3430 (N_3430,In_995,In_1250);
nor U3431 (N_3431,In_1050,In_1069);
or U3432 (N_3432,In_711,In_47);
nand U3433 (N_3433,In_1484,In_449);
and U3434 (N_3434,In_1148,In_1476);
and U3435 (N_3435,In_25,In_1046);
nor U3436 (N_3436,In_1356,In_754);
and U3437 (N_3437,In_1450,In_811);
or U3438 (N_3438,In_865,In_454);
xor U3439 (N_3439,In_658,In_889);
and U3440 (N_3440,In_284,In_1003);
xor U3441 (N_3441,In_1485,In_1272);
nor U3442 (N_3442,In_929,In_401);
nor U3443 (N_3443,In_1300,In_1459);
and U3444 (N_3444,In_140,In_467);
or U3445 (N_3445,In_1259,In_1449);
nand U3446 (N_3446,In_331,In_125);
nor U3447 (N_3447,In_146,In_1134);
nor U3448 (N_3448,In_275,In_716);
nand U3449 (N_3449,In_1169,In_292);
and U3450 (N_3450,In_754,In_453);
nand U3451 (N_3451,In_128,In_683);
and U3452 (N_3452,In_137,In_1077);
nand U3453 (N_3453,In_390,In_707);
or U3454 (N_3454,In_432,In_1140);
and U3455 (N_3455,In_1095,In_854);
xor U3456 (N_3456,In_490,In_266);
and U3457 (N_3457,In_622,In_1117);
or U3458 (N_3458,In_1253,In_1194);
nand U3459 (N_3459,In_985,In_56);
nand U3460 (N_3460,In_498,In_1104);
nor U3461 (N_3461,In_935,In_776);
nor U3462 (N_3462,In_250,In_384);
xnor U3463 (N_3463,In_512,In_843);
or U3464 (N_3464,In_396,In_1186);
and U3465 (N_3465,In_819,In_220);
xnor U3466 (N_3466,In_710,In_846);
nor U3467 (N_3467,In_81,In_623);
and U3468 (N_3468,In_1482,In_793);
xor U3469 (N_3469,In_1183,In_326);
or U3470 (N_3470,In_230,In_163);
or U3471 (N_3471,In_97,In_338);
or U3472 (N_3472,In_393,In_478);
and U3473 (N_3473,In_26,In_210);
nor U3474 (N_3474,In_507,In_1029);
and U3475 (N_3475,In_532,In_905);
nand U3476 (N_3476,In_387,In_1131);
nor U3477 (N_3477,In_953,In_545);
nand U3478 (N_3478,In_131,In_296);
or U3479 (N_3479,In_1202,In_406);
nor U3480 (N_3480,In_670,In_1404);
nand U3481 (N_3481,In_371,In_232);
and U3482 (N_3482,In_63,In_1005);
and U3483 (N_3483,In_553,In_1331);
xnor U3484 (N_3484,In_23,In_386);
nor U3485 (N_3485,In_1391,In_1073);
and U3486 (N_3486,In_464,In_1160);
and U3487 (N_3487,In_781,In_1481);
xor U3488 (N_3488,In_992,In_1366);
xnor U3489 (N_3489,In_448,In_531);
or U3490 (N_3490,In_951,In_318);
and U3491 (N_3491,In_49,In_683);
nor U3492 (N_3492,In_399,In_753);
nand U3493 (N_3493,In_1321,In_1061);
nor U3494 (N_3494,In_1146,In_580);
xnor U3495 (N_3495,In_1080,In_53);
and U3496 (N_3496,In_561,In_1478);
and U3497 (N_3497,In_1309,In_455);
nor U3498 (N_3498,In_838,In_370);
or U3499 (N_3499,In_914,In_1015);
or U3500 (N_3500,In_644,In_1338);
or U3501 (N_3501,In_1325,In_955);
nand U3502 (N_3502,In_537,In_1044);
nor U3503 (N_3503,In_1453,In_1339);
or U3504 (N_3504,In_799,In_101);
nand U3505 (N_3505,In_741,In_1481);
and U3506 (N_3506,In_949,In_0);
or U3507 (N_3507,In_1374,In_970);
nand U3508 (N_3508,In_1454,In_947);
and U3509 (N_3509,In_326,In_246);
xor U3510 (N_3510,In_1394,In_1367);
nor U3511 (N_3511,In_1134,In_1092);
nor U3512 (N_3512,In_565,In_164);
or U3513 (N_3513,In_976,In_816);
and U3514 (N_3514,In_790,In_1066);
xnor U3515 (N_3515,In_578,In_1052);
nor U3516 (N_3516,In_800,In_11);
nand U3517 (N_3517,In_1349,In_1384);
nand U3518 (N_3518,In_178,In_1273);
and U3519 (N_3519,In_1414,In_826);
or U3520 (N_3520,In_651,In_1258);
nand U3521 (N_3521,In_1113,In_1330);
nor U3522 (N_3522,In_1011,In_622);
xnor U3523 (N_3523,In_300,In_1382);
and U3524 (N_3524,In_344,In_414);
nor U3525 (N_3525,In_550,In_26);
nor U3526 (N_3526,In_1105,In_253);
and U3527 (N_3527,In_555,In_439);
nor U3528 (N_3528,In_560,In_24);
nand U3529 (N_3529,In_225,In_820);
nand U3530 (N_3530,In_308,In_1390);
or U3531 (N_3531,In_1289,In_538);
nor U3532 (N_3532,In_1250,In_1142);
and U3533 (N_3533,In_208,In_953);
or U3534 (N_3534,In_518,In_892);
nor U3535 (N_3535,In_862,In_590);
or U3536 (N_3536,In_942,In_852);
and U3537 (N_3537,In_365,In_1059);
nor U3538 (N_3538,In_1397,In_817);
or U3539 (N_3539,In_227,In_1041);
xnor U3540 (N_3540,In_832,In_1434);
xnor U3541 (N_3541,In_679,In_1496);
and U3542 (N_3542,In_892,In_385);
nor U3543 (N_3543,In_1218,In_826);
nand U3544 (N_3544,In_290,In_30);
or U3545 (N_3545,In_421,In_809);
nor U3546 (N_3546,In_28,In_1495);
or U3547 (N_3547,In_593,In_1457);
and U3548 (N_3548,In_411,In_80);
or U3549 (N_3549,In_1465,In_306);
nand U3550 (N_3550,In_333,In_561);
and U3551 (N_3551,In_1161,In_176);
and U3552 (N_3552,In_251,In_210);
xor U3553 (N_3553,In_1465,In_353);
or U3554 (N_3554,In_334,In_24);
or U3555 (N_3555,In_930,In_730);
and U3556 (N_3556,In_1344,In_689);
or U3557 (N_3557,In_750,In_365);
xnor U3558 (N_3558,In_104,In_1416);
and U3559 (N_3559,In_230,In_698);
or U3560 (N_3560,In_173,In_34);
or U3561 (N_3561,In_372,In_1005);
or U3562 (N_3562,In_164,In_897);
nand U3563 (N_3563,In_920,In_474);
and U3564 (N_3564,In_918,In_444);
and U3565 (N_3565,In_600,In_1268);
nor U3566 (N_3566,In_493,In_345);
xor U3567 (N_3567,In_1490,In_1433);
or U3568 (N_3568,In_1334,In_1271);
xor U3569 (N_3569,In_859,In_142);
nand U3570 (N_3570,In_629,In_1214);
xor U3571 (N_3571,In_646,In_459);
nand U3572 (N_3572,In_646,In_1340);
nand U3573 (N_3573,In_469,In_1006);
or U3574 (N_3574,In_819,In_639);
or U3575 (N_3575,In_970,In_565);
nor U3576 (N_3576,In_363,In_29);
xnor U3577 (N_3577,In_440,In_214);
nor U3578 (N_3578,In_317,In_715);
xnor U3579 (N_3579,In_301,In_613);
or U3580 (N_3580,In_1234,In_135);
or U3581 (N_3581,In_274,In_1441);
or U3582 (N_3582,In_140,In_959);
xor U3583 (N_3583,In_1450,In_671);
nand U3584 (N_3584,In_698,In_259);
nor U3585 (N_3585,In_111,In_1402);
nor U3586 (N_3586,In_597,In_863);
or U3587 (N_3587,In_769,In_113);
or U3588 (N_3588,In_574,In_1389);
nor U3589 (N_3589,In_1286,In_1217);
and U3590 (N_3590,In_296,In_760);
xnor U3591 (N_3591,In_999,In_1038);
and U3592 (N_3592,In_1035,In_79);
nor U3593 (N_3593,In_355,In_96);
nand U3594 (N_3594,In_333,In_107);
and U3595 (N_3595,In_358,In_674);
nand U3596 (N_3596,In_780,In_330);
or U3597 (N_3597,In_869,In_125);
xor U3598 (N_3598,In_797,In_47);
or U3599 (N_3599,In_1098,In_701);
nor U3600 (N_3600,In_192,In_689);
or U3601 (N_3601,In_1406,In_774);
xor U3602 (N_3602,In_1449,In_381);
nand U3603 (N_3603,In_545,In_471);
and U3604 (N_3604,In_105,In_1165);
xor U3605 (N_3605,In_616,In_551);
and U3606 (N_3606,In_459,In_1332);
xnor U3607 (N_3607,In_558,In_199);
or U3608 (N_3608,In_31,In_1059);
xnor U3609 (N_3609,In_845,In_263);
xnor U3610 (N_3610,In_1314,In_696);
nand U3611 (N_3611,In_470,In_630);
nor U3612 (N_3612,In_597,In_582);
nor U3613 (N_3613,In_1198,In_86);
xnor U3614 (N_3614,In_1100,In_573);
or U3615 (N_3615,In_664,In_386);
nor U3616 (N_3616,In_93,In_868);
xor U3617 (N_3617,In_492,In_284);
nand U3618 (N_3618,In_803,In_331);
nor U3619 (N_3619,In_1304,In_1);
or U3620 (N_3620,In_364,In_1344);
nand U3621 (N_3621,In_13,In_989);
nor U3622 (N_3622,In_866,In_600);
nor U3623 (N_3623,In_74,In_544);
xnor U3624 (N_3624,In_912,In_723);
nor U3625 (N_3625,In_542,In_1275);
nand U3626 (N_3626,In_1171,In_345);
nand U3627 (N_3627,In_982,In_336);
xnor U3628 (N_3628,In_1298,In_905);
and U3629 (N_3629,In_706,In_1011);
or U3630 (N_3630,In_782,In_728);
and U3631 (N_3631,In_329,In_992);
xor U3632 (N_3632,In_358,In_846);
or U3633 (N_3633,In_728,In_848);
or U3634 (N_3634,In_1288,In_1317);
and U3635 (N_3635,In_737,In_221);
nand U3636 (N_3636,In_341,In_1389);
and U3637 (N_3637,In_329,In_194);
xor U3638 (N_3638,In_620,In_851);
or U3639 (N_3639,In_1021,In_399);
nor U3640 (N_3640,In_685,In_208);
or U3641 (N_3641,In_595,In_1489);
and U3642 (N_3642,In_512,In_1029);
or U3643 (N_3643,In_921,In_1130);
nand U3644 (N_3644,In_138,In_807);
and U3645 (N_3645,In_1177,In_135);
nor U3646 (N_3646,In_274,In_735);
and U3647 (N_3647,In_563,In_50);
or U3648 (N_3648,In_1094,In_1029);
or U3649 (N_3649,In_940,In_767);
xnor U3650 (N_3650,In_1405,In_120);
or U3651 (N_3651,In_27,In_568);
xor U3652 (N_3652,In_700,In_333);
nand U3653 (N_3653,In_1158,In_1374);
or U3654 (N_3654,In_713,In_1365);
xor U3655 (N_3655,In_521,In_1480);
and U3656 (N_3656,In_312,In_1208);
nor U3657 (N_3657,In_812,In_240);
nand U3658 (N_3658,In_470,In_1368);
xor U3659 (N_3659,In_332,In_1087);
or U3660 (N_3660,In_113,In_210);
or U3661 (N_3661,In_1493,In_788);
or U3662 (N_3662,In_341,In_1198);
nand U3663 (N_3663,In_176,In_1393);
or U3664 (N_3664,In_1368,In_1041);
or U3665 (N_3665,In_447,In_698);
xnor U3666 (N_3666,In_960,In_467);
and U3667 (N_3667,In_1200,In_679);
nor U3668 (N_3668,In_603,In_508);
nor U3669 (N_3669,In_854,In_735);
nand U3670 (N_3670,In_1412,In_977);
xor U3671 (N_3671,In_373,In_920);
nor U3672 (N_3672,In_804,In_80);
nor U3673 (N_3673,In_18,In_171);
or U3674 (N_3674,In_944,In_217);
nand U3675 (N_3675,In_388,In_93);
nand U3676 (N_3676,In_459,In_1384);
and U3677 (N_3677,In_230,In_1183);
nor U3678 (N_3678,In_946,In_1065);
and U3679 (N_3679,In_1012,In_1349);
and U3680 (N_3680,In_128,In_500);
nand U3681 (N_3681,In_849,In_750);
nand U3682 (N_3682,In_1117,In_530);
xor U3683 (N_3683,In_767,In_659);
xnor U3684 (N_3684,In_1182,In_1249);
nand U3685 (N_3685,In_1110,In_1482);
xnor U3686 (N_3686,In_1127,In_191);
nor U3687 (N_3687,In_723,In_525);
or U3688 (N_3688,In_1238,In_1462);
nand U3689 (N_3689,In_378,In_678);
or U3690 (N_3690,In_89,In_780);
xor U3691 (N_3691,In_445,In_922);
nor U3692 (N_3692,In_840,In_1322);
or U3693 (N_3693,In_385,In_760);
xnor U3694 (N_3694,In_978,In_314);
nand U3695 (N_3695,In_1016,In_128);
nor U3696 (N_3696,In_978,In_477);
nand U3697 (N_3697,In_894,In_453);
xor U3698 (N_3698,In_181,In_870);
nand U3699 (N_3699,In_160,In_753);
nor U3700 (N_3700,In_363,In_1087);
nand U3701 (N_3701,In_375,In_1103);
or U3702 (N_3702,In_1302,In_972);
or U3703 (N_3703,In_173,In_1338);
or U3704 (N_3704,In_1341,In_1497);
nor U3705 (N_3705,In_1317,In_1401);
and U3706 (N_3706,In_192,In_13);
nor U3707 (N_3707,In_508,In_292);
nand U3708 (N_3708,In_200,In_383);
and U3709 (N_3709,In_881,In_1075);
xor U3710 (N_3710,In_1154,In_62);
xnor U3711 (N_3711,In_278,In_459);
nor U3712 (N_3712,In_1462,In_61);
nand U3713 (N_3713,In_842,In_944);
xnor U3714 (N_3714,In_733,In_694);
and U3715 (N_3715,In_733,In_1432);
nor U3716 (N_3716,In_129,In_734);
and U3717 (N_3717,In_41,In_960);
and U3718 (N_3718,In_75,In_769);
and U3719 (N_3719,In_68,In_1001);
and U3720 (N_3720,In_520,In_143);
and U3721 (N_3721,In_800,In_686);
nor U3722 (N_3722,In_1161,In_24);
and U3723 (N_3723,In_920,In_1498);
or U3724 (N_3724,In_922,In_276);
nor U3725 (N_3725,In_1044,In_317);
xor U3726 (N_3726,In_1452,In_318);
xor U3727 (N_3727,In_1177,In_185);
or U3728 (N_3728,In_212,In_1141);
nor U3729 (N_3729,In_1452,In_1492);
and U3730 (N_3730,In_1364,In_1446);
and U3731 (N_3731,In_749,In_941);
nand U3732 (N_3732,In_862,In_1435);
nand U3733 (N_3733,In_176,In_800);
or U3734 (N_3734,In_1275,In_1103);
nand U3735 (N_3735,In_157,In_371);
and U3736 (N_3736,In_1108,In_1252);
xnor U3737 (N_3737,In_1321,In_1290);
nor U3738 (N_3738,In_1083,In_734);
or U3739 (N_3739,In_1271,In_713);
and U3740 (N_3740,In_1334,In_554);
xnor U3741 (N_3741,In_617,In_906);
nand U3742 (N_3742,In_899,In_1133);
nor U3743 (N_3743,In_431,In_562);
nand U3744 (N_3744,In_1010,In_540);
xnor U3745 (N_3745,In_237,In_409);
nand U3746 (N_3746,In_213,In_293);
or U3747 (N_3747,In_1477,In_106);
nor U3748 (N_3748,In_133,In_1370);
or U3749 (N_3749,In_1130,In_489);
or U3750 (N_3750,In_1347,In_292);
or U3751 (N_3751,In_750,In_390);
xor U3752 (N_3752,In_293,In_1293);
nand U3753 (N_3753,In_1294,In_821);
nor U3754 (N_3754,In_269,In_824);
nor U3755 (N_3755,In_1363,In_725);
nand U3756 (N_3756,In_70,In_852);
or U3757 (N_3757,In_470,In_1096);
and U3758 (N_3758,In_1453,In_1257);
nor U3759 (N_3759,In_1134,In_512);
and U3760 (N_3760,In_477,In_779);
xor U3761 (N_3761,In_596,In_167);
nor U3762 (N_3762,In_1061,In_856);
xor U3763 (N_3763,In_1146,In_473);
or U3764 (N_3764,In_758,In_761);
or U3765 (N_3765,In_1020,In_792);
nand U3766 (N_3766,In_625,In_815);
xnor U3767 (N_3767,In_996,In_909);
or U3768 (N_3768,In_85,In_623);
and U3769 (N_3769,In_1341,In_1049);
or U3770 (N_3770,In_348,In_682);
and U3771 (N_3771,In_861,In_1492);
nand U3772 (N_3772,In_1339,In_1149);
xnor U3773 (N_3773,In_621,In_370);
and U3774 (N_3774,In_990,In_1482);
xor U3775 (N_3775,In_2,In_883);
nand U3776 (N_3776,In_427,In_717);
nor U3777 (N_3777,In_188,In_771);
nand U3778 (N_3778,In_360,In_806);
nand U3779 (N_3779,In_895,In_1183);
nor U3780 (N_3780,In_647,In_1458);
or U3781 (N_3781,In_151,In_1481);
and U3782 (N_3782,In_379,In_138);
nor U3783 (N_3783,In_1359,In_1034);
nand U3784 (N_3784,In_764,In_27);
and U3785 (N_3785,In_962,In_252);
xnor U3786 (N_3786,In_1154,In_146);
nor U3787 (N_3787,In_776,In_710);
nor U3788 (N_3788,In_160,In_1276);
xnor U3789 (N_3789,In_1069,In_1065);
nand U3790 (N_3790,In_1058,In_475);
nand U3791 (N_3791,In_876,In_748);
xor U3792 (N_3792,In_132,In_1355);
or U3793 (N_3793,In_686,In_1333);
nor U3794 (N_3794,In_769,In_67);
nand U3795 (N_3795,In_104,In_333);
and U3796 (N_3796,In_731,In_151);
nand U3797 (N_3797,In_1228,In_997);
or U3798 (N_3798,In_581,In_60);
nor U3799 (N_3799,In_1044,In_283);
or U3800 (N_3800,In_30,In_1177);
or U3801 (N_3801,In_1023,In_1217);
or U3802 (N_3802,In_665,In_492);
and U3803 (N_3803,In_454,In_89);
xor U3804 (N_3804,In_350,In_1308);
or U3805 (N_3805,In_436,In_220);
nand U3806 (N_3806,In_706,In_961);
xor U3807 (N_3807,In_1351,In_122);
or U3808 (N_3808,In_1115,In_1413);
and U3809 (N_3809,In_1277,In_1474);
xor U3810 (N_3810,In_1140,In_752);
xor U3811 (N_3811,In_829,In_507);
xor U3812 (N_3812,In_1411,In_1177);
nor U3813 (N_3813,In_346,In_800);
xor U3814 (N_3814,In_246,In_244);
nand U3815 (N_3815,In_18,In_472);
xnor U3816 (N_3816,In_614,In_1192);
and U3817 (N_3817,In_77,In_602);
nor U3818 (N_3818,In_1213,In_358);
nand U3819 (N_3819,In_705,In_50);
or U3820 (N_3820,In_663,In_278);
nor U3821 (N_3821,In_268,In_358);
and U3822 (N_3822,In_1416,In_947);
or U3823 (N_3823,In_106,In_197);
nor U3824 (N_3824,In_1076,In_1256);
xor U3825 (N_3825,In_747,In_491);
nand U3826 (N_3826,In_1399,In_488);
xor U3827 (N_3827,In_524,In_17);
or U3828 (N_3828,In_632,In_407);
nand U3829 (N_3829,In_126,In_1459);
nand U3830 (N_3830,In_425,In_824);
or U3831 (N_3831,In_251,In_466);
xor U3832 (N_3832,In_945,In_843);
nor U3833 (N_3833,In_338,In_1196);
nor U3834 (N_3834,In_1256,In_1177);
nand U3835 (N_3835,In_1497,In_265);
and U3836 (N_3836,In_1340,In_1210);
nor U3837 (N_3837,In_1260,In_1284);
nor U3838 (N_3838,In_202,In_1227);
xnor U3839 (N_3839,In_237,In_168);
or U3840 (N_3840,In_242,In_607);
and U3841 (N_3841,In_639,In_1381);
nand U3842 (N_3842,In_670,In_492);
and U3843 (N_3843,In_517,In_1137);
xor U3844 (N_3844,In_369,In_984);
and U3845 (N_3845,In_235,In_813);
nand U3846 (N_3846,In_1234,In_1106);
nor U3847 (N_3847,In_384,In_978);
nand U3848 (N_3848,In_1,In_1453);
xor U3849 (N_3849,In_530,In_33);
xnor U3850 (N_3850,In_552,In_1182);
and U3851 (N_3851,In_586,In_232);
and U3852 (N_3852,In_1440,In_790);
and U3853 (N_3853,In_753,In_977);
nand U3854 (N_3854,In_991,In_501);
nor U3855 (N_3855,In_1011,In_1236);
nand U3856 (N_3856,In_122,In_743);
nor U3857 (N_3857,In_330,In_25);
nor U3858 (N_3858,In_1230,In_385);
xor U3859 (N_3859,In_1379,In_3);
xor U3860 (N_3860,In_611,In_715);
nand U3861 (N_3861,In_921,In_479);
nor U3862 (N_3862,In_1429,In_629);
nor U3863 (N_3863,In_1151,In_882);
nor U3864 (N_3864,In_945,In_1476);
and U3865 (N_3865,In_152,In_676);
or U3866 (N_3866,In_1112,In_1301);
xor U3867 (N_3867,In_607,In_685);
nor U3868 (N_3868,In_662,In_1045);
or U3869 (N_3869,In_422,In_925);
or U3870 (N_3870,In_386,In_991);
xnor U3871 (N_3871,In_1144,In_326);
nand U3872 (N_3872,In_1439,In_414);
nor U3873 (N_3873,In_1271,In_688);
or U3874 (N_3874,In_1041,In_303);
nor U3875 (N_3875,In_1107,In_1419);
or U3876 (N_3876,In_1190,In_659);
nand U3877 (N_3877,In_442,In_1465);
nand U3878 (N_3878,In_933,In_325);
and U3879 (N_3879,In_373,In_325);
nor U3880 (N_3880,In_1150,In_284);
xor U3881 (N_3881,In_851,In_1123);
nand U3882 (N_3882,In_504,In_313);
nor U3883 (N_3883,In_69,In_1226);
and U3884 (N_3884,In_539,In_1158);
or U3885 (N_3885,In_1175,In_1216);
nand U3886 (N_3886,In_707,In_1085);
nand U3887 (N_3887,In_911,In_597);
xor U3888 (N_3888,In_117,In_1285);
and U3889 (N_3889,In_430,In_740);
and U3890 (N_3890,In_839,In_560);
xnor U3891 (N_3891,In_1352,In_959);
or U3892 (N_3892,In_1174,In_186);
nand U3893 (N_3893,In_1065,In_1387);
nor U3894 (N_3894,In_996,In_677);
and U3895 (N_3895,In_666,In_985);
or U3896 (N_3896,In_1289,In_1249);
xnor U3897 (N_3897,In_984,In_158);
and U3898 (N_3898,In_1130,In_1239);
xnor U3899 (N_3899,In_1280,In_1213);
and U3900 (N_3900,In_1230,In_748);
nand U3901 (N_3901,In_146,In_439);
or U3902 (N_3902,In_859,In_538);
nor U3903 (N_3903,In_906,In_1128);
and U3904 (N_3904,In_1373,In_412);
xnor U3905 (N_3905,In_92,In_949);
or U3906 (N_3906,In_304,In_54);
nand U3907 (N_3907,In_1174,In_1483);
or U3908 (N_3908,In_1181,In_58);
xnor U3909 (N_3909,In_957,In_682);
or U3910 (N_3910,In_1374,In_713);
and U3911 (N_3911,In_290,In_115);
xor U3912 (N_3912,In_356,In_1461);
nand U3913 (N_3913,In_582,In_913);
or U3914 (N_3914,In_740,In_273);
nor U3915 (N_3915,In_988,In_568);
xor U3916 (N_3916,In_115,In_582);
nand U3917 (N_3917,In_1424,In_960);
xor U3918 (N_3918,In_1310,In_1164);
nor U3919 (N_3919,In_1245,In_961);
or U3920 (N_3920,In_670,In_260);
nor U3921 (N_3921,In_381,In_281);
or U3922 (N_3922,In_312,In_1146);
nand U3923 (N_3923,In_850,In_149);
nor U3924 (N_3924,In_252,In_384);
xnor U3925 (N_3925,In_779,In_36);
and U3926 (N_3926,In_766,In_1017);
and U3927 (N_3927,In_833,In_983);
nor U3928 (N_3928,In_768,In_1470);
xnor U3929 (N_3929,In_627,In_903);
or U3930 (N_3930,In_1176,In_244);
xnor U3931 (N_3931,In_449,In_939);
nor U3932 (N_3932,In_519,In_368);
nand U3933 (N_3933,In_1171,In_303);
nand U3934 (N_3934,In_453,In_669);
or U3935 (N_3935,In_435,In_37);
xor U3936 (N_3936,In_1212,In_283);
or U3937 (N_3937,In_1078,In_690);
or U3938 (N_3938,In_281,In_695);
and U3939 (N_3939,In_1474,In_924);
nor U3940 (N_3940,In_286,In_1079);
nand U3941 (N_3941,In_1415,In_1445);
and U3942 (N_3942,In_980,In_1018);
nor U3943 (N_3943,In_1209,In_1136);
xor U3944 (N_3944,In_846,In_558);
nor U3945 (N_3945,In_5,In_1394);
nor U3946 (N_3946,In_1368,In_1455);
nor U3947 (N_3947,In_1445,In_487);
xnor U3948 (N_3948,In_687,In_722);
or U3949 (N_3949,In_215,In_1007);
and U3950 (N_3950,In_233,In_1299);
nand U3951 (N_3951,In_772,In_1462);
nor U3952 (N_3952,In_777,In_1228);
nor U3953 (N_3953,In_146,In_1350);
and U3954 (N_3954,In_1291,In_1475);
and U3955 (N_3955,In_1307,In_949);
or U3956 (N_3956,In_1289,In_756);
nor U3957 (N_3957,In_1299,In_1456);
xor U3958 (N_3958,In_95,In_730);
nand U3959 (N_3959,In_715,In_789);
or U3960 (N_3960,In_37,In_1419);
and U3961 (N_3961,In_395,In_227);
nand U3962 (N_3962,In_1494,In_758);
xnor U3963 (N_3963,In_1154,In_1117);
nor U3964 (N_3964,In_547,In_638);
or U3965 (N_3965,In_548,In_1410);
and U3966 (N_3966,In_137,In_1142);
or U3967 (N_3967,In_1067,In_768);
xor U3968 (N_3968,In_1208,In_928);
xnor U3969 (N_3969,In_1422,In_154);
and U3970 (N_3970,In_477,In_1276);
or U3971 (N_3971,In_1110,In_742);
and U3972 (N_3972,In_697,In_740);
or U3973 (N_3973,In_332,In_734);
nor U3974 (N_3974,In_926,In_197);
and U3975 (N_3975,In_798,In_136);
nor U3976 (N_3976,In_1082,In_810);
nor U3977 (N_3977,In_759,In_1135);
nand U3978 (N_3978,In_921,In_938);
xor U3979 (N_3979,In_331,In_615);
xnor U3980 (N_3980,In_88,In_553);
nand U3981 (N_3981,In_935,In_556);
nor U3982 (N_3982,In_125,In_507);
nor U3983 (N_3983,In_493,In_497);
xor U3984 (N_3984,In_154,In_286);
and U3985 (N_3985,In_634,In_799);
or U3986 (N_3986,In_29,In_1272);
or U3987 (N_3987,In_1177,In_1484);
nor U3988 (N_3988,In_662,In_133);
nor U3989 (N_3989,In_730,In_993);
nor U3990 (N_3990,In_128,In_734);
nor U3991 (N_3991,In_781,In_750);
xor U3992 (N_3992,In_423,In_483);
or U3993 (N_3993,In_791,In_496);
or U3994 (N_3994,In_1341,In_111);
or U3995 (N_3995,In_787,In_304);
xor U3996 (N_3996,In_417,In_518);
nand U3997 (N_3997,In_343,In_700);
and U3998 (N_3998,In_278,In_556);
xor U3999 (N_3999,In_339,In_1356);
or U4000 (N_4000,In_1008,In_291);
nor U4001 (N_4001,In_184,In_39);
nor U4002 (N_4002,In_1361,In_949);
xnor U4003 (N_4003,In_814,In_1363);
nor U4004 (N_4004,In_1420,In_308);
and U4005 (N_4005,In_1493,In_579);
nand U4006 (N_4006,In_1065,In_461);
and U4007 (N_4007,In_1041,In_859);
nand U4008 (N_4008,In_27,In_101);
xor U4009 (N_4009,In_151,In_883);
xor U4010 (N_4010,In_285,In_417);
nor U4011 (N_4011,In_991,In_778);
nand U4012 (N_4012,In_874,In_827);
nor U4013 (N_4013,In_53,In_1372);
and U4014 (N_4014,In_1376,In_209);
xor U4015 (N_4015,In_388,In_611);
xor U4016 (N_4016,In_1283,In_1354);
nor U4017 (N_4017,In_125,In_1134);
and U4018 (N_4018,In_1357,In_632);
nand U4019 (N_4019,In_621,In_1489);
nor U4020 (N_4020,In_1346,In_1005);
and U4021 (N_4021,In_1040,In_508);
or U4022 (N_4022,In_283,In_202);
nor U4023 (N_4023,In_939,In_959);
or U4024 (N_4024,In_185,In_243);
nand U4025 (N_4025,In_1075,In_1053);
and U4026 (N_4026,In_983,In_1437);
nor U4027 (N_4027,In_892,In_1420);
xnor U4028 (N_4028,In_1074,In_764);
nor U4029 (N_4029,In_1404,In_1355);
and U4030 (N_4030,In_297,In_679);
or U4031 (N_4031,In_76,In_565);
nand U4032 (N_4032,In_1312,In_125);
nand U4033 (N_4033,In_765,In_1229);
or U4034 (N_4034,In_959,In_446);
nand U4035 (N_4035,In_1315,In_469);
nor U4036 (N_4036,In_1398,In_129);
nor U4037 (N_4037,In_382,In_570);
and U4038 (N_4038,In_702,In_517);
or U4039 (N_4039,In_1295,In_1122);
nor U4040 (N_4040,In_319,In_637);
nand U4041 (N_4041,In_351,In_330);
nand U4042 (N_4042,In_691,In_1483);
nand U4043 (N_4043,In_1297,In_1203);
xnor U4044 (N_4044,In_397,In_302);
or U4045 (N_4045,In_445,In_464);
nor U4046 (N_4046,In_1111,In_866);
nor U4047 (N_4047,In_1340,In_886);
xnor U4048 (N_4048,In_350,In_369);
nand U4049 (N_4049,In_321,In_879);
or U4050 (N_4050,In_408,In_1370);
xnor U4051 (N_4051,In_318,In_478);
xor U4052 (N_4052,In_13,In_1151);
and U4053 (N_4053,In_1361,In_687);
and U4054 (N_4054,In_275,In_132);
xor U4055 (N_4055,In_387,In_1162);
nand U4056 (N_4056,In_317,In_1192);
xnor U4057 (N_4057,In_183,In_442);
or U4058 (N_4058,In_736,In_1004);
nor U4059 (N_4059,In_82,In_1139);
or U4060 (N_4060,In_477,In_442);
or U4061 (N_4061,In_440,In_412);
and U4062 (N_4062,In_305,In_150);
nand U4063 (N_4063,In_1141,In_1192);
and U4064 (N_4064,In_759,In_1008);
or U4065 (N_4065,In_1318,In_35);
or U4066 (N_4066,In_654,In_134);
nand U4067 (N_4067,In_1102,In_980);
nor U4068 (N_4068,In_1312,In_554);
or U4069 (N_4069,In_279,In_902);
nor U4070 (N_4070,In_504,In_861);
and U4071 (N_4071,In_749,In_680);
nor U4072 (N_4072,In_270,In_1099);
nor U4073 (N_4073,In_1449,In_1213);
nor U4074 (N_4074,In_172,In_413);
nand U4075 (N_4075,In_327,In_391);
xnor U4076 (N_4076,In_747,In_435);
and U4077 (N_4077,In_569,In_492);
nor U4078 (N_4078,In_166,In_88);
xnor U4079 (N_4079,In_365,In_906);
xor U4080 (N_4080,In_813,In_1439);
and U4081 (N_4081,In_40,In_791);
xnor U4082 (N_4082,In_70,In_1223);
or U4083 (N_4083,In_840,In_811);
nand U4084 (N_4084,In_469,In_94);
or U4085 (N_4085,In_679,In_594);
xnor U4086 (N_4086,In_1050,In_5);
nand U4087 (N_4087,In_1138,In_399);
nor U4088 (N_4088,In_388,In_874);
nor U4089 (N_4089,In_624,In_802);
or U4090 (N_4090,In_394,In_278);
nor U4091 (N_4091,In_445,In_1158);
nor U4092 (N_4092,In_815,In_975);
xnor U4093 (N_4093,In_399,In_1159);
or U4094 (N_4094,In_1185,In_857);
nand U4095 (N_4095,In_983,In_214);
and U4096 (N_4096,In_187,In_529);
nor U4097 (N_4097,In_145,In_1219);
or U4098 (N_4098,In_385,In_94);
xnor U4099 (N_4099,In_748,In_1424);
or U4100 (N_4100,In_1480,In_372);
and U4101 (N_4101,In_826,In_186);
nand U4102 (N_4102,In_923,In_1097);
or U4103 (N_4103,In_1131,In_230);
nor U4104 (N_4104,In_1137,In_588);
nor U4105 (N_4105,In_984,In_17);
or U4106 (N_4106,In_972,In_1173);
nand U4107 (N_4107,In_666,In_538);
xnor U4108 (N_4108,In_1143,In_586);
nor U4109 (N_4109,In_1164,In_119);
and U4110 (N_4110,In_1272,In_1025);
nor U4111 (N_4111,In_418,In_296);
xor U4112 (N_4112,In_634,In_1255);
or U4113 (N_4113,In_114,In_1377);
nor U4114 (N_4114,In_667,In_104);
or U4115 (N_4115,In_1472,In_888);
nor U4116 (N_4116,In_524,In_514);
and U4117 (N_4117,In_445,In_747);
or U4118 (N_4118,In_1402,In_1110);
xor U4119 (N_4119,In_986,In_508);
nor U4120 (N_4120,In_774,In_885);
nand U4121 (N_4121,In_822,In_275);
and U4122 (N_4122,In_835,In_1314);
nor U4123 (N_4123,In_767,In_1228);
nand U4124 (N_4124,In_834,In_824);
or U4125 (N_4125,In_610,In_1446);
or U4126 (N_4126,In_1292,In_593);
xor U4127 (N_4127,In_1164,In_233);
nand U4128 (N_4128,In_1093,In_430);
and U4129 (N_4129,In_1468,In_100);
and U4130 (N_4130,In_741,In_34);
nor U4131 (N_4131,In_1088,In_995);
nand U4132 (N_4132,In_311,In_231);
and U4133 (N_4133,In_1113,In_1261);
xor U4134 (N_4134,In_114,In_343);
or U4135 (N_4135,In_853,In_1247);
nand U4136 (N_4136,In_1482,In_164);
or U4137 (N_4137,In_1013,In_77);
or U4138 (N_4138,In_452,In_391);
nor U4139 (N_4139,In_634,In_939);
nand U4140 (N_4140,In_1438,In_864);
and U4141 (N_4141,In_388,In_153);
nor U4142 (N_4142,In_1269,In_1450);
nor U4143 (N_4143,In_1229,In_1268);
or U4144 (N_4144,In_793,In_523);
or U4145 (N_4145,In_564,In_1141);
nor U4146 (N_4146,In_134,In_67);
or U4147 (N_4147,In_422,In_728);
nor U4148 (N_4148,In_956,In_476);
and U4149 (N_4149,In_1452,In_918);
or U4150 (N_4150,In_476,In_486);
or U4151 (N_4151,In_947,In_1385);
and U4152 (N_4152,In_766,In_981);
nand U4153 (N_4153,In_929,In_884);
and U4154 (N_4154,In_377,In_159);
nand U4155 (N_4155,In_1033,In_1343);
xor U4156 (N_4156,In_1436,In_280);
xnor U4157 (N_4157,In_902,In_458);
and U4158 (N_4158,In_480,In_83);
xor U4159 (N_4159,In_38,In_855);
or U4160 (N_4160,In_4,In_12);
or U4161 (N_4161,In_844,In_285);
nand U4162 (N_4162,In_430,In_16);
and U4163 (N_4163,In_700,In_1236);
and U4164 (N_4164,In_6,In_793);
nor U4165 (N_4165,In_314,In_68);
xor U4166 (N_4166,In_534,In_1376);
xor U4167 (N_4167,In_756,In_901);
nand U4168 (N_4168,In_756,In_1176);
xnor U4169 (N_4169,In_885,In_767);
xnor U4170 (N_4170,In_413,In_1003);
and U4171 (N_4171,In_586,In_171);
xnor U4172 (N_4172,In_1272,In_789);
and U4173 (N_4173,In_607,In_646);
nand U4174 (N_4174,In_673,In_15);
nand U4175 (N_4175,In_1227,In_1465);
xor U4176 (N_4176,In_505,In_1021);
xnor U4177 (N_4177,In_1082,In_1275);
and U4178 (N_4178,In_1083,In_504);
nand U4179 (N_4179,In_1422,In_988);
xnor U4180 (N_4180,In_1389,In_203);
or U4181 (N_4181,In_788,In_1067);
nand U4182 (N_4182,In_451,In_1268);
or U4183 (N_4183,In_1037,In_1462);
nand U4184 (N_4184,In_1323,In_1430);
and U4185 (N_4185,In_255,In_272);
xor U4186 (N_4186,In_1124,In_1070);
nand U4187 (N_4187,In_1283,In_1144);
nor U4188 (N_4188,In_1441,In_94);
nor U4189 (N_4189,In_49,In_959);
nand U4190 (N_4190,In_310,In_682);
or U4191 (N_4191,In_1164,In_914);
or U4192 (N_4192,In_755,In_1334);
and U4193 (N_4193,In_613,In_1252);
xnor U4194 (N_4194,In_1408,In_1312);
or U4195 (N_4195,In_399,In_754);
and U4196 (N_4196,In_1385,In_1426);
nor U4197 (N_4197,In_266,In_614);
xnor U4198 (N_4198,In_1221,In_1101);
or U4199 (N_4199,In_1482,In_344);
or U4200 (N_4200,In_771,In_1303);
nand U4201 (N_4201,In_1358,In_1079);
and U4202 (N_4202,In_223,In_710);
xor U4203 (N_4203,In_627,In_187);
xnor U4204 (N_4204,In_855,In_553);
xnor U4205 (N_4205,In_932,In_742);
nand U4206 (N_4206,In_1453,In_503);
and U4207 (N_4207,In_1117,In_524);
and U4208 (N_4208,In_206,In_116);
or U4209 (N_4209,In_1010,In_436);
nand U4210 (N_4210,In_1029,In_330);
xor U4211 (N_4211,In_413,In_1005);
or U4212 (N_4212,In_1090,In_1338);
xnor U4213 (N_4213,In_287,In_440);
and U4214 (N_4214,In_1247,In_1086);
xnor U4215 (N_4215,In_107,In_72);
nor U4216 (N_4216,In_1466,In_692);
nand U4217 (N_4217,In_433,In_1283);
nor U4218 (N_4218,In_859,In_517);
nor U4219 (N_4219,In_830,In_306);
and U4220 (N_4220,In_1153,In_1498);
xor U4221 (N_4221,In_245,In_1391);
and U4222 (N_4222,In_1069,In_315);
nor U4223 (N_4223,In_472,In_42);
or U4224 (N_4224,In_111,In_108);
nand U4225 (N_4225,In_946,In_1317);
nor U4226 (N_4226,In_748,In_145);
and U4227 (N_4227,In_500,In_690);
or U4228 (N_4228,In_814,In_46);
and U4229 (N_4229,In_1031,In_967);
xnor U4230 (N_4230,In_1283,In_1418);
nand U4231 (N_4231,In_1258,In_1379);
and U4232 (N_4232,In_363,In_452);
xnor U4233 (N_4233,In_1130,In_162);
xnor U4234 (N_4234,In_132,In_795);
or U4235 (N_4235,In_179,In_1238);
nor U4236 (N_4236,In_850,In_1305);
xor U4237 (N_4237,In_1131,In_16);
xor U4238 (N_4238,In_575,In_169);
nor U4239 (N_4239,In_600,In_1098);
xor U4240 (N_4240,In_96,In_644);
or U4241 (N_4241,In_141,In_1352);
nor U4242 (N_4242,In_1394,In_1222);
nand U4243 (N_4243,In_31,In_529);
xor U4244 (N_4244,In_860,In_1368);
xnor U4245 (N_4245,In_239,In_0);
nor U4246 (N_4246,In_760,In_579);
and U4247 (N_4247,In_746,In_476);
xor U4248 (N_4248,In_193,In_1180);
nand U4249 (N_4249,In_609,In_1101);
nand U4250 (N_4250,In_53,In_219);
and U4251 (N_4251,In_1292,In_616);
and U4252 (N_4252,In_35,In_387);
or U4253 (N_4253,In_579,In_584);
or U4254 (N_4254,In_1425,In_1483);
nand U4255 (N_4255,In_1089,In_1458);
xor U4256 (N_4256,In_1284,In_647);
nor U4257 (N_4257,In_203,In_1393);
nand U4258 (N_4258,In_710,In_133);
nand U4259 (N_4259,In_32,In_226);
and U4260 (N_4260,In_1232,In_933);
or U4261 (N_4261,In_183,In_371);
xor U4262 (N_4262,In_706,In_1084);
nor U4263 (N_4263,In_246,In_742);
or U4264 (N_4264,In_489,In_1495);
and U4265 (N_4265,In_385,In_344);
and U4266 (N_4266,In_458,In_717);
nor U4267 (N_4267,In_659,In_68);
and U4268 (N_4268,In_1017,In_793);
or U4269 (N_4269,In_897,In_776);
nor U4270 (N_4270,In_355,In_517);
or U4271 (N_4271,In_1240,In_773);
and U4272 (N_4272,In_1202,In_1026);
or U4273 (N_4273,In_702,In_1195);
or U4274 (N_4274,In_1396,In_137);
nand U4275 (N_4275,In_673,In_559);
and U4276 (N_4276,In_1473,In_922);
nor U4277 (N_4277,In_489,In_851);
or U4278 (N_4278,In_604,In_575);
nor U4279 (N_4279,In_106,In_639);
xnor U4280 (N_4280,In_1267,In_214);
xor U4281 (N_4281,In_307,In_904);
and U4282 (N_4282,In_1137,In_79);
xor U4283 (N_4283,In_1464,In_440);
and U4284 (N_4284,In_1189,In_286);
xnor U4285 (N_4285,In_1347,In_1091);
and U4286 (N_4286,In_377,In_610);
and U4287 (N_4287,In_127,In_887);
nand U4288 (N_4288,In_576,In_1139);
xnor U4289 (N_4289,In_166,In_1464);
and U4290 (N_4290,In_1263,In_197);
or U4291 (N_4291,In_997,In_929);
and U4292 (N_4292,In_1217,In_1099);
nor U4293 (N_4293,In_1333,In_1472);
xor U4294 (N_4294,In_1019,In_1454);
xor U4295 (N_4295,In_1065,In_1179);
or U4296 (N_4296,In_1073,In_704);
and U4297 (N_4297,In_37,In_48);
nand U4298 (N_4298,In_354,In_589);
and U4299 (N_4299,In_526,In_420);
and U4300 (N_4300,In_1484,In_1181);
and U4301 (N_4301,In_71,In_571);
and U4302 (N_4302,In_676,In_997);
xnor U4303 (N_4303,In_187,In_513);
xor U4304 (N_4304,In_1130,In_447);
or U4305 (N_4305,In_515,In_1333);
nand U4306 (N_4306,In_219,In_895);
and U4307 (N_4307,In_968,In_1270);
and U4308 (N_4308,In_331,In_1036);
nand U4309 (N_4309,In_934,In_1434);
or U4310 (N_4310,In_1052,In_1279);
xnor U4311 (N_4311,In_522,In_35);
nor U4312 (N_4312,In_1065,In_562);
or U4313 (N_4313,In_275,In_340);
and U4314 (N_4314,In_254,In_372);
or U4315 (N_4315,In_636,In_275);
nor U4316 (N_4316,In_379,In_381);
xnor U4317 (N_4317,In_795,In_698);
nand U4318 (N_4318,In_1278,In_1478);
nor U4319 (N_4319,In_1455,In_1199);
and U4320 (N_4320,In_1287,In_1492);
and U4321 (N_4321,In_1270,In_91);
xor U4322 (N_4322,In_1317,In_232);
xnor U4323 (N_4323,In_990,In_963);
xor U4324 (N_4324,In_80,In_864);
or U4325 (N_4325,In_95,In_608);
or U4326 (N_4326,In_663,In_1090);
nor U4327 (N_4327,In_460,In_1168);
xnor U4328 (N_4328,In_1186,In_1179);
xor U4329 (N_4329,In_578,In_312);
nand U4330 (N_4330,In_1145,In_312);
nor U4331 (N_4331,In_1334,In_937);
xnor U4332 (N_4332,In_1155,In_123);
nor U4333 (N_4333,In_866,In_869);
xor U4334 (N_4334,In_340,In_415);
xnor U4335 (N_4335,In_166,In_1322);
xnor U4336 (N_4336,In_1334,In_367);
xor U4337 (N_4337,In_1364,In_135);
or U4338 (N_4338,In_1191,In_1419);
and U4339 (N_4339,In_320,In_738);
xor U4340 (N_4340,In_31,In_221);
and U4341 (N_4341,In_63,In_960);
nor U4342 (N_4342,In_359,In_21);
nor U4343 (N_4343,In_893,In_399);
or U4344 (N_4344,In_959,In_438);
or U4345 (N_4345,In_1471,In_750);
or U4346 (N_4346,In_1059,In_497);
xnor U4347 (N_4347,In_753,In_806);
nor U4348 (N_4348,In_3,In_1385);
nor U4349 (N_4349,In_502,In_691);
nand U4350 (N_4350,In_484,In_793);
xnor U4351 (N_4351,In_879,In_1188);
nand U4352 (N_4352,In_1221,In_171);
nor U4353 (N_4353,In_347,In_1079);
xor U4354 (N_4354,In_432,In_1429);
or U4355 (N_4355,In_1379,In_544);
xnor U4356 (N_4356,In_1042,In_1389);
xor U4357 (N_4357,In_120,In_1209);
nor U4358 (N_4358,In_616,In_375);
xnor U4359 (N_4359,In_1482,In_723);
or U4360 (N_4360,In_497,In_966);
nor U4361 (N_4361,In_1379,In_941);
xnor U4362 (N_4362,In_1309,In_467);
nor U4363 (N_4363,In_554,In_232);
or U4364 (N_4364,In_843,In_381);
and U4365 (N_4365,In_1271,In_435);
nand U4366 (N_4366,In_603,In_561);
xnor U4367 (N_4367,In_637,In_226);
nor U4368 (N_4368,In_7,In_323);
and U4369 (N_4369,In_1034,In_750);
nand U4370 (N_4370,In_263,In_247);
or U4371 (N_4371,In_59,In_797);
nand U4372 (N_4372,In_997,In_1087);
nand U4373 (N_4373,In_1204,In_831);
nor U4374 (N_4374,In_419,In_802);
or U4375 (N_4375,In_1157,In_963);
nand U4376 (N_4376,In_162,In_384);
xnor U4377 (N_4377,In_625,In_1273);
and U4378 (N_4378,In_565,In_1341);
or U4379 (N_4379,In_203,In_370);
or U4380 (N_4380,In_522,In_1112);
nor U4381 (N_4381,In_434,In_410);
nand U4382 (N_4382,In_925,In_913);
nand U4383 (N_4383,In_614,In_48);
nor U4384 (N_4384,In_329,In_351);
xor U4385 (N_4385,In_213,In_6);
and U4386 (N_4386,In_620,In_1379);
or U4387 (N_4387,In_1121,In_1213);
xor U4388 (N_4388,In_1074,In_439);
xor U4389 (N_4389,In_1211,In_786);
nor U4390 (N_4390,In_560,In_996);
or U4391 (N_4391,In_1116,In_293);
xor U4392 (N_4392,In_755,In_936);
xnor U4393 (N_4393,In_1234,In_1403);
xnor U4394 (N_4394,In_754,In_115);
and U4395 (N_4395,In_450,In_1357);
nand U4396 (N_4396,In_726,In_58);
or U4397 (N_4397,In_965,In_428);
nor U4398 (N_4398,In_94,In_161);
nand U4399 (N_4399,In_1430,In_1253);
or U4400 (N_4400,In_385,In_839);
and U4401 (N_4401,In_397,In_1181);
and U4402 (N_4402,In_435,In_1391);
or U4403 (N_4403,In_116,In_1106);
nand U4404 (N_4404,In_967,In_1115);
nand U4405 (N_4405,In_617,In_27);
and U4406 (N_4406,In_809,In_217);
or U4407 (N_4407,In_1138,In_571);
nor U4408 (N_4408,In_654,In_1218);
xnor U4409 (N_4409,In_1082,In_1099);
and U4410 (N_4410,In_967,In_1103);
xor U4411 (N_4411,In_1247,In_1331);
nor U4412 (N_4412,In_1045,In_654);
or U4413 (N_4413,In_172,In_883);
or U4414 (N_4414,In_644,In_1033);
and U4415 (N_4415,In_857,In_193);
xor U4416 (N_4416,In_1004,In_107);
nor U4417 (N_4417,In_532,In_486);
xnor U4418 (N_4418,In_958,In_1125);
xnor U4419 (N_4419,In_649,In_511);
nor U4420 (N_4420,In_443,In_369);
nor U4421 (N_4421,In_1059,In_1305);
nand U4422 (N_4422,In_62,In_926);
and U4423 (N_4423,In_118,In_160);
nand U4424 (N_4424,In_1008,In_302);
nand U4425 (N_4425,In_1143,In_1460);
nor U4426 (N_4426,In_1267,In_1427);
and U4427 (N_4427,In_1025,In_977);
nand U4428 (N_4428,In_241,In_152);
or U4429 (N_4429,In_655,In_435);
nand U4430 (N_4430,In_1474,In_108);
nor U4431 (N_4431,In_1018,In_1456);
xnor U4432 (N_4432,In_209,In_485);
xor U4433 (N_4433,In_1437,In_891);
and U4434 (N_4434,In_343,In_954);
nand U4435 (N_4435,In_989,In_585);
and U4436 (N_4436,In_101,In_1437);
xnor U4437 (N_4437,In_1423,In_1217);
nor U4438 (N_4438,In_619,In_484);
nand U4439 (N_4439,In_786,In_199);
and U4440 (N_4440,In_725,In_528);
and U4441 (N_4441,In_91,In_1256);
and U4442 (N_4442,In_783,In_221);
or U4443 (N_4443,In_780,In_619);
or U4444 (N_4444,In_644,In_990);
or U4445 (N_4445,In_405,In_456);
or U4446 (N_4446,In_531,In_1335);
and U4447 (N_4447,In_101,In_974);
nor U4448 (N_4448,In_1484,In_877);
xor U4449 (N_4449,In_966,In_306);
and U4450 (N_4450,In_406,In_18);
or U4451 (N_4451,In_1496,In_403);
nand U4452 (N_4452,In_350,In_1072);
nor U4453 (N_4453,In_487,In_894);
and U4454 (N_4454,In_711,In_324);
or U4455 (N_4455,In_435,In_101);
nor U4456 (N_4456,In_415,In_884);
and U4457 (N_4457,In_1295,In_637);
xor U4458 (N_4458,In_431,In_1283);
nand U4459 (N_4459,In_655,In_718);
xnor U4460 (N_4460,In_1308,In_1383);
and U4461 (N_4461,In_656,In_274);
or U4462 (N_4462,In_877,In_1088);
or U4463 (N_4463,In_824,In_759);
or U4464 (N_4464,In_296,In_339);
and U4465 (N_4465,In_1226,In_423);
nand U4466 (N_4466,In_818,In_369);
xor U4467 (N_4467,In_166,In_1483);
nor U4468 (N_4468,In_533,In_852);
nand U4469 (N_4469,In_488,In_750);
and U4470 (N_4470,In_267,In_1371);
and U4471 (N_4471,In_1421,In_814);
nand U4472 (N_4472,In_1486,In_567);
xor U4473 (N_4473,In_818,In_605);
nand U4474 (N_4474,In_944,In_194);
nor U4475 (N_4475,In_1140,In_101);
nor U4476 (N_4476,In_444,In_983);
and U4477 (N_4477,In_151,In_1318);
nor U4478 (N_4478,In_1039,In_480);
xor U4479 (N_4479,In_69,In_1189);
or U4480 (N_4480,In_1449,In_746);
xnor U4481 (N_4481,In_63,In_91);
and U4482 (N_4482,In_1499,In_940);
nor U4483 (N_4483,In_235,In_884);
nor U4484 (N_4484,In_352,In_185);
xnor U4485 (N_4485,In_1358,In_650);
nor U4486 (N_4486,In_1088,In_88);
nor U4487 (N_4487,In_213,In_803);
nor U4488 (N_4488,In_471,In_1149);
nor U4489 (N_4489,In_9,In_531);
and U4490 (N_4490,In_60,In_790);
nor U4491 (N_4491,In_1424,In_1305);
xnor U4492 (N_4492,In_443,In_67);
xor U4493 (N_4493,In_883,In_881);
nand U4494 (N_4494,In_547,In_625);
nand U4495 (N_4495,In_526,In_123);
or U4496 (N_4496,In_976,In_649);
xnor U4497 (N_4497,In_1087,In_1050);
or U4498 (N_4498,In_1276,In_9);
xnor U4499 (N_4499,In_282,In_228);
and U4500 (N_4500,In_653,In_585);
or U4501 (N_4501,In_17,In_604);
nor U4502 (N_4502,In_1348,In_1047);
nor U4503 (N_4503,In_645,In_993);
nor U4504 (N_4504,In_1400,In_857);
xor U4505 (N_4505,In_587,In_985);
or U4506 (N_4506,In_503,In_466);
nor U4507 (N_4507,In_812,In_1480);
and U4508 (N_4508,In_1114,In_134);
and U4509 (N_4509,In_214,In_865);
nor U4510 (N_4510,In_800,In_738);
xnor U4511 (N_4511,In_1295,In_606);
nand U4512 (N_4512,In_126,In_1085);
nand U4513 (N_4513,In_303,In_1328);
or U4514 (N_4514,In_1108,In_1095);
xor U4515 (N_4515,In_369,In_1145);
and U4516 (N_4516,In_287,In_554);
and U4517 (N_4517,In_306,In_599);
or U4518 (N_4518,In_1320,In_968);
and U4519 (N_4519,In_482,In_780);
nand U4520 (N_4520,In_46,In_1319);
nand U4521 (N_4521,In_689,In_947);
nand U4522 (N_4522,In_3,In_1244);
nand U4523 (N_4523,In_975,In_1272);
nand U4524 (N_4524,In_1441,In_1171);
or U4525 (N_4525,In_48,In_109);
or U4526 (N_4526,In_326,In_1123);
xor U4527 (N_4527,In_641,In_812);
nor U4528 (N_4528,In_528,In_1299);
or U4529 (N_4529,In_293,In_1408);
xnor U4530 (N_4530,In_1043,In_577);
nor U4531 (N_4531,In_725,In_974);
nand U4532 (N_4532,In_1377,In_892);
or U4533 (N_4533,In_147,In_1154);
and U4534 (N_4534,In_344,In_1427);
xnor U4535 (N_4535,In_1399,In_1078);
nand U4536 (N_4536,In_1425,In_1258);
xnor U4537 (N_4537,In_163,In_1107);
or U4538 (N_4538,In_1169,In_193);
and U4539 (N_4539,In_1060,In_1356);
nand U4540 (N_4540,In_745,In_1044);
nor U4541 (N_4541,In_1132,In_1406);
nand U4542 (N_4542,In_940,In_1132);
and U4543 (N_4543,In_704,In_386);
and U4544 (N_4544,In_1486,In_382);
and U4545 (N_4545,In_1324,In_810);
and U4546 (N_4546,In_1338,In_1047);
nand U4547 (N_4547,In_1268,In_1309);
nand U4548 (N_4548,In_1325,In_1022);
or U4549 (N_4549,In_20,In_1409);
xnor U4550 (N_4550,In_702,In_941);
xnor U4551 (N_4551,In_1435,In_596);
nor U4552 (N_4552,In_472,In_38);
nand U4553 (N_4553,In_781,In_127);
xnor U4554 (N_4554,In_603,In_1403);
and U4555 (N_4555,In_984,In_216);
and U4556 (N_4556,In_1175,In_1351);
or U4557 (N_4557,In_377,In_1178);
and U4558 (N_4558,In_632,In_183);
xnor U4559 (N_4559,In_269,In_410);
or U4560 (N_4560,In_493,In_1195);
xnor U4561 (N_4561,In_336,In_15);
or U4562 (N_4562,In_1197,In_666);
nor U4563 (N_4563,In_711,In_162);
and U4564 (N_4564,In_428,In_1052);
nand U4565 (N_4565,In_985,In_1131);
nor U4566 (N_4566,In_1373,In_1315);
xnor U4567 (N_4567,In_399,In_180);
and U4568 (N_4568,In_21,In_343);
and U4569 (N_4569,In_514,In_991);
nand U4570 (N_4570,In_1028,In_152);
or U4571 (N_4571,In_202,In_20);
nor U4572 (N_4572,In_1050,In_754);
and U4573 (N_4573,In_417,In_830);
nand U4574 (N_4574,In_556,In_1091);
and U4575 (N_4575,In_793,In_1460);
nor U4576 (N_4576,In_46,In_771);
nand U4577 (N_4577,In_1147,In_39);
nand U4578 (N_4578,In_1134,In_1410);
and U4579 (N_4579,In_1003,In_501);
xnor U4580 (N_4580,In_519,In_849);
and U4581 (N_4581,In_450,In_1402);
and U4582 (N_4582,In_715,In_79);
or U4583 (N_4583,In_392,In_280);
or U4584 (N_4584,In_1379,In_850);
or U4585 (N_4585,In_603,In_68);
and U4586 (N_4586,In_528,In_133);
or U4587 (N_4587,In_768,In_170);
nand U4588 (N_4588,In_1238,In_988);
xnor U4589 (N_4589,In_336,In_1429);
nand U4590 (N_4590,In_1070,In_573);
nor U4591 (N_4591,In_214,In_236);
xor U4592 (N_4592,In_965,In_1111);
nor U4593 (N_4593,In_193,In_533);
nor U4594 (N_4594,In_358,In_104);
or U4595 (N_4595,In_346,In_571);
nor U4596 (N_4596,In_1159,In_100);
and U4597 (N_4597,In_272,In_1048);
or U4598 (N_4598,In_1277,In_982);
nand U4599 (N_4599,In_582,In_1260);
or U4600 (N_4600,In_721,In_387);
nor U4601 (N_4601,In_877,In_286);
or U4602 (N_4602,In_351,In_1325);
and U4603 (N_4603,In_762,In_1301);
nor U4604 (N_4604,In_1494,In_870);
nor U4605 (N_4605,In_993,In_71);
or U4606 (N_4606,In_1202,In_596);
nand U4607 (N_4607,In_1384,In_1171);
nor U4608 (N_4608,In_415,In_169);
xor U4609 (N_4609,In_578,In_666);
or U4610 (N_4610,In_1401,In_1125);
xnor U4611 (N_4611,In_1389,In_916);
and U4612 (N_4612,In_961,In_1092);
xnor U4613 (N_4613,In_1104,In_1314);
nor U4614 (N_4614,In_57,In_56);
xnor U4615 (N_4615,In_321,In_813);
xnor U4616 (N_4616,In_942,In_926);
and U4617 (N_4617,In_1103,In_270);
nor U4618 (N_4618,In_354,In_1198);
xor U4619 (N_4619,In_1036,In_783);
nor U4620 (N_4620,In_1311,In_214);
xnor U4621 (N_4621,In_843,In_773);
xor U4622 (N_4622,In_227,In_1047);
and U4623 (N_4623,In_1267,In_1452);
nor U4624 (N_4624,In_557,In_1376);
or U4625 (N_4625,In_106,In_109);
xnor U4626 (N_4626,In_572,In_1249);
xor U4627 (N_4627,In_520,In_1112);
nor U4628 (N_4628,In_1432,In_1206);
nor U4629 (N_4629,In_799,In_1361);
or U4630 (N_4630,In_365,In_444);
nor U4631 (N_4631,In_492,In_221);
xor U4632 (N_4632,In_432,In_293);
xor U4633 (N_4633,In_514,In_942);
nand U4634 (N_4634,In_959,In_202);
xnor U4635 (N_4635,In_999,In_1463);
or U4636 (N_4636,In_1022,In_118);
and U4637 (N_4637,In_1408,In_583);
nand U4638 (N_4638,In_180,In_302);
nor U4639 (N_4639,In_922,In_1458);
nor U4640 (N_4640,In_3,In_1139);
and U4641 (N_4641,In_1129,In_932);
or U4642 (N_4642,In_1444,In_29);
nand U4643 (N_4643,In_205,In_232);
nor U4644 (N_4644,In_1179,In_1);
nand U4645 (N_4645,In_290,In_1022);
and U4646 (N_4646,In_308,In_514);
and U4647 (N_4647,In_945,In_1399);
nand U4648 (N_4648,In_1185,In_1112);
nand U4649 (N_4649,In_427,In_158);
and U4650 (N_4650,In_1063,In_836);
nor U4651 (N_4651,In_811,In_1495);
and U4652 (N_4652,In_293,In_69);
or U4653 (N_4653,In_1306,In_1395);
nor U4654 (N_4654,In_631,In_162);
nand U4655 (N_4655,In_481,In_1157);
and U4656 (N_4656,In_1228,In_1423);
xor U4657 (N_4657,In_1033,In_595);
nor U4658 (N_4658,In_335,In_599);
or U4659 (N_4659,In_1395,In_670);
and U4660 (N_4660,In_399,In_650);
or U4661 (N_4661,In_213,In_304);
and U4662 (N_4662,In_1126,In_849);
xnor U4663 (N_4663,In_871,In_273);
xor U4664 (N_4664,In_590,In_1431);
nor U4665 (N_4665,In_1047,In_697);
xnor U4666 (N_4666,In_116,In_671);
nand U4667 (N_4667,In_1226,In_416);
and U4668 (N_4668,In_798,In_20);
nor U4669 (N_4669,In_183,In_353);
nand U4670 (N_4670,In_969,In_1404);
and U4671 (N_4671,In_14,In_556);
and U4672 (N_4672,In_960,In_92);
nor U4673 (N_4673,In_1157,In_116);
xnor U4674 (N_4674,In_989,In_932);
nor U4675 (N_4675,In_258,In_463);
xor U4676 (N_4676,In_231,In_1371);
nor U4677 (N_4677,In_798,In_1141);
and U4678 (N_4678,In_1170,In_696);
nand U4679 (N_4679,In_1249,In_960);
and U4680 (N_4680,In_98,In_180);
or U4681 (N_4681,In_1354,In_985);
nor U4682 (N_4682,In_31,In_901);
xor U4683 (N_4683,In_299,In_1438);
or U4684 (N_4684,In_538,In_1383);
xor U4685 (N_4685,In_1284,In_654);
nand U4686 (N_4686,In_1163,In_68);
or U4687 (N_4687,In_272,In_610);
and U4688 (N_4688,In_438,In_621);
or U4689 (N_4689,In_1403,In_1176);
and U4690 (N_4690,In_1345,In_1431);
nor U4691 (N_4691,In_1101,In_957);
and U4692 (N_4692,In_40,In_1044);
nor U4693 (N_4693,In_346,In_368);
or U4694 (N_4694,In_1384,In_1118);
or U4695 (N_4695,In_1190,In_532);
and U4696 (N_4696,In_456,In_559);
or U4697 (N_4697,In_674,In_431);
nor U4698 (N_4698,In_1022,In_3);
nand U4699 (N_4699,In_442,In_549);
nor U4700 (N_4700,In_148,In_1354);
or U4701 (N_4701,In_871,In_948);
nor U4702 (N_4702,In_868,In_539);
nor U4703 (N_4703,In_236,In_143);
or U4704 (N_4704,In_1429,In_664);
nor U4705 (N_4705,In_1377,In_870);
nor U4706 (N_4706,In_563,In_1353);
nand U4707 (N_4707,In_723,In_774);
nand U4708 (N_4708,In_436,In_446);
nor U4709 (N_4709,In_341,In_508);
and U4710 (N_4710,In_975,In_1429);
xor U4711 (N_4711,In_1024,In_701);
nand U4712 (N_4712,In_778,In_813);
nor U4713 (N_4713,In_1032,In_1294);
and U4714 (N_4714,In_875,In_95);
nor U4715 (N_4715,In_267,In_250);
and U4716 (N_4716,In_951,In_550);
nor U4717 (N_4717,In_984,In_726);
nor U4718 (N_4718,In_362,In_325);
xor U4719 (N_4719,In_1488,In_13);
nand U4720 (N_4720,In_1485,In_905);
xnor U4721 (N_4721,In_1115,In_259);
or U4722 (N_4722,In_138,In_1247);
nand U4723 (N_4723,In_126,In_641);
nand U4724 (N_4724,In_1157,In_893);
or U4725 (N_4725,In_497,In_1068);
nor U4726 (N_4726,In_862,In_110);
or U4727 (N_4727,In_1346,In_453);
or U4728 (N_4728,In_66,In_43);
or U4729 (N_4729,In_853,In_142);
and U4730 (N_4730,In_1326,In_268);
and U4731 (N_4731,In_655,In_1082);
xnor U4732 (N_4732,In_549,In_343);
xnor U4733 (N_4733,In_972,In_608);
or U4734 (N_4734,In_758,In_251);
or U4735 (N_4735,In_595,In_966);
nor U4736 (N_4736,In_543,In_229);
nor U4737 (N_4737,In_860,In_48);
xor U4738 (N_4738,In_67,In_382);
or U4739 (N_4739,In_253,In_917);
xor U4740 (N_4740,In_349,In_92);
or U4741 (N_4741,In_614,In_944);
and U4742 (N_4742,In_104,In_1373);
and U4743 (N_4743,In_767,In_778);
nor U4744 (N_4744,In_727,In_1466);
or U4745 (N_4745,In_1164,In_814);
nor U4746 (N_4746,In_828,In_1005);
and U4747 (N_4747,In_1457,In_1434);
xor U4748 (N_4748,In_503,In_1147);
and U4749 (N_4749,In_1216,In_508);
xnor U4750 (N_4750,In_606,In_1167);
or U4751 (N_4751,In_1147,In_1385);
nor U4752 (N_4752,In_657,In_459);
xnor U4753 (N_4753,In_379,In_217);
nand U4754 (N_4754,In_1252,In_729);
xnor U4755 (N_4755,In_1105,In_307);
nand U4756 (N_4756,In_333,In_569);
nor U4757 (N_4757,In_142,In_274);
nor U4758 (N_4758,In_1007,In_32);
nand U4759 (N_4759,In_1195,In_242);
or U4760 (N_4760,In_1174,In_244);
and U4761 (N_4761,In_1223,In_1045);
and U4762 (N_4762,In_326,In_1487);
nand U4763 (N_4763,In_813,In_1240);
nor U4764 (N_4764,In_251,In_1056);
or U4765 (N_4765,In_280,In_31);
nor U4766 (N_4766,In_1016,In_370);
and U4767 (N_4767,In_1258,In_1067);
xnor U4768 (N_4768,In_1279,In_702);
nand U4769 (N_4769,In_651,In_1002);
nor U4770 (N_4770,In_925,In_1105);
nand U4771 (N_4771,In_1070,In_351);
nand U4772 (N_4772,In_1436,In_159);
nand U4773 (N_4773,In_1483,In_716);
nand U4774 (N_4774,In_70,In_490);
and U4775 (N_4775,In_468,In_800);
xor U4776 (N_4776,In_409,In_865);
and U4777 (N_4777,In_1178,In_960);
and U4778 (N_4778,In_240,In_138);
nor U4779 (N_4779,In_482,In_699);
xnor U4780 (N_4780,In_1002,In_672);
or U4781 (N_4781,In_870,In_436);
nor U4782 (N_4782,In_901,In_1179);
and U4783 (N_4783,In_1165,In_735);
nand U4784 (N_4784,In_387,In_1214);
or U4785 (N_4785,In_436,In_875);
nand U4786 (N_4786,In_443,In_1497);
or U4787 (N_4787,In_552,In_180);
nor U4788 (N_4788,In_700,In_1020);
nor U4789 (N_4789,In_207,In_708);
and U4790 (N_4790,In_1419,In_1299);
or U4791 (N_4791,In_33,In_696);
nand U4792 (N_4792,In_208,In_456);
or U4793 (N_4793,In_1002,In_1053);
and U4794 (N_4794,In_723,In_629);
xor U4795 (N_4795,In_1033,In_189);
nor U4796 (N_4796,In_961,In_37);
nor U4797 (N_4797,In_1230,In_465);
and U4798 (N_4798,In_987,In_133);
nor U4799 (N_4799,In_48,In_1066);
nand U4800 (N_4800,In_1185,In_1452);
or U4801 (N_4801,In_1305,In_1401);
and U4802 (N_4802,In_482,In_10);
xor U4803 (N_4803,In_307,In_837);
xnor U4804 (N_4804,In_241,In_95);
nor U4805 (N_4805,In_602,In_201);
nor U4806 (N_4806,In_1337,In_1150);
or U4807 (N_4807,In_1272,In_549);
nor U4808 (N_4808,In_859,In_994);
or U4809 (N_4809,In_100,In_1078);
and U4810 (N_4810,In_1400,In_106);
nor U4811 (N_4811,In_130,In_756);
nand U4812 (N_4812,In_1104,In_726);
or U4813 (N_4813,In_1391,In_1265);
nor U4814 (N_4814,In_1448,In_481);
nand U4815 (N_4815,In_204,In_237);
nand U4816 (N_4816,In_1364,In_469);
nand U4817 (N_4817,In_1395,In_173);
and U4818 (N_4818,In_1361,In_449);
or U4819 (N_4819,In_70,In_404);
nor U4820 (N_4820,In_998,In_544);
nand U4821 (N_4821,In_451,In_1444);
or U4822 (N_4822,In_128,In_453);
nor U4823 (N_4823,In_325,In_323);
nand U4824 (N_4824,In_794,In_706);
xnor U4825 (N_4825,In_910,In_580);
nor U4826 (N_4826,In_205,In_690);
nand U4827 (N_4827,In_404,In_808);
and U4828 (N_4828,In_658,In_66);
or U4829 (N_4829,In_906,In_236);
and U4830 (N_4830,In_1075,In_350);
nand U4831 (N_4831,In_1255,In_928);
or U4832 (N_4832,In_420,In_570);
nand U4833 (N_4833,In_260,In_966);
xor U4834 (N_4834,In_56,In_1433);
or U4835 (N_4835,In_722,In_137);
xor U4836 (N_4836,In_1148,In_560);
nand U4837 (N_4837,In_14,In_200);
nand U4838 (N_4838,In_19,In_1137);
nand U4839 (N_4839,In_599,In_649);
nor U4840 (N_4840,In_196,In_90);
and U4841 (N_4841,In_368,In_145);
and U4842 (N_4842,In_507,In_423);
or U4843 (N_4843,In_1439,In_452);
nand U4844 (N_4844,In_235,In_461);
and U4845 (N_4845,In_1303,In_1384);
or U4846 (N_4846,In_442,In_153);
xor U4847 (N_4847,In_997,In_99);
or U4848 (N_4848,In_1036,In_674);
nand U4849 (N_4849,In_786,In_317);
xor U4850 (N_4850,In_325,In_696);
nand U4851 (N_4851,In_1484,In_539);
nand U4852 (N_4852,In_635,In_581);
xnor U4853 (N_4853,In_162,In_485);
nand U4854 (N_4854,In_260,In_1025);
nand U4855 (N_4855,In_1388,In_510);
nor U4856 (N_4856,In_486,In_648);
nand U4857 (N_4857,In_826,In_386);
and U4858 (N_4858,In_296,In_1384);
nor U4859 (N_4859,In_17,In_1089);
xnor U4860 (N_4860,In_294,In_328);
or U4861 (N_4861,In_417,In_530);
and U4862 (N_4862,In_317,In_184);
nand U4863 (N_4863,In_492,In_1413);
nor U4864 (N_4864,In_779,In_116);
nor U4865 (N_4865,In_1362,In_1314);
nor U4866 (N_4866,In_25,In_793);
and U4867 (N_4867,In_1082,In_1222);
xnor U4868 (N_4868,In_473,In_527);
and U4869 (N_4869,In_300,In_321);
nand U4870 (N_4870,In_768,In_176);
nor U4871 (N_4871,In_645,In_1365);
xor U4872 (N_4872,In_751,In_1382);
xnor U4873 (N_4873,In_934,In_124);
or U4874 (N_4874,In_239,In_197);
or U4875 (N_4875,In_977,In_811);
or U4876 (N_4876,In_245,In_29);
nor U4877 (N_4877,In_1041,In_1325);
and U4878 (N_4878,In_356,In_371);
nor U4879 (N_4879,In_152,In_1414);
or U4880 (N_4880,In_1405,In_1489);
nor U4881 (N_4881,In_877,In_260);
xor U4882 (N_4882,In_97,In_41);
or U4883 (N_4883,In_1418,In_569);
and U4884 (N_4884,In_207,In_1116);
xnor U4885 (N_4885,In_217,In_885);
nor U4886 (N_4886,In_685,In_917);
and U4887 (N_4887,In_1243,In_504);
xor U4888 (N_4888,In_1211,In_1407);
or U4889 (N_4889,In_119,In_1020);
and U4890 (N_4890,In_359,In_220);
and U4891 (N_4891,In_158,In_903);
nand U4892 (N_4892,In_34,In_178);
or U4893 (N_4893,In_222,In_1069);
nand U4894 (N_4894,In_998,In_374);
nor U4895 (N_4895,In_1485,In_288);
nor U4896 (N_4896,In_1393,In_612);
xor U4897 (N_4897,In_42,In_1098);
xor U4898 (N_4898,In_106,In_825);
nand U4899 (N_4899,In_343,In_461);
and U4900 (N_4900,In_354,In_1352);
or U4901 (N_4901,In_1439,In_638);
nor U4902 (N_4902,In_922,In_1068);
nor U4903 (N_4903,In_1042,In_1285);
and U4904 (N_4904,In_414,In_1298);
nand U4905 (N_4905,In_520,In_578);
nor U4906 (N_4906,In_1421,In_752);
nor U4907 (N_4907,In_988,In_95);
or U4908 (N_4908,In_521,In_191);
xnor U4909 (N_4909,In_1182,In_1233);
and U4910 (N_4910,In_865,In_388);
nand U4911 (N_4911,In_1131,In_463);
xor U4912 (N_4912,In_172,In_1231);
and U4913 (N_4913,In_385,In_1211);
and U4914 (N_4914,In_357,In_43);
and U4915 (N_4915,In_105,In_1471);
nand U4916 (N_4916,In_542,In_498);
nor U4917 (N_4917,In_1033,In_708);
and U4918 (N_4918,In_1157,In_629);
and U4919 (N_4919,In_51,In_1479);
and U4920 (N_4920,In_1388,In_348);
xor U4921 (N_4921,In_1063,In_1286);
or U4922 (N_4922,In_1430,In_634);
or U4923 (N_4923,In_538,In_1406);
nor U4924 (N_4924,In_1410,In_666);
xor U4925 (N_4925,In_153,In_729);
or U4926 (N_4926,In_1024,In_914);
and U4927 (N_4927,In_809,In_723);
nor U4928 (N_4928,In_124,In_73);
and U4929 (N_4929,In_999,In_1402);
and U4930 (N_4930,In_1187,In_344);
nor U4931 (N_4931,In_21,In_1174);
and U4932 (N_4932,In_540,In_778);
nand U4933 (N_4933,In_1090,In_618);
xnor U4934 (N_4934,In_583,In_1243);
or U4935 (N_4935,In_1251,In_916);
nand U4936 (N_4936,In_541,In_27);
nand U4937 (N_4937,In_1168,In_1319);
and U4938 (N_4938,In_1049,In_477);
nor U4939 (N_4939,In_692,In_703);
xor U4940 (N_4940,In_70,In_101);
and U4941 (N_4941,In_39,In_1351);
and U4942 (N_4942,In_941,In_963);
or U4943 (N_4943,In_616,In_855);
and U4944 (N_4944,In_504,In_784);
xnor U4945 (N_4945,In_1075,In_1107);
xor U4946 (N_4946,In_763,In_1268);
and U4947 (N_4947,In_1058,In_285);
and U4948 (N_4948,In_418,In_647);
and U4949 (N_4949,In_1077,In_160);
or U4950 (N_4950,In_316,In_819);
xnor U4951 (N_4951,In_307,In_12);
nand U4952 (N_4952,In_1162,In_1083);
and U4953 (N_4953,In_946,In_597);
xnor U4954 (N_4954,In_1449,In_940);
nor U4955 (N_4955,In_1473,In_1326);
nand U4956 (N_4956,In_852,In_382);
nand U4957 (N_4957,In_26,In_1040);
nand U4958 (N_4958,In_657,In_285);
xnor U4959 (N_4959,In_679,In_198);
xor U4960 (N_4960,In_1046,In_711);
nand U4961 (N_4961,In_1308,In_344);
nor U4962 (N_4962,In_623,In_1463);
xor U4963 (N_4963,In_921,In_337);
nor U4964 (N_4964,In_209,In_562);
xnor U4965 (N_4965,In_1288,In_263);
nor U4966 (N_4966,In_791,In_167);
xor U4967 (N_4967,In_451,In_1092);
nor U4968 (N_4968,In_806,In_623);
xor U4969 (N_4969,In_1235,In_606);
or U4970 (N_4970,In_771,In_96);
nand U4971 (N_4971,In_1352,In_1168);
or U4972 (N_4972,In_765,In_443);
and U4973 (N_4973,In_270,In_788);
xnor U4974 (N_4974,In_821,In_353);
nor U4975 (N_4975,In_678,In_1321);
nor U4976 (N_4976,In_568,In_1297);
nand U4977 (N_4977,In_1104,In_1485);
nand U4978 (N_4978,In_83,In_1379);
nor U4979 (N_4979,In_388,In_1400);
and U4980 (N_4980,In_862,In_847);
and U4981 (N_4981,In_1287,In_58);
nand U4982 (N_4982,In_527,In_91);
xor U4983 (N_4983,In_908,In_1298);
or U4984 (N_4984,In_768,In_52);
nor U4985 (N_4985,In_78,In_541);
or U4986 (N_4986,In_1183,In_1108);
xor U4987 (N_4987,In_1195,In_1069);
nor U4988 (N_4988,In_1299,In_376);
nand U4989 (N_4989,In_445,In_148);
nor U4990 (N_4990,In_456,In_249);
xor U4991 (N_4991,In_466,In_228);
and U4992 (N_4992,In_1354,In_252);
nor U4993 (N_4993,In_115,In_391);
nor U4994 (N_4994,In_1281,In_1094);
xor U4995 (N_4995,In_5,In_324);
and U4996 (N_4996,In_354,In_32);
or U4997 (N_4997,In_652,In_602);
or U4998 (N_4998,In_183,In_837);
and U4999 (N_4999,In_1180,In_657);
and U5000 (N_5000,N_4413,N_2054);
xnor U5001 (N_5001,N_480,N_1933);
xnor U5002 (N_5002,N_4453,N_681);
nand U5003 (N_5003,N_4577,N_3079);
or U5004 (N_5004,N_1468,N_2278);
or U5005 (N_5005,N_2340,N_1415);
nor U5006 (N_5006,N_4858,N_686);
nand U5007 (N_5007,N_733,N_4472);
xnor U5008 (N_5008,N_1740,N_2099);
nor U5009 (N_5009,N_3826,N_1019);
xor U5010 (N_5010,N_3934,N_3739);
nor U5011 (N_5011,N_4836,N_3236);
and U5012 (N_5012,N_795,N_1767);
and U5013 (N_5013,N_812,N_4828);
nand U5014 (N_5014,N_2265,N_4385);
xor U5015 (N_5015,N_1881,N_876);
xor U5016 (N_5016,N_1481,N_927);
nand U5017 (N_5017,N_2722,N_4661);
nand U5018 (N_5018,N_3450,N_4485);
or U5019 (N_5019,N_1062,N_4639);
or U5020 (N_5020,N_775,N_4144);
nor U5021 (N_5021,N_2080,N_2495);
nand U5022 (N_5022,N_2146,N_3539);
nor U5023 (N_5023,N_4040,N_994);
nand U5024 (N_5024,N_1986,N_4308);
xnor U5025 (N_5025,N_4362,N_3312);
nand U5026 (N_5026,N_4424,N_2548);
nor U5027 (N_5027,N_4408,N_383);
xnor U5028 (N_5028,N_1696,N_3777);
nor U5029 (N_5029,N_4437,N_4082);
nand U5030 (N_5030,N_3086,N_3679);
xor U5031 (N_5031,N_749,N_1266);
nor U5032 (N_5032,N_785,N_1935);
xor U5033 (N_5033,N_168,N_4815);
nand U5034 (N_5034,N_902,N_765);
and U5035 (N_5035,N_2177,N_474);
xor U5036 (N_5036,N_1279,N_719);
nand U5037 (N_5037,N_111,N_3);
or U5038 (N_5038,N_913,N_3230);
and U5039 (N_5039,N_266,N_4176);
nand U5040 (N_5040,N_2403,N_717);
nor U5041 (N_5041,N_1204,N_2275);
xor U5042 (N_5042,N_107,N_2151);
or U5043 (N_5043,N_1046,N_2853);
or U5044 (N_5044,N_536,N_4683);
nand U5045 (N_5045,N_4099,N_2685);
or U5046 (N_5046,N_260,N_4831);
nor U5047 (N_5047,N_4512,N_2978);
and U5048 (N_5048,N_4244,N_2163);
or U5049 (N_5049,N_1825,N_557);
or U5050 (N_5050,N_4714,N_2726);
xor U5051 (N_5051,N_4026,N_2824);
or U5052 (N_5052,N_3529,N_360);
xnor U5053 (N_5053,N_1229,N_1166);
nand U5054 (N_5054,N_2704,N_81);
and U5055 (N_5055,N_2680,N_933);
xor U5056 (N_5056,N_583,N_2964);
xnor U5057 (N_5057,N_3921,N_4295);
or U5058 (N_5058,N_3518,N_864);
nand U5059 (N_5059,N_2049,N_4280);
and U5060 (N_5060,N_143,N_2349);
or U5061 (N_5061,N_3725,N_1960);
xor U5062 (N_5062,N_4880,N_3639);
nand U5063 (N_5063,N_3972,N_4536);
nor U5064 (N_5064,N_3856,N_199);
and U5065 (N_5065,N_4812,N_2612);
and U5066 (N_5066,N_4998,N_712);
or U5067 (N_5067,N_1234,N_1367);
nand U5068 (N_5068,N_3806,N_2191);
or U5069 (N_5069,N_2221,N_3437);
or U5070 (N_5070,N_3272,N_715);
or U5071 (N_5071,N_4234,N_1450);
and U5072 (N_5072,N_3609,N_3495);
and U5073 (N_5073,N_3906,N_297);
nor U5074 (N_5074,N_357,N_1514);
nand U5075 (N_5075,N_4595,N_836);
xor U5076 (N_5076,N_2208,N_842);
and U5077 (N_5077,N_3748,N_1555);
xnor U5078 (N_5078,N_4618,N_2679);
and U5079 (N_5079,N_2481,N_4327);
nand U5080 (N_5080,N_1303,N_2381);
xor U5081 (N_5081,N_2241,N_308);
or U5082 (N_5082,N_1274,N_2476);
nor U5083 (N_5083,N_2709,N_4449);
nor U5084 (N_5084,N_2107,N_2301);
xor U5085 (N_5085,N_3107,N_3523);
and U5086 (N_5086,N_4563,N_4587);
or U5087 (N_5087,N_181,N_1969);
xnor U5088 (N_5088,N_2172,N_4523);
and U5089 (N_5089,N_2098,N_548);
xnor U5090 (N_5090,N_1871,N_1714);
xnor U5091 (N_5091,N_3218,N_4283);
and U5092 (N_5092,N_2423,N_2510);
nand U5093 (N_5093,N_1212,N_4252);
xnor U5094 (N_5094,N_607,N_4692);
xnor U5095 (N_5095,N_643,N_4636);
nand U5096 (N_5096,N_4111,N_130);
nand U5097 (N_5097,N_1444,N_2549);
or U5098 (N_5098,N_2259,N_3543);
nor U5099 (N_5099,N_665,N_1943);
nand U5100 (N_5100,N_3515,N_1717);
nor U5101 (N_5101,N_2742,N_4046);
and U5102 (N_5102,N_907,N_2977);
nor U5103 (N_5103,N_696,N_4415);
nor U5104 (N_5104,N_1895,N_4806);
or U5105 (N_5105,N_2834,N_2916);
xnor U5106 (N_5106,N_1656,N_2619);
or U5107 (N_5107,N_3187,N_3492);
or U5108 (N_5108,N_568,N_75);
and U5109 (N_5109,N_3728,N_4717);
or U5110 (N_5110,N_2856,N_2696);
or U5111 (N_5111,N_1894,N_4411);
nand U5112 (N_5112,N_1304,N_4544);
xnor U5113 (N_5113,N_1693,N_2527);
nor U5114 (N_5114,N_1498,N_998);
nor U5115 (N_5115,N_1256,N_2184);
and U5116 (N_5116,N_3783,N_3595);
and U5117 (N_5117,N_3167,N_3546);
or U5118 (N_5118,N_2991,N_2873);
nor U5119 (N_5119,N_4432,N_1971);
or U5120 (N_5120,N_3519,N_4552);
nor U5121 (N_5121,N_1025,N_3023);
and U5122 (N_5122,N_1064,N_115);
or U5123 (N_5123,N_1194,N_1168);
and U5124 (N_5124,N_4063,N_1829);
and U5125 (N_5125,N_3036,N_3105);
nor U5126 (N_5126,N_125,N_3306);
nand U5127 (N_5127,N_4316,N_2953);
nand U5128 (N_5128,N_3397,N_3724);
and U5129 (N_5129,N_1142,N_2186);
or U5130 (N_5130,N_4266,N_3102);
nor U5131 (N_5131,N_4827,N_4072);
or U5132 (N_5132,N_1100,N_2695);
nand U5133 (N_5133,N_4065,N_2229);
and U5134 (N_5134,N_4908,N_3302);
nor U5135 (N_5135,N_3096,N_4312);
or U5136 (N_5136,N_2993,N_179);
nor U5137 (N_5137,N_4669,N_4750);
nor U5138 (N_5138,N_2321,N_611);
and U5139 (N_5139,N_2712,N_2963);
nor U5140 (N_5140,N_3235,N_2001);
nand U5141 (N_5141,N_2741,N_829);
or U5142 (N_5142,N_889,N_1078);
nand U5143 (N_5143,N_1283,N_3034);
nand U5144 (N_5144,N_3224,N_1698);
xor U5145 (N_5145,N_798,N_4925);
nor U5146 (N_5146,N_4937,N_1753);
xor U5147 (N_5147,N_310,N_2504);
nor U5148 (N_5148,N_4582,N_1291);
and U5149 (N_5149,N_755,N_2546);
nor U5150 (N_5150,N_1086,N_3172);
nor U5151 (N_5151,N_3173,N_2684);
xor U5152 (N_5152,N_4906,N_1772);
or U5153 (N_5153,N_1382,N_370);
or U5154 (N_5154,N_791,N_1116);
xor U5155 (N_5155,N_4110,N_2708);
or U5156 (N_5156,N_493,N_3415);
nor U5157 (N_5157,N_1954,N_24);
xnor U5158 (N_5158,N_1582,N_513);
nand U5159 (N_5159,N_1118,N_764);
nand U5160 (N_5160,N_4975,N_1641);
xnor U5161 (N_5161,N_4678,N_3967);
xnor U5162 (N_5162,N_3249,N_2567);
and U5163 (N_5163,N_4477,N_3401);
nor U5164 (N_5164,N_211,N_546);
nor U5165 (N_5165,N_2036,N_1667);
nor U5166 (N_5166,N_3631,N_2813);
and U5167 (N_5167,N_534,N_102);
or U5168 (N_5168,N_948,N_649);
and U5169 (N_5169,N_379,N_3900);
nor U5170 (N_5170,N_4847,N_3115);
xor U5171 (N_5171,N_591,N_1319);
nand U5172 (N_5172,N_1126,N_3993);
nand U5173 (N_5173,N_159,N_952);
nor U5174 (N_5174,N_641,N_1195);
nor U5175 (N_5175,N_1316,N_1040);
nor U5176 (N_5176,N_2234,N_2204);
nor U5177 (N_5177,N_1542,N_1685);
nor U5178 (N_5178,N_1818,N_1694);
nand U5179 (N_5179,N_2297,N_3720);
or U5180 (N_5180,N_2884,N_3222);
and U5181 (N_5181,N_3947,N_4374);
nand U5182 (N_5182,N_3267,N_2985);
xor U5183 (N_5183,N_1965,N_1742);
or U5184 (N_5184,N_2390,N_4301);
nor U5185 (N_5185,N_149,N_3380);
and U5186 (N_5186,N_4429,N_1392);
xnor U5187 (N_5187,N_4033,N_243);
nor U5188 (N_5188,N_3031,N_3298);
nand U5189 (N_5189,N_1573,N_589);
or U5190 (N_5190,N_4541,N_4599);
xnor U5191 (N_5191,N_1037,N_1006);
nand U5192 (N_5192,N_1684,N_3866);
xor U5193 (N_5193,N_1606,N_2595);
or U5194 (N_5194,N_2176,N_70);
nor U5195 (N_5195,N_232,N_3367);
or U5196 (N_5196,N_3727,N_4042);
nand U5197 (N_5197,N_858,N_27);
and U5198 (N_5198,N_3038,N_1120);
or U5199 (N_5199,N_3955,N_3604);
xor U5200 (N_5200,N_3000,N_4859);
nand U5201 (N_5201,N_2825,N_106);
nor U5202 (N_5202,N_1524,N_1587);
or U5203 (N_5203,N_4874,N_737);
xnor U5204 (N_5204,N_2010,N_3558);
and U5205 (N_5205,N_4410,N_3371);
and U5206 (N_5206,N_4835,N_2168);
nor U5207 (N_5207,N_3333,N_581);
and U5208 (N_5208,N_1646,N_1403);
nor U5209 (N_5209,N_3124,N_571);
nor U5210 (N_5210,N_3001,N_1790);
or U5211 (N_5211,N_4212,N_4559);
nand U5212 (N_5212,N_869,N_986);
and U5213 (N_5213,N_3471,N_277);
xnor U5214 (N_5214,N_1512,N_3636);
nand U5215 (N_5215,N_4565,N_4237);
or U5216 (N_5216,N_3940,N_4751);
nor U5217 (N_5217,N_2996,N_3088);
xor U5218 (N_5218,N_2909,N_2669);
nand U5219 (N_5219,N_4757,N_909);
xnor U5220 (N_5220,N_3575,N_3910);
nor U5221 (N_5221,N_1292,N_2430);
nand U5222 (N_5222,N_2921,N_76);
and U5223 (N_5223,N_2109,N_3688);
nand U5224 (N_5224,N_4753,N_4337);
nand U5225 (N_5225,N_1855,N_4579);
nor U5226 (N_5226,N_2749,N_4960);
xor U5227 (N_5227,N_1664,N_3773);
nor U5228 (N_5228,N_2250,N_2769);
nand U5229 (N_5229,N_1617,N_2694);
and U5230 (N_5230,N_4100,N_153);
nand U5231 (N_5231,N_1087,N_3328);
nand U5232 (N_5232,N_3377,N_1690);
nand U5233 (N_5233,N_1349,N_3442);
nor U5234 (N_5234,N_3532,N_3851);
nand U5235 (N_5235,N_3629,N_1243);
xnor U5236 (N_5236,N_2744,N_2795);
nor U5237 (N_5237,N_4359,N_414);
nand U5238 (N_5238,N_3412,N_547);
nand U5239 (N_5239,N_293,N_1830);
and U5240 (N_5240,N_2243,N_1858);
or U5241 (N_5241,N_3895,N_4175);
and U5242 (N_5242,N_1501,N_2920);
or U5243 (N_5243,N_3308,N_3952);
xnor U5244 (N_5244,N_1278,N_2473);
and U5245 (N_5245,N_567,N_1550);
and U5246 (N_5246,N_1788,N_1675);
nor U5247 (N_5247,N_4824,N_2106);
nor U5248 (N_5248,N_3215,N_3880);
xor U5249 (N_5249,N_4759,N_3689);
or U5250 (N_5250,N_1936,N_1074);
nand U5251 (N_5251,N_1990,N_999);
or U5252 (N_5252,N_2550,N_1668);
nor U5253 (N_5253,N_4606,N_2863);
nand U5254 (N_5254,N_4353,N_3081);
and U5255 (N_5255,N_1504,N_1624);
nand U5256 (N_5256,N_804,N_1532);
nor U5257 (N_5257,N_2335,N_1370);
nand U5258 (N_5258,N_1576,N_2118);
xnor U5259 (N_5259,N_714,N_1133);
and U5260 (N_5260,N_2526,N_4401);
nand U5261 (N_5261,N_387,N_1336);
or U5262 (N_5262,N_2312,N_3391);
or U5263 (N_5263,N_1193,N_3445);
nand U5264 (N_5264,N_4896,N_4241);
nand U5265 (N_5265,N_821,N_3787);
xor U5266 (N_5266,N_3290,N_3123);
nand U5267 (N_5267,N_273,N_2809);
nand U5268 (N_5268,N_1955,N_1779);
nand U5269 (N_5269,N_4917,N_3127);
nor U5270 (N_5270,N_1391,N_4631);
or U5271 (N_5271,N_2427,N_1785);
and U5272 (N_5272,N_1534,N_3907);
or U5273 (N_5273,N_3411,N_205);
nor U5274 (N_5274,N_1994,N_4628);
nand U5275 (N_5275,N_3231,N_3602);
or U5276 (N_5276,N_2268,N_947);
or U5277 (N_5277,N_4687,N_659);
nand U5278 (N_5278,N_1063,N_1160);
xnor U5279 (N_5279,N_4010,N_1502);
or U5280 (N_5280,N_3588,N_2305);
or U5281 (N_5281,N_4403,N_3920);
nand U5282 (N_5282,N_2511,N_2435);
and U5283 (N_5283,N_2363,N_3845);
nor U5284 (N_5284,N_3987,N_1096);
nor U5285 (N_5285,N_967,N_3911);
xnor U5286 (N_5286,N_295,N_875);
xnor U5287 (N_5287,N_3619,N_66);
nor U5288 (N_5288,N_904,N_332);
nand U5289 (N_5289,N_4774,N_2911);
xor U5290 (N_5290,N_3019,N_2564);
nand U5291 (N_5291,N_1977,N_21);
or U5292 (N_5292,N_2678,N_4138);
or U5293 (N_5293,N_4288,N_2458);
and U5294 (N_5294,N_4557,N_306);
and U5295 (N_5295,N_1932,N_940);
or U5296 (N_5296,N_1929,N_2617);
and U5297 (N_5297,N_2030,N_4643);
nand U5298 (N_5298,N_1163,N_2665);
and U5299 (N_5299,N_2491,N_4166);
or U5300 (N_5300,N_2521,N_4701);
or U5301 (N_5301,N_4293,N_3646);
nor U5302 (N_5302,N_3563,N_3622);
and U5303 (N_5303,N_3140,N_2952);
or U5304 (N_5304,N_1334,N_209);
nor U5305 (N_5305,N_3875,N_3175);
and U5306 (N_5306,N_2757,N_1378);
xnor U5307 (N_5307,N_3944,N_3072);
nand U5308 (N_5308,N_1672,N_3663);
nor U5309 (N_5309,N_1429,N_3058);
nand U5310 (N_5310,N_3590,N_4603);
xor U5311 (N_5311,N_4051,N_1139);
xnor U5312 (N_5312,N_2577,N_2868);
xnor U5313 (N_5313,N_741,N_3159);
nand U5314 (N_5314,N_1080,N_406);
and U5315 (N_5315,N_1101,N_1591);
or U5316 (N_5316,N_2707,N_2981);
nand U5317 (N_5317,N_2497,N_2506);
xnor U5318 (N_5318,N_4270,N_3672);
xor U5319 (N_5319,N_1431,N_1456);
nand U5320 (N_5320,N_207,N_2072);
or U5321 (N_5321,N_4676,N_915);
or U5322 (N_5322,N_2675,N_3100);
xor U5323 (N_5323,N_1903,N_1230);
or U5324 (N_5324,N_2671,N_4043);
and U5325 (N_5325,N_4102,N_3419);
nor U5326 (N_5326,N_3149,N_3796);
nand U5327 (N_5327,N_169,N_1622);
xor U5328 (N_5328,N_1457,N_3174);
xor U5329 (N_5329,N_4470,N_2998);
xor U5330 (N_5330,N_4963,N_2202);
or U5331 (N_5331,N_2426,N_1776);
xnor U5332 (N_5332,N_3744,N_362);
nor U5333 (N_5333,N_3007,N_3449);
and U5334 (N_5334,N_2294,N_4145);
nor U5335 (N_5335,N_1615,N_2345);
or U5336 (N_5336,N_1518,N_1688);
and U5337 (N_5337,N_3094,N_4200);
nor U5338 (N_5338,N_2289,N_708);
and U5339 (N_5339,N_4133,N_704);
nor U5340 (N_5340,N_4348,N_3797);
nor U5341 (N_5341,N_955,N_818);
or U5342 (N_5342,N_827,N_1173);
xor U5343 (N_5343,N_3014,N_4648);
or U5344 (N_5344,N_3476,N_978);
xnor U5345 (N_5345,N_4224,N_2195);
nand U5346 (N_5346,N_3627,N_1511);
nor U5347 (N_5347,N_2732,N_1143);
nor U5348 (N_5348,N_2496,N_1655);
xor U5349 (N_5349,N_4141,N_3360);
nand U5350 (N_5350,N_3238,N_3786);
nor U5351 (N_5351,N_3112,N_1397);
and U5352 (N_5352,N_3747,N_3752);
xnor U5353 (N_5353,N_2849,N_442);
nor U5354 (N_5354,N_753,N_122);
or U5355 (N_5355,N_3586,N_4814);
or U5356 (N_5356,N_3370,N_2810);
nand U5357 (N_5357,N_202,N_2892);
or U5358 (N_5358,N_1738,N_1595);
xor U5359 (N_5359,N_516,N_3067);
xnor U5360 (N_5360,N_910,N_1566);
nand U5361 (N_5361,N_3152,N_4131);
nor U5362 (N_5362,N_109,N_1634);
nor U5363 (N_5363,N_2645,N_3745);
or U5364 (N_5364,N_4510,N_3489);
or U5365 (N_5365,N_809,N_1343);
xor U5366 (N_5366,N_2083,N_1347);
nor U5367 (N_5367,N_4656,N_338);
xor U5368 (N_5368,N_4089,N_428);
xor U5369 (N_5369,N_403,N_3874);
nand U5370 (N_5370,N_3779,N_3559);
nor U5371 (N_5371,N_2937,N_1232);
or U5372 (N_5372,N_4018,N_4671);
nand U5373 (N_5373,N_4402,N_4736);
nand U5374 (N_5374,N_185,N_2091);
or U5375 (N_5375,N_1540,N_3999);
and U5376 (N_5376,N_4689,N_1048);
and U5377 (N_5377,N_238,N_3362);
xnor U5378 (N_5378,N_2125,N_3686);
nor U5379 (N_5379,N_4733,N_2999);
nor U5380 (N_5380,N_2563,N_2216);
nor U5381 (N_5381,N_1997,N_2288);
nor U5382 (N_5382,N_3894,N_2950);
or U5383 (N_5383,N_3936,N_3035);
nor U5384 (N_5384,N_4808,N_4680);
nand U5385 (N_5385,N_1843,N_826);
and U5386 (N_5386,N_1081,N_1546);
nor U5387 (N_5387,N_3042,N_2943);
nand U5388 (N_5388,N_4549,N_3835);
or U5389 (N_5389,N_3300,N_1433);
or U5390 (N_5390,N_31,N_3441);
or U5391 (N_5391,N_738,N_490);
xnor U5392 (N_5392,N_2651,N_326);
xor U5393 (N_5393,N_459,N_1743);
nand U5394 (N_5394,N_650,N_4872);
or U5395 (N_5395,N_1306,N_42);
or U5396 (N_5396,N_4706,N_1221);
xnor U5397 (N_5397,N_4467,N_3690);
xor U5398 (N_5398,N_2702,N_3811);
nand U5399 (N_5399,N_3871,N_2011);
xnor U5400 (N_5400,N_3110,N_4497);
or U5401 (N_5401,N_2697,N_2634);
nor U5402 (N_5402,N_2314,N_4526);
nand U5403 (N_5403,N_289,N_3253);
and U5404 (N_5404,N_1642,N_3956);
or U5405 (N_5405,N_543,N_823);
nand U5406 (N_5406,N_3439,N_4041);
and U5407 (N_5407,N_2362,N_4807);
or U5408 (N_5408,N_4354,N_285);
or U5409 (N_5409,N_3567,N_119);
or U5410 (N_5410,N_227,N_4179);
and U5411 (N_5411,N_386,N_2328);
and U5412 (N_5412,N_3012,N_2487);
nor U5413 (N_5413,N_4129,N_2479);
and U5414 (N_5414,N_2846,N_3633);
nand U5415 (N_5415,N_1891,N_901);
nand U5416 (N_5416,N_3760,N_3403);
and U5417 (N_5417,N_2734,N_2185);
xor U5418 (N_5418,N_2637,N_815);
xor U5419 (N_5419,N_4527,N_355);
and U5420 (N_5420,N_4967,N_4002);
xor U5421 (N_5421,N_1596,N_1928);
nand U5422 (N_5422,N_3615,N_814);
nor U5423 (N_5423,N_863,N_4634);
and U5424 (N_5424,N_2572,N_1909);
nor U5425 (N_5425,N_54,N_240);
or U5426 (N_5426,N_3497,N_438);
nand U5427 (N_5427,N_2592,N_311);
nor U5428 (N_5428,N_3425,N_1366);
nor U5429 (N_5429,N_4162,N_2207);
nand U5430 (N_5430,N_1209,N_4588);
or U5431 (N_5431,N_71,N_1774);
or U5432 (N_5432,N_3057,N_4773);
or U5433 (N_5433,N_3004,N_186);
and U5434 (N_5434,N_478,N_391);
nor U5435 (N_5435,N_3183,N_544);
or U5436 (N_5436,N_2596,N_4001);
nor U5437 (N_5437,N_679,N_2962);
nand U5438 (N_5438,N_1148,N_800);
or U5439 (N_5439,N_4772,N_4848);
or U5440 (N_5440,N_2253,N_898);
nand U5441 (N_5441,N_2533,N_1913);
or U5442 (N_5442,N_2640,N_92);
nand U5443 (N_5443,N_4275,N_1578);
nor U5444 (N_5444,N_4954,N_1381);
nand U5445 (N_5445,N_1477,N_1927);
and U5446 (N_5446,N_661,N_3821);
and U5447 (N_5447,N_4620,N_2615);
nor U5448 (N_5448,N_4537,N_1666);
xor U5449 (N_5449,N_4853,N_4192);
and U5450 (N_5450,N_2635,N_4899);
or U5451 (N_5451,N_1710,N_2974);
nand U5452 (N_5452,N_3277,N_3220);
xor U5453 (N_5453,N_1842,N_1439);
and U5454 (N_5454,N_4292,N_1333);
or U5455 (N_5455,N_3201,N_4747);
nor U5456 (N_5456,N_2382,N_3706);
or U5457 (N_5457,N_203,N_699);
and U5458 (N_5458,N_1594,N_2747);
nor U5459 (N_5459,N_4818,N_540);
nor U5460 (N_5460,N_2105,N_2966);
nor U5461 (N_5461,N_1763,N_4418);
xnor U5462 (N_5462,N_3374,N_1547);
and U5463 (N_5463,N_2832,N_1991);
nor U5464 (N_5464,N_239,N_2193);
nor U5465 (N_5465,N_4343,N_359);
or U5466 (N_5466,N_89,N_4115);
and U5467 (N_5467,N_1470,N_1270);
xor U5468 (N_5468,N_1376,N_1409);
or U5469 (N_5469,N_2965,N_283);
nand U5470 (N_5470,N_3087,N_3202);
or U5471 (N_5471,N_1228,N_4276);
nand U5472 (N_5472,N_4877,N_577);
xor U5473 (N_5473,N_1389,N_1105);
nand U5474 (N_5474,N_3015,N_4381);
nand U5475 (N_5475,N_4699,N_3073);
xor U5476 (N_5476,N_2598,N_4990);
and U5477 (N_5477,N_3251,N_2555);
and U5478 (N_5478,N_3553,N_4457);
nand U5479 (N_5479,N_1325,N_1886);
nor U5480 (N_5480,N_2318,N_729);
xnor U5481 (N_5481,N_2814,N_4569);
nor U5482 (N_5482,N_2463,N_20);
nor U5483 (N_5483,N_2837,N_4630);
xor U5484 (N_5484,N_2958,N_3592);
or U5485 (N_5485,N_1338,N_4048);
nor U5486 (N_5486,N_3775,N_1926);
and U5487 (N_5487,N_2446,N_3343);
nor U5488 (N_5488,N_1357,N_757);
or U5489 (N_5489,N_3054,N_1159);
xnor U5490 (N_5490,N_3628,N_2175);
or U5491 (N_5491,N_158,N_4261);
or U5492 (N_5492,N_236,N_2225);
nor U5493 (N_5493,N_843,N_477);
xnor U5494 (N_5494,N_3893,N_3276);
and U5495 (N_5495,N_4361,N_363);
nand U5496 (N_5496,N_3454,N_1888);
nand U5497 (N_5497,N_4328,N_3765);
or U5498 (N_5498,N_2095,N_1307);
xor U5499 (N_5499,N_446,N_4199);
or U5500 (N_5500,N_4345,N_4688);
and U5501 (N_5501,N_3060,N_4834);
nor U5502 (N_5502,N_3256,N_3984);
nand U5503 (N_5503,N_4326,N_4097);
nand U5504 (N_5504,N_1869,N_1205);
xor U5505 (N_5505,N_2475,N_4518);
xor U5506 (N_5506,N_1419,N_824);
nor U5507 (N_5507,N_885,N_2941);
or U5508 (N_5508,N_3550,N_1180);
nand U5509 (N_5509,N_249,N_4704);
nor U5510 (N_5510,N_3157,N_4551);
and U5511 (N_5511,N_514,N_114);
nand U5512 (N_5512,N_499,N_3062);
xor U5513 (N_5513,N_1027,N_2343);
or U5514 (N_5514,N_1032,N_1358);
nand U5515 (N_5515,N_1531,N_4330);
or U5516 (N_5516,N_4163,N_44);
xnor U5517 (N_5517,N_4466,N_1261);
xor U5518 (N_5518,N_3802,N_1733);
or U5519 (N_5519,N_3985,N_280);
and U5520 (N_5520,N_1302,N_2706);
and U5521 (N_5521,N_2513,N_3331);
nor U5522 (N_5522,N_1823,N_4594);
or U5523 (N_5523,N_3650,N_1979);
xnor U5524 (N_5524,N_2111,N_1169);
nor U5525 (N_5525,N_1156,N_4916);
nor U5526 (N_5526,N_3712,N_524);
or U5527 (N_5527,N_1645,N_3841);
xor U5528 (N_5528,N_2663,N_3847);
and U5529 (N_5529,N_3467,N_3463);
nor U5530 (N_5530,N_323,N_258);
xnor U5531 (N_5531,N_1390,N_3196);
or U5532 (N_5532,N_3506,N_1122);
nor U5533 (N_5533,N_793,N_1762);
or U5534 (N_5534,N_2097,N_1360);
and U5535 (N_5535,N_3462,N_2251);
xor U5536 (N_5536,N_4813,N_2448);
and U5537 (N_5537,N_1420,N_4318);
or U5538 (N_5538,N_69,N_284);
xor U5539 (N_5539,N_2461,N_4304);
nor U5540 (N_5540,N_2575,N_3191);
nor U5541 (N_5541,N_464,N_0);
nor U5542 (N_5542,N_4392,N_1041);
nand U5543 (N_5543,N_519,N_445);
nor U5544 (N_5544,N_2051,N_86);
and U5545 (N_5545,N_3192,N_1179);
nand U5546 (N_5546,N_1070,N_3862);
nand U5547 (N_5547,N_3116,N_3407);
and U5548 (N_5548,N_1993,N_1387);
xnor U5549 (N_5549,N_1052,N_1736);
nand U5550 (N_5550,N_790,N_2532);
and U5551 (N_5551,N_1912,N_2215);
or U5552 (N_5552,N_3171,N_2078);
nand U5553 (N_5553,N_1149,N_4169);
nor U5554 (N_5554,N_3368,N_2529);
or U5555 (N_5555,N_2059,N_3842);
xnor U5556 (N_5556,N_4448,N_710);
nand U5557 (N_5557,N_2517,N_4185);
or U5558 (N_5558,N_4339,N_1964);
or U5559 (N_5559,N_4171,N_1545);
and U5560 (N_5560,N_37,N_364);
nand U5561 (N_5561,N_835,N_4795);
nor U5562 (N_5562,N_2124,N_2071);
and U5563 (N_5563,N_3017,N_4600);
nor U5564 (N_5564,N_1893,N_2027);
xor U5565 (N_5565,N_412,N_4104);
xor U5566 (N_5566,N_3453,N_555);
or U5567 (N_5567,N_4832,N_3348);
xor U5568 (N_5568,N_2857,N_724);
nand U5569 (N_5569,N_3074,N_1090);
xnor U5570 (N_5570,N_2258,N_882);
xor U5571 (N_5571,N_3660,N_682);
nand U5572 (N_5572,N_3061,N_4965);
xor U5573 (N_5573,N_4481,N_2248);
or U5574 (N_5574,N_3820,N_1183);
or U5575 (N_5575,N_4784,N_166);
xor U5576 (N_5576,N_396,N_3898);
nand U5577 (N_5577,N_4785,N_2500);
nor U5578 (N_5578,N_2299,N_4039);
and U5579 (N_5579,N_1764,N_4977);
or U5580 (N_5580,N_1188,N_4395);
and U5581 (N_5581,N_3026,N_1388);
xnor U5582 (N_5582,N_4243,N_4576);
and U5583 (N_5583,N_960,N_2167);
and U5584 (N_5584,N_3424,N_1005);
xor U5585 (N_5585,N_4691,N_2067);
or U5586 (N_5586,N_52,N_4302);
and U5587 (N_5587,N_1992,N_4830);
nor U5588 (N_5588,N_436,N_4997);
nand U5589 (N_5589,N_99,N_3431);
nor U5590 (N_5590,N_98,N_217);
xnor U5591 (N_5591,N_854,N_4114);
nor U5592 (N_5592,N_4109,N_2724);
or U5593 (N_5593,N_2480,N_4780);
nor U5594 (N_5594,N_320,N_118);
xor U5595 (N_5595,N_4289,N_3098);
xor U5596 (N_5596,N_2584,N_2926);
nand U5597 (N_5597,N_2206,N_2662);
xnor U5598 (N_5598,N_2609,N_3941);
or U5599 (N_5599,N_2807,N_1520);
nand U5600 (N_5600,N_601,N_1554);
nand U5601 (N_5601,N_4438,N_615);
and U5602 (N_5602,N_315,N_1970);
or U5603 (N_5603,N_4249,N_695);
or U5604 (N_5604,N_2025,N_1571);
nand U5605 (N_5605,N_175,N_3965);
and U5606 (N_5606,N_2398,N_2599);
nand U5607 (N_5607,N_1597,N_806);
xnor U5608 (N_5608,N_2073,N_2400);
or U5609 (N_5609,N_874,N_1809);
or U5610 (N_5610,N_3613,N_1327);
nor U5611 (N_5611,N_1161,N_3053);
nand U5612 (N_5612,N_3358,N_2838);
or U5613 (N_5613,N_3134,N_2470);
and U5614 (N_5614,N_3458,N_2121);
or U5615 (N_5615,N_3204,N_4371);
and U5616 (N_5616,N_2134,N_2303);
xor U5617 (N_5617,N_1784,N_888);
and U5618 (N_5618,N_148,N_2131);
and U5619 (N_5619,N_1589,N_1987);
nor U5620 (N_5620,N_4355,N_4073);
and U5621 (N_5621,N_3687,N_4779);
or U5622 (N_5622,N_3357,N_4913);
xor U5623 (N_5623,N_1022,N_3280);
and U5624 (N_5624,N_4324,N_2954);
nand U5625 (N_5625,N_1904,N_1985);
nor U5626 (N_5626,N_1791,N_4044);
nand U5627 (N_5627,N_2714,N_3071);
and U5628 (N_5628,N_2751,N_4882);
nor U5629 (N_5629,N_381,N_3194);
and U5630 (N_5630,N_1013,N_1421);
nand U5631 (N_5631,N_4851,N_903);
or U5632 (N_5632,N_196,N_1883);
nand U5633 (N_5633,N_2782,N_3466);
or U5634 (N_5634,N_4732,N_3540);
nand U5635 (N_5635,N_1846,N_3982);
or U5636 (N_5636,N_4868,N_1569);
xnor U5637 (N_5637,N_2160,N_4311);
nor U5638 (N_5638,N_4742,N_1284);
nor U5639 (N_5639,N_3438,N_1890);
xnor U5640 (N_5640,N_2906,N_4098);
nand U5641 (N_5641,N_3596,N_4781);
nand U5642 (N_5642,N_4493,N_1459);
or U5643 (N_5643,N_2273,N_4974);
and U5644 (N_5644,N_847,N_1920);
and U5645 (N_5645,N_2016,N_4981);
nand U5646 (N_5646,N_1604,N_2703);
or U5647 (N_5647,N_3581,N_2942);
or U5648 (N_5648,N_1586,N_3742);
or U5649 (N_5649,N_4034,N_4357);
nand U5650 (N_5650,N_2731,N_4180);
nand U5651 (N_5651,N_3582,N_819);
or U5652 (N_5652,N_1908,N_3951);
or U5653 (N_5653,N_4695,N_2983);
xor U5654 (N_5654,N_3214,N_971);
or U5655 (N_5655,N_1240,N_1771);
and U5656 (N_5656,N_157,N_2945);
or U5657 (N_5657,N_2456,N_2325);
nand U5658 (N_5658,N_395,N_2292);
nor U5659 (N_5659,N_2740,N_4649);
xor U5660 (N_5660,N_3286,N_3521);
or U5661 (N_5661,N_1900,N_1043);
xor U5662 (N_5662,N_1811,N_559);
nor U5663 (N_5663,N_200,N_668);
nand U5664 (N_5664,N_2483,N_3764);
and U5665 (N_5665,N_222,N_3028);
and U5666 (N_5666,N_3738,N_4804);
nor U5667 (N_5667,N_1737,N_144);
nand U5668 (N_5668,N_291,N_1065);
and U5669 (N_5669,N_597,N_4627);
or U5670 (N_5670,N_3507,N_4794);
xor U5671 (N_5671,N_1757,N_1454);
xor U5672 (N_5672,N_3990,N_1405);
nor U5673 (N_5673,N_3055,N_3937);
or U5674 (N_5674,N_4668,N_4979);
xor U5675 (N_5675,N_1925,N_1907);
or U5676 (N_5676,N_3321,N_747);
or U5677 (N_5677,N_3647,N_3526);
xnor U5678 (N_5678,N_1852,N_598);
and U5679 (N_5679,N_4760,N_1581);
nor U5680 (N_5680,N_2603,N_3669);
nand U5681 (N_5681,N_2009,N_425);
nand U5682 (N_5682,N_60,N_4486);
nor U5683 (N_5683,N_347,N_931);
xor U5684 (N_5684,N_2159,N_4153);
and U5685 (N_5685,N_164,N_1787);
or U5686 (N_5686,N_1305,N_272);
or U5687 (N_5687,N_3163,N_2686);
or U5688 (N_5688,N_1689,N_2725);
nor U5689 (N_5689,N_2844,N_2930);
nor U5690 (N_5690,N_4118,N_2624);
nand U5691 (N_5691,N_4826,N_1982);
nand U5692 (N_5692,N_675,N_3954);
and U5693 (N_5693,N_3778,N_4658);
and U5694 (N_5694,N_4269,N_3133);
nor U5695 (N_5695,N_1215,N_163);
and U5696 (N_5696,N_2804,N_2041);
xnor U5697 (N_5697,N_957,N_4650);
or U5698 (N_5698,N_26,N_3997);
nor U5699 (N_5699,N_669,N_1677);
or U5700 (N_5700,N_2785,N_2307);
xnor U5701 (N_5701,N_772,N_2753);
nand U5702 (N_5702,N_993,N_84);
nor U5703 (N_5703,N_868,N_4329);
or U5704 (N_5704,N_1248,N_3114);
and U5705 (N_5705,N_3808,N_2787);
and U5706 (N_5706,N_3638,N_3460);
and U5707 (N_5707,N_1486,N_4740);
and U5708 (N_5708,N_632,N_2554);
and U5709 (N_5709,N_2994,N_3491);
and U5710 (N_5710,N_3483,N_2762);
and U5711 (N_5711,N_3696,N_4309);
xor U5712 (N_5712,N_1868,N_1475);
nand U5713 (N_5713,N_1451,N_2558);
or U5714 (N_5714,N_1111,N_4883);
nor U5715 (N_5715,N_2447,N_1735);
or U5716 (N_5716,N_873,N_2103);
or U5717 (N_5717,N_3465,N_1057);
or U5718 (N_5718,N_3427,N_4495);
and U5719 (N_5719,N_4801,N_1598);
nand U5720 (N_5720,N_4980,N_2076);
nor U5721 (N_5721,N_213,N_636);
xnor U5722 (N_5722,N_2794,N_4746);
xor U5723 (N_5723,N_663,N_3104);
and U5724 (N_5724,N_4028,N_1626);
nor U5725 (N_5725,N_3713,N_2110);
nand U5726 (N_5726,N_4870,N_1956);
and U5727 (N_5727,N_685,N_2478);
and U5728 (N_5728,N_4800,N_3927);
and U5729 (N_5729,N_2728,N_4654);
nand U5730 (N_5730,N_3776,N_3258);
nor U5731 (N_5731,N_1637,N_2431);
and U5732 (N_5732,N_1076,N_692);
and U5733 (N_5733,N_1329,N_3430);
and U5734 (N_5734,N_4238,N_2551);
or U5735 (N_5735,N_3657,N_4463);
and U5736 (N_5736,N_2501,N_2571);
xnor U5737 (N_5737,N_4286,N_2784);
nor U5738 (N_5738,N_4014,N_4011);
and U5739 (N_5739,N_3278,N_1245);
xnor U5740 (N_5740,N_4623,N_1264);
nor U5741 (N_5741,N_3846,N_1515);
xnor U5742 (N_5742,N_525,N_4564);
nand U5743 (N_5743,N_2976,N_2075);
xor U5744 (N_5744,N_4890,N_2329);
or U5745 (N_5745,N_2848,N_4589);
and U5746 (N_5746,N_1946,N_25);
nor U5747 (N_5747,N_2171,N_588);
and U5748 (N_5748,N_2621,N_4196);
or U5749 (N_5749,N_774,N_3899);
or U5750 (N_5750,N_496,N_2780);
nand U5751 (N_5751,N_3011,N_1789);
xor U5752 (N_5752,N_4284,N_684);
nand U5753 (N_5753,N_470,N_341);
xor U5754 (N_5754,N_2247,N_2452);
and U5755 (N_5755,N_2149,N_2581);
or U5756 (N_5756,N_575,N_2606);
or U5757 (N_5757,N_49,N_1508);
or U5758 (N_5758,N_1374,N_3117);
nand U5759 (N_5759,N_3305,N_2910);
nand U5760 (N_5760,N_3858,N_3968);
nor U5761 (N_5761,N_94,N_3544);
nor U5762 (N_5762,N_4513,N_739);
and U5763 (N_5763,N_2944,N_1247);
nand U5764 (N_5764,N_4667,N_1769);
nand U5765 (N_5765,N_1017,N_4031);
nand U5766 (N_5766,N_1945,N_4325);
xor U5767 (N_5767,N_3800,N_447);
or U5768 (N_5768,N_2039,N_87);
nor U5769 (N_5769,N_3237,N_3584);
and U5770 (N_5770,N_2210,N_2627);
xor U5771 (N_5771,N_2142,N_3184);
and U5772 (N_5772,N_4958,N_1466);
nor U5773 (N_5773,N_3313,N_1469);
and U5774 (N_5774,N_1782,N_1238);
xnor U5775 (N_5775,N_2409,N_1460);
nor U5776 (N_5776,N_1246,N_2138);
xnor U5777 (N_5777,N_4542,N_2045);
xor U5778 (N_5778,N_4067,N_3576);
nand U5779 (N_5779,N_4397,N_3502);
xor U5780 (N_5780,N_2182,N_2949);
or U5781 (N_5781,N_1165,N_3434);
nor U5782 (N_5782,N_2897,N_2642);
xnor U5783 (N_5783,N_2047,N_1961);
or U5784 (N_5784,N_3537,N_954);
nand U5785 (N_5785,N_4186,N_2068);
or U5786 (N_5786,N_3197,N_430);
or U5787 (N_5787,N_2862,N_1094);
xnor U5788 (N_5788,N_561,N_2372);
xnor U5789 (N_5789,N_3699,N_4013);
or U5790 (N_5790,N_392,N_1375);
or U5791 (N_5791,N_964,N_2279);
or U5792 (N_5792,N_4156,N_2765);
xnor U5793 (N_5793,N_393,N_4534);
and U5794 (N_5794,N_984,N_2560);
and U5795 (N_5795,N_3794,N_2383);
xor U5796 (N_5796,N_4455,N_3138);
and U5797 (N_5797,N_2494,N_2688);
nand U5798 (N_5798,N_1449,N_1797);
nand U5799 (N_5799,N_1732,N_4547);
and U5800 (N_5800,N_2629,N_4985);
nor U5801 (N_5801,N_1384,N_2360);
xnor U5802 (N_5802,N_3528,N_1286);
and U5803 (N_5803,N_1827,N_4948);
nand U5804 (N_5804,N_2165,N_1543);
and U5805 (N_5805,N_1172,N_4993);
nand U5806 (N_5806,N_856,N_3243);
nand U5807 (N_5807,N_1004,N_1792);
nor U5808 (N_5808,N_2387,N_4912);
nor U5809 (N_5809,N_2326,N_3912);
and U5810 (N_5810,N_1214,N_3285);
or U5811 (N_5811,N_110,N_528);
nor U5812 (N_5812,N_1798,N_4024);
or U5813 (N_5813,N_2647,N_1923);
xor U5814 (N_5814,N_1813,N_1372);
or U5815 (N_5815,N_14,N_3593);
and U5816 (N_5816,N_4617,N_2670);
and U5817 (N_5817,N_2819,N_274);
nor U5818 (N_5818,N_4020,N_4754);
and U5819 (N_5819,N_2630,N_3643);
and U5820 (N_5820,N_2267,N_3793);
nand U5821 (N_5821,N_2718,N_2768);
or U5822 (N_5822,N_4991,N_1355);
nor U5823 (N_5823,N_4764,N_1008);
and U5824 (N_5824,N_693,N_1609);
or U5825 (N_5825,N_4503,N_664);
nor U5826 (N_5826,N_2552,N_3978);
xor U5827 (N_5827,N_2342,N_4675);
nor U5828 (N_5828,N_1750,N_3281);
xnor U5829 (N_5829,N_4,N_1584);
or U5830 (N_5830,N_2775,N_991);
nor U5831 (N_5831,N_1012,N_2287);
nand U5832 (N_5832,N_78,N_1562);
or U5833 (N_5833,N_4528,N_184);
and U5834 (N_5834,N_2139,N_621);
xnor U5835 (N_5835,N_2874,N_1084);
or U5836 (N_5836,N_4112,N_2060);
or U5837 (N_5837,N_469,N_3991);
xor U5838 (N_5838,N_3435,N_3946);
nand U5839 (N_5839,N_2143,N_2455);
nand U5840 (N_5840,N_4147,N_1224);
or U5841 (N_5841,N_4282,N_526);
nand U5842 (N_5842,N_4632,N_1579);
xnor U5843 (N_5843,N_2386,N_2536);
nor U5844 (N_5844,N_4665,N_966);
and U5845 (N_5845,N_3926,N_587);
or U5846 (N_5846,N_2137,N_505);
xnor U5847 (N_5847,N_4021,N_3473);
and U5848 (N_5848,N_4203,N_2852);
xor U5849 (N_5849,N_1443,N_4837);
and U5850 (N_5850,N_2192,N_2436);
or U5851 (N_5851,N_2374,N_1699);
nor U5852 (N_5852,N_593,N_3510);
or U5853 (N_5853,N_374,N_483);
nor U5854 (N_5854,N_2956,N_3327);
or U5855 (N_5855,N_2189,N_4614);
nand U5856 (N_5856,N_3387,N_2424);
or U5857 (N_5857,N_4624,N_4427);
or U5858 (N_5858,N_3612,N_3212);
or U5859 (N_5859,N_3585,N_2233);
xor U5860 (N_5860,N_2065,N_4182);
nor U5861 (N_5861,N_299,N_3022);
or U5862 (N_5862,N_3361,N_3265);
nand U5863 (N_5863,N_3625,N_943);
or U5864 (N_5864,N_2925,N_4718);
xor U5865 (N_5865,N_742,N_2960);
or U5866 (N_5866,N_797,N_4277);
xor U5867 (N_5867,N_1836,N_3853);
nor U5868 (N_5868,N_3527,N_2767);
nand U5869 (N_5869,N_4502,N_2705);
nor U5870 (N_5870,N_2667,N_2031);
and U5871 (N_5871,N_4856,N_3132);
xnor U5872 (N_5872,N_3994,N_4451);
xor U5873 (N_5873,N_1354,N_2120);
xnor U5874 (N_5874,N_3410,N_3064);
nand U5875 (N_5875,N_1225,N_3877);
nand U5876 (N_5876,N_2681,N_2344);
or U5877 (N_5877,N_3525,N_3538);
nand U5878 (N_5878,N_1446,N_783);
or U5879 (N_5879,N_479,N_1931);
xnor U5880 (N_5880,N_3804,N_4529);
nor U5881 (N_5881,N_3013,N_1200);
xor U5882 (N_5882,N_2397,N_2044);
or U5883 (N_5883,N_1073,N_380);
or U5884 (N_5884,N_3447,N_2058);
or U5885 (N_5885,N_1644,N_640);
and U5886 (N_5886,N_602,N_1709);
or U5887 (N_5887,N_2057,N_2022);
or U5888 (N_5888,N_1255,N_2745);
nand U5889 (N_5889,N_4254,N_3971);
or U5890 (N_5890,N_225,N_4479);
and U5891 (N_5891,N_619,N_197);
nand U5892 (N_5892,N_2141,N_214);
xor U5893 (N_5893,N_4307,N_2291);
xor U5894 (N_5894,N_825,N_317);
or U5895 (N_5895,N_3252,N_3966);
nor U5896 (N_5896,N_752,N_4996);
xnor U5897 (N_5897,N_3388,N_3766);
or U5898 (N_5898,N_4568,N_4217);
and U5899 (N_5899,N_1494,N_1190);
xnor U5900 (N_5900,N_1507,N_2348);
or U5901 (N_5901,N_4953,N_1140);
nor U5902 (N_5902,N_4135,N_4514);
or U5903 (N_5903,N_2691,N_1975);
nand U5904 (N_5904,N_1452,N_475);
and U5905 (N_5905,N_4334,N_278);
xnor U5906 (N_5906,N_294,N_3816);
and U5907 (N_5907,N_2990,N_3605);
or U5908 (N_5908,N_319,N_4183);
nand U5909 (N_5909,N_997,N_2338);
xor U5910 (N_5910,N_4860,N_3219);
or U5911 (N_5911,N_453,N_257);
and U5912 (N_5912,N_1069,N_3618);
and U5913 (N_5913,N_3145,N_3069);
or U5914 (N_5914,N_2132,N_2201);
nor U5915 (N_5915,N_366,N_2384);
nor U5916 (N_5916,N_1348,N_969);
and U5917 (N_5917,N_4879,N_1847);
or U5918 (N_5918,N_2419,N_3048);
or U5919 (N_5919,N_64,N_1721);
xor U5920 (N_5920,N_3645,N_3840);
and U5921 (N_5921,N_2604,N_2922);
and U5922 (N_5922,N_570,N_541);
and U5923 (N_5923,N_653,N_12);
nand U5924 (N_5924,N_2444,N_508);
xnor U5925 (N_5925,N_4670,N_3326);
nand U5926 (N_5926,N_4077,N_2070);
and U5927 (N_5927,N_4376,N_2553);
nand U5928 (N_5928,N_433,N_2212);
or U5929 (N_5929,N_3279,N_635);
nand U5930 (N_5930,N_3574,N_4703);
and U5931 (N_5931,N_3746,N_3176);
or U5932 (N_5932,N_3683,N_4439);
nand U5933 (N_5933,N_4005,N_1417);
or U5934 (N_5934,N_2245,N_23);
and U5935 (N_5935,N_1748,N_990);
and U5936 (N_5936,N_1132,N_2004);
nor U5937 (N_5937,N_4070,N_1269);
nand U5938 (N_5938,N_3490,N_2227);
xnor U5939 (N_5939,N_2842,N_2885);
nand U5940 (N_5940,N_334,N_417);
or U5941 (N_5941,N_4936,N_2727);
or U5942 (N_5942,N_4285,N_4862);
nand U5943 (N_5943,N_4084,N_2485);
nor U5944 (N_5944,N_39,N_3771);
or U5945 (N_5945,N_877,N_4009);
nand U5946 (N_5946,N_1425,N_4105);
or U5947 (N_5947,N_4075,N_963);
or U5948 (N_5948,N_4820,N_1259);
or U5949 (N_5949,N_3177,N_4640);
and U5950 (N_5950,N_2464,N_916);
xnor U5951 (N_5951,N_3030,N_146);
xor U5952 (N_5952,N_3478,N_1839);
or U5953 (N_5953,N_263,N_1669);
or U5954 (N_5954,N_2525,N_2559);
and U5955 (N_5955,N_3637,N_4638);
and U5956 (N_5956,N_1647,N_3977);
nor U5957 (N_5957,N_2908,N_2224);
and U5958 (N_5958,N_1135,N_3642);
nor U5959 (N_5959,N_2119,N_4365);
xor U5960 (N_5960,N_2271,N_788);
and U5961 (N_5961,N_4064,N_2228);
or U5962 (N_5962,N_2907,N_2285);
or U5963 (N_5963,N_2796,N_2433);
and U5964 (N_5964,N_2898,N_865);
or U5965 (N_5965,N_2579,N_2147);
or U5966 (N_5966,N_2823,N_1356);
xor U5967 (N_5967,N_2927,N_614);
or U5968 (N_5968,N_1337,N_3029);
nor U5969 (N_5969,N_2002,N_2389);
nor U5970 (N_5970,N_594,N_4697);
xor U5971 (N_5971,N_3950,N_3754);
nor U5972 (N_5972,N_728,N_688);
nand U5973 (N_5973,N_2023,N_4842);
and U5974 (N_5974,N_4928,N_3288);
or U5975 (N_5975,N_1150,N_4735);
nor U5976 (N_5976,N_219,N_3671);
or U5977 (N_5977,N_1102,N_1244);
or U5978 (N_5978,N_4711,N_1692);
or U5979 (N_5979,N_3733,N_2240);
xor U5980 (N_5980,N_343,N_1632);
nand U5981 (N_5981,N_4914,N_689);
nor U5982 (N_5982,N_1487,N_911);
and U5983 (N_5983,N_2593,N_4663);
and U5984 (N_5984,N_4484,N_3420);
nor U5985 (N_5985,N_1223,N_4350);
nor U5986 (N_5986,N_3913,N_2940);
nor U5987 (N_5987,N_3517,N_2352);
xor U5988 (N_5988,N_1768,N_4641);
xnor U5989 (N_5989,N_85,N_3336);
and U5990 (N_5990,N_3557,N_4442);
and U5991 (N_5991,N_155,N_330);
or U5992 (N_5992,N_2817,N_3137);
nor U5993 (N_5993,N_4412,N_3472);
or U5994 (N_5994,N_2839,N_760);
nor U5995 (N_5995,N_1072,N_1289);
xor U5996 (N_5996,N_345,N_4770);
or U5997 (N_5997,N_1,N_1060);
nand U5998 (N_5998,N_2129,N_958);
nand U5999 (N_5999,N_4875,N_2449);
or U6000 (N_6000,N_418,N_3591);
or U6001 (N_6001,N_462,N_662);
nand U6002 (N_6002,N_2465,N_435);
or U6003 (N_6003,N_4150,N_3398);
nand U6004 (N_6004,N_3099,N_2006);
or U6005 (N_6005,N_2017,N_4776);
nor U6006 (N_6006,N_1535,N_4867);
and U6007 (N_6007,N_4236,N_351);
or U6008 (N_6008,N_402,N_150);
or U6009 (N_6009,N_1557,N_4315);
nor U6010 (N_6010,N_4900,N_2689);
or U6011 (N_6011,N_3661,N_2539);
or U6012 (N_6012,N_3170,N_1155);
nand U6013 (N_6013,N_1497,N_4478);
xor U6014 (N_6014,N_212,N_147);
xnor U6015 (N_6015,N_2364,N_1174);
and U6016 (N_6016,N_3359,N_4206);
xnor U6017 (N_6017,N_750,N_134);
xor U6018 (N_6018,N_4127,N_3077);
xnor U6019 (N_6019,N_807,N_4905);
and U6020 (N_6020,N_2763,N_1471);
xnor U6021 (N_6021,N_4811,N_234);
nand U6022 (N_6022,N_3772,N_3049);
nand U6023 (N_6023,N_457,N_740);
nor U6024 (N_6024,N_773,N_3046);
nand U6025 (N_6025,N_4629,N_2882);
xnor U6026 (N_6026,N_3324,N_2905);
nand U6027 (N_6027,N_30,N_3963);
and U6028 (N_6028,N_572,N_3935);
nor U6029 (N_6029,N_3254,N_4132);
and U6030 (N_6030,N_389,N_658);
nor U6031 (N_6031,N_884,N_4939);
or U6032 (N_6032,N_4423,N_1882);
nor U6033 (N_6033,N_2190,N_810);
and U6034 (N_6034,N_4498,N_4368);
nor U6035 (N_6035,N_3542,N_3423);
and U6036 (N_6036,N_3468,N_549);
nor U6037 (N_6037,N_886,N_1082);
or U6038 (N_6038,N_3995,N_4108);
and U6039 (N_6039,N_4918,N_2498);
xnor U6040 (N_6040,N_2429,N_3710);
or U6041 (N_6041,N_1817,N_4876);
or U6042 (N_6042,N_2355,N_4961);
xor U6043 (N_6043,N_1455,N_2438);
or U6044 (N_6044,N_4578,N_1780);
or U6045 (N_6045,N_4471,N_625);
and U6046 (N_6046,N_4710,N_3788);
and U6047 (N_6047,N_4885,N_3719);
nand U6048 (N_6048,N_1461,N_4933);
and U6049 (N_6049,N_2719,N_4050);
nor U6050 (N_6050,N_4988,N_983);
nor U6051 (N_6051,N_2237,N_88);
xnor U6052 (N_6052,N_4226,N_962);
nor U6053 (N_6053,N_1235,N_288);
or U6054 (N_6054,N_709,N_2490);
or U6055 (N_6055,N_781,N_3734);
xnor U6056 (N_6056,N_1976,N_3653);
nand U6057 (N_6057,N_4737,N_637);
nand U6058 (N_6058,N_4298,N_1530);
or U6059 (N_6059,N_4494,N_1423);
nand U6060 (N_6060,N_104,N_2122);
or U6061 (N_6061,N_612,N_2056);
nand U6062 (N_6062,N_4673,N_565);
nor U6063 (N_6063,N_2200,N_3901);
and U6064 (N_6064,N_899,N_3352);
or U6065 (N_6065,N_3810,N_275);
or U6066 (N_6066,N_4393,N_4940);
xor U6067 (N_6067,N_2808,N_4931);
nand U6068 (N_6068,N_3662,N_3318);
nand U6069 (N_6069,N_2802,N_11);
or U6070 (N_6070,N_1203,N_498);
nor U6071 (N_6071,N_2242,N_1777);
or U6072 (N_6072,N_2029,N_584);
nand U6073 (N_6073,N_500,N_4849);
or U6074 (N_6074,N_4725,N_4755);
nor U6075 (N_6075,N_2337,N_4321);
or U6076 (N_6076,N_3908,N_247);
and U6077 (N_6077,N_509,N_3109);
xnor U6078 (N_6078,N_346,N_3155);
nor U6079 (N_6079,N_3774,N_427);
nor U6080 (N_6080,N_3799,N_4038);
and U6081 (N_6081,N_1350,N_3338);
nor U6082 (N_6082,N_1114,N_1024);
nand U6083 (N_6083,N_1175,N_3700);
or U6084 (N_6084,N_4989,N_3758);
or U6085 (N_6085,N_2583,N_4702);
or U6086 (N_6086,N_313,N_3803);
and U6087 (N_6087,N_3801,N_617);
and U6088 (N_6088,N_3680,N_4889);
and U6089 (N_6089,N_4609,N_4344);
nand U6090 (N_6090,N_3905,N_1482);
nor U6091 (N_6091,N_2035,N_2987);
nor U6092 (N_6092,N_1629,N_3698);
xnor U6093 (N_6093,N_2088,N_1123);
or U6094 (N_6094,N_1523,N_1134);
or U6095 (N_6095,N_2093,N_3715);
xnor U6096 (N_6096,N_4682,N_1092);
or U6097 (N_6097,N_1055,N_1910);
or U6098 (N_6098,N_3781,N_206);
nor U6099 (N_6099,N_2636,N_4262);
or U6100 (N_6100,N_4342,N_2096);
and U6101 (N_6101,N_2652,N_1988);
nor U6102 (N_6102,N_4722,N_1572);
and U6103 (N_6103,N_1199,N_1401);
xor U6104 (N_6104,N_3217,N_3487);
and U6105 (N_6105,N_1653,N_4198);
nor U6106 (N_6106,N_3342,N_1686);
and U6107 (N_6107,N_2020,N_4999);
nor U6108 (N_6108,N_705,N_2079);
nor U6109 (N_6109,N_4778,N_3976);
nand U6110 (N_6110,N_3291,N_563);
or U6111 (N_6111,N_488,N_4333);
or U6112 (N_6112,N_987,N_3697);
nor U6113 (N_6113,N_1630,N_1435);
or U6114 (N_6114,N_4601,N_473);
nand U6115 (N_6115,N_3161,N_1770);
and U6116 (N_6116,N_644,N_920);
nor U6117 (N_6117,N_3319,N_4341);
or U6118 (N_6118,N_2019,N_1484);
nor U6119 (N_6119,N_3334,N_1402);
nand U6120 (N_6120,N_925,N_3731);
or U6121 (N_6121,N_3833,N_3040);
nor U6122 (N_6122,N_922,N_1241);
nor U6123 (N_6123,N_1258,N_3143);
or U6124 (N_6124,N_4969,N_4531);
or U6125 (N_6125,N_2407,N_2876);
nor U6126 (N_6126,N_4854,N_2735);
nand U6127 (N_6127,N_93,N_4758);
nor U6128 (N_6128,N_3973,N_2140);
or U6129 (N_6129,N_180,N_1196);
nor U6130 (N_6130,N_4866,N_2347);
xnor U6131 (N_6131,N_2815,N_1537);
and U6132 (N_6132,N_3730,N_4022);
nor U6133 (N_6133,N_3942,N_1311);
xor U6134 (N_6134,N_2580,N_4106);
or U6135 (N_6135,N_1643,N_4802);
nor U6136 (N_6136,N_1445,N_2466);
nor U6137 (N_6137,N_3130,N_2406);
nand U6138 (N_6138,N_3924,N_463);
and U6139 (N_6139,N_1036,N_1636);
and U6140 (N_6140,N_2414,N_850);
nor U6141 (N_6141,N_2350,N_4090);
xnor U6142 (N_6142,N_318,N_680);
and U6143 (N_6143,N_1924,N_3075);
or U6144 (N_6144,N_136,N_1003);
xnor U6145 (N_6145,N_906,N_1538);
or U6146 (N_6146,N_2845,N_2902);
nor U6147 (N_6147,N_2388,N_3608);
or U6148 (N_6148,N_1066,N_1973);
nand U6149 (N_6149,N_552,N_4789);
nand U6150 (N_6150,N_4347,N_3785);
or U6151 (N_6151,N_4360,N_735);
nor U6152 (N_6152,N_2557,N_1039);
and U6153 (N_6153,N_2266,N_1720);
nand U6154 (N_6154,N_1079,N_700);
nor U6155 (N_6155,N_1411,N_1054);
or U6156 (N_6156,N_718,N_3379);
nand U6157 (N_6157,N_972,N_1496);
and U6158 (N_6158,N_1803,N_4490);
xnor U6159 (N_6159,N_2144,N_19);
xor U6160 (N_6160,N_1773,N_1300);
nand U6161 (N_6161,N_3885,N_481);
xor U6162 (N_6162,N_4398,N_2183);
xor U6163 (N_6163,N_4336,N_3753);
or U6164 (N_6164,N_595,N_2951);
nor U6165 (N_6165,N_455,N_3455);
nor U6166 (N_6166,N_4274,N_4581);
xnor U6167 (N_6167,N_4142,N_1705);
xor U6168 (N_6168,N_4677,N_4299);
nor U6169 (N_6169,N_3198,N_4574);
nand U6170 (N_6170,N_3860,N_2737);
and U6171 (N_6171,N_2367,N_976);
nor U6172 (N_6172,N_397,N_4092);
nand U6173 (N_6173,N_2783,N_2957);
nor U6174 (N_6174,N_4926,N_754);
xnor U6175 (N_6175,N_138,N_4468);
xnor U6176 (N_6176,N_252,N_2672);
xor U6177 (N_6177,N_2412,N_1365);
nor U6178 (N_6178,N_3101,N_2368);
and U6179 (N_6179,N_3451,N_3135);
nor U6180 (N_6180,N_763,N_2760);
xor U6181 (N_6181,N_4817,N_1724);
or U6182 (N_6182,N_2967,N_2432);
or U6183 (N_6183,N_2833,N_303);
xor U6184 (N_6184,N_2366,N_1754);
nor U6185 (N_6185,N_4506,N_929);
xor U6186 (N_6186,N_1422,N_4267);
nand U6187 (N_6187,N_2113,N_4621);
nor U6188 (N_6188,N_4396,N_1317);
xnor U6189 (N_6189,N_2104,N_2931);
xnor U6190 (N_6190,N_941,N_4763);
and U6191 (N_6191,N_4509,N_2639);
nor U6192 (N_6192,N_2633,N_3571);
nor U6193 (N_6193,N_1682,N_881);
nand U6194 (N_6194,N_870,N_3422);
nor U6195 (N_6195,N_1297,N_454);
and U6196 (N_6196,N_3844,N_352);
xor U6197 (N_6197,N_2040,N_1963);
or U6198 (N_6198,N_1660,N_307);
and U6199 (N_6199,N_4646,N_3208);
xor U6200 (N_6200,N_905,N_95);
xnor U6201 (N_6201,N_3242,N_368);
or U6202 (N_6202,N_4272,N_4672);
nor U6203 (N_6203,N_1583,N_2442);
nand U6204 (N_6204,N_1109,N_3839);
and U6205 (N_6205,N_3757,N_2084);
nand U6206 (N_6206,N_4708,N_3006);
or U6207 (N_6207,N_4543,N_2378);
or U6208 (N_6208,N_1275,N_4263);
nor U6209 (N_6209,N_253,N_959);
nor U6210 (N_6210,N_4214,N_1751);
or U6211 (N_6211,N_3429,N_676);
nand U6212 (N_6212,N_4645,N_4964);
nand U6213 (N_6213,N_3234,N_3392);
nand U6214 (N_6214,N_1765,N_2082);
or U6215 (N_6215,N_4081,N_2330);
or U6216 (N_6216,N_4436,N_890);
nand U6217 (N_6217,N_3005,N_2472);
nor U6218 (N_6218,N_1362,N_1919);
nand U6219 (N_6219,N_3169,N_2585);
and U6220 (N_6220,N_3945,N_3599);
or U6221 (N_6221,N_423,N_2788);
nor U6222 (N_6222,N_2173,N_1377);
nand U6223 (N_6223,N_2597,N_2437);
xnor U6224 (N_6224,N_1290,N_4946);
and U6225 (N_6225,N_1901,N_1028);
nand U6226 (N_6226,N_2453,N_2915);
or U6227 (N_6227,N_2257,N_3182);
nand U6228 (N_6228,N_4943,N_3943);
nor U6229 (N_6229,N_2015,N_4612);
xnor U6230 (N_6230,N_2323,N_68);
or U6231 (N_6231,N_4567,N_4491);
xor U6232 (N_6232,N_3207,N_400);
xor U6233 (N_6233,N_2766,N_1564);
nor U6234 (N_6234,N_1217,N_3037);
nand U6235 (N_6235,N_4898,N_2602);
nor U6236 (N_6236,N_1885,N_1472);
xor U6237 (N_6237,N_123,N_3050);
nand U6238 (N_6238,N_1236,N_935);
and U6239 (N_6239,N_1210,N_1967);
or U6240 (N_6240,N_161,N_1448);
nor U6241 (N_6241,N_3394,N_622);
xnor U6242 (N_6242,N_642,N_3178);
or U6243 (N_6243,N_4036,N_1309);
xor U6244 (N_6244,N_3656,N_731);
xnor U6245 (N_6245,N_3228,N_4739);
xnor U6246 (N_6246,N_4364,N_4061);
xnor U6247 (N_6247,N_2451,N_2379);
and U6248 (N_6248,N_429,N_2777);
and U6249 (N_6249,N_4786,N_721);
xor U6250 (N_6250,N_1321,N_3349);
nor U6251 (N_6251,N_4239,N_4113);
or U6252 (N_6252,N_4585,N_3503);
and U6253 (N_6253,N_4154,N_2524);
nand U6254 (N_6254,N_3355,N_3154);
xor U6255 (N_6255,N_2866,N_3817);
or U6256 (N_6256,N_1730,N_892);
xnor U6257 (N_6257,N_2188,N_2790);
nor U6258 (N_6258,N_1093,N_3784);
or U6259 (N_6259,N_4087,N_727);
and U6260 (N_6260,N_746,N_2537);
and U6261 (N_6261,N_816,N_327);
and U6262 (N_6262,N_1231,N_2196);
xor U6263 (N_6263,N_2912,N_2733);
and U6264 (N_6264,N_4666,N_2576);
and U6265 (N_6265,N_520,N_3923);
or U6266 (N_6266,N_2890,N_2778);
nor U6267 (N_6267,N_2754,N_4146);
nand U6268 (N_6268,N_3651,N_4235);
nor U6269 (N_6269,N_2933,N_399);
xor U6270 (N_6270,N_4462,N_512);
nand U6271 (N_6271,N_4095,N_762);
nor U6272 (N_6272,N_3381,N_2867);
nand U6273 (N_6273,N_3879,N_305);
or U6274 (N_6274,N_328,N_3287);
or U6275 (N_6275,N_3385,N_569);
or U6276 (N_6276,N_833,N_2371);
or U6277 (N_6277,N_3045,N_1222);
xnor U6278 (N_6278,N_3828,N_3310);
nand U6279 (N_6279,N_3275,N_1351);
or U6280 (N_6280,N_1144,N_2565);
or U6281 (N_6281,N_456,N_4349);
and U6282 (N_6282,N_4290,N_296);
nand U6283 (N_6283,N_4181,N_1820);
or U6284 (N_6284,N_4566,N_3888);
or U6285 (N_6285,N_4532,N_1208);
and U6286 (N_6286,N_782,N_2717);
nand U6287 (N_6287,N_4873,N_1186);
or U6288 (N_6288,N_1260,N_2484);
nor U6289 (N_6289,N_4798,N_1310);
nor U6290 (N_6290,N_4027,N_3992);
xor U6291 (N_6291,N_2781,N_776);
or U6292 (N_6292,N_3823,N_2300);
and U6293 (N_6293,N_4158,N_4571);
nor U6294 (N_6294,N_2812,N_3436);
nand U6295 (N_6295,N_618,N_2673);
and U6296 (N_6296,N_3790,N_4085);
or U6297 (N_6297,N_1599,N_195);
nor U6298 (N_6298,N_4178,N_373);
xnor U6299 (N_6299,N_631,N_3917);
xnor U6300 (N_6300,N_564,N_2608);
nand U6301 (N_6301,N_1216,N_382);
or U6302 (N_6302,N_489,N_4517);
nor U6303 (N_6303,N_4047,N_652);
and U6304 (N_6304,N_2033,N_2457);
xnor U6305 (N_6305,N_2613,N_982);
nand U6306 (N_6306,N_4487,N_2486);
and U6307 (N_6307,N_2850,N_4787);
xor U6308 (N_6308,N_1840,N_1130);
nand U6309 (N_6309,N_1320,N_4562);
and U6310 (N_6310,N_2198,N_4358);
xor U6311 (N_6311,N_792,N_350);
and U6312 (N_6312,N_4372,N_4749);
nand U6313 (N_6313,N_2542,N_407);
and U6314 (N_6314,N_4399,N_3870);
or U6315 (N_6315,N_1807,N_208);
nor U6316 (N_6316,N_716,N_2443);
nor U6317 (N_6317,N_1860,N_3477);
xnor U6318 (N_6318,N_2739,N_2730);
nor U6319 (N_6319,N_2924,N_1015);
xor U6320 (N_6320,N_4465,N_4209);
or U6321 (N_6321,N_1009,N_975);
or U6322 (N_6322,N_1399,N_2646);
or U6323 (N_6323,N_3859,N_3246);
or U6324 (N_6324,N_1808,N_1539);
nand U6325 (N_6325,N_4983,N_3814);
or U6326 (N_6326,N_4433,N_4300);
and U6327 (N_6327,N_324,N_1616);
xor U6328 (N_6328,N_1326,N_853);
xor U6329 (N_6329,N_1734,N_605);
or U6330 (N_6330,N_2454,N_2774);
xor U6331 (N_6331,N_221,N_4955);
and U6332 (N_6332,N_2801,N_2904);
nor U6333 (N_6333,N_1363,N_2214);
or U6334 (N_6334,N_558,N_1272);
xnor U6335 (N_6335,N_2298,N_3792);
and U6336 (N_6336,N_2254,N_3825);
nand U6337 (N_6337,N_4000,N_1603);
nor U6338 (N_6338,N_141,N_2230);
nor U6339 (N_6339,N_4161,N_1262);
xor U6340 (N_6340,N_408,N_3354);
nor U6341 (N_6341,N_4450,N_3389);
nand U6342 (N_6342,N_1483,N_3206);
nor U6343 (N_6343,N_4406,N_492);
xnor U6344 (N_6344,N_3459,N_131);
and U6345 (N_6345,N_451,N_3587);
nor U6346 (N_6346,N_4271,N_3827);
nand U6347 (N_6347,N_4769,N_74);
nor U6348 (N_6348,N_2108,N_1819);
and U6349 (N_6349,N_3807,N_2365);
xor U6350 (N_6350,N_4454,N_2743);
nor U6351 (N_6351,N_101,N_48);
or U6352 (N_6352,N_1628,N_517);
and U6353 (N_6353,N_2100,N_1407);
and U6354 (N_6354,N_1663,N_3259);
and U6355 (N_6355,N_4407,N_50);
nor U6356 (N_6356,N_2786,N_1548);
nor U6357 (N_6357,N_1058,N_3047);
xor U6358 (N_6358,N_2923,N_4314);
xnor U6359 (N_6359,N_292,N_2066);
nor U6360 (N_6360,N_942,N_4741);
and U6361 (N_6361,N_596,N_2413);
nor U6362 (N_6362,N_4888,N_2050);
and U6363 (N_6363,N_1342,N_2827);
or U6364 (N_6364,N_3223,N_4157);
or U6365 (N_6365,N_3677,N_562);
or U6366 (N_6366,N_623,N_339);
xor U6367 (N_6367,N_9,N_2133);
nand U6368 (N_6368,N_848,N_609);
and U6369 (N_6369,N_4972,N_2736);
or U6370 (N_6370,N_1379,N_1727);
or U6371 (N_6371,N_3166,N_1237);
and U6372 (N_6372,N_316,N_2008);
or U6373 (N_6373,N_302,N_2509);
nand U6374 (N_6374,N_1426,N_2811);
and U6375 (N_6375,N_2209,N_2135);
nor U6376 (N_6376,N_944,N_1056);
nand U6377 (N_6377,N_1145,N_3095);
nor U6378 (N_6378,N_3919,N_2544);
xnor U6379 (N_6379,N_4170,N_3239);
and U6380 (N_6380,N_3032,N_3498);
or U6381 (N_6381,N_4079,N_4204);
nor U6382 (N_6382,N_3479,N_2779);
nor U6383 (N_6383,N_3652,N_671);
or U6384 (N_6384,N_1011,N_28);
nor U6385 (N_6385,N_268,N_3402);
or U6386 (N_6386,N_3514,N_3446);
nor U6387 (N_6387,N_2720,N_1670);
nand U6388 (N_6388,N_1373,N_4545);
and U6389 (N_6389,N_2631,N_62);
nor U6390 (N_6390,N_1220,N_3873);
nand U6391 (N_6391,N_2231,N_4066);
nor U6392 (N_6392,N_4049,N_1657);
or U6393 (N_6393,N_3089,N_486);
nor U6394 (N_6394,N_4642,N_2756);
nor U6395 (N_6395,N_2605,N_2361);
xnor U6396 (N_6396,N_4260,N_4096);
and U6397 (N_6397,N_1683,N_2840);
nand U6398 (N_6398,N_51,N_3512);
or U6399 (N_6399,N_3448,N_3904);
or U6400 (N_6400,N_3283,N_3233);
xor U6401 (N_6401,N_4230,N_2569);
xnor U6402 (N_6402,N_504,N_1887);
and U6403 (N_6403,N_4530,N_4952);
nor U6404 (N_6404,N_2968,N_4558);
nor U6405 (N_6405,N_4535,N_1983);
nor U6406 (N_6406,N_3511,N_1639);
nor U6407 (N_6407,N_1089,N_4591);
nor U6408 (N_6408,N_590,N_1299);
and U6409 (N_6409,N_3534,N_2375);
or U6410 (N_6410,N_2573,N_1713);
nand U6411 (N_6411,N_767,N_3723);
xnor U6412 (N_6412,N_537,N_3616);
and U6413 (N_6413,N_1884,N_1430);
or U6414 (N_6414,N_4738,N_2055);
or U6415 (N_6415,N_3769,N_2148);
xnor U6416 (N_6416,N_3837,N_3809);
and U6417 (N_6417,N_4707,N_2826);
nor U6418 (N_6418,N_3399,N_298);
xnor U6419 (N_6419,N_808,N_2919);
nand U6420 (N_6420,N_372,N_894);
or U6421 (N_6421,N_4139,N_3186);
nand U6422 (N_6422,N_3988,N_1323);
nor U6423 (N_6423,N_461,N_503);
or U6424 (N_6424,N_4730,N_3363);
and U6425 (N_6425,N_1050,N_4611);
and U6426 (N_6426,N_3125,N_409);
and U6427 (N_6427,N_187,N_41);
nand U6428 (N_6428,N_1611,N_3068);
or U6429 (N_6429,N_2855,N_3836);
nor U6430 (N_6430,N_4584,N_690);
xor U6431 (N_6431,N_3717,N_3464);
nand U6432 (N_6432,N_828,N_121);
and U6433 (N_6433,N_3931,N_4743);
xnor U6434 (N_6434,N_1091,N_162);
or U6435 (N_6435,N_2462,N_2395);
and U6436 (N_6436,N_1077,N_3383);
xnor U6437 (N_6437,N_878,N_2961);
nor U6438 (N_6438,N_4363,N_460);
nand U6439 (N_6439,N_3024,N_4793);
and U6440 (N_6440,N_2818,N_1213);
or U6441 (N_6441,N_1127,N_2610);
and U6442 (N_6442,N_1344,N_2311);
xor U6443 (N_6443,N_4496,N_108);
nor U6444 (N_6444,N_2090,N_4383);
and U6445 (N_6445,N_2281,N_4409);
and U6446 (N_6446,N_2793,N_3548);
xor U6447 (N_6447,N_3882,N_1000);
xnor U6448 (N_6448,N_1786,N_1201);
or U6449 (N_6449,N_1892,N_604);
xnor U6450 (N_6450,N_2408,N_2042);
xnor U6451 (N_6451,N_4644,N_2698);
nor U6452 (N_6452,N_1558,N_1211);
and U6453 (N_6453,N_2582,N_3297);
nor U6454 (N_6454,N_1865,N_4553);
or U6455 (N_6455,N_3741,N_3093);
nor U6456 (N_6456,N_4586,N_585);
nand U6457 (N_6457,N_768,N_1661);
xnor U6458 (N_6458,N_1725,N_1897);
or U6459 (N_6459,N_2331,N_840);
xnor U6460 (N_6460,N_1896,N_573);
nand U6461 (N_6461,N_2166,N_342);
xor U6462 (N_6462,N_1138,N_620);
and U6463 (N_6463,N_918,N_720);
nor U6464 (N_6464,N_38,N_1989);
or U6465 (N_6465,N_4825,N_2562);
nand U6466 (N_6466,N_112,N_3891);
or U6467 (N_6467,N_450,N_3791);
or U6468 (N_6468,N_1522,N_77);
and U6469 (N_6469,N_189,N_2864);
and U6470 (N_6470,N_4259,N_3829);
and U6471 (N_6471,N_1854,N_988);
or U6472 (N_6472,N_2591,N_554);
or U6473 (N_6473,N_4941,N_3505);
xnor U6474 (N_6474,N_1525,N_1778);
or U6475 (N_6475,N_3918,N_218);
nor U6476 (N_6476,N_103,N_1293);
xor U6477 (N_6477,N_1361,N_448);
or U6478 (N_6478,N_4278,N_2588);
nand U6479 (N_6479,N_1526,N_3889);
and U6480 (N_6480,N_2164,N_624);
and U6481 (N_6481,N_2280,N_4556);
nand U6482 (N_6482,N_4007,N_4766);
nor U6483 (N_6483,N_1680,N_441);
or U6484 (N_6484,N_2252,N_3721);
nor U6485 (N_6485,N_259,N_678);
or U6486 (N_6486,N_3666,N_1493);
or U6487 (N_6487,N_3335,N_3039);
xor U6488 (N_6488,N_3560,N_1034);
nor U6489 (N_6489,N_1838,N_3142);
nand U6490 (N_6490,N_1257,N_2600);
nor U6491 (N_6491,N_1613,N_1793);
or U6492 (N_6492,N_2676,N_2087);
nor U6493 (N_6493,N_4539,N_3240);
nand U6494 (N_6494,N_2393,N_2973);
and U6495 (N_6495,N_2831,N_4083);
nor U6496 (N_6496,N_1162,N_4322);
nor U6497 (N_6497,N_702,N_1164);
or U6498 (N_6498,N_832,N_1462);
or U6499 (N_6499,N_2805,N_3621);
and U6500 (N_6500,N_2013,N_2286);
xnor U6501 (N_6501,N_1905,N_4008);
and U6502 (N_6502,N_375,N_2037);
or U6503 (N_6503,N_4053,N_3648);
nor U6504 (N_6504,N_1601,N_3887);
or U6505 (N_6505,N_4626,N_4475);
xnor U6506 (N_6506,N_4790,N_3406);
nor U6507 (N_6507,N_3705,N_1335);
xor U6508 (N_6508,N_4057,N_3482);
nand U6509 (N_6509,N_3375,N_1527);
or U6510 (N_6510,N_2411,N_2656);
nor U6511 (N_6511,N_1580,N_276);
and U6512 (N_6512,N_1412,N_2894);
xnor U6513 (N_6513,N_1029,N_1136);
nor U6514 (N_6514,N_2789,N_2376);
nand U6515 (N_6515,N_1075,N_2607);
or U6516 (N_6516,N_3209,N_4622);
nor U6517 (N_6517,N_3617,N_4838);
nand U6518 (N_6518,N_4071,N_1821);
and U6519 (N_6519,N_96,N_286);
nand U6520 (N_6520,N_4982,N_1729);
xor U6521 (N_6521,N_845,N_4511);
nand U6522 (N_6522,N_3440,N_646);
xor U6523 (N_6523,N_579,N_246);
xnor U6524 (N_6524,N_861,N_4456);
nand U6525 (N_6525,N_2643,N_1612);
nor U6526 (N_6526,N_312,N_813);
or U6527 (N_6527,N_4752,N_2211);
and U6528 (N_6528,N_4035,N_3329);
xor U6529 (N_6529,N_4431,N_4346);
nor U6530 (N_6530,N_4227,N_4422);
nand U6531 (N_6531,N_170,N_2261);
xnor U6532 (N_6532,N_371,N_4524);
xor U6533 (N_6533,N_655,N_244);
and U6534 (N_6534,N_4173,N_3248);
nor U6535 (N_6535,N_2531,N_2515);
nor U6536 (N_6536,N_4674,N_177);
xor U6537 (N_6537,N_4625,N_4744);
or U6538 (N_6538,N_2711,N_1620);
xor U6539 (N_6539,N_3589,N_3162);
nor U6540 (N_6540,N_336,N_4869);
nand U6541 (N_6541,N_2979,N_3770);
xor U6542 (N_6542,N_3881,N_3925);
or U6543 (N_6543,N_4320,N_979);
nand U6544 (N_6544,N_4103,N_262);
or U6545 (N_6545,N_1921,N_4492);
nand U6546 (N_6546,N_4069,N_2632);
xnor U6547 (N_6547,N_4078,N_4886);
xor U6548 (N_6548,N_751,N_137);
nor U6549 (N_6549,N_3340,N_981);
nand U6550 (N_6550,N_3113,N_1083);
nor U6551 (N_6551,N_2878,N_2161);
or U6552 (N_6552,N_3292,N_1424);
or U6553 (N_6553,N_4930,N_3232);
nor U6554 (N_6554,N_2396,N_2063);
xnor U6555 (N_6555,N_80,N_443);
nand U6556 (N_6556,N_2946,N_2263);
and U6557 (N_6557,N_3577,N_56);
or U6558 (N_6558,N_3384,N_3644);
and U6559 (N_6559,N_1227,N_3701);
xnor U6560 (N_6560,N_2000,N_4756);
and U6561 (N_6561,N_1758,N_2545);
nand U6562 (N_6562,N_1590,N_4560);
nor U6563 (N_6563,N_4987,N_193);
nand U6564 (N_6564,N_506,N_4602);
nand U6565 (N_6565,N_3520,N_4809);
nor U6566 (N_6566,N_204,N_178);
nand U6567 (N_6567,N_2324,N_432);
nor U6568 (N_6568,N_2255,N_706);
or U6569 (N_6569,N_4590,N_4125);
nor U6570 (N_6570,N_2959,N_424);
and U6571 (N_6571,N_1857,N_1059);
and U6572 (N_6572,N_2313,N_2046);
xnor U6573 (N_6573,N_613,N_3722);
xor U6574 (N_6574,N_4653,N_1152);
or U6575 (N_6575,N_4901,N_1042);
nor U6576 (N_6576,N_1117,N_1950);
xnor U6577 (N_6577,N_2332,N_1783);
xnor U6578 (N_6578,N_449,N_610);
nor U6579 (N_6579,N_2797,N_4605);
nand U6580 (N_6580,N_4777,N_4331);
xnor U6581 (N_6581,N_1185,N_1250);
nor U6582 (N_6582,N_3501,N_3128);
nand U6583 (N_6583,N_4187,N_4935);
and U6584 (N_6584,N_2556,N_434);
xor U6585 (N_6585,N_3457,N_3654);
nor U6586 (N_6586,N_4694,N_1849);
nand U6587 (N_6587,N_1020,N_4635);
xnor U6588 (N_6588,N_4233,N_4116);
or U6589 (N_6589,N_730,N_803);
nor U6590 (N_6590,N_2181,N_3195);
and U6591 (N_6591,N_4384,N_4119);
and U6592 (N_6592,N_2404,N_1331);
xnor U6593 (N_6593,N_4121,N_626);
nor U6594 (N_6594,N_2975,N_3059);
nor U6595 (N_6595,N_897,N_4910);
and U6596 (N_6596,N_1045,N_3372);
or U6597 (N_6597,N_4726,N_309);
or U6598 (N_6598,N_2538,N_2939);
nand U6599 (N_6599,N_629,N_1654);
or U6600 (N_6600,N_2203,N_4546);
nand U6601 (N_6601,N_949,N_3848);
nor U6602 (N_6602,N_4459,N_3513);
xnor U6603 (N_6603,N_4126,N_817);
xnor U6604 (N_6604,N_3953,N_2700);
xor U6605 (N_6605,N_1119,N_1478);
and U6606 (N_6606,N_1981,N_1761);
xor U6607 (N_6607,N_1739,N_1509);
xor U6608 (N_6608,N_127,N_3916);
xnor U6609 (N_6609,N_1851,N_1848);
and U6610 (N_6610,N_697,N_2178);
nand U6611 (N_6611,N_1575,N_4029);
or U6612 (N_6612,N_4819,N_4222);
nand U6613 (N_6613,N_1202,N_1181);
nor U6614 (N_6614,N_4728,N_532);
nand U6615 (N_6615,N_4184,N_4201);
nand U6616 (N_6616,N_523,N_1756);
nand U6617 (N_6617,N_1124,N_3052);
nand U6618 (N_6618,N_3831,N_2471);
xnor U6619 (N_6619,N_1182,N_893);
xor U6620 (N_6620,N_2869,N_4356);
nand U6621 (N_6621,N_4580,N_3740);
nor U6622 (N_6622,N_4500,N_908);
nor U6623 (N_6623,N_3216,N_3396);
or U6624 (N_6624,N_3813,N_551);
nor U6625 (N_6625,N_4390,N_4655);
xor U6626 (N_6626,N_1556,N_1352);
xnor U6627 (N_6627,N_3025,N_4782);
nor U6628 (N_6628,N_2488,N_1110);
and U6629 (N_6629,N_4934,N_3962);
nor U6630 (N_6630,N_4059,N_4483);
nand U6631 (N_6631,N_2169,N_3080);
or U6632 (N_6632,N_3332,N_2535);
nand U6633 (N_6633,N_3568,N_4256);
nor U6634 (N_6634,N_1567,N_2128);
or U6635 (N_6635,N_4923,N_2622);
xnor U6636 (N_6636,N_566,N_2764);
or U6637 (N_6637,N_2649,N_3597);
or U6638 (N_6638,N_3735,N_1280);
and U6639 (N_6639,N_3729,N_3961);
or U6640 (N_6640,N_491,N_4287);
nor U6641 (N_6641,N_4037,N_1810);
and U6642 (N_6642,N_4306,N_2858);
xor U6643 (N_6643,N_3909,N_934);
or U6644 (N_6644,N_4074,N_2213);
and U6645 (N_6645,N_608,N_384);
xor U6646 (N_6646,N_2628,N_3179);
nand U6647 (N_6647,N_3078,N_3682);
xor U6648 (N_6648,N_1984,N_1623);
nand U6649 (N_6649,N_4003,N_3443);
xnor U6650 (N_6650,N_171,N_603);
xnor U6651 (N_6651,N_3337,N_3076);
nor U6652 (N_6652,N_1801,N_1621);
nor U6653 (N_6653,N_3579,N_4821);
or U6654 (N_6654,N_4911,N_1400);
or U6655 (N_6655,N_2085,N_3640);
or U6656 (N_6656,N_4504,N_287);
nand U6657 (N_6657,N_2199,N_896);
and U6658 (N_6658,N_2032,N_2401);
and U6659 (N_6659,N_3634,N_4903);
nor U6660 (N_6660,N_4434,N_3255);
or U6661 (N_6661,N_1602,N_1832);
or U6662 (N_6662,N_2877,N_1678);
and U6663 (N_6663,N_2716,N_3404);
or U6664 (N_6664,N_786,N_132);
and U6665 (N_6665,N_4771,N_530);
xnor U6666 (N_6666,N_4387,N_3180);
nor U6667 (N_6667,N_2474,N_2154);
nor U6668 (N_6668,N_40,N_388);
and U6669 (N_6669,N_3759,N_2821);
or U6670 (N_6670,N_367,N_3678);
and U6671 (N_6671,N_4945,N_183);
xnor U6672 (N_6672,N_670,N_2101);
and U6673 (N_6673,N_2750,N_4056);
nor U6674 (N_6674,N_1368,N_65);
or U6675 (N_6675,N_535,N_533);
or U6676 (N_6676,N_996,N_2460);
xnor U6677 (N_6677,N_2543,N_545);
nor U6678 (N_6678,N_2938,N_3980);
nor U6679 (N_6679,N_3865,N_3583);
nor U6680 (N_6680,N_3126,N_2601);
and U6681 (N_6681,N_759,N_4995);
nor U6682 (N_6682,N_1814,N_2638);
nor U6683 (N_6683,N_4829,N_2914);
or U6684 (N_6684,N_4414,N_3345);
nand U6685 (N_6685,N_2074,N_1345);
and U6686 (N_6686,N_45,N_3226);
nor U6687 (N_6687,N_1406,N_139);
nand U6688 (N_6688,N_79,N_4197);
and U6689 (N_6689,N_1804,N_1383);
xor U6690 (N_6690,N_4143,N_2270);
and U6691 (N_6691,N_4970,N_3085);
and U6692 (N_6692,N_3213,N_3824);
or U6693 (N_6693,N_2441,N_3668);
xor U6694 (N_6694,N_1658,N_3554);
and U6695 (N_6695,N_2887,N_3635);
nor U6696 (N_6696,N_1911,N_2130);
nor U6697 (N_6697,N_2162,N_4685);
nand U6698 (N_6698,N_683,N_502);
or U6699 (N_6699,N_3749,N_3933);
nor U6700 (N_6700,N_3704,N_3611);
or U6701 (N_6701,N_4305,N_3928);
or U6702 (N_6702,N_2872,N_2034);
xor U6703 (N_6703,N_152,N_4844);
nor U6704 (N_6704,N_281,N_1282);
xor U6705 (N_6705,N_2982,N_3151);
nand U6706 (N_6706,N_4208,N_3782);
nand U6707 (N_6707,N_2816,N_3762);
and U6708 (N_6708,N_580,N_2392);
or U6709 (N_6709,N_4473,N_3667);
nor U6710 (N_6710,N_3317,N_348);
nor U6711 (N_6711,N_4094,N_1872);
xor U6712 (N_6712,N_2568,N_223);
and U6713 (N_6713,N_701,N_1061);
or U6714 (N_6714,N_4062,N_1659);
nor U6715 (N_6715,N_4152,N_4944);
or U6716 (N_6716,N_1607,N_233);
nor U6717 (N_6717,N_1364,N_4693);
or U6718 (N_6718,N_129,N_4927);
or U6719 (N_6719,N_29,N_215);
and U6720 (N_6720,N_1314,N_33);
and U6721 (N_6721,N_4218,N_1948);
or U6722 (N_6722,N_97,N_1191);
or U6723 (N_6723,N_4017,N_1568);
xor U6724 (N_6724,N_2069,N_4216);
or U6725 (N_6725,N_3996,N_2320);
or U6726 (N_6726,N_4592,N_4231);
nand U6727 (N_6727,N_3598,N_1917);
nand U6728 (N_6728,N_723,N_156);
nand U6729 (N_6729,N_4748,N_4845);
nand U6730 (N_6730,N_3304,N_1853);
nand U6731 (N_6731,N_3494,N_4968);
nand U6732 (N_6732,N_4855,N_794);
nand U6733 (N_6733,N_1154,N_582);
nand U6734 (N_6734,N_2701,N_1447);
or U6735 (N_6735,N_1018,N_1251);
or U6736 (N_6736,N_3884,N_1649);
or U6737 (N_6737,N_1553,N_1489);
and U6738 (N_6738,N_1341,N_4745);
xnor U6739 (N_6739,N_1197,N_329);
or U6740 (N_6740,N_789,N_2729);
nand U6741 (N_6741,N_900,N_3869);
nor U6742 (N_6742,N_1436,N_2903);
or U6743 (N_6743,N_1288,N_2830);
and U6744 (N_6744,N_4921,N_1030);
xor U6745 (N_6745,N_4907,N_3732);
and U6746 (N_6746,N_160,N_1476);
nor U6747 (N_6747,N_2502,N_4922);
xor U6748 (N_6748,N_3830,N_4317);
or U6749 (N_6749,N_4555,N_4370);
nor U6750 (N_6750,N_2625,N_831);
and U6751 (N_6751,N_3718,N_4593);
nand U6752 (N_6752,N_2540,N_279);
or U6753 (N_6753,N_4460,N_413);
and U6754 (N_6754,N_1016,N_1794);
or U6755 (N_6755,N_1700,N_1465);
xnor U6756 (N_6756,N_2776,N_1002);
and U6757 (N_6757,N_3168,N_15);
and U6758 (N_6758,N_482,N_4942);
xnor U6759 (N_6759,N_1995,N_2156);
and U6760 (N_6760,N_485,N_2659);
nor U6761 (N_6761,N_4947,N_4177);
or U6762 (N_6762,N_3270,N_3555);
or U6763 (N_6763,N_2493,N_980);
nor U6764 (N_6764,N_2308,N_801);
nor U6765 (N_6765,N_1816,N_4823);
and U6766 (N_6766,N_2012,N_4296);
or U6767 (N_6767,N_1021,N_3314);
and U6768 (N_6768,N_113,N_265);
and U6769 (N_6769,N_1395,N_578);
and U6770 (N_6770,N_2399,N_59);
nor U6771 (N_6771,N_2534,N_2713);
nor U6772 (N_6772,N_4168,N_3153);
nor U6773 (N_6773,N_4799,N_1781);
xor U6774 (N_6774,N_3027,N_3789);
xor U6775 (N_6775,N_1437,N_4660);
and U6776 (N_6776,N_3572,N_4919);
nor U6777 (N_6777,N_3461,N_420);
nor U6778 (N_6778,N_3426,N_2503);
nor U6779 (N_6779,N_1371,N_1834);
or U6780 (N_6780,N_83,N_4080);
xor U6781 (N_6781,N_3957,N_1146);
nand U6782 (N_6782,N_3561,N_1014);
xor U6783 (N_6783,N_1665,N_2126);
xnor U6784 (N_6784,N_471,N_1131);
xor U6785 (N_6785,N_1824,N_2102);
or U6786 (N_6786,N_495,N_2334);
xnor U6787 (N_6787,N_2992,N_4446);
xor U6788 (N_6788,N_3892,N_1404);
or U6789 (N_6789,N_4724,N_666);
and U6790 (N_6790,N_1726,N_3189);
nor U6791 (N_6791,N_2410,N_2792);
xnor U6792 (N_6792,N_4575,N_4684);
nor U6793 (N_6793,N_639,N_2155);
or U6794 (N_6794,N_1007,N_10);
or U6795 (N_6795,N_1815,N_314);
or U6796 (N_6796,N_1467,N_4554);
and U6797 (N_6797,N_3630,N_4647);
nand U6798 (N_6798,N_4215,N_2315);
nand U6799 (N_6799,N_2422,N_651);
nor U6800 (N_6800,N_2984,N_4388);
and U6801 (N_6801,N_2094,N_2219);
nor U6802 (N_6802,N_2309,N_1474);
or U6803 (N_6803,N_4843,N_172);
nor U6804 (N_6804,N_3041,N_1495);
xnor U6805 (N_6805,N_2574,N_2654);
xor U6806 (N_6806,N_58,N_3998);
and U6807 (N_6807,N_711,N_2690);
nor U6808 (N_6808,N_3008,N_1752);
or U6809 (N_6809,N_2970,N_1394);
xor U6810 (N_6810,N_3989,N_1473);
nand U6811 (N_6811,N_862,N_1625);
or U6812 (N_6812,N_820,N_4570);
nor U6813 (N_6813,N_1218,N_3676);
nand U6814 (N_6814,N_1108,N_928);
nor U6815 (N_6815,N_1071,N_744);
nor U6816 (N_6816,N_2244,N_1541);
nand U6817 (N_6817,N_1980,N_2043);
or U6818 (N_6818,N_930,N_4698);
xnor U6819 (N_6819,N_4193,N_4957);
nand U6820 (N_6820,N_2589,N_3365);
nor U6821 (N_6821,N_2522,N_3607);
or U6822 (N_6822,N_4291,N_2117);
nand U6823 (N_6823,N_887,N_1999);
or U6824 (N_6824,N_756,N_2955);
nand U6825 (N_6825,N_2277,N_1863);
and U6826 (N_6826,N_1633,N_467);
nand U6827 (N_6827,N_3185,N_2092);
nand U6828 (N_6828,N_1744,N_3970);
and U6829 (N_6829,N_3271,N_3541);
nor U6830 (N_6830,N_1147,N_1233);
xor U6831 (N_6831,N_977,N_839);
or U6832 (N_6832,N_1563,N_3508);
and U6833 (N_6833,N_645,N_4352);
nand U6834 (N_6834,N_1551,N_188);
nor U6835 (N_6835,N_3610,N_254);
xnor U6836 (N_6836,N_100,N_4310);
and U6837 (N_6837,N_4573,N_3414);
nand U6838 (N_6838,N_261,N_198);
xnor U6839 (N_6839,N_3570,N_4839);
nor U6840 (N_6840,N_3193,N_3188);
nor U6841 (N_6841,N_2061,N_3229);
nor U6842 (N_6842,N_3350,N_4727);
nor U6843 (N_6843,N_891,N_1359);
nor U6844 (N_6844,N_192,N_4430);
or U6845 (N_6845,N_1850,N_3703);
xor U6846 (N_6846,N_687,N_3262);
xor U6847 (N_6847,N_4379,N_1206);
nor U6848 (N_6848,N_1049,N_784);
xor U6849 (N_6849,N_3854,N_3929);
nand U6850 (N_6850,N_2870,N_713);
and U6851 (N_6851,N_2327,N_2028);
and U6852 (N_6852,N_3606,N_4474);
or U6853 (N_6853,N_855,N_165);
xnor U6854 (N_6854,N_2468,N_4950);
nand U6855 (N_6855,N_1844,N_1396);
or U6856 (N_6856,N_860,N_2520);
or U6857 (N_6857,N_1189,N_560);
and U6858 (N_6858,N_2997,N_3623);
xor U6859 (N_6859,N_3981,N_1353);
nor U6860 (N_6860,N_228,N_4713);
nand U6861 (N_6861,N_4762,N_4242);
xor U6862 (N_6862,N_3914,N_2623);
nor U6863 (N_6863,N_3244,N_2587);
nor U6864 (N_6864,N_1719,N_322);
and U6865 (N_6865,N_4561,N_1914);
xnor U6866 (N_6866,N_4709,N_3818);
nand U6867 (N_6867,N_1268,N_3373);
nand U6868 (N_6868,N_872,N_1170);
xnor U6869 (N_6869,N_4225,N_3665);
and U6870 (N_6870,N_2062,N_770);
or U6871 (N_6871,N_1480,N_703);
nand U6872 (N_6872,N_1697,N_452);
and U6873 (N_6873,N_4651,N_4248);
and U6874 (N_6874,N_4323,N_2889);
nand U6875 (N_6875,N_2518,N_1922);
or U6876 (N_6876,N_3043,N_73);
and U6877 (N_6877,N_3382,N_2508);
or U6878 (N_6878,N_4681,N_4213);
or U6879 (N_6879,N_377,N_1346);
and U6880 (N_6880,N_3556,N_2677);
nand U6881 (N_6881,N_3264,N_3227);
xor U6882 (N_6882,N_3122,N_3573);
nand U6883 (N_6883,N_4240,N_2380);
xnor U6884 (N_6884,N_726,N_3433);
nand U6885 (N_6885,N_2746,N_4816);
or U6886 (N_6886,N_2917,N_2528);
and U6887 (N_6887,N_4615,N_4664);
and U6888 (N_6888,N_2428,N_1828);
nand U6889 (N_6889,N_2820,N_2723);
or U6890 (N_6890,N_3958,N_4416);
or U6891 (N_6891,N_1608,N_2370);
nor U6892 (N_6892,N_3761,N_2482);
xnor U6893 (N_6893,N_2871,N_4765);
nor U6894 (N_6894,N_3974,N_2664);
or U6895 (N_6895,N_3535,N_1151);
and U6896 (N_6896,N_542,N_416);
nor U6897 (N_6897,N_3603,N_2861);
nand U6898 (N_6898,N_3205,N_4878);
or U6899 (N_6899,N_1862,N_4444);
or U6900 (N_6900,N_1067,N_2418);
nor U6901 (N_6901,N_226,N_1731);
nor U6902 (N_6902,N_3852,N_4984);
or U6903 (N_6903,N_2274,N_2194);
nand U6904 (N_6904,N_4279,N_3347);
nand U6905 (N_6905,N_4616,N_3755);
and U6906 (N_6906,N_282,N_3120);
nand U6907 (N_6907,N_4420,N_2304);
and U6908 (N_6908,N_1676,N_771);
xnor U6909 (N_6909,N_951,N_1708);
xnor U6910 (N_6910,N_3516,N_799);
xnor U6911 (N_6911,N_2256,N_883);
xor U6912 (N_6912,N_1051,N_556);
or U6913 (N_6913,N_787,N_3504);
nor U6914 (N_6914,N_1380,N_2322);
and U6915 (N_6915,N_2369,N_3299);
xnor U6916 (N_6916,N_4389,N_1528);
or U6917 (N_6917,N_2657,N_1318);
nor U6918 (N_6918,N_3707,N_4207);
or U6919 (N_6919,N_1044,N_4160);
nor U6920 (N_6920,N_4404,N_3211);
nor U6921 (N_6921,N_3417,N_2218);
xor U6922 (N_6922,N_1941,N_4505);
xnor U6923 (N_6923,N_4172,N_3691);
xnor U6924 (N_6924,N_2699,N_511);
or U6925 (N_6925,N_3118,N_4124);
or U6926 (N_6926,N_766,N_4696);
or U6927 (N_6927,N_4489,N_4452);
nand U6928 (N_6928,N_2405,N_358);
xnor U6929 (N_6929,N_3737,N_1864);
and U6930 (N_6930,N_431,N_3649);
nor U6931 (N_6931,N_1035,N_2995);
and U6932 (N_6932,N_3692,N_3044);
xnor U6933 (N_6933,N_2052,N_1242);
xnor U6934 (N_6934,N_3456,N_3684);
xor U6935 (N_6935,N_2798,N_1648);
nor U6936 (N_6936,N_879,N_337);
xor U6937 (N_6937,N_834,N_4091);
xnor U6938 (N_6938,N_4480,N_3273);
and U6939 (N_6939,N_4223,N_61);
or U6940 (N_6940,N_3139,N_4633);
xnor U6941 (N_6941,N_4775,N_4189);
nor U6942 (N_6942,N_1957,N_1088);
xor U6943 (N_6943,N_1805,N_3857);
or U6944 (N_6944,N_2829,N_4519);
nand U6945 (N_6945,N_4375,N_4891);
nor U6946 (N_6946,N_1845,N_2007);
or U6947 (N_6947,N_3549,N_4613);
nand U6948 (N_6948,N_2879,N_1939);
and U6949 (N_6949,N_4191,N_3405);
or U6950 (N_6950,N_3129,N_2674);
nor U6951 (N_6951,N_3150,N_4729);
and U6952 (N_6952,N_2077,N_2980);
nand U6953 (N_6953,N_2116,N_4810);
and U6954 (N_6954,N_4540,N_1760);
and U6955 (N_6955,N_1640,N_3547);
xnor U6956 (N_6956,N_301,N_2566);
xor U6957 (N_6957,N_1313,N_777);
nand U6958 (N_6958,N_269,N_201);
xor U6959 (N_6959,N_3509,N_3545);
nor U6960 (N_6960,N_344,N_116);
xnor U6961 (N_6961,N_1287,N_1942);
nand U6962 (N_6962,N_3432,N_4421);
xnor U6963 (N_6963,N_3250,N_1038);
nand U6964 (N_6964,N_3726,N_2514);
xor U6965 (N_6965,N_1918,N_2687);
nand U6966 (N_6966,N_4992,N_4268);
and U6967 (N_6967,N_1877,N_3376);
and U6968 (N_6968,N_3474,N_6);
nor U6969 (N_6969,N_1095,N_748);
and U6970 (N_6970,N_2865,N_4264);
xor U6971 (N_6971,N_4508,N_3795);
nor U6972 (N_6972,N_2260,N_1500);
and U6973 (N_6973,N_1673,N_3296);
nand U6974 (N_6974,N_1239,N_1651);
nor U6975 (N_6975,N_4120,N_410);
xor U6976 (N_6976,N_1902,N_1866);
or U6977 (N_6977,N_1723,N_1570);
nor U6978 (N_6978,N_2988,N_2586);
nand U6979 (N_6979,N_3344,N_3416);
and U6980 (N_6980,N_4045,N_4137);
and U6981 (N_6981,N_2394,N_2112);
or U6982 (N_6982,N_4619,N_946);
nor U6983 (N_6983,N_4712,N_3594);
xnor U6984 (N_6984,N_1711,N_3867);
nor U6985 (N_6985,N_1427,N_2174);
nand U6986 (N_6986,N_2339,N_2220);
xor U6987 (N_6987,N_4864,N_656);
nand U6988 (N_6988,N_3485,N_354);
and U6989 (N_6989,N_3341,N_1506);
nor U6990 (N_6990,N_2969,N_2618);
and U6991 (N_6991,N_4101,N_2620);
nor U6992 (N_6992,N_576,N_1799);
nor U6993 (N_6993,N_627,N_1588);
xnor U6994 (N_6994,N_674,N_398);
nor U6995 (N_6995,N_2928,N_3311);
nor U6996 (N_6996,N_2972,N_3670);
and U6997 (N_6997,N_992,N_1631);
nor U6998 (N_6998,N_1867,N_3551);
nor U6999 (N_6999,N_1585,N_1835);
and U7000 (N_7000,N_769,N_1674);
and U7001 (N_7001,N_732,N_117);
nand U7002 (N_7002,N_2469,N_1295);
nand U7003 (N_7003,N_4533,N_1128);
xnor U7004 (N_7004,N_2402,N_349);
xnor U7005 (N_7005,N_1627,N_3855);
nor U7006 (N_7006,N_4659,N_3241);
and U7007 (N_7007,N_1434,N_2641);
xnor U7008 (N_7008,N_3949,N_1112);
nand U7009 (N_7009,N_4734,N_4857);
and U7010 (N_7010,N_3018,N_2901);
nand U7011 (N_7011,N_1605,N_1265);
nor U7012 (N_7012,N_1441,N_2239);
xor U7013 (N_7013,N_1870,N_600);
nand U7014 (N_7014,N_1889,N_3499);
xor U7015 (N_7015,N_923,N_3675);
and U7016 (N_7016,N_1559,N_3063);
nor U7017 (N_7017,N_245,N_1953);
or U7018 (N_7018,N_2269,N_2748);
or U7019 (N_7019,N_476,N_4720);
nor U7020 (N_7020,N_1701,N_1414);
and U7021 (N_7021,N_3626,N_586);
and U7022 (N_7022,N_472,N_2947);
nand U7023 (N_7023,N_1277,N_2710);
or U7024 (N_7024,N_4657,N_857);
nor U7025 (N_7025,N_4194,N_4366);
or U7026 (N_7026,N_1192,N_1226);
nand U7027 (N_7027,N_4425,N_3872);
nand U7028 (N_7028,N_1652,N_2450);
nand U7029 (N_7029,N_2799,N_2170);
and U7030 (N_7030,N_3309,N_4165);
nand U7031 (N_7031,N_3896,N_2682);
and U7032 (N_7032,N_3330,N_1085);
or U7033 (N_7033,N_2351,N_1614);
and U7034 (N_7034,N_2770,N_63);
or U7035 (N_7035,N_4881,N_1859);
or U7036 (N_7036,N_4250,N_2806);
and U7037 (N_7037,N_4679,N_4924);
xor U7038 (N_7038,N_912,N_4902);
nand U7039 (N_7039,N_3263,N_4865);
and U7040 (N_7040,N_2721,N_3136);
xor U7041 (N_7041,N_2822,N_2835);
nand U7042 (N_7042,N_4164,N_616);
nor U7043 (N_7043,N_2843,N_2284);
or U7044 (N_7044,N_2235,N_4340);
or U7045 (N_7045,N_1312,N_82);
nand U7046 (N_7046,N_1516,N_4841);
and U7047 (N_7047,N_1273,N_2693);
nand U7048 (N_7048,N_2773,N_3056);
or U7049 (N_7049,N_439,N_4417);
xor U7050 (N_7050,N_2541,N_3938);
or U7051 (N_7051,N_2752,N_1715);
nor U7052 (N_7052,N_4253,N_3144);
or U7053 (N_7053,N_1157,N_133);
and U7054 (N_7054,N_1103,N_1837);
or U7055 (N_7055,N_4686,N_1428);
and U7056 (N_7056,N_722,N_378);
nor U7057 (N_7057,N_1898,N_376);
or U7058 (N_7058,N_419,N_2377);
and U7059 (N_7059,N_2,N_369);
nor U7060 (N_7060,N_3148,N_973);
or U7061 (N_7061,N_2755,N_3969);
nand U7062 (N_7062,N_4232,N_2205);
or U7063 (N_7063,N_3805,N_1746);
xor U7064 (N_7064,N_290,N_2492);
or U7065 (N_7065,N_895,N_361);
or U7066 (N_7066,N_1544,N_4400);
nand U7067 (N_7067,N_3119,N_1171);
nand U7068 (N_7068,N_3418,N_404);
or U7069 (N_7069,N_2758,N_2276);
and U7070 (N_7070,N_1972,N_1340);
or U7071 (N_7071,N_938,N_3210);
or U7072 (N_7072,N_4715,N_3708);
nor U7073 (N_7073,N_1826,N_5);
nor U7074 (N_7074,N_1298,N_780);
xor U7075 (N_7075,N_3301,N_3566);
nor U7076 (N_7076,N_4956,N_1453);
and U7077 (N_7077,N_4461,N_16);
or U7078 (N_7078,N_4210,N_194);
or U7079 (N_7079,N_1722,N_67);
xnor U7080 (N_7080,N_4058,N_91);
nand U7081 (N_7081,N_2791,N_970);
xor U7082 (N_7082,N_3530,N_2127);
xor U7083 (N_7083,N_422,N_1978);
nor U7084 (N_7084,N_2086,N_4840);
nor U7085 (N_7085,N_1463,N_3452);
and U7086 (N_7086,N_1158,N_1561);
or U7087 (N_7087,N_654,N_105);
or U7088 (N_7088,N_3850,N_3261);
nor U7089 (N_7089,N_1184,N_3021);
and U7090 (N_7090,N_950,N_2880);
nand U7091 (N_7091,N_1940,N_4229);
nand U7092 (N_7092,N_3356,N_3033);
and U7093 (N_7093,N_4850,N_2547);
xor U7094 (N_7094,N_190,N_2888);
and U7095 (N_7095,N_3066,N_1339);
nor U7096 (N_7096,N_830,N_1593);
xnor U7097 (N_7097,N_1958,N_3421);
nand U7098 (N_7098,N_2530,N_2293);
nor U7099 (N_7099,N_2668,N_2197);
and U7100 (N_7100,N_3320,N_1113);
xnor U7101 (N_7101,N_2038,N_2570);
or U7102 (N_7102,N_985,N_3260);
nor U7103 (N_7103,N_3366,N_229);
or U7104 (N_7104,N_3564,N_3051);
xnor U7105 (N_7105,N_4378,N_220);
and U7106 (N_7106,N_3890,N_3486);
nor U7107 (N_7107,N_4155,N_4117);
nor U7108 (N_7108,N_2660,N_4959);
xnor U7109 (N_7109,N_1879,N_1418);
nand U7110 (N_7110,N_4538,N_507);
or U7111 (N_7111,N_1068,N_2319);
xor U7112 (N_7112,N_4373,N_1841);
xor U7113 (N_7113,N_4822,N_538);
or U7114 (N_7114,N_4909,N_2018);
nand U7115 (N_7115,N_4338,N_3002);
or U7116 (N_7116,N_3861,N_1393);
and U7117 (N_7117,N_4211,N_1438);
nor U7118 (N_7118,N_3247,N_440);
xor U7119 (N_7119,N_1198,N_1741);
xnor U7120 (N_7120,N_4796,N_3481);
or U7121 (N_7121,N_256,N_4662);
and U7122 (N_7122,N_518,N_1490);
or U7123 (N_7123,N_1802,N_3849);
nand U7124 (N_7124,N_55,N_1831);
xor U7125 (N_7125,N_1167,N_4994);
xnor U7126 (N_7126,N_1099,N_3655);
or U7127 (N_7127,N_3641,N_2157);
xor U7128 (N_7128,N_2282,N_4016);
or U7129 (N_7129,N_2477,N_3832);
nand U7130 (N_7130,N_837,N_3293);
or U7131 (N_7131,N_1806,N_3475);
and U7132 (N_7132,N_3147,N_142);
nand U7133 (N_7133,N_880,N_2290);
or U7134 (N_7134,N_725,N_3480);
nand U7135 (N_7135,N_1745,N_3020);
or U7136 (N_7136,N_3190,N_3393);
nand U7137 (N_7137,N_335,N_2333);
and U7138 (N_7138,N_4167,N_1271);
and U7139 (N_7139,N_4149,N_4195);
nor U7140 (N_7140,N_3876,N_182);
xnor U7141 (N_7141,N_2358,N_4894);
and U7142 (N_7142,N_3565,N_2123);
nor U7143 (N_7143,N_1759,N_1001);
or U7144 (N_7144,N_4025,N_3736);
nand U7145 (N_7145,N_1410,N_2499);
and U7146 (N_7146,N_521,N_2800);
xor U7147 (N_7147,N_3325,N_1638);
and U7148 (N_7148,N_1254,N_2467);
xnor U7149 (N_7149,N_914,N_4297);
and U7150 (N_7150,N_3496,N_4515);
or U7151 (N_7151,N_3614,N_1267);
xnor U7152 (N_7152,N_224,N_4783);
xor U7153 (N_7153,N_3922,N_2302);
and U7154 (N_7154,N_4507,N_3903);
or U7155 (N_7155,N_394,N_2854);
nand U7156 (N_7156,N_231,N_32);
nor U7157 (N_7157,N_1219,N_2935);
nand U7158 (N_7158,N_3307,N_2683);
or U7159 (N_7159,N_4159,N_2692);
and U7160 (N_7160,N_4637,N_2771);
xor U7161 (N_7161,N_2158,N_932);
and U7162 (N_7162,N_2391,N_628);
or U7163 (N_7163,N_1492,N_2489);
nor U7164 (N_7164,N_1533,N_1679);
nor U7165 (N_7165,N_4791,N_510);
xor U7166 (N_7166,N_2803,N_2152);
or U7167 (N_7167,N_4019,N_3878);
xor U7168 (N_7168,N_4130,N_2715);
nor U7169 (N_7169,N_4863,N_3010);
or U7170 (N_7170,N_965,N_2841);
xor U7171 (N_7171,N_3902,N_1104);
and U7172 (N_7172,N_4895,N_2986);
nand U7173 (N_7173,N_1795,N_2180);
nor U7174 (N_7174,N_4054,N_4205);
and U7175 (N_7175,N_4030,N_2440);
and U7176 (N_7176,N_871,N_3569);
xor U7177 (N_7177,N_3108,N_3695);
and U7178 (N_7178,N_1930,N_235);
nand U7179 (N_7179,N_2272,N_1398);
xnor U7180 (N_7180,N_4255,N_4469);
and U7181 (N_7181,N_2896,N_3369);
nand U7182 (N_7182,N_3400,N_1178);
nor U7183 (N_7183,N_550,N_3160);
nor U7184 (N_7184,N_1650,N_3493);
xnor U7185 (N_7185,N_592,N_4805);
or U7186 (N_7186,N_2851,N_2772);
nand U7187 (N_7187,N_1822,N_4221);
and U7188 (N_7188,N_4852,N_867);
nor U7189 (N_7189,N_3103,N_1413);
and U7190 (N_7190,N_926,N_4313);
or U7191 (N_7191,N_2505,N_3339);
nand U7192 (N_7192,N_3084,N_691);
or U7193 (N_7193,N_1687,N_210);
nand U7194 (N_7194,N_3470,N_1491);
xor U7195 (N_7195,N_124,N_3364);
nand U7196 (N_7196,N_90,N_3257);
nand U7197 (N_7197,N_2899,N_4482);
and U7198 (N_7198,N_1097,N_3768);
nand U7199 (N_7199,N_1505,N_3751);
xnor U7200 (N_7200,N_4419,N_2238);
and U7201 (N_7201,N_822,N_4273);
nor U7202 (N_7202,N_539,N_3694);
and U7203 (N_7203,N_3533,N_2936);
or U7204 (N_7204,N_4257,N_3121);
xnor U7205 (N_7205,N_1369,N_2354);
and U7206 (N_7206,N_2616,N_2971);
nand U7207 (N_7207,N_1023,N_3822);
and U7208 (N_7208,N_2003,N_4369);
and U7209 (N_7209,N_271,N_531);
and U7210 (N_7210,N_4391,N_796);
and U7211 (N_7211,N_18,N_1552);
or U7212 (N_7212,N_1285,N_3578);
and U7213 (N_7213,N_2283,N_2150);
nor U7214 (N_7214,N_3863,N_1386);
or U7215 (N_7215,N_939,N_3659);
nand U7216 (N_7216,N_1281,N_1294);
or U7217 (N_7217,N_4476,N_3983);
and U7218 (N_7218,N_501,N_3346);
xnor U7219 (N_7219,N_167,N_1107);
nor U7220 (N_7220,N_1549,N_2561);
and U7221 (N_7221,N_527,N_365);
nand U7222 (N_7222,N_3181,N_851);
xor U7223 (N_7223,N_145,N_3624);
or U7224 (N_7224,N_3282,N_2836);
xor U7225 (N_7225,N_2883,N_2236);
nand U7226 (N_7226,N_415,N_1141);
nor U7227 (N_7227,N_3562,N_989);
nor U7228 (N_7228,N_2512,N_3289);
and U7229 (N_7229,N_3798,N_2353);
nor U7230 (N_7230,N_3522,N_2048);
nand U7231 (N_7231,N_2523,N_140);
nand U7232 (N_7232,N_1252,N_8);
or U7233 (N_7233,N_736,N_57);
nand U7234 (N_7234,N_3322,N_1574);
xor U7235 (N_7235,N_3620,N_2445);
and U7236 (N_7236,N_3702,N_2223);
xnor U7237 (N_7237,N_1106,N_3111);
nor U7238 (N_7238,N_3834,N_4012);
nand U7239 (N_7239,N_1249,N_2232);
nor U7240 (N_7240,N_4458,N_4335);
and U7241 (N_7241,N_2578,N_1315);
or U7242 (N_7242,N_4971,N_3673);
or U7243 (N_7243,N_1513,N_1276);
and U7244 (N_7244,N_1704,N_3390);
or U7245 (N_7245,N_36,N_3812);
or U7246 (N_7246,N_1949,N_4394);
nor U7247 (N_7247,N_3531,N_4973);
nand U7248 (N_7248,N_2989,N_2217);
nand U7249 (N_7249,N_4228,N_1565);
nand U7250 (N_7250,N_4220,N_1728);
or U7251 (N_7251,N_4596,N_4440);
or U7252 (N_7252,N_4652,N_707);
and U7253 (N_7253,N_3323,N_3316);
or U7254 (N_7254,N_4871,N_1959);
xnor U7255 (N_7255,N_4251,N_191);
xor U7256 (N_7256,N_174,N_3664);
and U7257 (N_7257,N_2246,N_4445);
and U7258 (N_7258,N_2385,N_465);
and U7259 (N_7259,N_4351,N_4148);
and U7260 (N_7260,N_4188,N_1115);
nor U7261 (N_7261,N_4607,N_2341);
or U7262 (N_7262,N_2153,N_3948);
and U7263 (N_7263,N_151,N_3199);
nand U7264 (N_7264,N_1153,N_4140);
xnor U7265 (N_7265,N_2295,N_3351);
or U7266 (N_7266,N_4803,N_953);
xnor U7267 (N_7267,N_4915,N_2421);
nand U7268 (N_7268,N_4258,N_3685);
nand U7269 (N_7269,N_1695,N_120);
nor U7270 (N_7270,N_4006,N_4929);
nand U7271 (N_7271,N_1440,N_2893);
or U7272 (N_7272,N_4032,N_497);
xnor U7273 (N_7273,N_4122,N_1706);
nor U7274 (N_7274,N_264,N_3164);
or U7275 (N_7275,N_3268,N_4377);
and U7276 (N_7276,N_3065,N_1458);
nor U7277 (N_7277,N_1962,N_2666);
xnor U7278 (N_7278,N_3915,N_4294);
xor U7279 (N_7279,N_3716,N_2222);
or U7280 (N_7280,N_3975,N_4608);
xor U7281 (N_7281,N_4405,N_2434);
nand U7282 (N_7282,N_4904,N_4319);
or U7283 (N_7283,N_1510,N_2357);
nand U7284 (N_7284,N_2226,N_250);
and U7285 (N_7285,N_673,N_4788);
nand U7286 (N_7286,N_4004,N_3886);
or U7287 (N_7287,N_1610,N_1812);
or U7288 (N_7288,N_13,N_1938);
nor U7289 (N_7289,N_4897,N_4464);
or U7290 (N_7290,N_672,N_4572);
and U7291 (N_7291,N_3131,N_4520);
and U7292 (N_7292,N_3284,N_1681);
nand U7293 (N_7293,N_4986,N_300);
and U7294 (N_7294,N_2881,N_3266);
or U7295 (N_7295,N_1031,N_1968);
and U7296 (N_7296,N_4768,N_2900);
nor U7297 (N_7297,N_411,N_248);
and U7298 (N_7298,N_1187,N_852);
and U7299 (N_7299,N_1385,N_1937);
nor U7300 (N_7300,N_779,N_1747);
nor U7301 (N_7301,N_4731,N_3146);
or U7302 (N_7302,N_1047,N_2886);
nand U7303 (N_7303,N_421,N_694);
xnor U7304 (N_7304,N_734,N_1878);
and U7305 (N_7305,N_444,N_2145);
and U7306 (N_7306,N_2738,N_4174);
nand U7307 (N_7307,N_647,N_35);
and U7308 (N_7308,N_270,N_2932);
nand U7309 (N_7309,N_4443,N_2759);
or U7310 (N_7310,N_3225,N_1856);
nor U7311 (N_7311,N_2658,N_2346);
or U7312 (N_7312,N_3092,N_4597);
or U7313 (N_7313,N_3819,N_4949);
or U7314 (N_7314,N_1577,N_633);
xnor U7315 (N_7315,N_128,N_961);
and U7316 (N_7316,N_2373,N_1053);
and U7317 (N_7317,N_3658,N_1873);
nand U7318 (N_7318,N_4447,N_1324);
nand U7319 (N_7319,N_458,N_135);
xnor U7320 (N_7320,N_2114,N_484);
or U7321 (N_7321,N_1662,N_3156);
xor U7322 (N_7322,N_7,N_3295);
xnor U7323 (N_7323,N_4134,N_2415);
xor U7324 (N_7324,N_4548,N_3986);
nor U7325 (N_7325,N_1635,N_2053);
nand U7326 (N_7326,N_53,N_846);
and U7327 (N_7327,N_4068,N_1880);
nor U7328 (N_7328,N_2306,N_866);
or U7329 (N_7329,N_1207,N_1121);
xor U7330 (N_7330,N_3500,N_2948);
and U7331 (N_7331,N_1125,N_17);
nor U7332 (N_7332,N_1800,N_1521);
or U7333 (N_7333,N_743,N_4265);
and U7334 (N_7334,N_3203,N_1479);
or U7335 (N_7335,N_4767,N_1944);
nor U7336 (N_7336,N_1671,N_426);
and U7337 (N_7337,N_4721,N_1619);
and U7338 (N_7338,N_4435,N_4893);
and U7339 (N_7339,N_2650,N_3009);
and U7340 (N_7340,N_353,N_4382);
and U7341 (N_7341,N_1408,N_2026);
and U7342 (N_7342,N_1536,N_2264);
xnor U7343 (N_7343,N_3600,N_4076);
and U7344 (N_7344,N_2648,N_2614);
nand U7345 (N_7345,N_1833,N_4380);
and U7346 (N_7346,N_841,N_4303);
nand U7347 (N_7347,N_574,N_1308);
nor U7348 (N_7348,N_2416,N_4501);
nor U7349 (N_7349,N_995,N_4966);
nand U7350 (N_7350,N_1691,N_3750);
or U7351 (N_7351,N_1098,N_4052);
nor U7352 (N_7352,N_2847,N_3979);
and U7353 (N_7353,N_3158,N_1702);
and U7354 (N_7354,N_3413,N_945);
nor U7355 (N_7355,N_2859,N_4887);
or U7356 (N_7356,N_1263,N_1600);
and U7357 (N_7357,N_4861,N_1033);
xnor U7358 (N_7358,N_4723,N_3756);
nand U7359 (N_7359,N_251,N_4086);
xnor U7360 (N_7360,N_3488,N_3883);
nand U7361 (N_7361,N_340,N_1996);
xor U7362 (N_7362,N_3294,N_126);
or U7363 (N_7363,N_173,N_2913);
and U7364 (N_7364,N_4107,N_216);
or U7365 (N_7365,N_1026,N_2024);
nand U7366 (N_7366,N_3693,N_1296);
nand U7367 (N_7367,N_4700,N_4367);
or U7368 (N_7368,N_4792,N_2644);
xnor U7369 (N_7369,N_4060,N_3959);
and U7370 (N_7370,N_4202,N_2089);
nand U7371 (N_7371,N_849,N_3469);
xor U7372 (N_7372,N_838,N_2594);
nor U7373 (N_7373,N_2296,N_2420);
or U7374 (N_7374,N_3082,N_4123);
nand U7375 (N_7375,N_937,N_2187);
or U7376 (N_7376,N_802,N_1519);
nand U7377 (N_7377,N_1712,N_1010);
nand U7378 (N_7378,N_4604,N_304);
and U7379 (N_7379,N_529,N_4219);
nor U7380 (N_7380,N_667,N_4833);
and U7381 (N_7381,N_4920,N_4716);
nor U7382 (N_7382,N_1529,N_1560);
nor U7383 (N_7383,N_3709,N_3083);
nand U7384 (N_7384,N_3386,N_4525);
or U7385 (N_7385,N_4151,N_3353);
xor U7386 (N_7386,N_241,N_1766);
xnor U7387 (N_7387,N_2014,N_2507);
nor U7388 (N_7388,N_4892,N_2356);
nand U7389 (N_7389,N_4690,N_919);
and U7390 (N_7390,N_230,N_3408);
xor U7391 (N_7391,N_4521,N_1464);
and U7392 (N_7392,N_325,N_2761);
xor U7393 (N_7393,N_660,N_1707);
and U7394 (N_7394,N_522,N_333);
nand U7395 (N_7395,N_805,N_72);
and U7396 (N_7396,N_3165,N_2115);
nor U7397 (N_7397,N_3580,N_3681);
nand U7398 (N_7398,N_634,N_4136);
nand U7399 (N_7399,N_1485,N_936);
or U7400 (N_7400,N_4428,N_466);
or U7401 (N_7401,N_2934,N_2653);
or U7402 (N_7402,N_1703,N_1749);
or U7403 (N_7403,N_2310,N_1998);
and U7404 (N_7404,N_1915,N_3315);
nand U7405 (N_7405,N_468,N_4386);
or U7406 (N_7406,N_2249,N_4610);
nor U7407 (N_7407,N_2626,N_4088);
xor U7408 (N_7408,N_638,N_154);
or U7409 (N_7409,N_3378,N_4246);
nand U7410 (N_7410,N_4583,N_1755);
nor U7411 (N_7411,N_331,N_2081);
nand U7412 (N_7412,N_1442,N_3780);
nand U7413 (N_7413,N_1618,N_2064);
or U7414 (N_7414,N_401,N_3815);
nor U7415 (N_7415,N_4441,N_494);
nor U7416 (N_7416,N_758,N_3141);
nor U7417 (N_7417,N_3930,N_4245);
nor U7418 (N_7418,N_390,N_4522);
and U7419 (N_7419,N_956,N_1499);
and U7420 (N_7420,N_553,N_515);
or U7421 (N_7421,N_255,N_2516);
nor U7422 (N_7422,N_4488,N_4093);
nor U7423 (N_7423,N_4797,N_487);
nor U7424 (N_7424,N_1137,N_606);
xnor U7425 (N_7425,N_3106,N_968);
and U7426 (N_7426,N_3632,N_2439);
nor U7427 (N_7427,N_4055,N_2875);
and U7428 (N_7428,N_3409,N_1875);
nor U7429 (N_7429,N_1899,N_46);
and U7430 (N_7430,N_1716,N_1328);
and U7431 (N_7431,N_4938,N_2005);
xnor U7432 (N_7432,N_2179,N_2590);
nand U7433 (N_7433,N_1517,N_2828);
nand U7434 (N_7434,N_4247,N_3868);
nor U7435 (N_7435,N_3444,N_1416);
or U7436 (N_7436,N_2895,N_4426);
or U7437 (N_7437,N_2655,N_4978);
and U7438 (N_7438,N_3221,N_917);
and U7439 (N_7439,N_3601,N_3763);
or U7440 (N_7440,N_3303,N_2519);
xnor U7441 (N_7441,N_2136,N_2021);
xor U7442 (N_7442,N_3428,N_4598);
xor U7443 (N_7443,N_3097,N_3484);
xor U7444 (N_7444,N_698,N_3864);
and U7445 (N_7445,N_1951,N_1775);
or U7446 (N_7446,N_3091,N_1966);
nand U7447 (N_7447,N_1322,N_3090);
nor U7448 (N_7448,N_3711,N_1916);
nor U7449 (N_7449,N_2918,N_237);
or U7450 (N_7450,N_2317,N_1934);
nand U7451 (N_7451,N_1488,N_3714);
or U7452 (N_7452,N_1253,N_242);
nand U7453 (N_7453,N_648,N_2359);
xnor U7454 (N_7454,N_4023,N_3939);
nor U7455 (N_7455,N_3395,N_4976);
or U7456 (N_7456,N_437,N_3070);
nand U7457 (N_7457,N_356,N_4281);
nor U7458 (N_7458,N_924,N_2661);
and U7459 (N_7459,N_599,N_4190);
xor U7460 (N_7460,N_859,N_4719);
xor U7461 (N_7461,N_2929,N_2316);
and U7462 (N_7462,N_1592,N_3274);
and U7463 (N_7463,N_1876,N_321);
and U7464 (N_7464,N_1330,N_3964);
xor U7465 (N_7465,N_2417,N_1176);
and U7466 (N_7466,N_1906,N_3245);
nand U7467 (N_7467,N_405,N_2425);
and U7468 (N_7468,N_778,N_3743);
xnor U7469 (N_7469,N_2860,N_2336);
or U7470 (N_7470,N_4705,N_761);
or U7471 (N_7471,N_3767,N_1432);
and U7472 (N_7472,N_1947,N_3524);
nor U7473 (N_7473,N_974,N_657);
or U7474 (N_7474,N_3200,N_844);
and U7475 (N_7475,N_4884,N_1952);
xor U7476 (N_7476,N_3552,N_1796);
nand U7477 (N_7477,N_4962,N_921);
and U7478 (N_7478,N_4550,N_630);
xor U7479 (N_7479,N_3843,N_4332);
and U7480 (N_7480,N_43,N_4015);
or U7481 (N_7481,N_22,N_3838);
xnor U7482 (N_7482,N_677,N_3003);
xor U7483 (N_7483,N_2459,N_176);
nand U7484 (N_7484,N_3536,N_4516);
or U7485 (N_7485,N_1861,N_4951);
and U7486 (N_7486,N_1974,N_1503);
and U7487 (N_7487,N_1718,N_1129);
nand U7488 (N_7488,N_2611,N_4761);
or U7489 (N_7489,N_3960,N_1177);
nand U7490 (N_7490,N_267,N_1332);
and U7491 (N_7491,N_4499,N_4128);
and U7492 (N_7492,N_2891,N_1301);
or U7493 (N_7493,N_3269,N_3932);
xnor U7494 (N_7494,N_745,N_4932);
xor U7495 (N_7495,N_3016,N_4846);
nor U7496 (N_7496,N_1874,N_811);
nand U7497 (N_7497,N_3897,N_2262);
xor U7498 (N_7498,N_3674,N_34);
xnor U7499 (N_7499,N_47,N_385);
xor U7500 (N_7500,N_4214,N_672);
xnor U7501 (N_7501,N_4597,N_4890);
and U7502 (N_7502,N_1671,N_2390);
nor U7503 (N_7503,N_3807,N_986);
xor U7504 (N_7504,N_251,N_482);
or U7505 (N_7505,N_342,N_1873);
and U7506 (N_7506,N_3380,N_3553);
xor U7507 (N_7507,N_792,N_260);
or U7508 (N_7508,N_2713,N_500);
and U7509 (N_7509,N_4302,N_668);
nor U7510 (N_7510,N_2811,N_2018);
or U7511 (N_7511,N_2627,N_4799);
nor U7512 (N_7512,N_977,N_1331);
nor U7513 (N_7513,N_3142,N_393);
xnor U7514 (N_7514,N_3070,N_1006);
xnor U7515 (N_7515,N_991,N_4083);
and U7516 (N_7516,N_631,N_1604);
and U7517 (N_7517,N_1332,N_3463);
or U7518 (N_7518,N_1982,N_809);
or U7519 (N_7519,N_3486,N_1342);
and U7520 (N_7520,N_2473,N_4438);
xor U7521 (N_7521,N_1350,N_589);
xnor U7522 (N_7522,N_2659,N_268);
nand U7523 (N_7523,N_2091,N_257);
xnor U7524 (N_7524,N_189,N_3589);
or U7525 (N_7525,N_1644,N_3066);
nor U7526 (N_7526,N_1080,N_247);
or U7527 (N_7527,N_1941,N_4189);
nand U7528 (N_7528,N_1144,N_3755);
or U7529 (N_7529,N_3378,N_597);
and U7530 (N_7530,N_2782,N_2227);
or U7531 (N_7531,N_3605,N_4860);
xor U7532 (N_7532,N_4928,N_2100);
and U7533 (N_7533,N_4358,N_3442);
nand U7534 (N_7534,N_3531,N_3455);
nor U7535 (N_7535,N_1495,N_1449);
xnor U7536 (N_7536,N_1434,N_1070);
and U7537 (N_7537,N_3499,N_488);
nand U7538 (N_7538,N_1573,N_492);
and U7539 (N_7539,N_4460,N_2258);
xnor U7540 (N_7540,N_697,N_4207);
and U7541 (N_7541,N_3389,N_1502);
xnor U7542 (N_7542,N_2451,N_2564);
and U7543 (N_7543,N_295,N_1578);
or U7544 (N_7544,N_2331,N_1910);
nor U7545 (N_7545,N_62,N_3159);
and U7546 (N_7546,N_4684,N_3094);
nand U7547 (N_7547,N_1190,N_2969);
nand U7548 (N_7548,N_4050,N_2301);
or U7549 (N_7549,N_2403,N_84);
xor U7550 (N_7550,N_4519,N_1401);
and U7551 (N_7551,N_1559,N_1358);
nor U7552 (N_7552,N_980,N_1986);
nor U7553 (N_7553,N_3246,N_4286);
or U7554 (N_7554,N_301,N_720);
nor U7555 (N_7555,N_4149,N_2666);
xor U7556 (N_7556,N_2141,N_2225);
nor U7557 (N_7557,N_4384,N_4637);
and U7558 (N_7558,N_2409,N_4106);
xnor U7559 (N_7559,N_456,N_2778);
xnor U7560 (N_7560,N_2120,N_565);
nand U7561 (N_7561,N_3705,N_728);
nor U7562 (N_7562,N_3348,N_3630);
or U7563 (N_7563,N_4656,N_3619);
nand U7564 (N_7564,N_443,N_3105);
or U7565 (N_7565,N_329,N_4397);
xnor U7566 (N_7566,N_482,N_1074);
and U7567 (N_7567,N_4741,N_4726);
nand U7568 (N_7568,N_3920,N_3255);
or U7569 (N_7569,N_3567,N_4656);
or U7570 (N_7570,N_1206,N_2774);
or U7571 (N_7571,N_2431,N_847);
and U7572 (N_7572,N_4006,N_4126);
nand U7573 (N_7573,N_4648,N_47);
and U7574 (N_7574,N_2549,N_1405);
and U7575 (N_7575,N_1905,N_2423);
xnor U7576 (N_7576,N_1662,N_4698);
or U7577 (N_7577,N_4731,N_2626);
or U7578 (N_7578,N_421,N_2148);
nor U7579 (N_7579,N_541,N_4650);
and U7580 (N_7580,N_3537,N_887);
nand U7581 (N_7581,N_3244,N_1419);
xor U7582 (N_7582,N_3492,N_3434);
and U7583 (N_7583,N_101,N_907);
or U7584 (N_7584,N_656,N_3558);
nor U7585 (N_7585,N_1978,N_1407);
nor U7586 (N_7586,N_2537,N_624);
and U7587 (N_7587,N_3490,N_805);
and U7588 (N_7588,N_507,N_1420);
or U7589 (N_7589,N_2001,N_4215);
nand U7590 (N_7590,N_4998,N_2672);
xnor U7591 (N_7591,N_1808,N_396);
and U7592 (N_7592,N_3118,N_1765);
and U7593 (N_7593,N_406,N_4173);
nor U7594 (N_7594,N_2479,N_1306);
or U7595 (N_7595,N_119,N_1722);
nand U7596 (N_7596,N_414,N_1645);
nand U7597 (N_7597,N_3637,N_1820);
xnor U7598 (N_7598,N_2223,N_2644);
and U7599 (N_7599,N_4471,N_474);
nor U7600 (N_7600,N_1120,N_1377);
and U7601 (N_7601,N_2608,N_932);
nand U7602 (N_7602,N_3045,N_1535);
nor U7603 (N_7603,N_2472,N_2763);
xor U7604 (N_7604,N_4517,N_1354);
and U7605 (N_7605,N_2074,N_371);
nor U7606 (N_7606,N_1644,N_1173);
nor U7607 (N_7607,N_3329,N_3204);
and U7608 (N_7608,N_1107,N_4299);
nor U7609 (N_7609,N_4040,N_2222);
nand U7610 (N_7610,N_4970,N_3394);
or U7611 (N_7611,N_1148,N_950);
nor U7612 (N_7612,N_444,N_4233);
nor U7613 (N_7613,N_3320,N_1682);
xnor U7614 (N_7614,N_1854,N_1016);
and U7615 (N_7615,N_699,N_4739);
xor U7616 (N_7616,N_4244,N_3217);
and U7617 (N_7617,N_539,N_2540);
nand U7618 (N_7618,N_4700,N_1807);
and U7619 (N_7619,N_3501,N_4939);
or U7620 (N_7620,N_1507,N_732);
and U7621 (N_7621,N_4680,N_1357);
nand U7622 (N_7622,N_3056,N_1133);
nor U7623 (N_7623,N_1328,N_2492);
nor U7624 (N_7624,N_3615,N_2309);
and U7625 (N_7625,N_1864,N_2747);
and U7626 (N_7626,N_3587,N_2458);
or U7627 (N_7627,N_181,N_4429);
xor U7628 (N_7628,N_1292,N_4210);
nor U7629 (N_7629,N_4440,N_2442);
nor U7630 (N_7630,N_3732,N_3649);
nor U7631 (N_7631,N_2859,N_1299);
or U7632 (N_7632,N_3840,N_3715);
and U7633 (N_7633,N_4434,N_2292);
and U7634 (N_7634,N_4996,N_2107);
nand U7635 (N_7635,N_4368,N_1351);
xor U7636 (N_7636,N_243,N_2318);
nor U7637 (N_7637,N_4056,N_2614);
nand U7638 (N_7638,N_3864,N_771);
xnor U7639 (N_7639,N_895,N_4593);
xnor U7640 (N_7640,N_1338,N_1995);
or U7641 (N_7641,N_1595,N_373);
nand U7642 (N_7642,N_2214,N_3220);
nor U7643 (N_7643,N_62,N_3259);
nand U7644 (N_7644,N_4147,N_4123);
nand U7645 (N_7645,N_1072,N_649);
xnor U7646 (N_7646,N_3919,N_3792);
or U7647 (N_7647,N_3908,N_3289);
and U7648 (N_7648,N_868,N_643);
and U7649 (N_7649,N_3999,N_4085);
nand U7650 (N_7650,N_3618,N_2995);
nand U7651 (N_7651,N_242,N_4258);
xnor U7652 (N_7652,N_595,N_3187);
nand U7653 (N_7653,N_3835,N_3594);
nor U7654 (N_7654,N_535,N_3383);
nor U7655 (N_7655,N_3045,N_926);
and U7656 (N_7656,N_176,N_1628);
and U7657 (N_7657,N_969,N_1448);
nand U7658 (N_7658,N_4331,N_436);
xnor U7659 (N_7659,N_3559,N_698);
xor U7660 (N_7660,N_1204,N_3652);
or U7661 (N_7661,N_921,N_4358);
or U7662 (N_7662,N_2870,N_1517);
nand U7663 (N_7663,N_4638,N_622);
and U7664 (N_7664,N_1230,N_2654);
nand U7665 (N_7665,N_153,N_276);
nor U7666 (N_7666,N_4103,N_3854);
nor U7667 (N_7667,N_1791,N_1652);
or U7668 (N_7668,N_4807,N_3371);
nor U7669 (N_7669,N_1011,N_1739);
and U7670 (N_7670,N_862,N_2062);
or U7671 (N_7671,N_1059,N_29);
xor U7672 (N_7672,N_611,N_3657);
xor U7673 (N_7673,N_110,N_2268);
nand U7674 (N_7674,N_2323,N_1862);
nor U7675 (N_7675,N_1315,N_3552);
or U7676 (N_7676,N_3130,N_2567);
nand U7677 (N_7677,N_1172,N_3499);
nand U7678 (N_7678,N_1046,N_667);
and U7679 (N_7679,N_1122,N_3818);
nand U7680 (N_7680,N_1312,N_1210);
xor U7681 (N_7681,N_671,N_1926);
nand U7682 (N_7682,N_4405,N_994);
nor U7683 (N_7683,N_1416,N_1844);
and U7684 (N_7684,N_2619,N_2059);
nand U7685 (N_7685,N_345,N_3639);
or U7686 (N_7686,N_1583,N_1690);
or U7687 (N_7687,N_3412,N_305);
xnor U7688 (N_7688,N_184,N_3608);
nor U7689 (N_7689,N_745,N_3898);
nor U7690 (N_7690,N_3619,N_3279);
or U7691 (N_7691,N_3215,N_2148);
nor U7692 (N_7692,N_634,N_1981);
nand U7693 (N_7693,N_2221,N_3527);
nor U7694 (N_7694,N_3090,N_2772);
nand U7695 (N_7695,N_996,N_560);
and U7696 (N_7696,N_2368,N_443);
xnor U7697 (N_7697,N_3723,N_734);
and U7698 (N_7698,N_2553,N_2804);
xnor U7699 (N_7699,N_541,N_2093);
nor U7700 (N_7700,N_4499,N_1125);
nor U7701 (N_7701,N_4877,N_4939);
or U7702 (N_7702,N_3129,N_880);
nand U7703 (N_7703,N_2685,N_4436);
nand U7704 (N_7704,N_2830,N_1248);
nor U7705 (N_7705,N_2566,N_4592);
and U7706 (N_7706,N_2987,N_2184);
xor U7707 (N_7707,N_2148,N_2096);
or U7708 (N_7708,N_4369,N_3668);
or U7709 (N_7709,N_34,N_4600);
xor U7710 (N_7710,N_4283,N_875);
xor U7711 (N_7711,N_4995,N_1992);
nor U7712 (N_7712,N_2222,N_658);
xnor U7713 (N_7713,N_1381,N_472);
nand U7714 (N_7714,N_2465,N_3404);
xor U7715 (N_7715,N_880,N_4956);
and U7716 (N_7716,N_1198,N_2289);
xor U7717 (N_7717,N_956,N_4954);
nor U7718 (N_7718,N_2929,N_1533);
xor U7719 (N_7719,N_2932,N_2183);
and U7720 (N_7720,N_3913,N_2926);
nand U7721 (N_7721,N_4243,N_1838);
and U7722 (N_7722,N_4577,N_1072);
xor U7723 (N_7723,N_4546,N_1185);
nand U7724 (N_7724,N_3941,N_3278);
and U7725 (N_7725,N_3059,N_2747);
xor U7726 (N_7726,N_4585,N_2463);
nor U7727 (N_7727,N_2584,N_1791);
or U7728 (N_7728,N_1511,N_3186);
and U7729 (N_7729,N_630,N_3831);
or U7730 (N_7730,N_3423,N_3749);
xnor U7731 (N_7731,N_2871,N_1581);
and U7732 (N_7732,N_4198,N_1712);
or U7733 (N_7733,N_3822,N_3954);
or U7734 (N_7734,N_4411,N_3456);
nor U7735 (N_7735,N_374,N_974);
and U7736 (N_7736,N_1310,N_3635);
nand U7737 (N_7737,N_3852,N_4888);
or U7738 (N_7738,N_124,N_1070);
xor U7739 (N_7739,N_952,N_2198);
nand U7740 (N_7740,N_1179,N_4392);
nor U7741 (N_7741,N_3119,N_3754);
and U7742 (N_7742,N_3540,N_1534);
xor U7743 (N_7743,N_3251,N_2595);
and U7744 (N_7744,N_3615,N_901);
nor U7745 (N_7745,N_3208,N_777);
or U7746 (N_7746,N_2104,N_357);
or U7747 (N_7747,N_1521,N_2880);
and U7748 (N_7748,N_1612,N_3615);
nand U7749 (N_7749,N_3841,N_751);
or U7750 (N_7750,N_3104,N_2222);
and U7751 (N_7751,N_1016,N_1020);
or U7752 (N_7752,N_776,N_2873);
and U7753 (N_7753,N_2107,N_4693);
nand U7754 (N_7754,N_4284,N_3776);
xor U7755 (N_7755,N_1831,N_3773);
nor U7756 (N_7756,N_103,N_1018);
nand U7757 (N_7757,N_4051,N_4319);
nor U7758 (N_7758,N_2862,N_121);
or U7759 (N_7759,N_1499,N_4164);
nor U7760 (N_7760,N_3827,N_1864);
or U7761 (N_7761,N_3471,N_3146);
or U7762 (N_7762,N_1494,N_2031);
or U7763 (N_7763,N_2257,N_3192);
or U7764 (N_7764,N_1659,N_1044);
and U7765 (N_7765,N_1852,N_887);
or U7766 (N_7766,N_451,N_3706);
nand U7767 (N_7767,N_4525,N_1769);
xor U7768 (N_7768,N_378,N_4178);
nor U7769 (N_7769,N_1010,N_18);
xor U7770 (N_7770,N_2736,N_1831);
or U7771 (N_7771,N_2814,N_1274);
nor U7772 (N_7772,N_1499,N_1095);
nand U7773 (N_7773,N_4478,N_3860);
or U7774 (N_7774,N_538,N_2759);
and U7775 (N_7775,N_4363,N_2961);
xor U7776 (N_7776,N_3669,N_1103);
nor U7777 (N_7777,N_1612,N_3089);
or U7778 (N_7778,N_2375,N_4179);
or U7779 (N_7779,N_1026,N_3473);
and U7780 (N_7780,N_506,N_1067);
nor U7781 (N_7781,N_4736,N_2239);
xnor U7782 (N_7782,N_2588,N_103);
xnor U7783 (N_7783,N_588,N_624);
xor U7784 (N_7784,N_3614,N_3399);
and U7785 (N_7785,N_1660,N_4040);
nand U7786 (N_7786,N_2721,N_940);
or U7787 (N_7787,N_2478,N_4771);
xnor U7788 (N_7788,N_2280,N_2920);
nand U7789 (N_7789,N_1287,N_3000);
nand U7790 (N_7790,N_3459,N_1536);
nand U7791 (N_7791,N_2699,N_920);
or U7792 (N_7792,N_1266,N_3993);
nor U7793 (N_7793,N_3772,N_212);
and U7794 (N_7794,N_1361,N_3296);
nand U7795 (N_7795,N_709,N_4048);
nor U7796 (N_7796,N_1043,N_40);
or U7797 (N_7797,N_2221,N_430);
nand U7798 (N_7798,N_4704,N_2191);
or U7799 (N_7799,N_392,N_2509);
and U7800 (N_7800,N_3381,N_1800);
and U7801 (N_7801,N_2193,N_1819);
xnor U7802 (N_7802,N_3590,N_1089);
or U7803 (N_7803,N_1625,N_1882);
or U7804 (N_7804,N_3119,N_278);
and U7805 (N_7805,N_2474,N_3301);
and U7806 (N_7806,N_4696,N_3567);
nor U7807 (N_7807,N_760,N_1600);
nand U7808 (N_7808,N_1274,N_348);
xnor U7809 (N_7809,N_3925,N_222);
and U7810 (N_7810,N_236,N_1848);
nor U7811 (N_7811,N_4035,N_4847);
and U7812 (N_7812,N_2272,N_2976);
nor U7813 (N_7813,N_3615,N_859);
xnor U7814 (N_7814,N_4395,N_1163);
or U7815 (N_7815,N_2942,N_659);
nand U7816 (N_7816,N_3617,N_1773);
nand U7817 (N_7817,N_4709,N_210);
and U7818 (N_7818,N_4517,N_3212);
nor U7819 (N_7819,N_1911,N_3930);
or U7820 (N_7820,N_378,N_4386);
nor U7821 (N_7821,N_4612,N_2292);
nand U7822 (N_7822,N_4024,N_4394);
nor U7823 (N_7823,N_3038,N_4627);
nor U7824 (N_7824,N_577,N_3381);
nand U7825 (N_7825,N_4768,N_4975);
nand U7826 (N_7826,N_34,N_2160);
or U7827 (N_7827,N_3578,N_802);
and U7828 (N_7828,N_4688,N_4426);
and U7829 (N_7829,N_3493,N_1860);
xor U7830 (N_7830,N_1141,N_2207);
xnor U7831 (N_7831,N_4166,N_1093);
nand U7832 (N_7832,N_3976,N_1048);
and U7833 (N_7833,N_948,N_4317);
or U7834 (N_7834,N_1256,N_3053);
nand U7835 (N_7835,N_3886,N_3077);
nor U7836 (N_7836,N_50,N_1964);
or U7837 (N_7837,N_4823,N_772);
or U7838 (N_7838,N_4414,N_774);
nand U7839 (N_7839,N_4585,N_1087);
nor U7840 (N_7840,N_148,N_3753);
or U7841 (N_7841,N_957,N_4593);
nor U7842 (N_7842,N_2611,N_4851);
nor U7843 (N_7843,N_2658,N_1239);
nand U7844 (N_7844,N_4045,N_4588);
and U7845 (N_7845,N_2753,N_903);
and U7846 (N_7846,N_2139,N_3989);
xnor U7847 (N_7847,N_1675,N_1553);
nor U7848 (N_7848,N_3429,N_1167);
xnor U7849 (N_7849,N_3661,N_2058);
nor U7850 (N_7850,N_2175,N_530);
nor U7851 (N_7851,N_2859,N_227);
nand U7852 (N_7852,N_788,N_3878);
nor U7853 (N_7853,N_2848,N_2441);
nor U7854 (N_7854,N_2886,N_2789);
nand U7855 (N_7855,N_4572,N_1606);
or U7856 (N_7856,N_4424,N_3945);
and U7857 (N_7857,N_1666,N_850);
xnor U7858 (N_7858,N_1753,N_3682);
nor U7859 (N_7859,N_2725,N_3404);
nand U7860 (N_7860,N_3475,N_3270);
or U7861 (N_7861,N_1385,N_2109);
nand U7862 (N_7862,N_4092,N_2184);
nand U7863 (N_7863,N_1004,N_2358);
xor U7864 (N_7864,N_4850,N_3655);
and U7865 (N_7865,N_1688,N_643);
xor U7866 (N_7866,N_1659,N_395);
and U7867 (N_7867,N_4295,N_3580);
nand U7868 (N_7868,N_3474,N_924);
nand U7869 (N_7869,N_1384,N_4334);
nor U7870 (N_7870,N_1125,N_1561);
or U7871 (N_7871,N_3674,N_4805);
and U7872 (N_7872,N_4927,N_3307);
xnor U7873 (N_7873,N_362,N_1939);
nor U7874 (N_7874,N_4698,N_2231);
or U7875 (N_7875,N_199,N_821);
xnor U7876 (N_7876,N_4849,N_3814);
or U7877 (N_7877,N_1744,N_634);
nor U7878 (N_7878,N_1912,N_1778);
nand U7879 (N_7879,N_865,N_1375);
or U7880 (N_7880,N_3988,N_2945);
nand U7881 (N_7881,N_3056,N_3333);
or U7882 (N_7882,N_3846,N_624);
xnor U7883 (N_7883,N_3606,N_98);
nor U7884 (N_7884,N_505,N_480);
nor U7885 (N_7885,N_3427,N_2849);
or U7886 (N_7886,N_4511,N_235);
xor U7887 (N_7887,N_4842,N_3752);
nand U7888 (N_7888,N_3934,N_3479);
and U7889 (N_7889,N_4812,N_2341);
or U7890 (N_7890,N_2374,N_801);
and U7891 (N_7891,N_3835,N_3307);
or U7892 (N_7892,N_3040,N_2432);
or U7893 (N_7893,N_1194,N_4514);
and U7894 (N_7894,N_1974,N_206);
nor U7895 (N_7895,N_3062,N_4752);
nor U7896 (N_7896,N_4953,N_3899);
and U7897 (N_7897,N_4228,N_474);
nand U7898 (N_7898,N_4612,N_595);
or U7899 (N_7899,N_3102,N_3307);
nand U7900 (N_7900,N_2382,N_3722);
and U7901 (N_7901,N_2985,N_2452);
or U7902 (N_7902,N_912,N_2875);
nor U7903 (N_7903,N_2429,N_1501);
or U7904 (N_7904,N_4629,N_3899);
or U7905 (N_7905,N_2303,N_2704);
and U7906 (N_7906,N_4686,N_638);
xnor U7907 (N_7907,N_4271,N_4641);
nand U7908 (N_7908,N_3183,N_4554);
or U7909 (N_7909,N_2599,N_3863);
or U7910 (N_7910,N_4429,N_1294);
xor U7911 (N_7911,N_2332,N_4806);
and U7912 (N_7912,N_2459,N_1698);
nor U7913 (N_7913,N_1193,N_351);
xor U7914 (N_7914,N_3002,N_1053);
nand U7915 (N_7915,N_1789,N_2289);
xor U7916 (N_7916,N_438,N_4052);
and U7917 (N_7917,N_4912,N_1813);
nor U7918 (N_7918,N_146,N_1831);
nand U7919 (N_7919,N_735,N_1582);
xnor U7920 (N_7920,N_2544,N_3109);
xnor U7921 (N_7921,N_4176,N_3357);
or U7922 (N_7922,N_2977,N_3776);
nor U7923 (N_7923,N_1073,N_442);
or U7924 (N_7924,N_305,N_1868);
nor U7925 (N_7925,N_3553,N_1797);
and U7926 (N_7926,N_531,N_301);
xnor U7927 (N_7927,N_2180,N_819);
nand U7928 (N_7928,N_4198,N_4220);
and U7929 (N_7929,N_4961,N_1143);
xnor U7930 (N_7930,N_255,N_946);
and U7931 (N_7931,N_54,N_2837);
nand U7932 (N_7932,N_4899,N_3036);
or U7933 (N_7933,N_3653,N_792);
nor U7934 (N_7934,N_2743,N_675);
nand U7935 (N_7935,N_4976,N_642);
and U7936 (N_7936,N_3314,N_3703);
xor U7937 (N_7937,N_1427,N_3352);
or U7938 (N_7938,N_4481,N_27);
or U7939 (N_7939,N_3408,N_3927);
xnor U7940 (N_7940,N_669,N_3249);
or U7941 (N_7941,N_2230,N_4105);
and U7942 (N_7942,N_1686,N_3875);
nand U7943 (N_7943,N_985,N_2268);
nor U7944 (N_7944,N_4243,N_4017);
or U7945 (N_7945,N_145,N_3015);
xor U7946 (N_7946,N_1605,N_1208);
nand U7947 (N_7947,N_2539,N_1352);
nand U7948 (N_7948,N_522,N_1450);
or U7949 (N_7949,N_4674,N_1753);
xor U7950 (N_7950,N_447,N_39);
nand U7951 (N_7951,N_2650,N_3218);
nand U7952 (N_7952,N_324,N_3748);
xnor U7953 (N_7953,N_2339,N_809);
and U7954 (N_7954,N_3678,N_2484);
xnor U7955 (N_7955,N_3961,N_1126);
nand U7956 (N_7956,N_852,N_1830);
xnor U7957 (N_7957,N_2137,N_3768);
and U7958 (N_7958,N_743,N_783);
nor U7959 (N_7959,N_4188,N_61);
nand U7960 (N_7960,N_206,N_3240);
nand U7961 (N_7961,N_4389,N_3448);
and U7962 (N_7962,N_4226,N_379);
or U7963 (N_7963,N_1666,N_2887);
and U7964 (N_7964,N_297,N_1878);
xor U7965 (N_7965,N_2077,N_572);
nor U7966 (N_7966,N_59,N_3650);
and U7967 (N_7967,N_1753,N_2364);
nor U7968 (N_7968,N_4113,N_3237);
nand U7969 (N_7969,N_58,N_2562);
xor U7970 (N_7970,N_1424,N_4950);
nor U7971 (N_7971,N_3686,N_4421);
xor U7972 (N_7972,N_3431,N_3004);
or U7973 (N_7973,N_4613,N_939);
xnor U7974 (N_7974,N_1921,N_1520);
and U7975 (N_7975,N_4327,N_4275);
or U7976 (N_7976,N_4918,N_1732);
and U7977 (N_7977,N_4920,N_2350);
nand U7978 (N_7978,N_2739,N_564);
and U7979 (N_7979,N_4553,N_79);
nor U7980 (N_7980,N_3208,N_3654);
nor U7981 (N_7981,N_33,N_3602);
and U7982 (N_7982,N_1522,N_365);
nor U7983 (N_7983,N_303,N_2716);
nor U7984 (N_7984,N_128,N_903);
nor U7985 (N_7985,N_2454,N_158);
nor U7986 (N_7986,N_2624,N_659);
nor U7987 (N_7987,N_298,N_1316);
nand U7988 (N_7988,N_4221,N_1446);
nand U7989 (N_7989,N_308,N_2314);
xnor U7990 (N_7990,N_419,N_4219);
and U7991 (N_7991,N_4590,N_3983);
and U7992 (N_7992,N_3574,N_4162);
xnor U7993 (N_7993,N_1964,N_4816);
nand U7994 (N_7994,N_4523,N_826);
nor U7995 (N_7995,N_1118,N_2366);
xor U7996 (N_7996,N_2083,N_2376);
nand U7997 (N_7997,N_4326,N_3394);
nand U7998 (N_7998,N_451,N_1971);
nor U7999 (N_7999,N_1728,N_3194);
nand U8000 (N_8000,N_2045,N_3818);
nand U8001 (N_8001,N_676,N_886);
and U8002 (N_8002,N_1348,N_2385);
nor U8003 (N_8003,N_2074,N_2779);
nand U8004 (N_8004,N_1716,N_3698);
nor U8005 (N_8005,N_3951,N_25);
and U8006 (N_8006,N_4344,N_317);
or U8007 (N_8007,N_2728,N_2740);
or U8008 (N_8008,N_1328,N_991);
and U8009 (N_8009,N_1357,N_161);
or U8010 (N_8010,N_1752,N_3580);
nor U8011 (N_8011,N_2365,N_3201);
nor U8012 (N_8012,N_902,N_2340);
xor U8013 (N_8013,N_3839,N_697);
xor U8014 (N_8014,N_2117,N_1702);
xor U8015 (N_8015,N_3471,N_2479);
or U8016 (N_8016,N_3252,N_7);
xor U8017 (N_8017,N_3785,N_4719);
xor U8018 (N_8018,N_4053,N_1105);
or U8019 (N_8019,N_4578,N_704);
or U8020 (N_8020,N_3649,N_3340);
nor U8021 (N_8021,N_4083,N_68);
xor U8022 (N_8022,N_2624,N_3724);
xor U8023 (N_8023,N_3345,N_882);
nand U8024 (N_8024,N_2248,N_1970);
xnor U8025 (N_8025,N_2306,N_829);
or U8026 (N_8026,N_2797,N_4496);
xnor U8027 (N_8027,N_1557,N_3874);
and U8028 (N_8028,N_4389,N_2862);
or U8029 (N_8029,N_1631,N_2076);
nor U8030 (N_8030,N_2166,N_4696);
nor U8031 (N_8031,N_4127,N_4419);
xnor U8032 (N_8032,N_3129,N_4483);
and U8033 (N_8033,N_3189,N_1397);
nor U8034 (N_8034,N_1986,N_3700);
and U8035 (N_8035,N_1982,N_2182);
nor U8036 (N_8036,N_4061,N_3525);
nor U8037 (N_8037,N_4122,N_3918);
nand U8038 (N_8038,N_3717,N_2478);
nor U8039 (N_8039,N_1029,N_4288);
and U8040 (N_8040,N_3608,N_3814);
xnor U8041 (N_8041,N_2959,N_2052);
xor U8042 (N_8042,N_4016,N_2763);
or U8043 (N_8043,N_4617,N_3080);
xor U8044 (N_8044,N_4749,N_2796);
xor U8045 (N_8045,N_1089,N_4887);
and U8046 (N_8046,N_500,N_912);
or U8047 (N_8047,N_3326,N_1530);
xor U8048 (N_8048,N_814,N_1035);
nand U8049 (N_8049,N_1400,N_1117);
nand U8050 (N_8050,N_2793,N_2121);
or U8051 (N_8051,N_2292,N_981);
nand U8052 (N_8052,N_2216,N_4334);
and U8053 (N_8053,N_2895,N_856);
nand U8054 (N_8054,N_4320,N_3620);
or U8055 (N_8055,N_3054,N_4099);
nand U8056 (N_8056,N_4537,N_29);
and U8057 (N_8057,N_159,N_3668);
or U8058 (N_8058,N_2026,N_2059);
or U8059 (N_8059,N_2698,N_4211);
xnor U8060 (N_8060,N_3540,N_395);
nand U8061 (N_8061,N_3252,N_321);
xnor U8062 (N_8062,N_4392,N_2314);
and U8063 (N_8063,N_1650,N_2841);
nor U8064 (N_8064,N_3869,N_3523);
nand U8065 (N_8065,N_3212,N_3921);
and U8066 (N_8066,N_2211,N_4261);
nand U8067 (N_8067,N_4642,N_4338);
nand U8068 (N_8068,N_3411,N_2426);
nand U8069 (N_8069,N_1429,N_2670);
and U8070 (N_8070,N_570,N_1838);
or U8071 (N_8071,N_1240,N_126);
nor U8072 (N_8072,N_2927,N_4094);
nand U8073 (N_8073,N_4528,N_2059);
nor U8074 (N_8074,N_2555,N_2992);
or U8075 (N_8075,N_2142,N_3534);
and U8076 (N_8076,N_490,N_1807);
nor U8077 (N_8077,N_1149,N_3410);
or U8078 (N_8078,N_3076,N_2456);
nand U8079 (N_8079,N_3089,N_834);
and U8080 (N_8080,N_273,N_2559);
and U8081 (N_8081,N_4298,N_4601);
or U8082 (N_8082,N_918,N_3896);
nor U8083 (N_8083,N_785,N_3419);
nand U8084 (N_8084,N_1622,N_3866);
or U8085 (N_8085,N_3910,N_1573);
xnor U8086 (N_8086,N_3177,N_4688);
nand U8087 (N_8087,N_463,N_1368);
and U8088 (N_8088,N_496,N_3434);
nor U8089 (N_8089,N_2201,N_4592);
and U8090 (N_8090,N_1605,N_1671);
nand U8091 (N_8091,N_2063,N_1500);
nor U8092 (N_8092,N_1752,N_4751);
nand U8093 (N_8093,N_30,N_3969);
nand U8094 (N_8094,N_4682,N_2790);
or U8095 (N_8095,N_372,N_2317);
or U8096 (N_8096,N_2554,N_396);
and U8097 (N_8097,N_2930,N_2869);
nand U8098 (N_8098,N_3080,N_3188);
nand U8099 (N_8099,N_1828,N_82);
nand U8100 (N_8100,N_1125,N_488);
or U8101 (N_8101,N_1496,N_1679);
nand U8102 (N_8102,N_1713,N_5);
nand U8103 (N_8103,N_268,N_2179);
nor U8104 (N_8104,N_963,N_2361);
and U8105 (N_8105,N_1985,N_1756);
nor U8106 (N_8106,N_3397,N_764);
nand U8107 (N_8107,N_4590,N_2377);
nand U8108 (N_8108,N_4856,N_3945);
nand U8109 (N_8109,N_2023,N_3826);
nor U8110 (N_8110,N_3177,N_4811);
and U8111 (N_8111,N_1531,N_3544);
and U8112 (N_8112,N_2388,N_1002);
or U8113 (N_8113,N_3884,N_465);
nor U8114 (N_8114,N_501,N_592);
nand U8115 (N_8115,N_954,N_2127);
nor U8116 (N_8116,N_3275,N_4671);
nand U8117 (N_8117,N_4216,N_3859);
or U8118 (N_8118,N_4142,N_238);
nor U8119 (N_8119,N_3738,N_3150);
or U8120 (N_8120,N_2355,N_3722);
or U8121 (N_8121,N_295,N_3319);
nand U8122 (N_8122,N_2563,N_3220);
nor U8123 (N_8123,N_875,N_3340);
or U8124 (N_8124,N_2118,N_1937);
nor U8125 (N_8125,N_3042,N_453);
nor U8126 (N_8126,N_4101,N_2223);
or U8127 (N_8127,N_602,N_4225);
nand U8128 (N_8128,N_1953,N_996);
nor U8129 (N_8129,N_2017,N_1405);
nand U8130 (N_8130,N_1839,N_3160);
xor U8131 (N_8131,N_809,N_3938);
nand U8132 (N_8132,N_162,N_1517);
and U8133 (N_8133,N_3349,N_1872);
nand U8134 (N_8134,N_10,N_4335);
xnor U8135 (N_8135,N_3981,N_3375);
nand U8136 (N_8136,N_2604,N_543);
or U8137 (N_8137,N_2854,N_1889);
or U8138 (N_8138,N_4009,N_3826);
and U8139 (N_8139,N_4208,N_1252);
nor U8140 (N_8140,N_3964,N_3610);
nor U8141 (N_8141,N_1999,N_3979);
and U8142 (N_8142,N_1688,N_925);
and U8143 (N_8143,N_2185,N_662);
or U8144 (N_8144,N_1699,N_3904);
nor U8145 (N_8145,N_4780,N_1293);
nand U8146 (N_8146,N_1737,N_4916);
or U8147 (N_8147,N_1664,N_14);
nand U8148 (N_8148,N_4713,N_3410);
nor U8149 (N_8149,N_3098,N_1850);
and U8150 (N_8150,N_4522,N_3740);
and U8151 (N_8151,N_4159,N_83);
nor U8152 (N_8152,N_4965,N_117);
or U8153 (N_8153,N_2451,N_677);
and U8154 (N_8154,N_4544,N_4780);
nand U8155 (N_8155,N_1182,N_1710);
or U8156 (N_8156,N_2505,N_3652);
and U8157 (N_8157,N_1787,N_1164);
and U8158 (N_8158,N_3675,N_1368);
and U8159 (N_8159,N_2495,N_4293);
or U8160 (N_8160,N_2141,N_2291);
or U8161 (N_8161,N_419,N_4891);
xor U8162 (N_8162,N_1135,N_1209);
or U8163 (N_8163,N_555,N_2241);
xor U8164 (N_8164,N_1109,N_1589);
and U8165 (N_8165,N_554,N_2867);
nor U8166 (N_8166,N_1375,N_1223);
nor U8167 (N_8167,N_4321,N_3047);
nor U8168 (N_8168,N_142,N_1637);
nand U8169 (N_8169,N_3992,N_2178);
nand U8170 (N_8170,N_4801,N_3768);
nand U8171 (N_8171,N_4620,N_2587);
xnor U8172 (N_8172,N_1871,N_1361);
xor U8173 (N_8173,N_407,N_4196);
nor U8174 (N_8174,N_4493,N_3561);
xnor U8175 (N_8175,N_2324,N_3350);
and U8176 (N_8176,N_2337,N_2138);
xnor U8177 (N_8177,N_3252,N_914);
or U8178 (N_8178,N_4540,N_3033);
and U8179 (N_8179,N_154,N_2537);
nand U8180 (N_8180,N_2710,N_1341);
nand U8181 (N_8181,N_2332,N_2438);
nor U8182 (N_8182,N_2084,N_1654);
nor U8183 (N_8183,N_1220,N_1275);
xor U8184 (N_8184,N_4570,N_395);
nand U8185 (N_8185,N_1249,N_4138);
or U8186 (N_8186,N_3813,N_668);
nor U8187 (N_8187,N_4179,N_2278);
xnor U8188 (N_8188,N_3209,N_3252);
or U8189 (N_8189,N_1732,N_1506);
nor U8190 (N_8190,N_4351,N_4929);
nor U8191 (N_8191,N_3519,N_1553);
and U8192 (N_8192,N_4951,N_3814);
xor U8193 (N_8193,N_1460,N_4103);
nor U8194 (N_8194,N_4766,N_242);
nand U8195 (N_8195,N_282,N_1433);
nand U8196 (N_8196,N_2425,N_1487);
and U8197 (N_8197,N_45,N_2463);
or U8198 (N_8198,N_2027,N_3881);
and U8199 (N_8199,N_3812,N_984);
nor U8200 (N_8200,N_3205,N_3770);
and U8201 (N_8201,N_2906,N_1549);
xnor U8202 (N_8202,N_1858,N_3704);
xor U8203 (N_8203,N_2736,N_3662);
xnor U8204 (N_8204,N_2931,N_822);
or U8205 (N_8205,N_1422,N_3072);
nor U8206 (N_8206,N_1817,N_2037);
or U8207 (N_8207,N_680,N_1008);
xnor U8208 (N_8208,N_135,N_2137);
or U8209 (N_8209,N_2505,N_2051);
nand U8210 (N_8210,N_1763,N_1663);
and U8211 (N_8211,N_4996,N_4701);
xor U8212 (N_8212,N_3953,N_1428);
and U8213 (N_8213,N_74,N_1833);
xnor U8214 (N_8214,N_827,N_845);
and U8215 (N_8215,N_4466,N_2268);
nor U8216 (N_8216,N_962,N_4635);
and U8217 (N_8217,N_3558,N_2568);
nand U8218 (N_8218,N_1158,N_3739);
xor U8219 (N_8219,N_159,N_2333);
or U8220 (N_8220,N_3532,N_4358);
or U8221 (N_8221,N_1154,N_4082);
xor U8222 (N_8222,N_1743,N_1818);
and U8223 (N_8223,N_3331,N_4934);
xnor U8224 (N_8224,N_1213,N_4965);
or U8225 (N_8225,N_3478,N_2848);
nor U8226 (N_8226,N_854,N_4190);
and U8227 (N_8227,N_1239,N_680);
and U8228 (N_8228,N_3956,N_2953);
and U8229 (N_8229,N_1903,N_2607);
nand U8230 (N_8230,N_2570,N_44);
nand U8231 (N_8231,N_3825,N_2735);
xnor U8232 (N_8232,N_774,N_2468);
xnor U8233 (N_8233,N_3732,N_3203);
or U8234 (N_8234,N_3058,N_4118);
xnor U8235 (N_8235,N_4054,N_3607);
and U8236 (N_8236,N_2772,N_4818);
nor U8237 (N_8237,N_1499,N_1176);
nand U8238 (N_8238,N_3025,N_735);
xnor U8239 (N_8239,N_1242,N_376);
nor U8240 (N_8240,N_1071,N_3141);
nand U8241 (N_8241,N_584,N_172);
or U8242 (N_8242,N_3898,N_4623);
xor U8243 (N_8243,N_2543,N_4740);
and U8244 (N_8244,N_1895,N_3598);
or U8245 (N_8245,N_1265,N_2828);
and U8246 (N_8246,N_4177,N_3971);
and U8247 (N_8247,N_4227,N_2941);
and U8248 (N_8248,N_2529,N_485);
xor U8249 (N_8249,N_1176,N_1077);
xnor U8250 (N_8250,N_2014,N_486);
and U8251 (N_8251,N_4836,N_2515);
xor U8252 (N_8252,N_1364,N_3250);
xnor U8253 (N_8253,N_1438,N_1014);
nor U8254 (N_8254,N_3752,N_4877);
xnor U8255 (N_8255,N_3012,N_3136);
nand U8256 (N_8256,N_4717,N_4636);
nor U8257 (N_8257,N_1977,N_1292);
and U8258 (N_8258,N_4,N_2709);
nand U8259 (N_8259,N_1878,N_3472);
nand U8260 (N_8260,N_1520,N_315);
or U8261 (N_8261,N_4147,N_2739);
nor U8262 (N_8262,N_717,N_2906);
or U8263 (N_8263,N_2830,N_3838);
and U8264 (N_8264,N_3980,N_982);
nand U8265 (N_8265,N_1686,N_395);
or U8266 (N_8266,N_3301,N_82);
or U8267 (N_8267,N_1053,N_3174);
and U8268 (N_8268,N_1540,N_4950);
xnor U8269 (N_8269,N_331,N_4615);
nor U8270 (N_8270,N_1582,N_4987);
nand U8271 (N_8271,N_2886,N_4810);
or U8272 (N_8272,N_1313,N_337);
nor U8273 (N_8273,N_4703,N_4924);
xor U8274 (N_8274,N_1159,N_1625);
xnor U8275 (N_8275,N_3594,N_336);
and U8276 (N_8276,N_3099,N_4398);
and U8277 (N_8277,N_1367,N_629);
nand U8278 (N_8278,N_4039,N_2497);
xnor U8279 (N_8279,N_619,N_3156);
nand U8280 (N_8280,N_3218,N_490);
and U8281 (N_8281,N_1015,N_699);
nor U8282 (N_8282,N_3889,N_3240);
and U8283 (N_8283,N_3760,N_1574);
and U8284 (N_8284,N_1443,N_2792);
nand U8285 (N_8285,N_4686,N_3915);
or U8286 (N_8286,N_4193,N_4192);
nand U8287 (N_8287,N_3065,N_883);
or U8288 (N_8288,N_491,N_2603);
and U8289 (N_8289,N_1374,N_2859);
nor U8290 (N_8290,N_3029,N_4445);
or U8291 (N_8291,N_2035,N_2969);
xor U8292 (N_8292,N_621,N_2360);
and U8293 (N_8293,N_1633,N_82);
nand U8294 (N_8294,N_3320,N_4783);
nand U8295 (N_8295,N_765,N_2949);
xor U8296 (N_8296,N_370,N_4134);
nand U8297 (N_8297,N_3151,N_1376);
nand U8298 (N_8298,N_1289,N_3663);
nand U8299 (N_8299,N_1066,N_4096);
and U8300 (N_8300,N_753,N_3365);
xnor U8301 (N_8301,N_2661,N_612);
and U8302 (N_8302,N_2910,N_1761);
or U8303 (N_8303,N_3469,N_3467);
xnor U8304 (N_8304,N_4028,N_2082);
xor U8305 (N_8305,N_2906,N_4841);
and U8306 (N_8306,N_4133,N_4693);
nand U8307 (N_8307,N_4117,N_1918);
xnor U8308 (N_8308,N_2601,N_3947);
nand U8309 (N_8309,N_1367,N_4626);
nor U8310 (N_8310,N_4274,N_1482);
and U8311 (N_8311,N_3525,N_4877);
xnor U8312 (N_8312,N_344,N_4191);
xor U8313 (N_8313,N_2058,N_3531);
nand U8314 (N_8314,N_1975,N_4201);
nand U8315 (N_8315,N_2834,N_2880);
and U8316 (N_8316,N_3843,N_3610);
or U8317 (N_8317,N_90,N_1790);
nand U8318 (N_8318,N_2280,N_2566);
and U8319 (N_8319,N_4727,N_1255);
nand U8320 (N_8320,N_3615,N_2904);
nand U8321 (N_8321,N_2647,N_3953);
or U8322 (N_8322,N_4748,N_1369);
xor U8323 (N_8323,N_2123,N_580);
xor U8324 (N_8324,N_358,N_4591);
nand U8325 (N_8325,N_4700,N_2556);
and U8326 (N_8326,N_2892,N_1865);
or U8327 (N_8327,N_2499,N_415);
or U8328 (N_8328,N_2405,N_1318);
or U8329 (N_8329,N_4016,N_2879);
or U8330 (N_8330,N_95,N_716);
or U8331 (N_8331,N_745,N_3273);
nor U8332 (N_8332,N_588,N_1474);
or U8333 (N_8333,N_1146,N_1162);
or U8334 (N_8334,N_2147,N_411);
nand U8335 (N_8335,N_3923,N_100);
xor U8336 (N_8336,N_931,N_4572);
or U8337 (N_8337,N_4179,N_2540);
nor U8338 (N_8338,N_4384,N_1024);
nand U8339 (N_8339,N_3460,N_876);
xor U8340 (N_8340,N_3385,N_3523);
nor U8341 (N_8341,N_4312,N_872);
or U8342 (N_8342,N_551,N_491);
nor U8343 (N_8343,N_1384,N_2022);
nand U8344 (N_8344,N_4758,N_1363);
xnor U8345 (N_8345,N_4649,N_1247);
or U8346 (N_8346,N_2454,N_4971);
or U8347 (N_8347,N_3352,N_167);
or U8348 (N_8348,N_4044,N_1183);
xor U8349 (N_8349,N_3998,N_3456);
nand U8350 (N_8350,N_4278,N_2087);
xor U8351 (N_8351,N_1444,N_3612);
nor U8352 (N_8352,N_669,N_2942);
and U8353 (N_8353,N_1335,N_3556);
xor U8354 (N_8354,N_223,N_2474);
xor U8355 (N_8355,N_1198,N_3169);
xor U8356 (N_8356,N_2192,N_1437);
xnor U8357 (N_8357,N_3099,N_1176);
or U8358 (N_8358,N_3819,N_2739);
and U8359 (N_8359,N_65,N_2104);
nand U8360 (N_8360,N_4086,N_3017);
or U8361 (N_8361,N_4535,N_3498);
nor U8362 (N_8362,N_2524,N_3298);
nand U8363 (N_8363,N_1782,N_3449);
and U8364 (N_8364,N_1271,N_2979);
nand U8365 (N_8365,N_3861,N_145);
xnor U8366 (N_8366,N_1443,N_4108);
nand U8367 (N_8367,N_2215,N_1625);
and U8368 (N_8368,N_3164,N_2304);
or U8369 (N_8369,N_1847,N_3847);
nor U8370 (N_8370,N_4943,N_71);
nor U8371 (N_8371,N_2815,N_1895);
nand U8372 (N_8372,N_4323,N_745);
nor U8373 (N_8373,N_1833,N_2155);
xor U8374 (N_8374,N_3091,N_2852);
or U8375 (N_8375,N_4393,N_3778);
nand U8376 (N_8376,N_3584,N_4621);
nor U8377 (N_8377,N_2578,N_877);
nand U8378 (N_8378,N_1960,N_2651);
and U8379 (N_8379,N_4790,N_1232);
and U8380 (N_8380,N_3344,N_1363);
or U8381 (N_8381,N_2893,N_4225);
or U8382 (N_8382,N_2916,N_285);
nor U8383 (N_8383,N_4937,N_1122);
xor U8384 (N_8384,N_956,N_872);
nor U8385 (N_8385,N_1048,N_138);
and U8386 (N_8386,N_4225,N_4320);
and U8387 (N_8387,N_2794,N_4577);
and U8388 (N_8388,N_1480,N_3376);
and U8389 (N_8389,N_789,N_4330);
nand U8390 (N_8390,N_3802,N_1368);
xnor U8391 (N_8391,N_3949,N_1120);
nand U8392 (N_8392,N_2579,N_3514);
and U8393 (N_8393,N_737,N_444);
and U8394 (N_8394,N_1142,N_2254);
xor U8395 (N_8395,N_2289,N_692);
xnor U8396 (N_8396,N_3707,N_3947);
nand U8397 (N_8397,N_386,N_2089);
nor U8398 (N_8398,N_3720,N_3782);
nor U8399 (N_8399,N_3853,N_980);
nor U8400 (N_8400,N_3844,N_3259);
nor U8401 (N_8401,N_1265,N_2050);
or U8402 (N_8402,N_909,N_3361);
xor U8403 (N_8403,N_1867,N_2132);
and U8404 (N_8404,N_1619,N_4294);
and U8405 (N_8405,N_3539,N_1245);
nor U8406 (N_8406,N_4062,N_1837);
nand U8407 (N_8407,N_1680,N_2283);
and U8408 (N_8408,N_2507,N_1874);
nand U8409 (N_8409,N_120,N_4506);
and U8410 (N_8410,N_3600,N_2640);
and U8411 (N_8411,N_548,N_904);
and U8412 (N_8412,N_938,N_427);
xnor U8413 (N_8413,N_1756,N_4998);
xnor U8414 (N_8414,N_4833,N_3856);
and U8415 (N_8415,N_2470,N_1589);
or U8416 (N_8416,N_2646,N_1342);
xnor U8417 (N_8417,N_3673,N_954);
or U8418 (N_8418,N_2121,N_1339);
and U8419 (N_8419,N_479,N_836);
nand U8420 (N_8420,N_147,N_2216);
nand U8421 (N_8421,N_616,N_2763);
nand U8422 (N_8422,N_3873,N_590);
nor U8423 (N_8423,N_4227,N_2696);
nand U8424 (N_8424,N_2520,N_3716);
nand U8425 (N_8425,N_1442,N_3602);
nand U8426 (N_8426,N_1318,N_2862);
xnor U8427 (N_8427,N_4327,N_2458);
and U8428 (N_8428,N_2667,N_2944);
and U8429 (N_8429,N_1352,N_607);
nor U8430 (N_8430,N_2507,N_4984);
and U8431 (N_8431,N_4397,N_4538);
xnor U8432 (N_8432,N_2296,N_4881);
or U8433 (N_8433,N_4472,N_63);
nand U8434 (N_8434,N_2222,N_1854);
and U8435 (N_8435,N_607,N_579);
nor U8436 (N_8436,N_4470,N_2697);
or U8437 (N_8437,N_4146,N_1465);
or U8438 (N_8438,N_3446,N_1847);
xnor U8439 (N_8439,N_3679,N_3399);
nor U8440 (N_8440,N_1624,N_2192);
and U8441 (N_8441,N_3785,N_4268);
and U8442 (N_8442,N_4647,N_2116);
nor U8443 (N_8443,N_720,N_2313);
and U8444 (N_8444,N_4770,N_1419);
or U8445 (N_8445,N_3556,N_975);
xnor U8446 (N_8446,N_4200,N_3200);
or U8447 (N_8447,N_3058,N_1963);
nand U8448 (N_8448,N_4849,N_2104);
nand U8449 (N_8449,N_2823,N_2325);
xor U8450 (N_8450,N_1894,N_4427);
nand U8451 (N_8451,N_496,N_3649);
and U8452 (N_8452,N_4707,N_497);
xnor U8453 (N_8453,N_1239,N_679);
xor U8454 (N_8454,N_2008,N_2066);
xor U8455 (N_8455,N_1530,N_3503);
nand U8456 (N_8456,N_2865,N_4295);
nor U8457 (N_8457,N_3932,N_4088);
and U8458 (N_8458,N_2159,N_300);
xor U8459 (N_8459,N_4752,N_4012);
xor U8460 (N_8460,N_1401,N_3161);
and U8461 (N_8461,N_3242,N_4363);
nor U8462 (N_8462,N_2267,N_821);
or U8463 (N_8463,N_174,N_559);
nand U8464 (N_8464,N_4342,N_600);
nor U8465 (N_8465,N_310,N_1104);
nor U8466 (N_8466,N_2651,N_1245);
and U8467 (N_8467,N_2813,N_4699);
and U8468 (N_8468,N_1212,N_4388);
xnor U8469 (N_8469,N_1647,N_2688);
nor U8470 (N_8470,N_577,N_2892);
nor U8471 (N_8471,N_195,N_79);
nor U8472 (N_8472,N_2182,N_3653);
xor U8473 (N_8473,N_4813,N_3503);
and U8474 (N_8474,N_744,N_1522);
or U8475 (N_8475,N_3765,N_2348);
nor U8476 (N_8476,N_1528,N_697);
or U8477 (N_8477,N_1080,N_2986);
nand U8478 (N_8478,N_4482,N_963);
or U8479 (N_8479,N_1889,N_3051);
xor U8480 (N_8480,N_3049,N_4860);
or U8481 (N_8481,N_2342,N_1726);
and U8482 (N_8482,N_4603,N_1629);
nand U8483 (N_8483,N_1423,N_4635);
and U8484 (N_8484,N_2253,N_485);
nand U8485 (N_8485,N_4116,N_4428);
nor U8486 (N_8486,N_2051,N_994);
xnor U8487 (N_8487,N_3584,N_3412);
nor U8488 (N_8488,N_1026,N_3739);
xnor U8489 (N_8489,N_3230,N_4432);
xnor U8490 (N_8490,N_3149,N_366);
xnor U8491 (N_8491,N_2913,N_3262);
nor U8492 (N_8492,N_4628,N_1765);
and U8493 (N_8493,N_573,N_2330);
nand U8494 (N_8494,N_2146,N_3769);
and U8495 (N_8495,N_4826,N_4866);
and U8496 (N_8496,N_2930,N_294);
nand U8497 (N_8497,N_3051,N_3563);
nand U8498 (N_8498,N_2726,N_261);
nand U8499 (N_8499,N_411,N_4309);
nor U8500 (N_8500,N_4939,N_2190);
nor U8501 (N_8501,N_1387,N_977);
or U8502 (N_8502,N_3216,N_2425);
xor U8503 (N_8503,N_1808,N_2043);
and U8504 (N_8504,N_233,N_3608);
or U8505 (N_8505,N_4285,N_1441);
or U8506 (N_8506,N_2275,N_2450);
and U8507 (N_8507,N_128,N_4168);
xnor U8508 (N_8508,N_3824,N_661);
or U8509 (N_8509,N_1790,N_3509);
xnor U8510 (N_8510,N_3293,N_3075);
and U8511 (N_8511,N_1610,N_3358);
and U8512 (N_8512,N_1860,N_845);
and U8513 (N_8513,N_2856,N_2343);
or U8514 (N_8514,N_841,N_4605);
nor U8515 (N_8515,N_2920,N_4248);
and U8516 (N_8516,N_192,N_4272);
nor U8517 (N_8517,N_4276,N_2564);
nor U8518 (N_8518,N_1740,N_898);
or U8519 (N_8519,N_4259,N_3368);
xor U8520 (N_8520,N_3811,N_2263);
and U8521 (N_8521,N_3898,N_1437);
nand U8522 (N_8522,N_1408,N_3714);
xor U8523 (N_8523,N_2329,N_4135);
xor U8524 (N_8524,N_493,N_3540);
nand U8525 (N_8525,N_4629,N_318);
or U8526 (N_8526,N_3092,N_4284);
nor U8527 (N_8527,N_1716,N_4589);
xnor U8528 (N_8528,N_3605,N_4911);
xnor U8529 (N_8529,N_4258,N_3087);
and U8530 (N_8530,N_2224,N_4057);
or U8531 (N_8531,N_3192,N_791);
xor U8532 (N_8532,N_3461,N_3031);
xor U8533 (N_8533,N_1124,N_2121);
nor U8534 (N_8534,N_4671,N_3838);
or U8535 (N_8535,N_3001,N_2596);
xnor U8536 (N_8536,N_2773,N_1);
xor U8537 (N_8537,N_2180,N_4711);
xor U8538 (N_8538,N_4755,N_441);
and U8539 (N_8539,N_635,N_629);
or U8540 (N_8540,N_3674,N_3197);
and U8541 (N_8541,N_3092,N_1997);
or U8542 (N_8542,N_1299,N_4561);
nor U8543 (N_8543,N_1778,N_608);
nand U8544 (N_8544,N_3573,N_908);
xnor U8545 (N_8545,N_1750,N_3611);
nand U8546 (N_8546,N_1485,N_1069);
or U8547 (N_8547,N_1490,N_3504);
and U8548 (N_8548,N_4213,N_1890);
and U8549 (N_8549,N_4667,N_264);
nand U8550 (N_8550,N_2883,N_684);
nor U8551 (N_8551,N_3126,N_4415);
and U8552 (N_8552,N_46,N_1207);
nand U8553 (N_8553,N_4630,N_2164);
or U8554 (N_8554,N_3159,N_3838);
nor U8555 (N_8555,N_4111,N_3382);
xor U8556 (N_8556,N_2087,N_1352);
nand U8557 (N_8557,N_741,N_724);
nor U8558 (N_8558,N_3100,N_2560);
nand U8559 (N_8559,N_3478,N_1976);
nor U8560 (N_8560,N_1475,N_4498);
nor U8561 (N_8561,N_2243,N_3636);
nor U8562 (N_8562,N_2963,N_2402);
nor U8563 (N_8563,N_813,N_3349);
and U8564 (N_8564,N_4805,N_157);
nand U8565 (N_8565,N_2314,N_853);
nor U8566 (N_8566,N_3686,N_3775);
and U8567 (N_8567,N_1666,N_4783);
nor U8568 (N_8568,N_1675,N_4319);
xor U8569 (N_8569,N_2684,N_3420);
and U8570 (N_8570,N_3081,N_557);
xnor U8571 (N_8571,N_3155,N_865);
or U8572 (N_8572,N_4941,N_3446);
xnor U8573 (N_8573,N_3926,N_4573);
and U8574 (N_8574,N_2786,N_3934);
xor U8575 (N_8575,N_4398,N_2688);
or U8576 (N_8576,N_1888,N_784);
or U8577 (N_8577,N_1907,N_535);
or U8578 (N_8578,N_4263,N_3654);
or U8579 (N_8579,N_79,N_2783);
xnor U8580 (N_8580,N_4536,N_2816);
and U8581 (N_8581,N_4509,N_3643);
and U8582 (N_8582,N_375,N_4866);
nand U8583 (N_8583,N_3983,N_851);
xor U8584 (N_8584,N_2759,N_898);
and U8585 (N_8585,N_2715,N_3327);
nand U8586 (N_8586,N_161,N_2093);
nor U8587 (N_8587,N_1823,N_631);
xnor U8588 (N_8588,N_4944,N_2782);
nand U8589 (N_8589,N_1080,N_3490);
nand U8590 (N_8590,N_3036,N_2798);
xor U8591 (N_8591,N_4056,N_1339);
xor U8592 (N_8592,N_525,N_1125);
xnor U8593 (N_8593,N_2864,N_2791);
xnor U8594 (N_8594,N_2899,N_3831);
and U8595 (N_8595,N_3534,N_777);
nor U8596 (N_8596,N_2097,N_2854);
nor U8597 (N_8597,N_3653,N_2646);
and U8598 (N_8598,N_4598,N_250);
nor U8599 (N_8599,N_4084,N_1383);
xnor U8600 (N_8600,N_930,N_3988);
xor U8601 (N_8601,N_2074,N_4075);
nand U8602 (N_8602,N_4902,N_1572);
and U8603 (N_8603,N_1330,N_2609);
and U8604 (N_8604,N_2141,N_3158);
or U8605 (N_8605,N_1380,N_2525);
or U8606 (N_8606,N_2188,N_2891);
nand U8607 (N_8607,N_3571,N_2320);
nand U8608 (N_8608,N_1793,N_269);
nand U8609 (N_8609,N_3609,N_3130);
or U8610 (N_8610,N_263,N_1546);
nor U8611 (N_8611,N_2175,N_2443);
nand U8612 (N_8612,N_4822,N_1579);
nand U8613 (N_8613,N_3926,N_2596);
xnor U8614 (N_8614,N_3414,N_419);
nand U8615 (N_8615,N_1977,N_1698);
xor U8616 (N_8616,N_3378,N_1224);
xor U8617 (N_8617,N_3417,N_213);
xnor U8618 (N_8618,N_3891,N_3134);
and U8619 (N_8619,N_1221,N_371);
nand U8620 (N_8620,N_1796,N_1846);
and U8621 (N_8621,N_3928,N_4947);
xnor U8622 (N_8622,N_634,N_1798);
and U8623 (N_8623,N_3887,N_3927);
nand U8624 (N_8624,N_1385,N_1355);
xor U8625 (N_8625,N_3054,N_540);
xnor U8626 (N_8626,N_1508,N_2015);
nand U8627 (N_8627,N_2535,N_435);
nor U8628 (N_8628,N_513,N_2217);
or U8629 (N_8629,N_2221,N_38);
nand U8630 (N_8630,N_2932,N_2134);
or U8631 (N_8631,N_521,N_514);
and U8632 (N_8632,N_3430,N_327);
nand U8633 (N_8633,N_3492,N_1627);
xor U8634 (N_8634,N_2406,N_4330);
nand U8635 (N_8635,N_4589,N_490);
nand U8636 (N_8636,N_3007,N_4431);
nor U8637 (N_8637,N_2925,N_4683);
and U8638 (N_8638,N_1880,N_1580);
nand U8639 (N_8639,N_2466,N_1516);
xor U8640 (N_8640,N_3528,N_4795);
and U8641 (N_8641,N_635,N_2893);
nor U8642 (N_8642,N_1276,N_3024);
nor U8643 (N_8643,N_2613,N_1644);
or U8644 (N_8644,N_4921,N_550);
and U8645 (N_8645,N_710,N_1333);
xnor U8646 (N_8646,N_2753,N_1524);
xnor U8647 (N_8647,N_4259,N_4301);
and U8648 (N_8648,N_4384,N_1132);
nor U8649 (N_8649,N_3053,N_2382);
nand U8650 (N_8650,N_2029,N_3777);
or U8651 (N_8651,N_258,N_4613);
nand U8652 (N_8652,N_1557,N_3646);
and U8653 (N_8653,N_573,N_2348);
nand U8654 (N_8654,N_4794,N_1978);
or U8655 (N_8655,N_2717,N_2272);
xor U8656 (N_8656,N_1669,N_102);
or U8657 (N_8657,N_3824,N_2314);
or U8658 (N_8658,N_2463,N_157);
and U8659 (N_8659,N_4634,N_1201);
nor U8660 (N_8660,N_640,N_1474);
or U8661 (N_8661,N_414,N_3246);
nand U8662 (N_8662,N_2671,N_1727);
nor U8663 (N_8663,N_4893,N_2576);
and U8664 (N_8664,N_3691,N_2993);
or U8665 (N_8665,N_82,N_145);
nand U8666 (N_8666,N_582,N_3822);
nor U8667 (N_8667,N_2323,N_1024);
and U8668 (N_8668,N_4947,N_1449);
nand U8669 (N_8669,N_3478,N_3342);
xor U8670 (N_8670,N_1445,N_2737);
xnor U8671 (N_8671,N_3851,N_4778);
nand U8672 (N_8672,N_1152,N_4140);
nor U8673 (N_8673,N_595,N_2843);
nor U8674 (N_8674,N_3309,N_1817);
nand U8675 (N_8675,N_3168,N_830);
and U8676 (N_8676,N_3969,N_866);
nor U8677 (N_8677,N_3941,N_2028);
nand U8678 (N_8678,N_3709,N_28);
xnor U8679 (N_8679,N_1208,N_1781);
nand U8680 (N_8680,N_3175,N_2279);
nor U8681 (N_8681,N_2094,N_3594);
or U8682 (N_8682,N_690,N_819);
or U8683 (N_8683,N_4650,N_1162);
xor U8684 (N_8684,N_3773,N_2489);
xor U8685 (N_8685,N_2040,N_2894);
or U8686 (N_8686,N_3090,N_3515);
nor U8687 (N_8687,N_72,N_3455);
or U8688 (N_8688,N_9,N_1271);
and U8689 (N_8689,N_880,N_307);
or U8690 (N_8690,N_722,N_130);
nand U8691 (N_8691,N_4558,N_2502);
nor U8692 (N_8692,N_769,N_3666);
or U8693 (N_8693,N_1763,N_2161);
and U8694 (N_8694,N_4542,N_2841);
or U8695 (N_8695,N_3119,N_4168);
xor U8696 (N_8696,N_4974,N_2380);
nor U8697 (N_8697,N_3574,N_4701);
or U8698 (N_8698,N_15,N_2228);
or U8699 (N_8699,N_4063,N_2138);
nand U8700 (N_8700,N_800,N_1240);
and U8701 (N_8701,N_2173,N_3103);
nand U8702 (N_8702,N_2020,N_1772);
xnor U8703 (N_8703,N_1513,N_2937);
nor U8704 (N_8704,N_1038,N_4167);
or U8705 (N_8705,N_2188,N_4077);
or U8706 (N_8706,N_1064,N_1794);
xnor U8707 (N_8707,N_3269,N_3727);
nand U8708 (N_8708,N_3376,N_697);
nor U8709 (N_8709,N_596,N_4709);
or U8710 (N_8710,N_2539,N_2997);
nand U8711 (N_8711,N_2680,N_2856);
xor U8712 (N_8712,N_251,N_2014);
and U8713 (N_8713,N_4715,N_4281);
or U8714 (N_8714,N_2267,N_4776);
nor U8715 (N_8715,N_4683,N_2262);
xnor U8716 (N_8716,N_4329,N_1539);
or U8717 (N_8717,N_1079,N_3559);
nand U8718 (N_8718,N_1797,N_369);
and U8719 (N_8719,N_4848,N_4194);
and U8720 (N_8720,N_3995,N_4617);
or U8721 (N_8721,N_1568,N_3889);
nor U8722 (N_8722,N_2473,N_3161);
or U8723 (N_8723,N_2453,N_1079);
nor U8724 (N_8724,N_3451,N_2526);
xor U8725 (N_8725,N_3314,N_3948);
xnor U8726 (N_8726,N_2873,N_4472);
or U8727 (N_8727,N_3194,N_524);
nor U8728 (N_8728,N_153,N_2479);
and U8729 (N_8729,N_42,N_3542);
nand U8730 (N_8730,N_1506,N_1544);
or U8731 (N_8731,N_16,N_230);
xnor U8732 (N_8732,N_2955,N_3280);
or U8733 (N_8733,N_3596,N_2652);
or U8734 (N_8734,N_1487,N_2209);
or U8735 (N_8735,N_4047,N_4730);
nand U8736 (N_8736,N_4427,N_4820);
nor U8737 (N_8737,N_1760,N_320);
xnor U8738 (N_8738,N_628,N_2120);
or U8739 (N_8739,N_4395,N_3503);
nand U8740 (N_8740,N_3985,N_3163);
nor U8741 (N_8741,N_3661,N_1720);
and U8742 (N_8742,N_4344,N_3734);
or U8743 (N_8743,N_4321,N_731);
nor U8744 (N_8744,N_4680,N_4127);
and U8745 (N_8745,N_1435,N_3733);
nor U8746 (N_8746,N_2905,N_738);
and U8747 (N_8747,N_4516,N_4937);
xnor U8748 (N_8748,N_191,N_3753);
xor U8749 (N_8749,N_4507,N_1435);
nand U8750 (N_8750,N_1485,N_2321);
nand U8751 (N_8751,N_1924,N_1545);
nand U8752 (N_8752,N_4226,N_2260);
xor U8753 (N_8753,N_3724,N_95);
nand U8754 (N_8754,N_303,N_1632);
nand U8755 (N_8755,N_3522,N_974);
nand U8756 (N_8756,N_3846,N_1942);
nor U8757 (N_8757,N_458,N_2126);
nand U8758 (N_8758,N_770,N_1525);
xnor U8759 (N_8759,N_3396,N_4492);
nor U8760 (N_8760,N_1851,N_2451);
or U8761 (N_8761,N_448,N_3978);
xnor U8762 (N_8762,N_3301,N_3109);
nand U8763 (N_8763,N_3357,N_2449);
nand U8764 (N_8764,N_2408,N_1618);
nand U8765 (N_8765,N_3275,N_3580);
xnor U8766 (N_8766,N_665,N_3496);
and U8767 (N_8767,N_67,N_3278);
nand U8768 (N_8768,N_1173,N_3762);
or U8769 (N_8769,N_1489,N_3046);
xnor U8770 (N_8770,N_4317,N_1785);
and U8771 (N_8771,N_4134,N_3026);
nor U8772 (N_8772,N_1759,N_4783);
and U8773 (N_8773,N_1046,N_4726);
nor U8774 (N_8774,N_3066,N_1829);
nor U8775 (N_8775,N_4905,N_910);
nand U8776 (N_8776,N_3402,N_760);
nand U8777 (N_8777,N_1856,N_4420);
and U8778 (N_8778,N_3373,N_1351);
nand U8779 (N_8779,N_1368,N_994);
and U8780 (N_8780,N_3198,N_3204);
xnor U8781 (N_8781,N_746,N_3201);
or U8782 (N_8782,N_3265,N_2609);
nand U8783 (N_8783,N_3539,N_3083);
or U8784 (N_8784,N_1689,N_2420);
xor U8785 (N_8785,N_2612,N_4909);
and U8786 (N_8786,N_83,N_1497);
and U8787 (N_8787,N_3995,N_1249);
xor U8788 (N_8788,N_1776,N_1333);
or U8789 (N_8789,N_3423,N_4693);
or U8790 (N_8790,N_1570,N_1851);
and U8791 (N_8791,N_3200,N_1443);
xor U8792 (N_8792,N_4395,N_1059);
and U8793 (N_8793,N_3048,N_3356);
and U8794 (N_8794,N_4525,N_1515);
or U8795 (N_8795,N_4829,N_1333);
nand U8796 (N_8796,N_257,N_2261);
nor U8797 (N_8797,N_507,N_1993);
xor U8798 (N_8798,N_1121,N_395);
nor U8799 (N_8799,N_994,N_4052);
or U8800 (N_8800,N_4236,N_3265);
nor U8801 (N_8801,N_1273,N_3327);
xor U8802 (N_8802,N_1824,N_720);
nand U8803 (N_8803,N_1610,N_602);
and U8804 (N_8804,N_3807,N_785);
xnor U8805 (N_8805,N_2098,N_353);
and U8806 (N_8806,N_684,N_4392);
nand U8807 (N_8807,N_2667,N_2391);
nand U8808 (N_8808,N_4437,N_3190);
and U8809 (N_8809,N_3288,N_1357);
or U8810 (N_8810,N_4823,N_2811);
or U8811 (N_8811,N_4548,N_3307);
nor U8812 (N_8812,N_635,N_877);
nor U8813 (N_8813,N_2687,N_1277);
or U8814 (N_8814,N_2220,N_344);
xnor U8815 (N_8815,N_4601,N_4024);
nand U8816 (N_8816,N_3833,N_2888);
nand U8817 (N_8817,N_1329,N_821);
nand U8818 (N_8818,N_1234,N_3682);
xor U8819 (N_8819,N_1042,N_4580);
nor U8820 (N_8820,N_883,N_3991);
and U8821 (N_8821,N_4147,N_2981);
and U8822 (N_8822,N_436,N_793);
xnor U8823 (N_8823,N_2400,N_406);
nand U8824 (N_8824,N_4731,N_1118);
and U8825 (N_8825,N_3423,N_3048);
xor U8826 (N_8826,N_198,N_792);
or U8827 (N_8827,N_2815,N_1300);
and U8828 (N_8828,N_4121,N_118);
nand U8829 (N_8829,N_2684,N_864);
xor U8830 (N_8830,N_2318,N_3607);
nor U8831 (N_8831,N_1163,N_1957);
or U8832 (N_8832,N_3163,N_1257);
or U8833 (N_8833,N_1331,N_4867);
and U8834 (N_8834,N_1537,N_1662);
nand U8835 (N_8835,N_3055,N_3751);
xor U8836 (N_8836,N_3530,N_4598);
and U8837 (N_8837,N_4105,N_2958);
xnor U8838 (N_8838,N_3883,N_5);
nor U8839 (N_8839,N_1762,N_399);
xor U8840 (N_8840,N_2134,N_2803);
nor U8841 (N_8841,N_2375,N_1343);
nor U8842 (N_8842,N_2022,N_755);
xor U8843 (N_8843,N_3632,N_2161);
nor U8844 (N_8844,N_1110,N_162);
nor U8845 (N_8845,N_2266,N_837);
xnor U8846 (N_8846,N_504,N_3785);
and U8847 (N_8847,N_2273,N_3638);
xnor U8848 (N_8848,N_2090,N_4196);
nor U8849 (N_8849,N_1107,N_2133);
xor U8850 (N_8850,N_1125,N_4190);
and U8851 (N_8851,N_4957,N_4280);
or U8852 (N_8852,N_4313,N_4087);
and U8853 (N_8853,N_4818,N_4821);
nor U8854 (N_8854,N_1854,N_2610);
and U8855 (N_8855,N_297,N_3848);
nor U8856 (N_8856,N_2228,N_89);
xor U8857 (N_8857,N_2256,N_1811);
and U8858 (N_8858,N_3823,N_1727);
nor U8859 (N_8859,N_1491,N_4303);
or U8860 (N_8860,N_3280,N_4433);
xor U8861 (N_8861,N_3748,N_1343);
nand U8862 (N_8862,N_3923,N_1211);
and U8863 (N_8863,N_4165,N_510);
or U8864 (N_8864,N_2425,N_2294);
xnor U8865 (N_8865,N_2713,N_4134);
or U8866 (N_8866,N_2912,N_1143);
nand U8867 (N_8867,N_3014,N_920);
xor U8868 (N_8868,N_557,N_3009);
xnor U8869 (N_8869,N_1627,N_1089);
or U8870 (N_8870,N_4,N_3777);
or U8871 (N_8871,N_4474,N_4391);
nand U8872 (N_8872,N_4343,N_4665);
nand U8873 (N_8873,N_3617,N_4171);
nand U8874 (N_8874,N_2666,N_4327);
and U8875 (N_8875,N_1889,N_1079);
or U8876 (N_8876,N_4853,N_4293);
or U8877 (N_8877,N_4591,N_1125);
or U8878 (N_8878,N_2678,N_409);
nand U8879 (N_8879,N_4982,N_1310);
and U8880 (N_8880,N_4717,N_1903);
and U8881 (N_8881,N_2159,N_4422);
xnor U8882 (N_8882,N_3990,N_1372);
or U8883 (N_8883,N_2201,N_3821);
and U8884 (N_8884,N_4848,N_897);
or U8885 (N_8885,N_4696,N_2249);
xnor U8886 (N_8886,N_4554,N_4274);
xor U8887 (N_8887,N_2941,N_465);
nand U8888 (N_8888,N_2104,N_1060);
or U8889 (N_8889,N_1368,N_3804);
nand U8890 (N_8890,N_3882,N_2255);
or U8891 (N_8891,N_2105,N_854);
nor U8892 (N_8892,N_350,N_2412);
or U8893 (N_8893,N_3062,N_3681);
and U8894 (N_8894,N_1523,N_2142);
nor U8895 (N_8895,N_1157,N_287);
or U8896 (N_8896,N_3712,N_1826);
nor U8897 (N_8897,N_1835,N_585);
xnor U8898 (N_8898,N_4959,N_168);
nand U8899 (N_8899,N_2258,N_1254);
nor U8900 (N_8900,N_2494,N_3624);
nand U8901 (N_8901,N_2202,N_1169);
or U8902 (N_8902,N_1311,N_3214);
and U8903 (N_8903,N_2836,N_4797);
or U8904 (N_8904,N_624,N_1211);
nand U8905 (N_8905,N_3134,N_3225);
nor U8906 (N_8906,N_2168,N_1357);
or U8907 (N_8907,N_3498,N_4488);
and U8908 (N_8908,N_1384,N_4792);
nand U8909 (N_8909,N_4183,N_1984);
xor U8910 (N_8910,N_3479,N_3682);
and U8911 (N_8911,N_3298,N_4829);
or U8912 (N_8912,N_2423,N_3919);
nand U8913 (N_8913,N_1677,N_4485);
nor U8914 (N_8914,N_4301,N_4224);
xnor U8915 (N_8915,N_2760,N_526);
nand U8916 (N_8916,N_377,N_2036);
nand U8917 (N_8917,N_812,N_3451);
or U8918 (N_8918,N_2995,N_1086);
nand U8919 (N_8919,N_4075,N_2757);
nor U8920 (N_8920,N_297,N_763);
or U8921 (N_8921,N_3855,N_1315);
or U8922 (N_8922,N_716,N_39);
or U8923 (N_8923,N_365,N_4959);
and U8924 (N_8924,N_473,N_818);
xor U8925 (N_8925,N_1826,N_818);
nand U8926 (N_8926,N_2866,N_4141);
nor U8927 (N_8927,N_2043,N_3391);
nand U8928 (N_8928,N_1796,N_3693);
nand U8929 (N_8929,N_2157,N_1928);
nand U8930 (N_8930,N_4892,N_2676);
nand U8931 (N_8931,N_3786,N_2945);
or U8932 (N_8932,N_343,N_3491);
or U8933 (N_8933,N_4613,N_3249);
xor U8934 (N_8934,N_1328,N_4236);
or U8935 (N_8935,N_663,N_3665);
or U8936 (N_8936,N_3691,N_3377);
nand U8937 (N_8937,N_3055,N_1859);
xor U8938 (N_8938,N_4214,N_4292);
or U8939 (N_8939,N_3075,N_1608);
nor U8940 (N_8940,N_3641,N_3743);
or U8941 (N_8941,N_169,N_4875);
and U8942 (N_8942,N_1309,N_1223);
nor U8943 (N_8943,N_2390,N_3080);
and U8944 (N_8944,N_287,N_1142);
or U8945 (N_8945,N_2653,N_3438);
and U8946 (N_8946,N_3177,N_4754);
nand U8947 (N_8947,N_153,N_2042);
nor U8948 (N_8948,N_4104,N_3656);
and U8949 (N_8949,N_935,N_4226);
or U8950 (N_8950,N_2174,N_4646);
or U8951 (N_8951,N_3153,N_1084);
and U8952 (N_8952,N_2518,N_3260);
or U8953 (N_8953,N_1495,N_4604);
nor U8954 (N_8954,N_2698,N_3775);
nor U8955 (N_8955,N_1420,N_4352);
nor U8956 (N_8956,N_3204,N_4336);
nand U8957 (N_8957,N_2137,N_4783);
and U8958 (N_8958,N_3656,N_2242);
nor U8959 (N_8959,N_2484,N_2556);
and U8960 (N_8960,N_3861,N_2785);
and U8961 (N_8961,N_4887,N_2579);
nor U8962 (N_8962,N_4361,N_2384);
and U8963 (N_8963,N_981,N_952);
nor U8964 (N_8964,N_1937,N_3991);
nand U8965 (N_8965,N_3624,N_3155);
nor U8966 (N_8966,N_4217,N_3418);
nor U8967 (N_8967,N_679,N_1125);
nand U8968 (N_8968,N_683,N_1759);
nand U8969 (N_8969,N_225,N_4245);
and U8970 (N_8970,N_832,N_3010);
and U8971 (N_8971,N_4847,N_731);
and U8972 (N_8972,N_230,N_2695);
nand U8973 (N_8973,N_4898,N_4685);
and U8974 (N_8974,N_1258,N_3710);
xor U8975 (N_8975,N_427,N_2208);
xnor U8976 (N_8976,N_919,N_4906);
nor U8977 (N_8977,N_2710,N_1038);
nor U8978 (N_8978,N_1005,N_3494);
nand U8979 (N_8979,N_1273,N_3073);
or U8980 (N_8980,N_1677,N_4034);
or U8981 (N_8981,N_4161,N_2646);
nand U8982 (N_8982,N_3993,N_3120);
xor U8983 (N_8983,N_574,N_2324);
and U8984 (N_8984,N_2590,N_4788);
nand U8985 (N_8985,N_3403,N_2125);
or U8986 (N_8986,N_65,N_2545);
xor U8987 (N_8987,N_4507,N_1831);
nor U8988 (N_8988,N_2611,N_741);
nor U8989 (N_8989,N_2676,N_1368);
and U8990 (N_8990,N_223,N_3182);
or U8991 (N_8991,N_4632,N_1796);
and U8992 (N_8992,N_2221,N_203);
xor U8993 (N_8993,N_536,N_559);
xnor U8994 (N_8994,N_2935,N_451);
or U8995 (N_8995,N_3011,N_943);
and U8996 (N_8996,N_3001,N_1348);
or U8997 (N_8997,N_1355,N_4596);
nor U8998 (N_8998,N_2031,N_3241);
and U8999 (N_8999,N_1000,N_883);
and U9000 (N_9000,N_1995,N_2610);
and U9001 (N_9001,N_2061,N_3540);
and U9002 (N_9002,N_1171,N_2379);
nand U9003 (N_9003,N_2775,N_3149);
and U9004 (N_9004,N_2812,N_2941);
nand U9005 (N_9005,N_747,N_3004);
and U9006 (N_9006,N_900,N_4007);
and U9007 (N_9007,N_2966,N_3853);
nand U9008 (N_9008,N_2774,N_2530);
or U9009 (N_9009,N_198,N_4697);
nand U9010 (N_9010,N_1107,N_1937);
or U9011 (N_9011,N_1681,N_445);
nand U9012 (N_9012,N_344,N_24);
or U9013 (N_9013,N_2955,N_854);
and U9014 (N_9014,N_3344,N_1284);
nand U9015 (N_9015,N_1554,N_229);
or U9016 (N_9016,N_3461,N_2805);
nor U9017 (N_9017,N_612,N_712);
xnor U9018 (N_9018,N_2927,N_2811);
xor U9019 (N_9019,N_1811,N_824);
or U9020 (N_9020,N_1015,N_2781);
nand U9021 (N_9021,N_581,N_3691);
xnor U9022 (N_9022,N_1431,N_2032);
nand U9023 (N_9023,N_1283,N_1687);
or U9024 (N_9024,N_116,N_445);
nor U9025 (N_9025,N_2704,N_4891);
nand U9026 (N_9026,N_531,N_11);
nor U9027 (N_9027,N_1873,N_2172);
or U9028 (N_9028,N_2894,N_3878);
or U9029 (N_9029,N_3659,N_3520);
and U9030 (N_9030,N_1684,N_1429);
and U9031 (N_9031,N_198,N_2453);
and U9032 (N_9032,N_4547,N_1565);
and U9033 (N_9033,N_755,N_3645);
xnor U9034 (N_9034,N_2086,N_2700);
nor U9035 (N_9035,N_4392,N_1519);
nand U9036 (N_9036,N_4315,N_772);
nor U9037 (N_9037,N_936,N_4020);
nand U9038 (N_9038,N_1893,N_298);
xnor U9039 (N_9039,N_4511,N_4177);
or U9040 (N_9040,N_236,N_1980);
or U9041 (N_9041,N_3634,N_1683);
xor U9042 (N_9042,N_291,N_2692);
and U9043 (N_9043,N_1535,N_4401);
nand U9044 (N_9044,N_600,N_649);
or U9045 (N_9045,N_1559,N_808);
nand U9046 (N_9046,N_921,N_1612);
nor U9047 (N_9047,N_397,N_3616);
and U9048 (N_9048,N_698,N_3192);
xnor U9049 (N_9049,N_794,N_558);
or U9050 (N_9050,N_2464,N_4045);
or U9051 (N_9051,N_4788,N_2871);
nand U9052 (N_9052,N_229,N_1201);
and U9053 (N_9053,N_2946,N_2292);
xnor U9054 (N_9054,N_3370,N_3728);
xor U9055 (N_9055,N_1644,N_574);
nand U9056 (N_9056,N_1497,N_1391);
xor U9057 (N_9057,N_1051,N_4817);
xnor U9058 (N_9058,N_1707,N_3262);
nor U9059 (N_9059,N_1224,N_1124);
nand U9060 (N_9060,N_2867,N_1216);
and U9061 (N_9061,N_2644,N_2491);
nor U9062 (N_9062,N_961,N_52);
nor U9063 (N_9063,N_2911,N_1198);
xnor U9064 (N_9064,N_248,N_4948);
nand U9065 (N_9065,N_323,N_3146);
nor U9066 (N_9066,N_1201,N_1820);
nor U9067 (N_9067,N_4025,N_2272);
and U9068 (N_9068,N_3055,N_843);
and U9069 (N_9069,N_1125,N_1941);
xnor U9070 (N_9070,N_3224,N_4003);
and U9071 (N_9071,N_4031,N_3922);
or U9072 (N_9072,N_3122,N_220);
or U9073 (N_9073,N_1158,N_3007);
or U9074 (N_9074,N_580,N_4753);
nand U9075 (N_9075,N_3552,N_4417);
and U9076 (N_9076,N_499,N_3627);
xor U9077 (N_9077,N_3098,N_1910);
nand U9078 (N_9078,N_2812,N_4190);
or U9079 (N_9079,N_3225,N_105);
and U9080 (N_9080,N_714,N_84);
and U9081 (N_9081,N_105,N_4362);
nor U9082 (N_9082,N_3807,N_1099);
and U9083 (N_9083,N_4510,N_1065);
or U9084 (N_9084,N_2878,N_1139);
xor U9085 (N_9085,N_755,N_565);
nor U9086 (N_9086,N_4950,N_632);
or U9087 (N_9087,N_234,N_1473);
or U9088 (N_9088,N_3382,N_1016);
or U9089 (N_9089,N_1395,N_2160);
xnor U9090 (N_9090,N_1182,N_3106);
and U9091 (N_9091,N_2415,N_179);
xnor U9092 (N_9092,N_3653,N_3155);
or U9093 (N_9093,N_2498,N_3619);
xnor U9094 (N_9094,N_2528,N_4075);
xor U9095 (N_9095,N_778,N_1483);
nor U9096 (N_9096,N_106,N_1209);
xnor U9097 (N_9097,N_3277,N_640);
and U9098 (N_9098,N_666,N_4733);
and U9099 (N_9099,N_2473,N_3341);
nand U9100 (N_9100,N_3310,N_1669);
xor U9101 (N_9101,N_2886,N_574);
nand U9102 (N_9102,N_995,N_3068);
or U9103 (N_9103,N_554,N_1831);
nand U9104 (N_9104,N_2532,N_3470);
and U9105 (N_9105,N_2043,N_1074);
and U9106 (N_9106,N_1308,N_4067);
nand U9107 (N_9107,N_2001,N_2729);
xnor U9108 (N_9108,N_2699,N_2885);
nor U9109 (N_9109,N_3841,N_4223);
nor U9110 (N_9110,N_2644,N_1998);
nor U9111 (N_9111,N_4407,N_1130);
nor U9112 (N_9112,N_2558,N_4182);
or U9113 (N_9113,N_2254,N_4783);
and U9114 (N_9114,N_121,N_2356);
nand U9115 (N_9115,N_1736,N_1100);
xnor U9116 (N_9116,N_1309,N_2124);
nand U9117 (N_9117,N_4983,N_4868);
xnor U9118 (N_9118,N_1364,N_1154);
nor U9119 (N_9119,N_4644,N_3294);
nand U9120 (N_9120,N_3617,N_2122);
xnor U9121 (N_9121,N_3779,N_4959);
and U9122 (N_9122,N_2135,N_3324);
nor U9123 (N_9123,N_3371,N_2114);
nor U9124 (N_9124,N_4338,N_3516);
and U9125 (N_9125,N_3316,N_3994);
nand U9126 (N_9126,N_0,N_3884);
xnor U9127 (N_9127,N_3691,N_2051);
xor U9128 (N_9128,N_3318,N_105);
nor U9129 (N_9129,N_2598,N_528);
xnor U9130 (N_9130,N_3708,N_3679);
and U9131 (N_9131,N_866,N_2992);
nand U9132 (N_9132,N_4419,N_3916);
or U9133 (N_9133,N_834,N_3390);
nand U9134 (N_9134,N_684,N_1176);
nor U9135 (N_9135,N_4858,N_2265);
and U9136 (N_9136,N_2928,N_4829);
and U9137 (N_9137,N_376,N_766);
xnor U9138 (N_9138,N_4386,N_3760);
nand U9139 (N_9139,N_2484,N_4068);
nand U9140 (N_9140,N_256,N_2446);
or U9141 (N_9141,N_3502,N_1420);
nor U9142 (N_9142,N_760,N_3407);
xor U9143 (N_9143,N_451,N_4301);
nand U9144 (N_9144,N_2751,N_4388);
and U9145 (N_9145,N_1594,N_654);
nor U9146 (N_9146,N_764,N_3421);
and U9147 (N_9147,N_1286,N_3905);
nand U9148 (N_9148,N_1924,N_1980);
or U9149 (N_9149,N_1927,N_695);
or U9150 (N_9150,N_238,N_2537);
nor U9151 (N_9151,N_1259,N_2798);
nor U9152 (N_9152,N_1286,N_2554);
and U9153 (N_9153,N_3294,N_247);
and U9154 (N_9154,N_3581,N_2284);
xnor U9155 (N_9155,N_4531,N_745);
xnor U9156 (N_9156,N_3494,N_4558);
or U9157 (N_9157,N_2662,N_3571);
xnor U9158 (N_9158,N_3403,N_3326);
nor U9159 (N_9159,N_3786,N_1297);
nand U9160 (N_9160,N_1355,N_1792);
nand U9161 (N_9161,N_1026,N_3996);
nor U9162 (N_9162,N_2909,N_2845);
or U9163 (N_9163,N_4911,N_4375);
or U9164 (N_9164,N_3713,N_1824);
or U9165 (N_9165,N_4518,N_2350);
nor U9166 (N_9166,N_3514,N_1137);
or U9167 (N_9167,N_4730,N_828);
nor U9168 (N_9168,N_3418,N_2954);
and U9169 (N_9169,N_3146,N_1988);
or U9170 (N_9170,N_3214,N_2826);
nor U9171 (N_9171,N_2477,N_4558);
or U9172 (N_9172,N_3642,N_471);
and U9173 (N_9173,N_2438,N_2594);
xnor U9174 (N_9174,N_4923,N_4659);
and U9175 (N_9175,N_2707,N_910);
and U9176 (N_9176,N_1204,N_3542);
nor U9177 (N_9177,N_4281,N_3618);
nor U9178 (N_9178,N_4844,N_1609);
nor U9179 (N_9179,N_3395,N_6);
xnor U9180 (N_9180,N_3963,N_3065);
nor U9181 (N_9181,N_1459,N_4276);
xnor U9182 (N_9182,N_1917,N_4739);
nand U9183 (N_9183,N_3718,N_3357);
or U9184 (N_9184,N_4229,N_3121);
and U9185 (N_9185,N_385,N_118);
nor U9186 (N_9186,N_4212,N_4387);
nand U9187 (N_9187,N_2860,N_2121);
and U9188 (N_9188,N_31,N_439);
nand U9189 (N_9189,N_976,N_22);
nand U9190 (N_9190,N_4216,N_1500);
nand U9191 (N_9191,N_4793,N_2498);
nand U9192 (N_9192,N_2400,N_3180);
nand U9193 (N_9193,N_2963,N_3713);
or U9194 (N_9194,N_80,N_3845);
or U9195 (N_9195,N_803,N_2409);
xnor U9196 (N_9196,N_4175,N_4233);
or U9197 (N_9197,N_4844,N_1278);
xor U9198 (N_9198,N_357,N_3769);
nand U9199 (N_9199,N_2893,N_1145);
or U9200 (N_9200,N_4637,N_1069);
xnor U9201 (N_9201,N_1605,N_67);
nand U9202 (N_9202,N_4643,N_1439);
nor U9203 (N_9203,N_1868,N_1690);
nor U9204 (N_9204,N_940,N_3914);
and U9205 (N_9205,N_2393,N_2533);
and U9206 (N_9206,N_2225,N_267);
or U9207 (N_9207,N_4611,N_3545);
xnor U9208 (N_9208,N_2888,N_1000);
and U9209 (N_9209,N_3070,N_4471);
nor U9210 (N_9210,N_1308,N_2264);
or U9211 (N_9211,N_2697,N_3644);
nand U9212 (N_9212,N_3908,N_3489);
or U9213 (N_9213,N_995,N_2831);
or U9214 (N_9214,N_3552,N_4252);
xor U9215 (N_9215,N_637,N_1121);
nand U9216 (N_9216,N_3111,N_1231);
nor U9217 (N_9217,N_4404,N_1574);
and U9218 (N_9218,N_3108,N_415);
nand U9219 (N_9219,N_3002,N_2093);
nor U9220 (N_9220,N_3807,N_331);
nor U9221 (N_9221,N_881,N_1038);
xor U9222 (N_9222,N_1916,N_3224);
nor U9223 (N_9223,N_4250,N_2071);
nand U9224 (N_9224,N_1007,N_737);
nor U9225 (N_9225,N_4279,N_4559);
xor U9226 (N_9226,N_3625,N_4767);
and U9227 (N_9227,N_1086,N_2919);
or U9228 (N_9228,N_615,N_3322);
and U9229 (N_9229,N_1603,N_738);
xnor U9230 (N_9230,N_1437,N_3713);
or U9231 (N_9231,N_2361,N_2791);
nor U9232 (N_9232,N_618,N_2178);
or U9233 (N_9233,N_4010,N_675);
xor U9234 (N_9234,N_3832,N_1809);
nand U9235 (N_9235,N_4295,N_681);
xor U9236 (N_9236,N_1431,N_1083);
nand U9237 (N_9237,N_1124,N_699);
and U9238 (N_9238,N_1071,N_4037);
nor U9239 (N_9239,N_2932,N_3794);
xor U9240 (N_9240,N_3859,N_3714);
and U9241 (N_9241,N_2549,N_4882);
and U9242 (N_9242,N_4807,N_686);
or U9243 (N_9243,N_3236,N_2483);
or U9244 (N_9244,N_445,N_3396);
xnor U9245 (N_9245,N_3598,N_344);
xnor U9246 (N_9246,N_4641,N_91);
or U9247 (N_9247,N_843,N_481);
nand U9248 (N_9248,N_3878,N_3722);
nand U9249 (N_9249,N_4040,N_1274);
xor U9250 (N_9250,N_93,N_2546);
and U9251 (N_9251,N_4163,N_1764);
xnor U9252 (N_9252,N_2191,N_1752);
nand U9253 (N_9253,N_4086,N_2604);
and U9254 (N_9254,N_1554,N_1530);
xor U9255 (N_9255,N_1914,N_1638);
nor U9256 (N_9256,N_3868,N_3471);
nor U9257 (N_9257,N_240,N_688);
nor U9258 (N_9258,N_1822,N_3554);
or U9259 (N_9259,N_3043,N_2174);
xnor U9260 (N_9260,N_2890,N_3452);
and U9261 (N_9261,N_3258,N_1620);
and U9262 (N_9262,N_2916,N_211);
nor U9263 (N_9263,N_4323,N_4364);
nor U9264 (N_9264,N_1395,N_607);
and U9265 (N_9265,N_2608,N_1954);
xor U9266 (N_9266,N_4831,N_670);
nand U9267 (N_9267,N_505,N_247);
nand U9268 (N_9268,N_2778,N_3475);
xor U9269 (N_9269,N_1931,N_1602);
and U9270 (N_9270,N_3250,N_1489);
nand U9271 (N_9271,N_1961,N_2460);
xor U9272 (N_9272,N_4404,N_4460);
and U9273 (N_9273,N_1437,N_1885);
nand U9274 (N_9274,N_2349,N_4720);
nor U9275 (N_9275,N_367,N_4003);
and U9276 (N_9276,N_4497,N_1278);
xnor U9277 (N_9277,N_4980,N_2599);
nor U9278 (N_9278,N_316,N_2014);
xor U9279 (N_9279,N_1574,N_1336);
nor U9280 (N_9280,N_429,N_4841);
nand U9281 (N_9281,N_2655,N_3455);
xnor U9282 (N_9282,N_3725,N_3145);
xnor U9283 (N_9283,N_4289,N_1876);
xor U9284 (N_9284,N_743,N_440);
nor U9285 (N_9285,N_1500,N_1621);
and U9286 (N_9286,N_1916,N_349);
nand U9287 (N_9287,N_2012,N_4738);
or U9288 (N_9288,N_2337,N_2994);
xnor U9289 (N_9289,N_4680,N_4634);
nand U9290 (N_9290,N_1122,N_4283);
nand U9291 (N_9291,N_4277,N_997);
xnor U9292 (N_9292,N_86,N_2386);
and U9293 (N_9293,N_2420,N_3469);
nor U9294 (N_9294,N_578,N_4122);
nand U9295 (N_9295,N_3619,N_2248);
xnor U9296 (N_9296,N_4764,N_1447);
and U9297 (N_9297,N_3698,N_2061);
and U9298 (N_9298,N_70,N_3603);
nor U9299 (N_9299,N_4270,N_4556);
and U9300 (N_9300,N_3653,N_1802);
nand U9301 (N_9301,N_4098,N_3374);
or U9302 (N_9302,N_1839,N_1454);
nand U9303 (N_9303,N_4815,N_276);
nand U9304 (N_9304,N_361,N_4918);
nor U9305 (N_9305,N_3646,N_1526);
nand U9306 (N_9306,N_1071,N_2941);
nor U9307 (N_9307,N_1329,N_2345);
nor U9308 (N_9308,N_3743,N_4654);
and U9309 (N_9309,N_1651,N_4425);
nand U9310 (N_9310,N_3464,N_4963);
or U9311 (N_9311,N_604,N_433);
xor U9312 (N_9312,N_290,N_1647);
nor U9313 (N_9313,N_3710,N_3596);
or U9314 (N_9314,N_1186,N_4910);
xor U9315 (N_9315,N_4712,N_4658);
xor U9316 (N_9316,N_3290,N_1367);
nand U9317 (N_9317,N_4216,N_675);
nand U9318 (N_9318,N_3464,N_2233);
or U9319 (N_9319,N_1276,N_3145);
xnor U9320 (N_9320,N_1313,N_3748);
and U9321 (N_9321,N_303,N_840);
or U9322 (N_9322,N_1614,N_2544);
nor U9323 (N_9323,N_1490,N_2730);
and U9324 (N_9324,N_2682,N_2106);
nand U9325 (N_9325,N_3199,N_4888);
and U9326 (N_9326,N_4741,N_3512);
xnor U9327 (N_9327,N_4043,N_4568);
xor U9328 (N_9328,N_3062,N_1156);
nand U9329 (N_9329,N_2409,N_2344);
or U9330 (N_9330,N_2792,N_3491);
or U9331 (N_9331,N_2193,N_4512);
nor U9332 (N_9332,N_4736,N_684);
nand U9333 (N_9333,N_4980,N_199);
xnor U9334 (N_9334,N_3021,N_2410);
xor U9335 (N_9335,N_3416,N_915);
or U9336 (N_9336,N_1891,N_4435);
nor U9337 (N_9337,N_4796,N_1560);
nor U9338 (N_9338,N_4572,N_870);
xnor U9339 (N_9339,N_3839,N_4496);
or U9340 (N_9340,N_4395,N_484);
nand U9341 (N_9341,N_4129,N_2534);
or U9342 (N_9342,N_3636,N_3905);
nor U9343 (N_9343,N_4182,N_1908);
nor U9344 (N_9344,N_889,N_2022);
xnor U9345 (N_9345,N_2030,N_3956);
and U9346 (N_9346,N_1790,N_4125);
and U9347 (N_9347,N_67,N_4306);
nor U9348 (N_9348,N_4123,N_1300);
xor U9349 (N_9349,N_1912,N_403);
and U9350 (N_9350,N_1930,N_4391);
nor U9351 (N_9351,N_1180,N_3306);
xor U9352 (N_9352,N_1433,N_2698);
or U9353 (N_9353,N_3092,N_4610);
xor U9354 (N_9354,N_4073,N_2179);
nor U9355 (N_9355,N_4566,N_1810);
or U9356 (N_9356,N_4433,N_3658);
nand U9357 (N_9357,N_1116,N_1531);
and U9358 (N_9358,N_3184,N_1278);
xnor U9359 (N_9359,N_198,N_2729);
nand U9360 (N_9360,N_2867,N_1481);
and U9361 (N_9361,N_4713,N_1630);
or U9362 (N_9362,N_1670,N_1256);
and U9363 (N_9363,N_3713,N_1626);
xor U9364 (N_9364,N_2592,N_1461);
nand U9365 (N_9365,N_1073,N_3973);
or U9366 (N_9366,N_353,N_4942);
nor U9367 (N_9367,N_4050,N_2867);
and U9368 (N_9368,N_527,N_4376);
nor U9369 (N_9369,N_1846,N_1708);
and U9370 (N_9370,N_2321,N_125);
nor U9371 (N_9371,N_2895,N_2357);
nor U9372 (N_9372,N_1285,N_2785);
and U9373 (N_9373,N_3906,N_3245);
nor U9374 (N_9374,N_1370,N_2137);
nand U9375 (N_9375,N_3755,N_695);
or U9376 (N_9376,N_1899,N_1497);
nand U9377 (N_9377,N_1243,N_3653);
or U9378 (N_9378,N_4786,N_304);
nor U9379 (N_9379,N_513,N_647);
nand U9380 (N_9380,N_4823,N_4385);
and U9381 (N_9381,N_3199,N_4439);
nor U9382 (N_9382,N_4045,N_2173);
or U9383 (N_9383,N_436,N_3942);
xor U9384 (N_9384,N_2009,N_1393);
nand U9385 (N_9385,N_81,N_1721);
nor U9386 (N_9386,N_2167,N_3244);
nand U9387 (N_9387,N_3706,N_3135);
or U9388 (N_9388,N_4318,N_3461);
nor U9389 (N_9389,N_146,N_3218);
or U9390 (N_9390,N_380,N_1790);
or U9391 (N_9391,N_3394,N_3898);
and U9392 (N_9392,N_3826,N_4956);
nand U9393 (N_9393,N_144,N_3912);
nand U9394 (N_9394,N_129,N_900);
nand U9395 (N_9395,N_2296,N_1665);
xnor U9396 (N_9396,N_864,N_3679);
nand U9397 (N_9397,N_3284,N_1163);
nor U9398 (N_9398,N_466,N_144);
xnor U9399 (N_9399,N_4474,N_1639);
and U9400 (N_9400,N_2933,N_158);
or U9401 (N_9401,N_614,N_2937);
nor U9402 (N_9402,N_1900,N_2883);
or U9403 (N_9403,N_3699,N_2995);
nand U9404 (N_9404,N_1755,N_3306);
xor U9405 (N_9405,N_1568,N_1239);
nor U9406 (N_9406,N_2285,N_18);
nand U9407 (N_9407,N_4644,N_506);
and U9408 (N_9408,N_3260,N_4296);
and U9409 (N_9409,N_4084,N_868);
and U9410 (N_9410,N_417,N_3018);
nand U9411 (N_9411,N_2898,N_4548);
or U9412 (N_9412,N_4398,N_1863);
or U9413 (N_9413,N_4883,N_762);
or U9414 (N_9414,N_2443,N_4200);
nand U9415 (N_9415,N_1263,N_4924);
xor U9416 (N_9416,N_2772,N_845);
and U9417 (N_9417,N_3067,N_1796);
and U9418 (N_9418,N_4119,N_204);
nor U9419 (N_9419,N_111,N_293);
and U9420 (N_9420,N_2100,N_3651);
and U9421 (N_9421,N_902,N_2705);
and U9422 (N_9422,N_3906,N_3808);
nor U9423 (N_9423,N_3259,N_2489);
xor U9424 (N_9424,N_703,N_955);
nor U9425 (N_9425,N_31,N_4642);
or U9426 (N_9426,N_2394,N_4862);
nor U9427 (N_9427,N_1133,N_1669);
nor U9428 (N_9428,N_2082,N_4103);
or U9429 (N_9429,N_25,N_410);
nor U9430 (N_9430,N_1352,N_3022);
or U9431 (N_9431,N_2905,N_1033);
nand U9432 (N_9432,N_4272,N_1571);
and U9433 (N_9433,N_1798,N_1548);
nor U9434 (N_9434,N_4820,N_2230);
nor U9435 (N_9435,N_1815,N_446);
nor U9436 (N_9436,N_1351,N_548);
nor U9437 (N_9437,N_1366,N_1299);
xnor U9438 (N_9438,N_2385,N_2893);
nand U9439 (N_9439,N_788,N_1833);
and U9440 (N_9440,N_2298,N_1145);
and U9441 (N_9441,N_4556,N_1233);
and U9442 (N_9442,N_2584,N_933);
and U9443 (N_9443,N_4268,N_3970);
nor U9444 (N_9444,N_2407,N_4892);
nor U9445 (N_9445,N_1489,N_2054);
nand U9446 (N_9446,N_1832,N_4766);
and U9447 (N_9447,N_306,N_158);
and U9448 (N_9448,N_241,N_1867);
and U9449 (N_9449,N_2199,N_4800);
and U9450 (N_9450,N_4934,N_353);
and U9451 (N_9451,N_3376,N_4080);
nor U9452 (N_9452,N_4539,N_3617);
nor U9453 (N_9453,N_2475,N_4015);
or U9454 (N_9454,N_253,N_4492);
or U9455 (N_9455,N_4040,N_383);
nor U9456 (N_9456,N_2637,N_2355);
or U9457 (N_9457,N_1490,N_226);
xor U9458 (N_9458,N_4937,N_506);
nand U9459 (N_9459,N_1074,N_2187);
and U9460 (N_9460,N_4463,N_1231);
and U9461 (N_9461,N_1980,N_4623);
nand U9462 (N_9462,N_4207,N_713);
nand U9463 (N_9463,N_4717,N_1174);
or U9464 (N_9464,N_4718,N_3174);
or U9465 (N_9465,N_1748,N_2029);
xor U9466 (N_9466,N_4525,N_2589);
or U9467 (N_9467,N_4463,N_567);
nor U9468 (N_9468,N_2633,N_4922);
or U9469 (N_9469,N_1119,N_1285);
nor U9470 (N_9470,N_1090,N_10);
or U9471 (N_9471,N_429,N_4193);
and U9472 (N_9472,N_3985,N_3368);
and U9473 (N_9473,N_3255,N_226);
nor U9474 (N_9474,N_969,N_182);
nand U9475 (N_9475,N_1405,N_1240);
xnor U9476 (N_9476,N_3480,N_3652);
xor U9477 (N_9477,N_1811,N_2957);
and U9478 (N_9478,N_1975,N_1850);
nor U9479 (N_9479,N_4685,N_1449);
nand U9480 (N_9480,N_2749,N_4631);
or U9481 (N_9481,N_956,N_1718);
or U9482 (N_9482,N_533,N_2877);
nand U9483 (N_9483,N_3414,N_2806);
and U9484 (N_9484,N_2660,N_1355);
nor U9485 (N_9485,N_1983,N_2802);
nand U9486 (N_9486,N_3028,N_2666);
nor U9487 (N_9487,N_4837,N_1870);
or U9488 (N_9488,N_1330,N_2619);
xnor U9489 (N_9489,N_194,N_1048);
or U9490 (N_9490,N_1713,N_4690);
or U9491 (N_9491,N_4671,N_226);
and U9492 (N_9492,N_1195,N_521);
and U9493 (N_9493,N_3434,N_2087);
or U9494 (N_9494,N_1104,N_3962);
and U9495 (N_9495,N_4644,N_1983);
nor U9496 (N_9496,N_611,N_1031);
or U9497 (N_9497,N_4693,N_1677);
nor U9498 (N_9498,N_2005,N_3646);
or U9499 (N_9499,N_3683,N_841);
or U9500 (N_9500,N_2151,N_3206);
nand U9501 (N_9501,N_1559,N_1584);
nor U9502 (N_9502,N_4943,N_1854);
nand U9503 (N_9503,N_53,N_1616);
nand U9504 (N_9504,N_3551,N_31);
xor U9505 (N_9505,N_1897,N_24);
and U9506 (N_9506,N_4177,N_1992);
nor U9507 (N_9507,N_4564,N_4369);
or U9508 (N_9508,N_1289,N_3787);
and U9509 (N_9509,N_4035,N_4971);
nor U9510 (N_9510,N_4422,N_1091);
and U9511 (N_9511,N_1908,N_673);
xor U9512 (N_9512,N_1863,N_2878);
or U9513 (N_9513,N_1789,N_2440);
and U9514 (N_9514,N_3238,N_4710);
and U9515 (N_9515,N_4675,N_3716);
or U9516 (N_9516,N_642,N_4070);
and U9517 (N_9517,N_4542,N_1107);
or U9518 (N_9518,N_1705,N_2737);
xnor U9519 (N_9519,N_1785,N_1224);
xnor U9520 (N_9520,N_1753,N_2077);
nor U9521 (N_9521,N_3396,N_394);
or U9522 (N_9522,N_2347,N_2658);
or U9523 (N_9523,N_3079,N_2671);
and U9524 (N_9524,N_1559,N_983);
or U9525 (N_9525,N_2272,N_3744);
nor U9526 (N_9526,N_3714,N_3890);
nor U9527 (N_9527,N_4879,N_637);
nor U9528 (N_9528,N_1655,N_1956);
nand U9529 (N_9529,N_3001,N_2968);
xnor U9530 (N_9530,N_4844,N_3577);
nand U9531 (N_9531,N_1526,N_107);
nor U9532 (N_9532,N_900,N_3707);
nand U9533 (N_9533,N_932,N_169);
xor U9534 (N_9534,N_1998,N_2108);
and U9535 (N_9535,N_4819,N_3043);
and U9536 (N_9536,N_4535,N_3863);
nor U9537 (N_9537,N_1071,N_1305);
xor U9538 (N_9538,N_4814,N_4018);
and U9539 (N_9539,N_3651,N_17);
and U9540 (N_9540,N_2965,N_2417);
and U9541 (N_9541,N_2714,N_4032);
nor U9542 (N_9542,N_1547,N_4166);
xor U9543 (N_9543,N_49,N_864);
or U9544 (N_9544,N_4234,N_22);
nor U9545 (N_9545,N_791,N_998);
nor U9546 (N_9546,N_2776,N_1203);
and U9547 (N_9547,N_1279,N_3769);
nor U9548 (N_9548,N_3256,N_2885);
or U9549 (N_9549,N_2454,N_2460);
nand U9550 (N_9550,N_3135,N_1529);
nor U9551 (N_9551,N_2416,N_3819);
and U9552 (N_9552,N_671,N_2244);
xnor U9553 (N_9553,N_4769,N_3799);
xnor U9554 (N_9554,N_3055,N_4554);
nor U9555 (N_9555,N_1798,N_4569);
and U9556 (N_9556,N_2680,N_3414);
xnor U9557 (N_9557,N_3153,N_3616);
or U9558 (N_9558,N_4401,N_4074);
nand U9559 (N_9559,N_3561,N_4105);
nor U9560 (N_9560,N_335,N_2199);
and U9561 (N_9561,N_3835,N_2109);
and U9562 (N_9562,N_4708,N_2846);
and U9563 (N_9563,N_2312,N_2844);
nand U9564 (N_9564,N_4656,N_1113);
nand U9565 (N_9565,N_937,N_2231);
and U9566 (N_9566,N_2140,N_979);
and U9567 (N_9567,N_4099,N_3678);
and U9568 (N_9568,N_2260,N_4461);
nor U9569 (N_9569,N_2672,N_607);
and U9570 (N_9570,N_384,N_497);
or U9571 (N_9571,N_2269,N_3827);
nor U9572 (N_9572,N_3607,N_47);
or U9573 (N_9573,N_367,N_2416);
or U9574 (N_9574,N_1600,N_3772);
and U9575 (N_9575,N_1014,N_341);
nand U9576 (N_9576,N_749,N_280);
xor U9577 (N_9577,N_4963,N_4707);
xnor U9578 (N_9578,N_1269,N_2263);
and U9579 (N_9579,N_982,N_2352);
or U9580 (N_9580,N_937,N_2299);
and U9581 (N_9581,N_1363,N_2205);
and U9582 (N_9582,N_791,N_438);
and U9583 (N_9583,N_1373,N_1599);
and U9584 (N_9584,N_3946,N_3042);
and U9585 (N_9585,N_1062,N_4085);
nor U9586 (N_9586,N_4721,N_4145);
or U9587 (N_9587,N_4232,N_4727);
or U9588 (N_9588,N_489,N_4521);
or U9589 (N_9589,N_2025,N_3470);
and U9590 (N_9590,N_15,N_1632);
xnor U9591 (N_9591,N_3455,N_1556);
and U9592 (N_9592,N_3465,N_4039);
nor U9593 (N_9593,N_1819,N_4325);
or U9594 (N_9594,N_2378,N_1439);
or U9595 (N_9595,N_4104,N_2556);
or U9596 (N_9596,N_2930,N_4428);
and U9597 (N_9597,N_2886,N_1860);
and U9598 (N_9598,N_2243,N_171);
nor U9599 (N_9599,N_2588,N_3608);
or U9600 (N_9600,N_1748,N_3271);
or U9601 (N_9601,N_144,N_867);
or U9602 (N_9602,N_3622,N_4283);
nor U9603 (N_9603,N_1240,N_4568);
xor U9604 (N_9604,N_2139,N_4171);
nand U9605 (N_9605,N_866,N_3971);
nand U9606 (N_9606,N_1805,N_1576);
xnor U9607 (N_9607,N_2530,N_2751);
xnor U9608 (N_9608,N_3092,N_4211);
nor U9609 (N_9609,N_445,N_1860);
nand U9610 (N_9610,N_2000,N_2416);
nand U9611 (N_9611,N_4359,N_436);
nand U9612 (N_9612,N_4842,N_2287);
xnor U9613 (N_9613,N_4068,N_1262);
or U9614 (N_9614,N_1077,N_2611);
and U9615 (N_9615,N_423,N_415);
nand U9616 (N_9616,N_1961,N_880);
and U9617 (N_9617,N_1528,N_320);
nand U9618 (N_9618,N_1453,N_1890);
xnor U9619 (N_9619,N_542,N_1040);
xor U9620 (N_9620,N_568,N_2157);
or U9621 (N_9621,N_3871,N_1472);
nor U9622 (N_9622,N_4750,N_1639);
and U9623 (N_9623,N_3549,N_1595);
and U9624 (N_9624,N_3625,N_3654);
and U9625 (N_9625,N_1011,N_3732);
and U9626 (N_9626,N_1139,N_2656);
and U9627 (N_9627,N_2851,N_3345);
xor U9628 (N_9628,N_2115,N_4114);
and U9629 (N_9629,N_2374,N_1005);
and U9630 (N_9630,N_2459,N_3921);
nor U9631 (N_9631,N_930,N_1591);
nand U9632 (N_9632,N_812,N_1390);
and U9633 (N_9633,N_4472,N_3381);
and U9634 (N_9634,N_1757,N_1507);
nor U9635 (N_9635,N_2611,N_2908);
xor U9636 (N_9636,N_958,N_3816);
nor U9637 (N_9637,N_752,N_4411);
xnor U9638 (N_9638,N_3164,N_3601);
or U9639 (N_9639,N_1732,N_1943);
nor U9640 (N_9640,N_1962,N_3433);
xor U9641 (N_9641,N_885,N_4778);
or U9642 (N_9642,N_2402,N_2542);
or U9643 (N_9643,N_2743,N_3016);
and U9644 (N_9644,N_1441,N_3209);
xor U9645 (N_9645,N_4196,N_3164);
nor U9646 (N_9646,N_3415,N_4137);
and U9647 (N_9647,N_2981,N_2697);
nor U9648 (N_9648,N_4093,N_2633);
and U9649 (N_9649,N_3528,N_424);
and U9650 (N_9650,N_40,N_1372);
xor U9651 (N_9651,N_1014,N_2976);
and U9652 (N_9652,N_4208,N_3114);
or U9653 (N_9653,N_1345,N_3115);
xnor U9654 (N_9654,N_1373,N_2950);
nor U9655 (N_9655,N_4973,N_1753);
xor U9656 (N_9656,N_3068,N_55);
and U9657 (N_9657,N_4682,N_1867);
nand U9658 (N_9658,N_4925,N_722);
and U9659 (N_9659,N_4899,N_4343);
or U9660 (N_9660,N_4535,N_4585);
or U9661 (N_9661,N_4511,N_3687);
nand U9662 (N_9662,N_2295,N_4308);
nor U9663 (N_9663,N_1908,N_4023);
nand U9664 (N_9664,N_385,N_3082);
and U9665 (N_9665,N_4701,N_4767);
or U9666 (N_9666,N_1443,N_1106);
nor U9667 (N_9667,N_3792,N_715);
nand U9668 (N_9668,N_3900,N_4906);
nand U9669 (N_9669,N_4211,N_848);
nor U9670 (N_9670,N_2876,N_926);
nor U9671 (N_9671,N_2929,N_1349);
xnor U9672 (N_9672,N_2207,N_3400);
nor U9673 (N_9673,N_195,N_3632);
and U9674 (N_9674,N_826,N_4412);
nand U9675 (N_9675,N_706,N_4215);
xor U9676 (N_9676,N_3522,N_1492);
or U9677 (N_9677,N_2634,N_2671);
nand U9678 (N_9678,N_2143,N_2822);
nor U9679 (N_9679,N_4004,N_1611);
nor U9680 (N_9680,N_3972,N_3758);
or U9681 (N_9681,N_2731,N_2738);
xor U9682 (N_9682,N_831,N_998);
or U9683 (N_9683,N_3330,N_1349);
nand U9684 (N_9684,N_2780,N_4145);
nand U9685 (N_9685,N_1508,N_3777);
xnor U9686 (N_9686,N_1011,N_1816);
and U9687 (N_9687,N_3105,N_2698);
or U9688 (N_9688,N_4498,N_402);
nor U9689 (N_9689,N_3257,N_4887);
xor U9690 (N_9690,N_4631,N_2913);
nand U9691 (N_9691,N_775,N_2530);
nor U9692 (N_9692,N_2059,N_2100);
nand U9693 (N_9693,N_2429,N_2844);
and U9694 (N_9694,N_1414,N_4726);
or U9695 (N_9695,N_98,N_1069);
nand U9696 (N_9696,N_1867,N_3663);
and U9697 (N_9697,N_3591,N_3744);
and U9698 (N_9698,N_2345,N_486);
nor U9699 (N_9699,N_4406,N_1851);
nand U9700 (N_9700,N_3416,N_1493);
nor U9701 (N_9701,N_3518,N_1883);
nor U9702 (N_9702,N_2651,N_4702);
and U9703 (N_9703,N_4268,N_2933);
and U9704 (N_9704,N_1612,N_2884);
nand U9705 (N_9705,N_3351,N_1988);
or U9706 (N_9706,N_2081,N_371);
xor U9707 (N_9707,N_1807,N_1053);
nor U9708 (N_9708,N_4591,N_1133);
nor U9709 (N_9709,N_1799,N_4069);
nand U9710 (N_9710,N_454,N_1642);
and U9711 (N_9711,N_3037,N_3957);
or U9712 (N_9712,N_559,N_4405);
nand U9713 (N_9713,N_185,N_335);
nand U9714 (N_9714,N_3036,N_4494);
or U9715 (N_9715,N_4218,N_2217);
or U9716 (N_9716,N_2882,N_205);
or U9717 (N_9717,N_330,N_2672);
nand U9718 (N_9718,N_2065,N_59);
nand U9719 (N_9719,N_1975,N_4121);
nand U9720 (N_9720,N_3938,N_2988);
nor U9721 (N_9721,N_3692,N_844);
xor U9722 (N_9722,N_865,N_1632);
nor U9723 (N_9723,N_1390,N_513);
xor U9724 (N_9724,N_2384,N_166);
and U9725 (N_9725,N_4834,N_431);
and U9726 (N_9726,N_1412,N_145);
nor U9727 (N_9727,N_247,N_2665);
nor U9728 (N_9728,N_1055,N_4065);
xnor U9729 (N_9729,N_3592,N_4309);
and U9730 (N_9730,N_4427,N_3575);
or U9731 (N_9731,N_1857,N_4982);
and U9732 (N_9732,N_4915,N_4024);
and U9733 (N_9733,N_1779,N_1299);
and U9734 (N_9734,N_4261,N_619);
and U9735 (N_9735,N_1089,N_4733);
nand U9736 (N_9736,N_2548,N_1770);
nand U9737 (N_9737,N_2668,N_2987);
and U9738 (N_9738,N_4255,N_1241);
or U9739 (N_9739,N_4957,N_3354);
nor U9740 (N_9740,N_4462,N_4517);
and U9741 (N_9741,N_356,N_1303);
nand U9742 (N_9742,N_3631,N_3840);
or U9743 (N_9743,N_3944,N_4797);
nor U9744 (N_9744,N_716,N_1573);
nor U9745 (N_9745,N_4777,N_1066);
and U9746 (N_9746,N_1023,N_1421);
nand U9747 (N_9747,N_3473,N_3634);
nand U9748 (N_9748,N_2483,N_2667);
nand U9749 (N_9749,N_4850,N_1111);
and U9750 (N_9750,N_4415,N_4878);
and U9751 (N_9751,N_620,N_3113);
nor U9752 (N_9752,N_129,N_2972);
nand U9753 (N_9753,N_4269,N_4118);
and U9754 (N_9754,N_1562,N_3577);
nor U9755 (N_9755,N_3824,N_1990);
xor U9756 (N_9756,N_1047,N_2629);
or U9757 (N_9757,N_3931,N_2206);
nand U9758 (N_9758,N_2963,N_2164);
nand U9759 (N_9759,N_4550,N_2541);
nor U9760 (N_9760,N_2655,N_7);
and U9761 (N_9761,N_2690,N_1161);
nand U9762 (N_9762,N_4789,N_2444);
nand U9763 (N_9763,N_4759,N_3267);
nand U9764 (N_9764,N_95,N_4613);
xnor U9765 (N_9765,N_257,N_3586);
xnor U9766 (N_9766,N_101,N_1692);
nand U9767 (N_9767,N_4461,N_1993);
or U9768 (N_9768,N_4090,N_1731);
or U9769 (N_9769,N_343,N_2879);
and U9770 (N_9770,N_2457,N_2701);
nor U9771 (N_9771,N_2485,N_3286);
nand U9772 (N_9772,N_125,N_973);
and U9773 (N_9773,N_3657,N_2987);
or U9774 (N_9774,N_1485,N_1587);
nor U9775 (N_9775,N_4184,N_2196);
nand U9776 (N_9776,N_53,N_1841);
xor U9777 (N_9777,N_796,N_2580);
nand U9778 (N_9778,N_49,N_4792);
and U9779 (N_9779,N_133,N_4528);
xor U9780 (N_9780,N_3882,N_968);
nand U9781 (N_9781,N_770,N_2419);
xor U9782 (N_9782,N_955,N_1903);
xnor U9783 (N_9783,N_3367,N_157);
or U9784 (N_9784,N_1200,N_74);
nand U9785 (N_9785,N_586,N_2814);
xor U9786 (N_9786,N_2111,N_3090);
or U9787 (N_9787,N_45,N_2015);
and U9788 (N_9788,N_1476,N_4266);
nand U9789 (N_9789,N_4675,N_1905);
xnor U9790 (N_9790,N_4920,N_3742);
nand U9791 (N_9791,N_699,N_2921);
or U9792 (N_9792,N_1751,N_1129);
nand U9793 (N_9793,N_151,N_4245);
nor U9794 (N_9794,N_4167,N_1858);
nor U9795 (N_9795,N_563,N_4625);
and U9796 (N_9796,N_3888,N_1878);
nand U9797 (N_9797,N_1962,N_4143);
nor U9798 (N_9798,N_520,N_1497);
xnor U9799 (N_9799,N_4700,N_755);
or U9800 (N_9800,N_1428,N_2735);
or U9801 (N_9801,N_1943,N_376);
and U9802 (N_9802,N_2820,N_2587);
xnor U9803 (N_9803,N_2790,N_554);
xor U9804 (N_9804,N_2928,N_1882);
nand U9805 (N_9805,N_4855,N_2943);
xnor U9806 (N_9806,N_904,N_1203);
or U9807 (N_9807,N_1385,N_1410);
nor U9808 (N_9808,N_3014,N_4);
nand U9809 (N_9809,N_4317,N_1197);
xor U9810 (N_9810,N_1577,N_1940);
nand U9811 (N_9811,N_1276,N_2936);
or U9812 (N_9812,N_7,N_2759);
nor U9813 (N_9813,N_845,N_3569);
or U9814 (N_9814,N_173,N_3290);
and U9815 (N_9815,N_584,N_3733);
or U9816 (N_9816,N_1717,N_2125);
nor U9817 (N_9817,N_4523,N_3629);
and U9818 (N_9818,N_25,N_4939);
nand U9819 (N_9819,N_2805,N_924);
nor U9820 (N_9820,N_4092,N_3880);
xor U9821 (N_9821,N_1106,N_2621);
nand U9822 (N_9822,N_4306,N_2905);
nand U9823 (N_9823,N_2126,N_4657);
and U9824 (N_9824,N_2419,N_2934);
nand U9825 (N_9825,N_2541,N_1331);
xnor U9826 (N_9826,N_4016,N_3153);
or U9827 (N_9827,N_1509,N_4300);
or U9828 (N_9828,N_2781,N_3927);
nor U9829 (N_9829,N_4001,N_4403);
or U9830 (N_9830,N_2747,N_3450);
nand U9831 (N_9831,N_1809,N_4789);
nand U9832 (N_9832,N_606,N_618);
or U9833 (N_9833,N_2742,N_4217);
or U9834 (N_9834,N_1150,N_1664);
or U9835 (N_9835,N_3988,N_4780);
nor U9836 (N_9836,N_3910,N_2486);
or U9837 (N_9837,N_4228,N_742);
nand U9838 (N_9838,N_2631,N_4284);
nor U9839 (N_9839,N_1859,N_1658);
or U9840 (N_9840,N_1680,N_1694);
and U9841 (N_9841,N_4705,N_1237);
or U9842 (N_9842,N_941,N_3157);
xnor U9843 (N_9843,N_2976,N_2801);
and U9844 (N_9844,N_355,N_3859);
xor U9845 (N_9845,N_4756,N_2074);
nand U9846 (N_9846,N_1669,N_89);
and U9847 (N_9847,N_3874,N_3551);
nor U9848 (N_9848,N_1429,N_4594);
and U9849 (N_9849,N_4621,N_2241);
xnor U9850 (N_9850,N_4392,N_3081);
or U9851 (N_9851,N_691,N_1165);
or U9852 (N_9852,N_3990,N_2775);
and U9853 (N_9853,N_3558,N_2220);
xor U9854 (N_9854,N_2909,N_3559);
or U9855 (N_9855,N_4393,N_4313);
and U9856 (N_9856,N_4542,N_1185);
and U9857 (N_9857,N_4274,N_3335);
and U9858 (N_9858,N_892,N_1324);
and U9859 (N_9859,N_2845,N_1785);
xor U9860 (N_9860,N_4391,N_1091);
or U9861 (N_9861,N_395,N_625);
xor U9862 (N_9862,N_4484,N_3428);
nand U9863 (N_9863,N_4444,N_4828);
and U9864 (N_9864,N_2062,N_4135);
and U9865 (N_9865,N_3502,N_4382);
nor U9866 (N_9866,N_2651,N_970);
and U9867 (N_9867,N_1186,N_2740);
and U9868 (N_9868,N_4403,N_4828);
and U9869 (N_9869,N_695,N_3768);
nand U9870 (N_9870,N_4054,N_4736);
xnor U9871 (N_9871,N_3173,N_3160);
or U9872 (N_9872,N_3769,N_2862);
nand U9873 (N_9873,N_1114,N_3174);
and U9874 (N_9874,N_3658,N_1114);
and U9875 (N_9875,N_2259,N_4303);
nand U9876 (N_9876,N_2879,N_4495);
xor U9877 (N_9877,N_4196,N_2501);
nand U9878 (N_9878,N_657,N_1158);
and U9879 (N_9879,N_4739,N_4357);
and U9880 (N_9880,N_4907,N_3130);
nand U9881 (N_9881,N_171,N_2877);
and U9882 (N_9882,N_594,N_1035);
nand U9883 (N_9883,N_598,N_4374);
nand U9884 (N_9884,N_1075,N_4525);
and U9885 (N_9885,N_1917,N_3031);
nand U9886 (N_9886,N_1965,N_4654);
xor U9887 (N_9887,N_4591,N_2039);
or U9888 (N_9888,N_1265,N_59);
xnor U9889 (N_9889,N_1112,N_3774);
xnor U9890 (N_9890,N_1721,N_4444);
nand U9891 (N_9891,N_673,N_3197);
and U9892 (N_9892,N_2039,N_4673);
nand U9893 (N_9893,N_1451,N_3728);
or U9894 (N_9894,N_3519,N_1027);
nor U9895 (N_9895,N_374,N_603);
nor U9896 (N_9896,N_1506,N_2305);
nor U9897 (N_9897,N_2312,N_3301);
nor U9898 (N_9898,N_964,N_232);
nor U9899 (N_9899,N_3059,N_3501);
nand U9900 (N_9900,N_4239,N_1993);
xor U9901 (N_9901,N_1111,N_3075);
or U9902 (N_9902,N_1895,N_4909);
nand U9903 (N_9903,N_356,N_4295);
and U9904 (N_9904,N_1111,N_1443);
xnor U9905 (N_9905,N_2029,N_4291);
nor U9906 (N_9906,N_3867,N_4775);
or U9907 (N_9907,N_166,N_182);
nand U9908 (N_9908,N_221,N_3687);
and U9909 (N_9909,N_3447,N_531);
or U9910 (N_9910,N_4320,N_284);
nand U9911 (N_9911,N_1937,N_1756);
nand U9912 (N_9912,N_225,N_2246);
nor U9913 (N_9913,N_3500,N_4586);
and U9914 (N_9914,N_1234,N_889);
or U9915 (N_9915,N_4275,N_1546);
nand U9916 (N_9916,N_2361,N_718);
nand U9917 (N_9917,N_267,N_2507);
xor U9918 (N_9918,N_4984,N_944);
and U9919 (N_9919,N_3924,N_2039);
nor U9920 (N_9920,N_3825,N_3913);
and U9921 (N_9921,N_1764,N_4260);
or U9922 (N_9922,N_2881,N_2905);
nor U9923 (N_9923,N_3033,N_1434);
xnor U9924 (N_9924,N_2573,N_2321);
xnor U9925 (N_9925,N_559,N_2392);
nand U9926 (N_9926,N_236,N_476);
and U9927 (N_9927,N_218,N_668);
xnor U9928 (N_9928,N_2104,N_2912);
and U9929 (N_9929,N_782,N_2675);
and U9930 (N_9930,N_3316,N_3609);
nand U9931 (N_9931,N_813,N_1974);
xnor U9932 (N_9932,N_4209,N_1783);
xnor U9933 (N_9933,N_54,N_2492);
nand U9934 (N_9934,N_3865,N_2876);
xnor U9935 (N_9935,N_1583,N_1403);
nor U9936 (N_9936,N_4710,N_4611);
and U9937 (N_9937,N_2252,N_843);
and U9938 (N_9938,N_237,N_2439);
nand U9939 (N_9939,N_293,N_1006);
xor U9940 (N_9940,N_1578,N_4684);
nand U9941 (N_9941,N_3899,N_1597);
or U9942 (N_9942,N_1173,N_3356);
nand U9943 (N_9943,N_3072,N_3465);
nand U9944 (N_9944,N_1427,N_59);
and U9945 (N_9945,N_1060,N_65);
xnor U9946 (N_9946,N_1748,N_3512);
or U9947 (N_9947,N_3856,N_2783);
and U9948 (N_9948,N_4750,N_2107);
and U9949 (N_9949,N_4861,N_2149);
and U9950 (N_9950,N_1752,N_1985);
or U9951 (N_9951,N_1946,N_301);
xnor U9952 (N_9952,N_2954,N_1898);
or U9953 (N_9953,N_3745,N_1613);
xor U9954 (N_9954,N_3067,N_1872);
and U9955 (N_9955,N_1242,N_1930);
xor U9956 (N_9956,N_4939,N_3059);
nor U9957 (N_9957,N_58,N_3314);
xnor U9958 (N_9958,N_4484,N_4935);
nor U9959 (N_9959,N_179,N_2456);
nor U9960 (N_9960,N_3802,N_16);
or U9961 (N_9961,N_2124,N_4288);
or U9962 (N_9962,N_830,N_2314);
xnor U9963 (N_9963,N_2121,N_4302);
nor U9964 (N_9964,N_3689,N_630);
xor U9965 (N_9965,N_1491,N_1712);
nor U9966 (N_9966,N_2964,N_2746);
nor U9967 (N_9967,N_1484,N_1409);
xor U9968 (N_9968,N_1623,N_1260);
and U9969 (N_9969,N_1749,N_205);
xnor U9970 (N_9970,N_3591,N_286);
nand U9971 (N_9971,N_4861,N_489);
nand U9972 (N_9972,N_3255,N_2900);
nor U9973 (N_9973,N_209,N_1166);
or U9974 (N_9974,N_1198,N_3063);
or U9975 (N_9975,N_2137,N_195);
or U9976 (N_9976,N_3420,N_3060);
or U9977 (N_9977,N_1720,N_15);
xnor U9978 (N_9978,N_2953,N_4474);
xnor U9979 (N_9979,N_523,N_3077);
or U9980 (N_9980,N_3451,N_2003);
nand U9981 (N_9981,N_3192,N_3593);
and U9982 (N_9982,N_2527,N_748);
xor U9983 (N_9983,N_3087,N_4553);
xor U9984 (N_9984,N_850,N_4996);
and U9985 (N_9985,N_3530,N_2840);
and U9986 (N_9986,N_1979,N_2779);
xnor U9987 (N_9987,N_4162,N_2592);
nand U9988 (N_9988,N_2959,N_4466);
nand U9989 (N_9989,N_2624,N_1114);
nor U9990 (N_9990,N_3382,N_926);
or U9991 (N_9991,N_1521,N_3944);
nand U9992 (N_9992,N_4021,N_2861);
xnor U9993 (N_9993,N_1235,N_2054);
xnor U9994 (N_9994,N_928,N_2775);
nand U9995 (N_9995,N_4241,N_2671);
xor U9996 (N_9996,N_2423,N_3258);
nand U9997 (N_9997,N_3070,N_784);
xnor U9998 (N_9998,N_2498,N_1287);
and U9999 (N_9999,N_3316,N_1215);
or U10000 (N_10000,N_5169,N_9780);
nand U10001 (N_10001,N_5813,N_6148);
nand U10002 (N_10002,N_8043,N_5080);
xor U10003 (N_10003,N_5258,N_7403);
xor U10004 (N_10004,N_5760,N_9008);
and U10005 (N_10005,N_6033,N_9803);
nor U10006 (N_10006,N_7881,N_7265);
xor U10007 (N_10007,N_8238,N_6832);
and U10008 (N_10008,N_6494,N_5215);
nand U10009 (N_10009,N_9342,N_7383);
or U10010 (N_10010,N_7351,N_7233);
nand U10011 (N_10011,N_7440,N_8645);
nand U10012 (N_10012,N_7199,N_9997);
or U10013 (N_10013,N_8656,N_7662);
xor U10014 (N_10014,N_8391,N_9636);
or U10015 (N_10015,N_6571,N_8558);
nor U10016 (N_10016,N_6594,N_9648);
and U10017 (N_10017,N_6060,N_5347);
and U10018 (N_10018,N_6253,N_8689);
or U10019 (N_10019,N_5402,N_5333);
nand U10020 (N_10020,N_7218,N_9778);
nand U10021 (N_10021,N_7311,N_9991);
or U10022 (N_10022,N_5996,N_6115);
and U10023 (N_10023,N_9515,N_6091);
nand U10024 (N_10024,N_5667,N_9125);
or U10025 (N_10025,N_5932,N_7807);
nor U10026 (N_10026,N_7045,N_8754);
and U10027 (N_10027,N_5617,N_9822);
nand U10028 (N_10028,N_9158,N_8577);
and U10029 (N_10029,N_9986,N_7399);
xnor U10030 (N_10030,N_6525,N_6291);
or U10031 (N_10031,N_9339,N_5535);
and U10032 (N_10032,N_6848,N_7847);
nor U10033 (N_10033,N_5806,N_5263);
or U10034 (N_10034,N_7945,N_8950);
and U10035 (N_10035,N_7359,N_5807);
or U10036 (N_10036,N_8234,N_9152);
or U10037 (N_10037,N_6849,N_7465);
and U10038 (N_10038,N_5107,N_5013);
nand U10039 (N_10039,N_7164,N_5508);
or U10040 (N_10040,N_9611,N_5057);
nand U10041 (N_10041,N_6282,N_5369);
xor U10042 (N_10042,N_9094,N_5443);
or U10043 (N_10043,N_9206,N_5550);
or U10044 (N_10044,N_5067,N_9500);
xnor U10045 (N_10045,N_8476,N_9977);
nand U10046 (N_10046,N_7350,N_5922);
and U10047 (N_10047,N_6995,N_6551);
nand U10048 (N_10048,N_8197,N_7735);
and U10049 (N_10049,N_6501,N_8755);
nand U10050 (N_10050,N_5558,N_6378);
nor U10051 (N_10051,N_7602,N_5995);
and U10052 (N_10052,N_5834,N_5121);
nor U10053 (N_10053,N_7939,N_5001);
or U10054 (N_10054,N_9316,N_9644);
nand U10055 (N_10055,N_6162,N_8627);
and U10056 (N_10056,N_8169,N_6924);
nor U10057 (N_10057,N_6829,N_7476);
and U10058 (N_10058,N_8768,N_6249);
and U10059 (N_10059,N_7170,N_8437);
xnor U10060 (N_10060,N_8341,N_8021);
or U10061 (N_10061,N_9848,N_8142);
nand U10062 (N_10062,N_7270,N_9556);
nand U10063 (N_10063,N_8521,N_5582);
nand U10064 (N_10064,N_6393,N_9261);
nand U10065 (N_10065,N_7979,N_6289);
nor U10066 (N_10066,N_8194,N_5909);
nor U10067 (N_10067,N_7365,N_7842);
or U10068 (N_10068,N_5038,N_8695);
and U10069 (N_10069,N_7690,N_6283);
and U10070 (N_10070,N_8574,N_9916);
nor U10071 (N_10071,N_9324,N_5661);
and U10072 (N_10072,N_5842,N_5585);
and U10073 (N_10073,N_5052,N_6363);
xnor U10074 (N_10074,N_5050,N_9197);
or U10075 (N_10075,N_7558,N_6508);
and U10076 (N_10076,N_5664,N_5359);
nand U10077 (N_10077,N_8412,N_8785);
xnor U10078 (N_10078,N_6660,N_6417);
nor U10079 (N_10079,N_7419,N_5492);
or U10080 (N_10080,N_6330,N_9940);
or U10081 (N_10081,N_6907,N_8339);
nand U10082 (N_10082,N_8293,N_9038);
and U10083 (N_10083,N_6547,N_8775);
xor U10084 (N_10084,N_7159,N_6220);
and U10085 (N_10085,N_8835,N_8429);
nand U10086 (N_10086,N_5607,N_8196);
xnor U10087 (N_10087,N_8546,N_5532);
or U10088 (N_10088,N_8108,N_8707);
nand U10089 (N_10089,N_5479,N_8924);
nor U10090 (N_10090,N_5660,N_5461);
nor U10091 (N_10091,N_7422,N_6809);
nand U10092 (N_10092,N_8143,N_5594);
xor U10093 (N_10093,N_8333,N_7243);
nand U10094 (N_10094,N_8311,N_7165);
nand U10095 (N_10095,N_8449,N_9494);
nand U10096 (N_10096,N_7434,N_6264);
xor U10097 (N_10097,N_9157,N_9689);
nand U10098 (N_10098,N_7734,N_8374);
nand U10099 (N_10099,N_6197,N_6325);
nand U10100 (N_10100,N_6214,N_8126);
nor U10101 (N_10101,N_7687,N_7982);
nor U10102 (N_10102,N_5068,N_7854);
and U10103 (N_10103,N_6134,N_5151);
nor U10104 (N_10104,N_8564,N_5383);
or U10105 (N_10105,N_7702,N_9815);
and U10106 (N_10106,N_5900,N_8064);
and U10107 (N_10107,N_5757,N_8532);
and U10108 (N_10108,N_6013,N_8618);
nand U10109 (N_10109,N_5738,N_6491);
nor U10110 (N_10110,N_6331,N_7418);
nor U10111 (N_10111,N_7241,N_8235);
nand U10112 (N_10112,N_5280,N_8591);
nand U10113 (N_10113,N_8807,N_5938);
nor U10114 (N_10114,N_6210,N_8895);
xor U10115 (N_10115,N_9132,N_5256);
nand U10116 (N_10116,N_7126,N_6655);
or U10117 (N_10117,N_5033,N_6123);
nor U10118 (N_10118,N_5487,N_5022);
nor U10119 (N_10119,N_8173,N_9052);
xor U10120 (N_10120,N_7193,N_7450);
or U10121 (N_10121,N_7720,N_8359);
nor U10122 (N_10122,N_7041,N_7666);
or U10123 (N_10123,N_5344,N_6954);
nand U10124 (N_10124,N_6304,N_8543);
and U10125 (N_10125,N_7230,N_7801);
nand U10126 (N_10126,N_5414,N_8252);
xnor U10127 (N_10127,N_7040,N_8943);
nand U10128 (N_10128,N_5094,N_9218);
nand U10129 (N_10129,N_5941,N_6349);
or U10130 (N_10130,N_8536,N_8296);
nand U10131 (N_10131,N_6744,N_7300);
nand U10132 (N_10132,N_6636,N_9584);
nand U10133 (N_10133,N_6733,N_6117);
xor U10134 (N_10134,N_6438,N_6640);
and U10135 (N_10135,N_5516,N_9974);
xor U10136 (N_10136,N_8134,N_7083);
nand U10137 (N_10137,N_8081,N_9066);
nand U10138 (N_10138,N_9424,N_9397);
or U10139 (N_10139,N_9200,N_9242);
or U10140 (N_10140,N_6429,N_9585);
xnor U10141 (N_10141,N_5673,N_5000);
nor U10142 (N_10142,N_6534,N_6958);
nor U10143 (N_10143,N_6410,N_5305);
nor U10144 (N_10144,N_9182,N_5166);
and U10145 (N_10145,N_6688,N_9393);
or U10146 (N_10146,N_7220,N_8080);
xor U10147 (N_10147,N_8060,N_9283);
or U10148 (N_10148,N_5631,N_8639);
and U10149 (N_10149,N_9361,N_8007);
or U10150 (N_10150,N_6173,N_9666);
and U10151 (N_10151,N_5522,N_5229);
xnor U10152 (N_10152,N_6896,N_9348);
xnor U10153 (N_10153,N_6423,N_6615);
nor U10154 (N_10154,N_9830,N_5575);
nor U10155 (N_10155,N_9475,N_9349);
nor U10156 (N_10156,N_6816,N_9405);
or U10157 (N_10157,N_5036,N_9659);
xnor U10158 (N_10158,N_8630,N_8839);
xnor U10159 (N_10159,N_8324,N_8770);
xnor U10160 (N_10160,N_7634,N_8127);
xnor U10161 (N_10161,N_8345,N_8482);
and U10162 (N_10162,N_8453,N_6165);
xor U10163 (N_10163,N_7693,N_9151);
or U10164 (N_10164,N_5720,N_8918);
or U10165 (N_10165,N_8692,N_7551);
nor U10166 (N_10166,N_6276,N_5940);
xnor U10167 (N_10167,N_9990,N_5471);
and U10168 (N_10168,N_6481,N_5355);
xnor U10169 (N_10169,N_7183,N_9435);
nand U10170 (N_10170,N_6384,N_7719);
or U10171 (N_10171,N_7084,N_5903);
nand U10172 (N_10172,N_9557,N_7313);
xor U10173 (N_10173,N_9322,N_7330);
xor U10174 (N_10174,N_9669,N_6053);
nand U10175 (N_10175,N_9371,N_8612);
xnor U10176 (N_10176,N_7969,N_5910);
or U10177 (N_10177,N_9967,N_6181);
xor U10178 (N_10178,N_9310,N_6087);
nand U10179 (N_10179,N_7884,N_5948);
xnor U10180 (N_10180,N_7466,N_6887);
nor U10181 (N_10181,N_7988,N_6564);
xnor U10182 (N_10182,N_5275,N_9612);
nor U10183 (N_10183,N_5827,N_8268);
nor U10184 (N_10184,N_6350,N_8939);
xnor U10185 (N_10185,N_7845,N_9297);
nor U10186 (N_10186,N_8610,N_9837);
or U10187 (N_10187,N_8363,N_5570);
and U10188 (N_10188,N_5884,N_9290);
and U10189 (N_10189,N_5482,N_5978);
and U10190 (N_10190,N_8410,N_5872);
xor U10191 (N_10191,N_5271,N_9482);
xor U10192 (N_10192,N_6372,N_8382);
or U10193 (N_10193,N_7732,N_8983);
xor U10194 (N_10194,N_7175,N_7508);
or U10195 (N_10195,N_7714,N_9089);
xnor U10196 (N_10196,N_5307,N_8748);
or U10197 (N_10197,N_6301,N_9683);
nand U10198 (N_10198,N_6175,N_8207);
or U10199 (N_10199,N_6799,N_9904);
and U10200 (N_10200,N_7948,N_7586);
xnor U10201 (N_10201,N_7857,N_5919);
nand U10202 (N_10202,N_6105,N_5826);
or U10203 (N_10203,N_6323,N_9718);
or U10204 (N_10204,N_9819,N_6144);
nor U10205 (N_10205,N_7708,N_8479);
nand U10206 (N_10206,N_7116,N_6647);
and U10207 (N_10207,N_5225,N_7420);
or U10208 (N_10208,N_5889,N_5090);
xor U10209 (N_10209,N_9220,N_5597);
xnor U10210 (N_10210,N_6020,N_6486);
xor U10211 (N_10211,N_9399,N_7906);
or U10212 (N_10212,N_6824,N_5767);
nor U10213 (N_10213,N_9672,N_7893);
xnor U10214 (N_10214,N_5066,N_5843);
and U10215 (N_10215,N_5200,N_5973);
nor U10216 (N_10216,N_7179,N_5891);
or U10217 (N_10217,N_6965,N_5386);
or U10218 (N_10218,N_9193,N_8248);
xor U10219 (N_10219,N_5274,N_9437);
xor U10220 (N_10220,N_8179,N_9995);
nand U10221 (N_10221,N_7860,N_7389);
or U10222 (N_10222,N_6387,N_7152);
or U10223 (N_10223,N_5981,N_6119);
or U10224 (N_10224,N_9390,N_6926);
or U10225 (N_10225,N_9364,N_9949);
xor U10226 (N_10226,N_5444,N_8094);
nor U10227 (N_10227,N_6539,N_5413);
and U10228 (N_10228,N_9484,N_5350);
nor U10229 (N_10229,N_5675,N_6913);
and U10230 (N_10230,N_6303,N_5221);
or U10231 (N_10231,N_9050,N_7636);
and U10232 (N_10232,N_7596,N_9620);
and U10233 (N_10233,N_9296,N_6388);
and U10234 (N_10234,N_5164,N_6879);
or U10235 (N_10235,N_8031,N_9506);
or U10236 (N_10236,N_7048,N_8537);
nand U10237 (N_10237,N_9600,N_8444);
nand U10238 (N_10238,N_6503,N_7205);
or U10239 (N_10239,N_5942,N_8866);
or U10240 (N_10240,N_9088,N_7562);
nand U10241 (N_10241,N_8705,N_6822);
and U10242 (N_10242,N_7938,N_9536);
nand U10243 (N_10243,N_8104,N_6813);
and U10244 (N_10244,N_7163,N_8411);
xor U10245 (N_10245,N_7812,N_5152);
xor U10246 (N_10246,N_7433,N_9546);
nand U10247 (N_10247,N_5543,N_8519);
nand U10248 (N_10248,N_5893,N_6591);
nand U10249 (N_10249,N_8029,N_6895);
nand U10250 (N_10250,N_7989,N_6500);
xnor U10251 (N_10251,N_8722,N_5791);
and U10252 (N_10252,N_7321,N_5929);
or U10253 (N_10253,N_5719,N_6274);
xor U10254 (N_10254,N_9899,N_6456);
nor U10255 (N_10255,N_5706,N_5247);
nand U10256 (N_10256,N_8124,N_5467);
nor U10257 (N_10257,N_9326,N_8829);
and U10258 (N_10258,N_9170,N_6544);
or U10259 (N_10259,N_7492,N_7649);
and U10260 (N_10260,N_9357,N_6897);
and U10261 (N_10261,N_6579,N_6306);
nor U10262 (N_10262,N_8459,N_5336);
nor U10263 (N_10263,N_6908,N_6703);
or U10264 (N_10264,N_6678,N_6127);
nor U10265 (N_10265,N_8135,N_6427);
xor U10266 (N_10266,N_8762,N_8713);
nand U10267 (N_10267,N_7851,N_6102);
and U10268 (N_10268,N_5387,N_5657);
and U10269 (N_10269,N_9623,N_5469);
xnor U10270 (N_10270,N_8096,N_6273);
nor U10271 (N_10271,N_6550,N_8316);
and U10272 (N_10272,N_7256,N_6042);
xnor U10273 (N_10273,N_8477,N_8505);
nor U10274 (N_10274,N_6161,N_7427);
nand U10275 (N_10275,N_9925,N_6770);
and U10276 (N_10276,N_8321,N_7984);
nand U10277 (N_10277,N_9449,N_8590);
nand U10278 (N_10278,N_7239,N_5670);
nand U10279 (N_10279,N_7122,N_8962);
xor U10280 (N_10280,N_7216,N_9791);
nor U10281 (N_10281,N_6198,N_5600);
and U10282 (N_10282,N_6802,N_7138);
nand U10283 (N_10283,N_7463,N_8146);
nor U10284 (N_10284,N_5954,N_7785);
nor U10285 (N_10285,N_7053,N_9504);
or U10286 (N_10286,N_8911,N_5574);
or U10287 (N_10287,N_5411,N_5084);
or U10288 (N_10288,N_6103,N_6110);
nand U10289 (N_10289,N_7306,N_5463);
nor U10290 (N_10290,N_8600,N_5253);
nor U10291 (N_10291,N_9709,N_8348);
nor U10292 (N_10292,N_9015,N_8704);
nand U10293 (N_10293,N_8077,N_8319);
and U10294 (N_10294,N_9141,N_9126);
or U10295 (N_10295,N_5724,N_7188);
xor U10296 (N_10296,N_7502,N_9201);
nand U10297 (N_10297,N_8944,N_5349);
nand U10298 (N_10298,N_7140,N_6269);
nor U10299 (N_10299,N_7987,N_5923);
xnor U10300 (N_10300,N_8020,N_9000);
xor U10301 (N_10301,N_5231,N_8865);
nand U10302 (N_10302,N_9468,N_5069);
xnor U10303 (N_10303,N_6729,N_7754);
nor U10304 (N_10304,N_6628,N_5410);
nand U10305 (N_10305,N_5282,N_7114);
and U10306 (N_10306,N_6588,N_9769);
nand U10307 (N_10307,N_9929,N_5245);
and U10308 (N_10308,N_6174,N_5939);
nor U10309 (N_10309,N_7160,N_8510);
nand U10310 (N_10310,N_5885,N_5301);
xor U10311 (N_10311,N_9702,N_5964);
nor U10312 (N_10312,N_7846,N_6243);
nor U10313 (N_10313,N_9915,N_6595);
nand U10314 (N_10314,N_8210,N_9277);
or U10315 (N_10315,N_5624,N_5750);
and U10316 (N_10316,N_6788,N_7637);
and U10317 (N_10317,N_9762,N_8162);
xor U10318 (N_10318,N_7632,N_7675);
nand U10319 (N_10319,N_8783,N_5306);
or U10320 (N_10320,N_7317,N_7749);
nor U10321 (N_10321,N_5408,N_7576);
nor U10322 (N_10322,N_9745,N_7814);
nand U10323 (N_10323,N_8436,N_6007);
or U10324 (N_10324,N_7825,N_8999);
nand U10325 (N_10325,N_7299,N_9870);
nand U10326 (N_10326,N_7780,N_8854);
or U10327 (N_10327,N_9686,N_9992);
nor U10328 (N_10328,N_6627,N_8264);
nand U10329 (N_10329,N_9024,N_5493);
or U10330 (N_10330,N_8709,N_6644);
nand U10331 (N_10331,N_8191,N_8718);
and U10332 (N_10332,N_5378,N_9120);
and U10333 (N_10333,N_8670,N_7699);
nand U10334 (N_10334,N_9651,N_7339);
or U10335 (N_10335,N_9380,N_7788);
nor U10336 (N_10336,N_7581,N_7294);
xor U10337 (N_10337,N_9843,N_8758);
and U10338 (N_10338,N_5525,N_9433);
or U10339 (N_10339,N_6354,N_7599);
or U10340 (N_10340,N_9954,N_5966);
nor U10341 (N_10341,N_5478,N_7328);
or U10342 (N_10342,N_5688,N_5395);
xnor U10343 (N_10343,N_9451,N_8352);
xor U10344 (N_10344,N_5105,N_6064);
and U10345 (N_10345,N_6370,N_6969);
nand U10346 (N_10346,N_9173,N_8902);
nor U10347 (N_10347,N_9035,N_9119);
nand U10348 (N_10348,N_7639,N_8513);
and U10349 (N_10349,N_6725,N_7534);
or U10350 (N_10350,N_5546,N_6467);
nor U10351 (N_10351,N_5262,N_8086);
or U10352 (N_10352,N_8034,N_8511);
and U10353 (N_10353,N_7976,N_7647);
and U10354 (N_10354,N_9597,N_7621);
and U10355 (N_10355,N_8102,N_5669);
xor U10356 (N_10356,N_8701,N_7951);
nand U10357 (N_10357,N_8953,N_7640);
nand U10358 (N_10358,N_6763,N_7725);
or U10359 (N_10359,N_6474,N_7268);
xnor U10360 (N_10360,N_8063,N_5591);
and U10361 (N_10361,N_5875,N_5208);
and U10362 (N_10362,N_6555,N_5722);
or U10363 (N_10363,N_9047,N_6662);
xnor U10364 (N_10364,N_8601,N_5542);
or U10365 (N_10365,N_7654,N_5437);
and U10366 (N_10366,N_9323,N_6019);
xor U10367 (N_10367,N_5985,N_8045);
or U10368 (N_10368,N_9540,N_7771);
nor U10369 (N_10369,N_5658,N_5639);
nand U10370 (N_10370,N_8228,N_7618);
nor U10371 (N_10371,N_9722,N_8766);
nor U10372 (N_10372,N_5743,N_9789);
and U10373 (N_10373,N_7828,N_7426);
xnor U10374 (N_10374,N_8066,N_7722);
or U10375 (N_10375,N_7407,N_5540);
xor U10376 (N_10376,N_6869,N_8786);
nor U10377 (N_10377,N_5962,N_7166);
and U10378 (N_10378,N_7697,N_7134);
nand U10379 (N_10379,N_6596,N_9490);
nor U10380 (N_10380,N_6866,N_5814);
nand U10381 (N_10381,N_7519,N_6724);
and U10382 (N_10382,N_5686,N_6233);
nor U10383 (N_10383,N_7819,N_6587);
and U10384 (N_10384,N_7743,N_7777);
nor U10385 (N_10385,N_5147,N_8605);
nor U10386 (N_10386,N_7423,N_7197);
or U10387 (N_10387,N_9099,N_5058);
nor U10388 (N_10388,N_8576,N_6096);
nor U10389 (N_10389,N_8430,N_6613);
nor U10390 (N_10390,N_5312,N_7102);
and U10391 (N_10391,N_9263,N_6754);
or U10392 (N_10392,N_7961,N_8567);
nor U10393 (N_10393,N_9571,N_7821);
or U10394 (N_10394,N_5273,N_6972);
or U10395 (N_10395,N_9496,N_8700);
or U10396 (N_10396,N_9978,N_9400);
or U10397 (N_10397,N_7966,N_6658);
nand U10398 (N_10398,N_8834,N_8621);
nand U10399 (N_10399,N_9419,N_7885);
or U10400 (N_10400,N_7630,N_8460);
nor U10401 (N_10401,N_5146,N_6346);
and U10402 (N_10402,N_5334,N_6505);
xnor U10403 (N_10403,N_7149,N_6648);
or U10404 (N_10404,N_7032,N_9278);
nor U10405 (N_10405,N_6009,N_8379);
nor U10406 (N_10406,N_5520,N_7751);
nand U10407 (N_10407,N_9391,N_7063);
nor U10408 (N_10408,N_5093,N_7024);
xor U10409 (N_10409,N_9521,N_8814);
and U10410 (N_10410,N_6069,N_6461);
or U10411 (N_10411,N_7895,N_8565);
xor U10412 (N_10412,N_8798,N_8681);
or U10413 (N_10413,N_7014,N_8467);
xor U10414 (N_10414,N_6842,N_6199);
and U10415 (N_10415,N_6889,N_6394);
or U10416 (N_10416,N_8815,N_6248);
and U10417 (N_10417,N_7658,N_5541);
nand U10418 (N_10418,N_6143,N_8934);
nor U10419 (N_10419,N_6736,N_9566);
and U10420 (N_10420,N_5569,N_6605);
or U10421 (N_10421,N_7817,N_7858);
and U10422 (N_10422,N_6141,N_6614);
xor U10423 (N_10423,N_9053,N_9721);
xor U10424 (N_10424,N_6135,N_6195);
xor U10425 (N_10425,N_9315,N_7054);
and U10426 (N_10426,N_9184,N_9591);
nor U10427 (N_10427,N_7594,N_8109);
or U10428 (N_10428,N_6334,N_5926);
nor U10429 (N_10429,N_7405,N_9905);
nor U10430 (N_10430,N_5871,N_5007);
or U10431 (N_10431,N_7681,N_7892);
and U10432 (N_10432,N_5979,N_6258);
xor U10433 (N_10433,N_9483,N_8544);
nand U10434 (N_10434,N_5445,N_7145);
and U10435 (N_10435,N_6845,N_6988);
and U10436 (N_10436,N_5040,N_6823);
or U10437 (N_10437,N_6840,N_6207);
and U10438 (N_10438,N_8559,N_6911);
nor U10439 (N_10439,N_7680,N_5142);
or U10440 (N_10440,N_5854,N_5841);
or U10441 (N_10441,N_9448,N_9956);
or U10442 (N_10442,N_8799,N_8885);
and U10443 (N_10443,N_9716,N_8957);
xor U10444 (N_10444,N_9828,N_9629);
and U10445 (N_10445,N_5890,N_5188);
nand U10446 (N_10446,N_5599,N_5140);
xnor U10447 (N_10447,N_8201,N_5201);
and U10448 (N_10448,N_5565,N_5392);
nor U10449 (N_10449,N_5020,N_9305);
nor U10450 (N_10450,N_5223,N_8904);
or U10451 (N_10451,N_7531,N_8781);
nor U10452 (N_10452,N_5583,N_5446);
nor U10453 (N_10453,N_5449,N_8492);
xnor U10454 (N_10454,N_7696,N_7673);
or U10455 (N_10455,N_5994,N_8737);
and U10456 (N_10456,N_7678,N_9059);
nand U10457 (N_10457,N_6239,N_8903);
nor U10458 (N_10458,N_6899,N_9331);
xnor U10459 (N_10459,N_6910,N_7043);
and U10460 (N_10460,N_8067,N_5718);
nand U10461 (N_10461,N_5832,N_7387);
nand U10462 (N_10462,N_9885,N_6499);
nor U10463 (N_10463,N_7308,N_9282);
nor U10464 (N_10464,N_8447,N_9523);
and U10465 (N_10465,N_9293,N_8255);
xor U10466 (N_10466,N_6205,N_8483);
xnor U10467 (N_10467,N_6685,N_5984);
nor U10468 (N_10468,N_7994,N_5866);
or U10469 (N_10469,N_5552,N_8730);
or U10470 (N_10470,N_9353,N_6782);
or U10471 (N_10471,N_8216,N_5296);
nor U10472 (N_10472,N_5037,N_9136);
nor U10473 (N_10473,N_9429,N_6399);
nand U10474 (N_10474,N_8392,N_9028);
or U10475 (N_10475,N_9985,N_9113);
and U10476 (N_10476,N_6671,N_6833);
nor U10477 (N_10477,N_5496,N_8190);
nand U10478 (N_10478,N_5965,N_5401);
nor U10479 (N_10479,N_5566,N_6738);
nand U10480 (N_10480,N_5298,N_8329);
nand U10481 (N_10481,N_5702,N_5666);
nand U10482 (N_10482,N_7577,N_6379);
or U10483 (N_10483,N_5742,N_7866);
and U10484 (N_10484,N_6032,N_9817);
or U10485 (N_10485,N_7093,N_8337);
and U10486 (N_10486,N_5785,N_7029);
nand U10487 (N_10487,N_6231,N_7004);
xor U10488 (N_10488,N_9846,N_9133);
xnor U10489 (N_10489,N_5441,N_6381);
or U10490 (N_10490,N_7815,N_6145);
nand U10491 (N_10491,N_9011,N_5427);
nand U10492 (N_10492,N_8236,N_6116);
nor U10493 (N_10493,N_8859,N_9514);
or U10494 (N_10494,N_8189,N_6956);
or U10495 (N_10495,N_7362,N_8914);
or U10496 (N_10496,N_9881,N_7499);
nand U10497 (N_10497,N_6044,N_9021);
and U10498 (N_10498,N_9004,N_9418);
or U10499 (N_10499,N_5377,N_6516);
and U10500 (N_10500,N_7291,N_5380);
and U10501 (N_10501,N_9734,N_9402);
and U10502 (N_10502,N_5616,N_6819);
xor U10503 (N_10503,N_8013,N_5709);
xnor U10504 (N_10504,N_6519,N_8290);
and U10505 (N_10505,N_5393,N_8362);
or U10506 (N_10506,N_5316,N_6196);
and U10507 (N_10507,N_8372,N_7865);
xor U10508 (N_10508,N_6536,N_5562);
nor U10509 (N_10509,N_7496,N_5091);
nor U10510 (N_10510,N_8752,N_8199);
or U10511 (N_10511,N_5815,N_9701);
nor U10512 (N_10512,N_5958,N_7598);
nor U10513 (N_10513,N_9933,N_6504);
xnor U10514 (N_10514,N_5353,N_8182);
or U10515 (N_10515,N_9215,N_5803);
xor U10516 (N_10516,N_5219,N_8661);
nor U10517 (N_10517,N_7302,N_7047);
and U10518 (N_10518,N_5944,N_5206);
or U10519 (N_10519,N_5568,N_9510);
nand U10520 (N_10520,N_5220,N_9602);
and U10521 (N_10521,N_6003,N_7880);
nor U10522 (N_10522,N_5032,N_7109);
and U10523 (N_10523,N_9381,N_9410);
or U10524 (N_10524,N_7028,N_6715);
and U10525 (N_10525,N_9345,N_9939);
and U10526 (N_10526,N_6675,N_5537);
nor U10527 (N_10527,N_5315,N_6633);
nand U10528 (N_10528,N_6098,N_8938);
xnor U10529 (N_10529,N_5907,N_6309);
xnor U10530 (N_10530,N_7007,N_7940);
xnor U10531 (N_10531,N_8133,N_6875);
or U10532 (N_10532,N_5250,N_7397);
and U10533 (N_10533,N_6679,N_6371);
or U10534 (N_10534,N_5733,N_5745);
or U10535 (N_10535,N_6230,N_9124);
nand U10536 (N_10536,N_5641,N_7318);
nor U10537 (N_10537,N_9083,N_9269);
or U10538 (N_10538,N_5125,N_6202);
nand U10539 (N_10539,N_6874,N_6170);
xnor U10540 (N_10540,N_9657,N_8304);
xnor U10541 (N_10541,N_7135,N_9930);
or U10542 (N_10542,N_7322,N_6669);
nor U10543 (N_10543,N_9031,N_7563);
nand U10544 (N_10544,N_7731,N_7030);
or U10545 (N_10545,N_7886,N_7898);
or U10546 (N_10546,N_7916,N_7257);
and U10547 (N_10547,N_8089,N_8231);
xor U10548 (N_10548,N_9441,N_7653);
xnor U10549 (N_10549,N_6320,N_7920);
nand U10550 (N_10550,N_9271,N_7019);
or U10551 (N_10551,N_8749,N_6772);
and U10552 (N_10552,N_7184,N_8742);
and U10553 (N_10553,N_6850,N_5524);
nor U10554 (N_10554,N_9526,N_7334);
or U10555 (N_10555,N_9866,N_5630);
and U10556 (N_10556,N_8330,N_9880);
or U10557 (N_10557,N_7401,N_5830);
nand U10558 (N_10558,N_7142,N_5210);
nand U10559 (N_10559,N_6192,N_6557);
or U10560 (N_10560,N_7784,N_6213);
nand U10561 (N_10561,N_7803,N_9927);
and U10562 (N_10562,N_8455,N_5287);
xnor U10563 (N_10563,N_5654,N_6830);
xnor U10564 (N_10564,N_7835,N_9516);
or U10565 (N_10565,N_6489,N_8582);
nand U10566 (N_10566,N_9343,N_9210);
xor U10567 (N_10567,N_6909,N_7572);
xnor U10568 (N_10568,N_5276,N_6812);
nor U10569 (N_10569,N_6089,N_8826);
nand U10570 (N_10570,N_9593,N_5357);
and U10571 (N_10571,N_6348,N_7739);
nand U10572 (N_10572,N_9604,N_7723);
or U10573 (N_10573,N_5589,N_5390);
and U10574 (N_10574,N_7765,N_9796);
xor U10575 (N_10575,N_8422,N_9581);
nor U10576 (N_10576,N_7904,N_5936);
and U10577 (N_10577,N_6817,N_5488);
nand U10578 (N_10578,N_9639,N_6209);
or U10579 (N_10579,N_9499,N_9445);
nor U10580 (N_10580,N_9610,N_8978);
and U10581 (N_10581,N_9776,N_5897);
and U10582 (N_10582,N_5764,N_9541);
xor U10583 (N_10583,N_8603,N_9570);
nand U10584 (N_10584,N_7022,N_8275);
nand U10585 (N_10585,N_7280,N_5855);
and U10586 (N_10586,N_5010,N_8280);
and U10587 (N_10587,N_5291,N_9898);
xnor U10588 (N_10588,N_5680,N_6290);
nor U10589 (N_10589,N_6700,N_8882);
nor U10590 (N_10590,N_6657,N_7622);
or U10591 (N_10591,N_7578,N_5230);
or U10592 (N_10592,N_8284,N_7887);
and U10593 (N_10593,N_9712,N_9725);
nand U10594 (N_10594,N_8679,N_7774);
xnor U10595 (N_10595,N_5376,N_5453);
nand U10596 (N_10596,N_5695,N_7655);
or U10597 (N_10597,N_7026,N_8852);
and U10598 (N_10598,N_7064,N_8030);
or U10599 (N_10599,N_8355,N_6645);
or U10600 (N_10600,N_5174,N_9900);
nor U10601 (N_10601,N_6319,N_8721);
nand U10602 (N_10602,N_5952,N_5886);
or U10603 (N_10603,N_5590,N_8971);
nand U10604 (N_10604,N_5823,N_9186);
xnor U10605 (N_10605,N_9144,N_5181);
nor U10606 (N_10606,N_5218,N_9492);
and U10607 (N_10607,N_5506,N_8847);
nor U10608 (N_10608,N_8192,N_6745);
nand U10609 (N_10609,N_6412,N_5526);
xor U10610 (N_10610,N_6413,N_5613);
nor U10611 (N_10611,N_9087,N_9829);
xor U10612 (N_10612,N_7511,N_9106);
and U10613 (N_10613,N_6635,N_7694);
or U10614 (N_10614,N_8286,N_5251);
and U10615 (N_10615,N_5465,N_8548);
or U10616 (N_10616,N_5295,N_7507);
or U10617 (N_10617,N_9036,N_9732);
and U10618 (N_10618,N_8972,N_9592);
and U10619 (N_10619,N_6178,N_6618);
nand U10620 (N_10620,N_9626,N_9811);
and U10621 (N_10621,N_8846,N_8926);
nand U10622 (N_10622,N_9251,N_9137);
xor U10623 (N_10623,N_9569,N_6963);
or U10624 (N_10624,N_7611,N_9159);
nor U10625 (N_10625,N_8383,N_6479);
or U10626 (N_10626,N_6245,N_7057);
or U10627 (N_10627,N_6353,N_7954);
and U10628 (N_10628,N_6801,N_6610);
xor U10629 (N_10629,N_6814,N_6728);
nor U10630 (N_10630,N_5405,N_7000);
xor U10631 (N_10631,N_5651,N_8103);
and U10632 (N_10632,N_8806,N_9498);
and U10633 (N_10633,N_9801,N_8308);
nand U10634 (N_10634,N_5026,N_5911);
or U10635 (N_10635,N_5224,N_5946);
and U10636 (N_10636,N_7174,N_9741);
or U10637 (N_10637,N_8481,N_5163);
xor U10638 (N_10638,N_7539,N_7279);
nand U10639 (N_10639,N_5730,N_5337);
and U10640 (N_10640,N_6886,N_9676);
or U10641 (N_10641,N_7663,N_5818);
or U10642 (N_10642,N_5254,N_7286);
nor U10643 (N_10643,N_7374,N_9199);
or U10644 (N_10644,N_9226,N_8325);
and U10645 (N_10645,N_6172,N_8778);
xor U10646 (N_10646,N_5849,N_7515);
nor U10647 (N_10647,N_6986,N_8004);
nand U10648 (N_10648,N_7570,N_7255);
xor U10649 (N_10649,N_6711,N_8421);
nor U10650 (N_10650,N_6002,N_7207);
nor U10651 (N_10651,N_6629,N_7020);
nor U10652 (N_10652,N_6904,N_7588);
nand U10653 (N_10653,N_8877,N_5551);
xnor U10654 (N_10654,N_9858,N_9831);
nand U10655 (N_10655,N_9426,N_9312);
nor U10656 (N_10656,N_6015,N_8131);
or U10657 (N_10657,N_9358,N_6490);
xnor U10658 (N_10658,N_9304,N_5732);
nor U10659 (N_10659,N_9275,N_5851);
or U10660 (N_10660,N_7176,N_7937);
nand U10661 (N_10661,N_9231,N_8106);
and U10662 (N_10662,N_6024,N_8837);
xor U10663 (N_10663,N_7242,N_8991);
and U10664 (N_10664,N_9601,N_5074);
xnor U10665 (N_10665,N_5863,N_7789);
and U10666 (N_10666,N_9427,N_9238);
xor U10667 (N_10667,N_9901,N_6598);
xor U10668 (N_10668,N_6771,N_6793);
nor U10669 (N_10669,N_9042,N_9987);
or U10670 (N_10670,N_8952,N_9300);
and U10671 (N_10671,N_8415,N_6735);
and U10672 (N_10672,N_5011,N_8560);
nor U10673 (N_10673,N_9664,N_7762);
xnor U10674 (N_10674,N_7971,N_7475);
nor U10675 (N_10675,N_8672,N_9708);
xor U10676 (N_10676,N_6208,N_6366);
or U10677 (N_10677,N_6878,N_8251);
xor U10678 (N_10678,N_5781,N_6402);
or U10679 (N_10679,N_8009,N_5100);
or U10680 (N_10680,N_9731,N_7728);
xor U10681 (N_10681,N_7050,N_7891);
nand U10682 (N_10682,N_7635,N_8514);
nor U10683 (N_10683,N_9757,N_6386);
and U10684 (N_10684,N_7326,N_9097);
nand U10685 (N_10685,N_6443,N_5793);
nand U10686 (N_10686,N_9049,N_8040);
or U10687 (N_10687,N_8003,N_8019);
or U10688 (N_10688,N_5880,N_8690);
nand U10689 (N_10689,N_7781,N_6803);
nor U10690 (N_10690,N_6260,N_7190);
or U10691 (N_10691,N_8178,N_9878);
and U10692 (N_10692,N_9549,N_7169);
or U10693 (N_10693,N_5114,N_6966);
nand U10694 (N_10694,N_8732,N_5554);
nor U10695 (N_10695,N_8153,N_8300);
nand U10696 (N_10696,N_8503,N_9208);
nor U10697 (N_10697,N_5132,N_8869);
or U10698 (N_10698,N_5644,N_7614);
nor U10699 (N_10699,N_9859,N_7101);
nand U10700 (N_10700,N_5458,N_8405);
nand U10701 (N_10701,N_5977,N_6293);
nand U10702 (N_10702,N_5993,N_8397);
xor U10703 (N_10703,N_5980,N_8174);
and U10704 (N_10704,N_7332,N_5848);
and U10705 (N_10705,N_7566,N_9440);
xnor U10706 (N_10706,N_6721,N_6155);
nor U10707 (N_10707,N_7608,N_9631);
nor U10708 (N_10708,N_6478,N_5189);
nor U10709 (N_10709,N_7480,N_5207);
and U10710 (N_10710,N_5003,N_7922);
xor U10711 (N_10711,N_5272,N_9459);
nand U10712 (N_10712,N_8160,N_6111);
nand U10713 (N_10713,N_8008,N_5580);
xor U10714 (N_10714,N_8912,N_7795);
or U10715 (N_10715,N_9627,N_9596);
and U10716 (N_10716,N_6025,N_6741);
nand U10717 (N_10717,N_5731,N_9847);
nor U10718 (N_10718,N_7429,N_6666);
nand U10719 (N_10719,N_8028,N_8326);
xor U10720 (N_10720,N_6834,N_5726);
nand U10721 (N_10721,N_6357,N_9382);
nor U10722 (N_10722,N_5527,N_8739);
nand U10723 (N_10723,N_9813,N_6507);
xnor U10724 (N_10724,N_6142,N_5048);
or U10725 (N_10725,N_7738,N_7117);
nor U10726 (N_10726,N_7144,N_7130);
and U10727 (N_10727,N_7607,N_6338);
and U10728 (N_10728,N_9336,N_9288);
or U10729 (N_10729,N_9491,N_7327);
xor U10730 (N_10730,N_6028,N_6789);
or U10731 (N_10731,N_6101,N_7882);
and U10732 (N_10732,N_8138,N_9633);
xor U10733 (N_10733,N_8738,N_7089);
nor U10734 (N_10734,N_7553,N_9756);
xnor U10735 (N_10735,N_7509,N_8589);
xor U10736 (N_10736,N_6574,N_6730);
nor U10737 (N_10737,N_9645,N_7449);
and U10738 (N_10738,N_5335,N_9041);
xor U10739 (N_10739,N_9554,N_9469);
nand U10740 (N_10740,N_7716,N_6470);
nor U10741 (N_10741,N_8056,N_6484);
nand U10742 (N_10742,N_7527,N_6699);
or U10743 (N_10743,N_9787,N_8091);
nand U10744 (N_10744,N_9781,N_6183);
xor U10745 (N_10745,N_9280,N_9910);
nor U10746 (N_10746,N_5433,N_5787);
nand U10747 (N_10747,N_6514,N_6885);
and U10748 (N_10748,N_6777,N_8703);
or U10749 (N_10749,N_6308,N_5736);
nor U10750 (N_10750,N_7107,N_9246);
nand U10751 (N_10751,N_9854,N_7215);
nor U10752 (N_10752,N_9700,N_6080);
and U10753 (N_10753,N_5480,N_9675);
and U10754 (N_10754,N_5416,N_9668);
or U10755 (N_10755,N_5447,N_5283);
nor U10756 (N_10756,N_9330,N_8006);
nand U10757 (N_10757,N_7005,N_6077);
xnor U10758 (N_10758,N_6341,N_6767);
nor U10759 (N_10759,N_6764,N_9594);
or U10760 (N_10760,N_9081,N_5829);
and U10761 (N_10761,N_7106,N_5518);
and U10762 (N_10762,N_6468,N_7461);
xnor U10763 (N_10763,N_7718,N_5232);
and U10764 (N_10764,N_5124,N_7909);
or U10765 (N_10765,N_6575,N_9658);
or U10766 (N_10766,N_7128,N_8295);
or U10767 (N_10767,N_8012,N_9387);
nor U10768 (N_10768,N_5899,N_8886);
xor U10769 (N_10769,N_6784,N_6776);
nand U10770 (N_10770,N_9307,N_8076);
nor U10771 (N_10771,N_5833,N_7849);
nand U10772 (N_10772,N_6820,N_7099);
and U10773 (N_10773,N_7472,N_7960);
and U10774 (N_10774,N_9972,N_9963);
nor U10775 (N_10775,N_6983,N_8658);
and U10776 (N_10776,N_6453,N_9643);
nand U10777 (N_10777,N_6404,N_5214);
xnor U10778 (N_10778,N_5747,N_9172);
nand U10779 (N_10779,N_8696,N_7357);
and U10780 (N_10780,N_5195,N_6176);
nor U10781 (N_10781,N_7146,N_9882);
nand U10782 (N_10782,N_8309,N_7331);
xor U10783 (N_10783,N_8569,N_8487);
nand U10784 (N_10784,N_9897,N_5346);
nand U10785 (N_10785,N_5477,N_9295);
or U10786 (N_10786,N_7729,N_8354);
or U10787 (N_10787,N_6425,N_6259);
nor U10788 (N_10788,N_5799,N_5213);
nand U10789 (N_10789,N_6808,N_8745);
nand U10790 (N_10790,N_9953,N_9495);
nand U10791 (N_10791,N_5735,N_6731);
xnor U10792 (N_10792,N_6751,N_5925);
xnor U10793 (N_10793,N_5073,N_5634);
and U10794 (N_10794,N_8328,N_8278);
nand U10795 (N_10795,N_6975,N_8729);
or U10796 (N_10796,N_6442,N_8128);
or U10797 (N_10797,N_7670,N_7441);
xnor U10798 (N_10798,N_6095,N_7345);
and U10799 (N_10799,N_6901,N_7616);
xnor U10800 (N_10800,N_8593,N_7501);
or U10801 (N_10801,N_5579,N_5005);
xor U10802 (N_10802,N_7477,N_9109);
xor U10803 (N_10803,N_5544,N_6948);
and U10804 (N_10804,N_5209,N_5820);
nand U10805 (N_10805,N_9761,N_5619);
nor U10806 (N_10806,N_5025,N_9733);
nand U10807 (N_10807,N_5852,N_7393);
and U10808 (N_10808,N_8581,N_6229);
or U10809 (N_10809,N_7874,N_9414);
xor U10810 (N_10810,N_7532,N_7371);
xnor U10811 (N_10811,N_8149,N_9947);
nand U10812 (N_10812,N_5304,N_9578);
nand U10813 (N_10813,N_6099,N_6906);
xnor U10814 (N_10814,N_8425,N_8198);
xor U10815 (N_10815,N_9267,N_5184);
xnor U10816 (N_10816,N_5883,N_5713);
nor U10817 (N_10817,N_7119,N_5332);
nor U10818 (N_10818,N_5060,N_6498);
nand U10819 (N_10819,N_6619,N_6112);
xnor U10820 (N_10820,N_6734,N_9299);
nand U10821 (N_10821,N_7153,N_8347);
nand U10822 (N_10822,N_7460,N_9853);
nor U10823 (N_10823,N_5268,N_5759);
nand U10824 (N_10824,N_6302,N_9347);
nand U10825 (N_10825,N_7439,N_9167);
and U10826 (N_10826,N_6791,N_8384);
nand U10827 (N_10827,N_8249,N_8152);
nor U10828 (N_10828,N_6753,N_6804);
or U10829 (N_10829,N_6779,N_6426);
nand U10830 (N_10830,N_7451,N_7021);
and U10831 (N_10831,N_8945,N_9385);
nand U10832 (N_10832,N_6698,N_5324);
nor U10833 (N_10833,N_5650,N_6710);
nand U10834 (N_10834,N_6224,N_8941);
or U10835 (N_10835,N_6858,N_6836);
or U10836 (N_10836,N_9074,N_5319);
nor U10837 (N_10837,N_7348,N_5085);
nand U10838 (N_10838,N_6905,N_7249);
nor U10839 (N_10839,N_8947,N_7385);
nand U10840 (N_10840,N_6888,N_7406);
and U10841 (N_10841,N_9487,N_5805);
or U10842 (N_10842,N_8970,N_7121);
or U10843 (N_10843,N_6298,N_6643);
and U10844 (N_10844,N_8155,N_9976);
nor U10845 (N_10845,N_6118,N_8523);
and U10846 (N_10846,N_9790,N_6179);
or U10847 (N_10847,N_9691,N_7016);
xor U10848 (N_10848,N_6473,N_6702);
and U10849 (N_10849,N_9852,N_7770);
or U10850 (N_10850,N_6414,N_8861);
or U10851 (N_10851,N_7447,N_7258);
or U10852 (N_10852,N_9232,N_9553);
or U10853 (N_10853,N_6634,N_7290);
and U10854 (N_10854,N_5111,N_5681);
xnor U10855 (N_10855,N_6185,N_9058);
or U10856 (N_10856,N_8011,N_8053);
nand U10857 (N_10857,N_8205,N_9753);
nor U10858 (N_10858,N_8026,N_6140);
xor U10859 (N_10859,N_5162,N_6872);
and U10860 (N_10860,N_6339,N_7200);
nor U10861 (N_10861,N_6482,N_5768);
or U10862 (N_10862,N_9574,N_8310);
and U10863 (N_10863,N_6459,N_6611);
or U10864 (N_10864,N_8140,N_6923);
nor U10865 (N_10865,N_7933,N_9577);
nor U10866 (N_10866,N_7319,N_9194);
nand U10867 (N_10867,N_9763,N_5148);
and U10868 (N_10868,N_8250,N_9653);
xor U10869 (N_10869,N_9759,N_7683);
or U10870 (N_10870,N_5618,N_6894);
and U10871 (N_10871,N_8242,N_5626);
and U10872 (N_10872,N_7262,N_6061);
xor U10873 (N_10873,N_7103,N_8409);
nor U10874 (N_10874,N_8659,N_7682);
xor U10875 (N_10875,N_5351,N_8212);
xnor U10876 (N_10876,N_8617,N_9966);
nor U10877 (N_10877,N_5424,N_7834);
nor U10878 (N_10878,N_8813,N_7805);
and U10879 (N_10879,N_5762,N_9559);
or U10880 (N_10880,N_6329,N_6405);
nor U10881 (N_10881,N_6765,N_7310);
nand U10882 (N_10882,N_8240,N_8206);
nand U10883 (N_10883,N_6520,N_8039);
or U10884 (N_10884,N_6674,N_9228);
and U10885 (N_10885,N_9009,N_7303);
nor U10886 (N_10886,N_7962,N_5629);
or U10887 (N_10887,N_9973,N_9196);
and U10888 (N_10888,N_5753,N_7816);
or U10889 (N_10889,N_9457,N_6951);
and U10890 (N_10890,N_5456,N_9924);
nand U10891 (N_10891,N_8915,N_7669);
nor U10892 (N_10892,N_8098,N_9568);
and U10893 (N_10893,N_6540,N_8181);
and U10894 (N_10894,N_8684,N_6300);
and U10895 (N_10895,N_9034,N_6389);
and U10896 (N_10896,N_7036,N_7436);
nor U10897 (N_10897,N_9533,N_6072);
xnor U10898 (N_10898,N_7112,N_5203);
nand U10899 (N_10899,N_9436,N_8157);
nor U10900 (N_10900,N_8664,N_7958);
nand U10901 (N_10901,N_5014,N_7528);
nor U10902 (N_10902,N_7364,N_9622);
or U10903 (N_10903,N_7444,N_6549);
xor U10904 (N_10904,N_8100,N_9372);
nand U10905 (N_10905,N_9872,N_9960);
or U10906 (N_10906,N_6530,N_5784);
xor U10907 (N_10907,N_9107,N_6989);
and U10908 (N_10908,N_9621,N_5329);
and U10909 (N_10909,N_9245,N_7070);
and U10910 (N_10910,N_6073,N_6996);
xor U10911 (N_10911,N_9816,N_5384);
xnor U10912 (N_10912,N_8297,N_7824);
xnor U10913 (N_10913,N_7727,N_6537);
or U10914 (N_10914,N_5517,N_6083);
xor U10915 (N_10915,N_9687,N_5035);
or U10916 (N_10916,N_6255,N_6810);
and U10917 (N_10917,N_6898,N_5264);
xor U10918 (N_10918,N_7790,N_5876);
nor U10919 (N_10919,N_5610,N_8269);
nor U10920 (N_10920,N_6382,N_9679);
nand U10921 (N_10921,N_6676,N_9022);
xor U10922 (N_10922,N_7533,N_6606);
nor U10923 (N_10923,N_6559,N_8433);
nand U10924 (N_10924,N_9713,N_6690);
or U10925 (N_10925,N_9752,N_5945);
nor U10926 (N_10926,N_6014,N_9524);
nand U10927 (N_10927,N_9988,N_5955);
nor U10928 (N_10928,N_6600,N_6766);
nor U10929 (N_10929,N_5077,N_6278);
and U10930 (N_10930,N_8812,N_7671);
xor U10931 (N_10931,N_9301,N_9189);
or U10932 (N_10932,N_5755,N_8342);
and U10933 (N_10933,N_8608,N_7006);
nor U10934 (N_10934,N_8343,N_7983);
xnor U10935 (N_10935,N_6310,N_9673);
or U10936 (N_10936,N_8353,N_6428);
and U10937 (N_10937,N_6477,N_9798);
and U10938 (N_10938,N_6631,N_7018);
or U10939 (N_10939,N_6203,N_5070);
xor U10940 (N_10940,N_9889,N_6705);
nand U10941 (N_10941,N_8177,N_7373);
or U10942 (N_10942,N_9517,N_5744);
nand U10943 (N_10943,N_5861,N_6177);
or U10944 (N_10944,N_6180,N_7747);
or U10945 (N_10945,N_8862,N_7617);
nor U10946 (N_10946,N_8185,N_6242);
and U10947 (N_10947,N_7361,N_9285);
xnor U10948 (N_10948,N_8906,N_5407);
xnor U10949 (N_10949,N_5783,N_7001);
xnor U10950 (N_10950,N_7236,N_8434);
nor U10951 (N_10951,N_6960,N_6835);
and U10952 (N_10952,N_5489,N_9014);
and U10953 (N_10953,N_8000,N_5691);
xor U10954 (N_10954,N_5679,N_9156);
xnor U10955 (N_10955,N_7162,N_8002);
or U10956 (N_10956,N_6131,N_7883);
xnor U10957 (N_10957,N_9785,N_7288);
nand U10958 (N_10958,N_8018,N_6190);
xor U10959 (N_10959,N_8055,N_8792);
xor U10960 (N_10960,N_7875,N_7307);
nor U10961 (N_10961,N_6533,N_5237);
xor U10962 (N_10962,N_6528,N_9851);
nand U10963 (N_10963,N_9287,N_6739);
or U10964 (N_10964,N_7034,N_6914);
and U10965 (N_10965,N_5648,N_5774);
nand U10966 (N_10966,N_5136,N_8263);
and U10967 (N_10967,N_8526,N_7224);
or U10968 (N_10968,N_5578,N_9247);
nand U10969 (N_10969,N_6576,N_9233);
or U10970 (N_10970,N_8753,N_5553);
xor U10971 (N_10971,N_9166,N_5472);
and U10972 (N_10972,N_8802,N_5041);
nand U10973 (N_10973,N_7042,N_7141);
xnor U10974 (N_10974,N_5913,N_9919);
nor U10975 (N_10975,N_7375,N_6030);
xor U10976 (N_10976,N_7997,N_5145);
nor U10977 (N_10977,N_7111,N_8288);
nand U10978 (N_10978,N_9647,N_8760);
nand U10979 (N_10979,N_7973,N_8539);
and U10980 (N_10980,N_9040,N_9968);
and U10981 (N_10981,N_5199,N_9415);
nand U10982 (N_10982,N_7457,N_8936);
or U10983 (N_10983,N_8653,N_7096);
nand U10984 (N_10984,N_5027,N_9582);
or U10985 (N_10985,N_9160,N_5608);
nor U10986 (N_10986,N_6376,N_9606);
nor U10987 (N_10987,N_6223,N_5640);
and U10988 (N_10988,N_7685,N_5462);
xor U10989 (N_10989,N_8871,N_9871);
and U10990 (N_10990,N_7180,N_5637);
nor U10991 (N_10991,N_6740,N_6432);
nand U10992 (N_10992,N_5459,N_8365);
or U10993 (N_10993,N_9356,N_6004);
and U10994 (N_10994,N_9758,N_8202);
and U10995 (N_10995,N_6927,N_8651);
or U10996 (N_10996,N_9443,N_9714);
and U10997 (N_10997,N_7629,N_6051);
nor U10998 (N_10998,N_6067,N_7737);
and U10999 (N_10999,N_7125,N_8118);
or U11000 (N_11000,N_9128,N_7137);
nor U11001 (N_11001,N_5935,N_6654);
and U11002 (N_11002,N_5794,N_8933);
nor U11003 (N_11003,N_9114,N_8527);
and U11004 (N_11004,N_8761,N_5150);
or U11005 (N_11005,N_8256,N_9378);
or U11006 (N_11006,N_5906,N_6139);
or U11007 (N_11007,N_5484,N_6356);
and U11008 (N_11008,N_5534,N_6944);
and U11009 (N_11009,N_7709,N_8797);
or U11010 (N_11010,N_9774,N_5233);
xor U11011 (N_11011,N_9912,N_6108);
nand U11012 (N_11012,N_6921,N_7237);
nand U11013 (N_11013,N_6561,N_6431);
nand U11014 (N_11014,N_8598,N_5586);
and U11015 (N_11015,N_9969,N_8079);
and U11016 (N_11016,N_5707,N_6138);
nor U11017 (N_11017,N_9070,N_5398);
and U11018 (N_11018,N_5143,N_8809);
nand U11019 (N_11019,N_8047,N_5450);
and U11020 (N_11020,N_8400,N_9174);
nand U11021 (N_11021,N_5588,N_9486);
nand U11022 (N_11022,N_7609,N_6457);
and U11023 (N_11023,N_7396,N_6637);
nand U11024 (N_11024,N_6228,N_8386);
or U11025 (N_11025,N_9359,N_5917);
or U11026 (N_11026,N_8475,N_5620);
xnor U11027 (N_11027,N_9063,N_6121);
xnor U11028 (N_11028,N_6696,N_7297);
and U11029 (N_11029,N_9032,N_6964);
or U11030 (N_11030,N_9529,N_5361);
and U11031 (N_11031,N_7446,N_8110);
xnor U11032 (N_11032,N_5677,N_8344);
and U11033 (N_11033,N_8763,N_5300);
or U11034 (N_11034,N_9253,N_9681);
nand U11035 (N_11035,N_6215,N_8587);
and U11036 (N_11036,N_5212,N_8992);
nand U11037 (N_11037,N_7133,N_7829);
nand U11038 (N_11038,N_6488,N_8461);
xnor U11039 (N_11039,N_7090,N_5877);
xor U11040 (N_11040,N_5693,N_5061);
nor U11041 (N_11041,N_5430,N_8338);
nand U11042 (N_11042,N_6659,N_8320);
or U11043 (N_11043,N_9209,N_5078);
xnor U11044 (N_11044,N_5019,N_9628);
or U11045 (N_11045,N_5536,N_5672);
nor U11046 (N_11046,N_5267,N_5079);
nand U11047 (N_11047,N_8183,N_6573);
xnor U11048 (N_11048,N_6890,N_5086);
xnor U11049 (N_11049,N_5509,N_7644);
nand U11050 (N_11050,N_6586,N_7315);
or U11051 (N_11051,N_9203,N_9660);
nor U11052 (N_11052,N_8801,N_8708);
xnor U11053 (N_11053,N_8463,N_9936);
and U11054 (N_11054,N_6194,N_6578);
and U11055 (N_11055,N_7818,N_8927);
nand U11056 (N_11056,N_6018,N_6147);
nor U11057 (N_11057,N_8816,N_6527);
or U11058 (N_11058,N_7347,N_5112);
or U11059 (N_11059,N_9887,N_8407);
xnor U11060 (N_11060,N_9255,N_7546);
or U11061 (N_11061,N_6673,N_7400);
nand U11062 (N_11062,N_7810,N_8323);
xor U11063 (N_11063,N_8557,N_6211);
xor U11064 (N_11064,N_9306,N_9420);
and U11065 (N_11065,N_5653,N_8154);
or U11066 (N_11066,N_9605,N_6439);
or U11067 (N_11067,N_6925,N_8782);
or U11068 (N_11068,N_6295,N_7206);
nand U11069 (N_11069,N_7841,N_6035);
xnor U11070 (N_11070,N_7701,N_7698);
and U11071 (N_11071,N_8426,N_8491);
or U11072 (N_11072,N_5615,N_5423);
or U11073 (N_11073,N_9821,N_9941);
and U11074 (N_11074,N_6164,N_8114);
or U11075 (N_11075,N_9886,N_9176);
or U11076 (N_11076,N_6225,N_6090);
nor U11077 (N_11077,N_8727,N_7672);
nand U11078 (N_11078,N_5308,N_9431);
and U11079 (N_11079,N_9862,N_7935);
nor U11080 (N_11080,N_8820,N_7398);
and U11081 (N_11081,N_9696,N_5059);
and U11082 (N_11082,N_8097,N_6458);
nor U11083 (N_11083,N_8509,N_8107);
nor U11084 (N_11084,N_5519,N_6762);
and U11085 (N_11085,N_6120,N_7076);
nand U11086 (N_11086,N_8230,N_7744);
xor U11087 (N_11087,N_7108,N_8318);
and U11088 (N_11088,N_9412,N_8443);
xor U11089 (N_11089,N_9931,N_6396);
xnor U11090 (N_11090,N_6222,N_7595);
and U11091 (N_11091,N_5912,N_5340);
nand U11092 (N_11092,N_5547,N_7623);
nor U11093 (N_11093,N_6057,N_6517);
xor U11094 (N_11094,N_8702,N_9051);
nand U11095 (N_11095,N_8517,N_7600);
nor U11096 (N_11096,N_7664,N_9565);
xnor U11097 (N_11097,N_5238,N_9694);
xnor U11098 (N_11098,N_9026,N_6263);
nor U11099 (N_11099,N_6922,N_7852);
nor U11100 (N_11100,N_8501,N_7888);
nand U11101 (N_11101,N_8825,N_7848);
and U11102 (N_11102,N_6460,N_7067);
nand U11103 (N_11103,N_9652,N_6773);
nand U11104 (N_11104,N_6792,N_7217);
or U11105 (N_11105,N_8973,N_6708);
or U11106 (N_11106,N_7044,N_7124);
xnor U11107 (N_11107,N_7791,N_7575);
and U11108 (N_11108,N_8499,N_8111);
and U11109 (N_11109,N_5028,N_7592);
or U11110 (N_11110,N_7748,N_6286);
nand U11111 (N_11111,N_7289,N_8161);
nor U11112 (N_11112,N_5845,N_7278);
xor U11113 (N_11113,N_7942,N_9171);
xnor U11114 (N_11114,N_9279,N_9188);
nor U11115 (N_11115,N_6807,N_7736);
xor U11116 (N_11116,N_9957,N_9131);
nand U11117 (N_11117,N_5817,N_9932);
nand U11118 (N_11118,N_5605,N_5769);
and U11119 (N_11119,N_6166,N_6351);
or U11120 (N_11120,N_9395,N_8960);
nand U11121 (N_11121,N_6418,N_8888);
nor U11122 (N_11122,N_5530,N_7567);
and U11123 (N_11123,N_5529,N_8376);
xor U11124 (N_11124,N_8662,N_6034);
or U11125 (N_11125,N_6450,N_8831);
xnor U11126 (N_11126,N_7972,N_8423);
nand U11127 (N_11127,N_9552,N_5714);
and U11128 (N_11128,N_8963,N_6967);
xnor U11129 (N_11129,N_8751,N_8092);
nor U11130 (N_11130,N_6601,N_9116);
and U11131 (N_11131,N_9408,N_6667);
or U11132 (N_11132,N_9810,N_9528);
and U11133 (N_11133,N_9352,N_9018);
and U11134 (N_11134,N_9360,N_8393);
and U11135 (N_11135,N_7915,N_8842);
and U11136 (N_11136,N_7855,N_5674);
or U11137 (N_11137,N_8594,N_8789);
or U11138 (N_11138,N_9497,N_5419);
nor U11139 (N_11139,N_9971,N_7015);
nand U11140 (N_11140,N_5432,N_9377);
nor U11141 (N_11141,N_6038,N_5265);
and U11142 (N_11142,N_5647,N_6081);
nor U11143 (N_11143,N_5991,N_7730);
and U11144 (N_11144,N_6465,N_6097);
and U11145 (N_11145,N_6485,N_6566);
and U11146 (N_11146,N_9237,N_9230);
nor U11147 (N_11147,N_6722,N_7704);
or U11148 (N_11148,N_9149,N_5999);
nor U11149 (N_11149,N_8474,N_7253);
or U11150 (N_11150,N_7402,N_7573);
nor U11151 (N_11151,N_7668,N_6168);
and U11152 (N_11152,N_7349,N_9735);
and U11153 (N_11153,N_6952,N_6863);
nor U11154 (N_11154,N_9654,N_7585);
nor U11155 (N_11155,N_5222,N_5576);
or U11156 (N_11156,N_7772,N_9632);
and U11157 (N_11157,N_6441,N_5749);
nor U11158 (N_11158,N_6857,N_8561);
nand U11159 (N_11159,N_7717,N_9265);
nand U11160 (N_11160,N_9926,N_8607);
xnor U11161 (N_11161,N_6085,N_8456);
nor U11162 (N_11162,N_8910,N_5371);
or U11163 (N_11163,N_7250,N_9234);
and U11164 (N_11164,N_9833,N_9056);
nand U11165 (N_11165,N_5663,N_8693);
nand U11166 (N_11166,N_6542,N_5507);
and U11167 (N_11167,N_6843,N_6860);
and U11168 (N_11168,N_9706,N_7808);
xnor U11169 (N_11169,N_9082,N_9959);
nand U11170 (N_11170,N_7862,N_8553);
and U11171 (N_11171,N_9470,N_5325);
xnor U11172 (N_11172,N_7225,N_9219);
or U11173 (N_11173,N_5987,N_8350);
xnor U11174 (N_11174,N_6826,N_9221);
nor U11175 (N_11175,N_5601,N_5840);
nand U11176 (N_11176,N_8913,N_8428);
nand U11177 (N_11177,N_8170,N_8049);
and U11178 (N_11178,N_5771,N_8652);
or U11179 (N_11179,N_6385,N_9085);
and U11180 (N_11180,N_7914,N_5404);
xnor U11181 (N_11181,N_7209,N_8698);
xnor U11182 (N_11182,N_5474,N_5528);
nand U11183 (N_11183,N_6987,N_5454);
or U11184 (N_11184,N_7012,N_8660);
xor U11185 (N_11185,N_9092,N_5701);
nand U11186 (N_11186,N_5108,N_8665);
nor U11187 (N_11187,N_5102,N_8883);
and U11188 (N_11188,N_7689,N_8314);
xnor U11189 (N_11189,N_6216,N_7543);
nor U11190 (N_11190,N_6511,N_8121);
and U11191 (N_11191,N_6998,N_5957);
xnor U11192 (N_11192,N_8168,N_9177);
nor U11193 (N_11193,N_6668,N_9879);
xnor U11194 (N_11194,N_5421,N_5244);
and U11195 (N_11195,N_7710,N_9369);
xnor U11196 (N_11196,N_6079,N_7148);
nor U11197 (N_11197,N_9513,N_8061);
or U11198 (N_11198,N_9938,N_8171);
nand U11199 (N_11199,N_5878,N_6761);
and U11200 (N_11200,N_9302,N_7917);
and U11201 (N_11201,N_8247,N_5895);
and U11202 (N_11202,N_7628,N_5959);
nor U11203 (N_11203,N_5409,N_6436);
nand U11204 (N_11204,N_5740,N_9576);
xor U11205 (N_11205,N_5563,N_7058);
or U11206 (N_11206,N_8283,N_7061);
nor U11207 (N_11207,N_6343,N_9045);
and U11208 (N_11208,N_8001,N_6532);
nand U11209 (N_11209,N_8580,N_6865);
nand U11210 (N_11210,N_9864,N_8995);
nor U11211 (N_11211,N_9662,N_8796);
and U11212 (N_11212,N_6768,N_5399);
nor U11213 (N_11213,N_6086,N_6358);
and U11214 (N_11214,N_9996,N_8984);
nand U11215 (N_11215,N_8864,N_6472);
and U11216 (N_11216,N_6769,N_5246);
and U11217 (N_11217,N_8050,N_6445);
or U11218 (N_11218,N_7282,N_5521);
nor U11219 (N_11219,N_6609,N_6811);
xor U11220 (N_11220,N_9548,N_7779);
nand U11221 (N_11221,N_9333,N_6677);
and U11222 (N_11222,N_7820,N_6434);
xor U11223 (N_11223,N_5083,N_6137);
nand U11224 (N_11224,N_6005,N_6623);
xnor U11225 (N_11225,N_5838,N_6169);
and U11226 (N_11226,N_8356,N_8634);
xnor U11227 (N_11227,N_8439,N_8900);
or U11228 (N_11228,N_8504,N_6267);
nor U11229 (N_11229,N_8438,N_6548);
xnor U11230 (N_11230,N_5788,N_6915);
xnor U11231 (N_11231,N_8136,N_8525);
nand U11232 (N_11232,N_5191,N_6234);
and U11233 (N_11233,N_6475,N_8291);
xnor U11234 (N_11234,N_7196,N_8529);
nand U11235 (N_11235,N_9294,N_8059);
or U11236 (N_11236,N_6526,N_6466);
xor U11237 (N_11237,N_8989,N_7902);
nor U11238 (N_11238,N_7338,N_5342);
and U11239 (N_11239,N_8044,N_6191);
xor U11240 (N_11240,N_7069,N_8949);
or U11241 (N_11241,N_5127,N_5326);
or U11242 (N_11242,N_6398,N_8637);
and U11243 (N_11243,N_7963,N_8166);
nand U11244 (N_11244,N_5646,N_8241);
or U11245 (N_11245,N_7591,N_7483);
nand U11246 (N_11246,N_8498,N_6720);
nand U11247 (N_11247,N_6125,N_9825);
nor U11248 (N_11248,N_7100,N_6837);
or U11249 (N_11249,N_9544,N_9807);
nand U11250 (N_11250,N_7275,N_6322);
xnor U11251 (N_11251,N_6217,N_7458);
xnor U11252 (N_11252,N_6292,N_8176);
or U11253 (N_11253,N_8123,N_6041);
nand U11254 (N_11254,N_9325,N_9067);
or U11255 (N_11255,N_5331,N_6590);
xnor U11256 (N_11256,N_5711,N_5205);
xor U11257 (N_11257,N_9746,N_5721);
xor U11258 (N_11258,N_5864,N_9227);
xnor U11259 (N_11259,N_6307,N_7993);
xnor U11260 (N_11260,N_7931,N_9334);
nand U11261 (N_11261,N_5096,N_9726);
or U11262 (N_11262,N_8759,N_9181);
and U11263 (N_11263,N_5017,N_9044);
xnor U11264 (N_11264,N_9434,N_5170);
nor U11265 (N_11265,N_8985,N_9453);
nand U11266 (N_11266,N_7356,N_6152);
xnor U11267 (N_11267,N_5770,N_9561);
and U11268 (N_11268,N_5499,N_9161);
xnor U11269 (N_11269,N_9589,N_5089);
or U11270 (N_11270,N_5403,N_6701);
nor U11271 (N_11271,N_6620,N_9284);
and U11272 (N_11272,N_9827,N_8093);
and U11273 (N_11273,N_8611,N_8334);
nand U11274 (N_11274,N_7226,N_9123);
nand U11275 (N_11275,N_7455,N_5879);
or U11276 (N_11276,N_7445,N_9562);
nand U11277 (N_11277,N_6156,N_9309);
and U11278 (N_11278,N_5780,N_7131);
nor U11279 (N_11279,N_9023,N_5614);
and U11280 (N_11280,N_9861,N_7478);
and U11281 (N_11281,N_6296,N_6831);
or U11282 (N_11282,N_8120,N_9190);
xnor U11283 (N_11283,N_9695,N_7792);
nand U11284 (N_11284,N_8572,N_5729);
nor U11285 (N_11285,N_5992,N_6071);
xnor U11286 (N_11286,N_5609,N_7554);
or U11287 (N_11287,N_8851,N_7305);
and U11288 (N_11288,N_8038,N_8530);
nor U11289 (N_11289,N_5248,N_6707);
or U11290 (N_11290,N_7323,N_7474);
and U11291 (N_11291,N_6314,N_5642);
and U11292 (N_11292,N_9311,N_6916);
or U11293 (N_11293,N_9077,N_7750);
nand U11294 (N_11294,N_7363,N_6128);
nand U11295 (N_11295,N_9321,N_6920);
nor U11296 (N_11296,N_6940,N_7489);
nor U11297 (N_11297,N_7650,N_6375);
nand U11298 (N_11298,N_5431,N_6962);
xnor U11299 (N_11299,N_6340,N_5294);
nor U11300 (N_11300,N_6287,N_9477);
nor U11301 (N_11301,N_5375,N_5126);
nor U11302 (N_11302,N_8929,N_8890);
or U11303 (N_11303,N_6244,N_9856);
nor U11304 (N_11304,N_9892,N_9240);
and U11305 (N_11305,N_8215,N_8402);
or U11306 (N_11306,N_6408,N_8180);
xor U11307 (N_11307,N_8631,N_8274);
xnor U11308 (N_11308,N_9076,N_8757);
nand U11309 (N_11309,N_8916,N_6280);
nor U11310 (N_11310,N_6049,N_9464);
nand U11311 (N_11311,N_8819,N_8394);
nor U11312 (N_11312,N_5193,N_7065);
nand U11313 (N_11313,N_7929,N_8959);
xnor U11314 (N_11314,N_9417,N_5235);
xor U11315 (N_11315,N_7946,N_6556);
xor U11316 (N_11316,N_9975,N_8803);
nor U11317 (N_11317,N_7806,N_8968);
nand U11318 (N_11318,N_6454,N_7296);
and U11319 (N_11319,N_5299,N_9637);
xor U11320 (N_11320,N_7524,N_7768);
and U11321 (N_11321,N_8735,N_6844);
and U11322 (N_11322,N_5930,N_9766);
and U11323 (N_11323,N_9579,N_8186);
or U11324 (N_11324,N_6367,N_7276);
xnor U11325 (N_11325,N_9473,N_5485);
xnor U11326 (N_11326,N_8298,N_5226);
or U11327 (N_11327,N_5372,N_8922);
or U11328 (N_11328,N_9432,N_6990);
or U11329 (N_11329,N_7198,N_9922);
nand U11330 (N_11330,N_8466,N_5049);
and U11331 (N_11331,N_7934,N_8697);
and U11332 (N_11332,N_6062,N_8302);
xor U11333 (N_11333,N_7484,N_6011);
xor U11334 (N_11334,N_6607,N_6780);
or U11335 (N_11335,N_7248,N_7388);
nor U11336 (N_11336,N_6717,N_9350);
or U11337 (N_11337,N_6313,N_5054);
nand U11338 (N_11338,N_7203,N_5896);
and U11339 (N_11339,N_6012,N_8604);
nand U11340 (N_11340,N_8540,N_5777);
nor U11341 (N_11341,N_6355,N_9646);
or U11342 (N_11342,N_6650,N_6078);
and U11343 (N_11343,N_7104,N_7187);
or U11344 (N_11344,N_8289,N_7550);
xnor U11345 (N_11345,N_9511,N_9794);
nor U11346 (N_11346,N_8987,N_6219);
and U11347 (N_11347,N_6691,N_9422);
nor U11348 (N_11348,N_7905,N_8901);
or U11349 (N_11349,N_6241,N_6928);
and U11350 (N_11350,N_9142,N_7523);
or U11351 (N_11351,N_5904,N_9187);
or U11352 (N_11352,N_7060,N_5982);
xor U11353 (N_11353,N_9914,N_9560);
nor U11354 (N_11354,N_9442,N_9308);
nor U11355 (N_11355,N_5239,N_9281);
or U11356 (N_11356,N_5712,N_7686);
xor U11357 (N_11357,N_7092,N_9586);
and U11358 (N_11358,N_7381,N_6981);
nand U11359 (N_11359,N_6483,N_7908);
and U11360 (N_11360,N_7659,N_8282);
nand U11361 (N_11361,N_8977,N_9613);
nor U11362 (N_11362,N_6563,N_5510);
and U11363 (N_11363,N_6821,N_9663);
nor U11364 (N_11364,N_8398,N_5775);
nor U11365 (N_11365,N_9071,N_8980);
nand U11366 (N_11366,N_7742,N_9692);
nor U11367 (N_11367,N_6433,N_6026);
and U11368 (N_11368,N_8746,N_6755);
or U11369 (N_11369,N_7382,N_8710);
xnor U11370 (N_11370,N_5612,N_9747);
nand U11371 (N_11371,N_5429,N_9213);
xor U11372 (N_11372,N_7560,N_7756);
and U11373 (N_11373,N_8246,N_5183);
or U11374 (N_11374,N_8147,N_6312);
and U11375 (N_11375,N_9241,N_7949);
or U11376 (N_11376,N_5339,N_8887);
xor U11377 (N_11377,N_8969,N_9603);
or U11378 (N_11378,N_6881,N_5081);
or U11379 (N_11379,N_5428,N_8573);
and U11380 (N_11380,N_7079,N_5548);
and U11381 (N_11381,N_8996,N_7453);
or U11382 (N_11382,N_9065,N_8141);
xor U11383 (N_11383,N_6599,N_7876);
nand U11384 (N_11384,N_8307,N_7913);
xor U11385 (N_11385,N_9274,N_8723);
nand U11386 (N_11386,N_8635,N_5426);
xnor U11387 (N_11387,N_7794,N_7467);
and U11388 (N_11388,N_9207,N_6572);
nand U11389 (N_11389,N_9908,N_5808);
nor U11390 (N_11390,N_6719,N_8867);
nand U11391 (N_11391,N_8262,N_9950);
or U11392 (N_11392,N_5611,N_8041);
xnor U11393 (N_11393,N_5157,N_5844);
and U11394 (N_11394,N_5129,N_7094);
and U11395 (N_11395,N_6727,N_7273);
or U11396 (N_11396,N_9439,N_5968);
nor U11397 (N_11397,N_8632,N_6737);
xnor U11398 (N_11398,N_7919,N_8366);
or U11399 (N_11399,N_8399,N_8406);
xor U11400 (N_11400,N_5915,N_7335);
xor U11401 (N_11401,N_7471,N_5690);
and U11402 (N_11402,N_6430,N_6403);
nand U11403 (N_11403,N_7259,N_9481);
nand U11404 (N_11404,N_8624,N_7186);
xor U11405 (N_11405,N_8015,N_8736);
or U11406 (N_11406,N_5652,N_5779);
and U11407 (N_11407,N_9563,N_7932);
nor U11408 (N_11408,N_6856,N_7631);
or U11409 (N_11409,N_6316,N_7923);
nor U11410 (N_11410,N_7504,N_5503);
or U11411 (N_11411,N_9697,N_5739);
and U11412 (N_11412,N_9425,N_8998);
or U11413 (N_11413,N_6455,N_8845);
xor U11414 (N_11414,N_5859,N_6082);
nor U11415 (N_11415,N_5438,N_5705);
nor U11416 (N_11416,N_5452,N_9641);
nor U11417 (N_11417,N_6039,N_6171);
xor U11418 (N_11418,N_5442,N_5698);
xnor U11419 (N_11419,N_6783,N_8893);
nand U11420 (N_11420,N_8287,N_5990);
nor U11421 (N_11421,N_8879,N_8346);
nand U11422 (N_11422,N_8961,N_5725);
or U11423 (N_11423,N_7154,N_5099);
or U11424 (N_11424,N_5931,N_7911);
and U11425 (N_11425,N_6235,N_5098);
and U11426 (N_11426,N_5887,N_7143);
nand U11427 (N_11427,N_6029,N_9707);
or U11428 (N_11428,N_8596,N_9411);
nand U11429 (N_11429,N_5249,N_6884);
xor U11430 (N_11430,N_5021,N_8791);
and U11431 (N_11431,N_7707,N_9625);
xor U11432 (N_11432,N_7077,N_8087);
and U11433 (N_11433,N_6746,N_6261);
and U11434 (N_11434,N_9951,N_7957);
nand U11435 (N_11435,N_6040,N_8579);
or U11436 (N_11436,N_9838,N_7267);
and U11437 (N_11437,N_5809,N_9688);
or U11438 (N_11438,N_5933,N_8116);
nand U11439 (N_11439,N_7136,N_6000);
and U11440 (N_11440,N_9567,N_7372);
nor U11441 (N_11441,N_6284,N_5451);
xor U11442 (N_11442,N_6994,N_6827);
nand U11443 (N_11443,N_8113,N_8920);
or U11444 (N_11444,N_6938,N_5888);
or U11445 (N_11445,N_9362,N_5434);
and U11446 (N_11446,N_7903,N_5687);
or U11447 (N_11447,N_5417,N_9178);
or U11448 (N_11448,N_8747,N_8595);
or U11449 (N_11449,N_5662,N_9060);
nand U11450 (N_11450,N_8638,N_9891);
nor U11451 (N_11451,N_8480,N_9108);
xor U11452 (N_11452,N_9661,N_8714);
and U11453 (N_11453,N_8908,N_7059);
nand U11454 (N_11454,N_7039,N_9534);
nand U11455 (N_11455,N_6407,N_6652);
and U11456 (N_11456,N_8776,N_8823);
xor U11457 (N_11457,N_7766,N_7204);
or U11458 (N_11458,N_9438,N_9029);
or U11459 (N_11459,N_7266,N_9797);
nand U11460 (N_11460,N_7526,N_5117);
xnor U11461 (N_11461,N_9298,N_5133);
and U11462 (N_11462,N_7031,N_7943);
nor U11463 (N_11463,N_9551,N_9105);
and U11464 (N_11464,N_9873,N_6232);
and U11465 (N_11465,N_5776,N_9575);
nor U11466 (N_11466,N_6859,N_7965);
or U11467 (N_11467,N_7157,N_9792);
and U11468 (N_11468,N_6630,N_7195);
and U11469 (N_11469,N_8419,N_5175);
nand U11470 (N_11470,N_5439,N_8117);
and U11471 (N_11471,N_9250,N_6937);
xnor U11472 (N_11472,N_9493,N_6800);
xor U11473 (N_11473,N_9680,N_7620);
or U11474 (N_11474,N_7522,N_6279);
and U11475 (N_11475,N_5343,N_5180);
nand U11476 (N_11476,N_5800,N_8292);
or U11477 (N_11477,N_6017,N_7610);
and U11478 (N_11478,N_8863,N_7799);
and U11479 (N_11479,N_6326,N_8547);
and U11480 (N_11480,N_8848,N_5400);
xor U11481 (N_11481,N_7529,N_7755);
nor U11482 (N_11482,N_5159,N_6852);
nand U11483 (N_11483,N_7705,N_6522);
or U11484 (N_11484,N_8649,N_8597);
or U11485 (N_11485,N_8203,N_9503);
xor U11486 (N_11486,N_5972,N_5391);
xnor U11487 (N_11487,N_9452,N_7861);
nand U11488 (N_11488,N_8853,N_8844);
and U11489 (N_11489,N_5812,N_6518);
nor U11490 (N_11490,N_7625,N_7013);
and U11491 (N_11491,N_9338,N_7452);
nor U11492 (N_11492,N_6693,N_7877);
nand U11493 (N_11493,N_7002,N_7990);
and U11494 (N_11494,N_7759,N_8716);
or U11495 (N_11495,N_6714,N_8769);
xor U11496 (N_11496,N_5924,N_6157);
nand U11497 (N_11497,N_7838,N_7490);
and U11498 (N_11498,N_6400,N_7139);
nor U11499 (N_11499,N_9902,N_8623);
xor U11500 (N_11500,N_7510,N_8777);
and U11501 (N_11501,N_7156,N_8966);
or U11502 (N_11502,N_6997,N_6184);
nand U11503 (N_11503,N_7804,N_8200);
or U11504 (N_11504,N_9256,N_5998);
or U11505 (N_11505,N_6686,N_7185);
nand U11506 (N_11506,N_5918,N_6132);
nand U11507 (N_11507,N_7214,N_5097);
and U11508 (N_11508,N_8259,N_7232);
and U11509 (N_11509,N_5364,N_7068);
xnor U11510 (N_11510,N_9478,N_9667);
nor U11511 (N_11511,N_6114,N_7390);
or U11512 (N_11512,N_6065,N_6977);
and U11513 (N_11513,N_5790,N_9055);
nor U11514 (N_11514,N_6947,N_9148);
nand U11515 (N_11515,N_8424,N_8836);
or U11516 (N_11516,N_6577,N_9134);
nor U11517 (N_11517,N_5204,N_9062);
or U11518 (N_11518,N_7046,N_7488);
nand U11519 (N_11519,N_6158,N_8258);
nand U11520 (N_11520,N_9027,N_7081);
nand U11521 (N_11521,N_5828,N_9145);
xnor U11522 (N_11522,N_8849,N_9329);
nand U11523 (N_11523,N_6463,N_9479);
xor U11524 (N_11524,N_7646,N_9580);
nor U11525 (N_11525,N_7896,N_7947);
and U11526 (N_11526,N_6868,N_9392);
nor U11527 (N_11527,N_6238,N_5549);
or U11528 (N_11528,N_6638,N_7412);
nand U11529 (N_11529,N_9690,N_7561);
or U11530 (N_11530,N_9409,N_8470);
xor U11531 (N_11531,N_5047,N_5746);
and U11532 (N_11532,N_8112,N_9805);
or U11533 (N_11533,N_5348,N_9289);
and U11534 (N_11534,N_6943,N_7384);
xor U11535 (N_11535,N_8609,N_7571);
nor U11536 (N_11536,N_9262,N_5868);
nand U11537 (N_11537,N_5322,N_8923);
nor U11538 (N_11538,N_5656,N_5475);
xnor U11539 (N_11539,N_6689,N_8669);
nor U11540 (N_11540,N_9328,N_5821);
nand U11541 (N_11541,N_6968,N_8615);
nor U11542 (N_11542,N_8780,N_5154);
nor U11543 (N_11543,N_9064,N_5063);
or U11544 (N_11544,N_6756,N_5360);
nand U11545 (N_11545,N_8784,N_6622);
and U11546 (N_11546,N_7624,N_5635);
or U11547 (N_11547,N_6871,N_8494);
xnor U11548 (N_11548,N_6569,N_5153);
nand U11549 (N_11549,N_5723,N_5281);
nor U11550 (N_11550,N_8554,N_8955);
or U11551 (N_11551,N_7565,N_7540);
and U11552 (N_11552,N_6695,N_8078);
xnor U11553 (N_11553,N_9572,N_9634);
or U11554 (N_11554,N_9224,N_8535);
nand U11555 (N_11555,N_7408,N_6146);
nor U11556 (N_11556,N_7417,N_7712);
nor U11557 (N_11557,N_8024,N_8874);
and U11558 (N_11558,N_5192,N_9743);
or U11559 (N_11559,N_5072,N_6380);
and U11560 (N_11560,N_9474,N_7549);
nor U11561 (N_11561,N_5470,N_7633);
xor U11562 (N_11562,N_9355,N_9558);
xnor U11563 (N_11563,N_7129,N_6626);
and U11564 (N_11564,N_6336,N_9460);
nand U11565 (N_11565,N_9550,N_7864);
and U11566 (N_11566,N_5137,N_8538);
or U11567 (N_11567,N_9530,N_7354);
or U11568 (N_11568,N_7298,N_9272);
or U11569 (N_11569,N_5795,N_5002);
and U11570 (N_11570,N_6270,N_6625);
and U11571 (N_11571,N_5497,N_5960);
nor U11572 (N_11572,N_7873,N_5155);
and U11573 (N_11573,N_5194,N_9587);
nor U11574 (N_11574,N_5765,N_8272);
nor U11575 (N_11575,N_6978,N_8369);
nor U11576 (N_11576,N_7667,N_8273);
or U11577 (N_11577,N_7691,N_9115);
nor U11578 (N_11578,N_9292,N_7516);
or U11579 (N_11579,N_5075,N_5481);
and U11580 (N_11580,N_6315,N_9314);
and U11581 (N_11581,N_7017,N_7392);
or U11582 (N_11582,N_5460,N_7867);
xor U11583 (N_11583,N_8271,N_9607);
nand U11584 (N_11584,N_9615,N_9970);
nand U11585 (N_11585,N_9006,N_6113);
and U11586 (N_11586,N_9814,N_5708);
or U11587 (N_11587,N_8370,N_8917);
and U11588 (N_11588,N_7769,N_6246);
nand U11589 (N_11589,N_7753,N_6961);
and U11590 (N_11590,N_9834,N_7813);
nand U11591 (N_11591,N_7557,N_8245);
and U11592 (N_11592,N_9388,N_7661);
nor U11593 (N_11593,N_8193,N_7521);
xor U11594 (N_11594,N_7537,N_5811);
nor U11595 (N_11595,N_6328,N_5045);
xnor U11596 (N_11596,N_5128,N_8793);
or U11597 (N_11597,N_7010,N_8810);
and U11598 (N_11598,N_8221,N_7775);
nor U11599 (N_11599,N_8485,N_8448);
nand U11600 (N_11600,N_6419,N_7928);
or U11601 (N_11601,N_5323,N_6010);
and U11602 (N_11602,N_6480,N_5717);
and U11603 (N_11603,N_8725,N_5367);
and U11604 (N_11604,N_8294,N_6529);
nor U11605 (N_11605,N_9340,N_6818);
or U11606 (N_11606,N_6973,N_6088);
and U11607 (N_11607,N_7431,N_9650);
nor U11608 (N_11608,N_8881,N_8566);
and U11609 (N_11609,N_7223,N_7830);
xor U11610 (N_11610,N_9952,N_6420);
nor U11611 (N_11611,N_8306,N_9723);
nor U11612 (N_11612,N_9981,N_9507);
nand U11613 (N_11613,N_8371,N_6369);
nor U11614 (N_11614,N_5975,N_8315);
and U11615 (N_11615,N_5356,N_9531);
nor U11616 (N_11616,N_8458,N_8728);
or U11617 (N_11617,N_8767,N_7870);
nand U11618 (N_11618,N_6167,N_5345);
xor U11619 (N_11619,N_7506,N_8644);
and U11620 (N_11620,N_6713,N_5062);
nand U11621 (N_11621,N_6593,N_6383);
and U11622 (N_11622,N_6045,N_5835);
and U11623 (N_11623,N_8678,N_8619);
xnor U11624 (N_11624,N_8165,N_7688);
or U11625 (N_11625,N_8562,N_8451);
nor U11626 (N_11626,N_8613,N_6538);
xnor U11627 (N_11627,N_8441,N_8990);
nand U11628 (N_11628,N_5831,N_8158);
and U11629 (N_11629,N_6151,N_6621);
nor U11630 (N_11630,N_5486,N_8027);
nand U11631 (N_11631,N_7222,N_8674);
and U11632 (N_11632,N_7240,N_5752);
nor U11633 (N_11633,N_6787,N_6257);
and U11634 (N_11634,N_7921,N_5716);
nor U11635 (N_11635,N_9446,N_6642);
or U11636 (N_11636,N_5592,N_5278);
and U11637 (N_11637,N_5327,N_9642);
nor U11638 (N_11638,N_5056,N_7247);
and U11639 (N_11639,N_5055,N_7395);
or U11640 (N_11640,N_9239,N_8935);
nand U11641 (N_11641,N_9983,N_9913);
nand U11642 (N_11642,N_6360,N_5412);
and U11643 (N_11643,N_8022,N_6437);
nand U11644 (N_11644,N_6815,N_5190);
xor U11645 (N_11645,N_9699,N_5949);
xor U11646 (N_11646,N_8981,N_9962);
xnor U11647 (N_11647,N_8380,N_6718);
or U11648 (N_11648,N_7836,N_7086);
and U11649 (N_11649,N_6186,N_7049);
nand U11650 (N_11650,N_7648,N_6447);
nand U11651 (N_11651,N_6991,N_7890);
nand U11652 (N_11652,N_7980,N_8930);
xor U11653 (N_11653,N_5494,N_8628);
nor U11654 (N_11654,N_6344,N_6585);
xnor U11655 (N_11655,N_8137,N_7072);
or U11656 (N_11656,N_5734,N_5571);
nand U11657 (N_11657,N_9649,N_5051);
or U11658 (N_11658,N_5425,N_9205);
nand U11659 (N_11659,N_8065,N_7228);
or U11660 (N_11660,N_9937,N_6022);
nand U11661 (N_11661,N_5802,N_9235);
or U11662 (N_11662,N_5290,N_8685);
nor U11663 (N_11663,N_5297,N_6716);
nand U11664 (N_11664,N_9454,N_8299);
or U11665 (N_11665,N_8226,N_9319);
and U11666 (N_11666,N_6288,N_9075);
xnor U11667 (N_11667,N_6333,N_6268);
nand U11668 (N_11668,N_9450,N_8188);
or U11669 (N_11669,N_8585,N_8717);
nor U11670 (N_11670,N_9244,N_8172);
or U11671 (N_11671,N_5311,N_5603);
nand U11672 (N_11672,N_5176,N_6882);
or U11673 (N_11673,N_9754,N_6632);
or U11674 (N_11674,N_6838,N_8446);
xor U11675 (N_11675,N_7544,N_5023);
nor U11676 (N_11676,N_7652,N_8896);
and U11677 (N_11677,N_7485,N_9192);
xor U11678 (N_11678,N_7470,N_6694);
nor U11679 (N_11679,N_7832,N_9823);
or U11680 (N_11680,N_6841,N_5798);
and U11681 (N_11681,N_7721,N_6006);
and U11682 (N_11682,N_5621,N_8156);
nor U11683 (N_11683,N_7095,N_9072);
nand U11684 (N_11684,N_5873,N_8640);
xnor U11685 (N_11685,N_5894,N_5216);
nor U11686 (N_11686,N_9624,N_8195);
or U11687 (N_11687,N_5185,N_8951);
and U11688 (N_11688,N_7925,N_9266);
xnor U11689 (N_11689,N_9335,N_9223);
nor U11690 (N_11690,N_9751,N_5751);
nand U11691 (N_11691,N_8534,N_7181);
nand U11692 (N_11692,N_7773,N_7978);
and U11693 (N_11693,N_9860,N_5255);
and U11694 (N_11694,N_9705,N_6697);
nor U11695 (N_11695,N_6129,N_7811);
or U11696 (N_11696,N_5466,N_6345);
and U11697 (N_11697,N_5870,N_8719);
xnor U11698 (N_11698,N_7443,N_6531);
nor U11699 (N_11699,N_5772,N_7482);
nor U11700 (N_11700,N_9730,N_7377);
and U11701 (N_11701,N_6133,N_7168);
nand U11702 (N_11702,N_7254,N_5905);
nor U11703 (N_11703,N_8800,N_8629);
nor U11704 (N_11704,N_9043,N_8774);
nand U11705 (N_11705,N_8095,N_7656);
nand U11706 (N_11706,N_8794,N_9519);
nor U11707 (N_11707,N_9394,N_6864);
or U11708 (N_11708,N_5584,N_9010);
nor U11709 (N_11709,N_5602,N_8655);
and U11710 (N_11710,N_9564,N_6391);
xnor U11711 (N_11711,N_7366,N_8150);
nand U11712 (N_11712,N_9068,N_5846);
and U11713 (N_11713,N_9808,N_6999);
nor U11714 (N_11714,N_9121,N_6324);
nand U11715 (N_11715,N_7437,N_7564);
and U11716 (N_11716,N_5435,N_5241);
or U11717 (N_11717,N_7869,N_8420);
nand U11718 (N_11718,N_6945,N_8688);
xor U11719 (N_11719,N_8336,N_9243);
nand U11720 (N_11720,N_7167,N_6469);
nor U11721 (N_11721,N_8285,N_5737);
nor U11722 (N_11722,N_6285,N_8876);
xnor U11723 (N_11723,N_5388,N_8520);
and U11724 (N_11724,N_6796,N_7473);
xnor U11725 (N_11725,N_5545,N_8857);
nor U11726 (N_11726,N_5217,N_5983);
nand U11727 (N_11727,N_6397,N_9961);
nor U11728 (N_11728,N_5293,N_6992);
xor U11729 (N_11729,N_9367,N_9502);
and U11730 (N_11730,N_7778,N_6786);
and U11731 (N_11731,N_7627,N_7724);
nor U11732 (N_11732,N_5328,N_5514);
and U11733 (N_11733,N_5523,N_6670);
and U11734 (N_11734,N_5139,N_8145);
nor U11735 (N_11735,N_6798,N_5950);
or U11736 (N_11736,N_9037,N_9229);
or U11737 (N_11737,N_7679,N_7910);
nor U11738 (N_11738,N_8687,N_5557);
or U11739 (N_11739,N_8357,N_5847);
nor U11740 (N_11740,N_8225,N_8144);
and U11741 (N_11741,N_6075,N_6982);
nor U11742 (N_11742,N_8257,N_5623);
xor U11743 (N_11743,N_7292,N_6861);
and U11744 (N_11744,N_6971,N_8993);
and U11745 (N_11745,N_9248,N_5259);
nor U11746 (N_11746,N_8253,N_5632);
nor U11747 (N_11747,N_9555,N_9447);
nand U11748 (N_11748,N_7764,N_5515);
and U11749 (N_11749,N_6066,N_8673);
or U11750 (N_11750,N_8378,N_8139);
xnor U11751 (N_11751,N_8880,N_8085);
and U11752 (N_11752,N_5110,N_9711);
or U11753 (N_11753,N_6853,N_8650);
nor U11754 (N_11754,N_7120,N_8870);
and U11755 (N_11755,N_9154,N_7840);
nand U11756 (N_11756,N_6204,N_9363);
xor U11757 (N_11757,N_9964,N_8075);
and U11758 (N_11758,N_8545,N_8233);
nor U11759 (N_11759,N_5455,N_9907);
xnor U11760 (N_11760,N_8740,N_8125);
and U11761 (N_11761,N_6892,N_7912);
nand U11762 (N_11762,N_9545,N_7284);
nand U11763 (N_11763,N_5448,N_5309);
nand U11764 (N_11764,N_6570,N_5123);
and U11765 (N_11765,N_5464,N_7556);
nor U11766 (N_11766,N_9260,N_7991);
nor U11767 (N_11767,N_8643,N_9100);
xor U11768 (N_11768,N_9080,N_7641);
and U11769 (N_11769,N_8373,N_7343);
or U11770 (N_11770,N_5595,N_6743);
xnor U11771 (N_11771,N_7555,N_7872);
nand U11772 (N_11772,N_5692,N_7545);
xor U11773 (N_11773,N_8488,N_6163);
or U11774 (N_11774,N_9783,N_7150);
xor U11775 (N_11775,N_8084,N_9135);
or U11776 (N_11776,N_6876,N_5989);
nand U11777 (N_11777,N_6337,N_9518);
and U11778 (N_11778,N_7325,N_7301);
or U11779 (N_11779,N_7868,N_9472);
xnor U11780 (N_11780,N_7035,N_5564);
xor U11781 (N_11781,N_8071,N_7626);
nor U11782 (N_11782,N_7098,N_9724);
or U11783 (N_11783,N_5197,N_8224);
xnor U11784 (N_11784,N_8301,N_6237);
nand U11785 (N_11785,N_8270,N_6068);
or U11786 (N_11786,N_7355,N_5352);
xor U11787 (N_11787,N_6352,N_7425);
and U11788 (N_11788,N_8830,N_6752);
nand U11789 (N_11789,N_5042,N_6247);
and U11790 (N_11790,N_8312,N_9984);
nand U11791 (N_11791,N_9291,N_9948);
and U11792 (N_11792,N_8667,N_5882);
xor U11793 (N_11793,N_9236,N_8218);
or U11794 (N_11794,N_7760,N_7959);
nor U11795 (N_11795,N_9090,N_8361);
or U11796 (N_11796,N_9195,N_9225);
or U11797 (N_11797,N_6188,N_6056);
nand U11798 (N_11798,N_8860,N_9911);
nor U11799 (N_11799,N_5468,N_6201);
and U11800 (N_11800,N_7123,N_8682);
xnor U11801 (N_11801,N_5685,N_9249);
xor U11802 (N_11802,N_8037,N_8462);
nand U11803 (N_11803,N_5167,N_6124);
xnor U11804 (N_11804,N_8360,N_6321);
nand U11805 (N_11805,N_6512,N_7464);
xnor U11806 (N_11806,N_5901,N_7271);
and U11807 (N_11807,N_6104,N_8921);
or U11808 (N_11808,N_7899,N_7033);
nor U11809 (N_11809,N_9444,N_9842);
or U11810 (N_11810,N_9896,N_8790);
or U11811 (N_11811,N_6839,N_6093);
or U11812 (N_11812,N_7469,N_5030);
and U11813 (N_11813,N_9303,N_9461);
nand U11814 (N_11814,N_9401,N_6063);
xor U11815 (N_11815,N_5997,N_5415);
and U11816 (N_11816,N_9782,N_5956);
and U11817 (N_11817,N_5572,N_6929);
or U11818 (N_11818,N_7548,N_8486);
xor U11819 (N_11819,N_5261,N_6612);
or U11820 (N_11820,N_6589,N_6870);
xor U11821 (N_11821,N_9800,N_5748);
or U11822 (N_11822,N_8686,N_9185);
xor U11823 (N_11823,N_9320,N_5161);
or U11824 (N_11824,N_5710,N_9341);
or U11825 (N_11825,N_6226,N_9693);
nor U11826 (N_11826,N_8388,N_7353);
nor U11827 (N_11827,N_6021,N_8928);
xor U11828 (N_11828,N_5538,N_9698);
nor U11829 (N_11829,N_7999,N_5567);
nand U11830 (N_11830,N_6446,N_6362);
nand U11831 (N_11831,N_8648,N_6931);
nor U11832 (N_11832,N_6495,N_5819);
xor U11833 (N_11833,N_5362,N_8083);
nand U11834 (N_11834,N_8633,N_9876);
nand U11835 (N_11835,N_7530,N_9033);
xor U11836 (N_11836,N_7191,N_6936);
nor U11837 (N_11837,N_9489,N_8555);
xnor U11838 (N_11838,N_9078,N_9098);
xnor U11839 (N_11839,N_5178,N_9117);
and U11840 (N_11840,N_5902,N_9874);
or U11841 (N_11841,N_9421,N_6401);
and U11842 (N_11842,N_7210,N_5087);
nor U11843 (N_11843,N_7711,N_6335);
nand U11844 (N_11844,N_7843,N_6153);
xnor U11845 (N_11845,N_6930,N_8764);
nor U11846 (N_11846,N_9989,N_6373);
nand U11847 (N_11847,N_6665,N_7900);
nor U11848 (N_11848,N_6160,N_8005);
nor U11849 (N_11849,N_6706,N_5625);
nand U11850 (N_11850,N_7105,N_9183);
xor U11851 (N_11851,N_8937,N_7462);
xor U11852 (N_11852,N_8054,N_9091);
xnor U11853 (N_11853,N_8367,N_8377);
xnor U11854 (N_11854,N_7493,N_9386);
nor U11855 (N_11855,N_5160,N_6311);
and U11856 (N_11856,N_9110,N_8979);
and U11857 (N_11857,N_5505,N_6513);
and U11858 (N_11858,N_5671,N_5288);
nor U11859 (N_11859,N_7110,N_8349);
or U11860 (N_11860,N_7155,N_5303);
and U11861 (N_11861,N_9404,N_5498);
xor U11862 (N_11862,N_8417,N_8062);
xor U11863 (N_11863,N_7380,N_9935);
xor U11864 (N_11864,N_5754,N_7097);
or U11865 (N_11865,N_7487,N_7414);
or U11866 (N_11866,N_6552,N_8368);
or U11867 (N_11867,N_7800,N_7003);
nor U11868 (N_11868,N_5236,N_8734);
xnor U11869 (N_11869,N_5076,N_7177);
and U11870 (N_11870,N_9906,N_7783);
or U11871 (N_11871,N_6854,N_6435);
nand U11872 (N_11872,N_8070,N_8069);
xor U11873 (N_11873,N_9346,N_7505);
or U11874 (N_11874,N_8889,N_6704);
nand U11875 (N_11875,N_7574,N_9788);
nand U11876 (N_11876,N_7368,N_8541);
xnor U11877 (N_11877,N_6883,N_7827);
nor U11878 (N_11878,N_5365,N_6126);
nor U11879 (N_11879,N_8408,N_7645);
nor U11880 (N_11880,N_9153,N_9750);
nor U11881 (N_11881,N_6774,N_7235);
nor U11882 (N_11882,N_9079,N_9909);
nand U11883 (N_11883,N_8469,N_9139);
or U11884 (N_11884,N_6918,N_7559);
or U11885 (N_11885,N_9007,N_6748);
or U11886 (N_11886,N_7260,N_9982);
nand U11887 (N_11887,N_8431,N_6797);
nor U11888 (N_11888,N_5683,N_7304);
nand U11889 (N_11889,N_5029,N_6682);
nor U11890 (N_11890,N_6094,N_5138);
nor U11891 (N_11891,N_9944,N_5103);
nand U11892 (N_11892,N_8683,N_8907);
nor U11893 (N_11893,N_8715,N_5286);
or U11894 (N_11894,N_8808,N_6560);
xor U11895 (N_11895,N_9463,N_5156);
or U11896 (N_11896,N_9772,N_6959);
nand U11897 (N_11897,N_7590,N_9212);
xor U11898 (N_11898,N_5824,N_8454);
or U11899 (N_11899,N_5149,N_9802);
xnor U11900 (N_11900,N_5406,N_9180);
nand U11901 (N_11901,N_9685,N_5135);
nand U11902 (N_11902,N_9138,N_6584);
or U11903 (N_11903,N_7023,N_9456);
nand U11904 (N_11904,N_7584,N_5179);
or U11905 (N_11905,N_8478,N_9538);
nor U11906 (N_11906,N_6855,N_5898);
nor U11907 (N_11907,N_6934,N_8512);
and U11908 (N_11908,N_9222,N_8099);
or U11909 (N_11909,N_8942,N_8508);
xor U11910 (N_11910,N_9818,N_8389);
or U11911 (N_11911,N_5120,N_8148);
or U11912 (N_11912,N_8052,N_8058);
nor U11913 (N_11913,N_8575,N_5559);
nor U11914 (N_11914,N_5596,N_6750);
nand U11915 (N_11915,N_9508,N_7809);
nand U11916 (N_11916,N_7642,N_5792);
nor U11917 (N_11917,N_9264,N_9740);
xnor U11918 (N_11918,N_9670,N_7435);
or U11919 (N_11919,N_6392,N_6603);
or U11920 (N_11920,N_8657,N_7552);
or U11921 (N_11921,N_9767,N_6541);
nor U11922 (N_11922,N_6785,N_7535);
nor U11923 (N_11923,N_6806,N_5341);
nor U11924 (N_11924,N_6680,N_7438);
xor U11925 (N_11925,N_7428,N_5786);
xnor U11926 (N_11926,N_6900,N_8550);
or U11927 (N_11927,N_7344,N_9980);
or U11928 (N_11928,N_9039,N_9826);
and U11929 (N_11929,N_7977,N_9179);
nor U11930 (N_11930,N_7229,N_7227);
xnor U11931 (N_11931,N_7936,N_5970);
nor U11932 (N_11932,N_9370,N_9583);
or U11933 (N_11933,N_9254,N_9999);
and U11934 (N_11934,N_5758,N_5858);
xnor U11935 (N_11935,N_5837,N_7513);
xnor U11936 (N_11936,N_6781,N_8220);
nor U11937 (N_11937,N_5836,N_9599);
or U11938 (N_11938,N_9368,N_8516);
nand U11939 (N_11939,N_5182,N_7833);
xor U11940 (N_11940,N_8023,N_9030);
and U11941 (N_11941,N_5366,N_6122);
and U11942 (N_11942,N_9779,N_9770);
nor U11943 (N_11943,N_9590,N_7346);
xor U11944 (N_11944,N_9383,N_9840);
nor U11945 (N_11945,N_8832,N_9773);
xnor U11946 (N_11946,N_7674,N_5168);
and U11947 (N_11947,N_8305,N_6846);
xor U11948 (N_11948,N_9764,N_9760);
and U11949 (N_11949,N_9877,N_7261);
or U11950 (N_11950,N_6236,N_7619);
nand U11951 (N_11951,N_7897,N_5284);
xnor U11952 (N_11952,N_9993,N_9742);
or U11953 (N_11953,N_9728,N_6684);
nor U11954 (N_11954,N_7413,N_5187);
and U11955 (N_11955,N_8279,N_5643);
xnor U11956 (N_11956,N_6496,N_5228);
nand U11957 (N_11957,N_9480,N_6562);
or U11958 (N_11958,N_9351,N_9488);
nand U11959 (N_11959,N_7677,N_8787);
xor U11960 (N_11960,N_8772,N_9252);
and U11961 (N_11961,N_6206,N_8563);
nand U11962 (N_11962,N_6052,N_9883);
nor U11963 (N_11963,N_9428,N_8706);
xnor U11964 (N_11964,N_9337,N_8811);
or U11965 (N_11965,N_9820,N_7182);
xor U11966 (N_11966,N_5927,N_8401);
and U11967 (N_11967,N_6154,N_5092);
nand U11968 (N_11968,N_9002,N_5684);
and U11969 (N_11969,N_5697,N_9423);
xor U11970 (N_11970,N_7087,N_8167);
xnor U11971 (N_11971,N_5928,N_7692);
nor U11972 (N_11972,N_6250,N_9863);
xor U11973 (N_11973,N_6950,N_9017);
nand U11974 (N_11974,N_9162,N_9379);
xor U11975 (N_11975,N_5857,N_5043);
and U11976 (N_11976,N_5988,N_7333);
or U11977 (N_11977,N_7127,N_5242);
xnor U11978 (N_11978,N_5018,N_5689);
or U11979 (N_11979,N_6421,N_8932);
nor U11980 (N_11980,N_8261,N_7944);
or U11981 (N_11981,N_8396,N_6758);
or U11982 (N_11982,N_9165,N_6624);
xnor U11983 (N_11983,N_7410,N_8101);
nand U11984 (N_11984,N_6641,N_8868);
or U11985 (N_11985,N_5106,N_7541);
or U11986 (N_11986,N_7337,N_5969);
nor U11987 (N_11987,N_8016,N_8946);
or U11988 (N_11988,N_8340,N_6106);
nand U11989 (N_11989,N_7757,N_9942);
or U11990 (N_11990,N_7091,N_7974);
xor U11991 (N_11991,N_6509,N_8919);
xnor U11992 (N_11992,N_6742,N_5053);
nor U11993 (N_11993,N_9403,N_5379);
xnor U11994 (N_11994,N_7118,N_9003);
nor U11995 (N_11995,N_7853,N_8358);
or U11996 (N_11996,N_9635,N_8905);
nand U11997 (N_11997,N_8464,N_7367);
or U11998 (N_11998,N_8025,N_9458);
nor U11999 (N_11999,N_6649,N_6683);
and U12000 (N_12000,N_8375,N_8528);
or U12001 (N_12001,N_7580,N_9258);
or U12002 (N_12002,N_8578,N_5502);
xnor U12003 (N_12003,N_7924,N_6656);
and U12004 (N_12004,N_5134,N_9013);
or U12005 (N_12005,N_9509,N_8824);
or U12006 (N_12006,N_7651,N_9354);
xnor U12007 (N_12007,N_5260,N_8450);
and U12008 (N_12008,N_8500,N_6277);
xnor U12009 (N_12009,N_7071,N_7283);
or U12010 (N_12010,N_6070,N_9467);
or U12011 (N_12011,N_9595,N_8033);
or U12012 (N_12012,N_9799,N_5422);
xnor U12013 (N_12013,N_7008,N_9777);
nor U12014 (N_12014,N_5822,N_8671);
xnor U12015 (N_12015,N_8331,N_7085);
nand U12016 (N_12016,N_9286,N_9169);
nor U12017 (N_12017,N_9317,N_7995);
nor U12018 (N_12018,N_6545,N_9903);
xor U12019 (N_12019,N_6608,N_7212);
nor U12020 (N_12020,N_5606,N_6709);
nand U12021 (N_12021,N_8975,N_6031);
xor U12022 (N_12022,N_8636,N_5766);
and U12023 (N_12023,N_7831,N_9046);
xnor U12024 (N_12024,N_8743,N_8057);
xor U12025 (N_12025,N_6653,N_9717);
xor U12026 (N_12026,N_7758,N_6902);
and U12027 (N_12027,N_6919,N_8568);
nor U12028 (N_12028,N_7341,N_8332);
xor U12029 (N_12029,N_8223,N_5986);
and U12030 (N_12030,N_8925,N_8872);
nand U12031 (N_12031,N_6497,N_9198);
or U12032 (N_12032,N_9019,N_6521);
and U12033 (N_12033,N_9327,N_8571);
nor U12034 (N_12034,N_7797,N_8805);
nand U12035 (N_12035,N_6266,N_5008);
or U12036 (N_12036,N_6775,N_9270);
nor U12037 (N_12037,N_9744,N_6877);
nand U12038 (N_12038,N_6726,N_9845);
xnor U12039 (N_12039,N_7601,N_6189);
and U12040 (N_12040,N_5476,N_9955);
or U12041 (N_12041,N_5860,N_7907);
or U12042 (N_12042,N_7941,N_9095);
xor U12043 (N_12043,N_8163,N_5622);
and U12044 (N_12044,N_9127,N_9025);
or U12045 (N_12045,N_8088,N_9122);
nand U12046 (N_12046,N_6342,N_8542);
nand U12047 (N_12047,N_8115,N_5810);
nand U12048 (N_12048,N_9005,N_8858);
nor U12049 (N_12049,N_6581,N_8931);
nor U12050 (N_12050,N_8976,N_9061);
nand U12051 (N_12051,N_8909,N_6664);
and U12052 (N_12052,N_9836,N_7416);
or U12053 (N_12053,N_5440,N_5381);
nor U12054 (N_12054,N_8507,N_5943);
or U12055 (N_12055,N_8489,N_8773);
and U12056 (N_12056,N_8641,N_8843);
xnor U12057 (N_12057,N_7986,N_7221);
nor U12058 (N_12058,N_6374,N_9101);
or U12059 (N_12059,N_8606,N_9850);
or U12060 (N_12060,N_7038,N_9376);
xnor U12061 (N_12061,N_7761,N_6891);
and U12062 (N_12062,N_5581,N_5561);
nand U12063 (N_12063,N_8592,N_8675);
nand U12064 (N_12064,N_7073,N_7547);
nand U12065 (N_12065,N_9677,N_7251);
xor U12066 (N_12066,N_5071,N_9407);
and U12067 (N_12067,N_7542,N_9539);
or U12068 (N_12068,N_7953,N_5370);
xnor U12069 (N_12069,N_7967,N_9168);
nand U12070 (N_12070,N_7448,N_8726);
nand U12071 (N_12071,N_7459,N_9804);
or U12072 (N_12072,N_5728,N_9191);
nor U12073 (N_12073,N_6692,N_7370);
nor U12074 (N_12074,N_6583,N_8570);
nand U12075 (N_12075,N_9471,N_7285);
nor U12076 (N_12076,N_9466,N_8418);
and U12077 (N_12077,N_5285,N_5131);
xor U12078 (N_12078,N_5704,N_8948);
and U12079 (N_12079,N_9835,N_6043);
xnor U12080 (N_12080,N_9164,N_6565);
nor U12081 (N_12081,N_6903,N_5560);
nor U12082 (N_12082,N_6502,N_6805);
xor U12083 (N_12083,N_7011,N_7964);
nor U12084 (N_12084,N_5396,N_7950);
nand U12085 (N_12085,N_9465,N_5853);
or U12086 (N_12086,N_7442,N_8680);
xnor U12087 (N_12087,N_5628,N_9525);
xnor U12088 (N_12088,N_5782,N_7173);
xor U12089 (N_12089,N_5700,N_8496);
nand U12090 (N_12090,N_5801,N_7863);
xnor U12091 (N_12091,N_8335,N_6297);
and U12092 (N_12092,N_8642,N_6449);
nor U12093 (N_12093,N_5573,N_8894);
nand U12094 (N_12094,N_5039,N_7603);
nor U12095 (N_12095,N_8390,N_7536);
nor U12096 (N_12096,N_7587,N_8620);
and U12097 (N_12097,N_7703,N_9501);
xor U12098 (N_12098,N_7850,N_7272);
xor U12099 (N_12099,N_7787,N_7597);
and U12100 (N_12100,N_8404,N_8524);
nand U12101 (N_12101,N_8756,N_9527);
nor U12102 (N_12102,N_6448,N_7952);
and U12103 (N_12103,N_6976,N_5240);
or U12104 (N_12104,N_5031,N_8828);
nand U12105 (N_12105,N_6361,N_8875);
nand U12106 (N_12106,N_9888,N_5804);
nand U12107 (N_12107,N_7726,N_6933);
nand U12108 (N_12108,N_8322,N_9485);
nor U12109 (N_12109,N_8119,N_8654);
xnor U12110 (N_12110,N_8051,N_8584);
nand U12111 (N_12111,N_6535,N_5065);
nor U12112 (N_12112,N_9946,N_5318);
xor U12113 (N_12113,N_7996,N_6299);
nand U12114 (N_12114,N_9720,N_5513);
or U12115 (N_12115,N_6411,N_9202);
or U12116 (N_12116,N_9547,N_8522);
nor U12117 (N_12117,N_6262,N_8712);
or U12118 (N_12118,N_5598,N_6415);
nor U12119 (N_12119,N_9118,N_8239);
nand U12120 (N_12120,N_8074,N_8243);
and U12121 (N_12121,N_8129,N_8014);
nand U12122 (N_12122,N_7172,N_7582);
or U12123 (N_12123,N_8795,N_6873);
nor U12124 (N_12124,N_6506,N_7479);
or U12125 (N_12125,N_9617,N_5655);
nand U12126 (N_12126,N_7352,N_8164);
or U12127 (N_12127,N_5865,N_7500);
nor U12128 (N_12128,N_8956,N_9020);
or U12129 (N_12129,N_8130,N_8616);
and U12130 (N_12130,N_6955,N_7746);
nor U12131 (N_12131,N_8471,N_7192);
nor U12132 (N_12132,N_7741,N_9775);
nand U12133 (N_12133,N_5874,N_5368);
xor U12134 (N_12134,N_7878,N_6580);
xnor U12135 (N_12135,N_7415,N_9016);
nor U12136 (N_12136,N_9671,N_6979);
and U12137 (N_12137,N_7082,N_5015);
nor U12138 (N_12138,N_9130,N_7676);
xnor U12139 (N_12139,N_5699,N_5816);
or U12140 (N_12140,N_6395,N_9175);
xor U12141 (N_12141,N_6036,N_8556);
and U12142 (N_12142,N_8771,N_9884);
and U12143 (N_12143,N_6305,N_6240);
xor U12144 (N_12144,N_6317,N_5976);
and U12145 (N_12145,N_9958,N_6256);
nand U12146 (N_12146,N_5266,N_7606);
nor U12147 (N_12147,N_5490,N_8964);
nor U12148 (N_12148,N_5009,N_5211);
nor U12149 (N_12149,N_7763,N_9086);
xnor U12150 (N_12150,N_7219,N_8442);
or U12151 (N_12151,N_9522,N_6107);
and U12152 (N_12152,N_8175,N_6687);
xor U12153 (N_12153,N_8395,N_8048);
xor U12154 (N_12154,N_7238,N_6760);
and U12155 (N_12155,N_5310,N_7075);
nor U12156 (N_12156,N_8244,N_7074);
and U12157 (N_12157,N_8954,N_5659);
xnor U12158 (N_12158,N_5338,N_7468);
nand U12159 (N_12159,N_7269,N_8899);
or U12160 (N_12160,N_7263,N_5088);
xnor U12161 (N_12161,N_8385,N_5292);
xnor U12162 (N_12162,N_6444,N_9865);
and U12163 (N_12163,N_6523,N_9616);
nor U12164 (N_12164,N_6661,N_8733);
nand U12165 (N_12165,N_5016,N_6294);
and U12166 (N_12166,N_6281,N_8281);
and U12167 (N_12167,N_6939,N_5044);
nor U12168 (N_12168,N_9211,N_6227);
xnor U12169 (N_12169,N_5279,N_6440);
nor U12170 (N_12170,N_5436,N_9703);
nand U12171 (N_12171,N_5252,N_7901);
and U12172 (N_12172,N_7802,N_9268);
nand U12173 (N_12173,N_7839,N_6001);
nor U12174 (N_12174,N_8855,N_8724);
nand U12175 (N_12175,N_5034,N_8209);
or U12176 (N_12176,N_8381,N_5198);
nand U12177 (N_12177,N_7309,N_7066);
and U12178 (N_12178,N_6543,N_9867);
nand U12179 (N_12179,N_8838,N_9204);
and U12180 (N_12180,N_7968,N_6493);
nor U12181 (N_12181,N_7700,N_8892);
and U12182 (N_12182,N_7657,N_5277);
or U12183 (N_12183,N_6946,N_8822);
or U12184 (N_12184,N_8484,N_9923);
or U12185 (N_12185,N_6597,N_9684);
nor U12186 (N_12186,N_8472,N_5177);
and U12187 (N_12187,N_7051,N_5676);
nor U12188 (N_12188,N_8646,N_5165);
xor U12189 (N_12189,N_6993,N_8068);
and U12190 (N_12190,N_9373,N_8452);
xor U12191 (N_12191,N_7052,N_9054);
or U12192 (N_12192,N_6825,N_5418);
nand U12193 (N_12193,N_5916,N_6037);
nor U12194 (N_12194,N_9868,N_5727);
and U12195 (N_12195,N_6985,N_8266);
and U12196 (N_12196,N_8668,N_5172);
xnor U12197 (N_12197,N_9771,N_9318);
and U12198 (N_12198,N_6880,N_7409);
and U12199 (N_12199,N_9765,N_6074);
nand U12200 (N_12200,N_5963,N_9665);
nor U12201 (N_12201,N_9104,N_9398);
nand U12202 (N_12202,N_5389,N_5947);
or U12203 (N_12203,N_5539,N_9894);
or U12204 (N_12204,N_6047,N_7147);
nor U12205 (N_12205,N_7421,N_7589);
nand U12206 (N_12206,N_8073,N_7503);
or U12207 (N_12207,N_8614,N_9462);
or U12208 (N_12208,N_7378,N_5119);
nand U12209 (N_12209,N_9793,N_5317);
xnor U12210 (N_12210,N_6949,N_9736);
or U12211 (N_12211,N_8090,N_8010);
nor U12212 (N_12212,N_8533,N_6912);
nand U12213 (N_12213,N_7918,N_5243);
xnor U12214 (N_12214,N_8440,N_8473);
xor U12215 (N_12215,N_9710,N_8588);
nor U12216 (N_12216,N_5696,N_9618);
nand U12217 (N_12217,N_9259,N_7158);
nor U12218 (N_12218,N_7430,N_6582);
and U12219 (N_12219,N_7281,N_8965);
xnor U12220 (N_12220,N_6265,N_6092);
xor U12221 (N_12221,N_5483,N_9332);
and U12222 (N_12222,N_9313,N_7246);
nand U12223 (N_12223,N_6546,N_9537);
xnor U12224 (N_12224,N_6327,N_8036);
and U12225 (N_12225,N_5668,N_5555);
nand U12226 (N_12226,N_9374,N_6759);
nor U12227 (N_12227,N_5951,N_5636);
nand U12228 (N_12228,N_6059,N_8276);
or U12229 (N_12229,N_6359,N_8072);
xnor U12230 (N_12230,N_7244,N_9893);
xor U12231 (N_12231,N_9934,N_5234);
and U12232 (N_12232,N_8518,N_7009);
and U12233 (N_12233,N_8841,N_6893);
nand U12234 (N_12234,N_7161,N_7454);
nor U12235 (N_12235,N_7613,N_8327);
or U12236 (N_12236,N_7424,N_7342);
nand U12237 (N_12237,N_9809,N_5577);
nand U12238 (N_12238,N_7643,N_8313);
xnor U12239 (N_12239,N_6747,N_8151);
and U12240 (N_12240,N_9093,N_7583);
nand U12241 (N_12241,N_7752,N_7894);
nand U12242 (N_12242,N_7360,N_7295);
nand U12243 (N_12243,N_8219,N_9084);
nand U12244 (N_12244,N_8204,N_8232);
or U12245 (N_12245,N_5500,N_9598);
or U12246 (N_12246,N_6646,N_6851);
nor U12247 (N_12247,N_8818,N_7930);
and U12248 (N_12248,N_7822,N_8958);
nor U12249 (N_12249,N_9140,N_7132);
and U12250 (N_12250,N_6130,N_8122);
or U12251 (N_12251,N_6639,N_9476);
and U12252 (N_12252,N_9609,N_7615);
nand U12253 (N_12253,N_6406,N_7394);
xnor U12254 (N_12254,N_5892,N_8691);
nand U12255 (N_12255,N_7287,N_6100);
nor U12256 (N_12256,N_8986,N_7376);
xnor U12257 (N_12257,N_9965,N_7340);
nand U12258 (N_12258,N_5104,N_6942);
nor U12259 (N_12259,N_8435,N_7998);
xor U12260 (N_12260,N_6510,N_6464);
or U12261 (N_12261,N_5320,N_6604);
xnor U12262 (N_12262,N_8229,N_6212);
nand U12263 (N_12263,N_7312,N_9505);
nor U12264 (N_12264,N_6970,N_7055);
and U12265 (N_12265,N_5633,N_7889);
or U12266 (N_12266,N_9608,N_8159);
nor U12267 (N_12267,N_7975,N_7314);
nand U12268 (N_12268,N_8765,N_7171);
xnor U12269 (N_12269,N_9143,N_9150);
and U12270 (N_12270,N_6953,N_7660);
and U12271 (N_12271,N_8994,N_5144);
and U12272 (N_12272,N_8387,N_9216);
or U12273 (N_12273,N_5839,N_6416);
and U12274 (N_12274,N_7514,N_8035);
xor U12275 (N_12275,N_9630,N_9749);
and U12276 (N_12276,N_7231,N_6272);
xor U12277 (N_12277,N_6390,N_8416);
nor U12278 (N_12278,N_9146,N_8827);
nand U12279 (N_12279,N_9638,N_9396);
nor U12280 (N_12280,N_9413,N_8413);
xor U12281 (N_12281,N_9155,N_5394);
and U12282 (N_12282,N_8351,N_7638);
nor U12283 (N_12283,N_5109,N_8490);
xor U12284 (N_12284,N_5095,N_9257);
nor U12285 (N_12285,N_8599,N_5789);
xnor U12286 (N_12286,N_8187,N_9001);
nand U12287 (N_12287,N_7151,N_6364);
and U12288 (N_12288,N_8744,N_9737);
nand U12289 (N_12289,N_5012,N_6251);
xnor U12290 (N_12290,N_9943,N_8677);
or U12291 (N_12291,N_5064,N_8445);
nor U12292 (N_12292,N_5196,N_7404);
nand U12293 (N_12293,N_5374,N_8549);
xor U12294 (N_12294,N_9543,N_7985);
nor U12295 (N_12295,N_6592,N_5321);
nor U12296 (N_12296,N_6602,N_9875);
nand U12297 (N_12297,N_6271,N_8821);
or U12298 (N_12298,N_8647,N_9096);
and U12299 (N_12299,N_7080,N_9389);
nor U12300 (N_12300,N_7115,N_8213);
and U12301 (N_12301,N_9384,N_5908);
nand U12302 (N_12302,N_8046,N_7517);
nor U12303 (N_12303,N_5796,N_6150);
or U12304 (N_12304,N_7316,N_8741);
nor U12305 (N_12305,N_7879,N_6847);
nor U12306 (N_12306,N_7695,N_6048);
and U12307 (N_12307,N_5682,N_6008);
and U12308 (N_12308,N_7293,N_8997);
nor U12309 (N_12309,N_7211,N_9738);
or U12310 (N_12310,N_9824,N_6476);
or U12311 (N_12311,N_8184,N_9727);
or U12312 (N_12312,N_8493,N_5638);
nand U12313 (N_12313,N_6492,N_8211);
nand U12314 (N_12314,N_7955,N_9832);
xnor U12315 (N_12315,N_5953,N_6318);
nand U12316 (N_12316,N_7264,N_5289);
nand U12317 (N_12317,N_8465,N_9619);
nor U12318 (N_12318,N_7274,N_6084);
and U12319 (N_12319,N_8817,N_5118);
nor U12320 (N_12320,N_6663,N_7871);
or U12321 (N_12321,N_6749,N_7525);
nand U12322 (N_12322,N_8940,N_5082);
or U12323 (N_12323,N_7826,N_8626);
and U12324 (N_12324,N_6790,N_5385);
xnor U12325 (N_12325,N_8432,N_5363);
nand U12326 (N_12326,N_5703,N_6193);
nor U12327 (N_12327,N_7486,N_5382);
xnor U12328 (N_12328,N_9748,N_7178);
xor U12329 (N_12329,N_8583,N_6558);
nor U12330 (N_12330,N_8208,N_8856);
and U12331 (N_12331,N_9656,N_9276);
nor U12332 (N_12332,N_8720,N_6957);
xor U12333 (N_12333,N_6368,N_9918);
or U12334 (N_12334,N_7520,N_9739);
or U12335 (N_12335,N_5202,N_7497);
nand U12336 (N_12336,N_6524,N_5797);
or U12337 (N_12337,N_6187,N_9073);
and U12338 (N_12338,N_7713,N_5006);
or U12339 (N_12339,N_5867,N_7379);
or U12340 (N_12340,N_9147,N_6451);
xnor U12341 (N_12341,N_5678,N_7498);
and U12342 (N_12342,N_7859,N_8552);
and U12343 (N_12343,N_6046,N_6471);
nand U12344 (N_12344,N_6218,N_9869);
xnor U12345 (N_12345,N_6462,N_5354);
nand U12346 (N_12346,N_7786,N_7025);
or U12347 (N_12347,N_5115,N_5761);
or U12348 (N_12348,N_5495,N_5649);
and U12349 (N_12349,N_8265,N_7612);
nor U12350 (N_12350,N_9455,N_5694);
and U12351 (N_12351,N_8042,N_7927);
and U12352 (N_12352,N_8711,N_7518);
and U12353 (N_12353,N_6917,N_7411);
nand U12354 (N_12354,N_6778,N_5920);
or U12355 (N_12355,N_5665,N_9812);
or U12356 (N_12356,N_5122,N_9857);
nor U12357 (N_12357,N_9682,N_5921);
or U12358 (N_12358,N_7078,N_5715);
or U12359 (N_12359,N_6058,N_7605);
nand U12360 (N_12360,N_5881,N_8891);
xor U12361 (N_12361,N_5173,N_8840);
or U12362 (N_12362,N_5967,N_8260);
or U12363 (N_12363,N_8468,N_6136);
and U12364 (N_12364,N_8317,N_7512);
xnor U12365 (N_12365,N_6050,N_7956);
nand U12366 (N_12366,N_7992,N_7202);
nor U12367 (N_12367,N_6275,N_5171);
nand U12368 (N_12368,N_7481,N_5756);
nor U12369 (N_12369,N_7432,N_6867);
or U12370 (N_12370,N_8506,N_6553);
nor U12371 (N_12371,N_8694,N_8663);
and U12372 (N_12372,N_6254,N_6159);
and U12373 (N_12373,N_6016,N_8878);
xor U12374 (N_12374,N_9839,N_7088);
nor U12375 (N_12375,N_5856,N_6452);
nor U12376 (N_12376,N_5373,N_5504);
nand U12377 (N_12377,N_7538,N_9214);
xor U12378 (N_12378,N_5934,N_6862);
or U12379 (N_12379,N_7823,N_9057);
nor U12380 (N_12380,N_9729,N_8625);
nor U12381 (N_12381,N_5914,N_7245);
nor U12382 (N_12382,N_9217,N_7684);
xor U12383 (N_12383,N_9921,N_9512);
xor U12384 (N_12384,N_7336,N_9715);
and U12385 (N_12385,N_7844,N_6941);
nor U12386 (N_12386,N_6980,N_5778);
nand U12387 (N_12387,N_7456,N_8132);
or U12388 (N_12388,N_5587,N_7329);
or U12389 (N_12389,N_9640,N_5501);
or U12390 (N_12390,N_9344,N_5397);
xor U12391 (N_12391,N_7793,N_6554);
or U12392 (N_12392,N_6757,N_6617);
or U12393 (N_12393,N_8531,N_5116);
or U12394 (N_12394,N_7798,N_6424);
nor U12395 (N_12395,N_5971,N_7320);
and U12396 (N_12396,N_8403,N_9012);
and U12397 (N_12397,N_9920,N_9841);
xnor U12398 (N_12398,N_7981,N_7856);
and U12399 (N_12399,N_5825,N_8666);
nor U12400 (N_12400,N_9719,N_9365);
or U12401 (N_12401,N_7926,N_7391);
nor U12402 (N_12402,N_6651,N_9806);
and U12403 (N_12403,N_5257,N_6221);
xor U12404 (N_12404,N_5533,N_9917);
nand U12405 (N_12405,N_9112,N_6377);
nand U12406 (N_12406,N_8457,N_8804);
xnor U12407 (N_12407,N_6672,N_6027);
and U12408 (N_12408,N_7970,N_6794);
xnor U12409 (N_12409,N_9928,N_8227);
nor U12410 (N_12410,N_6712,N_9678);
or U12411 (N_12411,N_7386,N_5141);
nand U12412 (N_12412,N_7740,N_6732);
nor U12413 (N_12413,N_9945,N_6795);
nand U12414 (N_12414,N_5227,N_7495);
or U12415 (N_12415,N_7796,N_9998);
nor U12416 (N_12416,N_6252,N_9674);
xor U12417 (N_12417,N_9273,N_5457);
xnor U12418 (N_12418,N_5850,N_5512);
xnor U12419 (N_12419,N_9786,N_9614);
nor U12420 (N_12420,N_7234,N_8254);
nor U12421 (N_12421,N_7568,N_7837);
nand U12422 (N_12422,N_7189,N_9704);
and U12423 (N_12423,N_7037,N_8676);
and U12424 (N_12424,N_5763,N_6974);
and U12425 (N_12425,N_5511,N_5186);
nand U12426 (N_12426,N_9535,N_5974);
or U12427 (N_12427,N_5269,N_7782);
xnor U12428 (N_12428,N_5004,N_7579);
nor U12429 (N_12429,N_7201,N_9784);
nor U12430 (N_12430,N_7113,N_9163);
nand U12431 (N_12431,N_5593,N_7277);
and U12432 (N_12432,N_9844,N_7369);
xor U12433 (N_12433,N_9375,N_5741);
xnor U12434 (N_12434,N_6076,N_8364);
nand U12435 (N_12435,N_8303,N_9795);
nor U12436 (N_12436,N_9895,N_5862);
nand U12437 (N_12437,N_6109,N_9520);
xor U12438 (N_12438,N_6422,N_9994);
xnor U12439 (N_12439,N_9655,N_9406);
or U12440 (N_12440,N_6055,N_8277);
xor U12441 (N_12441,N_6332,N_8974);
or U12442 (N_12442,N_8699,N_6409);
xor U12443 (N_12443,N_5270,N_5302);
and U12444 (N_12444,N_5869,N_8414);
or U12445 (N_12445,N_8551,N_8586);
nor U12446 (N_12446,N_5113,N_6347);
or U12447 (N_12447,N_8502,N_7715);
nand U12448 (N_12448,N_5046,N_9048);
and U12449 (N_12449,N_8427,N_6182);
nand U12450 (N_12450,N_9416,N_7593);
nand U12451 (N_12451,N_7358,N_7252);
nor U12452 (N_12452,N_6932,N_9855);
xor U12453 (N_12453,N_5937,N_9111);
and U12454 (N_12454,N_5101,N_8222);
xor U12455 (N_12455,N_8873,N_7604);
or U12456 (N_12456,N_8850,N_9849);
and U12457 (N_12457,N_9979,N_9129);
xnor U12458 (N_12458,N_7494,N_8750);
nor U12459 (N_12459,N_8214,N_7569);
xor U12460 (N_12460,N_7062,N_5556);
or U12461 (N_12461,N_5130,N_7767);
nor U12462 (N_12462,N_6487,N_5473);
nor U12463 (N_12463,N_5313,N_8017);
and U12464 (N_12464,N_5627,N_7776);
nand U12465 (N_12465,N_6365,N_6054);
nor U12466 (N_12466,N_6023,N_6828);
or U12467 (N_12467,N_9768,N_5531);
xnor U12468 (N_12468,N_5314,N_8884);
nand U12469 (N_12469,N_6515,N_8982);
nand U12470 (N_12470,N_5358,N_7733);
or U12471 (N_12471,N_8082,N_5604);
nand U12472 (N_12472,N_7706,N_9755);
or U12473 (N_12473,N_7056,N_7213);
xnor U12474 (N_12474,N_6568,N_6567);
nand U12475 (N_12475,N_8032,N_8602);
nand U12476 (N_12476,N_7745,N_9069);
and U12477 (N_12477,N_6681,N_8267);
xnor U12478 (N_12478,N_9102,N_5158);
or U12479 (N_12479,N_9588,N_9532);
and U12480 (N_12480,N_9103,N_8497);
xnor U12481 (N_12481,N_6200,N_6149);
nor U12482 (N_12482,N_8515,N_9542);
xor U12483 (N_12483,N_5420,N_8495);
or U12484 (N_12484,N_5024,N_9430);
xor U12485 (N_12485,N_5961,N_9890);
xor U12486 (N_12486,N_8897,N_7194);
xor U12487 (N_12487,N_8217,N_9366);
and U12488 (N_12488,N_8779,N_9573);
nor U12489 (N_12489,N_8237,N_8898);
xnor U12490 (N_12490,N_6723,N_8788);
and U12491 (N_12491,N_7324,N_8731);
nand U12492 (N_12492,N_6984,N_6616);
xnor U12493 (N_12493,N_5773,N_7208);
or U12494 (N_12494,N_7027,N_8967);
or U12495 (N_12495,N_5330,N_6935);
and U12496 (N_12496,N_8622,N_8988);
or U12497 (N_12497,N_8833,N_8105);
nor U12498 (N_12498,N_7491,N_5645);
xor U12499 (N_12499,N_7665,N_5491);
xor U12500 (N_12500,N_6212,N_9181);
nand U12501 (N_12501,N_5557,N_8690);
and U12502 (N_12502,N_8484,N_5426);
nor U12503 (N_12503,N_7233,N_9204);
and U12504 (N_12504,N_9639,N_7162);
and U12505 (N_12505,N_9453,N_7463);
xnor U12506 (N_12506,N_6108,N_5864);
and U12507 (N_12507,N_7553,N_8210);
nor U12508 (N_12508,N_9317,N_7779);
nor U12509 (N_12509,N_6013,N_8443);
nor U12510 (N_12510,N_9778,N_8373);
and U12511 (N_12511,N_8512,N_6026);
and U12512 (N_12512,N_9424,N_7965);
nand U12513 (N_12513,N_7073,N_6650);
xor U12514 (N_12514,N_7076,N_7055);
xor U12515 (N_12515,N_8530,N_9707);
nor U12516 (N_12516,N_9941,N_5638);
nor U12517 (N_12517,N_5015,N_5161);
nand U12518 (N_12518,N_8826,N_8232);
nor U12519 (N_12519,N_8958,N_6578);
or U12520 (N_12520,N_9648,N_6303);
nor U12521 (N_12521,N_9230,N_5983);
xor U12522 (N_12522,N_9952,N_8143);
xnor U12523 (N_12523,N_6900,N_9984);
xnor U12524 (N_12524,N_7907,N_5018);
xor U12525 (N_12525,N_9023,N_8545);
nor U12526 (N_12526,N_7952,N_7289);
xor U12527 (N_12527,N_8473,N_5211);
or U12528 (N_12528,N_8747,N_6795);
or U12529 (N_12529,N_7524,N_6455);
xor U12530 (N_12530,N_5920,N_9591);
nand U12531 (N_12531,N_7752,N_6017);
and U12532 (N_12532,N_5449,N_5639);
xor U12533 (N_12533,N_9723,N_7423);
nand U12534 (N_12534,N_8996,N_5046);
and U12535 (N_12535,N_6326,N_6285);
nor U12536 (N_12536,N_8685,N_9693);
nand U12537 (N_12537,N_8061,N_8303);
and U12538 (N_12538,N_9281,N_6393);
and U12539 (N_12539,N_9710,N_5629);
and U12540 (N_12540,N_5925,N_9281);
nand U12541 (N_12541,N_8502,N_5962);
or U12542 (N_12542,N_7636,N_9339);
xnor U12543 (N_12543,N_5773,N_7541);
xnor U12544 (N_12544,N_9988,N_7166);
xor U12545 (N_12545,N_5008,N_9737);
nand U12546 (N_12546,N_5223,N_6303);
or U12547 (N_12547,N_7584,N_9911);
nand U12548 (N_12548,N_7682,N_8487);
xor U12549 (N_12549,N_5763,N_6423);
nand U12550 (N_12550,N_7355,N_9464);
nand U12551 (N_12551,N_7991,N_7118);
or U12552 (N_12552,N_5685,N_5487);
xnor U12553 (N_12553,N_9037,N_5510);
or U12554 (N_12554,N_9775,N_7750);
xnor U12555 (N_12555,N_8956,N_7228);
and U12556 (N_12556,N_6187,N_7287);
nor U12557 (N_12557,N_7959,N_8240);
xor U12558 (N_12558,N_8672,N_6112);
and U12559 (N_12559,N_6768,N_7673);
and U12560 (N_12560,N_9784,N_6417);
nand U12561 (N_12561,N_8720,N_8385);
or U12562 (N_12562,N_7491,N_7588);
and U12563 (N_12563,N_7948,N_5936);
and U12564 (N_12564,N_7671,N_7143);
and U12565 (N_12565,N_5735,N_6202);
and U12566 (N_12566,N_6566,N_7737);
xnor U12567 (N_12567,N_6784,N_9792);
or U12568 (N_12568,N_7616,N_9348);
xnor U12569 (N_12569,N_8558,N_5174);
or U12570 (N_12570,N_5328,N_7051);
nor U12571 (N_12571,N_6183,N_8271);
or U12572 (N_12572,N_9138,N_9508);
xnor U12573 (N_12573,N_9432,N_6625);
or U12574 (N_12574,N_9450,N_7547);
and U12575 (N_12575,N_5625,N_8960);
and U12576 (N_12576,N_5256,N_5911);
xnor U12577 (N_12577,N_8126,N_7754);
and U12578 (N_12578,N_7041,N_9956);
and U12579 (N_12579,N_8376,N_6287);
nand U12580 (N_12580,N_9912,N_8324);
and U12581 (N_12581,N_5712,N_8313);
and U12582 (N_12582,N_9410,N_5733);
or U12583 (N_12583,N_7812,N_9239);
nor U12584 (N_12584,N_6568,N_7001);
nand U12585 (N_12585,N_9029,N_8690);
or U12586 (N_12586,N_5559,N_8280);
and U12587 (N_12587,N_7959,N_7188);
xor U12588 (N_12588,N_7117,N_5131);
or U12589 (N_12589,N_9316,N_6105);
or U12590 (N_12590,N_9559,N_8276);
or U12591 (N_12591,N_6718,N_6254);
and U12592 (N_12592,N_7205,N_7099);
nor U12593 (N_12593,N_9063,N_5518);
or U12594 (N_12594,N_7791,N_9360);
nor U12595 (N_12595,N_6198,N_5887);
nand U12596 (N_12596,N_5398,N_8122);
nand U12597 (N_12597,N_6144,N_8243);
xor U12598 (N_12598,N_9279,N_6129);
nor U12599 (N_12599,N_7318,N_5190);
nand U12600 (N_12600,N_9367,N_9450);
or U12601 (N_12601,N_5466,N_9231);
and U12602 (N_12602,N_7341,N_9939);
xor U12603 (N_12603,N_9981,N_8842);
nor U12604 (N_12604,N_8744,N_7059);
or U12605 (N_12605,N_5859,N_8696);
or U12606 (N_12606,N_6701,N_7901);
and U12607 (N_12607,N_7887,N_9147);
and U12608 (N_12608,N_6572,N_6051);
or U12609 (N_12609,N_9399,N_9510);
or U12610 (N_12610,N_7539,N_8196);
nor U12611 (N_12611,N_9407,N_7709);
xor U12612 (N_12612,N_9803,N_7469);
nor U12613 (N_12613,N_9142,N_7798);
and U12614 (N_12614,N_9092,N_9426);
nor U12615 (N_12615,N_5570,N_7147);
and U12616 (N_12616,N_6469,N_5353);
xor U12617 (N_12617,N_7267,N_7093);
and U12618 (N_12618,N_6683,N_5979);
or U12619 (N_12619,N_8921,N_9442);
nor U12620 (N_12620,N_9027,N_9886);
nand U12621 (N_12621,N_5449,N_7806);
nand U12622 (N_12622,N_6021,N_8558);
xnor U12623 (N_12623,N_5334,N_6585);
xor U12624 (N_12624,N_5532,N_9605);
nand U12625 (N_12625,N_7742,N_7440);
and U12626 (N_12626,N_5667,N_6698);
nor U12627 (N_12627,N_8003,N_9787);
nand U12628 (N_12628,N_5593,N_8051);
xnor U12629 (N_12629,N_6863,N_7467);
nor U12630 (N_12630,N_8828,N_5972);
and U12631 (N_12631,N_5527,N_6011);
or U12632 (N_12632,N_7712,N_5105);
or U12633 (N_12633,N_6139,N_7633);
nand U12634 (N_12634,N_9506,N_8845);
xor U12635 (N_12635,N_9998,N_6100);
and U12636 (N_12636,N_9904,N_9852);
and U12637 (N_12637,N_5827,N_7778);
nor U12638 (N_12638,N_7364,N_8783);
nor U12639 (N_12639,N_6455,N_5150);
nand U12640 (N_12640,N_6309,N_5523);
and U12641 (N_12641,N_7345,N_5010);
xnor U12642 (N_12642,N_9644,N_9972);
or U12643 (N_12643,N_5371,N_6551);
or U12644 (N_12644,N_8506,N_9228);
nand U12645 (N_12645,N_9341,N_5411);
nor U12646 (N_12646,N_8389,N_6801);
nand U12647 (N_12647,N_6912,N_9296);
or U12648 (N_12648,N_8939,N_7097);
nand U12649 (N_12649,N_8885,N_8056);
and U12650 (N_12650,N_5783,N_9495);
nor U12651 (N_12651,N_8049,N_8294);
or U12652 (N_12652,N_8564,N_5013);
and U12653 (N_12653,N_6870,N_8571);
nand U12654 (N_12654,N_7328,N_9933);
xnor U12655 (N_12655,N_6303,N_9031);
xor U12656 (N_12656,N_9223,N_5808);
and U12657 (N_12657,N_9423,N_5231);
nand U12658 (N_12658,N_7606,N_6402);
xnor U12659 (N_12659,N_8871,N_5818);
xnor U12660 (N_12660,N_6470,N_7529);
nand U12661 (N_12661,N_5669,N_6634);
or U12662 (N_12662,N_8677,N_9200);
and U12663 (N_12663,N_8160,N_8180);
or U12664 (N_12664,N_5364,N_7012);
or U12665 (N_12665,N_9776,N_5597);
xnor U12666 (N_12666,N_7054,N_6797);
or U12667 (N_12667,N_9998,N_9930);
xnor U12668 (N_12668,N_5994,N_5475);
xor U12669 (N_12669,N_6471,N_8076);
xnor U12670 (N_12670,N_8018,N_8618);
xor U12671 (N_12671,N_5162,N_9855);
nor U12672 (N_12672,N_5519,N_7491);
nand U12673 (N_12673,N_7392,N_5939);
nor U12674 (N_12674,N_6952,N_7769);
nor U12675 (N_12675,N_5600,N_5800);
nand U12676 (N_12676,N_9620,N_6951);
nor U12677 (N_12677,N_5067,N_9804);
or U12678 (N_12678,N_6604,N_6512);
and U12679 (N_12679,N_9765,N_5088);
nor U12680 (N_12680,N_8217,N_6625);
xnor U12681 (N_12681,N_8373,N_5260);
or U12682 (N_12682,N_5207,N_7323);
nand U12683 (N_12683,N_6084,N_7607);
xor U12684 (N_12684,N_9956,N_6550);
xor U12685 (N_12685,N_6329,N_9777);
or U12686 (N_12686,N_8890,N_6648);
nor U12687 (N_12687,N_6140,N_8637);
xor U12688 (N_12688,N_6158,N_7252);
and U12689 (N_12689,N_8174,N_9169);
xor U12690 (N_12690,N_8653,N_9000);
nand U12691 (N_12691,N_9802,N_9585);
and U12692 (N_12692,N_7678,N_9773);
xnor U12693 (N_12693,N_7439,N_6578);
nor U12694 (N_12694,N_6709,N_7160);
nor U12695 (N_12695,N_8956,N_8454);
and U12696 (N_12696,N_9274,N_8217);
nand U12697 (N_12697,N_6317,N_8266);
nor U12698 (N_12698,N_5098,N_5557);
nor U12699 (N_12699,N_5699,N_9018);
nor U12700 (N_12700,N_5702,N_7541);
or U12701 (N_12701,N_8061,N_7944);
or U12702 (N_12702,N_5640,N_6320);
or U12703 (N_12703,N_5939,N_6980);
nor U12704 (N_12704,N_8689,N_8926);
nand U12705 (N_12705,N_5562,N_7296);
xor U12706 (N_12706,N_6009,N_8421);
nor U12707 (N_12707,N_6462,N_6963);
or U12708 (N_12708,N_8488,N_5100);
xor U12709 (N_12709,N_9991,N_6670);
nor U12710 (N_12710,N_7527,N_5680);
nor U12711 (N_12711,N_6906,N_9129);
nor U12712 (N_12712,N_8687,N_8583);
nor U12713 (N_12713,N_8912,N_9245);
nand U12714 (N_12714,N_7226,N_6394);
nand U12715 (N_12715,N_7405,N_9193);
nor U12716 (N_12716,N_6980,N_5462);
nand U12717 (N_12717,N_9254,N_7121);
xor U12718 (N_12718,N_8592,N_7293);
and U12719 (N_12719,N_5936,N_5970);
xnor U12720 (N_12720,N_6870,N_6285);
nor U12721 (N_12721,N_7616,N_7149);
nand U12722 (N_12722,N_5884,N_5592);
or U12723 (N_12723,N_6493,N_9855);
and U12724 (N_12724,N_8297,N_8066);
and U12725 (N_12725,N_7152,N_8886);
nor U12726 (N_12726,N_7074,N_6588);
or U12727 (N_12727,N_6812,N_5156);
or U12728 (N_12728,N_5876,N_7306);
and U12729 (N_12729,N_8194,N_8392);
nand U12730 (N_12730,N_5320,N_7167);
or U12731 (N_12731,N_7831,N_8977);
nand U12732 (N_12732,N_9015,N_9363);
and U12733 (N_12733,N_7553,N_5233);
nor U12734 (N_12734,N_5163,N_5981);
and U12735 (N_12735,N_7052,N_7867);
nor U12736 (N_12736,N_7101,N_5029);
and U12737 (N_12737,N_9555,N_5640);
or U12738 (N_12738,N_7502,N_8408);
nor U12739 (N_12739,N_8178,N_7906);
or U12740 (N_12740,N_9399,N_6020);
or U12741 (N_12741,N_5800,N_8702);
xor U12742 (N_12742,N_7979,N_7981);
nand U12743 (N_12743,N_8868,N_6784);
nand U12744 (N_12744,N_7829,N_6367);
or U12745 (N_12745,N_9670,N_6974);
nand U12746 (N_12746,N_6595,N_9124);
nand U12747 (N_12747,N_9912,N_7499);
nand U12748 (N_12748,N_9475,N_9253);
nor U12749 (N_12749,N_5461,N_5696);
and U12750 (N_12750,N_7416,N_6517);
or U12751 (N_12751,N_5186,N_7166);
nand U12752 (N_12752,N_7598,N_9376);
nor U12753 (N_12753,N_5761,N_9917);
and U12754 (N_12754,N_6962,N_5210);
and U12755 (N_12755,N_9822,N_5134);
nand U12756 (N_12756,N_7478,N_9190);
nor U12757 (N_12757,N_5881,N_6337);
xor U12758 (N_12758,N_9450,N_8845);
nand U12759 (N_12759,N_7303,N_7037);
or U12760 (N_12760,N_6692,N_6073);
xnor U12761 (N_12761,N_7139,N_6379);
xor U12762 (N_12762,N_8377,N_9112);
nand U12763 (N_12763,N_7360,N_6378);
xnor U12764 (N_12764,N_5222,N_9596);
and U12765 (N_12765,N_7819,N_9303);
and U12766 (N_12766,N_7334,N_8609);
or U12767 (N_12767,N_9081,N_8694);
or U12768 (N_12768,N_6999,N_5298);
xor U12769 (N_12769,N_5281,N_8996);
or U12770 (N_12770,N_5966,N_5548);
and U12771 (N_12771,N_8125,N_6375);
xnor U12772 (N_12772,N_7457,N_6584);
nand U12773 (N_12773,N_8392,N_5682);
nand U12774 (N_12774,N_7485,N_6190);
and U12775 (N_12775,N_6191,N_9091);
xnor U12776 (N_12776,N_8574,N_5673);
and U12777 (N_12777,N_8667,N_7389);
xnor U12778 (N_12778,N_6514,N_8872);
or U12779 (N_12779,N_9001,N_9465);
xor U12780 (N_12780,N_8307,N_9472);
nor U12781 (N_12781,N_7089,N_5497);
nand U12782 (N_12782,N_6299,N_6227);
xnor U12783 (N_12783,N_5606,N_6386);
or U12784 (N_12784,N_5663,N_6495);
or U12785 (N_12785,N_8531,N_6084);
or U12786 (N_12786,N_5299,N_9605);
nor U12787 (N_12787,N_5015,N_6535);
or U12788 (N_12788,N_6795,N_7574);
or U12789 (N_12789,N_8777,N_7581);
nand U12790 (N_12790,N_9778,N_6599);
xor U12791 (N_12791,N_9924,N_7804);
and U12792 (N_12792,N_9871,N_5926);
and U12793 (N_12793,N_7864,N_8866);
nand U12794 (N_12794,N_5137,N_8017);
xnor U12795 (N_12795,N_7518,N_5421);
nor U12796 (N_12796,N_9724,N_7927);
nand U12797 (N_12797,N_9876,N_7305);
or U12798 (N_12798,N_9360,N_9726);
nand U12799 (N_12799,N_5583,N_9631);
nand U12800 (N_12800,N_5069,N_5601);
xnor U12801 (N_12801,N_6860,N_5345);
nor U12802 (N_12802,N_8122,N_7479);
nor U12803 (N_12803,N_9332,N_6214);
or U12804 (N_12804,N_6464,N_6617);
nand U12805 (N_12805,N_9855,N_8445);
nand U12806 (N_12806,N_7905,N_5467);
and U12807 (N_12807,N_8241,N_8704);
xor U12808 (N_12808,N_6819,N_7472);
or U12809 (N_12809,N_7825,N_6406);
and U12810 (N_12810,N_8938,N_6398);
xnor U12811 (N_12811,N_9259,N_5198);
nor U12812 (N_12812,N_8413,N_6796);
xnor U12813 (N_12813,N_6565,N_8167);
nand U12814 (N_12814,N_6810,N_8766);
nand U12815 (N_12815,N_7933,N_8711);
or U12816 (N_12816,N_6878,N_9688);
or U12817 (N_12817,N_5562,N_6476);
and U12818 (N_12818,N_5939,N_7727);
and U12819 (N_12819,N_7874,N_9661);
or U12820 (N_12820,N_5646,N_8000);
nand U12821 (N_12821,N_7347,N_8809);
nand U12822 (N_12822,N_7958,N_5773);
nand U12823 (N_12823,N_7041,N_6514);
nor U12824 (N_12824,N_9534,N_5637);
or U12825 (N_12825,N_8458,N_7607);
nor U12826 (N_12826,N_9257,N_8883);
nor U12827 (N_12827,N_5186,N_6545);
xor U12828 (N_12828,N_5212,N_9491);
nor U12829 (N_12829,N_9164,N_7956);
xnor U12830 (N_12830,N_5854,N_7933);
or U12831 (N_12831,N_8843,N_9479);
and U12832 (N_12832,N_8663,N_5039);
nand U12833 (N_12833,N_8049,N_6420);
xnor U12834 (N_12834,N_6381,N_8489);
nand U12835 (N_12835,N_9404,N_6755);
and U12836 (N_12836,N_7198,N_7152);
xor U12837 (N_12837,N_8320,N_7544);
xnor U12838 (N_12838,N_8204,N_8268);
or U12839 (N_12839,N_5789,N_9561);
and U12840 (N_12840,N_5813,N_8308);
or U12841 (N_12841,N_5058,N_5543);
or U12842 (N_12842,N_5860,N_6856);
nor U12843 (N_12843,N_5046,N_9216);
nand U12844 (N_12844,N_9585,N_5826);
xnor U12845 (N_12845,N_6762,N_9345);
or U12846 (N_12846,N_5589,N_5610);
and U12847 (N_12847,N_8415,N_9829);
or U12848 (N_12848,N_5343,N_8090);
nor U12849 (N_12849,N_7324,N_7448);
and U12850 (N_12850,N_7697,N_7135);
xor U12851 (N_12851,N_9025,N_7906);
nand U12852 (N_12852,N_8928,N_6272);
and U12853 (N_12853,N_8685,N_6465);
nor U12854 (N_12854,N_5016,N_6184);
and U12855 (N_12855,N_6306,N_9508);
nor U12856 (N_12856,N_6345,N_5338);
xnor U12857 (N_12857,N_5130,N_6588);
xor U12858 (N_12858,N_7020,N_7224);
and U12859 (N_12859,N_5594,N_6999);
nor U12860 (N_12860,N_9896,N_9633);
or U12861 (N_12861,N_5364,N_9045);
nand U12862 (N_12862,N_8381,N_6135);
nor U12863 (N_12863,N_9629,N_5927);
and U12864 (N_12864,N_6722,N_9255);
nand U12865 (N_12865,N_8441,N_8335);
or U12866 (N_12866,N_6976,N_5611);
and U12867 (N_12867,N_5790,N_5177);
xnor U12868 (N_12868,N_6045,N_7807);
xnor U12869 (N_12869,N_6867,N_6260);
or U12870 (N_12870,N_8592,N_6864);
xnor U12871 (N_12871,N_8928,N_7590);
nor U12872 (N_12872,N_6643,N_7636);
nor U12873 (N_12873,N_8426,N_7213);
and U12874 (N_12874,N_6092,N_6644);
and U12875 (N_12875,N_8804,N_6024);
xor U12876 (N_12876,N_6947,N_6954);
nor U12877 (N_12877,N_8925,N_6553);
nand U12878 (N_12878,N_6095,N_7278);
or U12879 (N_12879,N_7700,N_6842);
nor U12880 (N_12880,N_7942,N_8211);
or U12881 (N_12881,N_9108,N_9318);
nor U12882 (N_12882,N_9679,N_9170);
nor U12883 (N_12883,N_5656,N_9513);
xor U12884 (N_12884,N_9655,N_5823);
xnor U12885 (N_12885,N_8642,N_6347);
nand U12886 (N_12886,N_5385,N_5599);
and U12887 (N_12887,N_7375,N_6456);
and U12888 (N_12888,N_9856,N_8701);
nand U12889 (N_12889,N_9789,N_5881);
or U12890 (N_12890,N_6459,N_5000);
nand U12891 (N_12891,N_7513,N_8584);
or U12892 (N_12892,N_6858,N_8986);
nor U12893 (N_12893,N_8260,N_7458);
and U12894 (N_12894,N_9430,N_8388);
nor U12895 (N_12895,N_7227,N_6697);
nand U12896 (N_12896,N_5746,N_6403);
and U12897 (N_12897,N_8847,N_9551);
nor U12898 (N_12898,N_5897,N_8634);
xor U12899 (N_12899,N_5697,N_9166);
nand U12900 (N_12900,N_6899,N_6852);
nor U12901 (N_12901,N_9043,N_6711);
or U12902 (N_12902,N_7205,N_7290);
nor U12903 (N_12903,N_9394,N_8291);
and U12904 (N_12904,N_9263,N_7569);
nand U12905 (N_12905,N_9239,N_6176);
or U12906 (N_12906,N_5977,N_9501);
nand U12907 (N_12907,N_7527,N_7273);
or U12908 (N_12908,N_8041,N_5646);
and U12909 (N_12909,N_8374,N_7984);
xor U12910 (N_12910,N_5864,N_8958);
and U12911 (N_12911,N_6999,N_5822);
or U12912 (N_12912,N_5149,N_7489);
nand U12913 (N_12913,N_7974,N_6618);
nor U12914 (N_12914,N_6739,N_6598);
nor U12915 (N_12915,N_7283,N_7278);
or U12916 (N_12916,N_9669,N_8340);
or U12917 (N_12917,N_8930,N_5480);
and U12918 (N_12918,N_8713,N_6188);
nand U12919 (N_12919,N_6279,N_6801);
nand U12920 (N_12920,N_9303,N_7394);
and U12921 (N_12921,N_9441,N_9223);
and U12922 (N_12922,N_5167,N_5986);
or U12923 (N_12923,N_6927,N_5933);
nor U12924 (N_12924,N_5892,N_7699);
nor U12925 (N_12925,N_8323,N_5860);
or U12926 (N_12926,N_7540,N_5642);
and U12927 (N_12927,N_6690,N_6539);
nand U12928 (N_12928,N_5724,N_9230);
xnor U12929 (N_12929,N_6464,N_5629);
nand U12930 (N_12930,N_7545,N_5879);
nand U12931 (N_12931,N_8626,N_9310);
nor U12932 (N_12932,N_7127,N_8917);
nor U12933 (N_12933,N_7114,N_9754);
and U12934 (N_12934,N_9971,N_8721);
xnor U12935 (N_12935,N_7564,N_7831);
nand U12936 (N_12936,N_7739,N_8354);
nor U12937 (N_12937,N_6961,N_6483);
and U12938 (N_12938,N_7799,N_9422);
xnor U12939 (N_12939,N_8603,N_9249);
nor U12940 (N_12940,N_7516,N_9388);
or U12941 (N_12941,N_8881,N_8486);
xnor U12942 (N_12942,N_8901,N_8360);
and U12943 (N_12943,N_5501,N_7159);
nand U12944 (N_12944,N_5687,N_5842);
or U12945 (N_12945,N_9444,N_7498);
nor U12946 (N_12946,N_9458,N_6193);
xnor U12947 (N_12947,N_7141,N_8069);
or U12948 (N_12948,N_9706,N_8328);
nor U12949 (N_12949,N_6332,N_5057);
nor U12950 (N_12950,N_6144,N_9365);
or U12951 (N_12951,N_5315,N_5322);
and U12952 (N_12952,N_7711,N_7713);
or U12953 (N_12953,N_8677,N_9032);
nand U12954 (N_12954,N_7359,N_6652);
or U12955 (N_12955,N_6735,N_8916);
nor U12956 (N_12956,N_9302,N_8937);
xnor U12957 (N_12957,N_6750,N_9245);
nor U12958 (N_12958,N_9732,N_7550);
xor U12959 (N_12959,N_8569,N_5720);
nand U12960 (N_12960,N_8465,N_6631);
nor U12961 (N_12961,N_8484,N_6771);
xor U12962 (N_12962,N_7451,N_7793);
or U12963 (N_12963,N_6965,N_7196);
nand U12964 (N_12964,N_7222,N_8989);
xor U12965 (N_12965,N_7242,N_9201);
xnor U12966 (N_12966,N_6368,N_7455);
or U12967 (N_12967,N_5520,N_5007);
or U12968 (N_12968,N_6067,N_8105);
xnor U12969 (N_12969,N_7534,N_6279);
and U12970 (N_12970,N_7831,N_8361);
and U12971 (N_12971,N_9194,N_7899);
xor U12972 (N_12972,N_7557,N_6930);
nand U12973 (N_12973,N_7562,N_9685);
or U12974 (N_12974,N_8279,N_9932);
nor U12975 (N_12975,N_6218,N_8154);
nand U12976 (N_12976,N_8272,N_7923);
xor U12977 (N_12977,N_9852,N_8829);
nand U12978 (N_12978,N_9109,N_5058);
nor U12979 (N_12979,N_5595,N_5066);
xor U12980 (N_12980,N_8131,N_9407);
nand U12981 (N_12981,N_6458,N_8796);
xor U12982 (N_12982,N_9210,N_6743);
nand U12983 (N_12983,N_5443,N_5481);
nand U12984 (N_12984,N_5348,N_7320);
nand U12985 (N_12985,N_7300,N_5801);
or U12986 (N_12986,N_5381,N_7746);
nor U12987 (N_12987,N_7820,N_6468);
nor U12988 (N_12988,N_9012,N_5769);
or U12989 (N_12989,N_5520,N_9088);
and U12990 (N_12990,N_6351,N_8476);
and U12991 (N_12991,N_7316,N_6972);
or U12992 (N_12992,N_8422,N_5005);
nand U12993 (N_12993,N_6584,N_8474);
nand U12994 (N_12994,N_6736,N_5480);
nor U12995 (N_12995,N_8976,N_5827);
xnor U12996 (N_12996,N_8041,N_9351);
nand U12997 (N_12997,N_6812,N_5027);
and U12998 (N_12998,N_7606,N_6005);
and U12999 (N_12999,N_8077,N_8384);
xor U13000 (N_13000,N_9774,N_9808);
xnor U13001 (N_13001,N_9105,N_8791);
and U13002 (N_13002,N_9286,N_5063);
or U13003 (N_13003,N_6312,N_8712);
nand U13004 (N_13004,N_6083,N_8858);
nand U13005 (N_13005,N_8341,N_6150);
xnor U13006 (N_13006,N_7418,N_7216);
nand U13007 (N_13007,N_5624,N_9873);
nand U13008 (N_13008,N_7281,N_5192);
or U13009 (N_13009,N_9216,N_8401);
or U13010 (N_13010,N_9179,N_6095);
or U13011 (N_13011,N_5978,N_9996);
and U13012 (N_13012,N_6774,N_8724);
or U13013 (N_13013,N_7335,N_8073);
xor U13014 (N_13014,N_7182,N_5463);
or U13015 (N_13015,N_6224,N_5641);
or U13016 (N_13016,N_9671,N_8523);
and U13017 (N_13017,N_8511,N_7975);
and U13018 (N_13018,N_6107,N_8102);
and U13019 (N_13019,N_9741,N_6512);
xor U13020 (N_13020,N_6843,N_5453);
and U13021 (N_13021,N_5812,N_5238);
or U13022 (N_13022,N_8164,N_5046);
nand U13023 (N_13023,N_5949,N_6744);
and U13024 (N_13024,N_6470,N_6062);
and U13025 (N_13025,N_9793,N_6226);
nand U13026 (N_13026,N_5650,N_6181);
xor U13027 (N_13027,N_9396,N_9197);
xor U13028 (N_13028,N_5247,N_6181);
and U13029 (N_13029,N_7885,N_8745);
xor U13030 (N_13030,N_7435,N_9112);
nor U13031 (N_13031,N_6886,N_9002);
or U13032 (N_13032,N_7746,N_7029);
or U13033 (N_13033,N_5443,N_6906);
or U13034 (N_13034,N_6087,N_8768);
nor U13035 (N_13035,N_9451,N_6823);
or U13036 (N_13036,N_9060,N_5703);
nor U13037 (N_13037,N_9189,N_7703);
and U13038 (N_13038,N_9898,N_9663);
and U13039 (N_13039,N_5161,N_8000);
nor U13040 (N_13040,N_9464,N_9766);
and U13041 (N_13041,N_5110,N_8141);
xnor U13042 (N_13042,N_8987,N_9176);
nor U13043 (N_13043,N_5326,N_7737);
or U13044 (N_13044,N_9007,N_7016);
xnor U13045 (N_13045,N_8656,N_7597);
and U13046 (N_13046,N_5298,N_7945);
xor U13047 (N_13047,N_7406,N_7423);
nand U13048 (N_13048,N_5380,N_7390);
or U13049 (N_13049,N_8779,N_6396);
nand U13050 (N_13050,N_9087,N_6727);
xor U13051 (N_13051,N_9044,N_7841);
xor U13052 (N_13052,N_7760,N_9874);
nand U13053 (N_13053,N_8388,N_6517);
xnor U13054 (N_13054,N_5031,N_6906);
xnor U13055 (N_13055,N_8409,N_8414);
or U13056 (N_13056,N_9595,N_5253);
nand U13057 (N_13057,N_7313,N_9335);
and U13058 (N_13058,N_9878,N_9704);
and U13059 (N_13059,N_8811,N_7063);
nand U13060 (N_13060,N_8739,N_9708);
xnor U13061 (N_13061,N_6764,N_7579);
xnor U13062 (N_13062,N_6167,N_7051);
nor U13063 (N_13063,N_7937,N_9344);
xor U13064 (N_13064,N_8489,N_7444);
nor U13065 (N_13065,N_7335,N_5422);
nor U13066 (N_13066,N_9734,N_7915);
or U13067 (N_13067,N_9357,N_7046);
and U13068 (N_13068,N_6748,N_8714);
nor U13069 (N_13069,N_9336,N_6976);
and U13070 (N_13070,N_8917,N_8541);
nor U13071 (N_13071,N_9721,N_8157);
and U13072 (N_13072,N_9763,N_7003);
nor U13073 (N_13073,N_5267,N_7539);
xnor U13074 (N_13074,N_8547,N_5946);
and U13075 (N_13075,N_8240,N_5874);
nor U13076 (N_13076,N_5938,N_7624);
xnor U13077 (N_13077,N_9755,N_9959);
xnor U13078 (N_13078,N_8746,N_9153);
or U13079 (N_13079,N_8433,N_8471);
nor U13080 (N_13080,N_8066,N_9210);
or U13081 (N_13081,N_8502,N_5687);
xor U13082 (N_13082,N_8299,N_8604);
and U13083 (N_13083,N_7503,N_9483);
nand U13084 (N_13084,N_9989,N_8707);
xor U13085 (N_13085,N_9955,N_9360);
and U13086 (N_13086,N_9300,N_5797);
nor U13087 (N_13087,N_7674,N_9849);
nand U13088 (N_13088,N_5677,N_6259);
nand U13089 (N_13089,N_8337,N_5263);
nor U13090 (N_13090,N_8634,N_5501);
nor U13091 (N_13091,N_5042,N_6719);
xnor U13092 (N_13092,N_6780,N_7196);
or U13093 (N_13093,N_6820,N_8495);
xnor U13094 (N_13094,N_5483,N_8969);
or U13095 (N_13095,N_6449,N_7170);
and U13096 (N_13096,N_9689,N_6346);
nor U13097 (N_13097,N_7522,N_5455);
and U13098 (N_13098,N_7606,N_5936);
and U13099 (N_13099,N_8057,N_9674);
and U13100 (N_13100,N_7360,N_9495);
nor U13101 (N_13101,N_7800,N_6799);
nand U13102 (N_13102,N_9730,N_6299);
or U13103 (N_13103,N_5439,N_5950);
or U13104 (N_13104,N_8269,N_8926);
nor U13105 (N_13105,N_5019,N_5989);
nand U13106 (N_13106,N_8285,N_6968);
and U13107 (N_13107,N_5428,N_7093);
nor U13108 (N_13108,N_8777,N_8743);
and U13109 (N_13109,N_7942,N_8445);
or U13110 (N_13110,N_6220,N_5853);
nor U13111 (N_13111,N_6977,N_7166);
nor U13112 (N_13112,N_9305,N_7377);
or U13113 (N_13113,N_9520,N_6947);
nand U13114 (N_13114,N_7689,N_9529);
xnor U13115 (N_13115,N_7180,N_8750);
or U13116 (N_13116,N_8802,N_5959);
xnor U13117 (N_13117,N_9853,N_8394);
nor U13118 (N_13118,N_7185,N_9663);
or U13119 (N_13119,N_8164,N_7033);
nor U13120 (N_13120,N_5989,N_8312);
or U13121 (N_13121,N_7296,N_7056);
nand U13122 (N_13122,N_5063,N_7608);
or U13123 (N_13123,N_6322,N_7795);
and U13124 (N_13124,N_7121,N_7115);
nor U13125 (N_13125,N_7907,N_7320);
or U13126 (N_13126,N_6344,N_8936);
and U13127 (N_13127,N_7474,N_5872);
nor U13128 (N_13128,N_6475,N_9909);
or U13129 (N_13129,N_9556,N_5848);
nor U13130 (N_13130,N_5752,N_6444);
nand U13131 (N_13131,N_8229,N_6259);
or U13132 (N_13132,N_7418,N_6487);
nand U13133 (N_13133,N_7105,N_9233);
nor U13134 (N_13134,N_5722,N_6160);
or U13135 (N_13135,N_9989,N_6734);
nand U13136 (N_13136,N_8288,N_9235);
nand U13137 (N_13137,N_5517,N_7053);
or U13138 (N_13138,N_9892,N_8290);
or U13139 (N_13139,N_6395,N_6353);
or U13140 (N_13140,N_6876,N_5217);
or U13141 (N_13141,N_7174,N_7273);
and U13142 (N_13142,N_5679,N_8078);
or U13143 (N_13143,N_6888,N_6079);
nand U13144 (N_13144,N_6795,N_8527);
and U13145 (N_13145,N_7857,N_5790);
or U13146 (N_13146,N_9878,N_5214);
or U13147 (N_13147,N_5786,N_7122);
xnor U13148 (N_13148,N_5242,N_5904);
nand U13149 (N_13149,N_8492,N_7067);
nand U13150 (N_13150,N_9735,N_8460);
and U13151 (N_13151,N_9899,N_6254);
nand U13152 (N_13152,N_7777,N_8510);
nand U13153 (N_13153,N_6508,N_8647);
and U13154 (N_13154,N_5590,N_5253);
nand U13155 (N_13155,N_8108,N_8203);
xnor U13156 (N_13156,N_5901,N_8793);
nand U13157 (N_13157,N_6608,N_6560);
or U13158 (N_13158,N_7333,N_5694);
nand U13159 (N_13159,N_8616,N_7037);
nand U13160 (N_13160,N_5567,N_9028);
or U13161 (N_13161,N_7343,N_7548);
or U13162 (N_13162,N_7264,N_5290);
nand U13163 (N_13163,N_6451,N_6510);
xor U13164 (N_13164,N_6150,N_6462);
xnor U13165 (N_13165,N_5293,N_9802);
nand U13166 (N_13166,N_9961,N_9585);
nor U13167 (N_13167,N_6559,N_8084);
xnor U13168 (N_13168,N_6504,N_7056);
and U13169 (N_13169,N_8794,N_6042);
nand U13170 (N_13170,N_9471,N_6746);
or U13171 (N_13171,N_5800,N_9172);
nor U13172 (N_13172,N_5266,N_5652);
and U13173 (N_13173,N_5121,N_7061);
or U13174 (N_13174,N_7120,N_8490);
and U13175 (N_13175,N_7545,N_6855);
nor U13176 (N_13176,N_8195,N_9077);
and U13177 (N_13177,N_8805,N_7914);
and U13178 (N_13178,N_6773,N_8803);
and U13179 (N_13179,N_9366,N_5941);
and U13180 (N_13180,N_7247,N_8211);
xnor U13181 (N_13181,N_6445,N_8166);
or U13182 (N_13182,N_5504,N_7404);
or U13183 (N_13183,N_5081,N_6272);
nand U13184 (N_13184,N_9130,N_5169);
or U13185 (N_13185,N_9733,N_5269);
nor U13186 (N_13186,N_6194,N_6286);
nor U13187 (N_13187,N_5430,N_8231);
nand U13188 (N_13188,N_9477,N_7286);
nand U13189 (N_13189,N_9924,N_6576);
or U13190 (N_13190,N_5320,N_8471);
nand U13191 (N_13191,N_6736,N_5919);
nand U13192 (N_13192,N_7319,N_7463);
xnor U13193 (N_13193,N_7809,N_7592);
nand U13194 (N_13194,N_7291,N_6274);
or U13195 (N_13195,N_7696,N_6188);
nand U13196 (N_13196,N_6525,N_8037);
nor U13197 (N_13197,N_9483,N_8755);
or U13198 (N_13198,N_7405,N_8599);
and U13199 (N_13199,N_7983,N_7306);
nand U13200 (N_13200,N_6891,N_6955);
nand U13201 (N_13201,N_5795,N_5034);
or U13202 (N_13202,N_5805,N_5771);
and U13203 (N_13203,N_5523,N_6859);
nor U13204 (N_13204,N_8463,N_7631);
or U13205 (N_13205,N_7220,N_6110);
and U13206 (N_13206,N_7389,N_5108);
nand U13207 (N_13207,N_6157,N_8438);
nand U13208 (N_13208,N_8503,N_7019);
nand U13209 (N_13209,N_7808,N_8836);
or U13210 (N_13210,N_8477,N_9636);
or U13211 (N_13211,N_6536,N_9805);
nor U13212 (N_13212,N_8230,N_9401);
or U13213 (N_13213,N_6999,N_6290);
nor U13214 (N_13214,N_8224,N_6848);
or U13215 (N_13215,N_6175,N_8978);
xnor U13216 (N_13216,N_8196,N_7776);
and U13217 (N_13217,N_7491,N_8977);
or U13218 (N_13218,N_7295,N_9522);
xor U13219 (N_13219,N_6359,N_9933);
nor U13220 (N_13220,N_8940,N_9280);
nand U13221 (N_13221,N_8663,N_8347);
or U13222 (N_13222,N_7803,N_8824);
or U13223 (N_13223,N_7945,N_9330);
and U13224 (N_13224,N_7260,N_8245);
or U13225 (N_13225,N_5034,N_7844);
xnor U13226 (N_13226,N_5942,N_8540);
nor U13227 (N_13227,N_5270,N_9961);
or U13228 (N_13228,N_9462,N_7929);
or U13229 (N_13229,N_5405,N_9504);
nor U13230 (N_13230,N_5142,N_8340);
xor U13231 (N_13231,N_8837,N_9400);
nand U13232 (N_13232,N_9758,N_6845);
nand U13233 (N_13233,N_8582,N_5221);
nor U13234 (N_13234,N_9410,N_7972);
nand U13235 (N_13235,N_6120,N_7028);
nor U13236 (N_13236,N_8377,N_7874);
xor U13237 (N_13237,N_5261,N_9102);
and U13238 (N_13238,N_7285,N_9504);
nand U13239 (N_13239,N_5108,N_9837);
and U13240 (N_13240,N_7803,N_7203);
or U13241 (N_13241,N_6234,N_7766);
nor U13242 (N_13242,N_6113,N_5081);
xor U13243 (N_13243,N_7816,N_7469);
nand U13244 (N_13244,N_5080,N_7605);
nor U13245 (N_13245,N_9040,N_9604);
and U13246 (N_13246,N_9913,N_7801);
or U13247 (N_13247,N_5515,N_8322);
or U13248 (N_13248,N_7244,N_7821);
and U13249 (N_13249,N_5018,N_9266);
and U13250 (N_13250,N_9083,N_8256);
xor U13251 (N_13251,N_9481,N_5544);
nor U13252 (N_13252,N_7950,N_7669);
nand U13253 (N_13253,N_7516,N_9888);
xnor U13254 (N_13254,N_8739,N_7188);
and U13255 (N_13255,N_6259,N_6657);
nand U13256 (N_13256,N_9700,N_6838);
or U13257 (N_13257,N_9967,N_8262);
nand U13258 (N_13258,N_8927,N_5057);
nor U13259 (N_13259,N_5972,N_7834);
nand U13260 (N_13260,N_6169,N_9246);
and U13261 (N_13261,N_6011,N_7695);
and U13262 (N_13262,N_7178,N_6478);
and U13263 (N_13263,N_6925,N_8318);
nand U13264 (N_13264,N_9292,N_7385);
or U13265 (N_13265,N_7223,N_5641);
and U13266 (N_13266,N_7288,N_6226);
xnor U13267 (N_13267,N_8843,N_8526);
nor U13268 (N_13268,N_5294,N_8694);
nor U13269 (N_13269,N_8300,N_6006);
nor U13270 (N_13270,N_6315,N_9692);
or U13271 (N_13271,N_9283,N_9046);
xor U13272 (N_13272,N_9324,N_6267);
and U13273 (N_13273,N_7402,N_6768);
nor U13274 (N_13274,N_5663,N_5755);
nand U13275 (N_13275,N_9453,N_9012);
nor U13276 (N_13276,N_8266,N_7276);
and U13277 (N_13277,N_5624,N_8359);
nor U13278 (N_13278,N_5863,N_8982);
nor U13279 (N_13279,N_8663,N_5032);
xnor U13280 (N_13280,N_9828,N_7617);
or U13281 (N_13281,N_9949,N_9290);
and U13282 (N_13282,N_6810,N_8410);
or U13283 (N_13283,N_7829,N_5535);
nor U13284 (N_13284,N_8474,N_6734);
nand U13285 (N_13285,N_8299,N_6060);
or U13286 (N_13286,N_9954,N_5690);
nand U13287 (N_13287,N_5950,N_6829);
xor U13288 (N_13288,N_7100,N_8523);
and U13289 (N_13289,N_9420,N_7325);
nor U13290 (N_13290,N_8997,N_5933);
xor U13291 (N_13291,N_8625,N_5942);
nand U13292 (N_13292,N_7611,N_9298);
or U13293 (N_13293,N_7087,N_7654);
xnor U13294 (N_13294,N_7649,N_6390);
nor U13295 (N_13295,N_8486,N_6353);
nand U13296 (N_13296,N_6510,N_8423);
nand U13297 (N_13297,N_6093,N_5557);
nand U13298 (N_13298,N_8240,N_6341);
nor U13299 (N_13299,N_9588,N_8347);
xnor U13300 (N_13300,N_9613,N_6408);
and U13301 (N_13301,N_6373,N_6981);
nor U13302 (N_13302,N_9789,N_6890);
nor U13303 (N_13303,N_5595,N_9297);
and U13304 (N_13304,N_5412,N_8389);
nand U13305 (N_13305,N_6055,N_7473);
and U13306 (N_13306,N_6189,N_8765);
xnor U13307 (N_13307,N_7760,N_7192);
and U13308 (N_13308,N_9426,N_6060);
xor U13309 (N_13309,N_8342,N_9449);
or U13310 (N_13310,N_7805,N_8874);
nor U13311 (N_13311,N_7366,N_5974);
xnor U13312 (N_13312,N_9781,N_8603);
nor U13313 (N_13313,N_7774,N_6557);
xor U13314 (N_13314,N_5587,N_9240);
nor U13315 (N_13315,N_5627,N_9773);
and U13316 (N_13316,N_6202,N_8833);
and U13317 (N_13317,N_5557,N_8480);
xnor U13318 (N_13318,N_6646,N_6943);
nor U13319 (N_13319,N_9258,N_6233);
nand U13320 (N_13320,N_8442,N_5050);
nand U13321 (N_13321,N_7419,N_9579);
nand U13322 (N_13322,N_8052,N_9504);
nand U13323 (N_13323,N_6167,N_6101);
xor U13324 (N_13324,N_6154,N_6148);
or U13325 (N_13325,N_9832,N_8458);
nor U13326 (N_13326,N_6971,N_5976);
nor U13327 (N_13327,N_6990,N_8609);
or U13328 (N_13328,N_5799,N_8551);
nand U13329 (N_13329,N_6563,N_8382);
xnor U13330 (N_13330,N_6785,N_5597);
nand U13331 (N_13331,N_5778,N_7099);
or U13332 (N_13332,N_8564,N_6035);
xor U13333 (N_13333,N_7094,N_8484);
xnor U13334 (N_13334,N_8561,N_9048);
xor U13335 (N_13335,N_5377,N_7745);
xor U13336 (N_13336,N_8344,N_6025);
nor U13337 (N_13337,N_7434,N_9926);
and U13338 (N_13338,N_6888,N_8204);
or U13339 (N_13339,N_8805,N_6410);
xor U13340 (N_13340,N_9752,N_9204);
nand U13341 (N_13341,N_8762,N_7532);
nor U13342 (N_13342,N_9272,N_5903);
and U13343 (N_13343,N_5491,N_5899);
nand U13344 (N_13344,N_9717,N_7185);
nor U13345 (N_13345,N_8196,N_8296);
nand U13346 (N_13346,N_7939,N_7387);
or U13347 (N_13347,N_5251,N_7093);
or U13348 (N_13348,N_7509,N_8005);
and U13349 (N_13349,N_9166,N_5437);
xor U13350 (N_13350,N_6858,N_7597);
and U13351 (N_13351,N_7367,N_9164);
nand U13352 (N_13352,N_7799,N_9896);
nor U13353 (N_13353,N_7813,N_5013);
nand U13354 (N_13354,N_7299,N_7954);
or U13355 (N_13355,N_5130,N_5631);
nand U13356 (N_13356,N_5486,N_7436);
xnor U13357 (N_13357,N_8891,N_9611);
nor U13358 (N_13358,N_6651,N_5889);
and U13359 (N_13359,N_9821,N_7411);
or U13360 (N_13360,N_5010,N_5914);
nor U13361 (N_13361,N_8553,N_9562);
or U13362 (N_13362,N_8372,N_5375);
and U13363 (N_13363,N_5466,N_5310);
nor U13364 (N_13364,N_6166,N_6301);
nor U13365 (N_13365,N_9010,N_9038);
or U13366 (N_13366,N_6239,N_6782);
xor U13367 (N_13367,N_9940,N_7126);
xor U13368 (N_13368,N_9010,N_8429);
nand U13369 (N_13369,N_6761,N_6812);
and U13370 (N_13370,N_6883,N_5821);
or U13371 (N_13371,N_7735,N_5847);
nand U13372 (N_13372,N_8433,N_6200);
nand U13373 (N_13373,N_6565,N_9460);
nor U13374 (N_13374,N_8855,N_6502);
xor U13375 (N_13375,N_5349,N_6105);
nand U13376 (N_13376,N_7131,N_7697);
and U13377 (N_13377,N_8022,N_7244);
nor U13378 (N_13378,N_8867,N_6066);
nor U13379 (N_13379,N_5366,N_8349);
or U13380 (N_13380,N_7183,N_8553);
or U13381 (N_13381,N_6029,N_5962);
and U13382 (N_13382,N_9901,N_9546);
nand U13383 (N_13383,N_9391,N_7834);
nor U13384 (N_13384,N_6044,N_9875);
xor U13385 (N_13385,N_9044,N_7167);
nand U13386 (N_13386,N_6396,N_6885);
nor U13387 (N_13387,N_5509,N_6946);
xnor U13388 (N_13388,N_8206,N_7926);
or U13389 (N_13389,N_9684,N_8261);
and U13390 (N_13390,N_6274,N_9892);
and U13391 (N_13391,N_6915,N_8749);
nand U13392 (N_13392,N_5840,N_5977);
nand U13393 (N_13393,N_7802,N_6065);
xnor U13394 (N_13394,N_9576,N_8157);
xor U13395 (N_13395,N_5332,N_5235);
nand U13396 (N_13396,N_6007,N_9669);
nand U13397 (N_13397,N_8308,N_8907);
and U13398 (N_13398,N_9834,N_5574);
nand U13399 (N_13399,N_7769,N_5585);
nor U13400 (N_13400,N_6299,N_5942);
and U13401 (N_13401,N_7333,N_9397);
nand U13402 (N_13402,N_8211,N_5530);
or U13403 (N_13403,N_8389,N_5606);
or U13404 (N_13404,N_6624,N_9071);
nor U13405 (N_13405,N_9500,N_7408);
xnor U13406 (N_13406,N_5177,N_6470);
and U13407 (N_13407,N_9777,N_7624);
xor U13408 (N_13408,N_6898,N_7138);
nand U13409 (N_13409,N_5326,N_9459);
and U13410 (N_13410,N_7937,N_6194);
xnor U13411 (N_13411,N_6384,N_6821);
nand U13412 (N_13412,N_9650,N_9896);
nand U13413 (N_13413,N_8921,N_5278);
nand U13414 (N_13414,N_5331,N_7838);
nor U13415 (N_13415,N_7146,N_7025);
nand U13416 (N_13416,N_8415,N_9819);
nor U13417 (N_13417,N_9785,N_7375);
and U13418 (N_13418,N_9082,N_6703);
nand U13419 (N_13419,N_7760,N_5392);
or U13420 (N_13420,N_5252,N_6122);
nand U13421 (N_13421,N_9257,N_9425);
xor U13422 (N_13422,N_5579,N_7016);
and U13423 (N_13423,N_5685,N_9269);
xor U13424 (N_13424,N_8127,N_8651);
and U13425 (N_13425,N_7923,N_5994);
nand U13426 (N_13426,N_7942,N_7503);
nor U13427 (N_13427,N_7502,N_5470);
and U13428 (N_13428,N_9752,N_6750);
nand U13429 (N_13429,N_9196,N_9504);
or U13430 (N_13430,N_8530,N_9751);
and U13431 (N_13431,N_6699,N_8994);
nand U13432 (N_13432,N_9983,N_6214);
or U13433 (N_13433,N_8305,N_7476);
nand U13434 (N_13434,N_5104,N_9998);
and U13435 (N_13435,N_6353,N_9928);
and U13436 (N_13436,N_7013,N_6504);
nor U13437 (N_13437,N_8802,N_5541);
and U13438 (N_13438,N_6657,N_8246);
or U13439 (N_13439,N_7113,N_5407);
nand U13440 (N_13440,N_9099,N_9106);
xor U13441 (N_13441,N_9622,N_5106);
xnor U13442 (N_13442,N_9244,N_7478);
xor U13443 (N_13443,N_7747,N_9023);
nor U13444 (N_13444,N_5831,N_8371);
or U13445 (N_13445,N_8324,N_6862);
or U13446 (N_13446,N_8736,N_5050);
nand U13447 (N_13447,N_7980,N_5635);
xnor U13448 (N_13448,N_6797,N_9944);
xor U13449 (N_13449,N_6168,N_5845);
nand U13450 (N_13450,N_5043,N_7262);
and U13451 (N_13451,N_7787,N_6758);
nor U13452 (N_13452,N_8392,N_8124);
and U13453 (N_13453,N_8379,N_6805);
xnor U13454 (N_13454,N_7748,N_6581);
nor U13455 (N_13455,N_8680,N_9071);
nand U13456 (N_13456,N_5466,N_5584);
xnor U13457 (N_13457,N_8192,N_8297);
and U13458 (N_13458,N_7543,N_5893);
and U13459 (N_13459,N_9987,N_6763);
nor U13460 (N_13460,N_8774,N_5159);
xnor U13461 (N_13461,N_9242,N_5420);
nand U13462 (N_13462,N_9326,N_6151);
nand U13463 (N_13463,N_6042,N_6564);
nor U13464 (N_13464,N_9729,N_7266);
nor U13465 (N_13465,N_7445,N_7888);
xor U13466 (N_13466,N_7925,N_8111);
nor U13467 (N_13467,N_9968,N_9855);
xnor U13468 (N_13468,N_9891,N_9602);
and U13469 (N_13469,N_7480,N_8887);
nor U13470 (N_13470,N_5471,N_7859);
nand U13471 (N_13471,N_6170,N_6835);
and U13472 (N_13472,N_6939,N_8403);
xor U13473 (N_13473,N_8744,N_6269);
nand U13474 (N_13474,N_7931,N_7276);
and U13475 (N_13475,N_9752,N_5546);
or U13476 (N_13476,N_6206,N_8355);
nor U13477 (N_13477,N_6907,N_6182);
nand U13478 (N_13478,N_6179,N_8731);
xnor U13479 (N_13479,N_8113,N_9097);
nor U13480 (N_13480,N_8025,N_7529);
or U13481 (N_13481,N_7322,N_7749);
nor U13482 (N_13482,N_6459,N_5635);
or U13483 (N_13483,N_6327,N_6951);
or U13484 (N_13484,N_7250,N_6477);
or U13485 (N_13485,N_6246,N_7591);
nor U13486 (N_13486,N_9069,N_9760);
nor U13487 (N_13487,N_9645,N_6044);
and U13488 (N_13488,N_6029,N_8569);
xnor U13489 (N_13489,N_7990,N_9595);
nand U13490 (N_13490,N_8779,N_6546);
nor U13491 (N_13491,N_9973,N_8742);
or U13492 (N_13492,N_5957,N_8235);
and U13493 (N_13493,N_6771,N_5109);
nand U13494 (N_13494,N_7063,N_7373);
nor U13495 (N_13495,N_6048,N_7232);
and U13496 (N_13496,N_9173,N_9977);
or U13497 (N_13497,N_7392,N_8932);
nand U13498 (N_13498,N_9018,N_7227);
xnor U13499 (N_13499,N_8593,N_7319);
and U13500 (N_13500,N_9921,N_6034);
nor U13501 (N_13501,N_9390,N_8603);
or U13502 (N_13502,N_9109,N_5667);
nor U13503 (N_13503,N_5444,N_5610);
and U13504 (N_13504,N_6075,N_6011);
nor U13505 (N_13505,N_6951,N_9778);
nand U13506 (N_13506,N_5423,N_6531);
nand U13507 (N_13507,N_5579,N_7117);
nor U13508 (N_13508,N_8258,N_9457);
nor U13509 (N_13509,N_5476,N_5578);
nor U13510 (N_13510,N_7133,N_9450);
nand U13511 (N_13511,N_6251,N_7715);
nand U13512 (N_13512,N_5054,N_6931);
nand U13513 (N_13513,N_5049,N_8337);
and U13514 (N_13514,N_8925,N_6412);
or U13515 (N_13515,N_9667,N_8155);
nor U13516 (N_13516,N_5033,N_8636);
and U13517 (N_13517,N_6699,N_5092);
or U13518 (N_13518,N_6445,N_7939);
nand U13519 (N_13519,N_5590,N_7284);
or U13520 (N_13520,N_7367,N_9014);
or U13521 (N_13521,N_7873,N_6530);
xor U13522 (N_13522,N_9893,N_7771);
and U13523 (N_13523,N_6053,N_7746);
xor U13524 (N_13524,N_6329,N_5406);
and U13525 (N_13525,N_7968,N_5195);
and U13526 (N_13526,N_6487,N_8796);
or U13527 (N_13527,N_9249,N_9889);
and U13528 (N_13528,N_9826,N_6253);
nor U13529 (N_13529,N_7123,N_6843);
and U13530 (N_13530,N_8537,N_9374);
nand U13531 (N_13531,N_9086,N_8572);
nand U13532 (N_13532,N_9052,N_8384);
nor U13533 (N_13533,N_9650,N_6600);
or U13534 (N_13534,N_5715,N_6028);
nand U13535 (N_13535,N_5947,N_6839);
or U13536 (N_13536,N_7259,N_6876);
and U13537 (N_13537,N_6813,N_9887);
nor U13538 (N_13538,N_8990,N_9319);
nand U13539 (N_13539,N_5441,N_5833);
xnor U13540 (N_13540,N_8835,N_8471);
nand U13541 (N_13541,N_5303,N_7939);
or U13542 (N_13542,N_9307,N_6160);
xor U13543 (N_13543,N_5438,N_7281);
nand U13544 (N_13544,N_7871,N_5548);
and U13545 (N_13545,N_7405,N_6929);
nand U13546 (N_13546,N_5762,N_7348);
xnor U13547 (N_13547,N_5369,N_5241);
nand U13548 (N_13548,N_8919,N_9015);
or U13549 (N_13549,N_9574,N_8565);
xor U13550 (N_13550,N_7357,N_8007);
nand U13551 (N_13551,N_5021,N_5211);
or U13552 (N_13552,N_7465,N_5810);
or U13553 (N_13553,N_9024,N_9472);
nor U13554 (N_13554,N_7623,N_6620);
nor U13555 (N_13555,N_5761,N_5535);
or U13556 (N_13556,N_8731,N_9607);
and U13557 (N_13557,N_5971,N_8536);
and U13558 (N_13558,N_6107,N_9175);
or U13559 (N_13559,N_6981,N_8597);
or U13560 (N_13560,N_9398,N_6407);
and U13561 (N_13561,N_7692,N_7139);
xnor U13562 (N_13562,N_9502,N_9058);
or U13563 (N_13563,N_8863,N_5035);
and U13564 (N_13564,N_7008,N_7987);
nand U13565 (N_13565,N_5318,N_6944);
nand U13566 (N_13566,N_7508,N_8288);
or U13567 (N_13567,N_8730,N_6087);
or U13568 (N_13568,N_5716,N_7689);
xnor U13569 (N_13569,N_8868,N_9489);
nor U13570 (N_13570,N_5768,N_6384);
xnor U13571 (N_13571,N_7981,N_6662);
nor U13572 (N_13572,N_6718,N_9334);
nand U13573 (N_13573,N_7556,N_6699);
nand U13574 (N_13574,N_6545,N_6216);
xnor U13575 (N_13575,N_9641,N_5399);
nand U13576 (N_13576,N_8264,N_7365);
or U13577 (N_13577,N_7042,N_8768);
or U13578 (N_13578,N_9026,N_9158);
nor U13579 (N_13579,N_8110,N_9906);
xnor U13580 (N_13580,N_8620,N_5673);
nor U13581 (N_13581,N_7986,N_7615);
nor U13582 (N_13582,N_7952,N_8701);
xnor U13583 (N_13583,N_9540,N_8753);
or U13584 (N_13584,N_5672,N_9805);
or U13585 (N_13585,N_8896,N_7074);
or U13586 (N_13586,N_6212,N_5731);
nand U13587 (N_13587,N_7209,N_9502);
or U13588 (N_13588,N_7584,N_6663);
nand U13589 (N_13589,N_7291,N_9100);
xnor U13590 (N_13590,N_6699,N_6556);
xor U13591 (N_13591,N_5249,N_7902);
and U13592 (N_13592,N_5003,N_6820);
or U13593 (N_13593,N_6540,N_8552);
nor U13594 (N_13594,N_6942,N_6852);
nand U13595 (N_13595,N_6257,N_7054);
nor U13596 (N_13596,N_9037,N_9588);
and U13597 (N_13597,N_5803,N_6864);
xor U13598 (N_13598,N_6937,N_5663);
xnor U13599 (N_13599,N_7647,N_6987);
xnor U13600 (N_13600,N_8175,N_9641);
and U13601 (N_13601,N_6134,N_6853);
nor U13602 (N_13602,N_6240,N_8926);
xor U13603 (N_13603,N_9343,N_8623);
nor U13604 (N_13604,N_7655,N_8449);
or U13605 (N_13605,N_7379,N_9078);
nor U13606 (N_13606,N_5277,N_8301);
or U13607 (N_13607,N_9515,N_6507);
and U13608 (N_13608,N_5945,N_9251);
xor U13609 (N_13609,N_7539,N_7029);
and U13610 (N_13610,N_6486,N_7051);
xor U13611 (N_13611,N_8702,N_9236);
nor U13612 (N_13612,N_8336,N_8330);
or U13613 (N_13613,N_7611,N_5018);
nor U13614 (N_13614,N_6779,N_9514);
xor U13615 (N_13615,N_8514,N_5971);
and U13616 (N_13616,N_9373,N_7852);
and U13617 (N_13617,N_6254,N_6167);
xor U13618 (N_13618,N_9810,N_6555);
xor U13619 (N_13619,N_5969,N_5464);
and U13620 (N_13620,N_9604,N_5747);
xnor U13621 (N_13621,N_6237,N_7284);
and U13622 (N_13622,N_8265,N_8272);
nand U13623 (N_13623,N_6879,N_6131);
nor U13624 (N_13624,N_7084,N_7153);
and U13625 (N_13625,N_7666,N_6459);
xnor U13626 (N_13626,N_5320,N_7938);
or U13627 (N_13627,N_8828,N_7237);
or U13628 (N_13628,N_7781,N_9082);
and U13629 (N_13629,N_5902,N_6640);
or U13630 (N_13630,N_5303,N_6953);
xor U13631 (N_13631,N_9027,N_6661);
nand U13632 (N_13632,N_7002,N_5166);
xnor U13633 (N_13633,N_9814,N_6239);
or U13634 (N_13634,N_9751,N_8339);
and U13635 (N_13635,N_7519,N_5764);
nand U13636 (N_13636,N_9792,N_7059);
and U13637 (N_13637,N_5888,N_5941);
xor U13638 (N_13638,N_9608,N_5555);
xor U13639 (N_13639,N_8892,N_9649);
or U13640 (N_13640,N_9838,N_9355);
xor U13641 (N_13641,N_6568,N_5176);
nand U13642 (N_13642,N_7254,N_8672);
nor U13643 (N_13643,N_8688,N_7132);
nand U13644 (N_13644,N_6867,N_5103);
xnor U13645 (N_13645,N_8743,N_9666);
and U13646 (N_13646,N_6281,N_6176);
nor U13647 (N_13647,N_5476,N_5316);
xnor U13648 (N_13648,N_9445,N_8459);
and U13649 (N_13649,N_6426,N_9055);
nor U13650 (N_13650,N_5647,N_5669);
nand U13651 (N_13651,N_7733,N_7136);
or U13652 (N_13652,N_8340,N_6091);
nor U13653 (N_13653,N_8454,N_8312);
nand U13654 (N_13654,N_6636,N_8330);
and U13655 (N_13655,N_8768,N_7370);
nor U13656 (N_13656,N_6602,N_8440);
and U13657 (N_13657,N_6499,N_9648);
nand U13658 (N_13658,N_5794,N_8580);
nand U13659 (N_13659,N_7648,N_7531);
nor U13660 (N_13660,N_5021,N_9345);
xor U13661 (N_13661,N_9914,N_7933);
and U13662 (N_13662,N_7658,N_8970);
nor U13663 (N_13663,N_7376,N_5268);
xor U13664 (N_13664,N_5588,N_9285);
xor U13665 (N_13665,N_6567,N_7466);
nand U13666 (N_13666,N_7705,N_5586);
or U13667 (N_13667,N_7854,N_5234);
xor U13668 (N_13668,N_8907,N_7785);
nand U13669 (N_13669,N_5950,N_9396);
and U13670 (N_13670,N_8777,N_8757);
nor U13671 (N_13671,N_9301,N_6537);
nand U13672 (N_13672,N_5889,N_7327);
xnor U13673 (N_13673,N_8891,N_8732);
xor U13674 (N_13674,N_7922,N_5154);
nand U13675 (N_13675,N_9675,N_9183);
nand U13676 (N_13676,N_8647,N_5864);
or U13677 (N_13677,N_6274,N_5226);
nand U13678 (N_13678,N_7689,N_8955);
and U13679 (N_13679,N_5160,N_6906);
and U13680 (N_13680,N_8311,N_5674);
or U13681 (N_13681,N_5316,N_8315);
or U13682 (N_13682,N_9716,N_5811);
nand U13683 (N_13683,N_8529,N_7815);
xnor U13684 (N_13684,N_5159,N_9280);
nor U13685 (N_13685,N_7762,N_8163);
nand U13686 (N_13686,N_8788,N_5028);
or U13687 (N_13687,N_9717,N_9458);
nor U13688 (N_13688,N_5823,N_9377);
and U13689 (N_13689,N_6139,N_5680);
nand U13690 (N_13690,N_7127,N_9264);
nor U13691 (N_13691,N_9209,N_6515);
nand U13692 (N_13692,N_6153,N_7045);
nand U13693 (N_13693,N_9639,N_5505);
xnor U13694 (N_13694,N_9419,N_6481);
or U13695 (N_13695,N_8011,N_7144);
nand U13696 (N_13696,N_7866,N_8489);
nor U13697 (N_13697,N_9424,N_8480);
nand U13698 (N_13698,N_5781,N_7460);
nor U13699 (N_13699,N_7783,N_7293);
nor U13700 (N_13700,N_6942,N_9941);
xnor U13701 (N_13701,N_8583,N_8554);
and U13702 (N_13702,N_8571,N_8984);
nand U13703 (N_13703,N_7976,N_8760);
nor U13704 (N_13704,N_9625,N_6873);
nor U13705 (N_13705,N_7833,N_7255);
nand U13706 (N_13706,N_8677,N_5228);
or U13707 (N_13707,N_7056,N_6953);
xnor U13708 (N_13708,N_7393,N_8780);
xnor U13709 (N_13709,N_7516,N_9621);
nor U13710 (N_13710,N_9151,N_5488);
and U13711 (N_13711,N_7940,N_7088);
xor U13712 (N_13712,N_5687,N_7326);
nor U13713 (N_13713,N_6845,N_8973);
xnor U13714 (N_13714,N_6102,N_5697);
or U13715 (N_13715,N_5805,N_5825);
nand U13716 (N_13716,N_9958,N_7395);
nand U13717 (N_13717,N_9040,N_5998);
nor U13718 (N_13718,N_7412,N_5975);
xor U13719 (N_13719,N_8597,N_7016);
and U13720 (N_13720,N_5903,N_5048);
xnor U13721 (N_13721,N_5241,N_9645);
or U13722 (N_13722,N_5999,N_5362);
nor U13723 (N_13723,N_6599,N_5200);
xor U13724 (N_13724,N_9192,N_7015);
nand U13725 (N_13725,N_5125,N_5873);
or U13726 (N_13726,N_7289,N_9948);
or U13727 (N_13727,N_6026,N_8430);
nor U13728 (N_13728,N_9396,N_8906);
nor U13729 (N_13729,N_9367,N_7824);
and U13730 (N_13730,N_9780,N_8658);
and U13731 (N_13731,N_5525,N_7717);
nand U13732 (N_13732,N_8641,N_7628);
nand U13733 (N_13733,N_5581,N_9284);
xnor U13734 (N_13734,N_9748,N_5782);
and U13735 (N_13735,N_5180,N_7322);
and U13736 (N_13736,N_8487,N_9233);
nor U13737 (N_13737,N_5609,N_6949);
or U13738 (N_13738,N_5854,N_6479);
and U13739 (N_13739,N_7939,N_6358);
nand U13740 (N_13740,N_5520,N_7745);
or U13741 (N_13741,N_5602,N_6663);
nand U13742 (N_13742,N_9162,N_7278);
and U13743 (N_13743,N_6630,N_7520);
or U13744 (N_13744,N_9348,N_5145);
nor U13745 (N_13745,N_9184,N_5337);
xnor U13746 (N_13746,N_7450,N_9584);
nor U13747 (N_13747,N_9568,N_9043);
or U13748 (N_13748,N_7188,N_7577);
and U13749 (N_13749,N_6449,N_9327);
or U13750 (N_13750,N_5075,N_5469);
nand U13751 (N_13751,N_9953,N_9562);
and U13752 (N_13752,N_6915,N_8991);
nand U13753 (N_13753,N_9112,N_9927);
and U13754 (N_13754,N_8066,N_6243);
nor U13755 (N_13755,N_9471,N_6768);
and U13756 (N_13756,N_5512,N_9604);
nor U13757 (N_13757,N_7862,N_5817);
nor U13758 (N_13758,N_8683,N_7073);
or U13759 (N_13759,N_6349,N_7304);
and U13760 (N_13760,N_6861,N_7617);
and U13761 (N_13761,N_6778,N_8399);
xnor U13762 (N_13762,N_8781,N_6899);
nor U13763 (N_13763,N_6058,N_8251);
nand U13764 (N_13764,N_5051,N_6710);
or U13765 (N_13765,N_9758,N_9810);
nand U13766 (N_13766,N_7075,N_7310);
nand U13767 (N_13767,N_5007,N_9650);
xnor U13768 (N_13768,N_8343,N_7577);
and U13769 (N_13769,N_8512,N_9635);
nand U13770 (N_13770,N_6131,N_9715);
nor U13771 (N_13771,N_8799,N_9568);
or U13772 (N_13772,N_5641,N_8802);
xnor U13773 (N_13773,N_7758,N_5840);
nor U13774 (N_13774,N_7776,N_9533);
nor U13775 (N_13775,N_8588,N_9789);
nor U13776 (N_13776,N_5185,N_5276);
nor U13777 (N_13777,N_6749,N_5756);
nand U13778 (N_13778,N_9064,N_8674);
nand U13779 (N_13779,N_6579,N_5711);
nor U13780 (N_13780,N_5475,N_6073);
and U13781 (N_13781,N_5608,N_7486);
xor U13782 (N_13782,N_7428,N_6664);
or U13783 (N_13783,N_6440,N_8441);
and U13784 (N_13784,N_6465,N_6853);
nor U13785 (N_13785,N_9075,N_8328);
nand U13786 (N_13786,N_9076,N_9810);
nand U13787 (N_13787,N_6782,N_7009);
nor U13788 (N_13788,N_8253,N_8659);
nand U13789 (N_13789,N_6231,N_9407);
nand U13790 (N_13790,N_8826,N_8430);
nor U13791 (N_13791,N_6675,N_6352);
and U13792 (N_13792,N_5515,N_8149);
xor U13793 (N_13793,N_5684,N_7544);
nor U13794 (N_13794,N_5409,N_6375);
or U13795 (N_13795,N_5171,N_6602);
nand U13796 (N_13796,N_5497,N_9850);
xor U13797 (N_13797,N_9085,N_8815);
xor U13798 (N_13798,N_6062,N_6360);
and U13799 (N_13799,N_6683,N_8552);
xnor U13800 (N_13800,N_7860,N_5364);
xor U13801 (N_13801,N_5028,N_6548);
and U13802 (N_13802,N_9422,N_6501);
and U13803 (N_13803,N_7210,N_9798);
nor U13804 (N_13804,N_5441,N_9010);
nor U13805 (N_13805,N_8565,N_8218);
or U13806 (N_13806,N_9381,N_8427);
or U13807 (N_13807,N_5548,N_9175);
or U13808 (N_13808,N_5358,N_8977);
nand U13809 (N_13809,N_6586,N_8247);
and U13810 (N_13810,N_7022,N_7673);
and U13811 (N_13811,N_6298,N_6997);
nor U13812 (N_13812,N_5522,N_8429);
nand U13813 (N_13813,N_8951,N_6851);
xor U13814 (N_13814,N_5809,N_8994);
or U13815 (N_13815,N_5884,N_9679);
or U13816 (N_13816,N_6816,N_5396);
or U13817 (N_13817,N_8461,N_8799);
nand U13818 (N_13818,N_9105,N_6027);
or U13819 (N_13819,N_9065,N_8722);
xnor U13820 (N_13820,N_5935,N_8170);
xnor U13821 (N_13821,N_7152,N_6203);
or U13822 (N_13822,N_8822,N_5746);
xnor U13823 (N_13823,N_7621,N_6289);
or U13824 (N_13824,N_9731,N_8060);
nor U13825 (N_13825,N_5848,N_7680);
nor U13826 (N_13826,N_8765,N_9926);
nor U13827 (N_13827,N_8839,N_8841);
or U13828 (N_13828,N_7413,N_7695);
and U13829 (N_13829,N_7042,N_6162);
xnor U13830 (N_13830,N_5831,N_5504);
or U13831 (N_13831,N_6292,N_5400);
nand U13832 (N_13832,N_5422,N_9412);
xor U13833 (N_13833,N_7282,N_5513);
or U13834 (N_13834,N_9002,N_7824);
nor U13835 (N_13835,N_6384,N_6614);
or U13836 (N_13836,N_9860,N_7131);
xor U13837 (N_13837,N_6794,N_6132);
xor U13838 (N_13838,N_8601,N_9112);
and U13839 (N_13839,N_6064,N_5529);
nor U13840 (N_13840,N_8102,N_8936);
nand U13841 (N_13841,N_6298,N_8724);
or U13842 (N_13842,N_5431,N_9171);
and U13843 (N_13843,N_8685,N_7347);
xor U13844 (N_13844,N_8331,N_7360);
xnor U13845 (N_13845,N_9589,N_6037);
xnor U13846 (N_13846,N_7770,N_7733);
nor U13847 (N_13847,N_7923,N_5211);
nand U13848 (N_13848,N_7721,N_8692);
and U13849 (N_13849,N_9036,N_5532);
and U13850 (N_13850,N_9951,N_8218);
nand U13851 (N_13851,N_7476,N_7928);
xnor U13852 (N_13852,N_7834,N_9862);
or U13853 (N_13853,N_9152,N_9624);
and U13854 (N_13854,N_7365,N_5088);
xor U13855 (N_13855,N_8010,N_5738);
nand U13856 (N_13856,N_7500,N_8140);
or U13857 (N_13857,N_5778,N_9517);
nand U13858 (N_13858,N_8309,N_7808);
or U13859 (N_13859,N_9195,N_7505);
nand U13860 (N_13860,N_9547,N_6455);
nand U13861 (N_13861,N_6838,N_6807);
and U13862 (N_13862,N_8694,N_6483);
nor U13863 (N_13863,N_8491,N_7352);
nor U13864 (N_13864,N_8247,N_5998);
and U13865 (N_13865,N_7734,N_5330);
xnor U13866 (N_13866,N_6703,N_5954);
and U13867 (N_13867,N_9607,N_7889);
or U13868 (N_13868,N_7857,N_8031);
or U13869 (N_13869,N_8500,N_5052);
or U13870 (N_13870,N_9283,N_8322);
or U13871 (N_13871,N_6121,N_8214);
or U13872 (N_13872,N_9797,N_7064);
and U13873 (N_13873,N_6156,N_6554);
or U13874 (N_13874,N_9352,N_6563);
nand U13875 (N_13875,N_8825,N_5373);
nand U13876 (N_13876,N_5956,N_5601);
nor U13877 (N_13877,N_5674,N_7334);
nor U13878 (N_13878,N_7964,N_6711);
and U13879 (N_13879,N_7440,N_9579);
and U13880 (N_13880,N_9083,N_8082);
xnor U13881 (N_13881,N_9203,N_8366);
nand U13882 (N_13882,N_9644,N_9680);
or U13883 (N_13883,N_7704,N_9856);
nor U13884 (N_13884,N_8555,N_9897);
and U13885 (N_13885,N_5314,N_7550);
xor U13886 (N_13886,N_5894,N_6201);
nor U13887 (N_13887,N_9372,N_7277);
or U13888 (N_13888,N_7069,N_6805);
or U13889 (N_13889,N_6421,N_6095);
and U13890 (N_13890,N_8926,N_9044);
or U13891 (N_13891,N_7487,N_9057);
nor U13892 (N_13892,N_8595,N_7024);
and U13893 (N_13893,N_7177,N_9378);
xor U13894 (N_13894,N_9328,N_9523);
nand U13895 (N_13895,N_7605,N_9488);
or U13896 (N_13896,N_9514,N_8098);
nor U13897 (N_13897,N_8736,N_5773);
and U13898 (N_13898,N_5342,N_6300);
nor U13899 (N_13899,N_8220,N_7361);
or U13900 (N_13900,N_9918,N_5491);
nor U13901 (N_13901,N_9558,N_9132);
or U13902 (N_13902,N_7440,N_9953);
xor U13903 (N_13903,N_7104,N_7697);
xnor U13904 (N_13904,N_7781,N_5708);
xor U13905 (N_13905,N_7011,N_7152);
nor U13906 (N_13906,N_7783,N_8633);
nand U13907 (N_13907,N_5982,N_6514);
nor U13908 (N_13908,N_7801,N_9834);
or U13909 (N_13909,N_9092,N_8692);
nor U13910 (N_13910,N_9315,N_8663);
or U13911 (N_13911,N_9582,N_7679);
or U13912 (N_13912,N_8253,N_8655);
or U13913 (N_13913,N_6183,N_5806);
xor U13914 (N_13914,N_9996,N_9193);
and U13915 (N_13915,N_6296,N_9898);
nor U13916 (N_13916,N_5335,N_6613);
or U13917 (N_13917,N_7946,N_8120);
nor U13918 (N_13918,N_9779,N_9511);
nand U13919 (N_13919,N_8550,N_5986);
and U13920 (N_13920,N_7290,N_5672);
and U13921 (N_13921,N_8655,N_8051);
or U13922 (N_13922,N_8952,N_9008);
or U13923 (N_13923,N_5715,N_9092);
nor U13924 (N_13924,N_8777,N_9698);
and U13925 (N_13925,N_7032,N_9854);
or U13926 (N_13926,N_8084,N_9384);
and U13927 (N_13927,N_5054,N_6412);
or U13928 (N_13928,N_8778,N_7728);
nand U13929 (N_13929,N_8874,N_9712);
xnor U13930 (N_13930,N_5260,N_8734);
xnor U13931 (N_13931,N_9751,N_6604);
xnor U13932 (N_13932,N_8479,N_9368);
nor U13933 (N_13933,N_9913,N_5631);
or U13934 (N_13934,N_5203,N_7703);
nand U13935 (N_13935,N_9238,N_5447);
nor U13936 (N_13936,N_5965,N_8957);
nand U13937 (N_13937,N_6634,N_6530);
nor U13938 (N_13938,N_7535,N_9597);
nor U13939 (N_13939,N_9643,N_8066);
nor U13940 (N_13940,N_8710,N_6907);
or U13941 (N_13941,N_9856,N_5863);
and U13942 (N_13942,N_6489,N_6686);
and U13943 (N_13943,N_7967,N_8300);
nor U13944 (N_13944,N_9720,N_5150);
or U13945 (N_13945,N_9881,N_5800);
and U13946 (N_13946,N_9828,N_6707);
and U13947 (N_13947,N_8557,N_7823);
or U13948 (N_13948,N_9707,N_9571);
xnor U13949 (N_13949,N_7614,N_9752);
or U13950 (N_13950,N_8734,N_6133);
and U13951 (N_13951,N_9437,N_5022);
or U13952 (N_13952,N_9090,N_8035);
and U13953 (N_13953,N_8523,N_6538);
or U13954 (N_13954,N_6051,N_7484);
nand U13955 (N_13955,N_6632,N_6792);
xnor U13956 (N_13956,N_7974,N_5460);
xor U13957 (N_13957,N_7957,N_8794);
or U13958 (N_13958,N_8025,N_9364);
or U13959 (N_13959,N_9549,N_9956);
nor U13960 (N_13960,N_9900,N_7889);
or U13961 (N_13961,N_7094,N_9592);
nand U13962 (N_13962,N_6316,N_6383);
xnor U13963 (N_13963,N_7469,N_9591);
and U13964 (N_13964,N_8561,N_5182);
and U13965 (N_13965,N_7930,N_7670);
nor U13966 (N_13966,N_8586,N_8343);
or U13967 (N_13967,N_7581,N_7865);
nor U13968 (N_13968,N_7448,N_6965);
and U13969 (N_13969,N_9506,N_5920);
xnor U13970 (N_13970,N_6979,N_5933);
xnor U13971 (N_13971,N_8508,N_8400);
nor U13972 (N_13972,N_7969,N_9506);
and U13973 (N_13973,N_9180,N_5900);
or U13974 (N_13974,N_7928,N_9917);
xnor U13975 (N_13975,N_9057,N_7400);
and U13976 (N_13976,N_9557,N_7170);
nor U13977 (N_13977,N_7752,N_8952);
and U13978 (N_13978,N_8901,N_6922);
or U13979 (N_13979,N_5602,N_8289);
nor U13980 (N_13980,N_5460,N_7169);
nand U13981 (N_13981,N_5926,N_7482);
and U13982 (N_13982,N_7389,N_7812);
xnor U13983 (N_13983,N_9100,N_5229);
xnor U13984 (N_13984,N_9362,N_9255);
xor U13985 (N_13985,N_5020,N_8718);
or U13986 (N_13986,N_5869,N_8182);
or U13987 (N_13987,N_6747,N_5687);
xnor U13988 (N_13988,N_7899,N_8633);
nor U13989 (N_13989,N_7972,N_6261);
and U13990 (N_13990,N_8771,N_8996);
nor U13991 (N_13991,N_6475,N_5308);
nand U13992 (N_13992,N_6072,N_7039);
xnor U13993 (N_13993,N_7791,N_7669);
nand U13994 (N_13994,N_8082,N_8184);
nor U13995 (N_13995,N_5127,N_7599);
or U13996 (N_13996,N_9543,N_8348);
xnor U13997 (N_13997,N_8681,N_5473);
nand U13998 (N_13998,N_9281,N_6643);
nor U13999 (N_13999,N_6525,N_9316);
nor U14000 (N_14000,N_7452,N_9025);
and U14001 (N_14001,N_9493,N_5535);
nor U14002 (N_14002,N_8641,N_8817);
xor U14003 (N_14003,N_5976,N_6953);
xnor U14004 (N_14004,N_8015,N_6317);
xor U14005 (N_14005,N_8370,N_5903);
nor U14006 (N_14006,N_7595,N_6975);
nand U14007 (N_14007,N_5645,N_5064);
nor U14008 (N_14008,N_6494,N_5283);
or U14009 (N_14009,N_6048,N_9912);
xor U14010 (N_14010,N_5754,N_6469);
nand U14011 (N_14011,N_7161,N_9519);
nand U14012 (N_14012,N_8331,N_5043);
xnor U14013 (N_14013,N_8324,N_9405);
nand U14014 (N_14014,N_5340,N_7124);
and U14015 (N_14015,N_6342,N_9367);
xor U14016 (N_14016,N_9230,N_8671);
xnor U14017 (N_14017,N_7316,N_9199);
nor U14018 (N_14018,N_9411,N_9003);
or U14019 (N_14019,N_5121,N_6505);
nand U14020 (N_14020,N_7914,N_7661);
xnor U14021 (N_14021,N_8886,N_6727);
or U14022 (N_14022,N_6744,N_5720);
xnor U14023 (N_14023,N_9510,N_8075);
and U14024 (N_14024,N_9851,N_9795);
or U14025 (N_14025,N_9184,N_6488);
or U14026 (N_14026,N_6798,N_7267);
and U14027 (N_14027,N_9337,N_8112);
nor U14028 (N_14028,N_6847,N_5649);
or U14029 (N_14029,N_6058,N_7722);
xor U14030 (N_14030,N_5115,N_5125);
nor U14031 (N_14031,N_9911,N_9717);
nor U14032 (N_14032,N_7180,N_9085);
or U14033 (N_14033,N_7963,N_5782);
nand U14034 (N_14034,N_6764,N_5276);
and U14035 (N_14035,N_7681,N_8557);
or U14036 (N_14036,N_9754,N_8791);
xnor U14037 (N_14037,N_7776,N_5382);
or U14038 (N_14038,N_6663,N_6571);
xor U14039 (N_14039,N_8710,N_5342);
nor U14040 (N_14040,N_7892,N_7775);
and U14041 (N_14041,N_9122,N_7903);
nand U14042 (N_14042,N_8575,N_8278);
or U14043 (N_14043,N_5808,N_7333);
or U14044 (N_14044,N_6217,N_5324);
xor U14045 (N_14045,N_7391,N_8893);
and U14046 (N_14046,N_5056,N_8061);
nor U14047 (N_14047,N_6650,N_9413);
or U14048 (N_14048,N_8316,N_8062);
or U14049 (N_14049,N_9545,N_5837);
and U14050 (N_14050,N_5087,N_6680);
xor U14051 (N_14051,N_9649,N_8705);
nor U14052 (N_14052,N_9604,N_9011);
or U14053 (N_14053,N_7894,N_5940);
nor U14054 (N_14054,N_9629,N_5656);
xnor U14055 (N_14055,N_8223,N_5989);
nand U14056 (N_14056,N_9600,N_7516);
nand U14057 (N_14057,N_7507,N_6330);
nand U14058 (N_14058,N_7256,N_8105);
or U14059 (N_14059,N_5206,N_6082);
and U14060 (N_14060,N_7870,N_9405);
nand U14061 (N_14061,N_5686,N_5720);
nor U14062 (N_14062,N_9883,N_5184);
nand U14063 (N_14063,N_7553,N_8537);
and U14064 (N_14064,N_8113,N_5569);
nor U14065 (N_14065,N_6261,N_9127);
xor U14066 (N_14066,N_8074,N_5781);
nor U14067 (N_14067,N_8185,N_7241);
and U14068 (N_14068,N_7720,N_9238);
or U14069 (N_14069,N_9500,N_6565);
and U14070 (N_14070,N_8331,N_5302);
nor U14071 (N_14071,N_8983,N_7798);
xor U14072 (N_14072,N_9666,N_8833);
xor U14073 (N_14073,N_9210,N_6403);
or U14074 (N_14074,N_5751,N_9276);
nor U14075 (N_14075,N_9991,N_9827);
xor U14076 (N_14076,N_9085,N_5763);
and U14077 (N_14077,N_8980,N_5258);
xor U14078 (N_14078,N_8689,N_5589);
nand U14079 (N_14079,N_7548,N_7067);
nand U14080 (N_14080,N_8308,N_5217);
nand U14081 (N_14081,N_8292,N_7632);
nor U14082 (N_14082,N_7019,N_5592);
nor U14083 (N_14083,N_5054,N_5222);
or U14084 (N_14084,N_6104,N_6394);
xnor U14085 (N_14085,N_6170,N_7461);
or U14086 (N_14086,N_9298,N_5576);
or U14087 (N_14087,N_9927,N_9454);
xnor U14088 (N_14088,N_6376,N_5319);
nand U14089 (N_14089,N_8550,N_9385);
nor U14090 (N_14090,N_7569,N_9608);
nand U14091 (N_14091,N_8113,N_6351);
or U14092 (N_14092,N_6074,N_9981);
xor U14093 (N_14093,N_9941,N_6314);
nand U14094 (N_14094,N_8477,N_8354);
and U14095 (N_14095,N_7983,N_6563);
nor U14096 (N_14096,N_6722,N_9292);
or U14097 (N_14097,N_7144,N_9238);
nor U14098 (N_14098,N_7704,N_9200);
and U14099 (N_14099,N_7539,N_8412);
nor U14100 (N_14100,N_8164,N_8893);
or U14101 (N_14101,N_8872,N_5944);
xor U14102 (N_14102,N_8235,N_7992);
nand U14103 (N_14103,N_5676,N_9895);
nand U14104 (N_14104,N_6327,N_9406);
nand U14105 (N_14105,N_7899,N_6156);
nand U14106 (N_14106,N_5512,N_5632);
nand U14107 (N_14107,N_8783,N_7274);
nand U14108 (N_14108,N_9128,N_9431);
nand U14109 (N_14109,N_9218,N_9773);
and U14110 (N_14110,N_5197,N_9526);
nor U14111 (N_14111,N_8025,N_9190);
or U14112 (N_14112,N_7935,N_8147);
or U14113 (N_14113,N_7892,N_5183);
nor U14114 (N_14114,N_8498,N_6222);
and U14115 (N_14115,N_8658,N_8966);
or U14116 (N_14116,N_6492,N_9137);
nor U14117 (N_14117,N_5722,N_9015);
nor U14118 (N_14118,N_8799,N_9887);
and U14119 (N_14119,N_8062,N_5093);
nand U14120 (N_14120,N_5063,N_7328);
nand U14121 (N_14121,N_8495,N_7387);
or U14122 (N_14122,N_5751,N_7327);
nor U14123 (N_14123,N_9352,N_6195);
nand U14124 (N_14124,N_7201,N_8377);
and U14125 (N_14125,N_7093,N_5756);
xor U14126 (N_14126,N_7504,N_8148);
and U14127 (N_14127,N_9473,N_8571);
nor U14128 (N_14128,N_8963,N_9807);
nand U14129 (N_14129,N_7136,N_8867);
nor U14130 (N_14130,N_8897,N_5336);
or U14131 (N_14131,N_7388,N_5462);
or U14132 (N_14132,N_8861,N_5031);
and U14133 (N_14133,N_6469,N_7900);
nand U14134 (N_14134,N_6887,N_6311);
nand U14135 (N_14135,N_6274,N_6920);
and U14136 (N_14136,N_8076,N_5281);
xnor U14137 (N_14137,N_8540,N_9484);
or U14138 (N_14138,N_9881,N_6861);
or U14139 (N_14139,N_8487,N_6625);
and U14140 (N_14140,N_7560,N_5238);
xnor U14141 (N_14141,N_9559,N_6233);
and U14142 (N_14142,N_9507,N_7792);
or U14143 (N_14143,N_7525,N_7079);
nand U14144 (N_14144,N_9811,N_7044);
nand U14145 (N_14145,N_6275,N_9331);
nor U14146 (N_14146,N_8621,N_7621);
or U14147 (N_14147,N_5803,N_9851);
nand U14148 (N_14148,N_7266,N_8071);
nor U14149 (N_14149,N_5641,N_6459);
xor U14150 (N_14150,N_8927,N_6410);
or U14151 (N_14151,N_5572,N_5721);
nand U14152 (N_14152,N_9641,N_7137);
or U14153 (N_14153,N_9038,N_6516);
or U14154 (N_14154,N_8026,N_7035);
or U14155 (N_14155,N_6908,N_8178);
xnor U14156 (N_14156,N_7187,N_6126);
and U14157 (N_14157,N_5652,N_7728);
nand U14158 (N_14158,N_9195,N_5041);
and U14159 (N_14159,N_9968,N_8277);
or U14160 (N_14160,N_7806,N_9575);
nand U14161 (N_14161,N_6989,N_8940);
and U14162 (N_14162,N_5151,N_7879);
nor U14163 (N_14163,N_9537,N_7614);
nand U14164 (N_14164,N_5869,N_8591);
xnor U14165 (N_14165,N_6639,N_8211);
xor U14166 (N_14166,N_7752,N_6353);
xnor U14167 (N_14167,N_8273,N_6339);
xor U14168 (N_14168,N_9156,N_7075);
xor U14169 (N_14169,N_5473,N_7972);
nor U14170 (N_14170,N_5063,N_6370);
or U14171 (N_14171,N_9260,N_8379);
xnor U14172 (N_14172,N_5348,N_8314);
and U14173 (N_14173,N_5125,N_7716);
nand U14174 (N_14174,N_5127,N_6048);
xor U14175 (N_14175,N_9770,N_6195);
nor U14176 (N_14176,N_5377,N_5937);
and U14177 (N_14177,N_8733,N_9430);
nor U14178 (N_14178,N_6026,N_8896);
or U14179 (N_14179,N_6448,N_6675);
xor U14180 (N_14180,N_7297,N_7891);
xor U14181 (N_14181,N_6979,N_5318);
or U14182 (N_14182,N_7827,N_6684);
xor U14183 (N_14183,N_7580,N_8105);
and U14184 (N_14184,N_8423,N_8835);
nor U14185 (N_14185,N_6560,N_9576);
nand U14186 (N_14186,N_9608,N_9657);
or U14187 (N_14187,N_6416,N_9101);
and U14188 (N_14188,N_8318,N_5704);
xor U14189 (N_14189,N_5728,N_9784);
and U14190 (N_14190,N_6553,N_5102);
nand U14191 (N_14191,N_5212,N_7501);
or U14192 (N_14192,N_6671,N_5663);
xor U14193 (N_14193,N_8139,N_6740);
nand U14194 (N_14194,N_8770,N_5265);
nand U14195 (N_14195,N_9593,N_6593);
nand U14196 (N_14196,N_9476,N_5823);
nand U14197 (N_14197,N_8494,N_9817);
and U14198 (N_14198,N_5075,N_6254);
nor U14199 (N_14199,N_6747,N_8153);
nand U14200 (N_14200,N_7849,N_7688);
or U14201 (N_14201,N_6689,N_9593);
or U14202 (N_14202,N_6132,N_5506);
and U14203 (N_14203,N_6602,N_9131);
and U14204 (N_14204,N_9067,N_8608);
xnor U14205 (N_14205,N_5715,N_7627);
or U14206 (N_14206,N_7710,N_5599);
nand U14207 (N_14207,N_9471,N_9084);
nor U14208 (N_14208,N_7906,N_9712);
nand U14209 (N_14209,N_9011,N_7115);
nor U14210 (N_14210,N_7495,N_6363);
nor U14211 (N_14211,N_8241,N_6064);
and U14212 (N_14212,N_9365,N_9582);
nor U14213 (N_14213,N_6850,N_9267);
and U14214 (N_14214,N_7832,N_9063);
or U14215 (N_14215,N_9784,N_8666);
or U14216 (N_14216,N_6358,N_8378);
or U14217 (N_14217,N_9768,N_9484);
nand U14218 (N_14218,N_5783,N_5019);
and U14219 (N_14219,N_8024,N_7689);
or U14220 (N_14220,N_7454,N_7143);
or U14221 (N_14221,N_7198,N_9833);
or U14222 (N_14222,N_8362,N_6722);
nand U14223 (N_14223,N_7742,N_6184);
nand U14224 (N_14224,N_7547,N_9756);
nand U14225 (N_14225,N_5247,N_7026);
xnor U14226 (N_14226,N_9839,N_7882);
and U14227 (N_14227,N_7844,N_9695);
nand U14228 (N_14228,N_9509,N_9699);
or U14229 (N_14229,N_8993,N_8290);
and U14230 (N_14230,N_5538,N_9330);
xnor U14231 (N_14231,N_5203,N_7447);
xor U14232 (N_14232,N_9026,N_9424);
or U14233 (N_14233,N_7355,N_7192);
nand U14234 (N_14234,N_6071,N_6710);
xor U14235 (N_14235,N_9109,N_8996);
nand U14236 (N_14236,N_5901,N_5574);
xor U14237 (N_14237,N_9941,N_9432);
and U14238 (N_14238,N_6158,N_8278);
nor U14239 (N_14239,N_9296,N_6777);
xnor U14240 (N_14240,N_9666,N_7530);
nand U14241 (N_14241,N_8627,N_7272);
and U14242 (N_14242,N_6694,N_6218);
nand U14243 (N_14243,N_8389,N_9135);
nand U14244 (N_14244,N_9265,N_7617);
xor U14245 (N_14245,N_7739,N_8456);
and U14246 (N_14246,N_8039,N_5102);
or U14247 (N_14247,N_8793,N_8788);
and U14248 (N_14248,N_5531,N_8708);
nor U14249 (N_14249,N_8778,N_9417);
nand U14250 (N_14250,N_8632,N_9527);
nand U14251 (N_14251,N_5704,N_6437);
nor U14252 (N_14252,N_8591,N_5733);
and U14253 (N_14253,N_8007,N_7749);
nand U14254 (N_14254,N_9777,N_9342);
or U14255 (N_14255,N_9989,N_6262);
nor U14256 (N_14256,N_5769,N_7091);
xnor U14257 (N_14257,N_6173,N_8159);
nand U14258 (N_14258,N_7543,N_8132);
nand U14259 (N_14259,N_6522,N_6078);
and U14260 (N_14260,N_7770,N_9673);
and U14261 (N_14261,N_9385,N_5899);
and U14262 (N_14262,N_5943,N_5078);
or U14263 (N_14263,N_6928,N_7615);
nand U14264 (N_14264,N_6629,N_8700);
and U14265 (N_14265,N_9894,N_9183);
nand U14266 (N_14266,N_6732,N_9541);
xor U14267 (N_14267,N_8881,N_8971);
and U14268 (N_14268,N_5565,N_9500);
xor U14269 (N_14269,N_5939,N_8320);
xor U14270 (N_14270,N_8048,N_7688);
nor U14271 (N_14271,N_9118,N_5731);
and U14272 (N_14272,N_5364,N_8109);
or U14273 (N_14273,N_8082,N_9943);
or U14274 (N_14274,N_7573,N_5854);
xnor U14275 (N_14275,N_7353,N_8370);
nand U14276 (N_14276,N_9936,N_7112);
nor U14277 (N_14277,N_9873,N_9375);
nand U14278 (N_14278,N_7287,N_6036);
nor U14279 (N_14279,N_6846,N_6136);
xnor U14280 (N_14280,N_7802,N_8786);
and U14281 (N_14281,N_5200,N_9193);
and U14282 (N_14282,N_8642,N_6197);
or U14283 (N_14283,N_8611,N_8095);
xnor U14284 (N_14284,N_5749,N_8960);
and U14285 (N_14285,N_9402,N_6374);
or U14286 (N_14286,N_8289,N_9542);
or U14287 (N_14287,N_9141,N_6458);
xor U14288 (N_14288,N_9015,N_8864);
and U14289 (N_14289,N_9284,N_6327);
xor U14290 (N_14290,N_5577,N_9876);
and U14291 (N_14291,N_9080,N_8727);
and U14292 (N_14292,N_8023,N_8597);
or U14293 (N_14293,N_8116,N_6474);
nand U14294 (N_14294,N_8274,N_5741);
nor U14295 (N_14295,N_8383,N_7704);
and U14296 (N_14296,N_5397,N_9711);
and U14297 (N_14297,N_6004,N_8973);
or U14298 (N_14298,N_9701,N_6263);
nor U14299 (N_14299,N_6429,N_6112);
or U14300 (N_14300,N_7509,N_7390);
or U14301 (N_14301,N_6149,N_6371);
and U14302 (N_14302,N_9298,N_5908);
xor U14303 (N_14303,N_6051,N_7515);
nor U14304 (N_14304,N_8148,N_5610);
xnor U14305 (N_14305,N_8822,N_9244);
xnor U14306 (N_14306,N_8196,N_8766);
nor U14307 (N_14307,N_5856,N_9892);
and U14308 (N_14308,N_8604,N_9121);
and U14309 (N_14309,N_8914,N_7354);
nand U14310 (N_14310,N_9599,N_9443);
and U14311 (N_14311,N_5000,N_7812);
nand U14312 (N_14312,N_6128,N_6194);
and U14313 (N_14313,N_8276,N_8661);
and U14314 (N_14314,N_6175,N_5667);
nor U14315 (N_14315,N_5047,N_6637);
or U14316 (N_14316,N_5468,N_5077);
xnor U14317 (N_14317,N_7674,N_7682);
nor U14318 (N_14318,N_7966,N_6538);
nor U14319 (N_14319,N_6183,N_9897);
nand U14320 (N_14320,N_8211,N_8477);
xnor U14321 (N_14321,N_8681,N_6935);
and U14322 (N_14322,N_6442,N_7000);
and U14323 (N_14323,N_5954,N_6629);
and U14324 (N_14324,N_8794,N_7492);
and U14325 (N_14325,N_9669,N_6435);
xor U14326 (N_14326,N_9077,N_6929);
or U14327 (N_14327,N_5898,N_7033);
or U14328 (N_14328,N_8299,N_9527);
or U14329 (N_14329,N_8402,N_5982);
nor U14330 (N_14330,N_8557,N_5752);
or U14331 (N_14331,N_9675,N_8924);
or U14332 (N_14332,N_7610,N_7428);
nand U14333 (N_14333,N_9184,N_5044);
and U14334 (N_14334,N_6477,N_6337);
or U14335 (N_14335,N_9231,N_9940);
and U14336 (N_14336,N_7072,N_5329);
nand U14337 (N_14337,N_7668,N_8756);
nand U14338 (N_14338,N_7038,N_7724);
xor U14339 (N_14339,N_6029,N_9684);
nand U14340 (N_14340,N_7019,N_8281);
nand U14341 (N_14341,N_8453,N_8009);
nor U14342 (N_14342,N_6759,N_6792);
or U14343 (N_14343,N_7577,N_8982);
nand U14344 (N_14344,N_5787,N_6318);
xor U14345 (N_14345,N_6276,N_7397);
or U14346 (N_14346,N_5341,N_9459);
and U14347 (N_14347,N_9240,N_5625);
nor U14348 (N_14348,N_6579,N_8016);
nand U14349 (N_14349,N_5709,N_9863);
xnor U14350 (N_14350,N_8151,N_9187);
nand U14351 (N_14351,N_9200,N_6112);
or U14352 (N_14352,N_6553,N_5038);
nand U14353 (N_14353,N_7446,N_7118);
nand U14354 (N_14354,N_8786,N_9652);
nand U14355 (N_14355,N_8525,N_8132);
xor U14356 (N_14356,N_8134,N_7405);
and U14357 (N_14357,N_7162,N_6395);
nor U14358 (N_14358,N_6279,N_7696);
nand U14359 (N_14359,N_5184,N_8628);
and U14360 (N_14360,N_7167,N_8449);
and U14361 (N_14361,N_5674,N_9549);
xor U14362 (N_14362,N_9405,N_7700);
xnor U14363 (N_14363,N_8934,N_7080);
nand U14364 (N_14364,N_9568,N_5222);
xnor U14365 (N_14365,N_9848,N_6845);
or U14366 (N_14366,N_7329,N_5896);
nand U14367 (N_14367,N_5805,N_7037);
nor U14368 (N_14368,N_8392,N_7512);
and U14369 (N_14369,N_7936,N_6044);
nand U14370 (N_14370,N_8779,N_6327);
nand U14371 (N_14371,N_9830,N_7779);
xor U14372 (N_14372,N_6343,N_5795);
or U14373 (N_14373,N_8112,N_5205);
nor U14374 (N_14374,N_7277,N_5742);
xnor U14375 (N_14375,N_8092,N_8240);
xor U14376 (N_14376,N_6038,N_6818);
nand U14377 (N_14377,N_7522,N_5718);
and U14378 (N_14378,N_7267,N_6866);
and U14379 (N_14379,N_9663,N_9265);
nand U14380 (N_14380,N_6688,N_6518);
xor U14381 (N_14381,N_9145,N_6337);
or U14382 (N_14382,N_7114,N_8261);
or U14383 (N_14383,N_9320,N_9271);
and U14384 (N_14384,N_8864,N_5208);
nand U14385 (N_14385,N_6947,N_8574);
and U14386 (N_14386,N_7154,N_5258);
and U14387 (N_14387,N_8345,N_5621);
and U14388 (N_14388,N_7597,N_5828);
nor U14389 (N_14389,N_8003,N_5911);
or U14390 (N_14390,N_7501,N_7986);
nor U14391 (N_14391,N_8507,N_8484);
nor U14392 (N_14392,N_7793,N_5707);
nor U14393 (N_14393,N_8082,N_5068);
and U14394 (N_14394,N_9936,N_8083);
nand U14395 (N_14395,N_7482,N_5038);
and U14396 (N_14396,N_6197,N_8378);
or U14397 (N_14397,N_9075,N_5340);
nand U14398 (N_14398,N_8508,N_6085);
xnor U14399 (N_14399,N_7874,N_8900);
xor U14400 (N_14400,N_6220,N_5362);
xnor U14401 (N_14401,N_5447,N_9150);
nor U14402 (N_14402,N_5674,N_8350);
nand U14403 (N_14403,N_8754,N_7074);
xor U14404 (N_14404,N_5998,N_5778);
xor U14405 (N_14405,N_6794,N_6597);
xnor U14406 (N_14406,N_6398,N_7497);
or U14407 (N_14407,N_7087,N_9439);
and U14408 (N_14408,N_8728,N_8438);
and U14409 (N_14409,N_7787,N_9074);
nand U14410 (N_14410,N_7896,N_9015);
xor U14411 (N_14411,N_7698,N_9867);
nor U14412 (N_14412,N_7713,N_8832);
or U14413 (N_14413,N_7604,N_5836);
and U14414 (N_14414,N_9093,N_7756);
nand U14415 (N_14415,N_5733,N_6245);
or U14416 (N_14416,N_6616,N_7357);
nor U14417 (N_14417,N_5960,N_8815);
or U14418 (N_14418,N_7990,N_8221);
nand U14419 (N_14419,N_8557,N_8260);
and U14420 (N_14420,N_7149,N_5665);
or U14421 (N_14421,N_9078,N_8740);
xnor U14422 (N_14422,N_5489,N_5901);
and U14423 (N_14423,N_9605,N_8622);
and U14424 (N_14424,N_6218,N_7910);
xnor U14425 (N_14425,N_6739,N_7043);
nand U14426 (N_14426,N_9797,N_5551);
nand U14427 (N_14427,N_5715,N_6081);
and U14428 (N_14428,N_5688,N_5811);
and U14429 (N_14429,N_9925,N_9110);
nand U14430 (N_14430,N_9173,N_7333);
xor U14431 (N_14431,N_9482,N_8470);
and U14432 (N_14432,N_9119,N_7332);
nor U14433 (N_14433,N_5304,N_6698);
and U14434 (N_14434,N_8391,N_7726);
nor U14435 (N_14435,N_6091,N_5259);
xor U14436 (N_14436,N_7117,N_5666);
nor U14437 (N_14437,N_7486,N_7492);
nor U14438 (N_14438,N_7577,N_9200);
nor U14439 (N_14439,N_8929,N_9684);
and U14440 (N_14440,N_7633,N_5216);
or U14441 (N_14441,N_5852,N_5764);
nand U14442 (N_14442,N_5531,N_5409);
or U14443 (N_14443,N_5679,N_6939);
xor U14444 (N_14444,N_9407,N_6756);
nand U14445 (N_14445,N_6858,N_9218);
and U14446 (N_14446,N_8178,N_9923);
nand U14447 (N_14447,N_9503,N_5048);
xor U14448 (N_14448,N_5884,N_8730);
and U14449 (N_14449,N_9770,N_8880);
xor U14450 (N_14450,N_9364,N_7600);
nand U14451 (N_14451,N_7378,N_6854);
nand U14452 (N_14452,N_5545,N_7959);
or U14453 (N_14453,N_8691,N_5443);
or U14454 (N_14454,N_5692,N_6951);
xor U14455 (N_14455,N_8827,N_7264);
nand U14456 (N_14456,N_8112,N_9646);
and U14457 (N_14457,N_9946,N_8165);
and U14458 (N_14458,N_7085,N_6085);
nand U14459 (N_14459,N_9112,N_7599);
nor U14460 (N_14460,N_9070,N_6781);
nand U14461 (N_14461,N_9914,N_8976);
xor U14462 (N_14462,N_9550,N_8222);
or U14463 (N_14463,N_8678,N_9845);
or U14464 (N_14464,N_5278,N_9991);
and U14465 (N_14465,N_6522,N_9406);
nor U14466 (N_14466,N_9392,N_5344);
nor U14467 (N_14467,N_9266,N_5998);
xor U14468 (N_14468,N_8307,N_9733);
nand U14469 (N_14469,N_7389,N_6787);
nand U14470 (N_14470,N_7650,N_7326);
nand U14471 (N_14471,N_6933,N_8598);
nand U14472 (N_14472,N_8999,N_5163);
xnor U14473 (N_14473,N_7446,N_8566);
and U14474 (N_14474,N_6362,N_5784);
xor U14475 (N_14475,N_7613,N_9685);
nand U14476 (N_14476,N_6508,N_9156);
nor U14477 (N_14477,N_7148,N_8131);
nor U14478 (N_14478,N_5722,N_6828);
nand U14479 (N_14479,N_7213,N_8537);
nor U14480 (N_14480,N_7660,N_9719);
nand U14481 (N_14481,N_9325,N_8646);
or U14482 (N_14482,N_6791,N_9944);
xor U14483 (N_14483,N_7682,N_9753);
or U14484 (N_14484,N_6107,N_7851);
and U14485 (N_14485,N_5837,N_7002);
nand U14486 (N_14486,N_9031,N_6351);
or U14487 (N_14487,N_6112,N_5958);
or U14488 (N_14488,N_9263,N_6836);
and U14489 (N_14489,N_5194,N_9423);
nor U14490 (N_14490,N_9247,N_6828);
and U14491 (N_14491,N_5415,N_5338);
or U14492 (N_14492,N_5717,N_5833);
nor U14493 (N_14493,N_5397,N_6154);
and U14494 (N_14494,N_9168,N_5110);
or U14495 (N_14495,N_9280,N_7479);
xor U14496 (N_14496,N_7607,N_7556);
nor U14497 (N_14497,N_5367,N_6547);
or U14498 (N_14498,N_5945,N_6130);
and U14499 (N_14499,N_5124,N_8188);
and U14500 (N_14500,N_7803,N_9394);
nand U14501 (N_14501,N_6751,N_7346);
nor U14502 (N_14502,N_8665,N_8815);
nor U14503 (N_14503,N_6116,N_8585);
or U14504 (N_14504,N_7069,N_7305);
xnor U14505 (N_14505,N_8811,N_6406);
and U14506 (N_14506,N_6320,N_5821);
xor U14507 (N_14507,N_9107,N_5254);
and U14508 (N_14508,N_8773,N_7448);
nand U14509 (N_14509,N_8874,N_8961);
nor U14510 (N_14510,N_8976,N_7622);
nor U14511 (N_14511,N_5910,N_5471);
xor U14512 (N_14512,N_9198,N_9839);
and U14513 (N_14513,N_5504,N_5821);
or U14514 (N_14514,N_5376,N_5865);
and U14515 (N_14515,N_7827,N_5346);
nand U14516 (N_14516,N_6359,N_5265);
xnor U14517 (N_14517,N_5472,N_6970);
and U14518 (N_14518,N_5953,N_8536);
nor U14519 (N_14519,N_6183,N_6025);
xor U14520 (N_14520,N_9581,N_7202);
nand U14521 (N_14521,N_5586,N_5311);
nor U14522 (N_14522,N_9962,N_6325);
or U14523 (N_14523,N_5255,N_9631);
nand U14524 (N_14524,N_7125,N_8941);
xor U14525 (N_14525,N_9809,N_9122);
and U14526 (N_14526,N_9806,N_6452);
or U14527 (N_14527,N_7513,N_9356);
nand U14528 (N_14528,N_9369,N_6863);
nand U14529 (N_14529,N_8080,N_9489);
nor U14530 (N_14530,N_5840,N_6957);
and U14531 (N_14531,N_5495,N_9271);
nor U14532 (N_14532,N_9731,N_7926);
nand U14533 (N_14533,N_9703,N_6423);
or U14534 (N_14534,N_7058,N_6926);
and U14535 (N_14535,N_9446,N_9460);
nand U14536 (N_14536,N_6512,N_5810);
xor U14537 (N_14537,N_7432,N_7880);
xor U14538 (N_14538,N_8252,N_7241);
and U14539 (N_14539,N_8225,N_7601);
or U14540 (N_14540,N_8062,N_8192);
nor U14541 (N_14541,N_7692,N_8823);
nor U14542 (N_14542,N_7956,N_8611);
or U14543 (N_14543,N_8874,N_8569);
and U14544 (N_14544,N_5648,N_9804);
xor U14545 (N_14545,N_8380,N_5540);
nor U14546 (N_14546,N_9784,N_6783);
and U14547 (N_14547,N_7565,N_6412);
nand U14548 (N_14548,N_8099,N_8950);
nor U14549 (N_14549,N_9511,N_8779);
xnor U14550 (N_14550,N_7950,N_6357);
or U14551 (N_14551,N_5411,N_9633);
or U14552 (N_14552,N_7231,N_6936);
nor U14553 (N_14553,N_9154,N_6000);
nor U14554 (N_14554,N_9105,N_8748);
nor U14555 (N_14555,N_8041,N_6860);
and U14556 (N_14556,N_8239,N_6190);
and U14557 (N_14557,N_8309,N_5456);
and U14558 (N_14558,N_7892,N_8217);
nand U14559 (N_14559,N_9859,N_6067);
xnor U14560 (N_14560,N_6661,N_6683);
or U14561 (N_14561,N_7048,N_5158);
xnor U14562 (N_14562,N_7723,N_6646);
or U14563 (N_14563,N_9968,N_5223);
nor U14564 (N_14564,N_7582,N_9238);
nor U14565 (N_14565,N_7013,N_5834);
xor U14566 (N_14566,N_8658,N_6091);
or U14567 (N_14567,N_5576,N_6185);
xor U14568 (N_14568,N_9307,N_5432);
nand U14569 (N_14569,N_6665,N_7216);
nand U14570 (N_14570,N_9716,N_5818);
nand U14571 (N_14571,N_8053,N_6369);
nand U14572 (N_14572,N_9623,N_8898);
xnor U14573 (N_14573,N_5733,N_9681);
and U14574 (N_14574,N_6907,N_5527);
and U14575 (N_14575,N_9254,N_5154);
xor U14576 (N_14576,N_8730,N_5033);
or U14577 (N_14577,N_7634,N_5836);
xor U14578 (N_14578,N_5005,N_7026);
or U14579 (N_14579,N_5581,N_8189);
nor U14580 (N_14580,N_8388,N_9992);
nor U14581 (N_14581,N_9426,N_8343);
and U14582 (N_14582,N_8059,N_6204);
and U14583 (N_14583,N_7466,N_7017);
and U14584 (N_14584,N_9503,N_8879);
or U14585 (N_14585,N_9600,N_8832);
nand U14586 (N_14586,N_9610,N_6419);
nor U14587 (N_14587,N_6031,N_7974);
nor U14588 (N_14588,N_8481,N_6741);
and U14589 (N_14589,N_8450,N_7039);
nand U14590 (N_14590,N_7039,N_6764);
or U14591 (N_14591,N_6732,N_7835);
or U14592 (N_14592,N_6502,N_9803);
and U14593 (N_14593,N_9562,N_7011);
or U14594 (N_14594,N_5813,N_9820);
or U14595 (N_14595,N_6843,N_9610);
or U14596 (N_14596,N_8291,N_9697);
xnor U14597 (N_14597,N_6845,N_9219);
nand U14598 (N_14598,N_5730,N_6091);
nand U14599 (N_14599,N_7425,N_6435);
and U14600 (N_14600,N_9060,N_8452);
xnor U14601 (N_14601,N_6043,N_5156);
nand U14602 (N_14602,N_7470,N_7737);
nor U14603 (N_14603,N_8800,N_6277);
and U14604 (N_14604,N_9063,N_5133);
xnor U14605 (N_14605,N_7093,N_9116);
nor U14606 (N_14606,N_8098,N_8997);
and U14607 (N_14607,N_6930,N_6380);
nor U14608 (N_14608,N_6726,N_7748);
and U14609 (N_14609,N_6830,N_6697);
nand U14610 (N_14610,N_9412,N_5850);
nor U14611 (N_14611,N_8897,N_7241);
or U14612 (N_14612,N_5950,N_7499);
or U14613 (N_14613,N_7196,N_9881);
nor U14614 (N_14614,N_9193,N_6484);
xnor U14615 (N_14615,N_9074,N_7672);
nor U14616 (N_14616,N_5479,N_5171);
nand U14617 (N_14617,N_5871,N_6034);
nand U14618 (N_14618,N_7087,N_8914);
and U14619 (N_14619,N_5250,N_6291);
or U14620 (N_14620,N_6787,N_7700);
and U14621 (N_14621,N_5965,N_5349);
and U14622 (N_14622,N_8657,N_8378);
and U14623 (N_14623,N_7724,N_6870);
nor U14624 (N_14624,N_8306,N_9634);
or U14625 (N_14625,N_8310,N_8460);
nand U14626 (N_14626,N_7531,N_7276);
or U14627 (N_14627,N_9001,N_5550);
or U14628 (N_14628,N_7922,N_7371);
nor U14629 (N_14629,N_6677,N_7790);
and U14630 (N_14630,N_7506,N_6605);
nor U14631 (N_14631,N_8229,N_9537);
nand U14632 (N_14632,N_6556,N_5240);
and U14633 (N_14633,N_9059,N_6109);
nand U14634 (N_14634,N_7889,N_9140);
xor U14635 (N_14635,N_8447,N_9187);
nand U14636 (N_14636,N_9727,N_9081);
nor U14637 (N_14637,N_5877,N_8376);
and U14638 (N_14638,N_5108,N_5006);
xnor U14639 (N_14639,N_5374,N_8765);
and U14640 (N_14640,N_5460,N_5742);
nand U14641 (N_14641,N_5432,N_9496);
xnor U14642 (N_14642,N_8050,N_9344);
and U14643 (N_14643,N_6291,N_7346);
and U14644 (N_14644,N_5086,N_6123);
xor U14645 (N_14645,N_9179,N_5957);
xor U14646 (N_14646,N_5122,N_5510);
xor U14647 (N_14647,N_9165,N_6930);
xor U14648 (N_14648,N_7317,N_6008);
and U14649 (N_14649,N_6153,N_8134);
xnor U14650 (N_14650,N_6327,N_8504);
nand U14651 (N_14651,N_8232,N_9802);
and U14652 (N_14652,N_5758,N_8790);
nand U14653 (N_14653,N_7718,N_8214);
nand U14654 (N_14654,N_9090,N_8927);
nand U14655 (N_14655,N_7808,N_7812);
or U14656 (N_14656,N_5104,N_9734);
nor U14657 (N_14657,N_7001,N_9079);
nor U14658 (N_14658,N_7629,N_5797);
nor U14659 (N_14659,N_5422,N_7931);
nor U14660 (N_14660,N_6091,N_5197);
and U14661 (N_14661,N_8788,N_6500);
xor U14662 (N_14662,N_5589,N_5447);
nor U14663 (N_14663,N_6088,N_8537);
xnor U14664 (N_14664,N_5761,N_8057);
nand U14665 (N_14665,N_9963,N_5613);
nand U14666 (N_14666,N_9336,N_9695);
or U14667 (N_14667,N_7300,N_9790);
and U14668 (N_14668,N_8715,N_7826);
or U14669 (N_14669,N_7222,N_6058);
nor U14670 (N_14670,N_9141,N_9143);
xnor U14671 (N_14671,N_6140,N_9402);
xnor U14672 (N_14672,N_7692,N_9904);
nand U14673 (N_14673,N_9226,N_9242);
and U14674 (N_14674,N_6162,N_6996);
nand U14675 (N_14675,N_8837,N_5650);
and U14676 (N_14676,N_5688,N_9878);
and U14677 (N_14677,N_6051,N_6479);
nor U14678 (N_14678,N_7546,N_6668);
and U14679 (N_14679,N_7243,N_5231);
xnor U14680 (N_14680,N_6871,N_6290);
xor U14681 (N_14681,N_8953,N_9968);
nor U14682 (N_14682,N_9357,N_5951);
or U14683 (N_14683,N_7246,N_5742);
xnor U14684 (N_14684,N_5157,N_6278);
xnor U14685 (N_14685,N_5944,N_7564);
and U14686 (N_14686,N_6666,N_6064);
nor U14687 (N_14687,N_5299,N_9026);
nand U14688 (N_14688,N_6315,N_6117);
nor U14689 (N_14689,N_6401,N_6241);
or U14690 (N_14690,N_9188,N_6383);
and U14691 (N_14691,N_7516,N_5981);
xnor U14692 (N_14692,N_7037,N_9932);
xnor U14693 (N_14693,N_6917,N_6014);
nand U14694 (N_14694,N_5460,N_8827);
or U14695 (N_14695,N_9672,N_7211);
or U14696 (N_14696,N_8562,N_5400);
xor U14697 (N_14697,N_7351,N_8271);
or U14698 (N_14698,N_7797,N_5147);
and U14699 (N_14699,N_5860,N_7536);
or U14700 (N_14700,N_6324,N_5630);
xor U14701 (N_14701,N_9705,N_7876);
nand U14702 (N_14702,N_5689,N_7464);
nor U14703 (N_14703,N_8706,N_9884);
xor U14704 (N_14704,N_7979,N_6791);
and U14705 (N_14705,N_9394,N_5254);
xor U14706 (N_14706,N_8891,N_7204);
or U14707 (N_14707,N_8660,N_9015);
and U14708 (N_14708,N_9286,N_8971);
nor U14709 (N_14709,N_9011,N_9681);
nand U14710 (N_14710,N_6275,N_5002);
nand U14711 (N_14711,N_7798,N_7976);
or U14712 (N_14712,N_6695,N_6534);
xnor U14713 (N_14713,N_6922,N_6312);
nor U14714 (N_14714,N_8916,N_5598);
nor U14715 (N_14715,N_8405,N_6618);
and U14716 (N_14716,N_6255,N_6248);
nor U14717 (N_14717,N_6927,N_5983);
nand U14718 (N_14718,N_5394,N_5628);
xnor U14719 (N_14719,N_7875,N_9615);
xor U14720 (N_14720,N_9583,N_8561);
or U14721 (N_14721,N_7130,N_7783);
xor U14722 (N_14722,N_7801,N_9999);
nor U14723 (N_14723,N_6069,N_8365);
nand U14724 (N_14724,N_5852,N_9796);
nand U14725 (N_14725,N_8879,N_5369);
and U14726 (N_14726,N_7978,N_7748);
nand U14727 (N_14727,N_8870,N_8781);
nor U14728 (N_14728,N_9495,N_5294);
xnor U14729 (N_14729,N_8674,N_6455);
and U14730 (N_14730,N_9569,N_5851);
nand U14731 (N_14731,N_8254,N_9356);
nor U14732 (N_14732,N_6220,N_9931);
or U14733 (N_14733,N_5070,N_8463);
xor U14734 (N_14734,N_8317,N_7541);
or U14735 (N_14735,N_9566,N_9242);
and U14736 (N_14736,N_5450,N_5492);
and U14737 (N_14737,N_5451,N_7167);
and U14738 (N_14738,N_8359,N_9322);
and U14739 (N_14739,N_7346,N_7944);
nor U14740 (N_14740,N_9393,N_6297);
xor U14741 (N_14741,N_7071,N_6456);
and U14742 (N_14742,N_7841,N_7346);
nand U14743 (N_14743,N_8494,N_6205);
nand U14744 (N_14744,N_7096,N_6048);
nor U14745 (N_14745,N_5858,N_9742);
and U14746 (N_14746,N_7282,N_7039);
xor U14747 (N_14747,N_9383,N_6227);
and U14748 (N_14748,N_6947,N_9993);
nand U14749 (N_14749,N_9798,N_9729);
nor U14750 (N_14750,N_5030,N_5813);
or U14751 (N_14751,N_7007,N_7869);
or U14752 (N_14752,N_9353,N_6490);
nand U14753 (N_14753,N_8293,N_5254);
and U14754 (N_14754,N_8727,N_8372);
and U14755 (N_14755,N_5988,N_8352);
or U14756 (N_14756,N_6922,N_6767);
xor U14757 (N_14757,N_7754,N_8284);
nor U14758 (N_14758,N_7032,N_9424);
nor U14759 (N_14759,N_7556,N_7904);
nand U14760 (N_14760,N_9005,N_7196);
nor U14761 (N_14761,N_6993,N_7479);
xnor U14762 (N_14762,N_8680,N_7962);
or U14763 (N_14763,N_7078,N_6775);
or U14764 (N_14764,N_6767,N_5137);
xor U14765 (N_14765,N_9163,N_7920);
or U14766 (N_14766,N_8977,N_5516);
nor U14767 (N_14767,N_9540,N_7062);
nor U14768 (N_14768,N_6678,N_5030);
nor U14769 (N_14769,N_6008,N_8763);
and U14770 (N_14770,N_6121,N_7231);
nand U14771 (N_14771,N_7123,N_9926);
xor U14772 (N_14772,N_5683,N_8553);
nor U14773 (N_14773,N_9934,N_5768);
or U14774 (N_14774,N_6182,N_6730);
nand U14775 (N_14775,N_6806,N_8459);
xor U14776 (N_14776,N_5803,N_8856);
nor U14777 (N_14777,N_5256,N_7295);
nand U14778 (N_14778,N_6101,N_5938);
or U14779 (N_14779,N_8395,N_8778);
xor U14780 (N_14780,N_5006,N_5171);
xnor U14781 (N_14781,N_7937,N_9951);
nor U14782 (N_14782,N_5514,N_6303);
or U14783 (N_14783,N_5656,N_6299);
and U14784 (N_14784,N_7551,N_9232);
nand U14785 (N_14785,N_6132,N_8349);
and U14786 (N_14786,N_7107,N_7873);
xor U14787 (N_14787,N_7282,N_9071);
nand U14788 (N_14788,N_6352,N_8402);
nor U14789 (N_14789,N_9957,N_8605);
nand U14790 (N_14790,N_8151,N_6144);
or U14791 (N_14791,N_9149,N_7022);
xor U14792 (N_14792,N_7703,N_5158);
or U14793 (N_14793,N_6602,N_5492);
nor U14794 (N_14794,N_9981,N_9232);
and U14795 (N_14795,N_8841,N_6391);
and U14796 (N_14796,N_7260,N_5329);
or U14797 (N_14797,N_9205,N_8434);
or U14798 (N_14798,N_9984,N_8105);
nor U14799 (N_14799,N_8644,N_9267);
xor U14800 (N_14800,N_8808,N_6849);
or U14801 (N_14801,N_6781,N_9620);
nand U14802 (N_14802,N_6232,N_6578);
or U14803 (N_14803,N_6799,N_9512);
and U14804 (N_14804,N_5851,N_7608);
nand U14805 (N_14805,N_7349,N_6362);
or U14806 (N_14806,N_9336,N_7701);
nor U14807 (N_14807,N_9341,N_9673);
and U14808 (N_14808,N_9323,N_5716);
nand U14809 (N_14809,N_7776,N_8652);
and U14810 (N_14810,N_5096,N_8704);
xor U14811 (N_14811,N_8987,N_7801);
nand U14812 (N_14812,N_5419,N_8908);
or U14813 (N_14813,N_5469,N_7653);
nor U14814 (N_14814,N_9758,N_6169);
nand U14815 (N_14815,N_8459,N_8208);
xnor U14816 (N_14816,N_9822,N_9615);
or U14817 (N_14817,N_5622,N_7405);
nand U14818 (N_14818,N_6762,N_6259);
xor U14819 (N_14819,N_9079,N_9338);
nand U14820 (N_14820,N_8757,N_8286);
and U14821 (N_14821,N_9979,N_8312);
and U14822 (N_14822,N_9475,N_5242);
or U14823 (N_14823,N_9681,N_9065);
nand U14824 (N_14824,N_8153,N_7419);
nand U14825 (N_14825,N_5723,N_8973);
nor U14826 (N_14826,N_6943,N_6775);
xor U14827 (N_14827,N_6404,N_9370);
nor U14828 (N_14828,N_8714,N_5240);
xnor U14829 (N_14829,N_5524,N_8771);
nor U14830 (N_14830,N_5847,N_6696);
nor U14831 (N_14831,N_5942,N_5667);
or U14832 (N_14832,N_7726,N_5318);
or U14833 (N_14833,N_5725,N_7176);
or U14834 (N_14834,N_6894,N_9795);
and U14835 (N_14835,N_5573,N_9036);
or U14836 (N_14836,N_5177,N_9754);
or U14837 (N_14837,N_7874,N_7622);
or U14838 (N_14838,N_7994,N_7577);
nor U14839 (N_14839,N_6813,N_5332);
and U14840 (N_14840,N_8075,N_9289);
nor U14841 (N_14841,N_5071,N_8187);
nand U14842 (N_14842,N_8490,N_7508);
nor U14843 (N_14843,N_7442,N_6602);
and U14844 (N_14844,N_6185,N_8229);
xor U14845 (N_14845,N_6300,N_9064);
xnor U14846 (N_14846,N_8456,N_7559);
nand U14847 (N_14847,N_8922,N_5834);
nor U14848 (N_14848,N_9510,N_9695);
nor U14849 (N_14849,N_8706,N_5606);
xor U14850 (N_14850,N_7924,N_9073);
xnor U14851 (N_14851,N_8930,N_7407);
nand U14852 (N_14852,N_8750,N_6896);
xor U14853 (N_14853,N_9080,N_9740);
nand U14854 (N_14854,N_9004,N_7935);
xnor U14855 (N_14855,N_5145,N_6345);
nor U14856 (N_14856,N_7562,N_5461);
or U14857 (N_14857,N_6752,N_6782);
or U14858 (N_14858,N_9627,N_7908);
xnor U14859 (N_14859,N_9893,N_7051);
and U14860 (N_14860,N_6402,N_9954);
and U14861 (N_14861,N_8367,N_6165);
nand U14862 (N_14862,N_7838,N_5375);
or U14863 (N_14863,N_8883,N_5372);
xnor U14864 (N_14864,N_6232,N_7178);
nand U14865 (N_14865,N_8357,N_5024);
xor U14866 (N_14866,N_9875,N_7333);
nor U14867 (N_14867,N_9975,N_8864);
or U14868 (N_14868,N_5991,N_6048);
and U14869 (N_14869,N_5343,N_5923);
nor U14870 (N_14870,N_8668,N_8458);
and U14871 (N_14871,N_8316,N_8878);
nor U14872 (N_14872,N_5337,N_6802);
or U14873 (N_14873,N_5409,N_8565);
nand U14874 (N_14874,N_8023,N_9249);
or U14875 (N_14875,N_8491,N_8371);
xnor U14876 (N_14876,N_5947,N_5287);
nor U14877 (N_14877,N_9943,N_7723);
nor U14878 (N_14878,N_6002,N_9346);
nand U14879 (N_14879,N_8206,N_5356);
nand U14880 (N_14880,N_7297,N_9947);
nand U14881 (N_14881,N_7043,N_9193);
and U14882 (N_14882,N_5071,N_5020);
nand U14883 (N_14883,N_6117,N_7818);
or U14884 (N_14884,N_5048,N_9426);
or U14885 (N_14885,N_7349,N_7779);
or U14886 (N_14886,N_5911,N_5208);
and U14887 (N_14887,N_6591,N_6769);
nand U14888 (N_14888,N_9564,N_8613);
nand U14889 (N_14889,N_8944,N_9266);
nor U14890 (N_14890,N_6505,N_9149);
nor U14891 (N_14891,N_5916,N_8927);
or U14892 (N_14892,N_6353,N_8798);
xnor U14893 (N_14893,N_9701,N_6673);
and U14894 (N_14894,N_6917,N_9074);
or U14895 (N_14895,N_8129,N_5754);
xor U14896 (N_14896,N_8800,N_6841);
nor U14897 (N_14897,N_7177,N_7121);
and U14898 (N_14898,N_9122,N_7500);
nand U14899 (N_14899,N_8932,N_9526);
or U14900 (N_14900,N_5530,N_7741);
xnor U14901 (N_14901,N_9798,N_5034);
or U14902 (N_14902,N_9466,N_5957);
or U14903 (N_14903,N_5891,N_5746);
nand U14904 (N_14904,N_7468,N_9287);
xnor U14905 (N_14905,N_8035,N_8565);
or U14906 (N_14906,N_6807,N_9741);
and U14907 (N_14907,N_6863,N_7128);
xor U14908 (N_14908,N_5510,N_8882);
nor U14909 (N_14909,N_7318,N_7930);
nand U14910 (N_14910,N_6168,N_8310);
or U14911 (N_14911,N_9555,N_9375);
or U14912 (N_14912,N_6007,N_6930);
xor U14913 (N_14913,N_5786,N_6617);
nor U14914 (N_14914,N_9305,N_5289);
nor U14915 (N_14915,N_7476,N_6772);
or U14916 (N_14916,N_8856,N_8329);
or U14917 (N_14917,N_8075,N_7500);
and U14918 (N_14918,N_6708,N_5991);
or U14919 (N_14919,N_9628,N_9469);
and U14920 (N_14920,N_7682,N_7826);
and U14921 (N_14921,N_7986,N_8710);
and U14922 (N_14922,N_8026,N_6037);
or U14923 (N_14923,N_8499,N_5720);
or U14924 (N_14924,N_5809,N_5914);
and U14925 (N_14925,N_5179,N_5583);
nand U14926 (N_14926,N_6480,N_8220);
nor U14927 (N_14927,N_7352,N_8777);
xor U14928 (N_14928,N_8211,N_6668);
nand U14929 (N_14929,N_7186,N_9294);
and U14930 (N_14930,N_7361,N_5125);
xnor U14931 (N_14931,N_9243,N_5084);
or U14932 (N_14932,N_8374,N_6486);
nor U14933 (N_14933,N_8293,N_5555);
and U14934 (N_14934,N_5462,N_8538);
nand U14935 (N_14935,N_8816,N_6303);
or U14936 (N_14936,N_8139,N_6642);
xor U14937 (N_14937,N_7415,N_9742);
nand U14938 (N_14938,N_8806,N_9906);
and U14939 (N_14939,N_9971,N_5399);
nand U14940 (N_14940,N_9114,N_8300);
nor U14941 (N_14941,N_6916,N_5978);
and U14942 (N_14942,N_8182,N_8861);
nor U14943 (N_14943,N_5532,N_6000);
xor U14944 (N_14944,N_9553,N_9480);
nand U14945 (N_14945,N_9709,N_5497);
or U14946 (N_14946,N_9804,N_7402);
nand U14947 (N_14947,N_6415,N_8216);
xor U14948 (N_14948,N_7721,N_7183);
nand U14949 (N_14949,N_6875,N_8553);
or U14950 (N_14950,N_5228,N_6962);
xnor U14951 (N_14951,N_7700,N_9696);
or U14952 (N_14952,N_7689,N_9047);
nand U14953 (N_14953,N_8096,N_8223);
or U14954 (N_14954,N_9251,N_5306);
xnor U14955 (N_14955,N_6835,N_7863);
and U14956 (N_14956,N_8507,N_6133);
and U14957 (N_14957,N_6070,N_7324);
and U14958 (N_14958,N_8546,N_7838);
nor U14959 (N_14959,N_9931,N_6203);
xnor U14960 (N_14960,N_8476,N_7209);
nor U14961 (N_14961,N_8928,N_9690);
xnor U14962 (N_14962,N_5471,N_9686);
or U14963 (N_14963,N_9911,N_7150);
nand U14964 (N_14964,N_5211,N_9994);
xnor U14965 (N_14965,N_8624,N_9051);
nor U14966 (N_14966,N_9731,N_9822);
and U14967 (N_14967,N_5589,N_7582);
nor U14968 (N_14968,N_9268,N_6242);
nand U14969 (N_14969,N_7499,N_8125);
nor U14970 (N_14970,N_5570,N_6050);
nand U14971 (N_14971,N_6473,N_9605);
and U14972 (N_14972,N_6333,N_8335);
or U14973 (N_14973,N_8478,N_7956);
xnor U14974 (N_14974,N_5101,N_8783);
nand U14975 (N_14975,N_9284,N_6020);
nand U14976 (N_14976,N_9786,N_8567);
nor U14977 (N_14977,N_8919,N_9375);
or U14978 (N_14978,N_5207,N_7207);
xor U14979 (N_14979,N_8382,N_9718);
nand U14980 (N_14980,N_6155,N_7000);
or U14981 (N_14981,N_7070,N_8988);
and U14982 (N_14982,N_6721,N_9250);
nor U14983 (N_14983,N_6892,N_6682);
xor U14984 (N_14984,N_8514,N_6234);
or U14985 (N_14985,N_8142,N_8619);
xnor U14986 (N_14986,N_5861,N_6315);
nor U14987 (N_14987,N_6041,N_5172);
nand U14988 (N_14988,N_9752,N_9774);
and U14989 (N_14989,N_9519,N_9945);
nor U14990 (N_14990,N_7552,N_6400);
xnor U14991 (N_14991,N_9118,N_5053);
nor U14992 (N_14992,N_7008,N_6465);
or U14993 (N_14993,N_6852,N_5969);
or U14994 (N_14994,N_9260,N_7780);
or U14995 (N_14995,N_8901,N_5427);
nor U14996 (N_14996,N_5365,N_6558);
and U14997 (N_14997,N_6219,N_7446);
nor U14998 (N_14998,N_7015,N_5994);
and U14999 (N_14999,N_9021,N_5166);
nand UO_0 (O_0,N_10446,N_10658);
nor UO_1 (O_1,N_12725,N_11030);
xnor UO_2 (O_2,N_11366,N_14082);
xor UO_3 (O_3,N_10227,N_12770);
nor UO_4 (O_4,N_14637,N_13595);
and UO_5 (O_5,N_12196,N_11902);
xnor UO_6 (O_6,N_14615,N_13089);
nor UO_7 (O_7,N_12663,N_10553);
nor UO_8 (O_8,N_12550,N_13724);
xnor UO_9 (O_9,N_13479,N_12349);
nand UO_10 (O_10,N_14681,N_14465);
nor UO_11 (O_11,N_14386,N_14289);
and UO_12 (O_12,N_14212,N_14422);
xnor UO_13 (O_13,N_10153,N_13933);
nor UO_14 (O_14,N_13426,N_14370);
and UO_15 (O_15,N_14135,N_13293);
nor UO_16 (O_16,N_11795,N_11690);
or UO_17 (O_17,N_11160,N_14474);
nand UO_18 (O_18,N_12575,N_13133);
or UO_19 (O_19,N_10890,N_14771);
or UO_20 (O_20,N_10091,N_12113);
or UO_21 (O_21,N_14137,N_12074);
nand UO_22 (O_22,N_10893,N_11357);
nor UO_23 (O_23,N_14551,N_11779);
and UO_24 (O_24,N_14004,N_14395);
nand UO_25 (O_25,N_11486,N_14248);
nor UO_26 (O_26,N_13387,N_11585);
nor UO_27 (O_27,N_14832,N_10858);
or UO_28 (O_28,N_10667,N_14697);
and UO_29 (O_29,N_14538,N_10229);
and UO_30 (O_30,N_10250,N_14099);
nor UO_31 (O_31,N_13333,N_10792);
or UO_32 (O_32,N_12237,N_12367);
xnor UO_33 (O_33,N_12556,N_14294);
xnor UO_34 (O_34,N_13557,N_11525);
nor UO_35 (O_35,N_13896,N_11359);
xor UO_36 (O_36,N_14504,N_10030);
xor UO_37 (O_37,N_13371,N_11345);
or UO_38 (O_38,N_10962,N_13540);
nand UO_39 (O_39,N_11023,N_13820);
or UO_40 (O_40,N_14316,N_12120);
and UO_41 (O_41,N_12202,N_13539);
nor UO_42 (O_42,N_14659,N_12332);
nor UO_43 (O_43,N_13869,N_11700);
nor UO_44 (O_44,N_13704,N_13608);
xor UO_45 (O_45,N_12793,N_14264);
nor UO_46 (O_46,N_10843,N_14893);
xor UO_47 (O_47,N_11260,N_10264);
xnor UO_48 (O_48,N_10562,N_13817);
xor UO_49 (O_49,N_13187,N_13812);
nand UO_50 (O_50,N_12404,N_13458);
xnor UO_51 (O_51,N_11860,N_12073);
xnor UO_52 (O_52,N_10850,N_14320);
or UO_53 (O_53,N_10717,N_11267);
nand UO_54 (O_54,N_12672,N_12827);
nor UO_55 (O_55,N_14895,N_11894);
nand UO_56 (O_56,N_11340,N_10711);
and UO_57 (O_57,N_12620,N_10088);
xor UO_58 (O_58,N_13946,N_10066);
nor UO_59 (O_59,N_13879,N_12699);
and UO_60 (O_60,N_13065,N_14518);
nor UO_61 (O_61,N_10151,N_14980);
xnor UO_62 (O_62,N_11174,N_10311);
nand UO_63 (O_63,N_13408,N_14463);
nand UO_64 (O_64,N_11342,N_13254);
xor UO_65 (O_65,N_11370,N_12723);
or UO_66 (O_66,N_11577,N_12278);
or UO_67 (O_67,N_12234,N_14159);
xnor UO_68 (O_68,N_13911,N_12121);
nor UO_69 (O_69,N_11104,N_11053);
and UO_70 (O_70,N_10539,N_14971);
nor UO_71 (O_71,N_14113,N_12433);
xnor UO_72 (O_72,N_10086,N_11048);
or UO_73 (O_73,N_11664,N_12402);
and UO_74 (O_74,N_14985,N_13437);
or UO_75 (O_75,N_12931,N_10732);
nand UO_76 (O_76,N_13576,N_13047);
and UO_77 (O_77,N_11094,N_10862);
and UO_78 (O_78,N_14715,N_11960);
xor UO_79 (O_79,N_10127,N_14675);
nand UO_80 (O_80,N_10125,N_10508);
and UO_81 (O_81,N_13234,N_14851);
xor UO_82 (O_82,N_13694,N_10874);
and UO_83 (O_83,N_13320,N_10304);
nand UO_84 (O_84,N_12316,N_11505);
or UO_85 (O_85,N_11316,N_12595);
or UO_86 (O_86,N_11974,N_11773);
nor UO_87 (O_87,N_11456,N_10406);
nand UO_88 (O_88,N_12938,N_14933);
and UO_89 (O_89,N_13581,N_10072);
or UO_90 (O_90,N_10137,N_11841);
and UO_91 (O_91,N_11776,N_11204);
xnor UO_92 (O_92,N_12884,N_10089);
nor UO_93 (O_93,N_10494,N_14567);
nor UO_94 (O_94,N_13265,N_13375);
or UO_95 (O_95,N_13490,N_12045);
and UO_96 (O_96,N_10260,N_14757);
nor UO_97 (O_97,N_10922,N_10338);
and UO_98 (O_98,N_10727,N_13406);
or UO_99 (O_99,N_12730,N_14695);
and UO_100 (O_100,N_13367,N_10369);
and UO_101 (O_101,N_12929,N_12114);
xnor UO_102 (O_102,N_10592,N_12634);
nor UO_103 (O_103,N_12221,N_12908);
and UO_104 (O_104,N_14952,N_10313);
and UO_105 (O_105,N_10768,N_13283);
xnor UO_106 (O_106,N_14270,N_12953);
xnor UO_107 (O_107,N_13097,N_10710);
nor UO_108 (O_108,N_12134,N_11077);
nor UO_109 (O_109,N_13229,N_14723);
or UO_110 (O_110,N_12739,N_11772);
or UO_111 (O_111,N_11872,N_11728);
or UO_112 (O_112,N_14534,N_10972);
nor UO_113 (O_113,N_13120,N_14399);
nand UO_114 (O_114,N_13685,N_12016);
or UO_115 (O_115,N_13693,N_14296);
nor UO_116 (O_116,N_12246,N_11828);
nand UO_117 (O_117,N_12690,N_11972);
and UO_118 (O_118,N_13448,N_13980);
nor UO_119 (O_119,N_13009,N_13649);
nor UO_120 (O_120,N_14600,N_12598);
nand UO_121 (O_121,N_12071,N_14634);
xor UO_122 (O_122,N_12506,N_12893);
and UO_123 (O_123,N_14136,N_14936);
xor UO_124 (O_124,N_13908,N_14578);
nor UO_125 (O_125,N_11521,N_13118);
xor UO_126 (O_126,N_13909,N_12366);
and UO_127 (O_127,N_12470,N_14444);
or UO_128 (O_128,N_11892,N_13793);
nand UO_129 (O_129,N_12662,N_10584);
or UO_130 (O_130,N_14792,N_10077);
and UO_131 (O_131,N_10484,N_13432);
nor UO_132 (O_132,N_12263,N_10943);
and UO_133 (O_133,N_14498,N_14947);
or UO_134 (O_134,N_13477,N_14139);
nor UO_135 (O_135,N_13252,N_12233);
and UO_136 (O_136,N_12297,N_12803);
nor UO_137 (O_137,N_11001,N_12849);
or UO_138 (O_138,N_11870,N_10546);
and UO_139 (O_139,N_11344,N_14245);
nand UO_140 (O_140,N_14674,N_13476);
and UO_141 (O_141,N_12386,N_11150);
nand UO_142 (O_142,N_14523,N_14312);
nand UO_143 (O_143,N_14736,N_10016);
xnor UO_144 (O_144,N_13904,N_13722);
nand UO_145 (O_145,N_10184,N_13082);
xnor UO_146 (O_146,N_11587,N_12606);
and UO_147 (O_147,N_10457,N_12306);
and UO_148 (O_148,N_12464,N_14722);
and UO_149 (O_149,N_12650,N_13369);
xor UO_150 (O_150,N_14494,N_13236);
nand UO_151 (O_151,N_11032,N_11284);
nor UO_152 (O_152,N_14220,N_12920);
and UO_153 (O_153,N_14999,N_11561);
nor UO_154 (O_154,N_12731,N_11371);
xnor UO_155 (O_155,N_14215,N_10513);
or UO_156 (O_156,N_13355,N_11068);
and UO_157 (O_157,N_11115,N_10693);
xor UO_158 (O_158,N_12219,N_10419);
and UO_159 (O_159,N_12062,N_10202);
nor UO_160 (O_160,N_12379,N_14271);
nor UO_161 (O_161,N_11998,N_11413);
nand UO_162 (O_162,N_11481,N_11081);
nand UO_163 (O_163,N_12945,N_10404);
or UO_164 (O_164,N_12815,N_10699);
nand UO_165 (O_165,N_10742,N_11881);
and UO_166 (O_166,N_12872,N_13891);
xnor UO_167 (O_167,N_11938,N_13150);
xnor UO_168 (O_168,N_11312,N_14188);
and UO_169 (O_169,N_13652,N_12549);
nor UO_170 (O_170,N_13261,N_10243);
nand UO_171 (O_171,N_14358,N_14731);
or UO_172 (O_172,N_13447,N_13174);
and UO_173 (O_173,N_12272,N_10538);
nand UO_174 (O_174,N_11515,N_14105);
or UO_175 (O_175,N_13565,N_14405);
nor UO_176 (O_176,N_13679,N_14291);
or UO_177 (O_177,N_13160,N_11825);
or UO_178 (O_178,N_10317,N_10359);
nand UO_179 (O_179,N_12696,N_14401);
or UO_180 (O_180,N_14599,N_12521);
and UO_181 (O_181,N_12830,N_10928);
nor UO_182 (O_182,N_10054,N_13951);
xor UO_183 (O_183,N_12504,N_11125);
or UO_184 (O_184,N_11114,N_12442);
xor UO_185 (O_185,N_11571,N_10236);
xnor UO_186 (O_186,N_10506,N_14944);
nor UO_187 (O_187,N_12804,N_12104);
nor UO_188 (O_188,N_13346,N_13262);
or UO_189 (O_189,N_13591,N_14191);
nand UO_190 (O_190,N_11350,N_14404);
nand UO_191 (O_191,N_10452,N_12511);
xnor UO_192 (O_192,N_13847,N_11328);
xor UO_193 (O_193,N_10174,N_11074);
nor UO_194 (O_194,N_11511,N_13184);
and UO_195 (O_195,N_10914,N_14882);
or UO_196 (O_196,N_12105,N_12972);
and UO_197 (O_197,N_12683,N_14862);
nand UO_198 (O_198,N_11476,N_14311);
nand UO_199 (O_199,N_11020,N_12664);
and UO_200 (O_200,N_12307,N_13073);
or UO_201 (O_201,N_14535,N_14066);
xnor UO_202 (O_202,N_13973,N_12888);
xnor UO_203 (O_203,N_10150,N_13952);
xnor UO_204 (O_204,N_12907,N_11672);
or UO_205 (O_205,N_11581,N_12096);
nand UO_206 (O_206,N_12239,N_12116);
or UO_207 (O_207,N_13528,N_13496);
xnor UO_208 (O_208,N_12837,N_13859);
nand UO_209 (O_209,N_14906,N_14920);
or UO_210 (O_210,N_10001,N_11411);
nor UO_211 (O_211,N_12279,N_13788);
and UO_212 (O_212,N_13579,N_11092);
or UO_213 (O_213,N_13526,N_14200);
nand UO_214 (O_214,N_14040,N_12314);
and UO_215 (O_215,N_11252,N_10087);
xnor UO_216 (O_216,N_14735,N_13706);
xnor UO_217 (O_217,N_14114,N_11372);
xnor UO_218 (O_218,N_10058,N_12578);
nand UO_219 (O_219,N_11172,N_11210);
nor UO_220 (O_220,N_10136,N_12553);
xnor UO_221 (O_221,N_11869,N_13950);
nor UO_222 (O_222,N_14322,N_13422);
or UO_223 (O_223,N_12626,N_12162);
nand UO_224 (O_224,N_10067,N_13143);
nand UO_225 (O_225,N_13942,N_10428);
and UO_226 (O_226,N_10547,N_10363);
nor UO_227 (O_227,N_10283,N_11736);
or UO_228 (O_228,N_12003,N_13006);
nor UO_229 (O_229,N_13041,N_13308);
or UO_230 (O_230,N_14282,N_10022);
nor UO_231 (O_231,N_10079,N_11853);
nor UO_232 (O_232,N_11464,N_11954);
nand UO_233 (O_233,N_10838,N_13961);
nor UO_234 (O_234,N_13030,N_10822);
and UO_235 (O_235,N_11228,N_14533);
xor UO_236 (O_236,N_10188,N_14861);
and UO_237 (O_237,N_10115,N_13807);
and UO_238 (O_238,N_12780,N_12401);
xor UO_239 (O_239,N_11043,N_13131);
nor UO_240 (O_240,N_14062,N_14480);
nor UO_241 (O_241,N_13483,N_10552);
nor UO_242 (O_242,N_10294,N_13749);
nand UO_243 (O_243,N_11673,N_13675);
xnor UO_244 (O_244,N_12310,N_10764);
nor UO_245 (O_245,N_12897,N_13099);
or UO_246 (O_246,N_12787,N_10724);
nor UO_247 (O_247,N_10622,N_11945);
nand UO_248 (O_248,N_14868,N_12478);
nand UO_249 (O_249,N_11769,N_12268);
nand UO_250 (O_250,N_10346,N_13596);
xnor UO_251 (O_251,N_12517,N_11531);
nor UO_252 (O_252,N_10314,N_14396);
nor UO_253 (O_253,N_12743,N_12603);
xnor UO_254 (O_254,N_10831,N_10726);
and UO_255 (O_255,N_11949,N_12127);
xnor UO_256 (O_256,N_10602,N_13395);
or UO_257 (O_257,N_11322,N_12789);
nand UO_258 (O_258,N_11638,N_13624);
or UO_259 (O_259,N_13948,N_11784);
xor UO_260 (O_260,N_12147,N_11814);
nand UO_261 (O_261,N_10305,N_11739);
xnor UO_262 (O_262,N_14773,N_12427);
and UO_263 (O_263,N_11497,N_11360);
or UO_264 (O_264,N_10374,N_12472);
or UO_265 (O_265,N_13148,N_14644);
or UO_266 (O_266,N_10706,N_14830);
and UO_267 (O_267,N_13113,N_13373);
nand UO_268 (O_268,N_11480,N_11494);
xor UO_269 (O_269,N_14487,N_13286);
xor UO_270 (O_270,N_10777,N_11304);
xnor UO_271 (O_271,N_11072,N_14261);
or UO_272 (O_272,N_11128,N_10950);
xnor UO_273 (O_273,N_11006,N_10154);
nor UO_274 (O_274,N_14173,N_13077);
nand UO_275 (O_275,N_13709,N_13342);
nand UO_276 (O_276,N_11642,N_14522);
nor UO_277 (O_277,N_10354,N_13469);
or UO_278 (O_278,N_12093,N_10210);
nor UO_279 (O_279,N_14647,N_13833);
and UO_280 (O_280,N_13992,N_11804);
nor UO_281 (O_281,N_11144,N_10275);
xnor UO_282 (O_282,N_11744,N_12960);
nor UO_283 (O_283,N_14158,N_14263);
nor UO_284 (O_284,N_10752,N_12227);
xnor UO_285 (O_285,N_13549,N_12516);
or UO_286 (O_286,N_14046,N_11012);
xnor UO_287 (O_287,N_11556,N_12777);
xnor UO_288 (O_288,N_11932,N_10099);
or UO_289 (O_289,N_13713,N_10980);
nor UO_290 (O_290,N_14127,N_10619);
nor UO_291 (O_291,N_14038,N_10495);
nor UO_292 (O_292,N_13000,N_11626);
nand UO_293 (O_293,N_14489,N_11948);
nor UO_294 (O_294,N_11962,N_13697);
nand UO_295 (O_295,N_12503,N_14355);
xnor UO_296 (O_296,N_12975,N_12412);
xor UO_297 (O_297,N_13383,N_12076);
nand UO_298 (O_298,N_12144,N_10686);
or UO_299 (O_299,N_11584,N_10011);
or UO_300 (O_300,N_10548,N_11156);
and UO_301 (O_301,N_10119,N_11601);
and UO_302 (O_302,N_14726,N_11545);
nand UO_303 (O_303,N_14157,N_11173);
nor UO_304 (O_304,N_14297,N_12824);
or UO_305 (O_305,N_14469,N_13248);
or UO_306 (O_306,N_12290,N_12496);
nor UO_307 (O_307,N_13520,N_10786);
and UO_308 (O_308,N_11047,N_11215);
xor UO_309 (O_309,N_14619,N_13877);
nor UO_310 (O_310,N_12860,N_13681);
or UO_311 (O_311,N_11829,N_14970);
xor UO_312 (O_312,N_12601,N_14515);
xor UO_313 (O_313,N_11586,N_12526);
nor UO_314 (O_314,N_14507,N_12749);
nor UO_315 (O_315,N_10676,N_13985);
or UO_316 (O_316,N_12557,N_14957);
nand UO_317 (O_317,N_11688,N_11615);
and UO_318 (O_318,N_12211,N_14905);
or UO_319 (O_319,N_11073,N_12056);
xnor UO_320 (O_320,N_12059,N_10945);
or UO_321 (O_321,N_14513,N_11105);
xnor UO_322 (O_322,N_14692,N_12179);
or UO_323 (O_323,N_12172,N_13943);
nor UO_324 (O_324,N_13389,N_14475);
or UO_325 (O_325,N_13474,N_10490);
or UO_326 (O_326,N_11031,N_14373);
nand UO_327 (O_327,N_11551,N_11165);
xor UO_328 (O_328,N_12189,N_11827);
xnor UO_329 (O_329,N_12936,N_13304);
nor UO_330 (O_330,N_10431,N_13835);
xnor UO_331 (O_331,N_13436,N_12429);
nand UO_332 (O_332,N_10672,N_11487);
and UO_333 (O_333,N_12173,N_14890);
nand UO_334 (O_334,N_10370,N_11588);
nand UO_335 (O_335,N_13802,N_14211);
xor UO_336 (O_336,N_11605,N_10300);
or UO_337 (O_337,N_13075,N_10319);
nand UO_338 (O_338,N_13332,N_12748);
nand UO_339 (O_339,N_12535,N_10761);
and UO_340 (O_340,N_10587,N_14198);
or UO_341 (O_341,N_10694,N_12154);
xnor UO_342 (O_342,N_11103,N_11489);
or UO_343 (O_343,N_11921,N_11106);
nand UO_344 (O_344,N_10519,N_13122);
nor UO_345 (O_345,N_14877,N_14255);
or UO_346 (O_346,N_12727,N_14164);
nor UO_347 (O_347,N_11708,N_13718);
or UO_348 (O_348,N_14817,N_11933);
nand UO_349 (O_349,N_12922,N_13809);
xnor UO_350 (O_350,N_13715,N_12984);
and UO_351 (O_351,N_13580,N_14718);
xor UO_352 (O_352,N_11130,N_14846);
xnor UO_353 (O_353,N_12653,N_10954);
or UO_354 (O_354,N_11448,N_12346);
nand UO_355 (O_355,N_14162,N_12705);
and UO_356 (O_356,N_12244,N_14299);
and UO_357 (O_357,N_13881,N_12102);
nor UO_358 (O_358,N_11694,N_11861);
and UO_359 (O_359,N_13860,N_13760);
nand UO_360 (O_360,N_11663,N_14176);
and UO_361 (O_361,N_14341,N_12085);
nand UO_362 (O_362,N_10292,N_12004);
and UO_363 (O_363,N_11253,N_11484);
or UO_364 (O_364,N_14709,N_14875);
xnor UO_365 (O_365,N_12281,N_12865);
nand UO_366 (O_366,N_12819,N_10781);
and UO_367 (O_367,N_13035,N_11537);
or UO_368 (O_368,N_11209,N_14627);
and UO_369 (O_369,N_10181,N_11468);
or UO_370 (O_370,N_11276,N_11710);
nand UO_371 (O_371,N_13049,N_13587);
and UO_372 (O_372,N_12274,N_11071);
and UO_373 (O_373,N_13863,N_12821);
xor UO_374 (O_374,N_13791,N_10074);
xor UO_375 (O_375,N_13277,N_13511);
and UO_376 (O_376,N_11713,N_14006);
nor UO_377 (O_377,N_10211,N_11242);
and UO_378 (O_378,N_13553,N_14887);
nor UO_379 (O_379,N_14897,N_13177);
xor UO_380 (O_380,N_14705,N_10216);
nor UO_381 (O_381,N_12585,N_12106);
and UO_382 (O_382,N_10564,N_14935);
xnor UO_383 (O_383,N_10223,N_12322);
or UO_384 (O_384,N_12487,N_14307);
or UO_385 (O_385,N_14761,N_10606);
nor UO_386 (O_386,N_10938,N_12761);
xor UO_387 (O_387,N_14630,N_12117);
nand UO_388 (O_388,N_12293,N_12707);
nor UO_389 (O_389,N_13363,N_14976);
nor UO_390 (O_390,N_12946,N_13305);
nand UO_391 (O_391,N_14411,N_14663);
or UO_392 (O_392,N_14978,N_13653);
nand UO_393 (O_393,N_14916,N_14845);
nor UO_394 (O_394,N_13127,N_12025);
xnor UO_395 (O_395,N_12288,N_13472);
nor UO_396 (O_396,N_14867,N_12836);
xnor UO_397 (O_397,N_13682,N_11166);
and UO_398 (O_398,N_14981,N_12457);
nor UO_399 (O_399,N_14326,N_13205);
or UO_400 (O_400,N_14783,N_12871);
xnor UO_401 (O_401,N_11361,N_12800);
xnor UO_402 (O_402,N_12423,N_10352);
nor UO_403 (O_403,N_13114,N_10436);
nor UO_404 (O_404,N_12782,N_14259);
or UO_405 (O_405,N_12843,N_11803);
nand UO_406 (O_406,N_11430,N_11665);
nor UO_407 (O_407,N_12976,N_12925);
or UO_408 (O_408,N_11850,N_12635);
nor UO_409 (O_409,N_11797,N_10621);
and UO_410 (O_410,N_11259,N_11654);
or UO_411 (O_411,N_14556,N_11611);
and UO_412 (O_412,N_11216,N_13707);
xnor UO_413 (O_413,N_13403,N_13180);
xnor UO_414 (O_414,N_10341,N_10647);
xor UO_415 (O_415,N_12674,N_14811);
and UO_416 (O_416,N_11376,N_10021);
nand UO_417 (O_417,N_13850,N_12477);
nand UO_418 (O_418,N_14754,N_12490);
nand UO_419 (O_419,N_12580,N_13413);
nor UO_420 (O_420,N_14413,N_14917);
xnor UO_421 (O_421,N_10217,N_13084);
or UO_422 (O_422,N_11681,N_11212);
and UO_423 (O_423,N_13884,N_13680);
xor UO_424 (O_424,N_12532,N_12941);
xor UO_425 (O_425,N_14602,N_10029);
nand UO_426 (O_426,N_13640,N_13917);
or UO_427 (O_427,N_13894,N_10521);
xor UO_428 (O_428,N_10634,N_11022);
nor UO_429 (O_429,N_14904,N_12767);
nor UO_430 (O_430,N_13121,N_13785);
and UO_431 (O_431,N_11186,N_11321);
xor UO_432 (O_432,N_12629,N_14934);
nor UO_433 (O_433,N_11786,N_10328);
or UO_434 (O_434,N_14560,N_14071);
and UO_435 (O_435,N_13773,N_12407);
nor UO_436 (O_436,N_13033,N_11810);
nand UO_437 (O_437,N_11646,N_12398);
and UO_438 (O_438,N_14298,N_10579);
and UO_439 (O_439,N_10665,N_13040);
xnor UO_440 (O_440,N_12303,N_12098);
and UO_441 (O_441,N_11683,N_14112);
xor UO_442 (O_442,N_10959,N_11002);
xor UO_443 (O_443,N_11830,N_13545);
xor UO_444 (O_444,N_14827,N_11433);
nand UO_445 (O_445,N_12013,N_14946);
nand UO_446 (O_446,N_13714,N_10801);
nand UO_447 (O_447,N_12124,N_14948);
nand UO_448 (O_448,N_13287,N_12924);
nor UO_449 (O_449,N_14601,N_12165);
xnor UO_450 (O_450,N_11879,N_11995);
or UO_451 (O_451,N_11265,N_14310);
and UO_452 (O_452,N_12861,N_13630);
or UO_453 (O_453,N_10303,N_13269);
nand UO_454 (O_454,N_11781,N_12594);
or UO_455 (O_455,N_13603,N_14884);
and UO_456 (O_456,N_11078,N_11465);
or UO_457 (O_457,N_12950,N_13329);
xnor UO_458 (O_458,N_11715,N_10480);
nor UO_459 (O_459,N_11753,N_14193);
xor UO_460 (O_460,N_12082,N_12757);
or UO_461 (O_461,N_11557,N_13771);
nand UO_462 (O_462,N_13656,N_10266);
xnor UO_463 (O_463,N_13240,N_12260);
and UO_464 (O_464,N_10025,N_14012);
nand UO_465 (O_465,N_11888,N_10718);
xor UO_466 (O_466,N_10094,N_10358);
or UO_467 (O_467,N_11573,N_14431);
nor UO_468 (O_468,N_14016,N_12686);
nand UO_469 (O_469,N_12832,N_12942);
or UO_470 (O_470,N_11332,N_13931);
xor UO_471 (O_471,N_10389,N_10868);
or UO_472 (O_472,N_11013,N_12063);
or UO_473 (O_473,N_12951,N_11908);
nor UO_474 (O_474,N_12600,N_10156);
or UO_475 (O_475,N_12033,N_10493);
nand UO_476 (O_476,N_13532,N_11457);
nand UO_477 (O_477,N_10098,N_14573);
or UO_478 (O_478,N_11183,N_13235);
nand UO_479 (O_479,N_10318,N_10785);
nor UO_480 (O_480,N_11288,N_12437);
and UO_481 (O_481,N_14870,N_12740);
nand UO_482 (O_482,N_14719,N_11000);
nand UO_483 (O_483,N_12151,N_13870);
nand UO_484 (O_484,N_10900,N_11059);
or UO_485 (O_485,N_11171,N_13101);
and UO_486 (O_486,N_14838,N_13944);
or UO_487 (O_487,N_12964,N_14241);
and UO_488 (O_488,N_12041,N_14554);
nand UO_489 (O_489,N_14967,N_10738);
xnor UO_490 (O_490,N_10267,N_12276);
xor UO_491 (O_491,N_14854,N_10971);
nor UO_492 (O_492,N_12869,N_13270);
nor UO_493 (O_493,N_11201,N_10155);
nor UO_494 (O_494,N_14635,N_11896);
nand UO_495 (O_495,N_13050,N_12681);
or UO_496 (O_496,N_12957,N_11129);
xnor UO_497 (O_497,N_14177,N_11597);
nand UO_498 (O_498,N_10297,N_11903);
or UO_499 (O_499,N_13027,N_10367);
and UO_500 (O_500,N_12387,N_13340);
or UO_501 (O_501,N_14168,N_13473);
and UO_502 (O_502,N_11471,N_11268);
xnor UO_503 (O_503,N_14045,N_11750);
nand UO_504 (O_504,N_12471,N_10878);
xnor UO_505 (O_505,N_11198,N_11575);
and UO_506 (O_506,N_11363,N_13146);
nand UO_507 (O_507,N_14238,N_14900);
xnor UO_508 (O_508,N_14865,N_11578);
and UO_509 (O_509,N_13699,N_14313);
nand UO_510 (O_510,N_10039,N_10209);
nand UO_511 (O_511,N_14666,N_10251);
and UO_512 (O_512,N_11927,N_14684);
and UO_513 (O_513,N_14711,N_10867);
and UO_514 (O_514,N_14956,N_13787);
nand UO_515 (O_515,N_11095,N_14691);
xnor UO_516 (O_516,N_12042,N_12344);
xnor UO_517 (O_517,N_12614,N_11261);
and UO_518 (O_518,N_14769,N_11056);
xor UO_519 (O_519,N_10837,N_11667);
and UO_520 (O_520,N_12395,N_14385);
or UO_521 (O_521,N_10438,N_13263);
or UO_522 (O_522,N_11333,N_14383);
or UO_523 (O_523,N_13119,N_14746);
and UO_524 (O_524,N_13210,N_14894);
and UO_525 (O_525,N_12271,N_12625);
nand UO_526 (O_526,N_14154,N_10169);
or UO_527 (O_527,N_10765,N_13783);
or UO_528 (O_528,N_13209,N_13423);
and UO_529 (O_529,N_11595,N_14325);
nor UO_530 (O_530,N_11939,N_14053);
and UO_531 (O_531,N_14017,N_13727);
or UO_532 (O_532,N_10121,N_10636);
nand UO_533 (O_533,N_13074,N_10486);
or UO_534 (O_534,N_13736,N_13466);
nor UO_535 (O_535,N_10459,N_13154);
nor UO_536 (O_536,N_12138,N_13751);
nor UO_537 (O_537,N_12505,N_14620);
nand UO_538 (O_538,N_12447,N_10002);
or UO_539 (O_539,N_14035,N_12502);
xor UO_540 (O_540,N_14067,N_14725);
nand UO_541 (O_541,N_13491,N_11819);
nand UO_542 (O_542,N_10810,N_12142);
and UO_543 (O_543,N_11550,N_14087);
nand UO_544 (O_544,N_10688,N_14055);
nand UO_545 (O_545,N_13615,N_13965);
and UO_546 (O_546,N_10505,N_10161);
nand UO_547 (O_547,N_14517,N_10532);
or UO_548 (O_548,N_12171,N_12011);
or UO_549 (O_549,N_14015,N_10609);
nand UO_550 (O_550,N_11099,N_14279);
nor UO_551 (O_551,N_11984,N_12898);
or UO_552 (O_552,N_13347,N_14586);
xor UO_553 (O_553,N_13307,N_13763);
nand UO_554 (O_554,N_13388,N_11682);
nor UO_555 (O_555,N_13060,N_10791);
nor UO_556 (O_556,N_11527,N_13368);
xor UO_557 (O_557,N_10458,N_10399);
nand UO_558 (O_558,N_14964,N_13501);
xnor UO_559 (O_559,N_10830,N_11865);
nand UO_560 (O_560,N_14959,N_12356);
xnor UO_561 (O_561,N_13551,N_10649);
nor UO_562 (O_562,N_14057,N_14876);
and UO_563 (O_563,N_13419,N_14488);
xor UO_564 (O_564,N_12879,N_12399);
xor UO_565 (O_565,N_10152,N_10158);
nor UO_566 (O_566,N_14954,N_12390);
or UO_567 (O_567,N_13356,N_12773);
nor UO_568 (O_568,N_11065,N_13231);
nor UO_569 (O_569,N_11247,N_12345);
or UO_570 (O_570,N_11976,N_11732);
nand UO_571 (O_571,N_11176,N_12564);
nor UO_572 (O_572,N_13586,N_13173);
nor UO_573 (O_573,N_12333,N_11788);
nor UO_574 (O_574,N_14252,N_11632);
xnor UO_575 (O_575,N_13854,N_13158);
xor UO_576 (O_576,N_12997,N_14614);
or UO_577 (O_577,N_13641,N_10872);
nand UO_578 (O_578,N_14078,N_10886);
xor UO_579 (O_579,N_12903,N_14756);
xor UO_580 (O_580,N_13384,N_11177);
and UO_581 (O_581,N_11379,N_12916);
nand UO_582 (O_582,N_13559,N_10368);
and UO_583 (O_583,N_13135,N_11631);
or UO_584 (O_584,N_13087,N_11514);
and UO_585 (O_585,N_11289,N_14568);
nor UO_586 (O_586,N_14858,N_13534);
or UO_587 (O_587,N_13670,N_14645);
and UO_588 (O_588,N_10704,N_10325);
nand UO_589 (O_589,N_14623,N_14423);
nand UO_590 (O_590,N_11309,N_14553);
nor UO_591 (O_591,N_14069,N_11124);
nor UO_592 (O_592,N_14618,N_14343);
and UO_593 (O_593,N_11529,N_10833);
xnor UO_594 (O_594,N_13291,N_12669);
xnor UO_595 (O_595,N_10048,N_13054);
or UO_596 (O_596,N_10163,N_10422);
nor UO_597 (O_597,N_13636,N_11017);
nand UO_598 (O_598,N_12992,N_12754);
and UO_599 (O_599,N_10424,N_14408);
xor UO_600 (O_600,N_13439,N_13902);
xnor UO_601 (O_601,N_14204,N_12520);
nor UO_602 (O_602,N_11441,N_13574);
and UO_603 (O_603,N_10109,N_11025);
xor UO_604 (O_604,N_13414,N_12193);
or UO_605 (O_605,N_11199,N_12195);
nor UO_606 (O_606,N_11439,N_11337);
and UO_607 (O_607,N_12498,N_10750);
xnor UO_608 (O_608,N_10741,N_11604);
nor UO_609 (O_609,N_14145,N_13848);
or UO_610 (O_610,N_10398,N_10082);
xnor UO_611 (O_611,N_10985,N_10835);
nor UO_612 (O_612,N_13001,N_14994);
or UO_613 (O_613,N_10682,N_12092);
nor UO_614 (O_614,N_13512,N_13947);
and UO_615 (O_615,N_13993,N_10178);
xor UO_616 (O_616,N_13949,N_10270);
xor UO_617 (O_617,N_10306,N_11392);
nor UO_618 (O_618,N_14775,N_11470);
or UO_619 (O_619,N_14254,N_14506);
and UO_620 (O_620,N_14428,N_11579);
nor UO_621 (O_621,N_14548,N_13141);
and UO_622 (O_622,N_11987,N_12695);
xor UO_623 (O_623,N_12587,N_11671);
and UO_624 (O_624,N_14278,N_13200);
xnor UO_625 (O_625,N_13871,N_14185);
or UO_626 (O_626,N_14643,N_11269);
nor UO_627 (O_627,N_12602,N_12514);
xnor UO_628 (O_628,N_10320,N_12583);
or UO_629 (O_629,N_13798,N_12776);
xor UO_630 (O_630,N_10269,N_13918);
nor UO_631 (O_631,N_10336,N_11218);
nor UO_632 (O_632,N_14076,N_14036);
nor UO_633 (O_633,N_10915,N_13522);
or UO_634 (O_634,N_13328,N_10451);
nand UO_635 (O_635,N_14700,N_12656);
or UO_636 (O_636,N_11524,N_14909);
nand UO_637 (O_637,N_10111,N_11859);
nor UO_638 (O_638,N_14471,N_11169);
or UO_639 (O_639,N_11330,N_14042);
xnor UO_640 (O_640,N_10515,N_12652);
or UO_641 (O_641,N_11978,N_12560);
nor UO_642 (O_642,N_10479,N_12524);
nand UO_643 (O_643,N_13326,N_12775);
xor UO_644 (O_644,N_11153,N_10946);
or UO_645 (O_645,N_14351,N_14892);
xor UO_646 (O_646,N_12055,N_13239);
and UO_647 (O_647,N_10228,N_12250);
nor UO_648 (O_648,N_14714,N_11832);
nand UO_649 (O_649,N_14789,N_10391);
xnor UO_650 (O_650,N_13316,N_13251);
or UO_651 (O_651,N_14669,N_14023);
nor UO_652 (O_652,N_11878,N_11175);
xnor UO_653 (O_653,N_11163,N_11274);
nor UO_654 (O_654,N_11543,N_12451);
xnor UO_655 (O_655,N_11542,N_12030);
xor UO_656 (O_656,N_10979,N_10612);
or UO_657 (O_657,N_14983,N_14651);
nand UO_658 (O_658,N_11458,N_10516);
and UO_659 (O_659,N_14485,N_11794);
nor UO_660 (O_660,N_11777,N_13245);
or UO_661 (O_661,N_11026,N_12068);
and UO_662 (O_662,N_12026,N_12388);
and UO_663 (O_663,N_14616,N_13220);
nor UO_664 (O_664,N_14340,N_12881);
and UO_665 (O_665,N_11447,N_14339);
or UO_666 (O_666,N_11622,N_13225);
and UO_667 (O_667,N_11603,N_14228);
nand UO_668 (O_668,N_10377,N_10416);
nand UO_669 (O_669,N_12050,N_14768);
and UO_670 (O_670,N_13811,N_10055);
or UO_671 (O_671,N_13669,N_12605);
nand UO_672 (O_672,N_13066,N_13563);
xor UO_673 (O_673,N_13607,N_14251);
nor UO_674 (O_674,N_13478,N_10282);
nor UO_675 (O_675,N_12518,N_14148);
nand UO_676 (O_676,N_11720,N_10393);
nand UO_677 (O_677,N_13351,N_10920);
and UO_678 (O_678,N_11237,N_13746);
and UO_679 (O_679,N_11785,N_14490);
nand UO_680 (O_680,N_13417,N_11054);
nand UO_681 (O_681,N_14587,N_11919);
xor UO_682 (O_682,N_10558,N_12621);
and UO_683 (O_683,N_10701,N_12905);
nor UO_684 (O_684,N_14764,N_12713);
xnor UO_685 (O_685,N_14989,N_10023);
nand UO_686 (O_686,N_14466,N_13916);
xor UO_687 (O_687,N_12611,N_10620);
xor UO_688 (O_688,N_10339,N_10241);
and UO_689 (O_689,N_11930,N_13010);
xnor UO_690 (O_690,N_12043,N_11137);
nand UO_691 (O_691,N_13444,N_11305);
xor UO_692 (O_692,N_13059,N_14108);
xor UO_693 (O_693,N_10105,N_10032);
xor UO_694 (O_694,N_14758,N_12900);
xnor UO_695 (O_695,N_14028,N_10755);
or UO_696 (O_696,N_11718,N_10237);
nor UO_697 (O_697,N_13416,N_10904);
nand UO_698 (O_698,N_13849,N_11809);
nor UO_699 (O_699,N_12873,N_10817);
and UO_700 (O_700,N_10455,N_10190);
nor UO_701 (O_701,N_10440,N_13392);
and UO_702 (O_702,N_11941,N_10614);
nand UO_703 (O_703,N_12543,N_11538);
and UO_704 (O_704,N_14810,N_12354);
or UO_705 (O_705,N_14359,N_13324);
nand UO_706 (O_706,N_11117,N_13632);
nand UO_707 (O_707,N_14486,N_14304);
and UO_708 (O_708,N_13726,N_10340);
xnor UO_709 (O_709,N_13354,N_11928);
nand UO_710 (O_710,N_12948,N_10905);
or UO_711 (O_711,N_11655,N_12236);
xor UO_712 (O_712,N_14380,N_10170);
nor UO_713 (O_713,N_12305,N_12548);
nand UO_714 (O_714,N_14536,N_10796);
and UO_715 (O_715,N_12413,N_12704);
or UO_716 (O_716,N_13267,N_14243);
nand UO_717 (O_717,N_12868,N_13079);
and UO_718 (O_718,N_14424,N_10660);
nor UO_719 (O_719,N_12528,N_13524);
xor UO_720 (O_720,N_14922,N_14720);
and UO_721 (O_721,N_11233,N_13435);
or UO_722 (O_722,N_12374,N_14740);
or UO_723 (O_723,N_14037,N_13191);
and UO_724 (O_724,N_13218,N_11628);
nand UO_725 (O_725,N_12565,N_14593);
nand UO_726 (O_726,N_12694,N_12842);
nor UO_727 (O_727,N_11668,N_13577);
or UO_728 (O_728,N_12988,N_12867);
and UO_729 (O_729,N_12440,N_14120);
and UO_730 (O_730,N_10757,N_10038);
and UO_731 (O_731,N_13558,N_10448);
nor UO_732 (O_732,N_11692,N_12654);
nor UO_733 (O_733,N_14041,N_10598);
and UO_734 (O_734,N_12207,N_12320);
or UO_735 (O_735,N_10734,N_12309);
xnor UO_736 (O_736,N_14555,N_13433);
nand UO_737 (O_737,N_10524,N_13634);
or UO_738 (O_738,N_14207,N_13564);
nor UO_739 (O_739,N_13815,N_11258);
xor UO_740 (O_740,N_12357,N_12183);
nor UO_741 (O_741,N_13988,N_14217);
and UO_742 (O_742,N_14384,N_10603);
or UO_743 (O_743,N_11912,N_10923);
and UO_744 (O_744,N_13430,N_12552);
or UO_745 (O_745,N_14996,N_11812);
nand UO_746 (O_746,N_12710,N_13208);
nor UO_747 (O_747,N_11724,N_13290);
nor UO_748 (O_748,N_14668,N_13939);
or UO_749 (O_749,N_14442,N_10925);
nand UO_750 (O_750,N_13901,N_14250);
xnor UO_751 (O_751,N_12641,N_10510);
or UO_752 (O_752,N_10050,N_10083);
and UO_753 (O_753,N_10182,N_14394);
xnor UO_754 (O_754,N_13588,N_12813);
nor UO_755 (O_755,N_14229,N_10235);
and UO_756 (O_756,N_12108,N_13381);
and UO_757 (O_757,N_12588,N_11262);
or UO_758 (O_758,N_13651,N_11206);
or UO_759 (O_759,N_12445,N_13214);
and UO_760 (O_760,N_13708,N_10259);
nor UO_761 (O_761,N_11303,N_13315);
nor UO_762 (O_762,N_14930,N_10324);
nor UO_763 (O_763,N_11569,N_10080);
nor UO_764 (O_764,N_12178,N_12220);
nand UO_765 (O_765,N_10487,N_14366);
or UO_766 (O_766,N_13314,N_10803);
or UO_767 (O_767,N_14338,N_10334);
and UO_768 (O_768,N_11485,N_11076);
or UO_769 (O_769,N_13966,N_13327);
nor UO_770 (O_770,N_14743,N_13212);
xor UO_771 (O_771,N_10031,N_10740);
nor UO_772 (O_772,N_10432,N_14794);
nor UO_773 (O_773,N_13936,N_13468);
or UO_774 (O_774,N_11424,N_14694);
xnor UO_775 (O_775,N_12508,N_13635);
or UO_776 (O_776,N_11844,N_12304);
xnor UO_777 (O_777,N_10581,N_13155);
xor UO_778 (O_778,N_11614,N_14190);
xor UO_779 (O_779,N_12177,N_11088);
nand UO_780 (O_780,N_11326,N_14334);
nand UO_781 (O_781,N_11857,N_10632);
and UO_782 (O_782,N_11817,N_11483);
and UO_783 (O_783,N_11985,N_12671);
nor UO_784 (O_784,N_12499,N_14737);
and UO_785 (O_785,N_11107,N_10529);
and UO_786 (O_786,N_14440,N_13541);
nor UO_787 (O_787,N_12329,N_14452);
xnor UO_788 (O_788,N_12958,N_10859);
xnor UO_789 (O_789,N_10051,N_11381);
nand UO_790 (O_790,N_10390,N_10882);
xnor UO_791 (O_791,N_14484,N_13297);
xnor UO_792 (O_792,N_13215,N_12655);
nor UO_793 (O_793,N_12110,N_14777);
or UO_794 (O_794,N_10355,N_13310);
nand UO_795 (O_795,N_10674,N_14392);
and UO_796 (O_796,N_14509,N_13194);
nor UO_797 (O_797,N_11594,N_13616);
nand UO_798 (O_798,N_10987,N_11905);
nand UO_799 (O_799,N_11134,N_14222);
nand UO_800 (O_800,N_11544,N_12525);
xor UO_801 (O_801,N_11648,N_14537);
nor UO_802 (O_802,N_13887,N_13509);
nand UO_803 (O_803,N_12160,N_11343);
nand UO_804 (O_804,N_11706,N_12628);
xor UO_805 (O_805,N_11666,N_10198);
nand UO_806 (O_806,N_10897,N_14805);
nand UO_807 (O_807,N_12462,N_10641);
xnor UO_808 (O_808,N_13770,N_13597);
nor UO_809 (O_809,N_11704,N_12939);
xor UO_810 (O_810,N_13450,N_14415);
or UO_811 (O_811,N_12576,N_12886);
nor UO_812 (O_812,N_14628,N_13167);
and UO_813 (O_813,N_13745,N_12712);
nor UO_814 (O_814,N_10968,N_12659);
xor UO_815 (O_815,N_11256,N_12251);
nor UO_816 (O_816,N_12507,N_14727);
or UO_817 (O_817,N_14448,N_14759);
and UO_818 (O_818,N_13043,N_11636);
or UO_819 (O_819,N_14688,N_12853);
nand UO_820 (O_820,N_10257,N_12986);
nand UO_821 (O_821,N_12820,N_14624);
or UO_822 (O_822,N_10183,N_10952);
or UO_823 (O_823,N_10735,N_14529);
nand UO_824 (O_824,N_11757,N_12212);
nand UO_825 (O_825,N_14309,N_10372);
xnor UO_826 (O_826,N_12796,N_10421);
and UO_827 (O_827,N_13407,N_13108);
and UO_828 (O_828,N_10852,N_14960);
or UO_829 (O_829,N_14595,N_10719);
nor UO_830 (O_830,N_12714,N_11623);
and UO_831 (O_831,N_11408,N_13926);
nor UO_832 (O_832,N_12698,N_14008);
and UO_833 (O_833,N_10991,N_13806);
xor UO_834 (O_834,N_13900,N_14224);
or UO_835 (O_835,N_13690,N_13888);
xnor UO_836 (O_836,N_14117,N_11299);
and UO_837 (O_837,N_12646,N_10522);
or UO_838 (O_838,N_13880,N_11661);
nor UO_839 (O_839,N_14840,N_12318);
xor UO_840 (O_840,N_10965,N_11365);
and UO_841 (O_841,N_14979,N_13280);
nand UO_842 (O_842,N_13128,N_14093);
nor UO_843 (O_843,N_10489,N_12031);
and UO_844 (O_844,N_10692,N_14019);
nand UO_845 (O_845,N_14505,N_14018);
or UO_846 (O_846,N_12579,N_10865);
or UO_847 (O_847,N_12228,N_11895);
xnor UO_848 (O_848,N_10623,N_10213);
nand UO_849 (O_849,N_11807,N_12831);
nor UO_850 (O_850,N_11098,N_14516);
and UO_851 (O_851,N_12644,N_13115);
and UO_852 (O_852,N_10035,N_14826);
xor UO_853 (O_853,N_13311,N_11552);
nand UO_854 (O_854,N_14594,N_14828);
and UO_855 (O_855,N_11118,N_11813);
xor UO_856 (O_856,N_11038,N_10230);
nand UO_857 (O_857,N_14290,N_11907);
and UO_858 (O_858,N_12491,N_10808);
nor UO_859 (O_859,N_11338,N_11775);
or UO_860 (O_860,N_12854,N_12218);
and UO_861 (O_861,N_10019,N_12802);
nand UO_862 (O_862,N_12167,N_11189);
nor UO_863 (O_863,N_13216,N_14133);
nor UO_864 (O_864,N_14991,N_10993);
and UO_865 (O_865,N_13779,N_10778);
nand UO_866 (O_866,N_13482,N_14665);
and UO_867 (O_867,N_14698,N_14102);
and UO_868 (O_868,N_12224,N_14696);
nand UO_869 (O_869,N_14083,N_13178);
xnor UO_870 (O_870,N_11145,N_13463);
xor UO_871 (O_871,N_11592,N_11730);
xnor UO_872 (O_872,N_10279,N_12750);
and UO_873 (O_873,N_14336,N_10176);
or UO_874 (O_874,N_12828,N_12285);
xnor UO_875 (O_875,N_13285,N_11635);
nor UO_876 (O_876,N_11417,N_13589);
xor UO_877 (O_877,N_13665,N_10060);
or UO_878 (O_878,N_14908,N_10684);
or UO_879 (O_879,N_14273,N_12161);
nand UO_880 (O_880,N_13192,N_13765);
or UO_881 (O_881,N_12909,N_10234);
and UO_882 (O_882,N_11738,N_10787);
xnor UO_883 (O_883,N_12005,N_12373);
xnor UO_884 (O_884,N_12981,N_12280);
xnor UO_885 (O_885,N_13730,N_13086);
and UO_886 (O_886,N_11493,N_10883);
nand UO_887 (O_887,N_12745,N_11358);
and UO_888 (O_888,N_12164,N_10671);
nor UO_889 (O_889,N_11695,N_12010);
and UO_890 (O_890,N_14151,N_14907);
and UO_891 (O_891,N_11558,N_12495);
nor UO_892 (O_892,N_12452,N_12061);
or UO_893 (O_893,N_11843,N_13038);
xnor UO_894 (O_894,N_11318,N_11801);
nand UO_895 (O_895,N_11385,N_10844);
and UO_896 (O_896,N_14796,N_11347);
nand UO_897 (O_897,N_10015,N_10697);
or UO_898 (O_898,N_10477,N_11834);
nor UO_899 (O_899,N_14945,N_10418);
nor UO_900 (O_900,N_10371,N_10625);
and UO_901 (O_901,N_13393,N_11004);
or UO_902 (O_902,N_13827,N_11876);
nor UO_903 (O_903,N_13207,N_10218);
nor UO_904 (O_904,N_14288,N_11999);
xnor UO_905 (O_905,N_10044,N_11737);
or UO_906 (O_906,N_10342,N_11598);
nor UO_907 (O_907,N_11816,N_13475);
and UO_908 (O_908,N_13814,N_11231);
or UO_909 (O_909,N_12155,N_11454);
or UO_910 (O_910,N_13922,N_10984);
nand UO_911 (O_911,N_13051,N_14765);
xnor UO_912 (O_912,N_14590,N_13055);
xor UO_913 (O_913,N_10716,N_11451);
nor UO_914 (O_914,N_13744,N_14940);
and UO_915 (O_915,N_14987,N_10316);
and UO_916 (O_916,N_11147,N_14530);
and UO_917 (O_917,N_13151,N_14589);
xor UO_918 (O_918,N_14526,N_14378);
nor UO_919 (O_919,N_12439,N_12428);
xor UO_920 (O_920,N_13622,N_12738);
xnor UO_921 (O_921,N_14708,N_13306);
or UO_922 (O_922,N_13031,N_14138);
or UO_923 (O_923,N_14377,N_10381);
and UO_924 (O_924,N_11207,N_12148);
and UO_925 (O_925,N_13825,N_11910);
xnor UO_926 (O_926,N_11727,N_11297);
or UO_927 (O_927,N_11627,N_12323);
or UO_928 (O_928,N_10131,N_12444);
nand UO_929 (O_929,N_12736,N_13317);
and UO_930 (O_930,N_13014,N_14857);
nor UO_931 (O_931,N_10554,N_10655);
and UO_932 (O_932,N_11346,N_14216);
xor UO_933 (O_933,N_11375,N_14673);
or UO_934 (O_934,N_12371,N_10895);
nor UO_935 (O_935,N_13008,N_12426);
nand UO_936 (O_936,N_10134,N_10805);
and UO_937 (O_937,N_10344,N_11963);
or UO_938 (O_938,N_12574,N_11740);
nand UO_939 (O_939,N_10397,N_11266);
nand UO_940 (O_940,N_11533,N_10160);
and UO_941 (O_941,N_12838,N_13222);
or UO_942 (O_942,N_10120,N_13962);
nand UO_943 (O_943,N_13978,N_11856);
nor UO_944 (O_944,N_12623,N_14859);
and UO_945 (O_945,N_11780,N_12079);
xor UO_946 (O_946,N_11179,N_10708);
xor UO_947 (O_947,N_14788,N_14558);
and UO_948 (O_948,N_14391,N_13517);
or UO_949 (O_949,N_11914,N_13039);
and UO_950 (O_950,N_11113,N_11534);
or UO_951 (O_951,N_10141,N_12779);
nor UO_952 (O_952,N_14267,N_11768);
or UO_953 (O_953,N_10807,N_13932);
nand UO_954 (O_954,N_13382,N_13162);
xnor UO_955 (O_955,N_11918,N_14799);
and UO_956 (O_956,N_10714,N_10449);
or UO_957 (O_957,N_12034,N_12531);
nand UO_958 (O_958,N_11570,N_12561);
nor UO_959 (O_959,N_13272,N_10729);
or UO_960 (O_960,N_10365,N_11637);
xor UO_961 (O_961,N_14293,N_11624);
and UO_962 (O_962,N_11139,N_14572);
nand UO_963 (O_963,N_13915,N_14234);
nor UO_964 (O_964,N_11021,N_13508);
and UO_965 (O_965,N_10930,N_10885);
nor UO_966 (O_966,N_14710,N_13613);
or UO_967 (O_967,N_13677,N_11419);
and UO_968 (O_968,N_11883,N_10435);
or UO_969 (O_969,N_14943,N_14201);
nand UO_970 (O_970,N_13503,N_12609);
and UO_971 (O_971,N_12956,N_10571);
nand UO_972 (O_972,N_12283,N_12129);
and UO_973 (O_973,N_13732,N_12359);
xor UO_974 (O_974,N_14420,N_14205);
nand UO_975 (O_975,N_12267,N_10917);
nand UO_976 (O_976,N_14381,N_13294);
and UO_977 (O_977,N_14549,N_14285);
nor UO_978 (O_978,N_13758,N_11818);
xnor UO_979 (O_979,N_13072,N_10986);
or UO_980 (O_980,N_11606,N_13830);
and UO_981 (O_981,N_13984,N_10219);
nand UO_982 (O_982,N_13510,N_13643);
xnor UO_983 (O_983,N_11478,N_12829);
or UO_984 (O_984,N_14266,N_14755);
or UO_985 (O_985,N_13938,N_11871);
and UO_986 (O_986,N_14079,N_13974);
xnor UO_987 (O_987,N_13700,N_12091);
nand UO_988 (O_988,N_14269,N_11230);
xor UO_989 (O_989,N_13689,N_14461);
or UO_990 (O_990,N_14111,N_14656);
and UO_991 (O_991,N_13910,N_10978);
nor UO_992 (O_992,N_10916,N_10836);
nor UO_993 (O_993,N_13007,N_14762);
nor UO_994 (O_994,N_14776,N_11406);
and UO_995 (O_995,N_13742,N_10140);
nand UO_996 (O_996,N_12302,N_10748);
xor UO_997 (O_997,N_10075,N_14100);
nor UO_998 (O_998,N_10499,N_10046);
xnor UO_999 (O_999,N_12624,N_13165);
nor UO_1000 (O_1000,N_12540,N_11887);
and UO_1001 (O_1001,N_10644,N_13767);
xnor UO_1002 (O_1002,N_13705,N_13350);
nand UO_1003 (O_1003,N_14770,N_12425);
xor UO_1004 (O_1004,N_10999,N_14202);
and UO_1005 (O_1005,N_13560,N_10194);
and UO_1006 (O_1006,N_11953,N_13592);
xor UO_1007 (O_1007,N_10507,N_13969);
nand UO_1008 (O_1008,N_14115,N_10642);
nand UO_1009 (O_1009,N_13928,N_11567);
xnor UO_1010 (O_1010,N_14323,N_11959);
or UO_1011 (O_1011,N_11915,N_13061);
and UO_1012 (O_1012,N_13897,N_14414);
xor UO_1013 (O_1013,N_10442,N_14641);
nor UO_1014 (O_1014,N_13132,N_14579);
nor UO_1015 (O_1015,N_12814,N_10309);
or UO_1016 (O_1016,N_12771,N_12737);
or UO_1017 (O_1017,N_14565,N_11070);
xnor UO_1018 (O_1018,N_14483,N_14503);
xor UO_1019 (O_1019,N_13489,N_13739);
or UO_1020 (O_1020,N_14437,N_13111);
or UO_1021 (O_1021,N_14349,N_12265);
nand UO_1022 (O_1022,N_12700,N_13243);
nor UO_1023 (O_1023,N_13840,N_11404);
xor UO_1024 (O_1024,N_10000,N_11323);
and UO_1025 (O_1025,N_12483,N_13836);
nor UO_1026 (O_1026,N_12238,N_13774);
nand UO_1027 (O_1027,N_14126,N_13445);
and UO_1028 (O_1028,N_10944,N_11302);
xnor UO_1029 (O_1029,N_11770,N_14998);
xor UO_1030 (O_1030,N_11248,N_14210);
and UO_1031 (O_1031,N_13914,N_10248);
or UO_1032 (O_1032,N_11446,N_14230);
xnor UO_1033 (O_1033,N_13668,N_14493);
or UO_1034 (O_1034,N_14231,N_11386);
xor UO_1035 (O_1035,N_14813,N_13189);
xor UO_1036 (O_1036,N_10345,N_14670);
nand UO_1037 (O_1037,N_14195,N_13018);
nand UO_1038 (O_1038,N_11610,N_12436);
nor UO_1039 (O_1039,N_13725,N_14150);
and UO_1040 (O_1040,N_12955,N_12570);
nor UO_1041 (O_1041,N_12866,N_10356);
nand UO_1042 (O_1042,N_13217,N_13921);
nand UO_1043 (O_1043,N_12512,N_14013);
or UO_1044 (O_1044,N_14679,N_11988);
xnor UO_1045 (O_1045,N_11778,N_12546);
nand UO_1046 (O_1046,N_10013,N_14849);
or UO_1047 (O_1047,N_14390,N_14281);
nor UO_1048 (O_1048,N_10293,N_14938);
nor UO_1049 (O_1049,N_13219,N_11036);
xnor UO_1050 (O_1050,N_12385,N_11120);
xor UO_1051 (O_1051,N_12990,N_12327);
nand UO_1052 (O_1052,N_12892,N_13246);
xnor UO_1053 (O_1053,N_13983,N_11349);
nor UO_1054 (O_1054,N_12060,N_12075);
nand UO_1055 (O_1055,N_14793,N_12785);
xor UO_1056 (O_1056,N_12315,N_11572);
and UO_1057 (O_1057,N_11197,N_12889);
xnor UO_1058 (O_1058,N_11644,N_11885);
nor UO_1059 (O_1059,N_11009,N_12636);
or UO_1060 (O_1060,N_10680,N_10961);
xor UO_1061 (O_1061,N_10107,N_11916);
nand UO_1062 (O_1062,N_10795,N_12415);
or UO_1063 (O_1063,N_10681,N_14961);
nor UO_1064 (O_1064,N_12857,N_11393);
nand UO_1065 (O_1065,N_10709,N_10881);
nor UO_1066 (O_1066,N_11924,N_11530);
or UO_1067 (O_1067,N_14209,N_11423);
and UO_1068 (O_1068,N_10559,N_10064);
xnor UO_1069 (O_1069,N_14128,N_12186);
or UO_1070 (O_1070,N_12206,N_11041);
nor UO_1071 (O_1071,N_11886,N_14314);
and UO_1072 (O_1072,N_14502,N_12067);
xor UO_1073 (O_1073,N_12987,N_14968);
xnor UO_1074 (O_1074,N_10474,N_10215);
and UO_1075 (O_1075,N_13673,N_13646);
and UO_1076 (O_1076,N_12299,N_10963);
or UO_1077 (O_1077,N_12396,N_12249);
nand UO_1078 (O_1078,N_13348,N_10003);
xor UO_1079 (O_1079,N_14495,N_10362);
or UO_1080 (O_1080,N_14441,N_14569);
nor UO_1081 (O_1081,N_12430,N_12443);
nand UO_1082 (O_1082,N_14966,N_14633);
or UO_1083 (O_1083,N_14477,N_12389);
or UO_1084 (O_1084,N_11820,N_10821);
nand UO_1085 (O_1085,N_10475,N_12264);
xor UO_1086 (O_1086,N_10375,N_13997);
or UO_1087 (O_1087,N_10588,N_13149);
and UO_1088 (O_1088,N_13826,N_10382);
nor UO_1089 (O_1089,N_10953,N_11469);
or UO_1090 (O_1090,N_13420,N_11526);
and UO_1091 (O_1091,N_13605,N_14443);
nand UO_1092 (O_1092,N_10126,N_14842);
or UO_1093 (O_1093,N_11213,N_14194);
xor UO_1094 (O_1094,N_11205,N_10700);
and UO_1095 (O_1095,N_11194,N_14607);
xnor UO_1096 (O_1096,N_11131,N_14187);
xor UO_1097 (O_1097,N_11583,N_12254);
and UO_1098 (O_1098,N_14056,N_13201);
or UO_1099 (O_1099,N_12979,N_11405);
and UO_1100 (O_1100,N_10145,N_13717);
nor UO_1101 (O_1101,N_10935,N_14372);
nand UO_1102 (O_1102,N_12703,N_12551);
nor UO_1103 (O_1103,N_11944,N_10100);
xnor UO_1104 (O_1104,N_10725,N_11566);
and UO_1105 (O_1105,N_12166,N_10364);
or UO_1106 (O_1106,N_13454,N_14014);
nand UO_1107 (O_1107,N_11705,N_10084);
and UO_1108 (O_1108,N_12959,N_14584);
nor UO_1109 (O_1109,N_13298,N_13044);
nor UO_1110 (O_1110,N_14246,N_12630);
nor UO_1111 (O_1111,N_10896,N_14803);
or UO_1112 (O_1112,N_11428,N_12209);
and UO_1113 (O_1113,N_10751,N_10263);
nor UO_1114 (O_1114,N_11851,N_13292);
and UO_1115 (O_1115,N_11656,N_14239);
xor UO_1116 (O_1116,N_14208,N_13536);
and UO_1117 (O_1117,N_13998,N_13766);
nor UO_1118 (O_1118,N_12797,N_12887);
nor UO_1119 (O_1119,N_13623,N_10617);
nand UO_1120 (O_1120,N_14077,N_11647);
nor UO_1121 (O_1121,N_13144,N_14308);
and UO_1122 (O_1122,N_11793,N_10887);
xor UO_1123 (O_1123,N_10613,N_10501);
nor UO_1124 (O_1124,N_13776,N_13455);
nor UO_1125 (O_1125,N_14661,N_11140);
nand UO_1126 (O_1126,N_11512,N_12027);
nor UO_1127 (O_1127,N_14435,N_10225);
nor UO_1128 (O_1128,N_11703,N_14244);
nand UO_1129 (O_1129,N_12331,N_10287);
nand UO_1130 (O_1130,N_11989,N_11355);
or UO_1131 (O_1131,N_10823,N_12809);
nand UO_1132 (O_1132,N_11119,N_13805);
xnor UO_1133 (O_1133,N_10659,N_10285);
nand UO_1134 (O_1134,N_12294,N_12915);
nand UO_1135 (O_1135,N_11940,N_10203);
nor UO_1136 (O_1136,N_11532,N_14007);
or UO_1137 (O_1137,N_11133,N_14425);
nand UO_1138 (O_1138,N_12613,N_10146);
or UO_1139 (O_1139,N_10491,N_13571);
nor UO_1140 (O_1140,N_12850,N_14433);
nand UO_1141 (O_1141,N_12128,N_11202);
or UO_1142 (O_1142,N_11991,N_12119);
nor UO_1143 (O_1143,N_12963,N_14889);
nor UO_1144 (O_1144,N_12994,N_10132);
and UO_1145 (O_1145,N_12355,N_11935);
and UO_1146 (O_1146,N_13959,N_10301);
and UO_1147 (O_1147,N_13832,N_10081);
xnor UO_1148 (O_1148,N_10043,N_14130);
and UO_1149 (O_1149,N_13400,N_13750);
nor UO_1150 (O_1150,N_14184,N_10464);
xnor UO_1151 (O_1151,N_10797,N_11965);
or UO_1152 (O_1152,N_13042,N_14937);
nand UO_1153 (O_1153,N_13964,N_13790);
and UO_1154 (O_1154,N_12633,N_13341);
or UO_1155 (O_1155,N_10222,N_13781);
or UO_1156 (O_1156,N_11158,N_12258);
and UO_1157 (O_1157,N_12993,N_10062);
xor UO_1158 (O_1158,N_10407,N_12012);
xor UO_1159 (O_1159,N_11295,N_10159);
or UO_1160 (O_1160,N_11040,N_10948);
xnor UO_1161 (O_1161,N_12014,N_14426);
nand UO_1162 (O_1162,N_11467,N_10988);
and UO_1163 (O_1163,N_10593,N_11600);
nand UO_1164 (O_1164,N_11509,N_12295);
and UO_1165 (O_1165,N_11384,N_11756);
and UO_1166 (O_1166,N_11504,N_12835);
nor UO_1167 (O_1167,N_14990,N_10802);
nand UO_1168 (O_1168,N_14472,N_10590);
and UO_1169 (O_1169,N_10976,N_12758);
nor UO_1170 (O_1170,N_10648,N_10949);
xor UO_1171 (O_1171,N_12755,N_13268);
and UO_1172 (O_1172,N_12660,N_14871);
nand UO_1173 (O_1173,N_10212,N_12541);
and UO_1174 (O_1174,N_12851,N_10130);
or UO_1175 (O_1175,N_10040,N_13572);
or UO_1176 (O_1176,N_14388,N_10857);
and UO_1177 (O_1177,N_11650,N_11010);
xnor UO_1178 (O_1178,N_14872,N_10308);
nor UO_1179 (O_1179,N_12480,N_11097);
nand UO_1180 (O_1180,N_12169,N_12665);
nor UO_1181 (O_1181,N_12648,N_10520);
nand UO_1182 (O_1182,N_14305,N_10595);
xor UO_1183 (O_1183,N_13056,N_10071);
and UO_1184 (O_1184,N_14460,N_11633);
and UO_1185 (O_1185,N_10577,N_10242);
nor UO_1186 (O_1186,N_13322,N_10193);
or UO_1187 (O_1187,N_11761,N_11539);
nor UO_1188 (O_1188,N_12242,N_13875);
and UO_1189 (O_1189,N_14347,N_10957);
and UO_1190 (O_1190,N_11223,N_13228);
xor UO_1191 (O_1191,N_13484,N_10628);
nand UO_1192 (O_1192,N_14801,N_14171);
nand UO_1193 (O_1193,N_11620,N_14625);
nand UO_1194 (O_1194,N_12592,N_11589);
or UO_1195 (O_1195,N_12421,N_14236);
nand UO_1196 (O_1196,N_11774,N_12021);
nand UO_1197 (O_1197,N_14481,N_10608);
nand UO_1198 (O_1198,N_11245,N_10447);
xor UO_1199 (O_1199,N_14559,N_10379);
nor UO_1200 (O_1200,N_13487,N_14932);
xnor UO_1201 (O_1201,N_12510,N_12376);
and UO_1202 (O_1202,N_11327,N_11714);
and UO_1203 (O_1203,N_11854,N_11970);
nor UO_1204 (O_1204,N_13604,N_12618);
nor UO_1205 (O_1205,N_14024,N_11893);
and UO_1206 (O_1206,N_12870,N_13747);
xor UO_1207 (O_1207,N_12019,N_12170);
and UO_1208 (O_1208,N_13507,N_13567);
and UO_1209 (O_1209,N_14219,N_11225);
or UO_1210 (O_1210,N_13578,N_12684);
or UO_1211 (O_1211,N_11255,N_10096);
nor UO_1212 (O_1212,N_10557,N_12522);
nor UO_1213 (O_1213,N_11353,N_12582);
and UO_1214 (O_1214,N_10164,N_14847);
nor UO_1215 (O_1215,N_14583,N_12759);
xor UO_1216 (O_1216,N_10138,N_11191);
and UO_1217 (O_1217,N_14886,N_11270);
or UO_1218 (O_1218,N_11214,N_10861);
xor UO_1219 (O_1219,N_10556,N_11612);
or UO_1220 (O_1220,N_11607,N_11599);
nand UO_1221 (O_1221,N_13975,N_12875);
or UO_1222 (O_1222,N_13903,N_11217);
nand UO_1223 (O_1223,N_13136,N_13857);
xnor UO_1224 (O_1224,N_13198,N_13838);
nor UO_1225 (O_1225,N_11689,N_13784);
xor UO_1226 (O_1226,N_12760,N_12145);
xnor UO_1227 (O_1227,N_10911,N_10353);
nor UO_1228 (O_1228,N_14436,N_10093);
and UO_1229 (O_1229,N_14575,N_11221);
xor UO_1230 (O_1230,N_12788,N_14375);
xnor UO_1231 (O_1231,N_13123,N_10366);
or UO_1232 (O_1232,N_10114,N_12383);
and UO_1233 (O_1233,N_13752,N_13876);
and UO_1234 (O_1234,N_12077,N_13584);
nand UO_1235 (O_1235,N_14606,N_12353);
or UO_1236 (O_1236,N_12417,N_12072);
xor UO_1237 (O_1237,N_13550,N_10958);
nor UO_1238 (O_1238,N_11608,N_12380);
and UO_1239 (O_1239,N_10966,N_12573);
nor UO_1240 (O_1240,N_12519,N_12716);
and UO_1241 (O_1241,N_12022,N_12537);
nor UO_1242 (O_1242,N_14873,N_11911);
or UO_1243 (O_1243,N_10461,N_12088);
nor UO_1244 (O_1244,N_10402,N_12678);
and UO_1245 (O_1245,N_14678,N_11067);
or UO_1246 (O_1246,N_14519,N_11559);
or UO_1247 (O_1247,N_10884,N_10274);
and UO_1248 (O_1248,N_13126,N_13492);
and UO_1249 (O_1249,N_12087,N_10469);
and UO_1250 (O_1250,N_12492,N_12479);
xnor UO_1251 (O_1251,N_12494,N_11058);
or UO_1252 (O_1252,N_11362,N_13264);
xnor UO_1253 (O_1253,N_11669,N_14268);
and UO_1254 (O_1254,N_12247,N_13190);
xnor UO_1255 (O_1255,N_12184,N_13134);
nor UO_1256 (O_1256,N_11460,N_11005);
nand UO_1257 (O_1257,N_13893,N_13206);
and UO_1258 (O_1258,N_14581,N_10869);
nor UO_1259 (O_1259,N_12168,N_10415);
and UO_1260 (O_1260,N_10411,N_14116);
or UO_1261 (O_1261,N_14701,N_11331);
xor UO_1262 (O_1262,N_10536,N_14636);
nand UO_1263 (O_1263,N_10839,N_14031);
nand UO_1264 (O_1264,N_13147,N_10057);
nand UO_1265 (O_1265,N_11993,N_11555);
and UO_1266 (O_1266,N_10463,N_10866);
and UO_1267 (O_1267,N_14896,N_11952);
xnor UO_1268 (O_1268,N_12718,N_14642);
and UO_1269 (O_1269,N_13628,N_11662);
or UO_1270 (O_1270,N_12312,N_13626);
or UO_1271 (O_1271,N_14576,N_11717);
nor UO_1272 (O_1272,N_10412,N_14047);
nor UO_1273 (O_1273,N_11491,N_11889);
and UO_1274 (O_1274,N_11507,N_12112);
xor UO_1275 (O_1275,N_12146,N_13401);
or UO_1276 (O_1276,N_10853,N_12989);
and UO_1277 (O_1277,N_13495,N_13464);
nor UO_1278 (O_1278,N_14213,N_14704);
nor UO_1279 (O_1279,N_10327,N_12921);
xor UO_1280 (O_1280,N_13090,N_13519);
xor UO_1281 (O_1281,N_13103,N_14010);
xnor UO_1282 (O_1282,N_13221,N_11148);
nand UO_1283 (O_1283,N_13546,N_11659);
nand UO_1284 (O_1284,N_11235,N_13769);
or UO_1285 (O_1285,N_14459,N_13547);
and UO_1286 (O_1286,N_10826,N_14084);
or UO_1287 (O_1287,N_10124,N_11135);
nor UO_1288 (O_1288,N_10784,N_11833);
and UO_1289 (O_1289,N_13823,N_13955);
nor UO_1290 (O_1290,N_10828,N_10723);
and UO_1291 (O_1291,N_12418,N_10527);
nor UO_1292 (O_1292,N_13016,N_13431);
and UO_1293 (O_1293,N_14550,N_10947);
xnor UO_1294 (O_1294,N_13004,N_12435);
or UO_1295 (O_1295,N_11246,N_10583);
or UO_1296 (O_1296,N_11463,N_13440);
nor UO_1297 (O_1297,N_10793,N_14476);
xor UO_1298 (O_1298,N_12597,N_14852);
nand UO_1299 (O_1299,N_13153,N_10814);
or UO_1300 (O_1300,N_11499,N_11313);
and UO_1301 (O_1301,N_14025,N_13425);
nor UO_1302 (O_1302,N_10466,N_13046);
xnor UO_1303 (O_1303,N_14081,N_13397);
or UO_1304 (O_1304,N_14525,N_12080);
nor UO_1305 (O_1305,N_14986,N_14969);
nor UO_1306 (O_1306,N_13394,N_12308);
or UO_1307 (O_1307,N_12049,N_12141);
nor UO_1308 (O_1308,N_11760,N_13494);
nand UO_1309 (O_1309,N_11164,N_10139);
nand UO_1310 (O_1310,N_12352,N_14662);
nand UO_1311 (O_1311,N_13036,N_13837);
nand UO_1312 (O_1312,N_11678,N_10041);
nor UO_1313 (O_1313,N_14570,N_11746);
xor UO_1314 (O_1314,N_13481,N_10498);
nor UO_1315 (O_1315,N_11061,N_14664);
xnor UO_1316 (O_1316,N_10871,N_10252);
and UO_1317 (O_1317,N_12637,N_13590);
or UO_1318 (O_1318,N_11990,N_14350);
nor UO_1319 (O_1319,N_10591,N_11141);
nor UO_1320 (O_1320,N_10296,N_10841);
nor UO_1321 (O_1321,N_10605,N_10703);
xor UO_1322 (O_1322,N_10800,N_13924);
or UO_1323 (O_1323,N_10488,N_10220);
or UO_1324 (O_1324,N_12095,N_13068);
nor UO_1325 (O_1325,N_12001,N_10434);
and UO_1326 (O_1326,N_11159,N_10615);
or UO_1327 (O_1327,N_10380,N_12400);
nor UO_1328 (O_1328,N_14763,N_13070);
nor UO_1329 (O_1329,N_14950,N_11111);
nand UO_1330 (O_1330,N_14807,N_11083);
nand UO_1331 (O_1331,N_13637,N_13022);
nor UO_1332 (O_1332,N_11015,N_13582);
nor UO_1333 (O_1333,N_14953,N_11808);
xnor UO_1334 (O_1334,N_13226,N_13017);
or UO_1335 (O_1335,N_12769,N_12450);
nand UO_1336 (O_1336,N_12422,N_14121);
and UO_1337 (O_1337,N_13872,N_14456);
nor UO_1338 (O_1338,N_13497,N_10478);
nand UO_1339 (O_1339,N_11540,N_12409);
nor UO_1340 (O_1340,N_11574,N_13618);
nor UO_1341 (O_1341,N_11222,N_13617);
nor UO_1342 (O_1342,N_10110,N_11394);
or UO_1343 (O_1343,N_13284,N_14406);
nand UO_1344 (O_1344,N_13789,N_13537);
nor UO_1345 (O_1345,N_11613,N_11192);
or UO_1346 (O_1346,N_13364,N_11979);
nand UO_1347 (O_1347,N_13172,N_14511);
nor UO_1348 (O_1348,N_14174,N_11649);
xnor UO_1349 (O_1349,N_11709,N_10901);
or UO_1350 (O_1350,N_11956,N_11877);
and UO_1351 (O_1351,N_13797,N_14161);
nand UO_1352 (O_1352,N_13281,N_12719);
nand UO_1353 (O_1353,N_13919,N_11275);
xor UO_1354 (O_1354,N_11315,N_11016);
nor UO_1355 (O_1355,N_10231,N_14197);
nor UO_1356 (O_1356,N_14240,N_11966);
xor UO_1357 (O_1357,N_13831,N_11443);
nand UO_1358 (O_1358,N_11280,N_12201);
nand UO_1359 (O_1359,N_14192,N_14911);
xnor UO_1360 (O_1360,N_12277,N_14650);
nor UO_1361 (O_1361,N_13967,N_12910);
xnor UO_1362 (O_1362,N_14276,N_14155);
nand UO_1363 (O_1363,N_11367,N_13609);
xnor UO_1364 (O_1364,N_10321,N_14541);
nand UO_1365 (O_1365,N_11195,N_10157);
or UO_1366 (O_1366,N_13048,N_13566);
xor UO_1367 (O_1367,N_11936,N_12406);
xor UO_1368 (O_1368,N_13953,N_12944);
and UO_1369 (O_1369,N_11388,N_10599);
nand UO_1370 (O_1370,N_13639,N_10076);
nand UO_1371 (O_1371,N_11591,N_14677);
and UO_1372 (O_1372,N_11731,N_14374);
and UO_1373 (O_1373,N_13960,N_11085);
nand UO_1374 (O_1374,N_14728,N_13019);
and UO_1375 (O_1375,N_11403,N_13612);
nand UO_1376 (O_1376,N_10485,N_14544);
nor UO_1377 (O_1377,N_12961,N_13786);
or UO_1378 (O_1378,N_12369,N_12756);
and UO_1379 (O_1379,N_13762,N_11824);
and UO_1380 (O_1380,N_11880,N_10907);
xnor UO_1381 (O_1381,N_12203,N_14856);
nor UO_1382 (O_1382,N_10929,N_10504);
or UO_1383 (O_1383,N_10967,N_10053);
or UO_1384 (O_1384,N_13349,N_12638);
xor UO_1385 (O_1385,N_14752,N_11596);
xor UO_1386 (O_1386,N_10090,N_14464);
nand UO_1387 (O_1387,N_13467,N_14344);
and UO_1388 (O_1388,N_14179,N_12970);
nand UO_1389 (O_1389,N_13140,N_12612);
and UO_1390 (O_1390,N_14610,N_12488);
nor UO_1391 (O_1391,N_10201,N_14098);
nor UO_1392 (O_1392,N_10940,N_11045);
or UO_1393 (O_1393,N_14473,N_10580);
or UO_1394 (O_1394,N_12137,N_11961);
or UO_1395 (O_1395,N_13864,N_12321);
nand UO_1396 (O_1396,N_14588,N_14795);
or UO_1397 (O_1397,N_12360,N_10026);
nor UO_1398 (O_1398,N_13037,N_13882);
nand UO_1399 (O_1399,N_13561,N_13258);
nor UO_1400 (O_1400,N_13107,N_11409);
xnor UO_1401 (O_1401,N_12132,N_12765);
nand UO_1402 (O_1402,N_10574,N_13045);
nand UO_1403 (O_1403,N_14721,N_14732);
nor UO_1404 (O_1404,N_11236,N_13161);
xor UO_1405 (O_1405,N_12726,N_11955);
or UO_1406 (O_1406,N_13457,N_10876);
xnor UO_1407 (O_1407,N_11969,N_12176);
or UO_1408 (O_1408,N_14512,N_12100);
nand UO_1409 (O_1409,N_11116,N_12679);
nand UO_1410 (O_1410,N_14617,N_13380);
or UO_1411 (O_1411,N_11167,N_10360);
nor UO_1412 (O_1412,N_10426,N_12231);
nor UO_1413 (O_1413,N_11208,N_10955);
xor UO_1414 (O_1414,N_14683,N_12965);
and UO_1415 (O_1415,N_13756,N_10772);
nand UO_1416 (O_1416,N_10969,N_12446);
and UO_1417 (O_1417,N_10472,N_10733);
and UO_1418 (O_1418,N_11368,N_10845);
nor UO_1419 (O_1419,N_13846,N_10239);
and UO_1420 (O_1420,N_10262,N_13780);
xnor UO_1421 (O_1421,N_14880,N_11858);
and UO_1422 (O_1422,N_11373,N_10653);
or UO_1423 (O_1423,N_11500,N_12015);
nor UO_1424 (O_1424,N_14032,N_12784);
nor UO_1425 (O_1425,N_11281,N_10052);
and UO_1426 (O_1426,N_11957,N_14982);
nand UO_1427 (O_1427,N_10226,N_10870);
nor UO_1428 (O_1428,N_11729,N_12515);
or UO_1429 (O_1429,N_13185,N_14455);
xor UO_1430 (O_1430,N_10240,N_13862);
nor UO_1431 (O_1431,N_12930,N_11616);
and UO_1432 (O_1432,N_12361,N_10690);
nand UO_1433 (O_1433,N_12806,N_12555);
nand UO_1434 (O_1434,N_11024,N_12899);
and UO_1435 (O_1435,N_10310,N_11725);
xnor UO_1436 (O_1436,N_10639,N_14324);
xnor UO_1437 (O_1437,N_13282,N_12126);
nor UO_1438 (O_1438,N_14225,N_13676);
or UO_1439 (O_1439,N_12542,N_10142);
nor UO_1440 (O_1440,N_13462,N_11378);
nand UO_1441 (O_1441,N_10818,N_14453);
xnor UO_1442 (O_1442,N_12130,N_13502);
nand UO_1443 (O_1443,N_12377,N_14778);
or UO_1444 (O_1444,N_13971,N_12969);
and UO_1445 (O_1445,N_10600,N_12926);
and UO_1446 (O_1446,N_13958,N_13204);
and UO_1447 (O_1447,N_14089,N_12065);
nor UO_1448 (O_1448,N_14733,N_12175);
nor UO_1449 (O_1449,N_11582,N_12962);
nor UO_1450 (O_1450,N_10627,N_11541);
nand UO_1451 (O_1451,N_11836,N_10108);
nor UO_1452 (O_1452,N_10683,N_12966);
nor UO_1453 (O_1453,N_11839,N_14808);
and UO_1454 (O_1454,N_10685,N_14814);
nor UO_1455 (O_1455,N_14354,N_10453);
nor UO_1456 (O_1456,N_14306,N_11272);
or UO_1457 (O_1457,N_14596,N_14995);
xor UO_1458 (O_1458,N_14690,N_13157);
xor UO_1459 (O_1459,N_10033,N_14931);
or UO_1460 (O_1460,N_11336,N_11069);
xnor UO_1461 (O_1461,N_14356,N_13721);
and UO_1462 (O_1462,N_13256,N_12500);
nor UO_1463 (O_1463,N_10329,N_10596);
or UO_1464 (O_1464,N_10350,N_13748);
or UO_1465 (O_1465,N_12791,N_11764);
and UO_1466 (O_1466,N_10939,N_10502);
nand UO_1467 (O_1467,N_10970,N_13175);
xnor UO_1468 (O_1468,N_12513,N_14640);
nand UO_1469 (O_1469,N_14160,N_11520);
and UO_1470 (O_1470,N_10573,N_14034);
or UO_1471 (O_1471,N_14131,N_11982);
xnor UO_1472 (O_1472,N_12136,N_11395);
nand UO_1473 (O_1473,N_13530,N_10611);
or UO_1474 (O_1474,N_10028,N_11711);
nor UO_1475 (O_1475,N_13230,N_14458);
nor UO_1476 (O_1476,N_10278,N_10167);
nor UO_1477 (O_1477,N_13843,N_11122);
xnor UO_1478 (O_1478,N_12364,N_12370);
nor UO_1479 (O_1479,N_12901,N_12668);
or UO_1480 (O_1480,N_11867,N_10483);
and UO_1481 (O_1481,N_11641,N_12270);
or UO_1482 (O_1482,N_13081,N_12372);
nor UO_1483 (O_1483,N_11400,N_11593);
or UO_1484 (O_1484,N_10172,N_11506);
xnor UO_1485 (O_1485,N_12282,N_14923);
xnor UO_1486 (O_1486,N_14482,N_13145);
and UO_1487 (O_1487,N_11014,N_13302);
xnor UO_1488 (O_1488,N_12035,N_14812);
xnor UO_1489 (O_1489,N_12289,N_11846);
and UO_1490 (O_1490,N_14649,N_13585);
and UO_1491 (O_1491,N_10912,N_12038);
nor UO_1492 (O_1492,N_10908,N_14839);
nor UO_1493 (O_1493,N_14809,N_11719);
or UO_1494 (O_1494,N_14095,N_11934);
nand UO_1495 (O_1495,N_14134,N_12078);
or UO_1496 (O_1496,N_13816,N_14949);
nor UO_1497 (O_1497,N_11862,N_13011);
or UO_1498 (O_1498,N_14178,N_12933);
nor UO_1499 (O_1499,N_11185,N_11702);
or UO_1500 (O_1500,N_10454,N_12057);
nand UO_1501 (O_1501,N_11279,N_10020);
and UO_1502 (O_1502,N_10753,N_14400);
nor UO_1503 (O_1503,N_12985,N_10288);
and UO_1504 (O_1504,N_14864,N_14364);
xor UO_1505 (O_1505,N_11311,N_10061);
nand UO_1506 (O_1506,N_14580,N_11722);
and UO_1507 (O_1507,N_12923,N_12083);
or UO_1508 (O_1508,N_10931,N_11758);
nand UO_1509 (O_1509,N_12688,N_13429);
and UO_1510 (O_1510,N_13661,N_11334);
xnor UO_1511 (O_1511,N_12094,N_12973);
and UO_1512 (O_1512,N_13506,N_12545);
xnor UO_1513 (O_1513,N_13852,N_11459);
or UO_1514 (O_1514,N_13385,N_13935);
nand UO_1515 (O_1515,N_10482,N_12982);
xor UO_1516 (O_1516,N_12466,N_11994);
nor UO_1517 (O_1517,N_10205,N_13296);
and UO_1518 (O_1518,N_10443,N_13678);
nand UO_1519 (O_1519,N_10832,N_10408);
or UO_1520 (O_1520,N_12649,N_12255);
xor UO_1521 (O_1521,N_11806,N_13647);
nand UO_1522 (O_1522,N_14760,N_11852);
or UO_1523 (O_1523,N_12590,N_12476);
or UO_1524 (O_1524,N_13176,N_14802);
nor UO_1525 (O_1525,N_13514,N_10425);
or UO_1526 (O_1526,N_14284,N_13288);
nand UO_1527 (O_1527,N_10008,N_10825);
xnor UO_1528 (O_1528,N_10017,N_11602);
nor UO_1529 (O_1529,N_14183,N_14510);
nand UO_1530 (O_1530,N_12240,N_14410);
or UO_1531 (O_1531,N_13535,N_13360);
or UO_1532 (O_1532,N_14734,N_12547);
or UO_1533 (O_1533,N_13427,N_14445);
xnor UO_1534 (O_1534,N_13186,N_10162);
nand UO_1535 (O_1535,N_13421,N_11110);
nand UO_1536 (O_1536,N_14398,N_11980);
xnor UO_1537 (O_1537,N_12182,N_12735);
and UO_1538 (O_1538,N_11374,N_14562);
nor UO_1539 (O_1539,N_10737,N_14492);
xor UO_1540 (O_1540,N_11190,N_11146);
nor UO_1541 (O_1541,N_12469,N_13731);
or UO_1542 (O_1542,N_14786,N_14478);
xnor UO_1543 (O_1543,N_11618,N_14454);
nand UO_1544 (O_1544,N_12408,N_13533);
nand UO_1545 (O_1545,N_12188,N_14699);
or UO_1546 (O_1546,N_10813,N_10208);
nand UO_1547 (O_1547,N_13516,N_14784);
nand UO_1548 (O_1548,N_13183,N_13460);
nand UO_1549 (O_1549,N_13569,N_11238);
and UO_1550 (O_1550,N_12217,N_11619);
xor UO_1551 (O_1551,N_13428,N_14412);
nand UO_1552 (O_1552,N_13456,N_10185);
and UO_1553 (O_1553,N_11735,N_14912);
or UO_1554 (O_1554,N_12935,N_13684);
and UO_1555 (O_1555,N_13735,N_10007);
nor UO_1556 (O_1556,N_11324,N_13804);
xor UO_1557 (O_1557,N_14277,N_14376);
xnor UO_1558 (O_1558,N_13247,N_11621);
and UO_1559 (O_1559,N_14528,N_12018);
and UO_1560 (O_1560,N_10445,N_14540);
nor UO_1561 (O_1561,N_10118,N_12348);
xor UO_1562 (O_1562,N_12458,N_14869);
nor UO_1563 (O_1563,N_10315,N_11314);
or UO_1564 (O_1564,N_12465,N_13486);
and UO_1565 (O_1565,N_11407,N_12020);
and UO_1566 (O_1566,N_12292,N_13667);
and UO_1567 (O_1567,N_13331,N_12584);
nand UO_1568 (O_1568,N_12774,N_13164);
nor UO_1569 (O_1569,N_14189,N_11162);
nor UO_1570 (O_1570,N_10276,N_11050);
or UO_1571 (O_1571,N_12904,N_12949);
nor UO_1572 (O_1572,N_11287,N_10514);
or UO_1573 (O_1573,N_12468,N_11835);
nand UO_1574 (O_1574,N_13865,N_13318);
xor UO_1575 (O_1575,N_10566,N_12241);
and UO_1576 (O_1576,N_12999,N_10281);
nand UO_1577 (O_1577,N_10460,N_13335);
and UO_1578 (O_1578,N_12917,N_14603);
xnor UO_1579 (O_1579,N_10204,N_10610);
nand UO_1580 (O_1580,N_13874,N_10541);
and UO_1581 (O_1581,N_13224,N_13598);
nand UO_1582 (O_1582,N_12081,N_11027);
nand UO_1583 (O_1583,N_10195,N_14514);
xnor UO_1584 (O_1584,N_13159,N_10103);
xor UO_1585 (O_1585,N_12883,N_12273);
xnor UO_1586 (O_1586,N_13845,N_11301);
or UO_1587 (O_1587,N_11875,N_13741);
or UO_1588 (O_1588,N_11906,N_14085);
and UO_1589 (O_1589,N_12762,N_14393);
nor UO_1590 (O_1590,N_12658,N_14779);
nand UO_1591 (O_1591,N_13855,N_12968);
nor UO_1592 (O_1592,N_14043,N_12732);
nand UO_1593 (O_1593,N_10809,N_12484);
nor UO_1594 (O_1594,N_11127,N_13069);
xnor UO_1595 (O_1595,N_12805,N_12918);
xor UO_1596 (O_1596,N_10572,N_11855);
or UO_1597 (O_1597,N_11382,N_14407);
and UO_1598 (O_1598,N_13994,N_11677);
xor UO_1599 (O_1599,N_10565,N_14180);
nand UO_1600 (O_1600,N_12225,N_14122);
xnor UO_1601 (O_1601,N_12708,N_12616);
or UO_1602 (O_1602,N_10569,N_11412);
xnor UO_1603 (O_1603,N_12567,N_12862);
nor UO_1604 (O_1604,N_13593,N_14766);
or UO_1605 (O_1605,N_14345,N_13052);
nand UO_1606 (O_1606,N_14993,N_14841);
nand UO_1607 (O_1607,N_11964,N_11522);
and UO_1608 (O_1608,N_12044,N_14280);
nand UO_1609 (O_1609,N_14295,N_10148);
xor UO_1610 (O_1610,N_14360,N_12895);
nand UO_1611 (O_1611,N_12101,N_11426);
or UO_1612 (O_1612,N_10123,N_13976);
nor UO_1613 (O_1613,N_14542,N_13666);
nand UO_1614 (O_1614,N_14972,N_14520);
xnor UO_1615 (O_1615,N_10956,N_10027);
xor UO_1616 (O_1616,N_14434,N_14800);
xor UO_1617 (O_1617,N_12210,N_12845);
nand UO_1618 (O_1618,N_11320,N_14143);
or UO_1619 (O_1619,N_10233,N_10913);
xor UO_1620 (O_1620,N_11564,N_11380);
or UO_1621 (O_1621,N_11101,N_11264);
and UO_1622 (O_1622,N_14748,N_10253);
or UO_1623 (O_1623,N_13925,N_12140);
nor UO_1624 (O_1624,N_13720,N_13868);
and UO_1625 (O_1625,N_11475,N_14048);
xor UO_1626 (O_1626,N_11925,N_11759);
nand UO_1627 (O_1627,N_12252,N_11562);
and UO_1628 (O_1628,N_11226,N_10540);
nand UO_1629 (O_1629,N_11290,N_14729);
or UO_1630 (O_1630,N_11306,N_14352);
nand UO_1631 (O_1631,N_13025,N_11062);
or UO_1632 (O_1632,N_10392,N_12721);
xor UO_1633 (O_1633,N_11922,N_14545);
and UO_1634 (O_1634,N_12823,N_11003);
nor UO_1635 (O_1635,N_13319,N_11687);
xnor UO_1636 (O_1636,N_13181,N_14072);
or UO_1637 (O_1637,N_14020,N_11007);
or UO_1638 (O_1638,N_13259,N_14001);
nand UO_1639 (O_1639,N_12977,N_11929);
or UO_1640 (O_1640,N_12174,N_12995);
xor UO_1641 (O_1641,N_13443,N_10856);
or UO_1642 (O_1642,N_11170,N_11112);
xor UO_1643 (O_1643,N_14327,N_13028);
nand UO_1644 (O_1644,N_10481,N_12204);
nand UO_1645 (O_1645,N_13930,N_11519);
nand UO_1646 (O_1646,N_10722,N_10749);
and UO_1647 (O_1647,N_12974,N_11080);
nand UO_1648 (O_1648,N_12291,N_13276);
nor UO_1649 (O_1649,N_12051,N_12149);
or UO_1650 (O_1650,N_10387,N_14910);
nand UO_1651 (O_1651,N_11291,N_13662);
or UO_1652 (O_1652,N_10004,N_12158);
nor UO_1653 (O_1653,N_14955,N_14292);
xor UO_1654 (O_1654,N_10934,N_13937);
nand UO_1655 (O_1655,N_11909,N_14029);
xor UO_1656 (O_1656,N_13867,N_12746);
and UO_1657 (O_1657,N_14798,N_14156);
nand UO_1658 (O_1658,N_13106,N_14879);
xnor UO_1659 (O_1659,N_12682,N_13105);
and UO_1660 (O_1660,N_12631,N_13142);
nor UO_1661 (O_1661,N_12768,N_11670);
nand UO_1662 (O_1662,N_12414,N_13117);
nor UO_1663 (O_1663,N_13601,N_11325);
or UO_1664 (O_1664,N_14050,N_10974);
xnor UO_1665 (O_1665,N_11782,N_12391);
or UO_1666 (O_1666,N_14059,N_13977);
nand UO_1667 (O_1667,N_10656,N_12880);
or UO_1668 (O_1668,N_12572,N_10441);
xor UO_1669 (O_1669,N_14152,N_14438);
and UO_1670 (O_1670,N_12326,N_12527);
nor UO_1671 (O_1671,N_11763,N_14574);
and UO_1672 (O_1672,N_11554,N_10624);
and UO_1673 (O_1673,N_14915,N_10936);
xnor UO_1674 (O_1674,N_13775,N_11292);
or UO_1675 (O_1675,N_12622,N_14730);
and UO_1676 (O_1676,N_14648,N_11821);
nand UO_1677 (O_1677,N_14140,N_14837);
or UO_1678 (O_1678,N_11548,N_11351);
xor UO_1679 (O_1679,N_10018,N_11219);
or UO_1680 (O_1680,N_11249,N_14361);
xor UO_1681 (O_1681,N_11783,N_12482);
and UO_1682 (O_1682,N_12133,N_10409);
or UO_1683 (O_1683,N_10005,N_13170);
xnor UO_1684 (O_1684,N_11184,N_10401);
xnor UO_1685 (O_1685,N_11653,N_11151);
xor UO_1686 (O_1686,N_14247,N_13139);
nand UO_1687 (O_1687,N_14497,N_13112);
nand UO_1688 (O_1688,N_12676,N_14591);
nor UO_1689 (O_1689,N_14592,N_12715);
xor UO_1690 (O_1690,N_14357,N_10745);
or UO_1691 (O_1691,N_11790,N_13633);
xor UO_1692 (O_1692,N_11913,N_12617);
xor UO_1693 (O_1693,N_12111,N_10560);
xnor UO_1694 (O_1694,N_10669,N_13866);
nor UO_1695 (O_1695,N_10892,N_13488);
and UO_1696 (O_1696,N_14608,N_10196);
xor UO_1697 (O_1697,N_11434,N_12790);
xnor UO_1698 (O_1698,N_13716,N_10265);
xor UO_1699 (O_1699,N_13330,N_11240);
xor UO_1700 (O_1700,N_10811,N_14106);
nand UO_1701 (O_1701,N_10941,N_10555);
nor UO_1702 (O_1702,N_11546,N_11942);
or UO_1703 (O_1703,N_12742,N_12058);
and UO_1704 (O_1704,N_11472,N_11898);
or UO_1705 (O_1705,N_11354,N_12848);
nand UO_1706 (O_1706,N_11926,N_13575);
xnor UO_1707 (O_1707,N_10349,N_10767);
or UO_1708 (O_1708,N_13645,N_13555);
xor UO_1709 (O_1709,N_11093,N_10788);
nor UO_1710 (O_1710,N_14214,N_10924);
and UO_1711 (O_1711,N_13064,N_12411);
xnor UO_1712 (O_1712,N_13313,N_11698);
xnor UO_1713 (O_1713,N_14546,N_12801);
and UO_1714 (O_1714,N_14500,N_11049);
and UO_1715 (O_1715,N_12734,N_14531);
nand UO_1716 (O_1716,N_14054,N_14632);
xnor UO_1717 (O_1717,N_14790,N_13729);
and UO_1718 (O_1718,N_12187,N_12876);
xor UO_1719 (O_1719,N_12571,N_14797);
xnor UO_1720 (O_1720,N_13402,N_11339);
xnor UO_1721 (O_1721,N_10604,N_13648);
and UO_1722 (O_1722,N_13754,N_13906);
or UO_1723 (O_1723,N_14439,N_10728);
xnor UO_1724 (O_1724,N_12798,N_12156);
nand UO_1725 (O_1725,N_14457,N_11422);
nand UO_1726 (O_1726,N_13080,N_11707);
nand UO_1727 (O_1727,N_10012,N_12298);
or UO_1728 (O_1728,N_14146,N_12632);
or UO_1729 (O_1729,N_11341,N_10224);
xnor UO_1730 (O_1730,N_12711,N_10192);
or UO_1731 (O_1731,N_14508,N_11900);
nor UO_1732 (O_1732,N_12262,N_14676);
and UO_1733 (O_1733,N_11317,N_13782);
or UO_1734 (O_1734,N_14829,N_13573);
and UO_1735 (O_1735,N_14003,N_14119);
nand UO_1736 (O_1736,N_14141,N_11973);
xnor UO_1737 (O_1737,N_11490,N_14685);
xor UO_1738 (O_1738,N_14022,N_10919);
and UO_1739 (O_1739,N_14258,N_13116);
xor UO_1740 (O_1740,N_11874,N_14265);
xnor UO_1741 (O_1741,N_10128,N_12538);
nand UO_1742 (O_1742,N_14597,N_11733);
nor UO_1743 (O_1743,N_11983,N_14446);
xnor UO_1744 (O_1744,N_10456,N_12300);
xor UO_1745 (O_1745,N_11651,N_13195);
xor UO_1746 (O_1746,N_14626,N_10129);
nor UO_1747 (O_1747,N_11178,N_12424);
and UO_1748 (O_1748,N_10664,N_11066);
and UO_1749 (O_1749,N_10756,N_11799);
or UO_1750 (O_1750,N_11263,N_13485);
xor UO_1751 (O_1751,N_10770,N_12786);
xnor UO_1752 (O_1752,N_10246,N_10395);
nand UO_1753 (O_1753,N_13343,N_11082);
nor UO_1754 (O_1754,N_10024,N_14218);
nor UO_1755 (O_1755,N_14646,N_10643);
nor UO_1756 (O_1756,N_12337,N_12639);
xor UO_1757 (O_1757,N_10165,N_14844);
or UO_1758 (O_1758,N_11701,N_10695);
nor UO_1759 (O_1759,N_13568,N_13094);
nand UO_1760 (O_1760,N_14973,N_14049);
xor UO_1761 (O_1761,N_12153,N_14163);
nor UO_1762 (O_1762,N_13499,N_14563);
nand UO_1763 (O_1763,N_12497,N_13583);
or UO_1764 (O_1764,N_14429,N_11946);
or UO_1765 (O_1765,N_10783,N_13338);
xnor UO_1766 (O_1766,N_11685,N_13996);
nand UO_1767 (O_1767,N_14963,N_14196);
nand UO_1768 (O_1768,N_12934,N_13654);
or UO_1769 (O_1769,N_10199,N_14132);
nand UO_1770 (O_1770,N_10631,N_13470);
and UO_1771 (O_1771,N_12086,N_11645);
nor UO_1772 (O_1772,N_13325,N_10909);
nor UO_1773 (O_1773,N_13822,N_13834);
or UO_1774 (O_1774,N_12751,N_14750);
nand UO_1775 (O_1775,N_12812,N_14988);
nand UO_1776 (O_1776,N_10689,N_13093);
or UO_1777 (O_1777,N_12852,N_12940);
nor UO_1778 (O_1778,N_14781,N_12673);
nand UO_1779 (O_1779,N_10207,N_14070);
and UO_1780 (O_1780,N_12419,N_13339);
and UO_1781 (O_1781,N_10189,N_12362);
nor UO_1782 (O_1782,N_10332,N_10771);
nand UO_1783 (O_1783,N_14123,N_12143);
and UO_1784 (O_1784,N_10691,N_13377);
xnor UO_1785 (O_1785,N_12319,N_14061);
or UO_1786 (O_1786,N_14368,N_12670);
and UO_1787 (O_1787,N_13372,N_13379);
and UO_1788 (O_1788,N_12781,N_10910);
nor UO_1789 (O_1789,N_12347,N_10383);
nor UO_1790 (O_1790,N_13761,N_11300);
nand UO_1791 (O_1791,N_12847,N_10798);
or UO_1792 (O_1792,N_12039,N_14742);
nand UO_1793 (O_1793,N_12152,N_11742);
nor UO_1794 (O_1794,N_12536,N_14706);
nand UO_1795 (O_1795,N_12693,N_12368);
nor UO_1796 (O_1796,N_11109,N_12448);
or UO_1797 (O_1797,N_11518,N_11755);
xor UO_1798 (O_1798,N_13137,N_14362);
nor UO_1799 (O_1799,N_10471,N_13244);
nand UO_1800 (O_1800,N_11462,N_11154);
and UO_1801 (O_1801,N_13740,N_11863);
xnor UO_1802 (O_1802,N_14064,N_11348);
and UO_1803 (O_1803,N_13034,N_11100);
nand UO_1804 (O_1804,N_13410,N_12717);
nand UO_1805 (O_1805,N_11791,N_12566);
nand UO_1806 (O_1806,N_11310,N_10286);
and UO_1807 (O_1807,N_10010,N_13570);
xnor UO_1808 (O_1808,N_10854,N_14330);
and UO_1809 (O_1809,N_11549,N_11680);
nor UO_1810 (O_1810,N_13376,N_10322);
xnor UO_1811 (O_1811,N_10179,N_10763);
and UO_1812 (O_1812,N_12028,N_14860);
and UO_1813 (O_1813,N_11060,N_12214);
nand UO_1814 (O_1814,N_14782,N_11138);
or UO_1815 (O_1815,N_10567,N_10766);
xor UO_1816 (O_1816,N_10670,N_14524);
nand UO_1817 (O_1817,N_11425,N_14785);
or UO_1818 (O_1818,N_12358,N_12343);
nor UO_1819 (O_1819,N_11414,N_11087);
nor UO_1820 (O_1820,N_14272,N_13821);
xnor UO_1821 (O_1821,N_13886,N_11089);
xnor UO_1822 (O_1822,N_13674,N_12455);
and UO_1823 (O_1823,N_11126,N_14899);
nand UO_1824 (O_1824,N_10570,N_10903);
or UO_1825 (O_1825,N_14039,N_13301);
or UO_1826 (O_1826,N_14598,N_11754);
nand UO_1827 (O_1827,N_13594,N_12378);
nand UO_1828 (O_1828,N_10534,N_11455);
xor UO_1829 (O_1829,N_10918,N_14073);
nor UO_1830 (O_1830,N_11352,N_11449);
nor UO_1831 (O_1831,N_11055,N_12666);
nand UO_1832 (O_1832,N_12795,N_10335);
nand UO_1833 (O_1833,N_13378,N_14682);
nor UO_1834 (O_1834,N_13794,N_10630);
xor UO_1835 (O_1835,N_14147,N_14977);
xnor UO_1836 (O_1836,N_11203,N_11438);
or UO_1837 (O_1837,N_11847,N_12311);
or UO_1838 (O_1838,N_12558,N_14891);
or UO_1839 (O_1839,N_11042,N_11296);
and UO_1840 (O_1840,N_11699,N_10289);
nor UO_1841 (O_1841,N_11227,N_12275);
and UO_1842 (O_1842,N_12568,N_12090);
xor UO_1843 (O_1843,N_10333,N_13299);
nand UO_1844 (O_1844,N_12896,N_10097);
or UO_1845 (O_1845,N_11640,N_13213);
or UO_1846 (O_1846,N_13600,N_13005);
and UO_1847 (O_1847,N_10989,N_13321);
nand UO_1848 (O_1848,N_13020,N_10736);
nand UO_1849 (O_1849,N_10646,N_13898);
or UO_1850 (O_1850,N_14604,N_13912);
xnor UO_1851 (O_1851,N_12811,N_12150);
xor UO_1852 (O_1852,N_12313,N_14223);
nor UO_1853 (O_1853,N_14337,N_12392);
nand UO_1854 (O_1854,N_12577,N_14101);
and UO_1855 (O_1855,N_12163,N_11977);
and UO_1856 (O_1856,N_12562,N_12301);
and UO_1857 (O_1857,N_13698,N_12839);
and UO_1858 (O_1858,N_11528,N_11079);
or UO_1859 (O_1859,N_12200,N_12894);
and UO_1860 (O_1860,N_10773,N_11884);
and UO_1861 (O_1861,N_11849,N_13664);
xnor UO_1862 (O_1862,N_14547,N_10973);
and UO_1863 (O_1863,N_10221,N_14527);
xor UO_1864 (O_1864,N_12983,N_14741);
nand UO_1865 (O_1865,N_10657,N_14658);
or UO_1866 (O_1866,N_11364,N_13515);
xor UO_1867 (O_1867,N_14739,N_12509);
xor UO_1868 (O_1868,N_11181,N_13085);
xor UO_1869 (O_1869,N_14712,N_11510);
xnor UO_1870 (O_1870,N_14843,N_12818);
nor UO_1871 (O_1871,N_14144,N_10068);
xor UO_1872 (O_1872,N_13743,N_13920);
nor UO_1873 (O_1873,N_12667,N_13544);
nand UO_1874 (O_1874,N_14707,N_12393);
nand UO_1875 (O_1875,N_14491,N_12441);
xnor UO_1876 (O_1876,N_11498,N_14927);
and UO_1877 (O_1877,N_13446,N_14566);
or UO_1878 (O_1878,N_12533,N_10731);
nor UO_1879 (O_1879,N_12539,N_12342);
and UO_1880 (O_1880,N_12733,N_10855);
nor UO_1881 (O_1881,N_10351,N_12047);
nand UO_1882 (O_1882,N_13979,N_11787);
xnor UO_1883 (O_1883,N_11444,N_12753);
xnor UO_1884 (O_1884,N_13357,N_10470);
and UO_1885 (O_1885,N_11161,N_14182);
and UO_1886 (O_1886,N_10713,N_14058);
nand UO_1887 (O_1887,N_12932,N_14753);
nand UO_1888 (O_1888,N_10290,N_13658);
or UO_1889 (O_1889,N_13365,N_12529);
nand UO_1890 (O_1890,N_12863,N_12032);
nand UO_1891 (O_1891,N_10512,N_14283);
nand UO_1892 (O_1892,N_13182,N_10678);
or UO_1893 (O_1893,N_10378,N_13688);
nand UO_1894 (O_1894,N_13345,N_10112);
xnor UO_1895 (O_1895,N_12230,N_14744);
nand UO_1896 (O_1896,N_11254,N_13130);
or UO_1897 (O_1897,N_13660,N_11868);
or UO_1898 (O_1898,N_11396,N_12069);
xor UO_1899 (O_1899,N_12198,N_10829);
nor UO_1900 (O_1900,N_10981,N_11842);
nand UO_1901 (O_1901,N_13692,N_11432);
nor UO_1902 (O_1902,N_14302,N_14571);
and UO_1903 (O_1903,N_10261,N_10760);
and UO_1904 (O_1904,N_13411,N_14287);
nand UO_1905 (O_1905,N_14962,N_12139);
nor UO_1906 (O_1906,N_10720,N_13063);
nor UO_1907 (O_1907,N_10330,N_11421);
or UO_1908 (O_1908,N_14353,N_10601);
nand UO_1909 (O_1909,N_13168,N_14672);
and UO_1910 (O_1910,N_12205,N_13396);
nor UO_1911 (O_1911,N_11243,N_13021);
xnor UO_1912 (O_1912,N_14068,N_13211);
xor UO_1913 (O_1913,N_14496,N_12000);
xnor UO_1914 (O_1914,N_13719,N_10994);
xnor UO_1915 (O_1915,N_12816,N_14379);
nor UO_1916 (O_1916,N_13657,N_11535);
xnor UO_1917 (O_1917,N_11132,N_10759);
nor UO_1918 (O_1918,N_14888,N_12213);
xor UO_1919 (O_1919,N_12651,N_14165);
and UO_1920 (O_1920,N_14703,N_12194);
nor UO_1921 (O_1921,N_13627,N_10467);
nor UO_1922 (O_1922,N_13353,N_11211);
nor UO_1923 (O_1923,N_10413,N_14421);
and UO_1924 (O_1924,N_11308,N_12523);
nor UO_1925 (O_1925,N_14687,N_13663);
xnor UO_1926 (O_1926,N_11391,N_13250);
or UO_1927 (O_1927,N_14153,N_12764);
nor UO_1928 (O_1928,N_12855,N_12657);
or UO_1929 (O_1929,N_11800,N_10575);
xnor UO_1930 (O_1930,N_11831,N_12215);
nand UO_1931 (O_1931,N_14652,N_10238);
xor UO_1932 (O_1932,N_11435,N_11046);
or UO_1933 (O_1933,N_11837,N_11693);
or UO_1934 (O_1934,N_14274,N_12610);
xor UO_1935 (O_1935,N_14226,N_10143);
nand UO_1936 (O_1936,N_14883,N_10834);
xor UO_1937 (O_1937,N_14557,N_10594);
nor UO_1938 (O_1938,N_14030,N_12350);
nand UO_1939 (O_1939,N_13334,N_10754);
xnor UO_1940 (O_1940,N_10247,N_13738);
nand UO_1941 (O_1941,N_11503,N_13405);
or UO_1942 (O_1942,N_12906,N_14419);
nand UO_1943 (O_1943,N_12591,N_14256);
xor UO_1944 (O_1944,N_12996,N_10992);
and UO_1945 (O_1945,N_12856,N_12325);
or UO_1946 (O_1946,N_11563,N_11745);
nand UO_1947 (O_1947,N_11437,N_14928);
and UO_1948 (O_1948,N_13163,N_11294);
nand UO_1949 (O_1949,N_13352,N_12449);
and UO_1950 (O_1950,N_12589,N_12967);
nand UO_1951 (O_1951,N_10180,N_13818);
nand UO_1952 (O_1952,N_13156,N_12287);
and UO_1953 (O_1953,N_13091,N_14403);
nand UO_1954 (O_1954,N_12501,N_12763);
nor UO_1955 (O_1955,N_11431,N_11450);
nand UO_1956 (O_1956,N_11143,N_11282);
and UO_1957 (O_1957,N_12645,N_10578);
and UO_1958 (O_1958,N_13266,N_11251);
xor UO_1959 (O_1959,N_12752,N_10135);
or UO_1960 (O_1960,N_11696,N_10561);
xor UO_1961 (O_1961,N_14552,N_13913);
xor UO_1962 (O_1962,N_13733,N_14997);
or UO_1963 (O_1963,N_14824,N_10047);
or UO_1964 (O_1964,N_12131,N_13841);
or UO_1965 (O_1965,N_11220,N_10535);
and UO_1966 (O_1966,N_12943,N_11943);
or UO_1967 (O_1967,N_13521,N_13238);
nand UO_1968 (O_1968,N_14992,N_14253);
nand UO_1969 (O_1969,N_13125,N_13828);
or UO_1970 (O_1970,N_10249,N_14002);
xnor UO_1971 (O_1971,N_11200,N_11697);
and UO_1972 (O_1972,N_13088,N_10414);
or UO_1973 (O_1973,N_12952,N_11474);
nand UO_1974 (O_1974,N_11429,N_11771);
and UO_1975 (O_1975,N_11149,N_12807);
and UO_1976 (O_1976,N_10302,N_10533);
xor UO_1977 (O_1977,N_14097,N_14689);
nand UO_1978 (O_1978,N_11250,N_13278);
and UO_1979 (O_1979,N_10280,N_13358);
and UO_1980 (O_1980,N_13441,N_11193);
or UO_1981 (O_1981,N_11904,N_14631);
nor UO_1982 (O_1982,N_10009,N_12599);
nand UO_1983 (O_1983,N_12844,N_10977);
nand UO_1984 (O_1984,N_13109,N_11466);
or UO_1985 (O_1985,N_12048,N_12125);
xor UO_1986 (O_1986,N_12109,N_12084);
nor UO_1987 (O_1987,N_10473,N_12913);
nor UO_1988 (O_1988,N_13102,N_12190);
xnor UO_1989 (O_1989,N_11899,N_14717);
and UO_1990 (O_1990,N_12680,N_14260);
or UO_1991 (O_1991,N_13523,N_10462);
or UO_1992 (O_1992,N_10607,N_14804);
and UO_1993 (O_1993,N_14300,N_11674);
xor UO_1994 (O_1994,N_12808,N_14622);
or UO_1995 (O_1995,N_14836,N_10430);
nand UO_1996 (O_1996,N_13851,N_11917);
nand UO_1997 (O_1997,N_10951,N_11123);
nand UO_1998 (O_1998,N_12675,N_12066);
nor UO_1999 (O_1999,N_11387,N_13629);
endmodule